module basic_1500_15000_2000_30_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_599,In_474);
xnor U1 (N_1,In_763,In_989);
nand U2 (N_2,In_929,In_809);
nand U3 (N_3,In_852,In_1055);
and U4 (N_4,In_456,In_1370);
xor U5 (N_5,In_412,In_1149);
and U6 (N_6,In_125,In_996);
nand U7 (N_7,In_638,In_111);
nand U8 (N_8,In_19,In_369);
or U9 (N_9,In_1223,In_1034);
nor U10 (N_10,In_1315,In_644);
nand U11 (N_11,In_202,In_287);
or U12 (N_12,In_484,In_908);
or U13 (N_13,In_281,In_52);
nand U14 (N_14,In_356,In_392);
xnor U15 (N_15,In_469,In_1440);
and U16 (N_16,In_967,In_733);
and U17 (N_17,In_548,In_846);
nor U18 (N_18,In_1265,In_537);
nor U19 (N_19,In_709,In_740);
and U20 (N_20,In_1270,In_1291);
xor U21 (N_21,In_1139,In_1129);
or U22 (N_22,In_396,In_1012);
and U23 (N_23,In_350,In_1080);
nand U24 (N_24,In_1249,In_785);
or U25 (N_25,In_152,In_1145);
and U26 (N_26,In_687,In_206);
or U27 (N_27,In_587,In_21);
or U28 (N_28,In_397,In_61);
xor U29 (N_29,In_1007,In_312);
nand U30 (N_30,In_895,In_909);
and U31 (N_31,In_930,In_843);
or U32 (N_32,In_209,In_535);
nand U33 (N_33,In_406,In_1352);
or U34 (N_34,In_945,In_1339);
nor U35 (N_35,In_1182,In_1446);
nand U36 (N_36,In_1138,In_1222);
nand U37 (N_37,In_76,In_1146);
and U38 (N_38,In_651,In_1165);
xnor U39 (N_39,In_906,In_575);
nor U40 (N_40,In_1389,In_1369);
nor U41 (N_41,In_1183,In_303);
or U42 (N_42,In_153,In_58);
nor U43 (N_43,In_1455,In_541);
and U44 (N_44,In_1075,In_1428);
xor U45 (N_45,In_1140,In_1022);
nand U46 (N_46,In_1303,In_1341);
or U47 (N_47,In_617,In_758);
or U48 (N_48,In_619,In_689);
or U49 (N_49,In_1326,In_1448);
and U50 (N_50,In_1136,In_1130);
or U51 (N_51,In_433,In_1027);
nor U52 (N_52,In_694,In_232);
xor U53 (N_53,In_864,In_316);
or U54 (N_54,In_530,In_378);
and U55 (N_55,In_635,In_566);
nor U56 (N_56,In_1392,In_308);
and U57 (N_57,In_868,In_804);
and U58 (N_58,In_1162,In_216);
or U59 (N_59,In_571,In_1091);
nor U60 (N_60,In_1131,In_509);
and U61 (N_61,In_821,In_1191);
and U62 (N_62,In_108,In_734);
and U63 (N_63,In_950,In_1148);
xnor U64 (N_64,In_1294,In_340);
nor U65 (N_65,In_873,In_245);
or U66 (N_66,In_521,In_1260);
nand U67 (N_67,In_1120,In_1090);
nand U68 (N_68,In_172,In_444);
xor U69 (N_69,In_164,In_1436);
and U70 (N_70,In_30,In_157);
and U71 (N_71,In_1362,In_1167);
or U72 (N_72,In_973,In_1304);
or U73 (N_73,In_855,In_600);
xnor U74 (N_74,In_344,In_1051);
and U75 (N_75,In_991,In_170);
or U76 (N_76,In_494,In_649);
nor U77 (N_77,In_815,In_28);
and U78 (N_78,In_552,In_1092);
or U79 (N_79,In_1403,In_1214);
and U80 (N_80,In_149,In_346);
nand U81 (N_81,In_425,In_724);
and U82 (N_82,In_1036,In_681);
and U83 (N_83,In_1283,In_1279);
or U84 (N_84,In_1324,In_673);
and U85 (N_85,In_15,In_215);
or U86 (N_86,In_191,In_1445);
nand U87 (N_87,In_1,In_313);
nand U88 (N_88,In_1390,In_579);
and U89 (N_89,In_1166,In_1156);
or U90 (N_90,In_761,In_831);
nand U91 (N_91,In_1499,In_289);
or U92 (N_92,In_1126,In_292);
or U93 (N_93,In_519,In_661);
xnor U94 (N_94,In_1382,In_1266);
or U95 (N_95,In_1234,In_1246);
and U96 (N_96,In_1132,In_6);
and U97 (N_97,In_1329,In_558);
xor U98 (N_98,In_175,In_326);
or U99 (N_99,In_163,In_631);
or U100 (N_100,In_1072,In_252);
nand U101 (N_101,In_64,In_1104);
nand U102 (N_102,In_293,In_940);
nor U103 (N_103,In_63,In_1231);
or U104 (N_104,In_105,In_1463);
nor U105 (N_105,In_89,In_595);
and U106 (N_106,In_630,In_1196);
nor U107 (N_107,In_976,In_739);
nor U108 (N_108,In_876,In_24);
or U109 (N_109,In_858,In_620);
nor U110 (N_110,In_35,In_961);
or U111 (N_111,In_539,In_389);
nand U112 (N_112,In_4,In_307);
and U113 (N_113,In_860,In_1275);
nor U114 (N_114,In_495,In_472);
nand U115 (N_115,In_233,In_1185);
or U116 (N_116,In_86,In_243);
xnor U117 (N_117,In_789,In_1255);
nor U118 (N_118,In_725,In_1037);
nand U119 (N_119,In_1331,In_602);
nand U120 (N_120,In_394,In_314);
nor U121 (N_121,In_590,In_1401);
nand U122 (N_122,In_641,In_576);
and U123 (N_123,In_1468,In_1006);
nor U124 (N_124,In_330,In_1084);
xor U125 (N_125,In_748,In_241);
or U126 (N_126,In_1487,In_880);
and U127 (N_127,In_791,In_1349);
nand U128 (N_128,In_1060,In_1374);
or U129 (N_129,In_918,In_1056);
nor U130 (N_130,In_388,In_606);
and U131 (N_131,In_914,In_975);
xor U132 (N_132,In_403,In_1114);
or U133 (N_133,In_555,In_547);
xnor U134 (N_134,In_672,In_165);
nand U135 (N_135,In_1258,In_954);
xnor U136 (N_136,In_557,In_705);
nand U137 (N_137,In_324,In_712);
xor U138 (N_138,In_656,In_290);
xnor U139 (N_139,In_1491,In_790);
nor U140 (N_140,In_1224,In_1202);
or U141 (N_141,In_743,In_449);
nand U142 (N_142,In_193,In_467);
xnor U143 (N_143,In_1267,In_1178);
and U144 (N_144,In_995,In_99);
xor U145 (N_145,In_890,In_1411);
nor U146 (N_146,In_792,In_483);
or U147 (N_147,In_1289,In_120);
nor U148 (N_148,In_1048,In_311);
and U149 (N_149,In_62,In_753);
and U150 (N_150,In_1099,In_933);
nand U151 (N_151,In_1274,In_910);
nor U152 (N_152,In_1313,In_1361);
nor U153 (N_153,In_1328,In_1016);
or U154 (N_154,In_488,In_382);
and U155 (N_155,In_702,In_710);
xnor U156 (N_156,In_1338,In_677);
or U157 (N_157,In_1251,In_794);
and U158 (N_158,In_911,In_26);
xor U159 (N_159,In_1197,In_1233);
nand U160 (N_160,In_113,In_124);
nand U161 (N_161,In_531,In_826);
or U162 (N_162,In_1187,In_140);
and U163 (N_163,In_865,In_65);
nand U164 (N_164,In_944,In_177);
or U165 (N_165,In_1128,In_1204);
nand U166 (N_166,In_1229,In_889);
and U167 (N_167,In_1282,In_1256);
or U168 (N_168,In_559,In_1212);
and U169 (N_169,In_112,In_1285);
xnor U170 (N_170,In_808,In_497);
xnor U171 (N_171,In_342,In_167);
nor U172 (N_172,In_665,In_185);
nand U173 (N_173,In_300,In_942);
or U174 (N_174,In_212,In_1317);
nor U175 (N_175,In_435,In_625);
xor U176 (N_176,In_383,In_956);
nand U177 (N_177,In_1239,In_1356);
nand U178 (N_178,In_331,In_1348);
or U179 (N_179,In_1035,In_1447);
and U180 (N_180,In_985,In_1474);
nor U181 (N_181,In_1142,In_742);
xor U182 (N_182,In_471,In_1453);
or U183 (N_183,In_390,In_82);
xnor U184 (N_184,In_1412,In_834);
nor U185 (N_185,In_91,In_1081);
nand U186 (N_186,In_772,In_87);
xnor U187 (N_187,In_1059,In_273);
and U188 (N_188,In_588,In_723);
xor U189 (N_189,In_399,In_1386);
nand U190 (N_190,In_1449,In_227);
nor U191 (N_191,In_250,In_714);
xor U192 (N_192,In_154,In_1323);
and U193 (N_193,In_1077,In_1300);
or U194 (N_194,In_887,In_376);
xnor U195 (N_195,In_1434,In_881);
and U196 (N_196,In_80,In_518);
nor U197 (N_197,In_1498,In_1330);
xnor U198 (N_198,In_1003,In_1497);
or U199 (N_199,In_213,In_74);
nor U200 (N_200,In_904,In_682);
nor U201 (N_201,In_1032,In_827);
xnor U202 (N_202,In_793,In_589);
xnor U203 (N_203,In_420,In_242);
xnor U204 (N_204,In_731,In_829);
xnor U205 (N_205,In_1040,In_132);
and U206 (N_206,In_458,In_1351);
and U207 (N_207,In_231,In_732);
nor U208 (N_208,In_1306,In_755);
nor U209 (N_209,In_837,In_1103);
nor U210 (N_210,In_1029,In_593);
nor U211 (N_211,In_1068,In_1444);
and U212 (N_212,In_1124,In_13);
or U213 (N_213,In_862,In_953);
and U214 (N_214,In_863,In_756);
or U215 (N_215,In_156,In_807);
xnor U216 (N_216,In_990,In_1049);
or U217 (N_217,In_114,In_1305);
and U218 (N_218,In_849,In_1226);
or U219 (N_219,In_278,In_782);
or U220 (N_220,In_424,In_452);
and U221 (N_221,In_1159,In_454);
xnor U222 (N_222,In_468,In_47);
nor U223 (N_223,In_173,In_370);
or U224 (N_224,In_722,In_1297);
or U225 (N_225,In_421,In_643);
and U226 (N_226,In_141,In_769);
or U227 (N_227,In_234,In_817);
xnor U228 (N_228,In_1050,In_1442);
and U229 (N_229,In_490,In_774);
nor U230 (N_230,In_607,In_393);
nor U231 (N_231,In_1121,In_11);
xnor U232 (N_232,In_1171,In_1096);
nor U233 (N_233,In_984,In_741);
xor U234 (N_234,In_249,In_1460);
or U235 (N_235,In_476,In_901);
nor U236 (N_236,In_151,In_43);
nand U237 (N_237,In_240,In_966);
xor U238 (N_238,In_253,In_1462);
nand U239 (N_239,In_1264,In_417);
xor U240 (N_240,In_200,In_1347);
or U241 (N_241,In_1409,In_1364);
nor U242 (N_242,In_1360,In_103);
xor U243 (N_243,In_459,In_1335);
or U244 (N_244,In_1344,In_338);
nor U245 (N_245,In_968,In_1465);
and U246 (N_246,In_894,In_219);
or U247 (N_247,In_912,In_1158);
or U248 (N_248,In_230,In_1414);
xnor U249 (N_249,In_500,In_1383);
and U250 (N_250,In_727,In_542);
nand U251 (N_251,In_546,In_135);
nor U252 (N_252,In_1109,In_288);
nand U253 (N_253,In_1367,In_1484);
and U254 (N_254,In_926,In_504);
xor U255 (N_255,In_441,In_1154);
nand U256 (N_256,In_134,In_72);
or U257 (N_257,In_1493,In_25);
and U258 (N_258,In_286,In_264);
xor U259 (N_259,In_1039,In_123);
nand U260 (N_260,In_309,In_982);
nor U261 (N_261,In_998,In_1477);
and U262 (N_262,In_1253,In_371);
and U263 (N_263,In_1230,In_419);
xor U264 (N_264,In_1295,In_1024);
nand U265 (N_265,In_128,In_413);
nand U266 (N_266,In_646,In_1451);
and U267 (N_267,In_691,In_964);
xor U268 (N_268,In_892,In_1026);
or U269 (N_269,In_489,In_357);
nand U270 (N_270,In_96,In_1107);
nand U271 (N_271,In_29,In_698);
nand U272 (N_272,In_1086,In_1398);
or U273 (N_273,In_1481,In_60);
and U274 (N_274,In_1227,In_1490);
and U275 (N_275,In_980,In_1061);
xnor U276 (N_276,In_1378,In_612);
nand U277 (N_277,In_695,In_1118);
or U278 (N_278,In_1280,In_1483);
and U279 (N_279,In_1371,In_629);
xnor U280 (N_280,In_805,In_594);
nor U281 (N_281,In_439,In_260);
and U282 (N_282,In_1046,In_121);
xor U283 (N_283,In_553,In_1473);
nor U284 (N_284,In_986,In_1175);
nor U285 (N_285,In_679,In_1495);
nand U286 (N_286,In_196,In_1134);
nor U287 (N_287,In_318,In_5);
xor U288 (N_288,In_328,In_948);
xnor U289 (N_289,In_655,In_1186);
xnor U290 (N_290,In_18,In_1209);
and U291 (N_291,In_190,In_499);
xnor U292 (N_292,In_1421,In_401);
and U293 (N_293,In_538,In_22);
nor U294 (N_294,In_582,In_122);
or U295 (N_295,In_783,In_615);
and U296 (N_296,In_1342,In_1419);
xnor U297 (N_297,In_487,In_845);
and U298 (N_298,In_1441,In_126);
and U299 (N_299,In_432,In_470);
xor U300 (N_300,In_1021,In_745);
or U301 (N_301,In_871,In_752);
nand U302 (N_302,In_398,In_343);
xor U303 (N_303,In_937,In_1064);
or U304 (N_304,In_1262,In_1277);
nand U305 (N_305,In_1108,In_147);
or U306 (N_306,In_1286,In_946);
nand U307 (N_307,In_1343,In_1248);
nand U308 (N_308,In_543,In_1438);
nand U309 (N_309,In_272,In_237);
xor U310 (N_310,In_1151,In_247);
xor U311 (N_311,In_94,In_465);
and U312 (N_312,In_1333,In_295);
and U313 (N_313,In_853,In_1170);
nand U314 (N_314,In_1492,In_701);
and U315 (N_315,In_68,In_222);
or U316 (N_316,In_983,In_1437);
xor U317 (N_317,In_71,In_992);
and U318 (N_318,In_762,In_426);
nand U319 (N_319,In_81,In_664);
xnor U320 (N_320,In_285,In_605);
nor U321 (N_321,In_201,In_818);
nor U322 (N_322,In_1079,In_296);
nand U323 (N_323,In_118,In_811);
xnor U324 (N_324,In_327,In_527);
nand U325 (N_325,In_1002,In_611);
or U326 (N_326,In_229,In_941);
nor U327 (N_327,In_508,In_1245);
nand U328 (N_328,In_115,In_776);
nor U329 (N_329,In_1115,In_1038);
nor U330 (N_330,In_276,In_1257);
nor U331 (N_331,In_1000,In_878);
nor U332 (N_332,In_56,In_997);
nand U333 (N_333,In_345,In_943);
nor U334 (N_334,In_585,In_886);
and U335 (N_335,In_628,In_438);
nor U336 (N_336,In_45,In_835);
nor U337 (N_337,In_757,In_1242);
nand U338 (N_338,In_1127,In_1357);
xnor U339 (N_339,In_766,In_728);
nand U340 (N_340,In_1416,In_1053);
nor U341 (N_341,In_102,In_1188);
or U342 (N_342,In_225,In_637);
nand U343 (N_343,In_1408,In_1346);
nand U344 (N_344,In_913,In_704);
xnor U345 (N_345,In_1388,In_1410);
nor U346 (N_346,In_246,In_720);
nand U347 (N_347,In_1232,In_529);
nand U348 (N_348,In_168,In_703);
nor U349 (N_349,In_564,In_1496);
nand U350 (N_350,In_1464,In_279);
or U351 (N_351,In_1396,In_280);
xnor U352 (N_352,In_528,In_1116);
nand U353 (N_353,In_1228,In_675);
nor U354 (N_354,In_738,In_491);
xnor U355 (N_355,In_298,In_699);
nand U356 (N_356,In_182,In_866);
xnor U357 (N_357,In_1469,In_988);
nor U358 (N_358,In_1017,In_604);
nor U359 (N_359,In_184,In_872);
and U360 (N_360,In_1311,In_197);
or U361 (N_361,In_806,In_372);
or U362 (N_362,In_78,In_37);
xor U363 (N_363,In_735,In_1194);
or U364 (N_364,In_999,In_1093);
nor U365 (N_365,In_1173,In_773);
nor U366 (N_366,In_457,In_522);
and U367 (N_367,In_51,In_1133);
or U368 (N_368,In_1045,In_798);
nand U369 (N_369,In_613,In_568);
xnor U370 (N_370,In_534,In_1161);
xor U371 (N_371,In_77,In_1152);
nor U372 (N_372,In_1377,In_884);
xnor U373 (N_373,In_799,In_493);
or U374 (N_374,In_647,In_31);
xnor U375 (N_375,In_315,In_377);
xor U376 (N_376,In_339,In_1095);
nor U377 (N_377,In_17,In_93);
and U378 (N_378,In_786,In_916);
or U379 (N_379,In_130,In_179);
nor U380 (N_380,In_532,In_797);
nor U381 (N_381,In_53,In_1100);
nand U382 (N_382,In_422,In_1206);
or U383 (N_383,In_931,In_442);
nor U384 (N_384,In_95,In_627);
or U385 (N_385,In_737,In_402);
nor U386 (N_386,In_648,In_1067);
or U387 (N_387,In_1458,In_387);
nor U388 (N_388,In_639,In_1433);
and U389 (N_389,In_959,In_416);
nand U390 (N_390,In_608,In_1314);
xor U391 (N_391,In_1236,In_696);
nand U392 (N_392,In_379,In_198);
xnor U393 (N_393,In_965,In_158);
or U394 (N_394,In_1259,In_780);
or U395 (N_395,In_501,In_634);
nor U396 (N_396,In_20,In_1254);
and U397 (N_397,In_429,In_255);
nand U398 (N_398,In_1088,In_847);
nor U399 (N_399,In_144,In_507);
and U400 (N_400,In_893,In_1147);
and U401 (N_401,In_1312,In_473);
nor U402 (N_402,In_978,In_1334);
nand U403 (N_403,In_10,In_92);
nor U404 (N_404,In_642,In_358);
nand U405 (N_405,In_1366,In_1405);
or U406 (N_406,In_1176,In_214);
or U407 (N_407,In_934,In_551);
or U408 (N_408,In_427,In_819);
xor U409 (N_409,In_258,In_917);
nand U410 (N_410,In_320,In_1423);
and U411 (N_411,In_957,In_1174);
nand U412 (N_412,In_657,In_1082);
xor U413 (N_413,In_877,In_1435);
and U414 (N_414,In_161,In_1117);
nand U415 (N_415,In_977,In_174);
and U416 (N_416,In_716,In_801);
or U417 (N_417,In_1425,In_869);
or U418 (N_418,In_1083,In_1023);
and U419 (N_419,In_692,In_668);
and U420 (N_420,In_771,In_1179);
nor U421 (N_421,In_485,In_261);
xor U422 (N_422,In_1047,In_256);
nor U423 (N_423,In_1296,In_1439);
and U424 (N_424,In_1135,In_970);
xnor U425 (N_425,In_359,In_455);
nand U426 (N_426,In_75,In_1387);
or U427 (N_427,In_479,In_1119);
nand U428 (N_428,In_3,In_795);
nor U429 (N_429,In_333,In_994);
nor U430 (N_430,In_1062,In_759);
and U431 (N_431,In_131,In_1244);
or U432 (N_432,In_351,In_554);
and U433 (N_433,In_1163,In_1144);
nor U434 (N_434,In_1391,In_217);
xnor U435 (N_435,In_409,In_1404);
nand U436 (N_436,In_428,In_1225);
and U437 (N_437,In_301,In_569);
nand U438 (N_438,In_833,In_1393);
xor U439 (N_439,In_584,In_574);
or U440 (N_440,In_875,In_1097);
or U441 (N_441,In_1177,In_573);
or U442 (N_442,In_840,In_836);
nor U443 (N_443,In_947,In_1052);
nor U444 (N_444,In_1033,In_561);
nor U445 (N_445,In_323,In_451);
nor U446 (N_446,In_1241,In_1293);
nor U447 (N_447,In_718,In_562);
nor U448 (N_448,In_971,In_563);
nor U449 (N_449,In_41,In_778);
or U450 (N_450,In_1071,In_1278);
or U451 (N_451,In_1431,In_1190);
nand U452 (N_452,In_100,In_1203);
nor U453 (N_453,In_1057,In_1384);
and U454 (N_454,In_110,In_129);
or U455 (N_455,In_73,In_768);
and U456 (N_456,In_16,In_431);
xnor U457 (N_457,In_317,In_700);
and U458 (N_458,In_659,In_171);
and U459 (N_459,In_1385,In_1089);
and U460 (N_460,In_199,In_1200);
nand U461 (N_461,In_736,In_70);
xnor U462 (N_462,In_1290,In_137);
nand U463 (N_463,In_730,In_14);
nor U464 (N_464,In_597,In_352);
or U465 (N_465,In_1168,In_1058);
nor U466 (N_466,In_787,In_400);
nor U467 (N_467,In_623,In_922);
and U468 (N_468,In_897,In_1213);
nor U469 (N_469,In_275,In_680);
nand U470 (N_470,In_502,In_1074);
xnor U471 (N_471,In_603,In_578);
nor U472 (N_472,In_962,In_79);
xnor U473 (N_473,In_1368,In_900);
nor U474 (N_474,In_48,In_824);
and U475 (N_475,In_751,In_192);
nor U476 (N_476,In_39,In_609);
nand U477 (N_477,In_662,In_1413);
nor U478 (N_478,In_903,In_706);
nand U479 (N_479,In_1426,In_1005);
xnor U480 (N_480,In_511,In_598);
and U481 (N_481,In_848,In_1210);
and U482 (N_482,In_437,In_1480);
nor U483 (N_483,In_1276,In_1044);
xor U484 (N_484,In_1112,In_373);
or U485 (N_485,In_879,In_586);
nand U486 (N_486,In_1430,In_1008);
xnor U487 (N_487,In_1308,In_44);
xnor U488 (N_488,In_1345,In_1054);
nor U489 (N_489,In_166,In_1143);
nor U490 (N_490,In_1063,In_674);
or U491 (N_491,In_244,In_1211);
nand U492 (N_492,In_33,In_1180);
xnor U493 (N_493,In_1350,In_353);
xor U494 (N_494,In_464,In_1319);
nand U495 (N_495,In_492,In_69);
nand U496 (N_496,In_27,In_1220);
and U497 (N_497,In_1070,In_1415);
or U498 (N_498,In_1069,In_155);
nand U499 (N_499,In_686,In_685);
or U500 (N_500,In_1272,N_106);
nand U501 (N_501,N_432,In_1028);
xor U502 (N_502,In_1269,N_255);
nor U503 (N_503,N_465,In_951);
nor U504 (N_504,N_439,In_236);
and U505 (N_505,N_350,In_188);
nor U506 (N_506,In_386,In_898);
xnor U507 (N_507,In_963,N_199);
and U508 (N_508,N_444,N_371);
or U509 (N_509,N_403,In_23);
and U510 (N_510,N_198,N_367);
nand U511 (N_511,In_828,In_204);
nor U512 (N_512,In_688,N_347);
or U513 (N_513,In_938,In_127);
nand U514 (N_514,In_670,N_31);
xor U515 (N_515,N_464,In_678);
and U516 (N_516,N_429,In_221);
nand U517 (N_517,In_1110,In_239);
nand U518 (N_518,N_69,In_38);
nand U519 (N_519,In_796,In_267);
nor U520 (N_520,In_857,N_478);
nor U521 (N_521,N_10,In_1395);
and U522 (N_522,N_492,In_119);
nor U523 (N_523,N_452,N_241);
nor U524 (N_524,N_254,N_153);
nor U525 (N_525,N_63,In_533);
or U526 (N_526,In_1247,N_411);
nand U527 (N_527,N_50,N_498);
nor U528 (N_528,In_90,In_1198);
nand U529 (N_529,N_384,N_156);
nor U530 (N_530,In_408,In_624);
nor U531 (N_531,N_321,In_1181);
nand U532 (N_532,In_802,In_1310);
or U533 (N_533,In_1325,In_266);
or U534 (N_534,N_377,N_318);
xor U535 (N_535,In_506,N_163);
xnor U536 (N_536,In_384,In_1372);
nand U537 (N_537,N_311,N_447);
nor U538 (N_538,N_74,In_650);
nor U539 (N_539,N_487,In_1065);
nor U540 (N_540,N_276,N_480);
nand U541 (N_541,N_326,In_891);
nand U542 (N_542,In_1201,N_18);
xor U543 (N_543,N_285,In_116);
and U544 (N_544,N_178,In_1215);
nor U545 (N_545,N_204,In_291);
nand U546 (N_546,In_1141,N_295);
xor U547 (N_547,In_1482,In_1150);
and U548 (N_548,N_23,In_974);
xnor U549 (N_549,N_64,N_190);
nand U550 (N_550,N_428,N_111);
and U551 (N_551,In_254,N_349);
and U552 (N_552,N_368,In_97);
nor U553 (N_553,In_347,In_305);
nand U554 (N_554,In_713,In_907);
or U555 (N_555,N_157,In_775);
or U556 (N_556,In_418,N_133);
nor U557 (N_557,In_764,N_192);
nand U558 (N_558,N_317,In_194);
or U559 (N_559,N_499,N_259);
or U560 (N_560,In_1073,N_107);
nand U561 (N_561,N_284,In_1252);
nand U562 (N_562,In_1240,N_258);
xnor U563 (N_563,N_485,In_368);
or U564 (N_564,N_3,N_414);
or U565 (N_565,N_183,In_109);
xnor U566 (N_566,N_116,In_1475);
and U567 (N_567,In_1018,In_1189);
and U568 (N_568,In_322,In_812);
xnor U569 (N_569,In_1470,N_59);
or U570 (N_570,In_667,In_1488);
and U571 (N_571,N_360,In_7);
xor U572 (N_572,In_1164,N_404);
and U573 (N_573,In_265,N_440);
xor U574 (N_574,N_450,N_474);
xnor U575 (N_575,In_1111,N_150);
or U576 (N_576,In_1307,In_414);
or U577 (N_577,In_284,In_580);
and U578 (N_578,N_271,In_850);
or U579 (N_579,In_583,N_427);
or U580 (N_580,N_108,N_421);
and U581 (N_581,N_82,In_1358);
nand U582 (N_582,N_324,N_152);
xor U583 (N_583,In_329,N_194);
nand U584 (N_584,N_379,N_328);
nor U585 (N_585,In_1459,In_1261);
nor U586 (N_586,In_777,In_1041);
and U587 (N_587,N_33,In_302);
and U588 (N_588,N_489,In_107);
or U589 (N_589,In_176,In_226);
and U590 (N_590,N_45,In_1169);
nand U591 (N_591,N_2,N_261);
nor U592 (N_592,N_305,In_1009);
and U593 (N_593,N_376,In_1281);
nand U594 (N_594,N_402,In_838);
or U595 (N_595,N_274,N_96);
or U596 (N_596,In_1155,N_296);
nor U597 (N_597,N_222,In_1085);
or U598 (N_598,N_177,In_407);
nor U599 (N_599,In_1288,In_1031);
xnor U600 (N_600,N_127,In_544);
nor U601 (N_601,N_84,N_331);
nor U602 (N_602,N_425,N_406);
nor U603 (N_603,N_236,N_209);
or U604 (N_604,In_512,N_313);
xnor U605 (N_605,In_1406,In_1066);
nor U606 (N_606,N_169,N_364);
nand U607 (N_607,In_784,In_921);
and U608 (N_608,In_549,N_456);
xor U609 (N_609,In_622,N_351);
or U610 (N_610,N_165,In_779);
and U611 (N_611,N_172,N_128);
xnor U612 (N_612,In_460,In_972);
xnor U613 (N_613,N_223,N_144);
xnor U614 (N_614,In_55,N_303);
xnor U615 (N_615,In_1102,In_211);
and U616 (N_616,N_378,In_269);
xor U617 (N_617,In_1087,N_4);
or U618 (N_618,In_478,In_341);
nor U619 (N_619,In_1122,N_265);
nand U620 (N_620,N_413,N_200);
nor U621 (N_621,In_932,In_1013);
or U622 (N_622,N_184,N_119);
nor U623 (N_623,N_47,N_308);
nor U624 (N_624,In_979,N_494);
or U625 (N_625,In_653,In_299);
nand U626 (N_626,In_545,N_55);
nor U627 (N_627,N_336,In_1327);
and U628 (N_628,In_1106,In_405);
or U629 (N_629,N_155,In_1015);
nand U630 (N_630,N_138,In_1380);
and U631 (N_631,N_85,N_345);
nor U632 (N_632,In_1250,N_80);
nand U633 (N_633,In_332,N_310);
or U634 (N_634,In_874,N_327);
xor U635 (N_635,In_645,N_216);
xor U636 (N_636,In_1373,N_0);
xor U637 (N_637,N_294,N_280);
nand U638 (N_638,N_417,In_683);
or U639 (N_639,In_749,In_1010);
nand U640 (N_640,N_160,N_139);
nor U641 (N_641,In_1457,N_176);
nand U642 (N_642,In_1218,In_1193);
nand U643 (N_643,In_1238,N_193);
and U644 (N_644,N_99,In_935);
and U645 (N_645,In_822,N_229);
nand U646 (N_646,N_179,In_496);
xnor U647 (N_647,N_353,In_1454);
nor U648 (N_648,In_660,N_112);
or U649 (N_649,In_1299,In_1485);
nand U650 (N_650,N_408,N_49);
xor U651 (N_651,N_479,N_297);
or U652 (N_652,N_182,N_468);
and U653 (N_653,N_34,In_1298);
nor U654 (N_654,In_1472,In_832);
nand U655 (N_655,N_391,In_693);
and U656 (N_656,In_1076,In_410);
xnor U657 (N_657,In_2,N_382);
xnor U658 (N_658,N_422,N_470);
xor U659 (N_659,N_81,N_48);
or U660 (N_660,In_1418,N_278);
nor U661 (N_661,N_231,N_338);
and U662 (N_662,In_203,N_466);
and U663 (N_663,N_197,In_259);
nor U664 (N_664,N_279,In_335);
xor U665 (N_665,In_813,In_106);
and U666 (N_666,N_30,In_708);
nor U667 (N_667,N_78,In_1292);
and U668 (N_668,In_636,In_707);
or U669 (N_669,N_245,In_1399);
nand U670 (N_670,In_1043,N_25);
nand U671 (N_671,N_214,N_400);
and U672 (N_672,In_1078,In_59);
and U673 (N_673,In_614,N_248);
and U674 (N_674,In_1098,In_321);
nand U675 (N_675,N_256,In_1025);
and U676 (N_676,N_235,In_717);
or U677 (N_677,In_803,N_307);
and U678 (N_678,N_252,In_101);
and U679 (N_679,In_228,N_292);
xor U680 (N_680,N_438,In_1363);
and U681 (N_681,N_443,In_32);
or U682 (N_682,N_221,In_729);
nand U683 (N_683,N_93,N_370);
and U684 (N_684,In_67,In_187);
nand U685 (N_685,N_185,In_374);
or U686 (N_686,In_1318,In_520);
or U687 (N_687,In_1268,N_94);
or U688 (N_688,N_14,In_726);
or U689 (N_689,In_1376,N_459);
nor U690 (N_690,In_355,In_870);
and U691 (N_691,N_394,In_960);
or U692 (N_692,N_120,In_334);
nor U693 (N_693,In_453,N_167);
or U694 (N_694,N_342,In_1489);
xor U695 (N_695,N_88,N_17);
xor U696 (N_696,In_924,In_711);
or U697 (N_697,In_861,In_1157);
and U698 (N_698,In_146,In_251);
nor U699 (N_699,In_830,In_1365);
or U700 (N_700,In_854,N_24);
xnor U701 (N_701,In_224,In_616);
or U702 (N_702,N_220,N_37);
and U703 (N_703,In_380,In_1417);
nor U704 (N_704,N_71,In_516);
xnor U705 (N_705,N_196,N_325);
or U706 (N_706,N_9,In_823);
or U707 (N_707,N_433,N_362);
and U708 (N_708,N_117,N_66);
nor U709 (N_709,In_525,In_306);
and U710 (N_710,In_767,In_770);
or U711 (N_711,In_440,N_39);
nor U712 (N_712,In_632,N_67);
nand U713 (N_713,N_475,In_993);
or U714 (N_714,In_510,N_344);
and U715 (N_715,In_1316,N_374);
nor U716 (N_716,In_621,In_844);
and U717 (N_717,N_335,N_282);
nand U718 (N_718,In_8,N_29);
nand U719 (N_719,N_20,N_314);
nand U720 (N_720,In_781,N_482);
nor U721 (N_721,N_363,In_747);
nor U722 (N_722,N_126,In_83);
and U723 (N_723,N_393,In_1001);
nor U724 (N_724,In_721,N_36);
nand U725 (N_725,N_334,N_109);
and U726 (N_726,N_287,In_411);
and U727 (N_727,In_180,N_442);
or U728 (N_728,In_765,N_113);
or U729 (N_729,N_419,In_160);
nor U730 (N_730,N_260,N_201);
nand U731 (N_731,N_385,N_215);
and U732 (N_732,In_375,In_626);
xnor U733 (N_733,N_124,In_40);
and U734 (N_734,N_340,N_356);
xnor U735 (N_735,In_1125,N_323);
and U736 (N_736,In_526,N_348);
and U737 (N_737,In_915,In_760);
or U738 (N_738,In_54,N_211);
or U739 (N_739,In_430,N_392);
nand U740 (N_740,In_1402,In_423);
xnor U741 (N_741,In_480,In_697);
nor U742 (N_742,In_1432,In_66);
nor U743 (N_743,In_825,In_482);
nand U744 (N_744,N_89,N_399);
xnor U745 (N_745,In_461,In_448);
xnor U746 (N_746,N_316,N_206);
or U747 (N_747,N_158,In_363);
nand U748 (N_748,N_268,N_416);
nand U749 (N_749,N_247,N_302);
or U750 (N_750,In_1105,In_885);
nand U751 (N_751,In_1217,In_36);
nor U752 (N_752,In_550,In_1476);
nor U753 (N_753,In_1359,N_398);
or U754 (N_754,N_135,In_189);
nand U755 (N_755,In_1456,N_44);
xor U756 (N_756,In_282,In_596);
nor U757 (N_757,In_820,In_207);
nor U758 (N_758,In_669,N_57);
xnor U759 (N_759,N_227,N_457);
nor U760 (N_760,N_86,In_263);
xor U761 (N_761,In_1020,N_46);
and U762 (N_762,In_744,In_360);
nor U763 (N_763,N_409,N_212);
and U764 (N_764,N_253,N_277);
nor U765 (N_765,N_180,In_117);
nand U766 (N_766,N_451,In_337);
or U767 (N_767,N_293,In_577);
xnor U768 (N_768,In_220,In_304);
xor U769 (N_769,N_463,In_446);
and U770 (N_770,N_110,N_6);
nor U771 (N_771,In_1375,N_224);
or U772 (N_772,In_142,In_514);
xnor U773 (N_773,N_15,In_283);
and U774 (N_774,In_354,N_481);
xnor U775 (N_775,N_51,In_486);
nor U776 (N_776,In_839,In_1263);
xor U777 (N_777,In_143,N_168);
and U778 (N_778,In_505,N_275);
and U779 (N_779,In_133,In_987);
nor U780 (N_780,N_161,In_601);
nand U781 (N_781,In_466,N_448);
or U782 (N_782,N_389,In_523);
nand U783 (N_783,In_859,In_565);
and U784 (N_784,In_186,In_477);
nand U785 (N_785,N_61,N_273);
or U786 (N_786,N_269,In_1302);
nand U787 (N_787,N_98,In_12);
nand U788 (N_788,N_175,In_42);
nand U789 (N_789,N_186,In_1397);
nand U790 (N_790,N_19,In_1332);
and U791 (N_791,N_130,In_297);
or U792 (N_792,In_98,N_154);
or U793 (N_793,N_396,In_1301);
nand U794 (N_794,N_435,N_92);
and U795 (N_795,N_309,N_52);
nand U796 (N_796,In_415,In_447);
nor U797 (N_797,N_125,N_242);
and U798 (N_798,N_497,N_170);
and U799 (N_799,N_387,N_251);
and U800 (N_800,N_380,N_12);
nand U801 (N_801,In_445,In_905);
or U802 (N_802,In_816,In_515);
and U803 (N_803,In_365,In_1427);
nand U804 (N_804,N_467,N_68);
or U805 (N_805,In_450,N_104);
xor U806 (N_806,N_257,In_1172);
nor U807 (N_807,N_208,N_121);
and U808 (N_808,N_441,In_362);
nand U809 (N_809,In_939,N_495);
xnor U810 (N_810,N_62,N_42);
xor U811 (N_811,In_205,In_367);
nor U812 (N_812,N_38,In_1429);
nand U813 (N_813,N_218,In_210);
xnor U814 (N_814,In_145,N_207);
nor U815 (N_815,In_1160,In_235);
xnor U816 (N_816,N_460,In_633);
nor U817 (N_817,N_486,N_202);
nand U818 (N_818,N_330,In_719);
and U819 (N_819,In_248,In_640);
and U820 (N_820,In_0,In_800);
nor U821 (N_821,In_238,In_436);
nor U822 (N_822,N_455,N_219);
xnor U823 (N_823,In_268,N_383);
nand U824 (N_824,N_137,In_592);
nor U825 (N_825,In_814,N_386);
and U826 (N_826,N_471,In_1004);
xor U827 (N_827,In_1113,N_237);
nand U828 (N_828,N_7,N_491);
nor U829 (N_829,In_888,In_46);
nor U830 (N_830,In_1101,N_75);
xnor U831 (N_831,N_476,N_332);
xnor U832 (N_832,In_925,N_449);
xnor U833 (N_833,N_21,In_50);
and U834 (N_834,N_239,In_498);
nor U835 (N_835,In_310,In_540);
or U836 (N_836,In_676,N_401);
nand U837 (N_837,In_395,N_355);
nand U838 (N_838,N_72,In_1322);
and U839 (N_839,N_203,N_381);
or U840 (N_840,N_73,In_381);
and U841 (N_841,N_164,N_372);
or U842 (N_842,N_267,In_513);
nor U843 (N_843,N_359,N_11);
xnor U844 (N_844,N_60,N_65);
or U845 (N_845,In_1271,In_136);
or U846 (N_846,N_143,N_304);
nor U847 (N_847,In_1422,In_1207);
and U848 (N_848,In_1219,In_923);
nand U849 (N_849,In_1014,In_658);
xor U850 (N_850,N_195,N_103);
xor U851 (N_851,In_366,N_420);
nor U852 (N_852,N_454,N_114);
nand U853 (N_853,In_1353,In_1407);
or U854 (N_854,In_955,In_654);
nor U855 (N_855,In_1461,N_228);
nand U856 (N_856,N_87,N_100);
or U857 (N_857,In_1284,In_663);
or U858 (N_858,N_397,N_418);
xnor U859 (N_859,In_85,N_249);
or U860 (N_860,In_364,In_1237);
nand U861 (N_861,N_5,N_244);
xnor U862 (N_862,N_188,In_1443);
or U863 (N_863,In_434,In_148);
nand U864 (N_864,N_390,In_572);
nand U865 (N_865,N_446,In_750);
xnor U866 (N_866,N_28,N_283);
xor U867 (N_867,N_35,In_1205);
and U868 (N_868,N_97,In_746);
nor U869 (N_869,N_306,In_1478);
xor U870 (N_870,In_1221,In_958);
or U871 (N_871,In_684,In_1400);
xor U872 (N_872,In_556,N_115);
nand U873 (N_873,In_208,N_477);
xor U874 (N_874,In_178,N_272);
or U875 (N_875,N_423,N_233);
and U876 (N_876,N_319,N_173);
and U877 (N_877,N_145,N_32);
nand U878 (N_878,In_443,N_246);
nand U879 (N_879,N_493,In_1354);
nand U880 (N_880,N_388,In_270);
nand U881 (N_881,In_1199,N_346);
xnor U882 (N_882,N_407,In_715);
and U883 (N_883,In_1216,N_16);
nand U884 (N_884,N_484,N_263);
and U885 (N_885,In_671,In_841);
nand U886 (N_886,N_95,N_105);
nor U887 (N_887,In_159,N_270);
xnor U888 (N_888,N_354,N_358);
and U889 (N_889,In_183,In_223);
xnor U890 (N_890,N_234,In_1471);
nand U891 (N_891,N_312,N_217);
nand U892 (N_892,N_122,In_899);
nor U893 (N_893,N_453,In_920);
nor U894 (N_894,In_49,In_325);
nand U895 (N_895,In_591,N_129);
and U896 (N_896,In_1011,N_166);
xnor U897 (N_897,In_348,N_462);
xor U898 (N_898,N_91,N_469);
or U899 (N_899,N_53,In_391);
and U900 (N_900,In_150,In_1450);
xor U901 (N_901,In_1030,N_286);
or U902 (N_902,In_1153,N_225);
or U903 (N_903,In_162,In_57);
nand U904 (N_904,N_369,In_536);
or U905 (N_905,N_434,In_274);
nor U906 (N_906,N_412,N_405);
and U907 (N_907,In_195,In_257);
xor U908 (N_908,N_210,In_1184);
nor U909 (N_909,N_70,In_84);
and U910 (N_910,In_883,N_232);
nand U911 (N_911,N_136,N_41);
or U912 (N_912,N_288,In_104);
xnor U913 (N_913,In_262,In_1243);
nor U914 (N_914,N_430,In_1235);
and U915 (N_915,N_230,N_373);
nor U916 (N_916,N_250,N_141);
or U917 (N_917,N_134,In_9);
and U918 (N_918,N_174,N_83);
and U919 (N_919,In_927,N_58);
nor U920 (N_920,N_77,N_361);
xnor U921 (N_921,N_90,N_79);
or U922 (N_922,In_1424,In_856);
nor U923 (N_923,In_462,In_481);
nand U924 (N_924,N_162,In_1467);
nand U925 (N_925,N_40,In_1340);
or U926 (N_926,N_76,N_262);
nor U927 (N_927,In_1379,N_473);
and U928 (N_928,N_123,In_1273);
nor U929 (N_929,In_1355,In_610);
and U930 (N_930,In_754,In_581);
and U931 (N_931,In_1042,In_277);
nand U932 (N_932,N_54,N_300);
and U933 (N_933,N_189,N_343);
xnor U934 (N_934,In_34,In_896);
nor U935 (N_935,N_264,N_329);
or U936 (N_936,In_690,In_981);
xor U937 (N_937,In_361,N_461);
and U938 (N_938,N_488,N_13);
or U939 (N_939,In_882,N_181);
and U940 (N_940,N_131,In_842);
nand U941 (N_941,N_315,In_1381);
and U942 (N_942,In_1494,N_226);
nor U943 (N_943,N_148,In_936);
and U944 (N_944,In_271,N_339);
or U945 (N_945,In_139,N_337);
or U946 (N_946,In_851,N_352);
or U947 (N_947,N_43,N_436);
and U948 (N_948,N_366,N_375);
xnor U949 (N_949,N_238,N_171);
xnor U950 (N_950,In_1394,In_1287);
nor U951 (N_951,In_1019,N_191);
nor U952 (N_952,In_1337,In_169);
nor U953 (N_953,N_243,In_88);
nor U954 (N_954,N_159,In_560);
nand U955 (N_955,In_1208,In_949);
xnor U956 (N_956,In_902,N_151);
or U957 (N_957,N_431,In_666);
or U958 (N_958,N_320,In_1195);
xor U959 (N_959,N_240,In_1466);
nand U960 (N_960,N_291,In_1420);
xor U961 (N_961,N_415,N_118);
xor U962 (N_962,In_1479,N_147);
xor U963 (N_963,N_290,N_365);
or U964 (N_964,N_101,In_952);
or U965 (N_965,N_142,In_1452);
nor U966 (N_966,In_1192,N_395);
or U967 (N_967,N_298,In_294);
nand U968 (N_968,N_357,N_281);
nand U969 (N_969,In_570,N_410);
nand U970 (N_970,In_1137,N_445);
or U971 (N_971,In_928,N_205);
xor U972 (N_972,N_496,In_517);
nand U973 (N_973,N_149,In_349);
nand U974 (N_974,N_187,In_1094);
or U975 (N_975,In_919,N_8);
nor U976 (N_976,N_341,N_299);
nand U977 (N_977,N_289,N_426);
or U978 (N_978,In_218,In_503);
or U979 (N_979,N_56,In_319);
nor U980 (N_980,In_1336,In_567);
xnor U981 (N_981,In_969,In_336);
and U982 (N_982,In_404,In_618);
or U983 (N_983,N_424,N_301);
and U984 (N_984,N_472,In_1123);
nand U985 (N_985,In_1309,In_138);
and U986 (N_986,In_810,N_132);
or U987 (N_987,N_22,N_333);
or U988 (N_988,In_385,N_102);
or U989 (N_989,In_867,N_483);
and U990 (N_990,N_266,N_213);
nor U991 (N_991,N_1,N_322);
xor U992 (N_992,In_463,In_652);
nand U993 (N_993,In_1486,In_1320);
or U994 (N_994,N_437,N_140);
nor U995 (N_995,In_475,N_27);
or U996 (N_996,In_788,In_181);
nand U997 (N_997,N_26,In_1321);
nor U998 (N_998,N_490,In_524);
or U999 (N_999,N_146,N_458);
xor U1000 (N_1000,N_536,N_914);
nand U1001 (N_1001,N_584,N_793);
and U1002 (N_1002,N_501,N_934);
nand U1003 (N_1003,N_818,N_560);
nand U1004 (N_1004,N_549,N_901);
or U1005 (N_1005,N_975,N_647);
or U1006 (N_1006,N_527,N_912);
xor U1007 (N_1007,N_814,N_736);
and U1008 (N_1008,N_553,N_844);
xnor U1009 (N_1009,N_625,N_713);
xnor U1010 (N_1010,N_548,N_731);
and U1011 (N_1011,N_869,N_595);
xor U1012 (N_1012,N_542,N_689);
nor U1013 (N_1013,N_999,N_730);
xnor U1014 (N_1014,N_760,N_623);
and U1015 (N_1015,N_950,N_575);
nor U1016 (N_1016,N_994,N_929);
xnor U1017 (N_1017,N_962,N_587);
or U1018 (N_1018,N_649,N_700);
nand U1019 (N_1019,N_905,N_770);
or U1020 (N_1020,N_969,N_831);
nand U1021 (N_1021,N_692,N_965);
nor U1022 (N_1022,N_617,N_616);
nand U1023 (N_1023,N_507,N_723);
nand U1024 (N_1024,N_634,N_669);
or U1025 (N_1025,N_932,N_976);
or U1026 (N_1026,N_897,N_904);
or U1027 (N_1027,N_956,N_676);
or U1028 (N_1028,N_528,N_907);
and U1029 (N_1029,N_564,N_534);
and U1030 (N_1030,N_550,N_555);
or U1031 (N_1031,N_574,N_985);
nand U1032 (N_1032,N_803,N_675);
xnor U1033 (N_1033,N_558,N_637);
and U1034 (N_1034,N_936,N_817);
nand U1035 (N_1035,N_571,N_748);
xor U1036 (N_1036,N_853,N_604);
xnor U1037 (N_1037,N_735,N_636);
xnor U1038 (N_1038,N_525,N_832);
xnor U1039 (N_1039,N_643,N_833);
nor U1040 (N_1040,N_543,N_761);
xnor U1041 (N_1041,N_751,N_513);
xnor U1042 (N_1042,N_737,N_658);
or U1043 (N_1043,N_910,N_695);
nor U1044 (N_1044,N_684,N_685);
nor U1045 (N_1045,N_615,N_997);
and U1046 (N_1046,N_876,N_955);
xnor U1047 (N_1047,N_709,N_742);
xnor U1048 (N_1048,N_576,N_788);
nand U1049 (N_1049,N_754,N_674);
xor U1050 (N_1050,N_570,N_941);
nand U1051 (N_1051,N_886,N_632);
nand U1052 (N_1052,N_820,N_919);
nor U1053 (N_1053,N_834,N_600);
nand U1054 (N_1054,N_593,N_728);
nor U1055 (N_1055,N_511,N_538);
xnor U1056 (N_1056,N_982,N_611);
nor U1057 (N_1057,N_644,N_772);
nor U1058 (N_1058,N_966,N_654);
nor U1059 (N_1059,N_948,N_890);
nand U1060 (N_1060,N_927,N_870);
nor U1061 (N_1061,N_628,N_924);
or U1062 (N_1062,N_992,N_752);
nand U1063 (N_1063,N_518,N_978);
and U1064 (N_1064,N_609,N_763);
and U1065 (N_1065,N_704,N_718);
nor U1066 (N_1066,N_896,N_509);
nand U1067 (N_1067,N_958,N_586);
xor U1068 (N_1068,N_638,N_865);
or U1069 (N_1069,N_660,N_579);
nor U1070 (N_1070,N_913,N_863);
and U1071 (N_1071,N_672,N_835);
nand U1072 (N_1072,N_783,N_755);
or U1073 (N_1073,N_724,N_727);
nand U1074 (N_1074,N_712,N_809);
nor U1075 (N_1075,N_830,N_597);
xor U1076 (N_1076,N_661,N_598);
and U1077 (N_1077,N_882,N_531);
and U1078 (N_1078,N_762,N_977);
nand U1079 (N_1079,N_603,N_627);
nand U1080 (N_1080,N_878,N_699);
xnor U1081 (N_1081,N_729,N_899);
nor U1082 (N_1082,N_665,N_562);
nand U1083 (N_1083,N_795,N_745);
and U1084 (N_1084,N_726,N_701);
xor U1085 (N_1085,N_590,N_565);
nor U1086 (N_1086,N_756,N_512);
nand U1087 (N_1087,N_650,N_959);
xor U1088 (N_1088,N_743,N_859);
xnor U1089 (N_1089,N_906,N_781);
nand U1090 (N_1090,N_851,N_871);
nor U1091 (N_1091,N_554,N_757);
or U1092 (N_1092,N_813,N_630);
or U1093 (N_1093,N_903,N_894);
and U1094 (N_1094,N_786,N_846);
xnor U1095 (N_1095,N_995,N_900);
or U1096 (N_1096,N_990,N_884);
nand U1097 (N_1097,N_662,N_891);
and U1098 (N_1098,N_867,N_629);
xnor U1099 (N_1099,N_670,N_708);
nand U1100 (N_1100,N_785,N_979);
nand U1101 (N_1101,N_552,N_522);
nor U1102 (N_1102,N_920,N_508);
and U1103 (N_1103,N_816,N_922);
nor U1104 (N_1104,N_721,N_860);
or U1105 (N_1105,N_688,N_697);
xnor U1106 (N_1106,N_987,N_502);
nor U1107 (N_1107,N_622,N_881);
nand U1108 (N_1108,N_974,N_691);
nor U1109 (N_1109,N_648,N_705);
or U1110 (N_1110,N_750,N_510);
nor U1111 (N_1111,N_917,N_961);
nand U1112 (N_1112,N_864,N_523);
and U1113 (N_1113,N_874,N_766);
or U1114 (N_1114,N_861,N_633);
nor U1115 (N_1115,N_696,N_848);
or U1116 (N_1116,N_799,N_779);
nor U1117 (N_1117,N_667,N_681);
xor U1118 (N_1118,N_946,N_619);
or U1119 (N_1119,N_892,N_624);
nand U1120 (N_1120,N_811,N_569);
nor U1121 (N_1121,N_559,N_828);
or U1122 (N_1122,N_812,N_521);
or U1123 (N_1123,N_725,N_690);
nand U1124 (N_1124,N_937,N_707);
and U1125 (N_1125,N_683,N_631);
and U1126 (N_1126,N_621,N_532);
nor U1127 (N_1127,N_592,N_953);
nand U1128 (N_1128,N_822,N_711);
and U1129 (N_1129,N_849,N_916);
nor U1130 (N_1130,N_767,N_942);
and U1131 (N_1131,N_952,N_773);
nor U1132 (N_1132,N_970,N_640);
nor U1133 (N_1133,N_939,N_957);
nor U1134 (N_1134,N_657,N_928);
xnor U1135 (N_1135,N_732,N_733);
or U1136 (N_1136,N_719,N_796);
or U1137 (N_1137,N_819,N_840);
nor U1138 (N_1138,N_734,N_666);
xnor U1139 (N_1139,N_653,N_971);
and U1140 (N_1140,N_545,N_673);
xor U1141 (N_1141,N_607,N_687);
or U1142 (N_1142,N_606,N_893);
or U1143 (N_1143,N_677,N_664);
and U1144 (N_1144,N_608,N_964);
nand U1145 (N_1145,N_854,N_573);
nand U1146 (N_1146,N_544,N_563);
nand U1147 (N_1147,N_949,N_626);
nor U1148 (N_1148,N_923,N_868);
and U1149 (N_1149,N_535,N_612);
xnor U1150 (N_1150,N_680,N_645);
and U1151 (N_1151,N_517,N_983);
xor U1152 (N_1152,N_682,N_506);
nor U1153 (N_1153,N_557,N_790);
nor U1154 (N_1154,N_533,N_710);
and U1155 (N_1155,N_826,N_940);
xnor U1156 (N_1156,N_850,N_614);
nor U1157 (N_1157,N_591,N_808);
and U1158 (N_1158,N_815,N_989);
nand U1159 (N_1159,N_679,N_663);
or U1160 (N_1160,N_872,N_561);
nor U1161 (N_1161,N_659,N_526);
nor U1162 (N_1162,N_519,N_769);
and U1163 (N_1163,N_778,N_858);
and U1164 (N_1164,N_933,N_739);
or U1165 (N_1165,N_980,N_596);
xor U1166 (N_1166,N_885,N_520);
nor U1167 (N_1167,N_879,N_837);
and U1168 (N_1168,N_960,N_702);
nand U1169 (N_1169,N_551,N_930);
nand U1170 (N_1170,N_805,N_524);
nand U1171 (N_1171,N_909,N_836);
nand U1172 (N_1172,N_856,N_798);
nor U1173 (N_1173,N_740,N_911);
xnor U1174 (N_1174,N_635,N_567);
xnor U1175 (N_1175,N_686,N_807);
xor U1176 (N_1176,N_541,N_988);
xnor U1177 (N_1177,N_577,N_503);
nand U1178 (N_1178,N_694,N_972);
nand U1179 (N_1179,N_852,N_986);
nor U1180 (N_1180,N_618,N_887);
and U1181 (N_1181,N_605,N_825);
nand U1182 (N_1182,N_540,N_877);
xnor U1183 (N_1183,N_866,N_505);
and U1184 (N_1184,N_652,N_578);
xnor U1185 (N_1185,N_973,N_599);
nand U1186 (N_1186,N_945,N_500);
and U1187 (N_1187,N_775,N_935);
nor U1188 (N_1188,N_791,N_824);
and U1189 (N_1189,N_780,N_529);
or U1190 (N_1190,N_749,N_610);
and U1191 (N_1191,N_698,N_847);
and U1192 (N_1192,N_585,N_794);
and U1193 (N_1193,N_880,N_537);
or U1194 (N_1194,N_895,N_806);
and U1195 (N_1195,N_855,N_993);
nor U1196 (N_1196,N_947,N_646);
or U1197 (N_1197,N_758,N_714);
or U1198 (N_1198,N_656,N_842);
xor U1199 (N_1199,N_589,N_804);
nor U1200 (N_1200,N_764,N_792);
nand U1201 (N_1201,N_841,N_642);
and U1202 (N_1202,N_668,N_944);
nor U1203 (N_1203,N_581,N_765);
and U1204 (N_1204,N_539,N_873);
and U1205 (N_1205,N_580,N_594);
nand U1206 (N_1206,N_991,N_801);
nand U1207 (N_1207,N_931,N_938);
nand U1208 (N_1208,N_921,N_898);
nor U1209 (N_1209,N_823,N_845);
nor U1210 (N_1210,N_883,N_514);
nand U1211 (N_1211,N_546,N_620);
nand U1212 (N_1212,N_918,N_703);
nor U1213 (N_1213,N_968,N_789);
and U1214 (N_1214,N_888,N_601);
xnor U1215 (N_1215,N_943,N_530);
nor U1216 (N_1216,N_821,N_715);
or U1217 (N_1217,N_588,N_777);
and U1218 (N_1218,N_744,N_768);
nand U1219 (N_1219,N_678,N_797);
xor U1220 (N_1220,N_515,N_655);
or U1221 (N_1221,N_613,N_504);
and U1222 (N_1222,N_566,N_651);
nor U1223 (N_1223,N_875,N_827);
and U1224 (N_1224,N_829,N_810);
nand U1225 (N_1225,N_902,N_720);
and U1226 (N_1226,N_753,N_926);
and U1227 (N_1227,N_717,N_641);
or U1228 (N_1228,N_889,N_784);
and U1229 (N_1229,N_954,N_747);
or U1230 (N_1230,N_963,N_925);
xnor U1231 (N_1231,N_996,N_516);
nor U1232 (N_1232,N_771,N_967);
or U1233 (N_1233,N_639,N_671);
nand U1234 (N_1234,N_547,N_843);
nand U1235 (N_1235,N_782,N_915);
nor U1236 (N_1236,N_706,N_759);
or U1237 (N_1237,N_568,N_602);
nand U1238 (N_1238,N_838,N_693);
or U1239 (N_1239,N_582,N_800);
or U1240 (N_1240,N_716,N_774);
nor U1241 (N_1241,N_908,N_746);
and U1242 (N_1242,N_572,N_981);
and U1243 (N_1243,N_787,N_776);
and U1244 (N_1244,N_722,N_839);
or U1245 (N_1245,N_738,N_984);
and U1246 (N_1246,N_802,N_583);
and U1247 (N_1247,N_741,N_556);
and U1248 (N_1248,N_862,N_998);
nand U1249 (N_1249,N_951,N_857);
xor U1250 (N_1250,N_892,N_941);
xor U1251 (N_1251,N_752,N_567);
nor U1252 (N_1252,N_573,N_655);
nor U1253 (N_1253,N_887,N_740);
nor U1254 (N_1254,N_937,N_761);
nand U1255 (N_1255,N_956,N_754);
nor U1256 (N_1256,N_522,N_538);
nor U1257 (N_1257,N_893,N_806);
nor U1258 (N_1258,N_631,N_675);
and U1259 (N_1259,N_572,N_952);
xor U1260 (N_1260,N_791,N_528);
nor U1261 (N_1261,N_652,N_558);
xor U1262 (N_1262,N_688,N_792);
xnor U1263 (N_1263,N_840,N_593);
nand U1264 (N_1264,N_730,N_833);
or U1265 (N_1265,N_675,N_846);
nand U1266 (N_1266,N_590,N_839);
or U1267 (N_1267,N_723,N_728);
or U1268 (N_1268,N_721,N_686);
xor U1269 (N_1269,N_926,N_908);
and U1270 (N_1270,N_631,N_855);
and U1271 (N_1271,N_575,N_937);
and U1272 (N_1272,N_993,N_990);
and U1273 (N_1273,N_653,N_798);
or U1274 (N_1274,N_641,N_580);
nand U1275 (N_1275,N_622,N_772);
and U1276 (N_1276,N_944,N_581);
xor U1277 (N_1277,N_597,N_956);
and U1278 (N_1278,N_859,N_536);
and U1279 (N_1279,N_588,N_738);
nand U1280 (N_1280,N_572,N_968);
nand U1281 (N_1281,N_798,N_759);
nor U1282 (N_1282,N_683,N_994);
and U1283 (N_1283,N_524,N_753);
nand U1284 (N_1284,N_765,N_981);
and U1285 (N_1285,N_647,N_825);
nand U1286 (N_1286,N_697,N_534);
or U1287 (N_1287,N_767,N_603);
nand U1288 (N_1288,N_838,N_529);
or U1289 (N_1289,N_925,N_507);
nor U1290 (N_1290,N_917,N_627);
and U1291 (N_1291,N_794,N_648);
and U1292 (N_1292,N_624,N_752);
nand U1293 (N_1293,N_899,N_620);
nand U1294 (N_1294,N_822,N_931);
xor U1295 (N_1295,N_662,N_674);
nor U1296 (N_1296,N_893,N_703);
or U1297 (N_1297,N_707,N_530);
nor U1298 (N_1298,N_996,N_565);
nand U1299 (N_1299,N_644,N_597);
or U1300 (N_1300,N_945,N_952);
nand U1301 (N_1301,N_858,N_741);
nand U1302 (N_1302,N_985,N_563);
and U1303 (N_1303,N_968,N_800);
or U1304 (N_1304,N_981,N_899);
xnor U1305 (N_1305,N_740,N_633);
xor U1306 (N_1306,N_682,N_975);
and U1307 (N_1307,N_991,N_800);
nor U1308 (N_1308,N_516,N_869);
and U1309 (N_1309,N_901,N_621);
and U1310 (N_1310,N_737,N_913);
or U1311 (N_1311,N_930,N_958);
xor U1312 (N_1312,N_952,N_707);
nor U1313 (N_1313,N_630,N_968);
nand U1314 (N_1314,N_591,N_684);
nand U1315 (N_1315,N_824,N_881);
nor U1316 (N_1316,N_845,N_851);
nand U1317 (N_1317,N_733,N_998);
and U1318 (N_1318,N_655,N_915);
nand U1319 (N_1319,N_715,N_975);
nor U1320 (N_1320,N_661,N_644);
xor U1321 (N_1321,N_633,N_702);
xor U1322 (N_1322,N_770,N_673);
nor U1323 (N_1323,N_713,N_608);
nand U1324 (N_1324,N_798,N_816);
or U1325 (N_1325,N_869,N_975);
and U1326 (N_1326,N_955,N_831);
or U1327 (N_1327,N_892,N_643);
nor U1328 (N_1328,N_970,N_527);
or U1329 (N_1329,N_934,N_836);
and U1330 (N_1330,N_718,N_590);
or U1331 (N_1331,N_681,N_722);
or U1332 (N_1332,N_611,N_861);
nor U1333 (N_1333,N_631,N_861);
or U1334 (N_1334,N_509,N_869);
or U1335 (N_1335,N_807,N_821);
nand U1336 (N_1336,N_966,N_920);
xor U1337 (N_1337,N_510,N_931);
nor U1338 (N_1338,N_550,N_776);
or U1339 (N_1339,N_967,N_964);
xor U1340 (N_1340,N_732,N_776);
and U1341 (N_1341,N_634,N_528);
xor U1342 (N_1342,N_564,N_622);
nand U1343 (N_1343,N_693,N_663);
and U1344 (N_1344,N_877,N_785);
nor U1345 (N_1345,N_648,N_734);
nor U1346 (N_1346,N_596,N_801);
or U1347 (N_1347,N_582,N_651);
or U1348 (N_1348,N_965,N_628);
or U1349 (N_1349,N_913,N_517);
nand U1350 (N_1350,N_741,N_941);
or U1351 (N_1351,N_538,N_821);
and U1352 (N_1352,N_948,N_872);
xnor U1353 (N_1353,N_520,N_584);
nor U1354 (N_1354,N_915,N_844);
nor U1355 (N_1355,N_759,N_904);
or U1356 (N_1356,N_615,N_573);
xnor U1357 (N_1357,N_949,N_699);
nor U1358 (N_1358,N_957,N_714);
xor U1359 (N_1359,N_664,N_693);
nor U1360 (N_1360,N_693,N_529);
or U1361 (N_1361,N_623,N_548);
or U1362 (N_1362,N_578,N_711);
and U1363 (N_1363,N_647,N_880);
and U1364 (N_1364,N_800,N_546);
and U1365 (N_1365,N_645,N_731);
or U1366 (N_1366,N_761,N_877);
or U1367 (N_1367,N_822,N_696);
nor U1368 (N_1368,N_795,N_986);
and U1369 (N_1369,N_962,N_691);
nor U1370 (N_1370,N_995,N_917);
and U1371 (N_1371,N_651,N_836);
and U1372 (N_1372,N_893,N_575);
nor U1373 (N_1373,N_545,N_979);
nand U1374 (N_1374,N_537,N_811);
and U1375 (N_1375,N_882,N_561);
nor U1376 (N_1376,N_899,N_887);
and U1377 (N_1377,N_595,N_836);
nor U1378 (N_1378,N_711,N_777);
xnor U1379 (N_1379,N_885,N_810);
or U1380 (N_1380,N_634,N_861);
xnor U1381 (N_1381,N_817,N_929);
and U1382 (N_1382,N_997,N_689);
nand U1383 (N_1383,N_811,N_953);
nor U1384 (N_1384,N_788,N_962);
nand U1385 (N_1385,N_553,N_669);
and U1386 (N_1386,N_773,N_673);
nor U1387 (N_1387,N_581,N_636);
nor U1388 (N_1388,N_994,N_960);
nor U1389 (N_1389,N_802,N_691);
nand U1390 (N_1390,N_795,N_779);
or U1391 (N_1391,N_592,N_706);
nor U1392 (N_1392,N_616,N_974);
nor U1393 (N_1393,N_707,N_951);
or U1394 (N_1394,N_904,N_755);
nand U1395 (N_1395,N_718,N_509);
nand U1396 (N_1396,N_717,N_533);
or U1397 (N_1397,N_977,N_594);
or U1398 (N_1398,N_501,N_514);
and U1399 (N_1399,N_537,N_856);
and U1400 (N_1400,N_948,N_673);
nand U1401 (N_1401,N_979,N_653);
and U1402 (N_1402,N_682,N_710);
xor U1403 (N_1403,N_710,N_915);
nor U1404 (N_1404,N_608,N_533);
and U1405 (N_1405,N_520,N_913);
or U1406 (N_1406,N_645,N_505);
or U1407 (N_1407,N_788,N_771);
xor U1408 (N_1408,N_794,N_996);
nor U1409 (N_1409,N_849,N_856);
xnor U1410 (N_1410,N_850,N_538);
and U1411 (N_1411,N_797,N_898);
nand U1412 (N_1412,N_849,N_502);
and U1413 (N_1413,N_558,N_778);
xor U1414 (N_1414,N_672,N_863);
nor U1415 (N_1415,N_988,N_536);
nor U1416 (N_1416,N_672,N_854);
nor U1417 (N_1417,N_614,N_812);
or U1418 (N_1418,N_539,N_865);
xor U1419 (N_1419,N_707,N_785);
or U1420 (N_1420,N_747,N_781);
nor U1421 (N_1421,N_787,N_708);
nor U1422 (N_1422,N_528,N_972);
nor U1423 (N_1423,N_567,N_648);
xor U1424 (N_1424,N_731,N_928);
nand U1425 (N_1425,N_915,N_862);
nor U1426 (N_1426,N_546,N_974);
xnor U1427 (N_1427,N_932,N_651);
nand U1428 (N_1428,N_884,N_815);
nor U1429 (N_1429,N_729,N_731);
nor U1430 (N_1430,N_968,N_643);
nand U1431 (N_1431,N_832,N_968);
nor U1432 (N_1432,N_870,N_686);
nor U1433 (N_1433,N_830,N_569);
and U1434 (N_1434,N_873,N_816);
nand U1435 (N_1435,N_536,N_996);
and U1436 (N_1436,N_741,N_887);
nand U1437 (N_1437,N_777,N_947);
xnor U1438 (N_1438,N_742,N_642);
nor U1439 (N_1439,N_638,N_527);
nor U1440 (N_1440,N_779,N_796);
nor U1441 (N_1441,N_891,N_569);
nor U1442 (N_1442,N_775,N_602);
xor U1443 (N_1443,N_975,N_796);
xor U1444 (N_1444,N_892,N_832);
and U1445 (N_1445,N_723,N_784);
and U1446 (N_1446,N_984,N_534);
nand U1447 (N_1447,N_939,N_630);
nor U1448 (N_1448,N_879,N_994);
xor U1449 (N_1449,N_831,N_657);
and U1450 (N_1450,N_571,N_896);
nand U1451 (N_1451,N_620,N_896);
or U1452 (N_1452,N_810,N_712);
xnor U1453 (N_1453,N_682,N_593);
or U1454 (N_1454,N_662,N_852);
nand U1455 (N_1455,N_918,N_621);
xor U1456 (N_1456,N_615,N_761);
nand U1457 (N_1457,N_759,N_589);
nand U1458 (N_1458,N_979,N_790);
nand U1459 (N_1459,N_580,N_549);
or U1460 (N_1460,N_909,N_989);
and U1461 (N_1461,N_908,N_843);
nor U1462 (N_1462,N_947,N_538);
and U1463 (N_1463,N_690,N_580);
nor U1464 (N_1464,N_991,N_782);
nor U1465 (N_1465,N_860,N_975);
and U1466 (N_1466,N_846,N_555);
and U1467 (N_1467,N_991,N_969);
nand U1468 (N_1468,N_775,N_850);
and U1469 (N_1469,N_732,N_804);
or U1470 (N_1470,N_747,N_822);
and U1471 (N_1471,N_974,N_640);
nand U1472 (N_1472,N_690,N_593);
xor U1473 (N_1473,N_926,N_833);
xnor U1474 (N_1474,N_571,N_910);
xor U1475 (N_1475,N_659,N_842);
or U1476 (N_1476,N_755,N_943);
and U1477 (N_1477,N_748,N_790);
nor U1478 (N_1478,N_832,N_548);
nor U1479 (N_1479,N_828,N_672);
and U1480 (N_1480,N_921,N_975);
xor U1481 (N_1481,N_937,N_999);
nor U1482 (N_1482,N_639,N_542);
xor U1483 (N_1483,N_540,N_901);
xor U1484 (N_1484,N_895,N_751);
nor U1485 (N_1485,N_695,N_732);
xor U1486 (N_1486,N_828,N_928);
xor U1487 (N_1487,N_742,N_614);
nor U1488 (N_1488,N_551,N_733);
xnor U1489 (N_1489,N_585,N_738);
nor U1490 (N_1490,N_921,N_508);
nand U1491 (N_1491,N_849,N_554);
xnor U1492 (N_1492,N_961,N_755);
and U1493 (N_1493,N_980,N_568);
nor U1494 (N_1494,N_736,N_833);
and U1495 (N_1495,N_792,N_844);
nor U1496 (N_1496,N_763,N_509);
and U1497 (N_1497,N_551,N_791);
and U1498 (N_1498,N_800,N_562);
or U1499 (N_1499,N_629,N_621);
nand U1500 (N_1500,N_1287,N_1474);
nor U1501 (N_1501,N_1019,N_1407);
or U1502 (N_1502,N_1368,N_1105);
and U1503 (N_1503,N_1208,N_1459);
nand U1504 (N_1504,N_1106,N_1126);
xnor U1505 (N_1505,N_1033,N_1216);
and U1506 (N_1506,N_1487,N_1274);
and U1507 (N_1507,N_1046,N_1427);
and U1508 (N_1508,N_1207,N_1484);
or U1509 (N_1509,N_1099,N_1113);
xor U1510 (N_1510,N_1316,N_1047);
nor U1511 (N_1511,N_1095,N_1074);
xnor U1512 (N_1512,N_1263,N_1029);
and U1513 (N_1513,N_1193,N_1058);
and U1514 (N_1514,N_1419,N_1417);
and U1515 (N_1515,N_1314,N_1203);
or U1516 (N_1516,N_1006,N_1110);
nor U1517 (N_1517,N_1009,N_1396);
or U1518 (N_1518,N_1444,N_1431);
xor U1519 (N_1519,N_1486,N_1433);
nand U1520 (N_1520,N_1172,N_1248);
nor U1521 (N_1521,N_1356,N_1189);
xor U1522 (N_1522,N_1461,N_1395);
or U1523 (N_1523,N_1082,N_1376);
or U1524 (N_1524,N_1219,N_1261);
nor U1525 (N_1525,N_1123,N_1155);
and U1526 (N_1526,N_1138,N_1390);
xnor U1527 (N_1527,N_1477,N_1035);
nor U1528 (N_1528,N_1100,N_1022);
or U1529 (N_1529,N_1323,N_1069);
xnor U1530 (N_1530,N_1067,N_1150);
nand U1531 (N_1531,N_1480,N_1363);
nor U1532 (N_1532,N_1247,N_1039);
nor U1533 (N_1533,N_1142,N_1490);
or U1534 (N_1534,N_1447,N_1340);
or U1535 (N_1535,N_1320,N_1332);
and U1536 (N_1536,N_1023,N_1346);
and U1537 (N_1537,N_1092,N_1278);
or U1538 (N_1538,N_1276,N_1239);
nor U1539 (N_1539,N_1204,N_1195);
nand U1540 (N_1540,N_1060,N_1124);
or U1541 (N_1541,N_1325,N_1233);
nor U1542 (N_1542,N_1385,N_1494);
and U1543 (N_1543,N_1334,N_1014);
xnor U1544 (N_1544,N_1243,N_1436);
or U1545 (N_1545,N_1168,N_1007);
and U1546 (N_1546,N_1202,N_1259);
nand U1547 (N_1547,N_1296,N_1107);
xor U1548 (N_1548,N_1299,N_1191);
and U1549 (N_1549,N_1140,N_1054);
nor U1550 (N_1550,N_1037,N_1045);
nor U1551 (N_1551,N_1442,N_1435);
or U1552 (N_1552,N_1268,N_1291);
and U1553 (N_1553,N_1463,N_1075);
or U1554 (N_1554,N_1430,N_1156);
nand U1555 (N_1555,N_1388,N_1324);
xnor U1556 (N_1556,N_1351,N_1429);
or U1557 (N_1557,N_1178,N_1416);
nand U1558 (N_1558,N_1297,N_1499);
or U1559 (N_1559,N_1042,N_1177);
nand U1560 (N_1560,N_1017,N_1162);
nand U1561 (N_1561,N_1311,N_1294);
xor U1562 (N_1562,N_1066,N_1224);
or U1563 (N_1563,N_1302,N_1098);
nand U1564 (N_1564,N_1111,N_1466);
or U1565 (N_1565,N_1222,N_1174);
nor U1566 (N_1566,N_1370,N_1031);
and U1567 (N_1567,N_1088,N_1161);
or U1568 (N_1568,N_1425,N_1212);
or U1569 (N_1569,N_1280,N_1115);
and U1570 (N_1570,N_1360,N_1049);
or U1571 (N_1571,N_1264,N_1437);
and U1572 (N_1572,N_1077,N_1192);
nand U1573 (N_1573,N_1364,N_1026);
nand U1574 (N_1574,N_1333,N_1218);
or U1575 (N_1575,N_1104,N_1375);
nor U1576 (N_1576,N_1227,N_1034);
and U1577 (N_1577,N_1257,N_1420);
and U1578 (N_1578,N_1310,N_1374);
nand U1579 (N_1579,N_1462,N_1167);
nor U1580 (N_1580,N_1065,N_1262);
xnor U1581 (N_1581,N_1496,N_1118);
or U1582 (N_1582,N_1116,N_1139);
nand U1583 (N_1583,N_1258,N_1186);
or U1584 (N_1584,N_1144,N_1488);
xnor U1585 (N_1585,N_1392,N_1336);
or U1586 (N_1586,N_1215,N_1093);
and U1587 (N_1587,N_1440,N_1321);
xor U1588 (N_1588,N_1358,N_1160);
nand U1589 (N_1589,N_1357,N_1322);
nand U1590 (N_1590,N_1331,N_1327);
and U1591 (N_1591,N_1483,N_1498);
or U1592 (N_1592,N_1415,N_1284);
and U1593 (N_1593,N_1032,N_1152);
nor U1594 (N_1594,N_1128,N_1410);
nor U1595 (N_1595,N_1236,N_1305);
and U1596 (N_1596,N_1256,N_1085);
nand U1597 (N_1597,N_1379,N_1101);
and U1598 (N_1598,N_1005,N_1412);
xnor U1599 (N_1599,N_1080,N_1306);
and U1600 (N_1600,N_1485,N_1328);
nand U1601 (N_1601,N_1438,N_1010);
nor U1602 (N_1602,N_1460,N_1478);
or U1603 (N_1603,N_1348,N_1362);
nand U1604 (N_1604,N_1073,N_1072);
or U1605 (N_1605,N_1000,N_1057);
and U1606 (N_1606,N_1345,N_1397);
nor U1607 (N_1607,N_1103,N_1163);
and U1608 (N_1608,N_1451,N_1063);
nand U1609 (N_1609,N_1076,N_1468);
nor U1610 (N_1610,N_1170,N_1350);
nor U1611 (N_1611,N_1020,N_1359);
and U1612 (N_1612,N_1381,N_1015);
xnor U1613 (N_1613,N_1176,N_1053);
and U1614 (N_1614,N_1183,N_1091);
xnor U1615 (N_1615,N_1024,N_1025);
nand U1616 (N_1616,N_1141,N_1120);
nor U1617 (N_1617,N_1471,N_1279);
nor U1618 (N_1618,N_1414,N_1282);
xor U1619 (N_1619,N_1040,N_1267);
and U1620 (N_1620,N_1454,N_1084);
or U1621 (N_1621,N_1181,N_1326);
nor U1622 (N_1622,N_1117,N_1179);
xnor U1623 (N_1623,N_1044,N_1151);
nand U1624 (N_1624,N_1081,N_1246);
and U1625 (N_1625,N_1145,N_1221);
xnor U1626 (N_1626,N_1061,N_1458);
nor U1627 (N_1627,N_1071,N_1289);
and U1628 (N_1628,N_1200,N_1241);
nor U1629 (N_1629,N_1226,N_1229);
and U1630 (N_1630,N_1411,N_1011);
nand U1631 (N_1631,N_1055,N_1197);
and U1632 (N_1632,N_1062,N_1249);
or U1633 (N_1633,N_1403,N_1021);
or U1634 (N_1634,N_1149,N_1109);
xor U1635 (N_1635,N_1122,N_1402);
and U1636 (N_1636,N_1406,N_1159);
nor U1637 (N_1637,N_1464,N_1030);
nor U1638 (N_1638,N_1232,N_1408);
nor U1639 (N_1639,N_1108,N_1309);
nor U1640 (N_1640,N_1255,N_1387);
nand U1641 (N_1641,N_1070,N_1449);
xnor U1642 (N_1642,N_1050,N_1409);
xor U1643 (N_1643,N_1421,N_1273);
and U1644 (N_1644,N_1231,N_1225);
xnor U1645 (N_1645,N_1335,N_1114);
xor U1646 (N_1646,N_1164,N_1377);
xnor U1647 (N_1647,N_1265,N_1016);
and U1648 (N_1648,N_1217,N_1426);
and U1649 (N_1649,N_1180,N_1173);
and U1650 (N_1650,N_1457,N_1295);
xor U1651 (N_1651,N_1389,N_1446);
nand U1652 (N_1652,N_1059,N_1251);
or U1653 (N_1653,N_1228,N_1441);
and U1654 (N_1654,N_1313,N_1254);
and U1655 (N_1655,N_1482,N_1018);
or U1656 (N_1656,N_1472,N_1079);
nor U1657 (N_1657,N_1382,N_1300);
nand U1658 (N_1658,N_1166,N_1384);
xnor U1659 (N_1659,N_1242,N_1004);
xnor U1660 (N_1660,N_1473,N_1234);
nand U1661 (N_1661,N_1450,N_1285);
or U1662 (N_1662,N_1354,N_1470);
and U1663 (N_1663,N_1400,N_1210);
nor U1664 (N_1664,N_1132,N_1068);
xor U1665 (N_1665,N_1272,N_1391);
and U1666 (N_1666,N_1148,N_1214);
and U1667 (N_1667,N_1373,N_1135);
nor U1668 (N_1668,N_1056,N_1143);
xnor U1669 (N_1669,N_1064,N_1428);
or U1670 (N_1670,N_1209,N_1318);
or U1671 (N_1671,N_1112,N_1393);
and U1672 (N_1672,N_1337,N_1130);
or U1673 (N_1673,N_1165,N_1489);
or U1674 (N_1674,N_1371,N_1423);
or U1675 (N_1675,N_1090,N_1290);
xor U1676 (N_1676,N_1157,N_1344);
or U1677 (N_1677,N_1001,N_1432);
and U1678 (N_1678,N_1308,N_1260);
or U1679 (N_1679,N_1078,N_1399);
or U1680 (N_1680,N_1292,N_1269);
and U1681 (N_1681,N_1422,N_1491);
nand U1682 (N_1682,N_1198,N_1244);
nor U1683 (N_1683,N_1252,N_1481);
nor U1684 (N_1684,N_1043,N_1086);
nor U1685 (N_1685,N_1154,N_1317);
nor U1686 (N_1686,N_1465,N_1394);
nor U1687 (N_1687,N_1127,N_1136);
and U1688 (N_1688,N_1052,N_1293);
and U1689 (N_1689,N_1190,N_1206);
nand U1690 (N_1690,N_1194,N_1250);
xor U1691 (N_1691,N_1089,N_1188);
nand U1692 (N_1692,N_1238,N_1187);
and U1693 (N_1693,N_1271,N_1448);
nor U1694 (N_1694,N_1418,N_1008);
xor U1695 (N_1695,N_1003,N_1083);
xor U1696 (N_1696,N_1213,N_1492);
and U1697 (N_1697,N_1230,N_1452);
nor U1698 (N_1698,N_1220,N_1121);
xor U1699 (N_1699,N_1288,N_1347);
nand U1700 (N_1700,N_1355,N_1240);
xor U1701 (N_1701,N_1469,N_1298);
or U1702 (N_1702,N_1479,N_1125);
nor U1703 (N_1703,N_1365,N_1352);
or U1704 (N_1704,N_1475,N_1286);
and U1705 (N_1705,N_1401,N_1038);
or U1706 (N_1706,N_1283,N_1405);
nand U1707 (N_1707,N_1319,N_1131);
or U1708 (N_1708,N_1361,N_1235);
xor U1709 (N_1709,N_1445,N_1372);
xor U1710 (N_1710,N_1378,N_1237);
and U1711 (N_1711,N_1341,N_1102);
nor U1712 (N_1712,N_1281,N_1369);
xor U1713 (N_1713,N_1199,N_1455);
xor U1714 (N_1714,N_1339,N_1367);
xnor U1715 (N_1715,N_1036,N_1002);
or U1716 (N_1716,N_1439,N_1366);
xor U1717 (N_1717,N_1424,N_1307);
and U1718 (N_1718,N_1497,N_1027);
xor U1719 (N_1719,N_1133,N_1182);
nor U1720 (N_1720,N_1129,N_1028);
or U1721 (N_1721,N_1146,N_1495);
xor U1722 (N_1722,N_1169,N_1349);
nand U1723 (N_1723,N_1223,N_1380);
nor U1724 (N_1724,N_1434,N_1051);
and U1725 (N_1725,N_1094,N_1353);
and U1726 (N_1726,N_1338,N_1443);
or U1727 (N_1727,N_1119,N_1303);
xnor U1728 (N_1728,N_1476,N_1386);
nor U1729 (N_1729,N_1205,N_1453);
xor U1730 (N_1730,N_1301,N_1041);
and U1731 (N_1731,N_1277,N_1383);
xor U1732 (N_1732,N_1196,N_1013);
nor U1733 (N_1733,N_1012,N_1171);
nand U1734 (N_1734,N_1097,N_1158);
nand U1735 (N_1735,N_1185,N_1404);
nand U1736 (N_1736,N_1201,N_1087);
xnor U1737 (N_1737,N_1096,N_1330);
and U1738 (N_1738,N_1493,N_1398);
or U1739 (N_1739,N_1413,N_1147);
and U1740 (N_1740,N_1270,N_1467);
nor U1741 (N_1741,N_1275,N_1153);
xnor U1742 (N_1742,N_1343,N_1266);
nand U1743 (N_1743,N_1315,N_1304);
or U1744 (N_1744,N_1456,N_1048);
xor U1745 (N_1745,N_1175,N_1184);
and U1746 (N_1746,N_1342,N_1312);
and U1747 (N_1747,N_1137,N_1134);
nor U1748 (N_1748,N_1245,N_1211);
xor U1749 (N_1749,N_1253,N_1329);
nor U1750 (N_1750,N_1142,N_1139);
xor U1751 (N_1751,N_1183,N_1037);
and U1752 (N_1752,N_1359,N_1055);
xnor U1753 (N_1753,N_1169,N_1235);
nand U1754 (N_1754,N_1118,N_1328);
or U1755 (N_1755,N_1170,N_1185);
nor U1756 (N_1756,N_1062,N_1180);
and U1757 (N_1757,N_1491,N_1257);
or U1758 (N_1758,N_1345,N_1031);
nor U1759 (N_1759,N_1276,N_1174);
nor U1760 (N_1760,N_1099,N_1416);
nor U1761 (N_1761,N_1374,N_1265);
nand U1762 (N_1762,N_1171,N_1275);
or U1763 (N_1763,N_1338,N_1161);
nand U1764 (N_1764,N_1314,N_1333);
xor U1765 (N_1765,N_1270,N_1360);
or U1766 (N_1766,N_1114,N_1112);
nand U1767 (N_1767,N_1011,N_1404);
nor U1768 (N_1768,N_1177,N_1159);
xnor U1769 (N_1769,N_1094,N_1051);
nand U1770 (N_1770,N_1133,N_1016);
xor U1771 (N_1771,N_1289,N_1219);
and U1772 (N_1772,N_1211,N_1005);
nor U1773 (N_1773,N_1121,N_1442);
xor U1774 (N_1774,N_1174,N_1293);
nor U1775 (N_1775,N_1024,N_1017);
nor U1776 (N_1776,N_1134,N_1437);
or U1777 (N_1777,N_1133,N_1024);
nand U1778 (N_1778,N_1267,N_1352);
or U1779 (N_1779,N_1274,N_1308);
nor U1780 (N_1780,N_1308,N_1250);
nor U1781 (N_1781,N_1045,N_1246);
nand U1782 (N_1782,N_1207,N_1477);
nand U1783 (N_1783,N_1317,N_1361);
nand U1784 (N_1784,N_1351,N_1396);
or U1785 (N_1785,N_1398,N_1391);
and U1786 (N_1786,N_1366,N_1378);
nand U1787 (N_1787,N_1440,N_1090);
nand U1788 (N_1788,N_1068,N_1207);
or U1789 (N_1789,N_1155,N_1146);
and U1790 (N_1790,N_1048,N_1187);
and U1791 (N_1791,N_1269,N_1393);
nor U1792 (N_1792,N_1174,N_1038);
or U1793 (N_1793,N_1409,N_1230);
xor U1794 (N_1794,N_1284,N_1499);
xnor U1795 (N_1795,N_1433,N_1050);
and U1796 (N_1796,N_1316,N_1381);
or U1797 (N_1797,N_1405,N_1399);
xnor U1798 (N_1798,N_1057,N_1338);
nor U1799 (N_1799,N_1145,N_1236);
and U1800 (N_1800,N_1255,N_1104);
or U1801 (N_1801,N_1474,N_1356);
nand U1802 (N_1802,N_1343,N_1253);
nor U1803 (N_1803,N_1317,N_1302);
or U1804 (N_1804,N_1209,N_1139);
and U1805 (N_1805,N_1354,N_1059);
or U1806 (N_1806,N_1115,N_1289);
nor U1807 (N_1807,N_1218,N_1362);
nand U1808 (N_1808,N_1119,N_1475);
and U1809 (N_1809,N_1292,N_1473);
and U1810 (N_1810,N_1399,N_1229);
nor U1811 (N_1811,N_1054,N_1044);
and U1812 (N_1812,N_1216,N_1419);
and U1813 (N_1813,N_1128,N_1346);
or U1814 (N_1814,N_1081,N_1459);
or U1815 (N_1815,N_1459,N_1020);
and U1816 (N_1816,N_1051,N_1107);
and U1817 (N_1817,N_1157,N_1094);
nor U1818 (N_1818,N_1215,N_1478);
or U1819 (N_1819,N_1096,N_1231);
nor U1820 (N_1820,N_1204,N_1068);
and U1821 (N_1821,N_1240,N_1065);
nor U1822 (N_1822,N_1476,N_1144);
nor U1823 (N_1823,N_1112,N_1315);
or U1824 (N_1824,N_1432,N_1095);
nand U1825 (N_1825,N_1204,N_1285);
and U1826 (N_1826,N_1045,N_1499);
or U1827 (N_1827,N_1082,N_1352);
nor U1828 (N_1828,N_1054,N_1092);
or U1829 (N_1829,N_1136,N_1252);
nand U1830 (N_1830,N_1160,N_1211);
nor U1831 (N_1831,N_1135,N_1242);
nand U1832 (N_1832,N_1286,N_1231);
xnor U1833 (N_1833,N_1058,N_1417);
and U1834 (N_1834,N_1351,N_1389);
xnor U1835 (N_1835,N_1149,N_1224);
and U1836 (N_1836,N_1077,N_1184);
nand U1837 (N_1837,N_1159,N_1334);
nand U1838 (N_1838,N_1244,N_1408);
nand U1839 (N_1839,N_1392,N_1020);
and U1840 (N_1840,N_1467,N_1230);
or U1841 (N_1841,N_1151,N_1167);
nand U1842 (N_1842,N_1187,N_1434);
nor U1843 (N_1843,N_1039,N_1449);
xnor U1844 (N_1844,N_1282,N_1301);
or U1845 (N_1845,N_1294,N_1463);
xor U1846 (N_1846,N_1037,N_1208);
xor U1847 (N_1847,N_1310,N_1498);
nand U1848 (N_1848,N_1464,N_1228);
nand U1849 (N_1849,N_1196,N_1256);
and U1850 (N_1850,N_1006,N_1434);
xnor U1851 (N_1851,N_1189,N_1308);
and U1852 (N_1852,N_1383,N_1230);
nand U1853 (N_1853,N_1044,N_1082);
nor U1854 (N_1854,N_1042,N_1371);
nand U1855 (N_1855,N_1281,N_1253);
nor U1856 (N_1856,N_1377,N_1158);
and U1857 (N_1857,N_1329,N_1277);
and U1858 (N_1858,N_1381,N_1444);
or U1859 (N_1859,N_1319,N_1360);
or U1860 (N_1860,N_1328,N_1482);
or U1861 (N_1861,N_1482,N_1038);
xor U1862 (N_1862,N_1149,N_1106);
nor U1863 (N_1863,N_1313,N_1391);
or U1864 (N_1864,N_1363,N_1306);
xor U1865 (N_1865,N_1292,N_1291);
nand U1866 (N_1866,N_1231,N_1356);
xnor U1867 (N_1867,N_1222,N_1143);
nand U1868 (N_1868,N_1159,N_1292);
or U1869 (N_1869,N_1459,N_1123);
xnor U1870 (N_1870,N_1362,N_1402);
nand U1871 (N_1871,N_1496,N_1373);
xor U1872 (N_1872,N_1137,N_1029);
and U1873 (N_1873,N_1323,N_1419);
xor U1874 (N_1874,N_1494,N_1176);
nor U1875 (N_1875,N_1076,N_1253);
xor U1876 (N_1876,N_1443,N_1179);
or U1877 (N_1877,N_1118,N_1337);
nor U1878 (N_1878,N_1414,N_1192);
nor U1879 (N_1879,N_1297,N_1188);
or U1880 (N_1880,N_1147,N_1298);
or U1881 (N_1881,N_1200,N_1456);
or U1882 (N_1882,N_1121,N_1044);
nor U1883 (N_1883,N_1258,N_1488);
nand U1884 (N_1884,N_1269,N_1209);
and U1885 (N_1885,N_1124,N_1183);
nand U1886 (N_1886,N_1329,N_1046);
xnor U1887 (N_1887,N_1100,N_1483);
or U1888 (N_1888,N_1065,N_1491);
or U1889 (N_1889,N_1354,N_1383);
or U1890 (N_1890,N_1023,N_1475);
xor U1891 (N_1891,N_1117,N_1094);
or U1892 (N_1892,N_1319,N_1262);
and U1893 (N_1893,N_1025,N_1203);
nor U1894 (N_1894,N_1111,N_1286);
or U1895 (N_1895,N_1426,N_1020);
nor U1896 (N_1896,N_1407,N_1117);
and U1897 (N_1897,N_1089,N_1176);
nand U1898 (N_1898,N_1229,N_1081);
xor U1899 (N_1899,N_1284,N_1113);
and U1900 (N_1900,N_1059,N_1208);
and U1901 (N_1901,N_1064,N_1181);
nor U1902 (N_1902,N_1210,N_1354);
or U1903 (N_1903,N_1149,N_1277);
and U1904 (N_1904,N_1478,N_1301);
xor U1905 (N_1905,N_1194,N_1117);
xor U1906 (N_1906,N_1402,N_1221);
xnor U1907 (N_1907,N_1034,N_1174);
xnor U1908 (N_1908,N_1210,N_1323);
nor U1909 (N_1909,N_1487,N_1225);
and U1910 (N_1910,N_1270,N_1067);
and U1911 (N_1911,N_1356,N_1055);
and U1912 (N_1912,N_1290,N_1048);
and U1913 (N_1913,N_1115,N_1439);
and U1914 (N_1914,N_1295,N_1425);
or U1915 (N_1915,N_1034,N_1364);
xor U1916 (N_1916,N_1197,N_1362);
or U1917 (N_1917,N_1113,N_1238);
nand U1918 (N_1918,N_1152,N_1176);
and U1919 (N_1919,N_1132,N_1170);
xnor U1920 (N_1920,N_1089,N_1275);
xor U1921 (N_1921,N_1166,N_1213);
nand U1922 (N_1922,N_1410,N_1036);
nand U1923 (N_1923,N_1196,N_1354);
nand U1924 (N_1924,N_1333,N_1250);
nor U1925 (N_1925,N_1267,N_1043);
and U1926 (N_1926,N_1124,N_1369);
or U1927 (N_1927,N_1246,N_1134);
or U1928 (N_1928,N_1160,N_1188);
or U1929 (N_1929,N_1111,N_1237);
nor U1930 (N_1930,N_1242,N_1234);
and U1931 (N_1931,N_1210,N_1129);
xnor U1932 (N_1932,N_1209,N_1357);
nor U1933 (N_1933,N_1327,N_1499);
and U1934 (N_1934,N_1439,N_1349);
or U1935 (N_1935,N_1189,N_1191);
nand U1936 (N_1936,N_1185,N_1225);
nand U1937 (N_1937,N_1275,N_1036);
nand U1938 (N_1938,N_1045,N_1113);
nand U1939 (N_1939,N_1066,N_1433);
xor U1940 (N_1940,N_1190,N_1184);
nor U1941 (N_1941,N_1108,N_1262);
xnor U1942 (N_1942,N_1166,N_1049);
nand U1943 (N_1943,N_1450,N_1232);
nor U1944 (N_1944,N_1393,N_1215);
xor U1945 (N_1945,N_1263,N_1138);
nor U1946 (N_1946,N_1255,N_1473);
xnor U1947 (N_1947,N_1167,N_1191);
or U1948 (N_1948,N_1379,N_1155);
or U1949 (N_1949,N_1077,N_1263);
nor U1950 (N_1950,N_1243,N_1412);
nor U1951 (N_1951,N_1156,N_1276);
nor U1952 (N_1952,N_1068,N_1334);
nor U1953 (N_1953,N_1390,N_1455);
nand U1954 (N_1954,N_1057,N_1376);
or U1955 (N_1955,N_1205,N_1227);
xnor U1956 (N_1956,N_1214,N_1410);
nand U1957 (N_1957,N_1388,N_1247);
xor U1958 (N_1958,N_1285,N_1449);
nand U1959 (N_1959,N_1378,N_1194);
nand U1960 (N_1960,N_1058,N_1138);
nand U1961 (N_1961,N_1099,N_1070);
and U1962 (N_1962,N_1049,N_1353);
and U1963 (N_1963,N_1194,N_1410);
and U1964 (N_1964,N_1108,N_1119);
nor U1965 (N_1965,N_1346,N_1392);
nor U1966 (N_1966,N_1106,N_1463);
nor U1967 (N_1967,N_1482,N_1086);
nor U1968 (N_1968,N_1211,N_1214);
nor U1969 (N_1969,N_1438,N_1427);
xor U1970 (N_1970,N_1034,N_1064);
or U1971 (N_1971,N_1309,N_1457);
xor U1972 (N_1972,N_1003,N_1076);
or U1973 (N_1973,N_1048,N_1405);
or U1974 (N_1974,N_1487,N_1108);
and U1975 (N_1975,N_1327,N_1125);
and U1976 (N_1976,N_1192,N_1234);
nand U1977 (N_1977,N_1059,N_1065);
xor U1978 (N_1978,N_1367,N_1356);
nor U1979 (N_1979,N_1366,N_1288);
nor U1980 (N_1980,N_1193,N_1367);
and U1981 (N_1981,N_1001,N_1459);
and U1982 (N_1982,N_1108,N_1274);
xnor U1983 (N_1983,N_1063,N_1196);
nor U1984 (N_1984,N_1048,N_1400);
or U1985 (N_1985,N_1243,N_1352);
nand U1986 (N_1986,N_1078,N_1384);
nand U1987 (N_1987,N_1425,N_1089);
nor U1988 (N_1988,N_1010,N_1456);
and U1989 (N_1989,N_1041,N_1129);
xor U1990 (N_1990,N_1234,N_1487);
nor U1991 (N_1991,N_1377,N_1476);
or U1992 (N_1992,N_1353,N_1437);
and U1993 (N_1993,N_1380,N_1016);
and U1994 (N_1994,N_1357,N_1435);
nand U1995 (N_1995,N_1319,N_1033);
xor U1996 (N_1996,N_1415,N_1363);
nand U1997 (N_1997,N_1047,N_1065);
nand U1998 (N_1998,N_1294,N_1117);
xnor U1999 (N_1999,N_1103,N_1016);
xor U2000 (N_2000,N_1730,N_1692);
nand U2001 (N_2001,N_1537,N_1626);
nand U2002 (N_2002,N_1829,N_1745);
xnor U2003 (N_2003,N_1785,N_1972);
or U2004 (N_2004,N_1546,N_1780);
nor U2005 (N_2005,N_1754,N_1635);
and U2006 (N_2006,N_1986,N_1932);
and U2007 (N_2007,N_1768,N_1636);
xnor U2008 (N_2008,N_1505,N_1755);
nand U2009 (N_2009,N_1543,N_1977);
nand U2010 (N_2010,N_1882,N_1989);
nor U2011 (N_2011,N_1616,N_1828);
nor U2012 (N_2012,N_1618,N_1840);
xnor U2013 (N_2013,N_1717,N_1594);
nor U2014 (N_2014,N_1883,N_1689);
nor U2015 (N_2015,N_1617,N_1819);
xor U2016 (N_2016,N_1707,N_1502);
xnor U2017 (N_2017,N_1836,N_1984);
or U2018 (N_2018,N_1578,N_1678);
xor U2019 (N_2019,N_1670,N_1593);
and U2020 (N_2020,N_1987,N_1838);
xnor U2021 (N_2021,N_1794,N_1753);
and U2022 (N_2022,N_1835,N_1807);
and U2023 (N_2023,N_1672,N_1607);
or U2024 (N_2024,N_1741,N_1605);
nor U2025 (N_2025,N_1500,N_1575);
or U2026 (N_2026,N_1936,N_1916);
or U2027 (N_2027,N_1708,N_1816);
nand U2028 (N_2028,N_1632,N_1731);
nor U2029 (N_2029,N_1899,N_1724);
and U2030 (N_2030,N_1948,N_1966);
and U2031 (N_2031,N_1850,N_1718);
nand U2032 (N_2032,N_1997,N_1530);
or U2033 (N_2033,N_1798,N_1778);
nor U2034 (N_2034,N_1845,N_1868);
or U2035 (N_2035,N_1705,N_1647);
xnor U2036 (N_2036,N_1784,N_1859);
xnor U2037 (N_2037,N_1957,N_1928);
nand U2038 (N_2038,N_1979,N_1676);
nand U2039 (N_2039,N_1574,N_1894);
nand U2040 (N_2040,N_1649,N_1969);
xor U2041 (N_2041,N_1914,N_1752);
xnor U2042 (N_2042,N_1934,N_1791);
xnor U2043 (N_2043,N_1517,N_1541);
nor U2044 (N_2044,N_1614,N_1803);
or U2045 (N_2045,N_1581,N_1657);
and U2046 (N_2046,N_1808,N_1540);
and U2047 (N_2047,N_1975,N_1521);
nor U2048 (N_2048,N_1596,N_1843);
and U2049 (N_2049,N_1786,N_1736);
nor U2050 (N_2050,N_1650,N_1851);
and U2051 (N_2051,N_1773,N_1527);
nor U2052 (N_2052,N_1503,N_1955);
and U2053 (N_2053,N_1652,N_1925);
and U2054 (N_2054,N_1766,N_1663);
or U2055 (N_2055,N_1522,N_1853);
and U2056 (N_2056,N_1841,N_1719);
xor U2057 (N_2057,N_1789,N_1613);
nand U2058 (N_2058,N_1556,N_1664);
and U2059 (N_2059,N_1974,N_1625);
nor U2060 (N_2060,N_1712,N_1589);
xor U2061 (N_2061,N_1886,N_1720);
nand U2062 (N_2062,N_1601,N_1747);
nor U2063 (N_2063,N_1535,N_1611);
and U2064 (N_2064,N_1976,N_1849);
and U2065 (N_2065,N_1529,N_1938);
xnor U2066 (N_2066,N_1864,N_1999);
xor U2067 (N_2067,N_1912,N_1861);
nand U2068 (N_2068,N_1534,N_1658);
nand U2069 (N_2069,N_1628,N_1603);
and U2070 (N_2070,N_1597,N_1715);
nor U2071 (N_2071,N_1901,N_1639);
and U2072 (N_2072,N_1690,N_1548);
xor U2073 (N_2073,N_1551,N_1743);
and U2074 (N_2074,N_1587,N_1895);
nor U2075 (N_2075,N_1532,N_1797);
and U2076 (N_2076,N_1848,N_1967);
or U2077 (N_2077,N_1508,N_1930);
and U2078 (N_2078,N_1509,N_1586);
nand U2079 (N_2079,N_1683,N_1788);
and U2080 (N_2080,N_1620,N_1760);
nand U2081 (N_2081,N_1837,N_1926);
nor U2082 (N_2082,N_1561,N_1777);
xor U2083 (N_2083,N_1641,N_1973);
and U2084 (N_2084,N_1876,N_1923);
or U2085 (N_2085,N_1640,N_1550);
and U2086 (N_2086,N_1834,N_1854);
nor U2087 (N_2087,N_1567,N_1554);
nor U2088 (N_2088,N_1629,N_1713);
or U2089 (N_2089,N_1638,N_1863);
nor U2090 (N_2090,N_1698,N_1951);
or U2091 (N_2091,N_1729,N_1891);
xnor U2092 (N_2092,N_1526,N_1949);
nand U2093 (N_2093,N_1893,N_1885);
and U2094 (N_2094,N_1790,N_1699);
and U2095 (N_2095,N_1523,N_1542);
xor U2096 (N_2096,N_1918,N_1959);
nor U2097 (N_2097,N_1595,N_1890);
nand U2098 (N_2098,N_1519,N_1598);
and U2099 (N_2099,N_1566,N_1547);
nand U2100 (N_2100,N_1824,N_1702);
and U2101 (N_2101,N_1763,N_1742);
xor U2102 (N_2102,N_1884,N_1878);
and U2103 (N_2103,N_1947,N_1538);
xnor U2104 (N_2104,N_1700,N_1668);
and U2105 (N_2105,N_1814,N_1818);
xnor U2106 (N_2106,N_1782,N_1653);
nor U2107 (N_2107,N_1703,N_1776);
or U2108 (N_2108,N_1659,N_1994);
and U2109 (N_2109,N_1911,N_1552);
xnor U2110 (N_2110,N_1706,N_1651);
nor U2111 (N_2111,N_1697,N_1813);
xnor U2112 (N_2112,N_1666,N_1665);
and U2113 (N_2113,N_1604,N_1919);
or U2114 (N_2114,N_1684,N_1902);
or U2115 (N_2115,N_1832,N_1783);
or U2116 (N_2116,N_1988,N_1802);
nor U2117 (N_2117,N_1946,N_1875);
and U2118 (N_2118,N_1671,N_1528);
nand U2119 (N_2119,N_1998,N_1565);
xnor U2120 (N_2120,N_1961,N_1648);
or U2121 (N_2121,N_1779,N_1661);
nand U2122 (N_2122,N_1759,N_1906);
or U2123 (N_2123,N_1660,N_1558);
or U2124 (N_2124,N_1709,N_1950);
and U2125 (N_2125,N_1583,N_1991);
and U2126 (N_2126,N_1515,N_1758);
xnor U2127 (N_2127,N_1872,N_1563);
xnor U2128 (N_2128,N_1960,N_1799);
or U2129 (N_2129,N_1680,N_1619);
nand U2130 (N_2130,N_1761,N_1996);
and U2131 (N_2131,N_1920,N_1858);
or U2132 (N_2132,N_1701,N_1591);
nor U2133 (N_2133,N_1856,N_1956);
xor U2134 (N_2134,N_1501,N_1811);
or U2135 (N_2135,N_1734,N_1900);
and U2136 (N_2136,N_1545,N_1716);
or U2137 (N_2137,N_1531,N_1965);
nor U2138 (N_2138,N_1922,N_1602);
xor U2139 (N_2139,N_1681,N_1822);
or U2140 (N_2140,N_1917,N_1504);
nand U2141 (N_2141,N_1564,N_1931);
nand U2142 (N_2142,N_1744,N_1568);
nor U2143 (N_2143,N_1874,N_1870);
nand U2144 (N_2144,N_1656,N_1963);
or U2145 (N_2145,N_1599,N_1748);
nand U2146 (N_2146,N_1855,N_1821);
and U2147 (N_2147,N_1622,N_1970);
and U2148 (N_2148,N_1944,N_1630);
nor U2149 (N_2149,N_1524,N_1817);
nand U2150 (N_2150,N_1775,N_1770);
and U2151 (N_2151,N_1533,N_1518);
nor U2152 (N_2152,N_1993,N_1806);
or U2153 (N_2153,N_1881,N_1787);
nor U2154 (N_2154,N_1512,N_1728);
xnor U2155 (N_2155,N_1710,N_1954);
or U2156 (N_2156,N_1711,N_1631);
or U2157 (N_2157,N_1990,N_1615);
xor U2158 (N_2158,N_1507,N_1769);
and U2159 (N_2159,N_1839,N_1643);
xor U2160 (N_2160,N_1726,N_1637);
nor U2161 (N_2161,N_1588,N_1669);
nor U2162 (N_2162,N_1933,N_1940);
or U2163 (N_2163,N_1582,N_1847);
xor U2164 (N_2164,N_1952,N_1609);
and U2165 (N_2165,N_1722,N_1655);
xor U2166 (N_2166,N_1675,N_1750);
or U2167 (N_2167,N_1871,N_1725);
or U2168 (N_2168,N_1907,N_1756);
and U2169 (N_2169,N_1516,N_1913);
nand U2170 (N_2170,N_1600,N_1572);
nand U2171 (N_2171,N_1737,N_1823);
xor U2172 (N_2172,N_1555,N_1585);
and U2173 (N_2173,N_1682,N_1879);
nand U2174 (N_2174,N_1800,N_1897);
nor U2175 (N_2175,N_1765,N_1714);
nor U2176 (N_2176,N_1506,N_1688);
nor U2177 (N_2177,N_1796,N_1757);
and U2178 (N_2178,N_1608,N_1852);
nand U2179 (N_2179,N_1921,N_1842);
and U2180 (N_2180,N_1514,N_1945);
and U2181 (N_2181,N_1612,N_1536);
nand U2182 (N_2182,N_1580,N_1621);
or U2183 (N_2183,N_1831,N_1721);
and U2184 (N_2184,N_1764,N_1887);
nor U2185 (N_2185,N_1584,N_1723);
nand U2186 (N_2186,N_1982,N_1792);
xnor U2187 (N_2187,N_1667,N_1746);
nor U2188 (N_2188,N_1691,N_1857);
xnor U2189 (N_2189,N_1772,N_1634);
and U2190 (N_2190,N_1910,N_1929);
or U2191 (N_2191,N_1781,N_1846);
xnor U2192 (N_2192,N_1510,N_1978);
xnor U2193 (N_2193,N_1696,N_1826);
nand U2194 (N_2194,N_1579,N_1962);
or U2195 (N_2195,N_1908,N_1662);
nor U2196 (N_2196,N_1801,N_1877);
nor U2197 (N_2197,N_1873,N_1880);
and U2198 (N_2198,N_1771,N_1869);
nand U2199 (N_2199,N_1898,N_1915);
nand U2200 (N_2200,N_1577,N_1860);
or U2201 (N_2201,N_1903,N_1767);
nor U2202 (N_2202,N_1610,N_1694);
xnor U2203 (N_2203,N_1693,N_1624);
nand U2204 (N_2204,N_1679,N_1673);
and U2205 (N_2205,N_1642,N_1815);
or U2206 (N_2206,N_1953,N_1654);
and U2207 (N_2207,N_1888,N_1985);
or U2208 (N_2208,N_1939,N_1825);
nor U2209 (N_2209,N_1844,N_1943);
or U2210 (N_2210,N_1562,N_1809);
nor U2211 (N_2211,N_1549,N_1576);
nand U2212 (N_2212,N_1751,N_1804);
xnor U2213 (N_2213,N_1889,N_1971);
and U2214 (N_2214,N_1674,N_1830);
or U2215 (N_2215,N_1559,N_1590);
and U2216 (N_2216,N_1866,N_1958);
xnor U2217 (N_2217,N_1738,N_1909);
nor U2218 (N_2218,N_1732,N_1827);
or U2219 (N_2219,N_1606,N_1941);
and U2220 (N_2220,N_1513,N_1644);
or U2221 (N_2221,N_1904,N_1695);
nand U2222 (N_2222,N_1569,N_1525);
nand U2223 (N_2223,N_1981,N_1740);
or U2224 (N_2224,N_1570,N_1520);
xor U2225 (N_2225,N_1685,N_1646);
nand U2226 (N_2226,N_1749,N_1937);
or U2227 (N_2227,N_1935,N_1686);
and U2228 (N_2228,N_1735,N_1964);
nor U2229 (N_2229,N_1795,N_1511);
nor U2230 (N_2230,N_1805,N_1539);
nor U2231 (N_2231,N_1905,N_1557);
nor U2232 (N_2232,N_1992,N_1833);
or U2233 (N_2233,N_1896,N_1704);
xnor U2234 (N_2234,N_1762,N_1793);
or U2235 (N_2235,N_1623,N_1995);
nand U2236 (N_2236,N_1820,N_1573);
nand U2237 (N_2237,N_1553,N_1812);
xor U2238 (N_2238,N_1733,N_1592);
and U2239 (N_2239,N_1677,N_1560);
or U2240 (N_2240,N_1862,N_1687);
xnor U2241 (N_2241,N_1727,N_1942);
or U2242 (N_2242,N_1865,N_1892);
xor U2243 (N_2243,N_1645,N_1774);
xor U2244 (N_2244,N_1739,N_1980);
and U2245 (N_2245,N_1968,N_1927);
or U2246 (N_2246,N_1924,N_1627);
nand U2247 (N_2247,N_1983,N_1544);
nor U2248 (N_2248,N_1571,N_1633);
and U2249 (N_2249,N_1810,N_1867);
nand U2250 (N_2250,N_1626,N_1842);
nand U2251 (N_2251,N_1943,N_1593);
nand U2252 (N_2252,N_1581,N_1826);
nor U2253 (N_2253,N_1996,N_1523);
or U2254 (N_2254,N_1563,N_1552);
or U2255 (N_2255,N_1923,N_1807);
or U2256 (N_2256,N_1590,N_1813);
nor U2257 (N_2257,N_1611,N_1603);
xnor U2258 (N_2258,N_1922,N_1817);
nand U2259 (N_2259,N_1627,N_1661);
or U2260 (N_2260,N_1843,N_1963);
nor U2261 (N_2261,N_1711,N_1968);
or U2262 (N_2262,N_1662,N_1898);
nand U2263 (N_2263,N_1709,N_1852);
and U2264 (N_2264,N_1939,N_1771);
nand U2265 (N_2265,N_1629,N_1760);
nand U2266 (N_2266,N_1678,N_1908);
nor U2267 (N_2267,N_1687,N_1708);
nor U2268 (N_2268,N_1985,N_1940);
or U2269 (N_2269,N_1661,N_1566);
or U2270 (N_2270,N_1856,N_1536);
and U2271 (N_2271,N_1921,N_1784);
and U2272 (N_2272,N_1689,N_1639);
xor U2273 (N_2273,N_1724,N_1547);
nand U2274 (N_2274,N_1934,N_1502);
nor U2275 (N_2275,N_1827,N_1961);
xnor U2276 (N_2276,N_1842,N_1663);
nor U2277 (N_2277,N_1648,N_1787);
xnor U2278 (N_2278,N_1584,N_1792);
nor U2279 (N_2279,N_1514,N_1520);
xor U2280 (N_2280,N_1998,N_1884);
nor U2281 (N_2281,N_1984,N_1794);
nand U2282 (N_2282,N_1590,N_1687);
xnor U2283 (N_2283,N_1736,N_1841);
nand U2284 (N_2284,N_1628,N_1641);
xor U2285 (N_2285,N_1950,N_1686);
nor U2286 (N_2286,N_1655,N_1846);
or U2287 (N_2287,N_1627,N_1721);
xnor U2288 (N_2288,N_1915,N_1733);
nor U2289 (N_2289,N_1555,N_1513);
and U2290 (N_2290,N_1736,N_1862);
nand U2291 (N_2291,N_1584,N_1853);
and U2292 (N_2292,N_1736,N_1800);
nand U2293 (N_2293,N_1742,N_1827);
nor U2294 (N_2294,N_1831,N_1962);
nand U2295 (N_2295,N_1570,N_1771);
nor U2296 (N_2296,N_1618,N_1944);
or U2297 (N_2297,N_1927,N_1828);
xor U2298 (N_2298,N_1562,N_1966);
nand U2299 (N_2299,N_1996,N_1669);
and U2300 (N_2300,N_1976,N_1776);
nand U2301 (N_2301,N_1653,N_1910);
nor U2302 (N_2302,N_1720,N_1975);
or U2303 (N_2303,N_1516,N_1519);
nand U2304 (N_2304,N_1568,N_1857);
or U2305 (N_2305,N_1839,N_1601);
nor U2306 (N_2306,N_1642,N_1665);
or U2307 (N_2307,N_1745,N_1652);
xnor U2308 (N_2308,N_1938,N_1818);
nor U2309 (N_2309,N_1671,N_1714);
nand U2310 (N_2310,N_1837,N_1714);
and U2311 (N_2311,N_1564,N_1603);
xor U2312 (N_2312,N_1642,N_1760);
xnor U2313 (N_2313,N_1794,N_1895);
or U2314 (N_2314,N_1953,N_1571);
xnor U2315 (N_2315,N_1560,N_1517);
xnor U2316 (N_2316,N_1658,N_1765);
nor U2317 (N_2317,N_1816,N_1560);
and U2318 (N_2318,N_1816,N_1577);
xnor U2319 (N_2319,N_1756,N_1590);
and U2320 (N_2320,N_1674,N_1914);
nor U2321 (N_2321,N_1936,N_1834);
nor U2322 (N_2322,N_1528,N_1935);
xnor U2323 (N_2323,N_1956,N_1809);
and U2324 (N_2324,N_1741,N_1638);
xnor U2325 (N_2325,N_1506,N_1992);
nand U2326 (N_2326,N_1740,N_1825);
nand U2327 (N_2327,N_1984,N_1863);
and U2328 (N_2328,N_1870,N_1535);
and U2329 (N_2329,N_1902,N_1891);
and U2330 (N_2330,N_1600,N_1905);
nor U2331 (N_2331,N_1562,N_1941);
and U2332 (N_2332,N_1549,N_1507);
nand U2333 (N_2333,N_1836,N_1849);
nand U2334 (N_2334,N_1706,N_1621);
nand U2335 (N_2335,N_1705,N_1514);
nor U2336 (N_2336,N_1585,N_1989);
or U2337 (N_2337,N_1764,N_1526);
nor U2338 (N_2338,N_1703,N_1925);
nor U2339 (N_2339,N_1624,N_1696);
or U2340 (N_2340,N_1721,N_1728);
and U2341 (N_2341,N_1509,N_1807);
and U2342 (N_2342,N_1844,N_1500);
nor U2343 (N_2343,N_1669,N_1727);
and U2344 (N_2344,N_1772,N_1776);
nor U2345 (N_2345,N_1764,N_1683);
nand U2346 (N_2346,N_1790,N_1551);
or U2347 (N_2347,N_1628,N_1507);
nand U2348 (N_2348,N_1724,N_1973);
nor U2349 (N_2349,N_1584,N_1562);
nor U2350 (N_2350,N_1961,N_1776);
xor U2351 (N_2351,N_1980,N_1622);
xnor U2352 (N_2352,N_1653,N_1941);
or U2353 (N_2353,N_1961,N_1519);
and U2354 (N_2354,N_1606,N_1626);
xor U2355 (N_2355,N_1530,N_1503);
nand U2356 (N_2356,N_1840,N_1795);
nand U2357 (N_2357,N_1834,N_1951);
and U2358 (N_2358,N_1990,N_1927);
xor U2359 (N_2359,N_1747,N_1834);
nor U2360 (N_2360,N_1690,N_1790);
nor U2361 (N_2361,N_1996,N_1527);
nand U2362 (N_2362,N_1593,N_1862);
nor U2363 (N_2363,N_1984,N_1675);
and U2364 (N_2364,N_1808,N_1765);
xor U2365 (N_2365,N_1767,N_1861);
or U2366 (N_2366,N_1756,N_1823);
nor U2367 (N_2367,N_1800,N_1602);
nand U2368 (N_2368,N_1933,N_1599);
and U2369 (N_2369,N_1578,N_1704);
nor U2370 (N_2370,N_1823,N_1888);
nand U2371 (N_2371,N_1828,N_1728);
xor U2372 (N_2372,N_1624,N_1564);
nor U2373 (N_2373,N_1683,N_1655);
nor U2374 (N_2374,N_1663,N_1532);
nor U2375 (N_2375,N_1900,N_1530);
and U2376 (N_2376,N_1709,N_1725);
nor U2377 (N_2377,N_1789,N_1631);
nor U2378 (N_2378,N_1761,N_1791);
and U2379 (N_2379,N_1777,N_1759);
nor U2380 (N_2380,N_1933,N_1569);
nor U2381 (N_2381,N_1940,N_1575);
xor U2382 (N_2382,N_1547,N_1731);
nor U2383 (N_2383,N_1646,N_1622);
or U2384 (N_2384,N_1767,N_1868);
or U2385 (N_2385,N_1762,N_1961);
and U2386 (N_2386,N_1776,N_1931);
xnor U2387 (N_2387,N_1708,N_1921);
nand U2388 (N_2388,N_1844,N_1549);
and U2389 (N_2389,N_1855,N_1897);
and U2390 (N_2390,N_1521,N_1856);
nor U2391 (N_2391,N_1958,N_1966);
and U2392 (N_2392,N_1786,N_1580);
nand U2393 (N_2393,N_1718,N_1805);
xor U2394 (N_2394,N_1822,N_1939);
or U2395 (N_2395,N_1761,N_1860);
nand U2396 (N_2396,N_1682,N_1762);
nor U2397 (N_2397,N_1602,N_1690);
and U2398 (N_2398,N_1597,N_1525);
nand U2399 (N_2399,N_1961,N_1721);
and U2400 (N_2400,N_1707,N_1913);
nor U2401 (N_2401,N_1848,N_1993);
and U2402 (N_2402,N_1926,N_1828);
xnor U2403 (N_2403,N_1980,N_1858);
nor U2404 (N_2404,N_1591,N_1547);
nand U2405 (N_2405,N_1797,N_1512);
or U2406 (N_2406,N_1774,N_1827);
nand U2407 (N_2407,N_1807,N_1695);
and U2408 (N_2408,N_1987,N_1527);
xnor U2409 (N_2409,N_1941,N_1764);
nor U2410 (N_2410,N_1722,N_1898);
nand U2411 (N_2411,N_1782,N_1849);
nand U2412 (N_2412,N_1731,N_1613);
xnor U2413 (N_2413,N_1606,N_1830);
nor U2414 (N_2414,N_1603,N_1613);
nor U2415 (N_2415,N_1957,N_1860);
and U2416 (N_2416,N_1761,N_1526);
nor U2417 (N_2417,N_1814,N_1800);
nor U2418 (N_2418,N_1784,N_1846);
nand U2419 (N_2419,N_1753,N_1632);
or U2420 (N_2420,N_1578,N_1705);
xor U2421 (N_2421,N_1684,N_1648);
or U2422 (N_2422,N_1938,N_1948);
nor U2423 (N_2423,N_1694,N_1706);
and U2424 (N_2424,N_1917,N_1967);
or U2425 (N_2425,N_1971,N_1778);
xor U2426 (N_2426,N_1909,N_1985);
xor U2427 (N_2427,N_1896,N_1681);
nand U2428 (N_2428,N_1568,N_1878);
and U2429 (N_2429,N_1607,N_1949);
nor U2430 (N_2430,N_1812,N_1630);
nor U2431 (N_2431,N_1962,N_1804);
xor U2432 (N_2432,N_1640,N_1954);
xnor U2433 (N_2433,N_1608,N_1940);
nor U2434 (N_2434,N_1843,N_1780);
and U2435 (N_2435,N_1888,N_1603);
nand U2436 (N_2436,N_1693,N_1679);
or U2437 (N_2437,N_1561,N_1799);
or U2438 (N_2438,N_1806,N_1991);
nand U2439 (N_2439,N_1621,N_1906);
and U2440 (N_2440,N_1819,N_1642);
nand U2441 (N_2441,N_1665,N_1699);
nand U2442 (N_2442,N_1841,N_1981);
nor U2443 (N_2443,N_1631,N_1527);
and U2444 (N_2444,N_1811,N_1665);
nor U2445 (N_2445,N_1885,N_1704);
xnor U2446 (N_2446,N_1690,N_1536);
or U2447 (N_2447,N_1647,N_1909);
xnor U2448 (N_2448,N_1692,N_1643);
and U2449 (N_2449,N_1739,N_1766);
nor U2450 (N_2450,N_1624,N_1827);
nor U2451 (N_2451,N_1592,N_1789);
xor U2452 (N_2452,N_1516,N_1925);
or U2453 (N_2453,N_1540,N_1736);
nor U2454 (N_2454,N_1913,N_1538);
and U2455 (N_2455,N_1742,N_1800);
or U2456 (N_2456,N_1707,N_1965);
nand U2457 (N_2457,N_1918,N_1642);
nor U2458 (N_2458,N_1834,N_1568);
xor U2459 (N_2459,N_1788,N_1718);
nor U2460 (N_2460,N_1879,N_1561);
or U2461 (N_2461,N_1693,N_1694);
or U2462 (N_2462,N_1780,N_1698);
nor U2463 (N_2463,N_1837,N_1959);
nand U2464 (N_2464,N_1551,N_1958);
nand U2465 (N_2465,N_1747,N_1941);
xnor U2466 (N_2466,N_1787,N_1804);
xnor U2467 (N_2467,N_1836,N_1733);
nand U2468 (N_2468,N_1512,N_1789);
or U2469 (N_2469,N_1511,N_1938);
nand U2470 (N_2470,N_1864,N_1764);
or U2471 (N_2471,N_1526,N_1653);
or U2472 (N_2472,N_1771,N_1729);
and U2473 (N_2473,N_1916,N_1950);
nand U2474 (N_2474,N_1677,N_1875);
and U2475 (N_2475,N_1868,N_1837);
nand U2476 (N_2476,N_1788,N_1797);
nand U2477 (N_2477,N_1896,N_1514);
and U2478 (N_2478,N_1722,N_1596);
and U2479 (N_2479,N_1612,N_1858);
nand U2480 (N_2480,N_1897,N_1976);
nand U2481 (N_2481,N_1807,N_1798);
or U2482 (N_2482,N_1678,N_1625);
and U2483 (N_2483,N_1990,N_1864);
nand U2484 (N_2484,N_1657,N_1950);
xor U2485 (N_2485,N_1675,N_1633);
and U2486 (N_2486,N_1651,N_1681);
or U2487 (N_2487,N_1706,N_1816);
xnor U2488 (N_2488,N_1892,N_1735);
nand U2489 (N_2489,N_1958,N_1732);
or U2490 (N_2490,N_1516,N_1948);
xnor U2491 (N_2491,N_1629,N_1718);
and U2492 (N_2492,N_1909,N_1778);
nor U2493 (N_2493,N_1562,N_1630);
nand U2494 (N_2494,N_1920,N_1708);
and U2495 (N_2495,N_1772,N_1611);
nand U2496 (N_2496,N_1666,N_1995);
and U2497 (N_2497,N_1567,N_1548);
and U2498 (N_2498,N_1735,N_1592);
and U2499 (N_2499,N_1740,N_1711);
nand U2500 (N_2500,N_2015,N_2009);
or U2501 (N_2501,N_2440,N_2164);
and U2502 (N_2502,N_2207,N_2161);
and U2503 (N_2503,N_2403,N_2071);
nand U2504 (N_2504,N_2464,N_2484);
and U2505 (N_2505,N_2360,N_2343);
nand U2506 (N_2506,N_2004,N_2355);
or U2507 (N_2507,N_2385,N_2014);
and U2508 (N_2508,N_2198,N_2177);
or U2509 (N_2509,N_2283,N_2433);
nor U2510 (N_2510,N_2390,N_2049);
or U2511 (N_2511,N_2087,N_2232);
nand U2512 (N_2512,N_2065,N_2341);
or U2513 (N_2513,N_2442,N_2496);
nor U2514 (N_2514,N_2294,N_2040);
nand U2515 (N_2515,N_2371,N_2259);
nor U2516 (N_2516,N_2061,N_2258);
nand U2517 (N_2517,N_2159,N_2081);
nand U2518 (N_2518,N_2261,N_2041);
nor U2519 (N_2519,N_2497,N_2115);
nand U2520 (N_2520,N_2270,N_2169);
and U2521 (N_2521,N_2451,N_2263);
and U2522 (N_2522,N_2375,N_2067);
xnor U2523 (N_2523,N_2483,N_2482);
or U2524 (N_2524,N_2361,N_2405);
xor U2525 (N_2525,N_2141,N_2091);
xnor U2526 (N_2526,N_2346,N_2447);
and U2527 (N_2527,N_2044,N_2367);
nand U2528 (N_2528,N_2195,N_2336);
or U2529 (N_2529,N_2284,N_2036);
nand U2530 (N_2530,N_2302,N_2053);
or U2531 (N_2531,N_2090,N_2264);
nand U2532 (N_2532,N_2325,N_2211);
xnor U2533 (N_2533,N_2292,N_2072);
nor U2534 (N_2534,N_2299,N_2022);
nand U2535 (N_2535,N_2012,N_2449);
xor U2536 (N_2536,N_2190,N_2391);
nand U2537 (N_2537,N_2202,N_2435);
and U2538 (N_2538,N_2303,N_2329);
or U2539 (N_2539,N_2382,N_2297);
or U2540 (N_2540,N_2013,N_2352);
nand U2541 (N_2541,N_2192,N_2338);
or U2542 (N_2542,N_2142,N_2278);
nand U2543 (N_2543,N_2281,N_2335);
nor U2544 (N_2544,N_2498,N_2250);
nor U2545 (N_2545,N_2466,N_2268);
xnor U2546 (N_2546,N_2314,N_2241);
nor U2547 (N_2547,N_2327,N_2117);
nor U2548 (N_2548,N_2468,N_2060);
and U2549 (N_2549,N_2016,N_2293);
and U2550 (N_2550,N_2409,N_2260);
xor U2551 (N_2551,N_2291,N_2046);
or U2552 (N_2552,N_2039,N_2461);
and U2553 (N_2553,N_2194,N_2453);
xor U2554 (N_2554,N_2369,N_2413);
nand U2555 (N_2555,N_2056,N_2062);
nor U2556 (N_2556,N_2025,N_2032);
nor U2557 (N_2557,N_2389,N_2020);
nor U2558 (N_2558,N_2140,N_2148);
or U2559 (N_2559,N_2388,N_2184);
xor U2560 (N_2560,N_2147,N_2132);
nor U2561 (N_2561,N_2310,N_2082);
or U2562 (N_2562,N_2018,N_2240);
nand U2563 (N_2563,N_2287,N_2489);
nand U2564 (N_2564,N_2394,N_2411);
or U2565 (N_2565,N_2155,N_2277);
nor U2566 (N_2566,N_2480,N_2476);
or U2567 (N_2567,N_2337,N_2017);
or U2568 (N_2568,N_2163,N_2055);
nor U2569 (N_2569,N_2216,N_2471);
and U2570 (N_2570,N_2379,N_2057);
and U2571 (N_2571,N_2478,N_2286);
or U2572 (N_2572,N_2135,N_2034);
nor U2573 (N_2573,N_2326,N_2324);
xnor U2574 (N_2574,N_2357,N_2000);
nand U2575 (N_2575,N_2331,N_2438);
and U2576 (N_2576,N_2351,N_2063);
or U2577 (N_2577,N_2199,N_2246);
and U2578 (N_2578,N_2054,N_2328);
nor U2579 (N_2579,N_2410,N_2069);
nor U2580 (N_2580,N_2064,N_2398);
nor U2581 (N_2581,N_2425,N_2348);
nor U2582 (N_2582,N_2358,N_2304);
and U2583 (N_2583,N_2455,N_2234);
xor U2584 (N_2584,N_2499,N_2474);
nand U2585 (N_2585,N_2076,N_2490);
or U2586 (N_2586,N_2058,N_2254);
or U2587 (N_2587,N_2365,N_2029);
xor U2588 (N_2588,N_2001,N_2295);
and U2589 (N_2589,N_2092,N_2030);
and U2590 (N_2590,N_2206,N_2288);
and U2591 (N_2591,N_2182,N_2154);
or U2592 (N_2592,N_2273,N_2187);
xnor U2593 (N_2593,N_2309,N_2179);
and U2594 (N_2594,N_2084,N_2350);
nand U2595 (N_2595,N_2423,N_2075);
xnor U2596 (N_2596,N_2083,N_2308);
xor U2597 (N_2597,N_2125,N_2021);
nand U2598 (N_2598,N_2005,N_2307);
and U2599 (N_2599,N_2196,N_2426);
and U2600 (N_2600,N_2276,N_2188);
or U2601 (N_2601,N_2248,N_2342);
xor U2602 (N_2602,N_2137,N_2472);
nand U2603 (N_2603,N_2218,N_2493);
and U2604 (N_2604,N_2235,N_2111);
nor U2605 (N_2605,N_2271,N_2123);
xor U2606 (N_2606,N_2395,N_2356);
or U2607 (N_2607,N_2372,N_2212);
or U2608 (N_2608,N_2122,N_2387);
xor U2609 (N_2609,N_2428,N_2150);
nor U2610 (N_2610,N_2446,N_2368);
or U2611 (N_2611,N_2006,N_2174);
nor U2612 (N_2612,N_2120,N_2253);
and U2613 (N_2613,N_2043,N_2363);
and U2614 (N_2614,N_2366,N_2401);
nor U2615 (N_2615,N_2168,N_2349);
xor U2616 (N_2616,N_2208,N_2220);
nor U2617 (N_2617,N_2024,N_2257);
or U2618 (N_2618,N_2439,N_2279);
or U2619 (N_2619,N_2093,N_2465);
and U2620 (N_2620,N_2492,N_2491);
or U2621 (N_2621,N_2215,N_2443);
or U2622 (N_2622,N_2079,N_2048);
or U2623 (N_2623,N_2101,N_2344);
nor U2624 (N_2624,N_2052,N_2045);
or U2625 (N_2625,N_2353,N_2485);
and U2626 (N_2626,N_2204,N_2186);
and U2627 (N_2627,N_2104,N_2116);
nand U2628 (N_2628,N_2010,N_2296);
xor U2629 (N_2629,N_2393,N_2422);
xnor U2630 (N_2630,N_2227,N_2033);
and U2631 (N_2631,N_2078,N_2432);
or U2632 (N_2632,N_2427,N_2272);
and U2633 (N_2633,N_2332,N_2031);
and U2634 (N_2634,N_2237,N_2097);
nand U2635 (N_2635,N_2239,N_2322);
and U2636 (N_2636,N_2473,N_2051);
or U2637 (N_2637,N_2238,N_2399);
xor U2638 (N_2638,N_2124,N_2495);
xor U2639 (N_2639,N_2330,N_2412);
nor U2640 (N_2640,N_2231,N_2225);
nand U2641 (N_2641,N_2417,N_2252);
nor U2642 (N_2642,N_2019,N_2255);
nand U2643 (N_2643,N_2305,N_2139);
or U2644 (N_2644,N_2318,N_2444);
and U2645 (N_2645,N_2089,N_2463);
or U2646 (N_2646,N_2450,N_2267);
and U2647 (N_2647,N_2378,N_2256);
xor U2648 (N_2648,N_2321,N_2103);
xnor U2649 (N_2649,N_2430,N_2200);
nand U2650 (N_2650,N_2138,N_2129);
or U2651 (N_2651,N_2477,N_2149);
or U2652 (N_2652,N_2441,N_2007);
nor U2653 (N_2653,N_2445,N_2152);
or U2654 (N_2654,N_2214,N_2153);
and U2655 (N_2655,N_2436,N_2404);
and U2656 (N_2656,N_2217,N_2136);
nor U2657 (N_2657,N_2066,N_2249);
nor U2658 (N_2658,N_2481,N_2300);
xor U2659 (N_2659,N_2157,N_2230);
nor U2660 (N_2660,N_2457,N_2128);
nand U2661 (N_2661,N_2362,N_2146);
or U2662 (N_2662,N_2080,N_2197);
nand U2663 (N_2663,N_2460,N_2143);
or U2664 (N_2664,N_2334,N_2158);
and U2665 (N_2665,N_2035,N_2429);
nor U2666 (N_2666,N_2203,N_2178);
or U2667 (N_2667,N_2345,N_2392);
and U2668 (N_2668,N_2437,N_2243);
nor U2669 (N_2669,N_2108,N_2320);
xor U2670 (N_2670,N_2201,N_2074);
nand U2671 (N_2671,N_2339,N_2088);
nand U2672 (N_2672,N_2047,N_2028);
nor U2673 (N_2673,N_2290,N_2133);
xnor U2674 (N_2674,N_2145,N_2402);
or U2675 (N_2675,N_2112,N_2377);
nand U2676 (N_2676,N_2319,N_2229);
or U2677 (N_2677,N_2347,N_2462);
nand U2678 (N_2678,N_2095,N_2121);
or U2679 (N_2679,N_2162,N_2173);
nand U2680 (N_2680,N_2233,N_2172);
xnor U2681 (N_2681,N_2301,N_2167);
nor U2682 (N_2682,N_2384,N_2488);
nand U2683 (N_2683,N_2381,N_2470);
nand U2684 (N_2684,N_2274,N_2397);
nor U2685 (N_2685,N_2285,N_2102);
nor U2686 (N_2686,N_2130,N_2364);
xnor U2687 (N_2687,N_2166,N_2113);
and U2688 (N_2688,N_2073,N_2306);
and U2689 (N_2689,N_2222,N_2494);
nor U2690 (N_2690,N_2096,N_2236);
xor U2691 (N_2691,N_2226,N_2408);
and U2692 (N_2692,N_2131,N_2386);
xnor U2693 (N_2693,N_2251,N_2244);
or U2694 (N_2694,N_2419,N_2396);
and U2695 (N_2695,N_2110,N_2099);
nor U2696 (N_2696,N_2175,N_2312);
xor U2697 (N_2697,N_2171,N_2156);
nor U2698 (N_2698,N_2106,N_2354);
or U2699 (N_2699,N_2059,N_2418);
or U2700 (N_2700,N_2340,N_2042);
and U2701 (N_2701,N_2100,N_2469);
xor U2702 (N_2702,N_2280,N_2003);
nor U2703 (N_2703,N_2209,N_2266);
nor U2704 (N_2704,N_2400,N_2380);
or U2705 (N_2705,N_2323,N_2370);
or U2706 (N_2706,N_2191,N_2118);
or U2707 (N_2707,N_2050,N_2210);
or U2708 (N_2708,N_2223,N_2383);
and U2709 (N_2709,N_2077,N_2224);
or U2710 (N_2710,N_2134,N_2406);
xnor U2711 (N_2711,N_2313,N_2085);
and U2712 (N_2712,N_2479,N_2262);
and U2713 (N_2713,N_2176,N_2298);
nand U2714 (N_2714,N_2424,N_2114);
xor U2715 (N_2715,N_2373,N_2359);
xor U2716 (N_2716,N_2487,N_2068);
xor U2717 (N_2717,N_2414,N_2170);
nor U2718 (N_2718,N_2269,N_2127);
and U2719 (N_2719,N_2205,N_2407);
or U2720 (N_2720,N_2475,N_2376);
xor U2721 (N_2721,N_2086,N_2144);
and U2722 (N_2722,N_2247,N_2448);
or U2723 (N_2723,N_2165,N_2242);
or U2724 (N_2724,N_2454,N_2180);
and U2725 (N_2725,N_2458,N_2160);
or U2726 (N_2726,N_2038,N_2316);
xor U2727 (N_2727,N_2185,N_2431);
and U2728 (N_2728,N_2026,N_2219);
nor U2729 (N_2729,N_2023,N_2008);
xor U2730 (N_2730,N_2221,N_2452);
xnor U2731 (N_2731,N_2126,N_2486);
or U2732 (N_2732,N_2421,N_2189);
nor U2733 (N_2733,N_2333,N_2317);
nand U2734 (N_2734,N_2420,N_2265);
and U2735 (N_2735,N_2109,N_2416);
nand U2736 (N_2736,N_2193,N_2181);
nor U2737 (N_2737,N_2228,N_2098);
nand U2738 (N_2738,N_2374,N_2027);
or U2739 (N_2739,N_2415,N_2434);
xnor U2740 (N_2740,N_2105,N_2315);
xnor U2741 (N_2741,N_2183,N_2037);
and U2742 (N_2742,N_2119,N_2107);
or U2743 (N_2743,N_2011,N_2456);
nand U2744 (N_2744,N_2151,N_2245);
and U2745 (N_2745,N_2002,N_2459);
or U2746 (N_2746,N_2289,N_2094);
nand U2747 (N_2747,N_2467,N_2070);
xnor U2748 (N_2748,N_2311,N_2282);
nor U2749 (N_2749,N_2275,N_2213);
nor U2750 (N_2750,N_2205,N_2156);
or U2751 (N_2751,N_2078,N_2151);
and U2752 (N_2752,N_2259,N_2402);
and U2753 (N_2753,N_2235,N_2483);
or U2754 (N_2754,N_2004,N_2351);
or U2755 (N_2755,N_2412,N_2134);
xor U2756 (N_2756,N_2425,N_2238);
xnor U2757 (N_2757,N_2498,N_2128);
or U2758 (N_2758,N_2315,N_2057);
nor U2759 (N_2759,N_2181,N_2007);
or U2760 (N_2760,N_2407,N_2147);
and U2761 (N_2761,N_2268,N_2392);
and U2762 (N_2762,N_2483,N_2271);
and U2763 (N_2763,N_2180,N_2489);
xor U2764 (N_2764,N_2230,N_2355);
or U2765 (N_2765,N_2174,N_2207);
or U2766 (N_2766,N_2047,N_2322);
nand U2767 (N_2767,N_2353,N_2110);
xor U2768 (N_2768,N_2469,N_2200);
or U2769 (N_2769,N_2278,N_2063);
nor U2770 (N_2770,N_2418,N_2066);
xnor U2771 (N_2771,N_2391,N_2243);
xor U2772 (N_2772,N_2438,N_2483);
or U2773 (N_2773,N_2339,N_2470);
nor U2774 (N_2774,N_2223,N_2454);
nor U2775 (N_2775,N_2448,N_2023);
or U2776 (N_2776,N_2269,N_2001);
and U2777 (N_2777,N_2400,N_2228);
and U2778 (N_2778,N_2341,N_2001);
xor U2779 (N_2779,N_2383,N_2208);
and U2780 (N_2780,N_2021,N_2282);
and U2781 (N_2781,N_2171,N_2367);
nor U2782 (N_2782,N_2119,N_2354);
nor U2783 (N_2783,N_2212,N_2274);
nand U2784 (N_2784,N_2460,N_2355);
nor U2785 (N_2785,N_2155,N_2419);
xnor U2786 (N_2786,N_2384,N_2464);
nor U2787 (N_2787,N_2311,N_2054);
or U2788 (N_2788,N_2270,N_2047);
xnor U2789 (N_2789,N_2371,N_2303);
or U2790 (N_2790,N_2343,N_2271);
nor U2791 (N_2791,N_2214,N_2445);
xor U2792 (N_2792,N_2320,N_2484);
and U2793 (N_2793,N_2371,N_2017);
and U2794 (N_2794,N_2291,N_2435);
xor U2795 (N_2795,N_2438,N_2482);
and U2796 (N_2796,N_2245,N_2045);
xor U2797 (N_2797,N_2473,N_2463);
nor U2798 (N_2798,N_2019,N_2240);
nor U2799 (N_2799,N_2168,N_2253);
nand U2800 (N_2800,N_2280,N_2091);
or U2801 (N_2801,N_2159,N_2073);
or U2802 (N_2802,N_2443,N_2048);
or U2803 (N_2803,N_2476,N_2440);
nand U2804 (N_2804,N_2472,N_2387);
nand U2805 (N_2805,N_2085,N_2146);
nor U2806 (N_2806,N_2129,N_2482);
nand U2807 (N_2807,N_2310,N_2115);
nand U2808 (N_2808,N_2473,N_2213);
nand U2809 (N_2809,N_2225,N_2283);
xor U2810 (N_2810,N_2399,N_2010);
xor U2811 (N_2811,N_2316,N_2143);
nor U2812 (N_2812,N_2345,N_2262);
nand U2813 (N_2813,N_2430,N_2316);
or U2814 (N_2814,N_2432,N_2131);
and U2815 (N_2815,N_2353,N_2073);
nor U2816 (N_2816,N_2239,N_2381);
xor U2817 (N_2817,N_2108,N_2146);
or U2818 (N_2818,N_2349,N_2299);
or U2819 (N_2819,N_2080,N_2342);
nand U2820 (N_2820,N_2203,N_2364);
nor U2821 (N_2821,N_2281,N_2022);
xor U2822 (N_2822,N_2268,N_2369);
nand U2823 (N_2823,N_2084,N_2020);
xor U2824 (N_2824,N_2080,N_2035);
or U2825 (N_2825,N_2068,N_2019);
nand U2826 (N_2826,N_2384,N_2400);
xnor U2827 (N_2827,N_2439,N_2164);
xor U2828 (N_2828,N_2080,N_2200);
nor U2829 (N_2829,N_2174,N_2204);
or U2830 (N_2830,N_2417,N_2432);
nand U2831 (N_2831,N_2094,N_2332);
or U2832 (N_2832,N_2209,N_2153);
or U2833 (N_2833,N_2063,N_2492);
xor U2834 (N_2834,N_2018,N_2274);
or U2835 (N_2835,N_2000,N_2164);
nor U2836 (N_2836,N_2155,N_2013);
and U2837 (N_2837,N_2288,N_2124);
nor U2838 (N_2838,N_2211,N_2171);
and U2839 (N_2839,N_2090,N_2366);
xor U2840 (N_2840,N_2242,N_2314);
and U2841 (N_2841,N_2405,N_2251);
nor U2842 (N_2842,N_2352,N_2184);
nand U2843 (N_2843,N_2099,N_2036);
xnor U2844 (N_2844,N_2137,N_2241);
or U2845 (N_2845,N_2095,N_2202);
nand U2846 (N_2846,N_2307,N_2197);
or U2847 (N_2847,N_2138,N_2397);
nand U2848 (N_2848,N_2013,N_2047);
xor U2849 (N_2849,N_2326,N_2406);
and U2850 (N_2850,N_2032,N_2046);
nor U2851 (N_2851,N_2113,N_2060);
nand U2852 (N_2852,N_2330,N_2335);
and U2853 (N_2853,N_2439,N_2230);
nand U2854 (N_2854,N_2022,N_2051);
nand U2855 (N_2855,N_2450,N_2301);
nand U2856 (N_2856,N_2272,N_2210);
nand U2857 (N_2857,N_2259,N_2050);
xnor U2858 (N_2858,N_2309,N_2083);
xor U2859 (N_2859,N_2423,N_2011);
nand U2860 (N_2860,N_2194,N_2336);
nor U2861 (N_2861,N_2422,N_2353);
or U2862 (N_2862,N_2284,N_2315);
nand U2863 (N_2863,N_2353,N_2415);
nand U2864 (N_2864,N_2244,N_2144);
and U2865 (N_2865,N_2335,N_2420);
xnor U2866 (N_2866,N_2402,N_2342);
xnor U2867 (N_2867,N_2092,N_2480);
and U2868 (N_2868,N_2261,N_2236);
or U2869 (N_2869,N_2176,N_2491);
or U2870 (N_2870,N_2207,N_2124);
nor U2871 (N_2871,N_2082,N_2385);
nor U2872 (N_2872,N_2149,N_2400);
xnor U2873 (N_2873,N_2131,N_2185);
nor U2874 (N_2874,N_2423,N_2120);
and U2875 (N_2875,N_2240,N_2186);
nand U2876 (N_2876,N_2020,N_2104);
and U2877 (N_2877,N_2186,N_2159);
and U2878 (N_2878,N_2281,N_2048);
xnor U2879 (N_2879,N_2349,N_2060);
nor U2880 (N_2880,N_2485,N_2028);
or U2881 (N_2881,N_2468,N_2273);
or U2882 (N_2882,N_2216,N_2401);
nand U2883 (N_2883,N_2005,N_2204);
nand U2884 (N_2884,N_2490,N_2162);
nor U2885 (N_2885,N_2244,N_2140);
nor U2886 (N_2886,N_2420,N_2286);
nor U2887 (N_2887,N_2336,N_2015);
nor U2888 (N_2888,N_2471,N_2072);
and U2889 (N_2889,N_2354,N_2486);
and U2890 (N_2890,N_2354,N_2076);
and U2891 (N_2891,N_2477,N_2041);
and U2892 (N_2892,N_2216,N_2083);
and U2893 (N_2893,N_2153,N_2210);
and U2894 (N_2894,N_2275,N_2402);
and U2895 (N_2895,N_2314,N_2219);
or U2896 (N_2896,N_2035,N_2247);
and U2897 (N_2897,N_2381,N_2102);
nand U2898 (N_2898,N_2480,N_2136);
and U2899 (N_2899,N_2147,N_2347);
xnor U2900 (N_2900,N_2214,N_2006);
and U2901 (N_2901,N_2391,N_2474);
xnor U2902 (N_2902,N_2021,N_2104);
nand U2903 (N_2903,N_2353,N_2346);
or U2904 (N_2904,N_2412,N_2283);
nand U2905 (N_2905,N_2319,N_2227);
nand U2906 (N_2906,N_2001,N_2301);
or U2907 (N_2907,N_2382,N_2143);
nand U2908 (N_2908,N_2137,N_2064);
nor U2909 (N_2909,N_2184,N_2214);
nor U2910 (N_2910,N_2360,N_2254);
and U2911 (N_2911,N_2221,N_2336);
nor U2912 (N_2912,N_2234,N_2173);
nand U2913 (N_2913,N_2409,N_2041);
and U2914 (N_2914,N_2413,N_2006);
nand U2915 (N_2915,N_2426,N_2096);
or U2916 (N_2916,N_2429,N_2012);
nor U2917 (N_2917,N_2364,N_2403);
and U2918 (N_2918,N_2429,N_2490);
nor U2919 (N_2919,N_2449,N_2492);
and U2920 (N_2920,N_2175,N_2030);
nand U2921 (N_2921,N_2411,N_2148);
nand U2922 (N_2922,N_2447,N_2491);
nand U2923 (N_2923,N_2490,N_2018);
xor U2924 (N_2924,N_2232,N_2230);
nor U2925 (N_2925,N_2490,N_2038);
and U2926 (N_2926,N_2030,N_2157);
or U2927 (N_2927,N_2174,N_2430);
and U2928 (N_2928,N_2157,N_2282);
and U2929 (N_2929,N_2044,N_2409);
or U2930 (N_2930,N_2289,N_2016);
xor U2931 (N_2931,N_2210,N_2452);
nand U2932 (N_2932,N_2189,N_2334);
nor U2933 (N_2933,N_2344,N_2460);
and U2934 (N_2934,N_2345,N_2247);
and U2935 (N_2935,N_2305,N_2112);
and U2936 (N_2936,N_2229,N_2372);
nor U2937 (N_2937,N_2086,N_2038);
and U2938 (N_2938,N_2205,N_2067);
or U2939 (N_2939,N_2401,N_2056);
nand U2940 (N_2940,N_2358,N_2086);
nor U2941 (N_2941,N_2156,N_2432);
and U2942 (N_2942,N_2449,N_2483);
nor U2943 (N_2943,N_2294,N_2086);
and U2944 (N_2944,N_2407,N_2428);
nand U2945 (N_2945,N_2329,N_2052);
and U2946 (N_2946,N_2076,N_2465);
or U2947 (N_2947,N_2291,N_2363);
and U2948 (N_2948,N_2028,N_2033);
xor U2949 (N_2949,N_2463,N_2232);
nand U2950 (N_2950,N_2391,N_2324);
or U2951 (N_2951,N_2134,N_2242);
or U2952 (N_2952,N_2293,N_2004);
or U2953 (N_2953,N_2402,N_2354);
xnor U2954 (N_2954,N_2414,N_2297);
or U2955 (N_2955,N_2345,N_2164);
nor U2956 (N_2956,N_2337,N_2116);
nor U2957 (N_2957,N_2279,N_2235);
xnor U2958 (N_2958,N_2061,N_2386);
xnor U2959 (N_2959,N_2489,N_2221);
nor U2960 (N_2960,N_2018,N_2045);
and U2961 (N_2961,N_2000,N_2376);
nand U2962 (N_2962,N_2397,N_2255);
or U2963 (N_2963,N_2304,N_2462);
and U2964 (N_2964,N_2345,N_2265);
or U2965 (N_2965,N_2372,N_2187);
and U2966 (N_2966,N_2163,N_2459);
and U2967 (N_2967,N_2020,N_2291);
nand U2968 (N_2968,N_2099,N_2383);
xnor U2969 (N_2969,N_2394,N_2418);
nor U2970 (N_2970,N_2215,N_2367);
or U2971 (N_2971,N_2488,N_2241);
xor U2972 (N_2972,N_2017,N_2126);
or U2973 (N_2973,N_2317,N_2314);
nor U2974 (N_2974,N_2022,N_2467);
nand U2975 (N_2975,N_2022,N_2011);
nor U2976 (N_2976,N_2463,N_2299);
and U2977 (N_2977,N_2148,N_2276);
xor U2978 (N_2978,N_2276,N_2133);
xor U2979 (N_2979,N_2108,N_2000);
and U2980 (N_2980,N_2451,N_2082);
xnor U2981 (N_2981,N_2082,N_2321);
and U2982 (N_2982,N_2063,N_2468);
nand U2983 (N_2983,N_2353,N_2467);
xor U2984 (N_2984,N_2092,N_2268);
nand U2985 (N_2985,N_2282,N_2069);
xor U2986 (N_2986,N_2210,N_2089);
or U2987 (N_2987,N_2381,N_2466);
and U2988 (N_2988,N_2225,N_2258);
and U2989 (N_2989,N_2110,N_2344);
nand U2990 (N_2990,N_2375,N_2349);
and U2991 (N_2991,N_2443,N_2183);
nor U2992 (N_2992,N_2090,N_2412);
and U2993 (N_2993,N_2067,N_2219);
nand U2994 (N_2994,N_2199,N_2021);
nand U2995 (N_2995,N_2412,N_2291);
xor U2996 (N_2996,N_2230,N_2408);
or U2997 (N_2997,N_2160,N_2494);
or U2998 (N_2998,N_2361,N_2448);
nor U2999 (N_2999,N_2128,N_2135);
and U3000 (N_3000,N_2634,N_2860);
or U3001 (N_3001,N_2770,N_2824);
nor U3002 (N_3002,N_2542,N_2889);
xnor U3003 (N_3003,N_2899,N_2747);
nand U3004 (N_3004,N_2769,N_2852);
nand U3005 (N_3005,N_2514,N_2718);
or U3006 (N_3006,N_2788,N_2954);
nand U3007 (N_3007,N_2555,N_2736);
xor U3008 (N_3008,N_2582,N_2951);
nor U3009 (N_3009,N_2746,N_2971);
and U3010 (N_3010,N_2898,N_2664);
or U3011 (N_3011,N_2610,N_2638);
or U3012 (N_3012,N_2503,N_2841);
nor U3013 (N_3013,N_2731,N_2932);
nand U3014 (N_3014,N_2957,N_2553);
xor U3015 (N_3015,N_2512,N_2533);
nand U3016 (N_3016,N_2984,N_2863);
and U3017 (N_3017,N_2600,N_2504);
nand U3018 (N_3018,N_2569,N_2843);
nor U3019 (N_3019,N_2689,N_2607);
nand U3020 (N_3020,N_2719,N_2847);
nand U3021 (N_3021,N_2619,N_2606);
nand U3022 (N_3022,N_2869,N_2922);
nand U3023 (N_3023,N_2727,N_2846);
or U3024 (N_3024,N_2953,N_2609);
nand U3025 (N_3025,N_2637,N_2868);
or U3026 (N_3026,N_2790,N_2945);
and U3027 (N_3027,N_2981,N_2862);
nor U3028 (N_3028,N_2982,N_2651);
nand U3029 (N_3029,N_2670,N_2848);
and U3030 (N_3030,N_2726,N_2837);
or U3031 (N_3031,N_2585,N_2732);
nand U3032 (N_3032,N_2884,N_2591);
and U3033 (N_3033,N_2743,N_2794);
nand U3034 (N_3034,N_2778,N_2567);
nor U3035 (N_3035,N_2818,N_2693);
or U3036 (N_3036,N_2784,N_2621);
or U3037 (N_3037,N_2574,N_2838);
or U3038 (N_3038,N_2738,N_2545);
and U3039 (N_3039,N_2825,N_2844);
nand U3040 (N_3040,N_2763,N_2781);
nand U3041 (N_3041,N_2717,N_2563);
and U3042 (N_3042,N_2723,N_2509);
and U3043 (N_3043,N_2827,N_2682);
nor U3044 (N_3044,N_2835,N_2686);
or U3045 (N_3045,N_2615,N_2766);
or U3046 (N_3046,N_2876,N_2739);
xor U3047 (N_3047,N_2668,N_2920);
and U3048 (N_3048,N_2614,N_2602);
and U3049 (N_3049,N_2928,N_2939);
or U3050 (N_3050,N_2687,N_2931);
nand U3051 (N_3051,N_2777,N_2677);
nand U3052 (N_3052,N_2640,N_2722);
xor U3053 (N_3053,N_2989,N_2887);
nand U3054 (N_3054,N_2660,N_2833);
nor U3055 (N_3055,N_2894,N_2577);
xor U3056 (N_3056,N_2879,N_2758);
xor U3057 (N_3057,N_2683,N_2870);
nor U3058 (N_3058,N_2537,N_2705);
nor U3059 (N_3059,N_2517,N_2978);
nor U3060 (N_3060,N_2720,N_2562);
xor U3061 (N_3061,N_2616,N_2901);
nor U3062 (N_3062,N_2776,N_2895);
xnor U3063 (N_3063,N_2923,N_2772);
xnor U3064 (N_3064,N_2699,N_2540);
xor U3065 (N_3065,N_2905,N_2930);
or U3066 (N_3066,N_2810,N_2539);
or U3067 (N_3067,N_2851,N_2696);
nand U3068 (N_3068,N_2821,N_2544);
nor U3069 (N_3069,N_2890,N_2783);
nand U3070 (N_3070,N_2855,N_2605);
nand U3071 (N_3071,N_2962,N_2815);
nand U3072 (N_3072,N_2710,N_2526);
and U3073 (N_3073,N_2673,N_2612);
and U3074 (N_3074,N_2633,N_2628);
nor U3075 (N_3075,N_2506,N_2875);
or U3076 (N_3076,N_2573,N_2775);
xor U3077 (N_3077,N_2538,N_2771);
and U3078 (N_3078,N_2749,N_2625);
nor U3079 (N_3079,N_2698,N_2589);
xor U3080 (N_3080,N_2636,N_2907);
nand U3081 (N_3081,N_2795,N_2976);
nand U3082 (N_3082,N_2566,N_2934);
nor U3083 (N_3083,N_2830,N_2631);
or U3084 (N_3084,N_2871,N_2762);
and U3085 (N_3085,N_2842,N_2571);
nand U3086 (N_3086,N_2532,N_2948);
and U3087 (N_3087,N_2613,N_2570);
and U3088 (N_3088,N_2946,N_2583);
or U3089 (N_3089,N_2801,N_2599);
nand U3090 (N_3090,N_2734,N_2992);
and U3091 (N_3091,N_2767,N_2867);
and U3092 (N_3092,N_2750,N_2950);
and U3093 (N_3093,N_2590,N_2858);
nand U3094 (N_3094,N_2888,N_2706);
xnor U3095 (N_3095,N_2961,N_2559);
nand U3096 (N_3096,N_2986,N_2617);
and U3097 (N_3097,N_2725,N_2697);
nor U3098 (N_3098,N_2803,N_2534);
and U3099 (N_3099,N_2715,N_2672);
or U3100 (N_3100,N_2845,N_2942);
or U3101 (N_3101,N_2787,N_2520);
xnor U3102 (N_3102,N_2754,N_2780);
nand U3103 (N_3103,N_2753,N_2941);
nand U3104 (N_3104,N_2740,N_2891);
nor U3105 (N_3105,N_2674,N_2756);
nor U3106 (N_3106,N_2565,N_2690);
and U3107 (N_3107,N_2505,N_2707);
and U3108 (N_3108,N_2921,N_2575);
or U3109 (N_3109,N_2759,N_2700);
nand U3110 (N_3110,N_2958,N_2635);
xor U3111 (N_3111,N_2949,N_2912);
or U3112 (N_3112,N_2695,N_2861);
and U3113 (N_3113,N_2798,N_2676);
or U3114 (N_3114,N_2712,N_2974);
nand U3115 (N_3115,N_2983,N_2659);
or U3116 (N_3116,N_2977,N_2938);
and U3117 (N_3117,N_2550,N_2704);
or U3118 (N_3118,N_2782,N_2935);
or U3119 (N_3119,N_2748,N_2850);
nand U3120 (N_3120,N_2998,N_2655);
nor U3121 (N_3121,N_2711,N_2521);
nand U3122 (N_3122,N_2987,N_2929);
or U3123 (N_3123,N_2530,N_2866);
xnor U3124 (N_3124,N_2880,N_2805);
xnor U3125 (N_3125,N_2502,N_2995);
nor U3126 (N_3126,N_2908,N_2709);
and U3127 (N_3127,N_2809,N_2996);
or U3128 (N_3128,N_2915,N_2856);
nor U3129 (N_3129,N_2630,N_2826);
nor U3130 (N_3130,N_2642,N_2701);
xnor U3131 (N_3131,N_2729,N_2812);
xnor U3132 (N_3132,N_2691,N_2800);
or U3133 (N_3133,N_2933,N_2873);
and U3134 (N_3134,N_2814,N_2947);
and U3135 (N_3135,N_2654,N_2904);
and U3136 (N_3136,N_2618,N_2593);
or U3137 (N_3137,N_2581,N_2797);
or U3138 (N_3138,N_2561,N_2597);
xnor U3139 (N_3139,N_2666,N_2528);
xnor U3140 (N_3140,N_2716,N_2808);
xnor U3141 (N_3141,N_2557,N_2546);
or U3142 (N_3142,N_2902,N_2822);
and U3143 (N_3143,N_2547,N_2745);
nand U3144 (N_3144,N_2556,N_2604);
xor U3145 (N_3145,N_2596,N_2598);
or U3146 (N_3146,N_2507,N_2874);
nor U3147 (N_3147,N_2737,N_2649);
or U3148 (N_3148,N_2807,N_2658);
and U3149 (N_3149,N_2892,N_2878);
and U3150 (N_3150,N_2603,N_2648);
or U3151 (N_3151,N_2911,N_2966);
nor U3152 (N_3152,N_2975,N_2688);
nand U3153 (N_3153,N_2882,N_2963);
and U3154 (N_3154,N_2518,N_2595);
and U3155 (N_3155,N_2973,N_2501);
nor U3156 (N_3156,N_2926,N_2587);
nand U3157 (N_3157,N_2955,N_2832);
or U3158 (N_3158,N_2681,N_2548);
and U3159 (N_3159,N_2900,N_2786);
and U3160 (N_3160,N_2624,N_2991);
and U3161 (N_3161,N_2968,N_2985);
nand U3162 (N_3162,N_2657,N_2647);
xor U3163 (N_3163,N_2853,N_2865);
nand U3164 (N_3164,N_2979,N_2760);
nand U3165 (N_3165,N_2755,N_2918);
nand U3166 (N_3166,N_2592,N_2529);
and U3167 (N_3167,N_2541,N_2831);
and U3168 (N_3168,N_2694,N_2924);
or U3169 (N_3169,N_2972,N_2988);
or U3170 (N_3170,N_2531,N_2993);
or U3171 (N_3171,N_2752,N_2936);
xor U3172 (N_3172,N_2857,N_2774);
nand U3173 (N_3173,N_2765,N_2910);
and U3174 (N_3174,N_2896,N_2644);
nand U3175 (N_3175,N_2646,N_2864);
and U3176 (N_3176,N_2836,N_2513);
xor U3177 (N_3177,N_2543,N_2943);
nor U3178 (N_3178,N_2669,N_2535);
and U3179 (N_3179,N_2632,N_2925);
or U3180 (N_3180,N_2940,N_2527);
xor U3181 (N_3181,N_2671,N_2956);
or U3182 (N_3182,N_2620,N_2588);
nand U3183 (N_3183,N_2714,N_2702);
or U3184 (N_3184,N_2703,N_2893);
and U3185 (N_3185,N_2761,N_2560);
or U3186 (N_3186,N_2576,N_2829);
nand U3187 (N_3187,N_2578,N_2508);
and U3188 (N_3188,N_2819,N_2802);
xor U3189 (N_3189,N_2713,N_2906);
nand U3190 (N_3190,N_2652,N_2653);
nand U3191 (N_3191,N_2735,N_2679);
nor U3192 (N_3192,N_2678,N_2629);
and U3193 (N_3193,N_2594,N_2622);
xor U3194 (N_3194,N_2849,N_2662);
and U3195 (N_3195,N_2627,N_2885);
nand U3196 (N_3196,N_2779,N_2515);
or U3197 (N_3197,N_2744,N_2913);
and U3198 (N_3198,N_2919,N_2584);
nand U3199 (N_3199,N_2708,N_2859);
xor U3200 (N_3200,N_2969,N_2768);
nand U3201 (N_3201,N_2680,N_2970);
nand U3202 (N_3202,N_2839,N_2959);
nand U3203 (N_3203,N_2645,N_2733);
xnor U3204 (N_3204,N_2917,N_2773);
nor U3205 (N_3205,N_2828,N_2523);
and U3206 (N_3206,N_2952,N_2967);
or U3207 (N_3207,N_2685,N_2536);
xnor U3208 (N_3208,N_2579,N_2823);
nand U3209 (N_3209,N_2611,N_2791);
and U3210 (N_3210,N_2785,N_2854);
nand U3211 (N_3211,N_2883,N_2927);
nor U3212 (N_3212,N_2564,N_2799);
and U3213 (N_3213,N_2751,N_2623);
or U3214 (N_3214,N_2549,N_2572);
and U3215 (N_3215,N_2840,N_2519);
and U3216 (N_3216,N_2516,N_2994);
or U3217 (N_3217,N_2554,N_2834);
or U3218 (N_3218,N_2813,N_2524);
or U3219 (N_3219,N_2764,N_2789);
and U3220 (N_3220,N_2999,N_2793);
nand U3221 (N_3221,N_2692,N_2684);
or U3222 (N_3222,N_2665,N_2881);
xnor U3223 (N_3223,N_2980,N_2663);
or U3224 (N_3224,N_2897,N_2990);
nand U3225 (N_3225,N_2656,N_2728);
and U3226 (N_3226,N_2960,N_2817);
and U3227 (N_3227,N_2877,N_2724);
nor U3228 (N_3228,N_2580,N_2650);
or U3229 (N_3229,N_2641,N_2558);
xnor U3230 (N_3230,N_2500,N_2742);
nor U3231 (N_3231,N_2804,N_2551);
and U3232 (N_3232,N_2552,N_2608);
nor U3233 (N_3233,N_2903,N_2997);
nor U3234 (N_3234,N_2820,N_2643);
and U3235 (N_3235,N_2510,N_2964);
and U3236 (N_3236,N_2872,N_2909);
and U3237 (N_3237,N_2916,N_2721);
or U3238 (N_3238,N_2937,N_2525);
nand U3239 (N_3239,N_2511,N_2586);
and U3240 (N_3240,N_2792,N_2811);
or U3241 (N_3241,N_2796,N_2667);
xnor U3242 (N_3242,N_2730,N_2522);
xor U3243 (N_3243,N_2675,N_2626);
nand U3244 (N_3244,N_2601,N_2639);
xor U3245 (N_3245,N_2886,N_2944);
nor U3246 (N_3246,N_2757,N_2661);
and U3247 (N_3247,N_2914,N_2741);
or U3248 (N_3248,N_2816,N_2965);
and U3249 (N_3249,N_2568,N_2806);
xor U3250 (N_3250,N_2766,N_2651);
nor U3251 (N_3251,N_2641,N_2849);
nand U3252 (N_3252,N_2567,N_2538);
nand U3253 (N_3253,N_2873,N_2681);
or U3254 (N_3254,N_2649,N_2789);
and U3255 (N_3255,N_2963,N_2590);
nand U3256 (N_3256,N_2767,N_2976);
xnor U3257 (N_3257,N_2787,N_2640);
xor U3258 (N_3258,N_2773,N_2653);
xnor U3259 (N_3259,N_2958,N_2640);
or U3260 (N_3260,N_2912,N_2679);
or U3261 (N_3261,N_2952,N_2759);
xnor U3262 (N_3262,N_2621,N_2737);
and U3263 (N_3263,N_2567,N_2777);
xor U3264 (N_3264,N_2527,N_2650);
and U3265 (N_3265,N_2656,N_2957);
and U3266 (N_3266,N_2501,N_2670);
xnor U3267 (N_3267,N_2659,N_2549);
or U3268 (N_3268,N_2926,N_2779);
nand U3269 (N_3269,N_2571,N_2898);
or U3270 (N_3270,N_2882,N_2918);
or U3271 (N_3271,N_2570,N_2607);
nor U3272 (N_3272,N_2506,N_2891);
and U3273 (N_3273,N_2643,N_2771);
nand U3274 (N_3274,N_2998,N_2625);
and U3275 (N_3275,N_2586,N_2516);
and U3276 (N_3276,N_2549,N_2545);
or U3277 (N_3277,N_2590,N_2900);
and U3278 (N_3278,N_2837,N_2869);
xnor U3279 (N_3279,N_2898,N_2838);
and U3280 (N_3280,N_2916,N_2524);
or U3281 (N_3281,N_2947,N_2527);
nand U3282 (N_3282,N_2504,N_2690);
or U3283 (N_3283,N_2684,N_2656);
and U3284 (N_3284,N_2685,N_2931);
nand U3285 (N_3285,N_2534,N_2617);
and U3286 (N_3286,N_2587,N_2745);
and U3287 (N_3287,N_2869,N_2606);
xor U3288 (N_3288,N_2720,N_2671);
xnor U3289 (N_3289,N_2910,N_2698);
xor U3290 (N_3290,N_2555,N_2527);
nor U3291 (N_3291,N_2708,N_2921);
and U3292 (N_3292,N_2781,N_2623);
and U3293 (N_3293,N_2723,N_2963);
nand U3294 (N_3294,N_2507,N_2558);
nor U3295 (N_3295,N_2504,N_2718);
nor U3296 (N_3296,N_2811,N_2862);
nand U3297 (N_3297,N_2523,N_2941);
nand U3298 (N_3298,N_2754,N_2736);
and U3299 (N_3299,N_2893,N_2681);
nor U3300 (N_3300,N_2984,N_2706);
xnor U3301 (N_3301,N_2843,N_2558);
or U3302 (N_3302,N_2763,N_2620);
xor U3303 (N_3303,N_2797,N_2644);
nor U3304 (N_3304,N_2612,N_2503);
nor U3305 (N_3305,N_2733,N_2958);
nand U3306 (N_3306,N_2868,N_2524);
and U3307 (N_3307,N_2687,N_2720);
xnor U3308 (N_3308,N_2903,N_2819);
xor U3309 (N_3309,N_2827,N_2757);
nand U3310 (N_3310,N_2691,N_2641);
nor U3311 (N_3311,N_2964,N_2547);
nor U3312 (N_3312,N_2691,N_2739);
xnor U3313 (N_3313,N_2932,N_2937);
or U3314 (N_3314,N_2665,N_2942);
and U3315 (N_3315,N_2928,N_2755);
nor U3316 (N_3316,N_2711,N_2883);
or U3317 (N_3317,N_2913,N_2609);
nand U3318 (N_3318,N_2695,N_2981);
or U3319 (N_3319,N_2703,N_2530);
and U3320 (N_3320,N_2895,N_2635);
nand U3321 (N_3321,N_2516,N_2530);
xor U3322 (N_3322,N_2961,N_2845);
and U3323 (N_3323,N_2887,N_2787);
nor U3324 (N_3324,N_2770,N_2903);
nor U3325 (N_3325,N_2715,N_2717);
and U3326 (N_3326,N_2898,N_2831);
or U3327 (N_3327,N_2910,N_2878);
nor U3328 (N_3328,N_2518,N_2777);
and U3329 (N_3329,N_2717,N_2519);
or U3330 (N_3330,N_2800,N_2980);
xor U3331 (N_3331,N_2615,N_2536);
and U3332 (N_3332,N_2897,N_2533);
or U3333 (N_3333,N_2983,N_2632);
nand U3334 (N_3334,N_2760,N_2696);
nor U3335 (N_3335,N_2534,N_2713);
nor U3336 (N_3336,N_2715,N_2923);
nand U3337 (N_3337,N_2790,N_2611);
nor U3338 (N_3338,N_2545,N_2539);
nand U3339 (N_3339,N_2802,N_2578);
or U3340 (N_3340,N_2826,N_2882);
xor U3341 (N_3341,N_2725,N_2717);
xor U3342 (N_3342,N_2652,N_2538);
or U3343 (N_3343,N_2588,N_2930);
nor U3344 (N_3344,N_2998,N_2588);
xor U3345 (N_3345,N_2720,N_2634);
nand U3346 (N_3346,N_2867,N_2511);
nor U3347 (N_3347,N_2748,N_2957);
nand U3348 (N_3348,N_2803,N_2888);
xnor U3349 (N_3349,N_2924,N_2508);
or U3350 (N_3350,N_2870,N_2618);
nand U3351 (N_3351,N_2744,N_2652);
xor U3352 (N_3352,N_2647,N_2565);
nor U3353 (N_3353,N_2557,N_2715);
nor U3354 (N_3354,N_2675,N_2917);
xnor U3355 (N_3355,N_2715,N_2809);
nand U3356 (N_3356,N_2643,N_2660);
xnor U3357 (N_3357,N_2700,N_2668);
xnor U3358 (N_3358,N_2837,N_2989);
and U3359 (N_3359,N_2988,N_2918);
and U3360 (N_3360,N_2555,N_2632);
xnor U3361 (N_3361,N_2637,N_2638);
xnor U3362 (N_3362,N_2843,N_2626);
nand U3363 (N_3363,N_2777,N_2534);
xnor U3364 (N_3364,N_2920,N_2937);
xnor U3365 (N_3365,N_2834,N_2804);
or U3366 (N_3366,N_2812,N_2837);
and U3367 (N_3367,N_2607,N_2947);
or U3368 (N_3368,N_2955,N_2538);
or U3369 (N_3369,N_2623,N_2678);
nand U3370 (N_3370,N_2598,N_2815);
or U3371 (N_3371,N_2856,N_2517);
and U3372 (N_3372,N_2798,N_2593);
nand U3373 (N_3373,N_2589,N_2696);
or U3374 (N_3374,N_2820,N_2985);
or U3375 (N_3375,N_2841,N_2737);
xor U3376 (N_3376,N_2973,N_2897);
nor U3377 (N_3377,N_2693,N_2528);
or U3378 (N_3378,N_2927,N_2546);
nand U3379 (N_3379,N_2561,N_2943);
nand U3380 (N_3380,N_2818,N_2780);
and U3381 (N_3381,N_2942,N_2893);
nor U3382 (N_3382,N_2992,N_2909);
nand U3383 (N_3383,N_2979,N_2748);
nor U3384 (N_3384,N_2824,N_2849);
nand U3385 (N_3385,N_2634,N_2653);
nor U3386 (N_3386,N_2747,N_2527);
or U3387 (N_3387,N_2772,N_2696);
or U3388 (N_3388,N_2528,N_2998);
nor U3389 (N_3389,N_2640,N_2676);
nor U3390 (N_3390,N_2904,N_2597);
xor U3391 (N_3391,N_2507,N_2746);
or U3392 (N_3392,N_2677,N_2728);
nand U3393 (N_3393,N_2889,N_2539);
nand U3394 (N_3394,N_2598,N_2790);
and U3395 (N_3395,N_2946,N_2528);
nor U3396 (N_3396,N_2594,N_2646);
xnor U3397 (N_3397,N_2985,N_2636);
nor U3398 (N_3398,N_2743,N_2822);
nand U3399 (N_3399,N_2791,N_2659);
nand U3400 (N_3400,N_2570,N_2869);
nor U3401 (N_3401,N_2880,N_2597);
nand U3402 (N_3402,N_2701,N_2727);
or U3403 (N_3403,N_2752,N_2730);
and U3404 (N_3404,N_2535,N_2747);
nor U3405 (N_3405,N_2603,N_2992);
nor U3406 (N_3406,N_2680,N_2668);
nand U3407 (N_3407,N_2550,N_2792);
xnor U3408 (N_3408,N_2733,N_2600);
and U3409 (N_3409,N_2747,N_2772);
nor U3410 (N_3410,N_2712,N_2744);
or U3411 (N_3411,N_2698,N_2671);
nor U3412 (N_3412,N_2833,N_2997);
nand U3413 (N_3413,N_2569,N_2967);
or U3414 (N_3414,N_2724,N_2800);
or U3415 (N_3415,N_2972,N_2829);
nor U3416 (N_3416,N_2798,N_2502);
xor U3417 (N_3417,N_2541,N_2784);
or U3418 (N_3418,N_2638,N_2891);
nor U3419 (N_3419,N_2802,N_2799);
and U3420 (N_3420,N_2609,N_2858);
nor U3421 (N_3421,N_2536,N_2575);
xor U3422 (N_3422,N_2792,N_2637);
nor U3423 (N_3423,N_2766,N_2561);
or U3424 (N_3424,N_2728,N_2823);
nand U3425 (N_3425,N_2680,N_2981);
and U3426 (N_3426,N_2544,N_2929);
nor U3427 (N_3427,N_2557,N_2501);
and U3428 (N_3428,N_2841,N_2878);
or U3429 (N_3429,N_2674,N_2601);
and U3430 (N_3430,N_2614,N_2918);
xor U3431 (N_3431,N_2835,N_2905);
xor U3432 (N_3432,N_2704,N_2930);
nor U3433 (N_3433,N_2532,N_2860);
and U3434 (N_3434,N_2951,N_2561);
or U3435 (N_3435,N_2927,N_2775);
nor U3436 (N_3436,N_2661,N_2731);
nor U3437 (N_3437,N_2762,N_2547);
or U3438 (N_3438,N_2892,N_2585);
xor U3439 (N_3439,N_2781,N_2777);
or U3440 (N_3440,N_2836,N_2639);
xor U3441 (N_3441,N_2618,N_2835);
xor U3442 (N_3442,N_2730,N_2525);
and U3443 (N_3443,N_2679,N_2658);
and U3444 (N_3444,N_2640,N_2564);
xor U3445 (N_3445,N_2649,N_2960);
and U3446 (N_3446,N_2930,N_2746);
and U3447 (N_3447,N_2643,N_2806);
xor U3448 (N_3448,N_2635,N_2823);
xnor U3449 (N_3449,N_2687,N_2518);
xor U3450 (N_3450,N_2940,N_2718);
xnor U3451 (N_3451,N_2603,N_2642);
and U3452 (N_3452,N_2947,N_2890);
nand U3453 (N_3453,N_2791,N_2976);
and U3454 (N_3454,N_2502,N_2884);
nand U3455 (N_3455,N_2741,N_2532);
nand U3456 (N_3456,N_2898,N_2597);
nand U3457 (N_3457,N_2808,N_2695);
and U3458 (N_3458,N_2547,N_2639);
nor U3459 (N_3459,N_2975,N_2520);
nor U3460 (N_3460,N_2782,N_2672);
or U3461 (N_3461,N_2613,N_2828);
xnor U3462 (N_3462,N_2796,N_2946);
xor U3463 (N_3463,N_2872,N_2857);
or U3464 (N_3464,N_2726,N_2886);
xnor U3465 (N_3465,N_2585,N_2993);
nand U3466 (N_3466,N_2717,N_2977);
or U3467 (N_3467,N_2519,N_2941);
nor U3468 (N_3468,N_2870,N_2651);
and U3469 (N_3469,N_2774,N_2834);
nand U3470 (N_3470,N_2792,N_2925);
nor U3471 (N_3471,N_2650,N_2657);
xor U3472 (N_3472,N_2710,N_2743);
xnor U3473 (N_3473,N_2663,N_2774);
and U3474 (N_3474,N_2592,N_2703);
or U3475 (N_3475,N_2917,N_2659);
nor U3476 (N_3476,N_2740,N_2618);
nand U3477 (N_3477,N_2768,N_2805);
xnor U3478 (N_3478,N_2724,N_2507);
nand U3479 (N_3479,N_2633,N_2643);
xnor U3480 (N_3480,N_2836,N_2953);
nor U3481 (N_3481,N_2981,N_2572);
and U3482 (N_3482,N_2838,N_2670);
nand U3483 (N_3483,N_2551,N_2910);
nand U3484 (N_3484,N_2633,N_2846);
and U3485 (N_3485,N_2557,N_2783);
nand U3486 (N_3486,N_2791,N_2977);
nand U3487 (N_3487,N_2845,N_2868);
nor U3488 (N_3488,N_2840,N_2849);
or U3489 (N_3489,N_2879,N_2539);
and U3490 (N_3490,N_2802,N_2759);
nand U3491 (N_3491,N_2681,N_2706);
nand U3492 (N_3492,N_2555,N_2694);
nor U3493 (N_3493,N_2534,N_2692);
or U3494 (N_3494,N_2777,N_2601);
nor U3495 (N_3495,N_2956,N_2753);
and U3496 (N_3496,N_2879,N_2850);
nand U3497 (N_3497,N_2760,N_2615);
and U3498 (N_3498,N_2622,N_2710);
and U3499 (N_3499,N_2522,N_2990);
or U3500 (N_3500,N_3246,N_3240);
and U3501 (N_3501,N_3045,N_3079);
xor U3502 (N_3502,N_3161,N_3227);
nand U3503 (N_3503,N_3044,N_3210);
and U3504 (N_3504,N_3352,N_3415);
nand U3505 (N_3505,N_3242,N_3299);
and U3506 (N_3506,N_3008,N_3357);
nand U3507 (N_3507,N_3050,N_3325);
xor U3508 (N_3508,N_3305,N_3365);
or U3509 (N_3509,N_3165,N_3324);
and U3510 (N_3510,N_3274,N_3424);
nor U3511 (N_3511,N_3173,N_3092);
or U3512 (N_3512,N_3326,N_3379);
or U3513 (N_3513,N_3082,N_3195);
nor U3514 (N_3514,N_3488,N_3059);
xnor U3515 (N_3515,N_3430,N_3482);
nand U3516 (N_3516,N_3064,N_3312);
and U3517 (N_3517,N_3018,N_3002);
nor U3518 (N_3518,N_3220,N_3039);
nor U3519 (N_3519,N_3143,N_3134);
nand U3520 (N_3520,N_3232,N_3267);
or U3521 (N_3521,N_3419,N_3056);
or U3522 (N_3522,N_3199,N_3159);
or U3523 (N_3523,N_3223,N_3499);
or U3524 (N_3524,N_3112,N_3071);
nor U3525 (N_3525,N_3114,N_3395);
or U3526 (N_3526,N_3275,N_3226);
nor U3527 (N_3527,N_3066,N_3036);
nand U3528 (N_3528,N_3089,N_3392);
xor U3529 (N_3529,N_3200,N_3411);
and U3530 (N_3530,N_3405,N_3054);
and U3531 (N_3531,N_3487,N_3048);
or U3532 (N_3532,N_3127,N_3407);
nand U3533 (N_3533,N_3495,N_3123);
or U3534 (N_3534,N_3128,N_3148);
or U3535 (N_3535,N_3179,N_3306);
nor U3536 (N_3536,N_3185,N_3260);
nand U3537 (N_3537,N_3025,N_3435);
xor U3538 (N_3538,N_3484,N_3279);
xor U3539 (N_3539,N_3063,N_3243);
nand U3540 (N_3540,N_3498,N_3027);
nand U3541 (N_3541,N_3087,N_3230);
and U3542 (N_3542,N_3021,N_3207);
nor U3543 (N_3543,N_3055,N_3351);
xnor U3544 (N_3544,N_3225,N_3014);
xnor U3545 (N_3545,N_3022,N_3409);
xnor U3546 (N_3546,N_3162,N_3080);
nand U3547 (N_3547,N_3007,N_3410);
nand U3548 (N_3548,N_3081,N_3190);
nor U3549 (N_3549,N_3035,N_3341);
xnor U3550 (N_3550,N_3170,N_3428);
nand U3551 (N_3551,N_3247,N_3286);
and U3552 (N_3552,N_3367,N_3318);
xor U3553 (N_3553,N_3203,N_3360);
or U3554 (N_3554,N_3145,N_3390);
nand U3555 (N_3555,N_3072,N_3213);
and U3556 (N_3556,N_3288,N_3024);
and U3557 (N_3557,N_3103,N_3317);
and U3558 (N_3558,N_3211,N_3294);
or U3559 (N_3559,N_3142,N_3403);
xnor U3560 (N_3560,N_3141,N_3216);
nand U3561 (N_3561,N_3358,N_3383);
xor U3562 (N_3562,N_3091,N_3344);
nand U3563 (N_3563,N_3239,N_3308);
nand U3564 (N_3564,N_3172,N_3368);
or U3565 (N_3565,N_3292,N_3125);
nor U3566 (N_3566,N_3010,N_3214);
or U3567 (N_3567,N_3437,N_3273);
nor U3568 (N_3568,N_3377,N_3444);
xor U3569 (N_3569,N_3062,N_3233);
nand U3570 (N_3570,N_3309,N_3122);
nand U3571 (N_3571,N_3468,N_3321);
nand U3572 (N_3572,N_3212,N_3353);
nand U3573 (N_3573,N_3492,N_3139);
nor U3574 (N_3574,N_3478,N_3238);
nand U3575 (N_3575,N_3003,N_3310);
nor U3576 (N_3576,N_3155,N_3315);
and U3577 (N_3577,N_3262,N_3337);
and U3578 (N_3578,N_3381,N_3389);
and U3579 (N_3579,N_3252,N_3327);
xnor U3580 (N_3580,N_3398,N_3400);
xnor U3581 (N_3581,N_3278,N_3263);
and U3582 (N_3582,N_3343,N_3158);
xor U3583 (N_3583,N_3303,N_3457);
or U3584 (N_3584,N_3277,N_3355);
nand U3585 (N_3585,N_3030,N_3194);
or U3586 (N_3586,N_3181,N_3284);
nand U3587 (N_3587,N_3470,N_3259);
or U3588 (N_3588,N_3058,N_3100);
nand U3589 (N_3589,N_3193,N_3297);
nand U3590 (N_3590,N_3333,N_3204);
xnor U3591 (N_3591,N_3493,N_3462);
nand U3592 (N_3592,N_3053,N_3023);
or U3593 (N_3593,N_3102,N_3329);
xnor U3594 (N_3594,N_3156,N_3130);
nand U3595 (N_3595,N_3174,N_3032);
xnor U3596 (N_3596,N_3154,N_3034);
or U3597 (N_3597,N_3241,N_3157);
nor U3598 (N_3598,N_3222,N_3300);
xor U3599 (N_3599,N_3219,N_3440);
and U3600 (N_3600,N_3146,N_3209);
nor U3601 (N_3601,N_3388,N_3132);
or U3602 (N_3602,N_3264,N_3319);
xor U3603 (N_3603,N_3422,N_3116);
or U3604 (N_3604,N_3004,N_3339);
or U3605 (N_3605,N_3373,N_3402);
nand U3606 (N_3606,N_3009,N_3332);
or U3607 (N_3607,N_3480,N_3370);
and U3608 (N_3608,N_3113,N_3236);
and U3609 (N_3609,N_3393,N_3095);
and U3610 (N_3610,N_3496,N_3295);
nor U3611 (N_3611,N_3497,N_3131);
nor U3612 (N_3612,N_3334,N_3245);
nand U3613 (N_3613,N_3117,N_3051);
xnor U3614 (N_3614,N_3472,N_3285);
or U3615 (N_3615,N_3429,N_3320);
and U3616 (N_3616,N_3192,N_3372);
nor U3617 (N_3617,N_3399,N_3396);
or U3618 (N_3618,N_3369,N_3012);
and U3619 (N_3619,N_3182,N_3414);
xnor U3620 (N_3620,N_3107,N_3140);
or U3621 (N_3621,N_3382,N_3234);
nand U3622 (N_3622,N_3331,N_3293);
or U3623 (N_3623,N_3153,N_3208);
xor U3624 (N_3624,N_3042,N_3198);
or U3625 (N_3625,N_3265,N_3416);
xnor U3626 (N_3626,N_3347,N_3442);
nor U3627 (N_3627,N_3166,N_3129);
xnor U3628 (N_3628,N_3160,N_3120);
nand U3629 (N_3629,N_3481,N_3137);
or U3630 (N_3630,N_3126,N_3350);
and U3631 (N_3631,N_3261,N_3178);
or U3632 (N_3632,N_3224,N_3272);
or U3633 (N_3633,N_3291,N_3463);
nor U3634 (N_3634,N_3426,N_3366);
and U3635 (N_3635,N_3412,N_3362);
nor U3636 (N_3636,N_3434,N_3460);
nand U3637 (N_3637,N_3423,N_3184);
and U3638 (N_3638,N_3201,N_3057);
and U3639 (N_3639,N_3401,N_3096);
nand U3640 (N_3640,N_3387,N_3016);
nand U3641 (N_3641,N_3380,N_3256);
or U3642 (N_3642,N_3026,N_3099);
or U3643 (N_3643,N_3356,N_3384);
or U3644 (N_3644,N_3283,N_3322);
nor U3645 (N_3645,N_3276,N_3404);
nor U3646 (N_3646,N_3485,N_3271);
nor U3647 (N_3647,N_3266,N_3421);
nand U3648 (N_3648,N_3255,N_3231);
xor U3649 (N_3649,N_3307,N_3237);
and U3650 (N_3650,N_3287,N_3342);
xor U3651 (N_3651,N_3374,N_3391);
nand U3652 (N_3652,N_3450,N_3186);
nor U3653 (N_3653,N_3065,N_3073);
and U3654 (N_3654,N_3152,N_3378);
xnor U3655 (N_3655,N_3475,N_3135);
nor U3656 (N_3656,N_3467,N_3465);
nor U3657 (N_3657,N_3354,N_3469);
and U3658 (N_3658,N_3486,N_3385);
or U3659 (N_3659,N_3202,N_3316);
or U3660 (N_3660,N_3005,N_3169);
nand U3661 (N_3661,N_3340,N_3408);
or U3662 (N_3662,N_3298,N_3477);
and U3663 (N_3663,N_3349,N_3070);
nand U3664 (N_3664,N_3364,N_3033);
nor U3665 (N_3665,N_3289,N_3168);
and U3666 (N_3666,N_3397,N_3443);
and U3667 (N_3667,N_3215,N_3150);
and U3668 (N_3668,N_3413,N_3138);
nor U3669 (N_3669,N_3453,N_3249);
xnor U3670 (N_3670,N_3253,N_3031);
nand U3671 (N_3671,N_3109,N_3013);
nand U3672 (N_3672,N_3175,N_3282);
and U3673 (N_3673,N_3136,N_3494);
and U3674 (N_3674,N_3346,N_3449);
nand U3675 (N_3675,N_3479,N_3177);
xnor U3676 (N_3676,N_3311,N_3459);
or U3677 (N_3677,N_3270,N_3115);
nand U3678 (N_3678,N_3432,N_3229);
nand U3679 (N_3679,N_3084,N_3455);
nor U3680 (N_3680,N_3197,N_3000);
nand U3681 (N_3681,N_3328,N_3029);
or U3682 (N_3682,N_3006,N_3043);
nor U3683 (N_3683,N_3098,N_3094);
xnor U3684 (N_3684,N_3205,N_3313);
and U3685 (N_3685,N_3376,N_3436);
or U3686 (N_3686,N_3068,N_3217);
xor U3687 (N_3687,N_3425,N_3188);
nand U3688 (N_3688,N_3218,N_3330);
nor U3689 (N_3689,N_3418,N_3304);
or U3690 (N_3690,N_3290,N_3471);
and U3691 (N_3691,N_3491,N_3083);
or U3692 (N_3692,N_3301,N_3020);
nand U3693 (N_3693,N_3335,N_3452);
or U3694 (N_3694,N_3076,N_3187);
xor U3695 (N_3695,N_3456,N_3281);
nand U3696 (N_3696,N_3086,N_3075);
nand U3697 (N_3697,N_3446,N_3119);
and U3698 (N_3698,N_3015,N_3067);
nor U3699 (N_3699,N_3438,N_3314);
nand U3700 (N_3700,N_3163,N_3483);
xor U3701 (N_3701,N_3250,N_3206);
nand U3702 (N_3702,N_3359,N_3133);
nor U3703 (N_3703,N_3077,N_3101);
nand U3704 (N_3704,N_3302,N_3108);
or U3705 (N_3705,N_3427,N_3124);
and U3706 (N_3706,N_3069,N_3268);
nand U3707 (N_3707,N_3149,N_3257);
or U3708 (N_3708,N_3451,N_3448);
nand U3709 (N_3709,N_3191,N_3041);
and U3710 (N_3710,N_3176,N_3061);
xor U3711 (N_3711,N_3454,N_3111);
or U3712 (N_3712,N_3164,N_3420);
nand U3713 (N_3713,N_3049,N_3441);
or U3714 (N_3714,N_3248,N_3280);
nor U3715 (N_3715,N_3431,N_3090);
nor U3716 (N_3716,N_3345,N_3336);
or U3717 (N_3717,N_3037,N_3251);
xor U3718 (N_3718,N_3348,N_3375);
or U3719 (N_3719,N_3489,N_3180);
nand U3720 (N_3720,N_3183,N_3361);
nand U3721 (N_3721,N_3147,N_3196);
or U3722 (N_3722,N_3001,N_3110);
xor U3723 (N_3723,N_3474,N_3417);
and U3724 (N_3724,N_3121,N_3104);
and U3725 (N_3725,N_3338,N_3235);
xor U3726 (N_3726,N_3047,N_3461);
nand U3727 (N_3727,N_3118,N_3167);
nand U3728 (N_3728,N_3363,N_3171);
or U3729 (N_3729,N_3105,N_3254);
or U3730 (N_3730,N_3371,N_3046);
or U3731 (N_3731,N_3097,N_3017);
nand U3732 (N_3732,N_3221,N_3144);
nand U3733 (N_3733,N_3011,N_3394);
and U3734 (N_3734,N_3052,N_3323);
nor U3735 (N_3735,N_3490,N_3019);
xnor U3736 (N_3736,N_3189,N_3093);
xnor U3737 (N_3737,N_3106,N_3244);
or U3738 (N_3738,N_3433,N_3078);
nand U3739 (N_3739,N_3445,N_3060);
or U3740 (N_3740,N_3296,N_3447);
nand U3741 (N_3741,N_3151,N_3074);
and U3742 (N_3742,N_3386,N_3228);
nand U3743 (N_3743,N_3269,N_3458);
or U3744 (N_3744,N_3088,N_3473);
or U3745 (N_3745,N_3476,N_3466);
nor U3746 (N_3746,N_3258,N_3406);
or U3747 (N_3747,N_3085,N_3028);
nor U3748 (N_3748,N_3040,N_3439);
xnor U3749 (N_3749,N_3038,N_3464);
or U3750 (N_3750,N_3132,N_3131);
nor U3751 (N_3751,N_3301,N_3037);
and U3752 (N_3752,N_3253,N_3330);
and U3753 (N_3753,N_3370,N_3139);
xnor U3754 (N_3754,N_3389,N_3179);
nor U3755 (N_3755,N_3011,N_3225);
and U3756 (N_3756,N_3486,N_3147);
nand U3757 (N_3757,N_3229,N_3235);
nand U3758 (N_3758,N_3457,N_3171);
and U3759 (N_3759,N_3236,N_3478);
or U3760 (N_3760,N_3278,N_3143);
nor U3761 (N_3761,N_3206,N_3418);
xor U3762 (N_3762,N_3103,N_3005);
nand U3763 (N_3763,N_3390,N_3444);
nand U3764 (N_3764,N_3425,N_3228);
and U3765 (N_3765,N_3194,N_3350);
or U3766 (N_3766,N_3039,N_3036);
xnor U3767 (N_3767,N_3241,N_3205);
or U3768 (N_3768,N_3037,N_3016);
or U3769 (N_3769,N_3077,N_3211);
and U3770 (N_3770,N_3134,N_3357);
and U3771 (N_3771,N_3097,N_3463);
and U3772 (N_3772,N_3298,N_3311);
xor U3773 (N_3773,N_3308,N_3161);
nand U3774 (N_3774,N_3001,N_3222);
or U3775 (N_3775,N_3378,N_3048);
or U3776 (N_3776,N_3215,N_3236);
nand U3777 (N_3777,N_3056,N_3456);
and U3778 (N_3778,N_3014,N_3135);
xor U3779 (N_3779,N_3162,N_3200);
xnor U3780 (N_3780,N_3056,N_3477);
nand U3781 (N_3781,N_3173,N_3201);
or U3782 (N_3782,N_3151,N_3139);
nand U3783 (N_3783,N_3243,N_3343);
nor U3784 (N_3784,N_3059,N_3259);
nand U3785 (N_3785,N_3384,N_3060);
nand U3786 (N_3786,N_3370,N_3172);
and U3787 (N_3787,N_3266,N_3390);
xor U3788 (N_3788,N_3420,N_3272);
nor U3789 (N_3789,N_3034,N_3242);
xor U3790 (N_3790,N_3065,N_3415);
xor U3791 (N_3791,N_3276,N_3281);
and U3792 (N_3792,N_3010,N_3471);
nor U3793 (N_3793,N_3041,N_3046);
nand U3794 (N_3794,N_3039,N_3191);
nor U3795 (N_3795,N_3173,N_3056);
nand U3796 (N_3796,N_3012,N_3466);
nand U3797 (N_3797,N_3125,N_3397);
nand U3798 (N_3798,N_3175,N_3459);
and U3799 (N_3799,N_3254,N_3094);
nor U3800 (N_3800,N_3198,N_3140);
xor U3801 (N_3801,N_3427,N_3434);
nor U3802 (N_3802,N_3338,N_3185);
nand U3803 (N_3803,N_3168,N_3434);
or U3804 (N_3804,N_3269,N_3190);
nor U3805 (N_3805,N_3428,N_3306);
and U3806 (N_3806,N_3174,N_3030);
nor U3807 (N_3807,N_3454,N_3260);
nor U3808 (N_3808,N_3121,N_3245);
nor U3809 (N_3809,N_3437,N_3448);
and U3810 (N_3810,N_3010,N_3479);
xnor U3811 (N_3811,N_3135,N_3175);
xor U3812 (N_3812,N_3271,N_3336);
or U3813 (N_3813,N_3441,N_3269);
and U3814 (N_3814,N_3374,N_3253);
xor U3815 (N_3815,N_3002,N_3168);
nor U3816 (N_3816,N_3021,N_3294);
xnor U3817 (N_3817,N_3064,N_3077);
nand U3818 (N_3818,N_3258,N_3387);
xor U3819 (N_3819,N_3222,N_3210);
xnor U3820 (N_3820,N_3020,N_3448);
nor U3821 (N_3821,N_3346,N_3486);
or U3822 (N_3822,N_3318,N_3269);
or U3823 (N_3823,N_3143,N_3238);
xor U3824 (N_3824,N_3405,N_3166);
nor U3825 (N_3825,N_3443,N_3007);
nor U3826 (N_3826,N_3462,N_3323);
nor U3827 (N_3827,N_3181,N_3319);
or U3828 (N_3828,N_3137,N_3388);
and U3829 (N_3829,N_3348,N_3100);
xor U3830 (N_3830,N_3069,N_3149);
and U3831 (N_3831,N_3106,N_3194);
or U3832 (N_3832,N_3128,N_3256);
and U3833 (N_3833,N_3322,N_3356);
nand U3834 (N_3834,N_3051,N_3287);
nor U3835 (N_3835,N_3266,N_3294);
xor U3836 (N_3836,N_3429,N_3239);
and U3837 (N_3837,N_3368,N_3112);
and U3838 (N_3838,N_3085,N_3319);
nor U3839 (N_3839,N_3263,N_3455);
nand U3840 (N_3840,N_3167,N_3232);
or U3841 (N_3841,N_3468,N_3151);
and U3842 (N_3842,N_3148,N_3375);
nor U3843 (N_3843,N_3286,N_3079);
nand U3844 (N_3844,N_3366,N_3090);
or U3845 (N_3845,N_3063,N_3431);
and U3846 (N_3846,N_3342,N_3138);
or U3847 (N_3847,N_3345,N_3379);
nand U3848 (N_3848,N_3015,N_3470);
nand U3849 (N_3849,N_3353,N_3149);
and U3850 (N_3850,N_3480,N_3067);
or U3851 (N_3851,N_3054,N_3446);
and U3852 (N_3852,N_3205,N_3038);
nand U3853 (N_3853,N_3339,N_3452);
xnor U3854 (N_3854,N_3381,N_3028);
and U3855 (N_3855,N_3457,N_3086);
and U3856 (N_3856,N_3219,N_3458);
nand U3857 (N_3857,N_3482,N_3292);
nand U3858 (N_3858,N_3217,N_3048);
and U3859 (N_3859,N_3380,N_3277);
or U3860 (N_3860,N_3191,N_3030);
or U3861 (N_3861,N_3479,N_3404);
nor U3862 (N_3862,N_3441,N_3147);
nand U3863 (N_3863,N_3183,N_3200);
xnor U3864 (N_3864,N_3141,N_3439);
nor U3865 (N_3865,N_3285,N_3314);
or U3866 (N_3866,N_3163,N_3449);
nor U3867 (N_3867,N_3351,N_3118);
or U3868 (N_3868,N_3206,N_3139);
and U3869 (N_3869,N_3490,N_3301);
or U3870 (N_3870,N_3393,N_3087);
nor U3871 (N_3871,N_3286,N_3425);
or U3872 (N_3872,N_3069,N_3189);
nand U3873 (N_3873,N_3138,N_3246);
nor U3874 (N_3874,N_3370,N_3416);
nor U3875 (N_3875,N_3074,N_3463);
and U3876 (N_3876,N_3008,N_3267);
nand U3877 (N_3877,N_3306,N_3432);
or U3878 (N_3878,N_3387,N_3211);
xor U3879 (N_3879,N_3458,N_3196);
and U3880 (N_3880,N_3040,N_3443);
or U3881 (N_3881,N_3359,N_3228);
nand U3882 (N_3882,N_3105,N_3499);
nor U3883 (N_3883,N_3115,N_3372);
and U3884 (N_3884,N_3240,N_3462);
xnor U3885 (N_3885,N_3495,N_3382);
and U3886 (N_3886,N_3153,N_3012);
xnor U3887 (N_3887,N_3045,N_3164);
nor U3888 (N_3888,N_3046,N_3293);
xnor U3889 (N_3889,N_3266,N_3152);
and U3890 (N_3890,N_3343,N_3088);
xnor U3891 (N_3891,N_3315,N_3353);
and U3892 (N_3892,N_3360,N_3399);
nand U3893 (N_3893,N_3338,N_3116);
nand U3894 (N_3894,N_3312,N_3342);
nor U3895 (N_3895,N_3414,N_3099);
xor U3896 (N_3896,N_3459,N_3105);
or U3897 (N_3897,N_3191,N_3306);
nand U3898 (N_3898,N_3053,N_3389);
nor U3899 (N_3899,N_3175,N_3482);
and U3900 (N_3900,N_3162,N_3248);
or U3901 (N_3901,N_3434,N_3377);
nor U3902 (N_3902,N_3182,N_3194);
and U3903 (N_3903,N_3382,N_3473);
or U3904 (N_3904,N_3001,N_3077);
nor U3905 (N_3905,N_3331,N_3123);
nand U3906 (N_3906,N_3214,N_3470);
nor U3907 (N_3907,N_3134,N_3495);
and U3908 (N_3908,N_3005,N_3079);
and U3909 (N_3909,N_3179,N_3387);
nor U3910 (N_3910,N_3392,N_3005);
or U3911 (N_3911,N_3140,N_3370);
nand U3912 (N_3912,N_3204,N_3300);
nor U3913 (N_3913,N_3470,N_3183);
and U3914 (N_3914,N_3191,N_3264);
or U3915 (N_3915,N_3444,N_3461);
or U3916 (N_3916,N_3444,N_3202);
xor U3917 (N_3917,N_3492,N_3177);
nand U3918 (N_3918,N_3058,N_3458);
xnor U3919 (N_3919,N_3491,N_3013);
nand U3920 (N_3920,N_3377,N_3335);
xnor U3921 (N_3921,N_3329,N_3012);
nor U3922 (N_3922,N_3309,N_3107);
nor U3923 (N_3923,N_3016,N_3334);
and U3924 (N_3924,N_3068,N_3266);
nor U3925 (N_3925,N_3338,N_3395);
nor U3926 (N_3926,N_3323,N_3376);
xor U3927 (N_3927,N_3402,N_3103);
or U3928 (N_3928,N_3144,N_3006);
or U3929 (N_3929,N_3332,N_3284);
xnor U3930 (N_3930,N_3005,N_3019);
nor U3931 (N_3931,N_3190,N_3060);
nand U3932 (N_3932,N_3042,N_3260);
nor U3933 (N_3933,N_3040,N_3321);
nand U3934 (N_3934,N_3436,N_3027);
xor U3935 (N_3935,N_3385,N_3430);
and U3936 (N_3936,N_3032,N_3413);
or U3937 (N_3937,N_3389,N_3471);
or U3938 (N_3938,N_3095,N_3083);
nand U3939 (N_3939,N_3081,N_3368);
xor U3940 (N_3940,N_3338,N_3253);
and U3941 (N_3941,N_3103,N_3408);
or U3942 (N_3942,N_3462,N_3439);
and U3943 (N_3943,N_3265,N_3104);
or U3944 (N_3944,N_3339,N_3381);
nor U3945 (N_3945,N_3113,N_3337);
and U3946 (N_3946,N_3298,N_3182);
nand U3947 (N_3947,N_3186,N_3486);
or U3948 (N_3948,N_3258,N_3020);
nand U3949 (N_3949,N_3124,N_3311);
xnor U3950 (N_3950,N_3312,N_3166);
nor U3951 (N_3951,N_3116,N_3084);
nand U3952 (N_3952,N_3162,N_3326);
nor U3953 (N_3953,N_3423,N_3280);
nand U3954 (N_3954,N_3240,N_3122);
nor U3955 (N_3955,N_3189,N_3475);
nor U3956 (N_3956,N_3047,N_3280);
and U3957 (N_3957,N_3259,N_3076);
nor U3958 (N_3958,N_3420,N_3044);
or U3959 (N_3959,N_3174,N_3088);
or U3960 (N_3960,N_3449,N_3379);
and U3961 (N_3961,N_3346,N_3423);
nor U3962 (N_3962,N_3462,N_3023);
nand U3963 (N_3963,N_3400,N_3068);
or U3964 (N_3964,N_3205,N_3181);
and U3965 (N_3965,N_3194,N_3165);
or U3966 (N_3966,N_3211,N_3436);
nand U3967 (N_3967,N_3447,N_3360);
nand U3968 (N_3968,N_3146,N_3238);
or U3969 (N_3969,N_3175,N_3327);
and U3970 (N_3970,N_3353,N_3013);
and U3971 (N_3971,N_3264,N_3188);
nand U3972 (N_3972,N_3191,N_3261);
or U3973 (N_3973,N_3075,N_3437);
and U3974 (N_3974,N_3072,N_3437);
nand U3975 (N_3975,N_3108,N_3283);
nor U3976 (N_3976,N_3473,N_3086);
nor U3977 (N_3977,N_3331,N_3358);
xor U3978 (N_3978,N_3280,N_3050);
and U3979 (N_3979,N_3412,N_3104);
and U3980 (N_3980,N_3131,N_3113);
and U3981 (N_3981,N_3053,N_3222);
nand U3982 (N_3982,N_3457,N_3261);
xnor U3983 (N_3983,N_3396,N_3429);
nand U3984 (N_3984,N_3325,N_3489);
or U3985 (N_3985,N_3421,N_3074);
and U3986 (N_3986,N_3024,N_3059);
xor U3987 (N_3987,N_3103,N_3172);
nand U3988 (N_3988,N_3200,N_3314);
nand U3989 (N_3989,N_3443,N_3171);
xnor U3990 (N_3990,N_3114,N_3249);
or U3991 (N_3991,N_3249,N_3372);
xnor U3992 (N_3992,N_3128,N_3168);
nor U3993 (N_3993,N_3464,N_3186);
nor U3994 (N_3994,N_3014,N_3115);
nand U3995 (N_3995,N_3271,N_3030);
and U3996 (N_3996,N_3204,N_3356);
nor U3997 (N_3997,N_3443,N_3325);
and U3998 (N_3998,N_3413,N_3068);
nor U3999 (N_3999,N_3393,N_3136);
and U4000 (N_4000,N_3515,N_3919);
nand U4001 (N_4001,N_3845,N_3668);
nand U4002 (N_4002,N_3976,N_3673);
nor U4003 (N_4003,N_3697,N_3662);
nor U4004 (N_4004,N_3785,N_3548);
nor U4005 (N_4005,N_3941,N_3572);
nor U4006 (N_4006,N_3539,N_3852);
or U4007 (N_4007,N_3898,N_3883);
xnor U4008 (N_4008,N_3937,N_3911);
or U4009 (N_4009,N_3925,N_3765);
nor U4010 (N_4010,N_3886,N_3955);
or U4011 (N_4011,N_3996,N_3602);
nor U4012 (N_4012,N_3866,N_3906);
or U4013 (N_4013,N_3727,N_3653);
xor U4014 (N_4014,N_3603,N_3899);
nand U4015 (N_4015,N_3848,N_3527);
nand U4016 (N_4016,N_3679,N_3760);
or U4017 (N_4017,N_3592,N_3728);
xor U4018 (N_4018,N_3874,N_3618);
or U4019 (N_4019,N_3676,N_3908);
or U4020 (N_4020,N_3770,N_3549);
and U4021 (N_4021,N_3702,N_3892);
nor U4022 (N_4022,N_3701,N_3684);
nand U4023 (N_4023,N_3950,N_3751);
and U4024 (N_4024,N_3945,N_3951);
or U4025 (N_4025,N_3789,N_3761);
nor U4026 (N_4026,N_3514,N_3520);
xnor U4027 (N_4027,N_3881,N_3759);
xnor U4028 (N_4028,N_3887,N_3717);
nand U4029 (N_4029,N_3862,N_3777);
or U4030 (N_4030,N_3624,N_3553);
nand U4031 (N_4031,N_3640,N_3667);
xor U4032 (N_4032,N_3860,N_3696);
nor U4033 (N_4033,N_3725,N_3829);
and U4034 (N_4034,N_3677,N_3913);
xor U4035 (N_4035,N_3985,N_3735);
nand U4036 (N_4036,N_3693,N_3509);
and U4037 (N_4037,N_3896,N_3987);
and U4038 (N_4038,N_3871,N_3587);
nand U4039 (N_4039,N_3629,N_3580);
and U4040 (N_4040,N_3816,N_3972);
nor U4041 (N_4041,N_3828,N_3570);
or U4042 (N_4042,N_3819,N_3656);
nor U4043 (N_4043,N_3821,N_3695);
nand U4044 (N_4044,N_3722,N_3512);
nor U4045 (N_4045,N_3675,N_3861);
xor U4046 (N_4046,N_3902,N_3754);
nor U4047 (N_4047,N_3646,N_3894);
or U4048 (N_4048,N_3960,N_3973);
and U4049 (N_4049,N_3655,N_3686);
nand U4050 (N_4050,N_3918,N_3975);
nand U4051 (N_4051,N_3837,N_3589);
xor U4052 (N_4052,N_3564,N_3762);
xor U4053 (N_4053,N_3547,N_3538);
xnor U4054 (N_4054,N_3663,N_3752);
or U4055 (N_4055,N_3801,N_3521);
and U4056 (N_4056,N_3631,N_3584);
xnor U4057 (N_4057,N_3875,N_3511);
xor U4058 (N_4058,N_3809,N_3659);
or U4059 (N_4059,N_3614,N_3510);
nor U4060 (N_4060,N_3968,N_3596);
xor U4061 (N_4061,N_3814,N_3608);
nand U4062 (N_4062,N_3648,N_3573);
nand U4063 (N_4063,N_3555,N_3732);
nor U4064 (N_4064,N_3786,N_3857);
or U4065 (N_4065,N_3856,N_3745);
and U4066 (N_4066,N_3713,N_3997);
nand U4067 (N_4067,N_3999,N_3737);
or U4068 (N_4068,N_3981,N_3849);
nor U4069 (N_4069,N_3827,N_3711);
nand U4070 (N_4070,N_3681,N_3634);
xor U4071 (N_4071,N_3712,N_3811);
and U4072 (N_4072,N_3780,N_3787);
nor U4073 (N_4073,N_3867,N_3579);
nand U4074 (N_4074,N_3726,N_3595);
nand U4075 (N_4075,N_3869,N_3800);
and U4076 (N_4076,N_3773,N_3774);
and U4077 (N_4077,N_3680,N_3844);
and U4078 (N_4078,N_3674,N_3891);
or U4079 (N_4079,N_3971,N_3781);
nand U4080 (N_4080,N_3628,N_3805);
nor U4081 (N_4081,N_3615,N_3958);
nand U4082 (N_4082,N_3657,N_3836);
and U4083 (N_4083,N_3823,N_3638);
xor U4084 (N_4084,N_3994,N_3565);
xor U4085 (N_4085,N_3914,N_3907);
nor U4086 (N_4086,N_3873,N_3879);
and U4087 (N_4087,N_3991,N_3636);
nor U4088 (N_4088,N_3778,N_3692);
and U4089 (N_4089,N_3621,N_3854);
or U4090 (N_4090,N_3792,N_3930);
nand U4091 (N_4091,N_3698,N_3915);
xnor U4092 (N_4092,N_3591,N_3586);
nor U4093 (N_4093,N_3834,N_3649);
and U4094 (N_4094,N_3885,N_3897);
or U4095 (N_4095,N_3808,N_3588);
nor U4096 (N_4096,N_3784,N_3912);
and U4097 (N_4097,N_3526,N_3948);
and U4098 (N_4098,N_3716,N_3544);
nand U4099 (N_4099,N_3926,N_3790);
xnor U4100 (N_4100,N_3576,N_3750);
and U4101 (N_4101,N_3893,N_3768);
nor U4102 (N_4102,N_3904,N_3536);
xor U4103 (N_4103,N_3884,N_3705);
xnor U4104 (N_4104,N_3643,N_3597);
xnor U4105 (N_4105,N_3590,N_3661);
or U4106 (N_4106,N_3970,N_3859);
nand U4107 (N_4107,N_3583,N_3870);
or U4108 (N_4108,N_3707,N_3942);
or U4109 (N_4109,N_3952,N_3910);
nand U4110 (N_4110,N_3822,N_3660);
and U4111 (N_4111,N_3833,N_3704);
and U4112 (N_4112,N_3804,N_3949);
xor U4113 (N_4113,N_3607,N_3645);
nand U4114 (N_4114,N_3637,N_3741);
xor U4115 (N_4115,N_3531,N_3835);
nand U4116 (N_4116,N_3766,N_3546);
and U4117 (N_4117,N_3715,N_3518);
or U4118 (N_4118,N_3775,N_3807);
or U4119 (N_4119,N_3795,N_3530);
xor U4120 (N_4120,N_3933,N_3909);
or U4121 (N_4121,N_3689,N_3936);
and U4122 (N_4122,N_3932,N_3609);
nor U4123 (N_4123,N_3758,N_3505);
xor U4124 (N_4124,N_3700,N_3502);
nand U4125 (N_4125,N_3810,N_3938);
xor U4126 (N_4126,N_3946,N_3563);
and U4127 (N_4127,N_3944,N_3923);
or U4128 (N_4128,N_3788,N_3642);
or U4129 (N_4129,N_3961,N_3578);
or U4130 (N_4130,N_3665,N_3990);
nand U4131 (N_4131,N_3503,N_3855);
nand U4132 (N_4132,N_3714,N_3507);
nor U4133 (N_4133,N_3710,N_3687);
nor U4134 (N_4134,N_3666,N_3776);
xnor U4135 (N_4135,N_3622,N_3683);
nand U4136 (N_4136,N_3734,N_3703);
xnor U4137 (N_4137,N_3993,N_3880);
xnor U4138 (N_4138,N_3922,N_3995);
xor U4139 (N_4139,N_3953,N_3635);
xnor U4140 (N_4140,N_3935,N_3820);
nor U4141 (N_4141,N_3605,N_3756);
or U4142 (N_4142,N_3818,N_3783);
xnor U4143 (N_4143,N_3947,N_3838);
and U4144 (N_4144,N_3562,N_3980);
nor U4145 (N_4145,N_3610,N_3619);
nor U4146 (N_4146,N_3832,N_3506);
xnor U4147 (N_4147,N_3957,N_3920);
xnor U4148 (N_4148,N_3682,N_3504);
xor U4149 (N_4149,N_3793,N_3889);
xnor U4150 (N_4150,N_3543,N_3977);
nor U4151 (N_4151,N_3989,N_3688);
nor U4152 (N_4152,N_3966,N_3963);
xnor U4153 (N_4153,N_3841,N_3747);
nor U4154 (N_4154,N_3812,N_3513);
and U4155 (N_4155,N_3529,N_3552);
or U4156 (N_4156,N_3882,N_3699);
xor U4157 (N_4157,N_3651,N_3630);
nor U4158 (N_4158,N_3633,N_3559);
nand U4159 (N_4159,N_3877,N_3658);
or U4160 (N_4160,N_3690,N_3962);
and U4161 (N_4161,N_3940,N_3718);
nor U4162 (N_4162,N_3522,N_3931);
or U4163 (N_4163,N_3782,N_3895);
xnor U4164 (N_4164,N_3921,N_3998);
xnor U4165 (N_4165,N_3523,N_3802);
nand U4166 (N_4166,N_3569,N_3974);
nand U4167 (N_4167,N_3545,N_3575);
or U4168 (N_4168,N_3813,N_3669);
xor U4169 (N_4169,N_3979,N_3983);
and U4170 (N_4170,N_3508,N_3541);
or U4171 (N_4171,N_3967,N_3825);
nor U4172 (N_4172,N_3731,N_3817);
nor U4173 (N_4173,N_3561,N_3740);
nand U4174 (N_4174,N_3890,N_3678);
or U4175 (N_4175,N_3830,N_3796);
and U4176 (N_4176,N_3542,N_3525);
nor U4177 (N_4177,N_3582,N_3672);
nand U4178 (N_4178,N_3654,N_3599);
xor U4179 (N_4179,N_3650,N_3566);
nor U4180 (N_4180,N_3550,N_3738);
or U4181 (N_4181,N_3901,N_3872);
or U4182 (N_4182,N_3685,N_3927);
xor U4183 (N_4183,N_3558,N_3519);
and U4184 (N_4184,N_3964,N_3798);
nand U4185 (N_4185,N_3905,N_3535);
xnor U4186 (N_4186,N_3986,N_3719);
nand U4187 (N_4187,N_3557,N_3641);
nor U4188 (N_4188,N_3721,N_3749);
and U4189 (N_4189,N_3620,N_3917);
and U4190 (N_4190,N_3791,N_3755);
nor U4191 (N_4191,N_3992,N_3694);
or U4192 (N_4192,N_3956,N_3839);
nand U4193 (N_4193,N_3652,N_3533);
and U4194 (N_4194,N_3863,N_3815);
nand U4195 (N_4195,N_3551,N_3824);
or U4196 (N_4196,N_3724,N_3611);
xor U4197 (N_4197,N_3772,N_3803);
or U4198 (N_4198,N_3601,N_3623);
nor U4199 (N_4199,N_3744,N_3560);
nor U4200 (N_4200,N_3743,N_3831);
nand U4201 (N_4201,N_3556,N_3501);
nand U4202 (N_4202,N_3939,N_3988);
nand U4203 (N_4203,N_3846,N_3691);
xor U4204 (N_4204,N_3644,N_3928);
nor U4205 (N_4205,N_3500,N_3799);
nand U4206 (N_4206,N_3806,N_3581);
nand U4207 (N_4207,N_3929,N_3585);
nand U4208 (N_4208,N_3598,N_3534);
and U4209 (N_4209,N_3954,N_3826);
or U4210 (N_4210,N_3528,N_3733);
and U4211 (N_4211,N_3764,N_3612);
nand U4212 (N_4212,N_3916,N_3554);
nor U4213 (N_4213,N_3794,N_3606);
nor U4214 (N_4214,N_3568,N_3878);
and U4215 (N_4215,N_3736,N_3571);
nor U4216 (N_4216,N_3729,N_3709);
or U4217 (N_4217,N_3594,N_3626);
or U4218 (N_4218,N_3708,N_3969);
nor U4219 (N_4219,N_3524,N_3753);
and U4220 (N_4220,N_3842,N_3748);
and U4221 (N_4221,N_3616,N_3617);
xor U4222 (N_4222,N_3763,N_3532);
nand U4223 (N_4223,N_3742,N_3851);
nand U4224 (N_4224,N_3537,N_3982);
or U4225 (N_4225,N_3730,N_3876);
nor U4226 (N_4226,N_3664,N_3903);
nor U4227 (N_4227,N_3613,N_3577);
xor U4228 (N_4228,N_3868,N_3847);
nor U4229 (N_4229,N_3706,N_3934);
and U4230 (N_4230,N_3647,N_3965);
and U4231 (N_4231,N_3864,N_3767);
or U4232 (N_4232,N_3769,N_3720);
and U4233 (N_4233,N_3625,N_3779);
or U4234 (N_4234,N_3757,N_3739);
nor U4235 (N_4235,N_3540,N_3858);
and U4236 (N_4236,N_3670,N_3924);
and U4237 (N_4237,N_3771,N_3843);
and U4238 (N_4238,N_3639,N_3604);
or U4239 (N_4239,N_3517,N_3900);
nand U4240 (N_4240,N_3984,N_3850);
or U4241 (N_4241,N_3959,N_3746);
nor U4242 (N_4242,N_3840,N_3865);
and U4243 (N_4243,N_3600,N_3627);
xnor U4244 (N_4244,N_3567,N_3723);
or U4245 (N_4245,N_3888,N_3671);
and U4246 (N_4246,N_3978,N_3943);
nor U4247 (N_4247,N_3797,N_3574);
or U4248 (N_4248,N_3853,N_3593);
nand U4249 (N_4249,N_3516,N_3632);
xor U4250 (N_4250,N_3990,N_3944);
and U4251 (N_4251,N_3662,N_3689);
or U4252 (N_4252,N_3719,N_3876);
xnor U4253 (N_4253,N_3633,N_3843);
nor U4254 (N_4254,N_3906,N_3833);
xor U4255 (N_4255,N_3723,N_3514);
or U4256 (N_4256,N_3930,N_3587);
xor U4257 (N_4257,N_3995,N_3866);
and U4258 (N_4258,N_3625,N_3544);
nand U4259 (N_4259,N_3730,N_3528);
nor U4260 (N_4260,N_3701,N_3637);
nor U4261 (N_4261,N_3865,N_3989);
nand U4262 (N_4262,N_3695,N_3993);
xor U4263 (N_4263,N_3773,N_3868);
xnor U4264 (N_4264,N_3567,N_3720);
or U4265 (N_4265,N_3876,N_3676);
and U4266 (N_4266,N_3503,N_3520);
and U4267 (N_4267,N_3550,N_3722);
nand U4268 (N_4268,N_3964,N_3597);
xnor U4269 (N_4269,N_3652,N_3944);
or U4270 (N_4270,N_3562,N_3785);
xor U4271 (N_4271,N_3791,N_3885);
nand U4272 (N_4272,N_3767,N_3665);
xor U4273 (N_4273,N_3578,N_3528);
or U4274 (N_4274,N_3644,N_3545);
or U4275 (N_4275,N_3767,N_3534);
nand U4276 (N_4276,N_3913,N_3864);
and U4277 (N_4277,N_3981,N_3944);
nor U4278 (N_4278,N_3567,N_3844);
or U4279 (N_4279,N_3739,N_3825);
xnor U4280 (N_4280,N_3684,N_3760);
xor U4281 (N_4281,N_3977,N_3610);
and U4282 (N_4282,N_3969,N_3569);
or U4283 (N_4283,N_3941,N_3695);
nor U4284 (N_4284,N_3852,N_3506);
nor U4285 (N_4285,N_3909,N_3517);
and U4286 (N_4286,N_3894,N_3976);
and U4287 (N_4287,N_3870,N_3884);
xnor U4288 (N_4288,N_3912,N_3703);
xor U4289 (N_4289,N_3713,N_3758);
and U4290 (N_4290,N_3973,N_3573);
or U4291 (N_4291,N_3582,N_3890);
xnor U4292 (N_4292,N_3716,N_3736);
xor U4293 (N_4293,N_3985,N_3972);
and U4294 (N_4294,N_3612,N_3680);
nor U4295 (N_4295,N_3940,N_3830);
nand U4296 (N_4296,N_3651,N_3855);
or U4297 (N_4297,N_3783,N_3718);
nand U4298 (N_4298,N_3644,N_3572);
and U4299 (N_4299,N_3683,N_3635);
and U4300 (N_4300,N_3750,N_3842);
xnor U4301 (N_4301,N_3996,N_3582);
and U4302 (N_4302,N_3684,N_3538);
nand U4303 (N_4303,N_3929,N_3760);
and U4304 (N_4304,N_3585,N_3640);
nand U4305 (N_4305,N_3773,N_3864);
nand U4306 (N_4306,N_3576,N_3852);
nor U4307 (N_4307,N_3708,N_3554);
or U4308 (N_4308,N_3959,N_3674);
xnor U4309 (N_4309,N_3680,N_3533);
and U4310 (N_4310,N_3698,N_3594);
xnor U4311 (N_4311,N_3987,N_3852);
xnor U4312 (N_4312,N_3553,N_3606);
or U4313 (N_4313,N_3691,N_3898);
and U4314 (N_4314,N_3755,N_3515);
and U4315 (N_4315,N_3520,N_3729);
or U4316 (N_4316,N_3954,N_3980);
xnor U4317 (N_4317,N_3976,N_3659);
or U4318 (N_4318,N_3820,N_3665);
nor U4319 (N_4319,N_3774,N_3970);
or U4320 (N_4320,N_3901,N_3703);
and U4321 (N_4321,N_3851,N_3651);
nand U4322 (N_4322,N_3747,N_3670);
and U4323 (N_4323,N_3906,N_3776);
xnor U4324 (N_4324,N_3513,N_3885);
nor U4325 (N_4325,N_3665,N_3867);
nor U4326 (N_4326,N_3919,N_3826);
nand U4327 (N_4327,N_3513,N_3939);
and U4328 (N_4328,N_3610,N_3770);
nand U4329 (N_4329,N_3848,N_3947);
and U4330 (N_4330,N_3519,N_3586);
nand U4331 (N_4331,N_3881,N_3999);
and U4332 (N_4332,N_3640,N_3744);
xor U4333 (N_4333,N_3847,N_3980);
nand U4334 (N_4334,N_3592,N_3690);
nand U4335 (N_4335,N_3810,N_3898);
and U4336 (N_4336,N_3545,N_3893);
nand U4337 (N_4337,N_3802,N_3938);
xor U4338 (N_4338,N_3869,N_3602);
nor U4339 (N_4339,N_3894,N_3954);
and U4340 (N_4340,N_3987,N_3600);
xnor U4341 (N_4341,N_3961,N_3646);
nor U4342 (N_4342,N_3595,N_3618);
nor U4343 (N_4343,N_3823,N_3982);
xnor U4344 (N_4344,N_3967,N_3719);
nor U4345 (N_4345,N_3766,N_3652);
and U4346 (N_4346,N_3531,N_3766);
nand U4347 (N_4347,N_3729,N_3787);
nand U4348 (N_4348,N_3564,N_3506);
or U4349 (N_4349,N_3920,N_3975);
xor U4350 (N_4350,N_3890,N_3865);
nor U4351 (N_4351,N_3550,N_3533);
and U4352 (N_4352,N_3633,N_3611);
nand U4353 (N_4353,N_3705,N_3869);
and U4354 (N_4354,N_3532,N_3607);
and U4355 (N_4355,N_3544,N_3796);
xnor U4356 (N_4356,N_3677,N_3534);
xnor U4357 (N_4357,N_3937,N_3693);
nand U4358 (N_4358,N_3874,N_3898);
nand U4359 (N_4359,N_3879,N_3584);
and U4360 (N_4360,N_3804,N_3722);
nor U4361 (N_4361,N_3770,N_3628);
nor U4362 (N_4362,N_3694,N_3775);
nand U4363 (N_4363,N_3582,N_3799);
xnor U4364 (N_4364,N_3584,N_3852);
xnor U4365 (N_4365,N_3519,N_3709);
nor U4366 (N_4366,N_3885,N_3612);
xor U4367 (N_4367,N_3791,N_3720);
nand U4368 (N_4368,N_3854,N_3863);
xor U4369 (N_4369,N_3859,N_3769);
xnor U4370 (N_4370,N_3819,N_3511);
and U4371 (N_4371,N_3916,N_3899);
xor U4372 (N_4372,N_3915,N_3765);
nand U4373 (N_4373,N_3549,N_3984);
nand U4374 (N_4374,N_3592,N_3520);
nor U4375 (N_4375,N_3744,N_3678);
nand U4376 (N_4376,N_3540,N_3671);
or U4377 (N_4377,N_3684,N_3988);
xor U4378 (N_4378,N_3560,N_3648);
xor U4379 (N_4379,N_3953,N_3864);
nor U4380 (N_4380,N_3679,N_3601);
or U4381 (N_4381,N_3999,N_3948);
or U4382 (N_4382,N_3942,N_3787);
or U4383 (N_4383,N_3667,N_3627);
xor U4384 (N_4384,N_3840,N_3732);
and U4385 (N_4385,N_3632,N_3560);
nor U4386 (N_4386,N_3857,N_3813);
xor U4387 (N_4387,N_3524,N_3508);
xnor U4388 (N_4388,N_3781,N_3661);
nand U4389 (N_4389,N_3938,N_3897);
xor U4390 (N_4390,N_3552,N_3895);
nand U4391 (N_4391,N_3540,N_3885);
xor U4392 (N_4392,N_3796,N_3585);
and U4393 (N_4393,N_3571,N_3971);
nor U4394 (N_4394,N_3844,N_3838);
nor U4395 (N_4395,N_3694,N_3642);
nor U4396 (N_4396,N_3950,N_3822);
or U4397 (N_4397,N_3532,N_3511);
and U4398 (N_4398,N_3974,N_3724);
nor U4399 (N_4399,N_3816,N_3898);
nor U4400 (N_4400,N_3562,N_3846);
xnor U4401 (N_4401,N_3763,N_3573);
nor U4402 (N_4402,N_3944,N_3629);
nand U4403 (N_4403,N_3610,N_3574);
xnor U4404 (N_4404,N_3691,N_3840);
xnor U4405 (N_4405,N_3715,N_3663);
nand U4406 (N_4406,N_3515,N_3806);
nand U4407 (N_4407,N_3595,N_3517);
nand U4408 (N_4408,N_3649,N_3661);
nand U4409 (N_4409,N_3978,N_3764);
nand U4410 (N_4410,N_3603,N_3956);
nor U4411 (N_4411,N_3740,N_3543);
and U4412 (N_4412,N_3773,N_3691);
or U4413 (N_4413,N_3618,N_3540);
nor U4414 (N_4414,N_3874,N_3664);
xnor U4415 (N_4415,N_3827,N_3943);
nand U4416 (N_4416,N_3769,N_3791);
nand U4417 (N_4417,N_3942,N_3875);
nor U4418 (N_4418,N_3749,N_3736);
nand U4419 (N_4419,N_3516,N_3640);
nor U4420 (N_4420,N_3687,N_3973);
or U4421 (N_4421,N_3983,N_3883);
nand U4422 (N_4422,N_3952,N_3693);
or U4423 (N_4423,N_3650,N_3943);
nor U4424 (N_4424,N_3887,N_3713);
xor U4425 (N_4425,N_3970,N_3817);
or U4426 (N_4426,N_3539,N_3985);
and U4427 (N_4427,N_3725,N_3734);
nand U4428 (N_4428,N_3548,N_3829);
and U4429 (N_4429,N_3537,N_3572);
xor U4430 (N_4430,N_3702,N_3574);
xnor U4431 (N_4431,N_3535,N_3759);
xor U4432 (N_4432,N_3647,N_3762);
and U4433 (N_4433,N_3716,N_3650);
or U4434 (N_4434,N_3610,N_3551);
nand U4435 (N_4435,N_3939,N_3998);
xor U4436 (N_4436,N_3806,N_3918);
or U4437 (N_4437,N_3967,N_3686);
nor U4438 (N_4438,N_3757,N_3894);
nor U4439 (N_4439,N_3601,N_3611);
and U4440 (N_4440,N_3580,N_3622);
and U4441 (N_4441,N_3872,N_3891);
and U4442 (N_4442,N_3546,N_3731);
or U4443 (N_4443,N_3704,N_3791);
nor U4444 (N_4444,N_3925,N_3888);
or U4445 (N_4445,N_3697,N_3611);
xor U4446 (N_4446,N_3655,N_3875);
nand U4447 (N_4447,N_3916,N_3993);
nor U4448 (N_4448,N_3714,N_3619);
and U4449 (N_4449,N_3970,N_3650);
and U4450 (N_4450,N_3693,N_3855);
nand U4451 (N_4451,N_3991,N_3866);
nand U4452 (N_4452,N_3828,N_3729);
nor U4453 (N_4453,N_3847,N_3747);
and U4454 (N_4454,N_3550,N_3866);
nand U4455 (N_4455,N_3987,N_3689);
nand U4456 (N_4456,N_3667,N_3883);
or U4457 (N_4457,N_3653,N_3529);
and U4458 (N_4458,N_3917,N_3929);
or U4459 (N_4459,N_3919,N_3701);
xnor U4460 (N_4460,N_3551,N_3683);
or U4461 (N_4461,N_3903,N_3619);
xor U4462 (N_4462,N_3868,N_3841);
nand U4463 (N_4463,N_3797,N_3917);
or U4464 (N_4464,N_3502,N_3907);
and U4465 (N_4465,N_3985,N_3876);
nand U4466 (N_4466,N_3848,N_3661);
nor U4467 (N_4467,N_3987,N_3508);
or U4468 (N_4468,N_3796,N_3759);
xnor U4469 (N_4469,N_3991,N_3981);
and U4470 (N_4470,N_3978,N_3996);
and U4471 (N_4471,N_3617,N_3926);
or U4472 (N_4472,N_3734,N_3901);
xor U4473 (N_4473,N_3739,N_3751);
nor U4474 (N_4474,N_3843,N_3933);
xor U4475 (N_4475,N_3612,N_3893);
nor U4476 (N_4476,N_3993,N_3691);
nor U4477 (N_4477,N_3620,N_3864);
nand U4478 (N_4478,N_3850,N_3819);
and U4479 (N_4479,N_3819,N_3870);
xor U4480 (N_4480,N_3576,N_3932);
or U4481 (N_4481,N_3724,N_3950);
nand U4482 (N_4482,N_3558,N_3675);
or U4483 (N_4483,N_3519,N_3890);
and U4484 (N_4484,N_3597,N_3559);
nand U4485 (N_4485,N_3514,N_3888);
nand U4486 (N_4486,N_3624,N_3625);
or U4487 (N_4487,N_3991,N_3749);
nand U4488 (N_4488,N_3786,N_3982);
or U4489 (N_4489,N_3641,N_3519);
and U4490 (N_4490,N_3805,N_3959);
nor U4491 (N_4491,N_3562,N_3515);
and U4492 (N_4492,N_3985,N_3629);
xor U4493 (N_4493,N_3951,N_3918);
or U4494 (N_4494,N_3827,N_3834);
and U4495 (N_4495,N_3669,N_3584);
xnor U4496 (N_4496,N_3929,N_3895);
nand U4497 (N_4497,N_3701,N_3571);
or U4498 (N_4498,N_3678,N_3916);
xor U4499 (N_4499,N_3558,N_3986);
xor U4500 (N_4500,N_4036,N_4261);
xor U4501 (N_4501,N_4146,N_4395);
and U4502 (N_4502,N_4030,N_4228);
and U4503 (N_4503,N_4086,N_4488);
xnor U4504 (N_4504,N_4266,N_4298);
and U4505 (N_4505,N_4370,N_4346);
or U4506 (N_4506,N_4489,N_4429);
nor U4507 (N_4507,N_4384,N_4037);
or U4508 (N_4508,N_4348,N_4357);
nand U4509 (N_4509,N_4262,N_4144);
nand U4510 (N_4510,N_4226,N_4212);
and U4511 (N_4511,N_4284,N_4127);
xnor U4512 (N_4512,N_4031,N_4277);
or U4513 (N_4513,N_4453,N_4013);
and U4514 (N_4514,N_4499,N_4297);
nand U4515 (N_4515,N_4256,N_4007);
xnor U4516 (N_4516,N_4179,N_4314);
xor U4517 (N_4517,N_4047,N_4498);
xor U4518 (N_4518,N_4033,N_4342);
and U4519 (N_4519,N_4358,N_4095);
xor U4520 (N_4520,N_4046,N_4341);
or U4521 (N_4521,N_4123,N_4045);
or U4522 (N_4522,N_4374,N_4068);
nand U4523 (N_4523,N_4232,N_4274);
or U4524 (N_4524,N_4057,N_4294);
or U4525 (N_4525,N_4288,N_4476);
nand U4526 (N_4526,N_4029,N_4072);
nor U4527 (N_4527,N_4461,N_4243);
xor U4528 (N_4528,N_4247,N_4380);
nor U4529 (N_4529,N_4382,N_4272);
xor U4530 (N_4530,N_4215,N_4299);
or U4531 (N_4531,N_4147,N_4471);
and U4532 (N_4532,N_4111,N_4181);
nand U4533 (N_4533,N_4309,N_4002);
or U4534 (N_4534,N_4157,N_4385);
or U4535 (N_4535,N_4455,N_4333);
xor U4536 (N_4536,N_4242,N_4217);
and U4537 (N_4537,N_4438,N_4016);
and U4538 (N_4538,N_4252,N_4414);
nand U4539 (N_4539,N_4244,N_4041);
nor U4540 (N_4540,N_4233,N_4108);
xor U4541 (N_4541,N_4220,N_4185);
or U4542 (N_4542,N_4081,N_4319);
nand U4543 (N_4543,N_4257,N_4289);
xnor U4544 (N_4544,N_4209,N_4365);
xnor U4545 (N_4545,N_4311,N_4375);
or U4546 (N_4546,N_4418,N_4308);
nor U4547 (N_4547,N_4109,N_4285);
and U4548 (N_4548,N_4315,N_4379);
or U4549 (N_4549,N_4145,N_4125);
or U4550 (N_4550,N_4313,N_4390);
nand U4551 (N_4551,N_4281,N_4135);
nand U4552 (N_4552,N_4022,N_4347);
nor U4553 (N_4553,N_4448,N_4473);
and U4554 (N_4554,N_4049,N_4408);
or U4555 (N_4555,N_4402,N_4059);
or U4556 (N_4556,N_4400,N_4351);
nand U4557 (N_4557,N_4103,N_4381);
nor U4558 (N_4558,N_4158,N_4080);
or U4559 (N_4559,N_4406,N_4106);
xnor U4560 (N_4560,N_4221,N_4097);
xor U4561 (N_4561,N_4337,N_4238);
and U4562 (N_4562,N_4100,N_4195);
nor U4563 (N_4563,N_4139,N_4492);
and U4564 (N_4564,N_4434,N_4339);
or U4565 (N_4565,N_4470,N_4409);
xor U4566 (N_4566,N_4330,N_4460);
nor U4567 (N_4567,N_4424,N_4441);
nor U4568 (N_4568,N_4457,N_4362);
nor U4569 (N_4569,N_4250,N_4287);
or U4570 (N_4570,N_4454,N_4343);
and U4571 (N_4571,N_4140,N_4273);
and U4572 (N_4572,N_4223,N_4203);
or U4573 (N_4573,N_4404,N_4128);
and U4574 (N_4574,N_4363,N_4474);
or U4575 (N_4575,N_4070,N_4051);
or U4576 (N_4576,N_4456,N_4464);
xor U4577 (N_4577,N_4138,N_4096);
and U4578 (N_4578,N_4486,N_4246);
nand U4579 (N_4579,N_4023,N_4304);
or U4580 (N_4580,N_4160,N_4075);
nand U4581 (N_4581,N_4387,N_4032);
nand U4582 (N_4582,N_4413,N_4151);
nand U4583 (N_4583,N_4446,N_4367);
and U4584 (N_4584,N_4172,N_4497);
nand U4585 (N_4585,N_4263,N_4323);
and U4586 (N_4586,N_4231,N_4324);
xor U4587 (N_4587,N_4234,N_4412);
or U4588 (N_4588,N_4401,N_4344);
nor U4589 (N_4589,N_4469,N_4089);
nor U4590 (N_4590,N_4276,N_4320);
xnor U4591 (N_4591,N_4329,N_4177);
nand U4592 (N_4592,N_4377,N_4165);
or U4593 (N_4593,N_4268,N_4042);
nand U4594 (N_4594,N_4201,N_4200);
nand U4595 (N_4595,N_4170,N_4431);
and U4596 (N_4596,N_4197,N_4194);
nor U4597 (N_4597,N_4468,N_4199);
and U4598 (N_4598,N_4087,N_4230);
and U4599 (N_4599,N_4118,N_4432);
and U4600 (N_4600,N_4301,N_4282);
nor U4601 (N_4601,N_4066,N_4105);
xnor U4602 (N_4602,N_4317,N_4187);
xnor U4603 (N_4603,N_4267,N_4480);
and U4604 (N_4604,N_4114,N_4227);
or U4605 (N_4605,N_4182,N_4117);
or U4606 (N_4606,N_4260,N_4248);
xnor U4607 (N_4607,N_4407,N_4010);
or U4608 (N_4608,N_4425,N_4153);
and U4609 (N_4609,N_4015,N_4475);
and U4610 (N_4610,N_4040,N_4419);
nor U4611 (N_4611,N_4161,N_4083);
or U4612 (N_4612,N_4442,N_4451);
xnor U4613 (N_4613,N_4316,N_4062);
xnor U4614 (N_4614,N_4044,N_4270);
xor U4615 (N_4615,N_4167,N_4206);
and U4616 (N_4616,N_4335,N_4079);
nor U4617 (N_4617,N_4265,N_4372);
nor U4618 (N_4618,N_4000,N_4026);
nand U4619 (N_4619,N_4447,N_4077);
or U4620 (N_4620,N_4011,N_4148);
xnor U4621 (N_4621,N_4477,N_4052);
nor U4622 (N_4622,N_4466,N_4411);
and U4623 (N_4623,N_4055,N_4112);
nor U4624 (N_4624,N_4091,N_4310);
xor U4625 (N_4625,N_4039,N_4050);
nand U4626 (N_4626,N_4130,N_4101);
and U4627 (N_4627,N_4071,N_4332);
and U4628 (N_4628,N_4229,N_4355);
and U4629 (N_4629,N_4137,N_4133);
nand U4630 (N_4630,N_4490,N_4099);
or U4631 (N_4631,N_4255,N_4162);
or U4632 (N_4632,N_4174,N_4249);
nand U4633 (N_4633,N_4110,N_4462);
xor U4634 (N_4634,N_4383,N_4222);
and U4635 (N_4635,N_4331,N_4378);
and U4636 (N_4636,N_4371,N_4038);
nor U4637 (N_4637,N_4305,N_4325);
or U4638 (N_4638,N_4364,N_4478);
nor U4639 (N_4639,N_4235,N_4073);
or U4640 (N_4640,N_4175,N_4394);
or U4641 (N_4641,N_4254,N_4184);
nand U4642 (N_4642,N_4218,N_4213);
nor U4643 (N_4643,N_4366,N_4445);
and U4644 (N_4644,N_4479,N_4143);
xnor U4645 (N_4645,N_4403,N_4420);
or U4646 (N_4646,N_4017,N_4024);
nand U4647 (N_4647,N_4426,N_4300);
nand U4648 (N_4648,N_4421,N_4004);
or U4649 (N_4649,N_4482,N_4043);
and U4650 (N_4650,N_4336,N_4020);
and U4651 (N_4651,N_4279,N_4159);
nor U4652 (N_4652,N_4345,N_4166);
or U4653 (N_4653,N_4190,N_4207);
and U4654 (N_4654,N_4208,N_4211);
and U4655 (N_4655,N_4417,N_4428);
nor U4656 (N_4656,N_4003,N_4481);
nand U4657 (N_4657,N_4094,N_4082);
or U4658 (N_4658,N_4107,N_4416);
nor U4659 (N_4659,N_4048,N_4435);
or U4660 (N_4660,N_4061,N_4350);
nand U4661 (N_4661,N_4065,N_4389);
or U4662 (N_4662,N_4369,N_4214);
xor U4663 (N_4663,N_4009,N_4126);
xnor U4664 (N_4664,N_4005,N_4034);
and U4665 (N_4665,N_4168,N_4439);
nor U4666 (N_4666,N_4318,N_4399);
nor U4667 (N_4667,N_4120,N_4458);
nor U4668 (N_4668,N_4092,N_4463);
nor U4669 (N_4669,N_4302,N_4253);
and U4670 (N_4670,N_4090,N_4271);
xnor U4671 (N_4671,N_4291,N_4129);
xor U4672 (N_4672,N_4236,N_4113);
nand U4673 (N_4673,N_4186,N_4307);
or U4674 (N_4674,N_4269,N_4465);
nand U4675 (N_4675,N_4021,N_4239);
nor U4676 (N_4676,N_4150,N_4115);
xor U4677 (N_4677,N_4121,N_4102);
and U4678 (N_4678,N_4322,N_4173);
or U4679 (N_4679,N_4422,N_4410);
nand U4680 (N_4680,N_4278,N_4405);
and U4681 (N_4681,N_4006,N_4224);
nand U4682 (N_4682,N_4303,N_4178);
and U4683 (N_4683,N_4074,N_4440);
nor U4684 (N_4684,N_4452,N_4035);
and U4685 (N_4685,N_4283,N_4001);
xor U4686 (N_4686,N_4376,N_4025);
xnor U4687 (N_4687,N_4056,N_4415);
nand U4688 (N_4688,N_4496,N_4423);
nor U4689 (N_4689,N_4237,N_4349);
xor U4690 (N_4690,N_4338,N_4334);
nor U4691 (N_4691,N_4204,N_4116);
and U4692 (N_4692,N_4196,N_4360);
and U4693 (N_4693,N_4134,N_4494);
nand U4694 (N_4694,N_4054,N_4210);
and U4695 (N_4695,N_4202,N_4176);
nand U4696 (N_4696,N_4264,N_4085);
or U4697 (N_4697,N_4306,N_4251);
nor U4698 (N_4698,N_4286,N_4493);
and U4699 (N_4699,N_4388,N_4436);
or U4700 (N_4700,N_4164,N_4027);
and U4701 (N_4701,N_4018,N_4241);
and U4702 (N_4702,N_4312,N_4205);
xor U4703 (N_4703,N_4012,N_4008);
nand U4704 (N_4704,N_4078,N_4354);
nor U4705 (N_4705,N_4245,N_4014);
nand U4706 (N_4706,N_4093,N_4398);
xnor U4707 (N_4707,N_4163,N_4141);
xnor U4708 (N_4708,N_4084,N_4136);
nand U4709 (N_4709,N_4443,N_4495);
xor U4710 (N_4710,N_4444,N_4327);
xor U4711 (N_4711,N_4368,N_4156);
nor U4712 (N_4712,N_4104,N_4225);
nor U4713 (N_4713,N_4028,N_4180);
nand U4714 (N_4714,N_4437,N_4491);
nor U4715 (N_4715,N_4149,N_4373);
or U4716 (N_4716,N_4122,N_4067);
and U4717 (N_4717,N_4188,N_4427);
nor U4718 (N_4718,N_4467,N_4359);
nor U4719 (N_4719,N_4392,N_4487);
nor U4720 (N_4720,N_4353,N_4290);
or U4721 (N_4721,N_4275,N_4433);
and U4722 (N_4722,N_4058,N_4098);
and U4723 (N_4723,N_4154,N_4019);
and U4724 (N_4724,N_4191,N_4459);
nand U4725 (N_4725,N_4060,N_4483);
and U4726 (N_4726,N_4280,N_4352);
xor U4727 (N_4727,N_4361,N_4189);
nand U4728 (N_4728,N_4142,N_4328);
and U4729 (N_4729,N_4219,N_4053);
nand U4730 (N_4730,N_4198,N_4192);
xnor U4731 (N_4731,N_4258,N_4295);
and U4732 (N_4732,N_4386,N_4183);
nor U4733 (N_4733,N_4063,N_4449);
or U4734 (N_4734,N_4484,N_4397);
nand U4735 (N_4735,N_4430,N_4485);
and U4736 (N_4736,N_4240,N_4396);
and U4737 (N_4737,N_4293,N_4132);
xnor U4738 (N_4738,N_4450,N_4076);
nor U4739 (N_4739,N_4119,N_4472);
and U4740 (N_4740,N_4292,N_4193);
nand U4741 (N_4741,N_4064,N_4393);
nand U4742 (N_4742,N_4259,N_4171);
or U4743 (N_4743,N_4321,N_4356);
and U4744 (N_4744,N_4155,N_4131);
nor U4745 (N_4745,N_4326,N_4216);
xor U4746 (N_4746,N_4124,N_4069);
and U4747 (N_4747,N_4391,N_4088);
and U4748 (N_4748,N_4340,N_4152);
or U4749 (N_4749,N_4296,N_4169);
nor U4750 (N_4750,N_4435,N_4238);
nand U4751 (N_4751,N_4062,N_4269);
or U4752 (N_4752,N_4148,N_4209);
and U4753 (N_4753,N_4253,N_4153);
and U4754 (N_4754,N_4194,N_4391);
or U4755 (N_4755,N_4493,N_4263);
nor U4756 (N_4756,N_4391,N_4364);
nor U4757 (N_4757,N_4322,N_4334);
or U4758 (N_4758,N_4485,N_4324);
or U4759 (N_4759,N_4272,N_4061);
and U4760 (N_4760,N_4109,N_4430);
nand U4761 (N_4761,N_4239,N_4296);
xnor U4762 (N_4762,N_4002,N_4399);
nor U4763 (N_4763,N_4096,N_4355);
nor U4764 (N_4764,N_4488,N_4045);
and U4765 (N_4765,N_4448,N_4016);
xnor U4766 (N_4766,N_4378,N_4285);
or U4767 (N_4767,N_4257,N_4210);
or U4768 (N_4768,N_4019,N_4486);
xnor U4769 (N_4769,N_4268,N_4287);
or U4770 (N_4770,N_4397,N_4372);
nand U4771 (N_4771,N_4356,N_4308);
nor U4772 (N_4772,N_4377,N_4403);
nor U4773 (N_4773,N_4490,N_4168);
nand U4774 (N_4774,N_4104,N_4074);
xor U4775 (N_4775,N_4371,N_4212);
or U4776 (N_4776,N_4089,N_4199);
nor U4777 (N_4777,N_4323,N_4013);
nand U4778 (N_4778,N_4132,N_4214);
and U4779 (N_4779,N_4446,N_4479);
and U4780 (N_4780,N_4233,N_4370);
or U4781 (N_4781,N_4154,N_4320);
nor U4782 (N_4782,N_4315,N_4257);
and U4783 (N_4783,N_4332,N_4230);
or U4784 (N_4784,N_4485,N_4377);
xnor U4785 (N_4785,N_4465,N_4187);
or U4786 (N_4786,N_4228,N_4048);
or U4787 (N_4787,N_4231,N_4439);
nor U4788 (N_4788,N_4282,N_4068);
nor U4789 (N_4789,N_4094,N_4175);
and U4790 (N_4790,N_4017,N_4000);
nor U4791 (N_4791,N_4427,N_4380);
and U4792 (N_4792,N_4215,N_4466);
xnor U4793 (N_4793,N_4190,N_4490);
nand U4794 (N_4794,N_4269,N_4170);
xnor U4795 (N_4795,N_4486,N_4237);
nor U4796 (N_4796,N_4295,N_4246);
nor U4797 (N_4797,N_4211,N_4429);
or U4798 (N_4798,N_4145,N_4187);
nand U4799 (N_4799,N_4498,N_4365);
xor U4800 (N_4800,N_4390,N_4198);
or U4801 (N_4801,N_4302,N_4027);
nor U4802 (N_4802,N_4063,N_4140);
and U4803 (N_4803,N_4341,N_4266);
nand U4804 (N_4804,N_4160,N_4065);
or U4805 (N_4805,N_4062,N_4356);
nor U4806 (N_4806,N_4168,N_4491);
and U4807 (N_4807,N_4142,N_4203);
xnor U4808 (N_4808,N_4434,N_4145);
or U4809 (N_4809,N_4113,N_4444);
or U4810 (N_4810,N_4141,N_4013);
or U4811 (N_4811,N_4409,N_4054);
or U4812 (N_4812,N_4167,N_4169);
xor U4813 (N_4813,N_4145,N_4103);
nor U4814 (N_4814,N_4044,N_4019);
nor U4815 (N_4815,N_4022,N_4255);
or U4816 (N_4816,N_4307,N_4092);
nor U4817 (N_4817,N_4013,N_4032);
nand U4818 (N_4818,N_4196,N_4320);
or U4819 (N_4819,N_4003,N_4170);
and U4820 (N_4820,N_4216,N_4378);
and U4821 (N_4821,N_4378,N_4199);
and U4822 (N_4822,N_4002,N_4073);
nand U4823 (N_4823,N_4461,N_4433);
and U4824 (N_4824,N_4064,N_4135);
and U4825 (N_4825,N_4285,N_4397);
and U4826 (N_4826,N_4435,N_4414);
xor U4827 (N_4827,N_4429,N_4037);
nand U4828 (N_4828,N_4382,N_4246);
xor U4829 (N_4829,N_4188,N_4049);
or U4830 (N_4830,N_4217,N_4399);
xnor U4831 (N_4831,N_4300,N_4327);
and U4832 (N_4832,N_4149,N_4471);
xor U4833 (N_4833,N_4486,N_4447);
nor U4834 (N_4834,N_4022,N_4476);
nand U4835 (N_4835,N_4323,N_4321);
nand U4836 (N_4836,N_4351,N_4379);
xor U4837 (N_4837,N_4344,N_4332);
nor U4838 (N_4838,N_4072,N_4230);
nand U4839 (N_4839,N_4129,N_4343);
nand U4840 (N_4840,N_4037,N_4166);
xnor U4841 (N_4841,N_4426,N_4247);
and U4842 (N_4842,N_4020,N_4169);
nor U4843 (N_4843,N_4125,N_4166);
xnor U4844 (N_4844,N_4434,N_4222);
nor U4845 (N_4845,N_4088,N_4095);
nand U4846 (N_4846,N_4166,N_4271);
nor U4847 (N_4847,N_4221,N_4413);
nor U4848 (N_4848,N_4493,N_4401);
nor U4849 (N_4849,N_4064,N_4224);
nor U4850 (N_4850,N_4344,N_4094);
nor U4851 (N_4851,N_4146,N_4330);
nor U4852 (N_4852,N_4311,N_4072);
or U4853 (N_4853,N_4405,N_4197);
nor U4854 (N_4854,N_4488,N_4067);
xnor U4855 (N_4855,N_4104,N_4233);
nor U4856 (N_4856,N_4279,N_4481);
nand U4857 (N_4857,N_4032,N_4404);
nor U4858 (N_4858,N_4309,N_4368);
or U4859 (N_4859,N_4002,N_4082);
and U4860 (N_4860,N_4433,N_4270);
xor U4861 (N_4861,N_4292,N_4006);
nor U4862 (N_4862,N_4229,N_4015);
nand U4863 (N_4863,N_4111,N_4348);
nor U4864 (N_4864,N_4322,N_4360);
or U4865 (N_4865,N_4145,N_4331);
nand U4866 (N_4866,N_4443,N_4245);
nand U4867 (N_4867,N_4084,N_4233);
xor U4868 (N_4868,N_4338,N_4331);
and U4869 (N_4869,N_4451,N_4268);
and U4870 (N_4870,N_4245,N_4090);
xnor U4871 (N_4871,N_4148,N_4455);
xor U4872 (N_4872,N_4488,N_4237);
xnor U4873 (N_4873,N_4037,N_4403);
or U4874 (N_4874,N_4161,N_4098);
nand U4875 (N_4875,N_4135,N_4422);
and U4876 (N_4876,N_4170,N_4439);
xnor U4877 (N_4877,N_4302,N_4301);
and U4878 (N_4878,N_4151,N_4133);
and U4879 (N_4879,N_4293,N_4256);
nor U4880 (N_4880,N_4426,N_4101);
xnor U4881 (N_4881,N_4100,N_4237);
nand U4882 (N_4882,N_4481,N_4455);
nand U4883 (N_4883,N_4137,N_4437);
xor U4884 (N_4884,N_4228,N_4398);
nor U4885 (N_4885,N_4470,N_4465);
and U4886 (N_4886,N_4088,N_4256);
nor U4887 (N_4887,N_4300,N_4200);
xor U4888 (N_4888,N_4398,N_4088);
or U4889 (N_4889,N_4362,N_4260);
and U4890 (N_4890,N_4004,N_4348);
nand U4891 (N_4891,N_4176,N_4053);
and U4892 (N_4892,N_4087,N_4459);
nand U4893 (N_4893,N_4319,N_4237);
nor U4894 (N_4894,N_4205,N_4234);
nor U4895 (N_4895,N_4201,N_4071);
xor U4896 (N_4896,N_4101,N_4475);
xor U4897 (N_4897,N_4179,N_4106);
xnor U4898 (N_4898,N_4244,N_4403);
nand U4899 (N_4899,N_4495,N_4105);
and U4900 (N_4900,N_4422,N_4079);
xnor U4901 (N_4901,N_4433,N_4398);
or U4902 (N_4902,N_4104,N_4332);
nand U4903 (N_4903,N_4280,N_4034);
and U4904 (N_4904,N_4249,N_4102);
or U4905 (N_4905,N_4183,N_4296);
and U4906 (N_4906,N_4445,N_4367);
or U4907 (N_4907,N_4205,N_4155);
and U4908 (N_4908,N_4319,N_4147);
or U4909 (N_4909,N_4424,N_4259);
xnor U4910 (N_4910,N_4361,N_4062);
and U4911 (N_4911,N_4472,N_4273);
xor U4912 (N_4912,N_4072,N_4080);
nor U4913 (N_4913,N_4078,N_4232);
nand U4914 (N_4914,N_4184,N_4027);
or U4915 (N_4915,N_4343,N_4256);
xnor U4916 (N_4916,N_4111,N_4488);
nand U4917 (N_4917,N_4420,N_4271);
nor U4918 (N_4918,N_4316,N_4109);
nand U4919 (N_4919,N_4305,N_4411);
or U4920 (N_4920,N_4341,N_4069);
nor U4921 (N_4921,N_4481,N_4461);
and U4922 (N_4922,N_4220,N_4290);
xnor U4923 (N_4923,N_4348,N_4449);
or U4924 (N_4924,N_4138,N_4459);
nand U4925 (N_4925,N_4165,N_4494);
or U4926 (N_4926,N_4381,N_4496);
xnor U4927 (N_4927,N_4357,N_4194);
nor U4928 (N_4928,N_4055,N_4143);
or U4929 (N_4929,N_4276,N_4180);
nor U4930 (N_4930,N_4323,N_4084);
nand U4931 (N_4931,N_4396,N_4203);
nand U4932 (N_4932,N_4226,N_4345);
or U4933 (N_4933,N_4452,N_4174);
xor U4934 (N_4934,N_4452,N_4047);
nand U4935 (N_4935,N_4305,N_4485);
or U4936 (N_4936,N_4427,N_4316);
nand U4937 (N_4937,N_4215,N_4382);
xnor U4938 (N_4938,N_4317,N_4017);
nor U4939 (N_4939,N_4403,N_4106);
and U4940 (N_4940,N_4288,N_4057);
or U4941 (N_4941,N_4162,N_4107);
and U4942 (N_4942,N_4088,N_4027);
or U4943 (N_4943,N_4112,N_4302);
xor U4944 (N_4944,N_4258,N_4004);
nand U4945 (N_4945,N_4203,N_4041);
or U4946 (N_4946,N_4068,N_4229);
or U4947 (N_4947,N_4215,N_4118);
nand U4948 (N_4948,N_4002,N_4437);
or U4949 (N_4949,N_4335,N_4330);
or U4950 (N_4950,N_4412,N_4027);
nor U4951 (N_4951,N_4258,N_4456);
and U4952 (N_4952,N_4366,N_4104);
xnor U4953 (N_4953,N_4396,N_4196);
nor U4954 (N_4954,N_4006,N_4167);
nand U4955 (N_4955,N_4096,N_4496);
or U4956 (N_4956,N_4207,N_4102);
nand U4957 (N_4957,N_4002,N_4225);
nand U4958 (N_4958,N_4179,N_4326);
and U4959 (N_4959,N_4225,N_4120);
nand U4960 (N_4960,N_4044,N_4131);
xnor U4961 (N_4961,N_4283,N_4341);
and U4962 (N_4962,N_4077,N_4400);
and U4963 (N_4963,N_4226,N_4492);
or U4964 (N_4964,N_4169,N_4048);
and U4965 (N_4965,N_4102,N_4399);
or U4966 (N_4966,N_4364,N_4351);
nor U4967 (N_4967,N_4252,N_4198);
or U4968 (N_4968,N_4050,N_4405);
nand U4969 (N_4969,N_4465,N_4102);
and U4970 (N_4970,N_4438,N_4351);
xor U4971 (N_4971,N_4029,N_4434);
nor U4972 (N_4972,N_4489,N_4211);
nand U4973 (N_4973,N_4415,N_4024);
nand U4974 (N_4974,N_4034,N_4168);
and U4975 (N_4975,N_4345,N_4106);
and U4976 (N_4976,N_4448,N_4009);
and U4977 (N_4977,N_4441,N_4061);
nor U4978 (N_4978,N_4096,N_4444);
and U4979 (N_4979,N_4281,N_4493);
and U4980 (N_4980,N_4473,N_4325);
and U4981 (N_4981,N_4199,N_4209);
nand U4982 (N_4982,N_4483,N_4124);
nor U4983 (N_4983,N_4087,N_4042);
and U4984 (N_4984,N_4489,N_4262);
nand U4985 (N_4985,N_4457,N_4451);
and U4986 (N_4986,N_4077,N_4027);
nand U4987 (N_4987,N_4210,N_4194);
xor U4988 (N_4988,N_4029,N_4291);
nand U4989 (N_4989,N_4484,N_4003);
nand U4990 (N_4990,N_4383,N_4057);
and U4991 (N_4991,N_4480,N_4045);
and U4992 (N_4992,N_4281,N_4238);
and U4993 (N_4993,N_4053,N_4091);
and U4994 (N_4994,N_4263,N_4476);
nor U4995 (N_4995,N_4404,N_4210);
and U4996 (N_4996,N_4279,N_4273);
and U4997 (N_4997,N_4264,N_4048);
and U4998 (N_4998,N_4110,N_4155);
and U4999 (N_4999,N_4269,N_4071);
xnor U5000 (N_5000,N_4908,N_4808);
and U5001 (N_5001,N_4733,N_4644);
nor U5002 (N_5002,N_4885,N_4829);
nor U5003 (N_5003,N_4870,N_4500);
and U5004 (N_5004,N_4887,N_4533);
nor U5005 (N_5005,N_4928,N_4797);
nor U5006 (N_5006,N_4941,N_4804);
or U5007 (N_5007,N_4691,N_4790);
nor U5008 (N_5008,N_4626,N_4554);
or U5009 (N_5009,N_4844,N_4562);
nand U5010 (N_5010,N_4613,N_4745);
nand U5011 (N_5011,N_4837,N_4523);
nor U5012 (N_5012,N_4712,N_4749);
xor U5013 (N_5013,N_4976,N_4738);
or U5014 (N_5014,N_4871,N_4549);
and U5015 (N_5015,N_4772,N_4728);
or U5016 (N_5016,N_4815,N_4710);
and U5017 (N_5017,N_4588,N_4722);
xor U5018 (N_5018,N_4996,N_4664);
xnor U5019 (N_5019,N_4542,N_4576);
nor U5020 (N_5020,N_4584,N_4913);
and U5021 (N_5021,N_4751,N_4930);
xor U5022 (N_5022,N_4938,N_4730);
nor U5023 (N_5023,N_4583,N_4592);
or U5024 (N_5024,N_4907,N_4971);
xnor U5025 (N_5025,N_4657,N_4964);
nor U5026 (N_5026,N_4902,N_4715);
or U5027 (N_5027,N_4690,N_4799);
or U5028 (N_5028,N_4606,N_4636);
or U5029 (N_5029,N_4561,N_4742);
nand U5030 (N_5030,N_4543,N_4527);
nand U5031 (N_5031,N_4944,N_4535);
xor U5032 (N_5032,N_4998,N_4640);
nand U5033 (N_5033,N_4882,N_4507);
xor U5034 (N_5034,N_4771,N_4858);
and U5035 (N_5035,N_4857,N_4571);
and U5036 (N_5036,N_4853,N_4696);
nand U5037 (N_5037,N_4748,N_4619);
xor U5038 (N_5038,N_4994,N_4973);
and U5039 (N_5039,N_4741,N_4635);
nand U5040 (N_5040,N_4925,N_4717);
or U5041 (N_5041,N_4982,N_4586);
or U5042 (N_5042,N_4631,N_4521);
or U5043 (N_5043,N_4823,N_4508);
and U5044 (N_5044,N_4598,N_4827);
and U5045 (N_5045,N_4660,N_4989);
nand U5046 (N_5046,N_4943,N_4750);
or U5047 (N_5047,N_4689,N_4628);
and U5048 (N_5048,N_4632,N_4517);
xnor U5049 (N_5049,N_4579,N_4642);
nand U5050 (N_5050,N_4623,N_4822);
or U5051 (N_5051,N_4604,N_4869);
nor U5052 (N_5052,N_4936,N_4630);
or U5053 (N_5053,N_4846,N_4716);
and U5054 (N_5054,N_4794,N_4565);
or U5055 (N_5055,N_4945,N_4686);
nand U5056 (N_5056,N_4924,N_4904);
and U5057 (N_5057,N_4911,N_4877);
nand U5058 (N_5058,N_4849,N_4843);
nor U5059 (N_5059,N_4610,N_4611);
or U5060 (N_5060,N_4891,N_4914);
and U5061 (N_5061,N_4793,N_4676);
nand U5062 (N_5062,N_4950,N_4530);
and U5063 (N_5063,N_4739,N_4693);
or U5064 (N_5064,N_4638,N_4939);
and U5065 (N_5065,N_4706,N_4672);
nand U5066 (N_5066,N_4569,N_4865);
nor U5067 (N_5067,N_4560,N_4556);
nand U5068 (N_5068,N_4627,N_4680);
nor U5069 (N_5069,N_4662,N_4677);
nor U5070 (N_5070,N_4667,N_4502);
or U5071 (N_5071,N_4724,N_4841);
xor U5072 (N_5072,N_4572,N_4697);
xnor U5073 (N_5073,N_4912,N_4951);
and U5074 (N_5074,N_4587,N_4983);
nand U5075 (N_5075,N_4819,N_4743);
nand U5076 (N_5076,N_4863,N_4949);
and U5077 (N_5077,N_4740,N_4605);
xnor U5078 (N_5078,N_4753,N_4889);
or U5079 (N_5079,N_4665,N_4763);
xnor U5080 (N_5080,N_4736,N_4504);
or U5081 (N_5081,N_4821,N_4634);
nand U5082 (N_5082,N_4616,N_4528);
and U5083 (N_5083,N_4931,N_4957);
and U5084 (N_5084,N_4558,N_4550);
nand U5085 (N_5085,N_4969,N_4537);
nand U5086 (N_5086,N_4608,N_4655);
or U5087 (N_5087,N_4895,N_4614);
nand U5088 (N_5088,N_4699,N_4834);
xor U5089 (N_5089,N_4862,N_4761);
or U5090 (N_5090,N_4591,N_4547);
nor U5091 (N_5091,N_4773,N_4835);
xnor U5092 (N_5092,N_4757,N_4780);
nor U5093 (N_5093,N_4568,N_4539);
or U5094 (N_5094,N_4702,N_4812);
xor U5095 (N_5095,N_4966,N_4932);
or U5096 (N_5096,N_4595,N_4621);
xnor U5097 (N_5097,N_4708,N_4714);
or U5098 (N_5098,N_4811,N_4776);
xnor U5099 (N_5099,N_4937,N_4501);
or U5100 (N_5100,N_4510,N_4816);
nor U5101 (N_5101,N_4511,N_4872);
and U5102 (N_5102,N_4593,N_4573);
or U5103 (N_5103,N_4555,N_4833);
and U5104 (N_5104,N_4884,N_4756);
nand U5105 (N_5105,N_4781,N_4639);
nand U5106 (N_5106,N_4775,N_4620);
and U5107 (N_5107,N_4876,N_4618);
xnor U5108 (N_5108,N_4786,N_4522);
nor U5109 (N_5109,N_4553,N_4727);
or U5110 (N_5110,N_4546,N_4955);
or U5111 (N_5111,N_4578,N_4997);
or U5112 (N_5112,N_4651,N_4836);
and U5113 (N_5113,N_4968,N_4653);
xnor U5114 (N_5114,N_4769,N_4585);
and U5115 (N_5115,N_4954,N_4903);
nand U5116 (N_5116,N_4525,N_4864);
xor U5117 (N_5117,N_4559,N_4852);
xnor U5118 (N_5118,N_4538,N_4762);
nand U5119 (N_5119,N_4881,N_4566);
xnor U5120 (N_5120,N_4652,N_4920);
nand U5121 (N_5121,N_4601,N_4946);
xnor U5122 (N_5122,N_4602,N_4734);
nor U5123 (N_5123,N_4529,N_4654);
or U5124 (N_5124,N_4892,N_4979);
xnor U5125 (N_5125,N_4807,N_4860);
xnor U5126 (N_5126,N_4959,N_4961);
xnor U5127 (N_5127,N_4866,N_4671);
or U5128 (N_5128,N_4596,N_4791);
nor U5129 (N_5129,N_4999,N_4802);
xor U5130 (N_5130,N_4935,N_4625);
or U5131 (N_5131,N_4970,N_4612);
or U5132 (N_5132,N_4540,N_4649);
and U5133 (N_5133,N_4993,N_4867);
xor U5134 (N_5134,N_4622,N_4894);
nor U5135 (N_5135,N_4806,N_4668);
and U5136 (N_5136,N_4766,N_4704);
and U5137 (N_5137,N_4544,N_4875);
nand U5138 (N_5138,N_4552,N_4800);
nor U5139 (N_5139,N_4603,N_4721);
or U5140 (N_5140,N_4956,N_4787);
xor U5141 (N_5141,N_4856,N_4792);
nor U5142 (N_5142,N_4770,N_4520);
or U5143 (N_5143,N_4942,N_4817);
and U5144 (N_5144,N_4624,N_4725);
xor U5145 (N_5145,N_4899,N_4893);
xor U5146 (N_5146,N_4980,N_4582);
and U5147 (N_5147,N_4851,N_4663);
nor U5148 (N_5148,N_4695,N_4838);
nor U5149 (N_5149,N_4915,N_4659);
and U5150 (N_5150,N_4709,N_4992);
or U5151 (N_5151,N_4617,N_4647);
nand U5152 (N_5152,N_4842,N_4607);
nor U5153 (N_5153,N_4990,N_4921);
and U5154 (N_5154,N_4754,N_4948);
nand U5155 (N_5155,N_4906,N_4813);
or U5156 (N_5156,N_4518,N_4633);
nor U5157 (N_5157,N_4952,N_4960);
nor U5158 (N_5158,N_4681,N_4703);
xor U5159 (N_5159,N_4995,N_4590);
xnor U5160 (N_5160,N_4683,N_4981);
or U5161 (N_5161,N_4927,N_4726);
nand U5162 (N_5162,N_4963,N_4958);
xor U5163 (N_5163,N_4803,N_4516);
xor U5164 (N_5164,N_4563,N_4880);
or U5165 (N_5165,N_4698,N_4720);
or U5166 (N_5166,N_4747,N_4735);
xnor U5167 (N_5167,N_4814,N_4809);
or U5168 (N_5168,N_4541,N_4929);
nor U5169 (N_5169,N_4861,N_4905);
or U5170 (N_5170,N_4953,N_4512);
nor U5171 (N_5171,N_4828,N_4599);
nor U5172 (N_5172,N_4637,N_4825);
or U5173 (N_5173,N_4922,N_4965);
and U5174 (N_5174,N_4755,N_4679);
nand U5175 (N_5175,N_4581,N_4645);
or U5176 (N_5176,N_4514,N_4707);
and U5177 (N_5177,N_4918,N_4675);
xor U5178 (N_5178,N_4847,N_4575);
and U5179 (N_5179,N_4705,N_4744);
nor U5180 (N_5180,N_4839,N_4685);
or U5181 (N_5181,N_4910,N_4687);
nand U5182 (N_5182,N_4701,N_4795);
nor U5183 (N_5183,N_4923,N_4629);
or U5184 (N_5184,N_4991,N_4919);
nand U5185 (N_5185,N_4656,N_4531);
xor U5186 (N_5186,N_4934,N_4641);
nor U5187 (N_5187,N_4767,N_4886);
nor U5188 (N_5188,N_4796,N_4896);
xor U5189 (N_5189,N_4580,N_4788);
nand U5190 (N_5190,N_4798,N_4758);
and U5191 (N_5191,N_4694,N_4732);
or U5192 (N_5192,N_4826,N_4848);
and U5193 (N_5193,N_4567,N_4783);
nand U5194 (N_5194,N_4832,N_4940);
nand U5195 (N_5195,N_4729,N_4840);
nor U5196 (N_5196,N_4805,N_4974);
nor U5197 (N_5197,N_4985,N_4972);
nor U5198 (N_5198,N_4897,N_4820);
and U5199 (N_5199,N_4678,N_4524);
and U5200 (N_5200,N_4977,N_4768);
nor U5201 (N_5201,N_4850,N_4615);
xor U5202 (N_5202,N_4987,N_4782);
and U5203 (N_5203,N_4682,N_4777);
and U5204 (N_5204,N_4845,N_4765);
or U5205 (N_5205,N_4532,N_4933);
nor U5206 (N_5206,N_4785,N_4648);
nor U5207 (N_5207,N_4711,N_4564);
or U5208 (N_5208,N_4661,N_4513);
and U5209 (N_5209,N_4673,N_4646);
and U5210 (N_5210,N_4688,N_4670);
or U5211 (N_5211,N_4574,N_4898);
xnor U5212 (N_5212,N_4926,N_4779);
xor U5213 (N_5213,N_4978,N_4669);
and U5214 (N_5214,N_4810,N_4774);
xnor U5215 (N_5215,N_4988,N_4570);
xnor U5216 (N_5216,N_4916,N_4986);
nand U5217 (N_5217,N_4890,N_4759);
or U5218 (N_5218,N_4909,N_4818);
xor U5219 (N_5219,N_4536,N_4883);
and U5220 (N_5220,N_4674,N_4548);
xor U5221 (N_5221,N_4878,N_4868);
nand U5222 (N_5222,N_4643,N_4594);
nor U5223 (N_5223,N_4984,N_4967);
nand U5224 (N_5224,N_4879,N_4515);
xor U5225 (N_5225,N_4719,N_4658);
nand U5226 (N_5226,N_4723,N_4874);
nand U5227 (N_5227,N_4713,N_4855);
nor U5228 (N_5228,N_4888,N_4503);
and U5229 (N_5229,N_4859,N_4505);
and U5230 (N_5230,N_4824,N_4551);
nor U5231 (N_5231,N_4917,N_4519);
nor U5232 (N_5232,N_4760,N_4597);
xor U5233 (N_5233,N_4650,N_4731);
nor U5234 (N_5234,N_4589,N_4526);
and U5235 (N_5235,N_4577,N_4778);
nand U5236 (N_5236,N_4509,N_4784);
or U5237 (N_5237,N_4600,N_4764);
nand U5238 (N_5238,N_4962,N_4801);
or U5239 (N_5239,N_4901,N_4789);
nor U5240 (N_5240,N_4700,N_4506);
and U5241 (N_5241,N_4752,N_4609);
and U5242 (N_5242,N_4684,N_4947);
nor U5243 (N_5243,N_4975,N_4666);
nand U5244 (N_5244,N_4746,N_4873);
xor U5245 (N_5245,N_4534,N_4718);
xor U5246 (N_5246,N_4545,N_4831);
nor U5247 (N_5247,N_4854,N_4900);
xnor U5248 (N_5248,N_4692,N_4557);
or U5249 (N_5249,N_4830,N_4737);
xnor U5250 (N_5250,N_4560,N_4678);
xor U5251 (N_5251,N_4760,N_4687);
nand U5252 (N_5252,N_4960,N_4890);
and U5253 (N_5253,N_4759,N_4825);
nor U5254 (N_5254,N_4588,N_4917);
xnor U5255 (N_5255,N_4938,N_4909);
nor U5256 (N_5256,N_4810,N_4750);
nor U5257 (N_5257,N_4929,N_4994);
xnor U5258 (N_5258,N_4870,N_4917);
xor U5259 (N_5259,N_4610,N_4952);
or U5260 (N_5260,N_4706,N_4943);
nand U5261 (N_5261,N_4834,N_4742);
nor U5262 (N_5262,N_4593,N_4899);
nor U5263 (N_5263,N_4820,N_4594);
and U5264 (N_5264,N_4702,N_4507);
and U5265 (N_5265,N_4661,N_4761);
nand U5266 (N_5266,N_4795,N_4676);
nor U5267 (N_5267,N_4597,N_4944);
nor U5268 (N_5268,N_4532,N_4797);
or U5269 (N_5269,N_4657,N_4703);
xor U5270 (N_5270,N_4989,N_4716);
or U5271 (N_5271,N_4965,N_4820);
or U5272 (N_5272,N_4770,N_4963);
nor U5273 (N_5273,N_4723,N_4938);
xnor U5274 (N_5274,N_4572,N_4617);
xor U5275 (N_5275,N_4649,N_4595);
or U5276 (N_5276,N_4909,N_4568);
nor U5277 (N_5277,N_4538,N_4500);
nand U5278 (N_5278,N_4633,N_4991);
or U5279 (N_5279,N_4676,N_4800);
nor U5280 (N_5280,N_4629,N_4958);
nand U5281 (N_5281,N_4560,N_4505);
and U5282 (N_5282,N_4697,N_4633);
nor U5283 (N_5283,N_4573,N_4621);
and U5284 (N_5284,N_4533,N_4995);
nor U5285 (N_5285,N_4850,N_4806);
nor U5286 (N_5286,N_4786,N_4933);
or U5287 (N_5287,N_4704,N_4750);
nand U5288 (N_5288,N_4953,N_4944);
and U5289 (N_5289,N_4618,N_4685);
xnor U5290 (N_5290,N_4862,N_4524);
xor U5291 (N_5291,N_4505,N_4835);
xnor U5292 (N_5292,N_4780,N_4546);
nor U5293 (N_5293,N_4717,N_4581);
xor U5294 (N_5294,N_4865,N_4898);
or U5295 (N_5295,N_4639,N_4769);
and U5296 (N_5296,N_4824,N_4523);
xor U5297 (N_5297,N_4944,N_4554);
nand U5298 (N_5298,N_4578,N_4823);
and U5299 (N_5299,N_4954,N_4906);
xor U5300 (N_5300,N_4965,N_4593);
nor U5301 (N_5301,N_4970,N_4501);
nor U5302 (N_5302,N_4571,N_4876);
and U5303 (N_5303,N_4686,N_4615);
nand U5304 (N_5304,N_4933,N_4684);
nand U5305 (N_5305,N_4893,N_4832);
nor U5306 (N_5306,N_4990,N_4854);
xor U5307 (N_5307,N_4751,N_4518);
xnor U5308 (N_5308,N_4680,N_4809);
and U5309 (N_5309,N_4975,N_4569);
or U5310 (N_5310,N_4561,N_4566);
or U5311 (N_5311,N_4557,N_4689);
nand U5312 (N_5312,N_4603,N_4860);
nor U5313 (N_5313,N_4995,N_4742);
nor U5314 (N_5314,N_4854,N_4650);
or U5315 (N_5315,N_4641,N_4667);
and U5316 (N_5316,N_4682,N_4616);
nand U5317 (N_5317,N_4783,N_4990);
nand U5318 (N_5318,N_4885,N_4680);
or U5319 (N_5319,N_4555,N_4574);
nor U5320 (N_5320,N_4567,N_4811);
nand U5321 (N_5321,N_4897,N_4642);
nor U5322 (N_5322,N_4980,N_4593);
and U5323 (N_5323,N_4688,N_4777);
or U5324 (N_5324,N_4992,N_4659);
xor U5325 (N_5325,N_4840,N_4969);
nand U5326 (N_5326,N_4567,N_4696);
xor U5327 (N_5327,N_4889,N_4974);
nor U5328 (N_5328,N_4603,N_4654);
nor U5329 (N_5329,N_4737,N_4695);
and U5330 (N_5330,N_4930,N_4771);
and U5331 (N_5331,N_4972,N_4663);
nor U5332 (N_5332,N_4749,N_4921);
xor U5333 (N_5333,N_4670,N_4723);
or U5334 (N_5334,N_4560,N_4703);
nor U5335 (N_5335,N_4792,N_4945);
nand U5336 (N_5336,N_4766,N_4599);
nand U5337 (N_5337,N_4595,N_4909);
or U5338 (N_5338,N_4542,N_4688);
xor U5339 (N_5339,N_4993,N_4909);
nand U5340 (N_5340,N_4759,N_4747);
nor U5341 (N_5341,N_4858,N_4548);
nand U5342 (N_5342,N_4589,N_4793);
nor U5343 (N_5343,N_4526,N_4613);
xor U5344 (N_5344,N_4695,N_4841);
nor U5345 (N_5345,N_4903,N_4811);
or U5346 (N_5346,N_4516,N_4645);
or U5347 (N_5347,N_4836,N_4753);
xor U5348 (N_5348,N_4904,N_4864);
nor U5349 (N_5349,N_4573,N_4550);
nor U5350 (N_5350,N_4834,N_4595);
and U5351 (N_5351,N_4745,N_4808);
or U5352 (N_5352,N_4835,N_4632);
and U5353 (N_5353,N_4533,N_4812);
nand U5354 (N_5354,N_4985,N_4644);
or U5355 (N_5355,N_4630,N_4538);
or U5356 (N_5356,N_4849,N_4713);
nand U5357 (N_5357,N_4851,N_4609);
nand U5358 (N_5358,N_4767,N_4782);
nand U5359 (N_5359,N_4987,N_4842);
and U5360 (N_5360,N_4730,N_4609);
and U5361 (N_5361,N_4818,N_4749);
or U5362 (N_5362,N_4687,N_4998);
nor U5363 (N_5363,N_4623,N_4675);
nor U5364 (N_5364,N_4751,N_4746);
or U5365 (N_5365,N_4634,N_4617);
nand U5366 (N_5366,N_4999,N_4703);
or U5367 (N_5367,N_4758,N_4677);
and U5368 (N_5368,N_4888,N_4762);
xnor U5369 (N_5369,N_4720,N_4546);
nor U5370 (N_5370,N_4565,N_4677);
xnor U5371 (N_5371,N_4972,N_4869);
and U5372 (N_5372,N_4980,N_4734);
nor U5373 (N_5373,N_4832,N_4629);
nand U5374 (N_5374,N_4662,N_4670);
and U5375 (N_5375,N_4700,N_4913);
nor U5376 (N_5376,N_4577,N_4608);
xnor U5377 (N_5377,N_4998,N_4671);
and U5378 (N_5378,N_4831,N_4724);
nor U5379 (N_5379,N_4739,N_4867);
nand U5380 (N_5380,N_4902,N_4937);
nand U5381 (N_5381,N_4861,N_4691);
and U5382 (N_5382,N_4902,N_4553);
nor U5383 (N_5383,N_4803,N_4993);
nor U5384 (N_5384,N_4819,N_4624);
or U5385 (N_5385,N_4658,N_4634);
xnor U5386 (N_5386,N_4904,N_4758);
xnor U5387 (N_5387,N_4763,N_4530);
xor U5388 (N_5388,N_4688,N_4775);
nor U5389 (N_5389,N_4617,N_4520);
or U5390 (N_5390,N_4928,N_4633);
nand U5391 (N_5391,N_4642,N_4777);
nor U5392 (N_5392,N_4509,N_4907);
nand U5393 (N_5393,N_4650,N_4746);
xor U5394 (N_5394,N_4620,N_4894);
nand U5395 (N_5395,N_4945,N_4952);
xor U5396 (N_5396,N_4613,N_4978);
or U5397 (N_5397,N_4999,N_4544);
or U5398 (N_5398,N_4895,N_4568);
and U5399 (N_5399,N_4649,N_4790);
nor U5400 (N_5400,N_4513,N_4599);
and U5401 (N_5401,N_4602,N_4797);
nor U5402 (N_5402,N_4807,N_4659);
nand U5403 (N_5403,N_4531,N_4744);
xor U5404 (N_5404,N_4708,N_4951);
xor U5405 (N_5405,N_4600,N_4919);
nand U5406 (N_5406,N_4903,N_4919);
and U5407 (N_5407,N_4998,N_4585);
nor U5408 (N_5408,N_4921,N_4852);
or U5409 (N_5409,N_4737,N_4523);
and U5410 (N_5410,N_4742,N_4784);
nor U5411 (N_5411,N_4861,N_4753);
xor U5412 (N_5412,N_4520,N_4598);
xor U5413 (N_5413,N_4944,N_4752);
and U5414 (N_5414,N_4967,N_4960);
nor U5415 (N_5415,N_4565,N_4843);
nand U5416 (N_5416,N_4532,N_4896);
and U5417 (N_5417,N_4561,N_4952);
or U5418 (N_5418,N_4790,N_4907);
xnor U5419 (N_5419,N_4943,N_4919);
and U5420 (N_5420,N_4768,N_4750);
nand U5421 (N_5421,N_4787,N_4978);
xor U5422 (N_5422,N_4836,N_4658);
nor U5423 (N_5423,N_4706,N_4975);
nand U5424 (N_5424,N_4872,N_4520);
xnor U5425 (N_5425,N_4537,N_4743);
xor U5426 (N_5426,N_4816,N_4953);
or U5427 (N_5427,N_4849,N_4897);
or U5428 (N_5428,N_4778,N_4726);
or U5429 (N_5429,N_4866,N_4931);
nand U5430 (N_5430,N_4808,N_4630);
or U5431 (N_5431,N_4506,N_4618);
nand U5432 (N_5432,N_4919,N_4956);
or U5433 (N_5433,N_4826,N_4542);
nor U5434 (N_5434,N_4742,N_4798);
nor U5435 (N_5435,N_4964,N_4982);
nand U5436 (N_5436,N_4714,N_4921);
and U5437 (N_5437,N_4603,N_4855);
nor U5438 (N_5438,N_4902,N_4836);
or U5439 (N_5439,N_4849,N_4814);
xnor U5440 (N_5440,N_4652,N_4604);
nand U5441 (N_5441,N_4883,N_4808);
nand U5442 (N_5442,N_4616,N_4605);
nor U5443 (N_5443,N_4655,N_4905);
or U5444 (N_5444,N_4795,N_4886);
xor U5445 (N_5445,N_4829,N_4614);
nand U5446 (N_5446,N_4804,N_4752);
nand U5447 (N_5447,N_4607,N_4569);
and U5448 (N_5448,N_4617,N_4809);
xnor U5449 (N_5449,N_4678,N_4906);
xnor U5450 (N_5450,N_4969,N_4612);
xor U5451 (N_5451,N_4640,N_4778);
nand U5452 (N_5452,N_4554,N_4931);
xor U5453 (N_5453,N_4689,N_4723);
xnor U5454 (N_5454,N_4601,N_4995);
and U5455 (N_5455,N_4838,N_4674);
and U5456 (N_5456,N_4874,N_4851);
nand U5457 (N_5457,N_4636,N_4857);
or U5458 (N_5458,N_4691,N_4932);
xnor U5459 (N_5459,N_4519,N_4689);
nor U5460 (N_5460,N_4811,N_4860);
or U5461 (N_5461,N_4968,N_4669);
nor U5462 (N_5462,N_4808,N_4814);
xnor U5463 (N_5463,N_4538,N_4809);
or U5464 (N_5464,N_4765,N_4953);
or U5465 (N_5465,N_4734,N_4505);
xnor U5466 (N_5466,N_4844,N_4717);
nor U5467 (N_5467,N_4727,N_4631);
or U5468 (N_5468,N_4969,N_4766);
nand U5469 (N_5469,N_4877,N_4765);
or U5470 (N_5470,N_4628,N_4729);
or U5471 (N_5471,N_4901,N_4527);
and U5472 (N_5472,N_4839,N_4951);
nor U5473 (N_5473,N_4517,N_4941);
xnor U5474 (N_5474,N_4858,N_4970);
and U5475 (N_5475,N_4660,N_4752);
and U5476 (N_5476,N_4931,N_4755);
nand U5477 (N_5477,N_4982,N_4617);
or U5478 (N_5478,N_4874,N_4508);
nand U5479 (N_5479,N_4640,N_4524);
and U5480 (N_5480,N_4949,N_4912);
xor U5481 (N_5481,N_4920,N_4783);
nor U5482 (N_5482,N_4595,N_4801);
and U5483 (N_5483,N_4769,N_4535);
nand U5484 (N_5484,N_4668,N_4666);
xor U5485 (N_5485,N_4718,N_4595);
or U5486 (N_5486,N_4757,N_4588);
nand U5487 (N_5487,N_4783,N_4848);
and U5488 (N_5488,N_4826,N_4675);
nand U5489 (N_5489,N_4857,N_4677);
nor U5490 (N_5490,N_4751,N_4679);
xor U5491 (N_5491,N_4987,N_4813);
nor U5492 (N_5492,N_4881,N_4645);
nor U5493 (N_5493,N_4527,N_4524);
and U5494 (N_5494,N_4951,N_4731);
xor U5495 (N_5495,N_4818,N_4893);
nor U5496 (N_5496,N_4812,N_4801);
or U5497 (N_5497,N_4838,N_4503);
nand U5498 (N_5498,N_4664,N_4896);
or U5499 (N_5499,N_4965,N_4843);
or U5500 (N_5500,N_5401,N_5479);
or U5501 (N_5501,N_5386,N_5013);
nor U5502 (N_5502,N_5200,N_5436);
nand U5503 (N_5503,N_5288,N_5142);
nand U5504 (N_5504,N_5480,N_5374);
or U5505 (N_5505,N_5080,N_5253);
xnor U5506 (N_5506,N_5129,N_5377);
and U5507 (N_5507,N_5381,N_5031);
or U5508 (N_5508,N_5462,N_5357);
nand U5509 (N_5509,N_5388,N_5495);
xnor U5510 (N_5510,N_5322,N_5182);
nand U5511 (N_5511,N_5092,N_5130);
and U5512 (N_5512,N_5299,N_5094);
xor U5513 (N_5513,N_5372,N_5148);
or U5514 (N_5514,N_5290,N_5348);
and U5515 (N_5515,N_5282,N_5280);
and U5516 (N_5516,N_5215,N_5447);
nor U5517 (N_5517,N_5435,N_5395);
nor U5518 (N_5518,N_5229,N_5276);
nand U5519 (N_5519,N_5360,N_5459);
or U5520 (N_5520,N_5050,N_5361);
xnor U5521 (N_5521,N_5057,N_5499);
or U5522 (N_5522,N_5373,N_5019);
nand U5523 (N_5523,N_5203,N_5431);
nand U5524 (N_5524,N_5305,N_5230);
and U5525 (N_5525,N_5392,N_5258);
or U5526 (N_5526,N_5359,N_5201);
xnor U5527 (N_5527,N_5303,N_5478);
nand U5528 (N_5528,N_5312,N_5400);
or U5529 (N_5529,N_5437,N_5457);
or U5530 (N_5530,N_5206,N_5167);
xor U5531 (N_5531,N_5012,N_5430);
or U5532 (N_5532,N_5150,N_5445);
nor U5533 (N_5533,N_5032,N_5036);
xor U5534 (N_5534,N_5110,N_5375);
nor U5535 (N_5535,N_5433,N_5325);
and U5536 (N_5536,N_5496,N_5185);
xor U5537 (N_5537,N_5407,N_5155);
and U5538 (N_5538,N_5293,N_5277);
nand U5539 (N_5539,N_5441,N_5053);
nand U5540 (N_5540,N_5465,N_5202);
nand U5541 (N_5541,N_5417,N_5298);
xor U5542 (N_5542,N_5389,N_5485);
or U5543 (N_5543,N_5027,N_5264);
nand U5544 (N_5544,N_5035,N_5390);
nand U5545 (N_5545,N_5368,N_5211);
nand U5546 (N_5546,N_5175,N_5404);
xnor U5547 (N_5547,N_5346,N_5428);
xnor U5548 (N_5548,N_5358,N_5052);
or U5549 (N_5549,N_5330,N_5331);
nand U5550 (N_5550,N_5335,N_5458);
or U5551 (N_5551,N_5158,N_5051);
nand U5552 (N_5552,N_5188,N_5168);
xnor U5553 (N_5553,N_5432,N_5444);
nor U5554 (N_5554,N_5213,N_5207);
nand U5555 (N_5555,N_5045,N_5272);
and U5556 (N_5556,N_5235,N_5310);
nand U5557 (N_5557,N_5145,N_5107);
nand U5558 (N_5558,N_5119,N_5010);
nand U5559 (N_5559,N_5149,N_5289);
nand U5560 (N_5560,N_5398,N_5038);
xnor U5561 (N_5561,N_5278,N_5486);
xnor U5562 (N_5562,N_5260,N_5197);
and U5563 (N_5563,N_5047,N_5232);
and U5564 (N_5564,N_5385,N_5065);
xnor U5565 (N_5565,N_5350,N_5328);
nor U5566 (N_5566,N_5384,N_5429);
nor U5567 (N_5567,N_5420,N_5251);
or U5568 (N_5568,N_5442,N_5214);
nand U5569 (N_5569,N_5466,N_5410);
or U5570 (N_5570,N_5091,N_5041);
and U5571 (N_5571,N_5326,N_5231);
and U5572 (N_5572,N_5128,N_5409);
and U5573 (N_5573,N_5406,N_5402);
or U5574 (N_5574,N_5237,N_5244);
xnor U5575 (N_5575,N_5489,N_5176);
xnor U5576 (N_5576,N_5339,N_5482);
and U5577 (N_5577,N_5367,N_5153);
and U5578 (N_5578,N_5008,N_5227);
or U5579 (N_5579,N_5252,N_5191);
nor U5580 (N_5580,N_5492,N_5306);
nand U5581 (N_5581,N_5140,N_5484);
xnor U5582 (N_5582,N_5240,N_5454);
nand U5583 (N_5583,N_5332,N_5068);
xnor U5584 (N_5584,N_5024,N_5297);
nor U5585 (N_5585,N_5069,N_5286);
and U5586 (N_5586,N_5029,N_5343);
or U5587 (N_5587,N_5085,N_5030);
nand U5588 (N_5588,N_5329,N_5313);
nand U5589 (N_5589,N_5151,N_5194);
xor U5590 (N_5590,N_5370,N_5104);
or U5591 (N_5591,N_5112,N_5355);
nor U5592 (N_5592,N_5247,N_5396);
nor U5593 (N_5593,N_5157,N_5004);
xor U5594 (N_5594,N_5204,N_5267);
nand U5595 (N_5595,N_5308,N_5311);
nand U5596 (N_5596,N_5379,N_5192);
xnor U5597 (N_5597,N_5452,N_5347);
and U5598 (N_5598,N_5169,N_5199);
nand U5599 (N_5599,N_5307,N_5451);
nor U5600 (N_5600,N_5382,N_5268);
xnor U5601 (N_5601,N_5131,N_5039);
and U5602 (N_5602,N_5111,N_5265);
and U5603 (N_5603,N_5042,N_5183);
nand U5604 (N_5604,N_5399,N_5271);
nor U5605 (N_5605,N_5234,N_5100);
nand U5606 (N_5606,N_5071,N_5037);
and U5607 (N_5607,N_5490,N_5195);
nand U5608 (N_5608,N_5022,N_5016);
nor U5609 (N_5609,N_5380,N_5143);
or U5610 (N_5610,N_5141,N_5446);
nand U5611 (N_5611,N_5021,N_5174);
xnor U5612 (N_5612,N_5172,N_5414);
nor U5613 (N_5613,N_5315,N_5471);
nand U5614 (N_5614,N_5095,N_5146);
nor U5615 (N_5615,N_5327,N_5295);
and U5616 (N_5616,N_5391,N_5285);
and U5617 (N_5617,N_5133,N_5048);
xor U5618 (N_5618,N_5256,N_5494);
nand U5619 (N_5619,N_5426,N_5043);
xnor U5620 (N_5620,N_5249,N_5002);
and U5621 (N_5621,N_5349,N_5114);
xnor U5622 (N_5622,N_5352,N_5317);
or U5623 (N_5623,N_5323,N_5000);
nor U5624 (N_5624,N_5424,N_5171);
or U5625 (N_5625,N_5166,N_5261);
or U5626 (N_5626,N_5493,N_5178);
and U5627 (N_5627,N_5070,N_5034);
or U5628 (N_5628,N_5090,N_5198);
nand U5629 (N_5629,N_5225,N_5170);
nor U5630 (N_5630,N_5003,N_5134);
nor U5631 (N_5631,N_5345,N_5109);
xor U5632 (N_5632,N_5106,N_5033);
nand U5633 (N_5633,N_5469,N_5217);
or U5634 (N_5634,N_5075,N_5063);
nor U5635 (N_5635,N_5470,N_5245);
xor U5636 (N_5636,N_5147,N_5284);
nand U5637 (N_5637,N_5044,N_5089);
nand U5638 (N_5638,N_5061,N_5221);
xnor U5639 (N_5639,N_5491,N_5011);
and U5640 (N_5640,N_5083,N_5113);
xor U5641 (N_5641,N_5023,N_5275);
nor U5642 (N_5642,N_5082,N_5309);
and U5643 (N_5643,N_5208,N_5412);
nor U5644 (N_5644,N_5383,N_5099);
xnor U5645 (N_5645,N_5269,N_5403);
and U5646 (N_5646,N_5314,N_5218);
or U5647 (N_5647,N_5179,N_5121);
or U5648 (N_5648,N_5005,N_5124);
and U5649 (N_5649,N_5394,N_5474);
and U5650 (N_5650,N_5196,N_5220);
nor U5651 (N_5651,N_5009,N_5257);
or U5652 (N_5652,N_5283,N_5259);
nand U5653 (N_5653,N_5255,N_5137);
nor U5654 (N_5654,N_5007,N_5097);
nand U5655 (N_5655,N_5073,N_5096);
nand U5656 (N_5656,N_5356,N_5448);
nand U5657 (N_5657,N_5294,N_5300);
nor U5658 (N_5658,N_5270,N_5304);
xor U5659 (N_5659,N_5223,N_5418);
xnor U5660 (N_5660,N_5076,N_5046);
nor U5661 (N_5661,N_5473,N_5318);
or U5662 (N_5662,N_5463,N_5321);
nand U5663 (N_5663,N_5324,N_5105);
nor U5664 (N_5664,N_5351,N_5405);
or U5665 (N_5665,N_5164,N_5262);
xnor U5666 (N_5666,N_5483,N_5084);
or U5667 (N_5667,N_5040,N_5205);
xor U5668 (N_5668,N_5246,N_5086);
or U5669 (N_5669,N_5236,N_5026);
and U5670 (N_5670,N_5273,N_5138);
xor U5671 (N_5671,N_5162,N_5122);
or U5672 (N_5672,N_5212,N_5415);
and U5673 (N_5673,N_5453,N_5001);
nor U5674 (N_5674,N_5425,N_5219);
xor U5675 (N_5675,N_5216,N_5460);
or U5676 (N_5676,N_5476,N_5116);
or U5677 (N_5677,N_5363,N_5060);
nor U5678 (N_5678,N_5127,N_5287);
or U5679 (N_5679,N_5369,N_5279);
nand U5680 (N_5680,N_5455,N_5281);
and U5681 (N_5681,N_5056,N_5018);
and U5682 (N_5682,N_5115,N_5180);
or U5683 (N_5683,N_5376,N_5487);
xnor U5684 (N_5684,N_5334,N_5366);
nor U5685 (N_5685,N_5165,N_5340);
xor U5686 (N_5686,N_5241,N_5296);
or U5687 (N_5687,N_5067,N_5411);
and U5688 (N_5688,N_5064,N_5419);
or U5689 (N_5689,N_5154,N_5126);
or U5690 (N_5690,N_5434,N_5224);
and U5691 (N_5691,N_5291,N_5344);
xnor U5692 (N_5692,N_5078,N_5371);
nor U5693 (N_5693,N_5152,N_5093);
xnor U5694 (N_5694,N_5364,N_5423);
nor U5695 (N_5695,N_5015,N_5181);
or U5696 (N_5696,N_5210,N_5413);
and U5697 (N_5697,N_5186,N_5450);
nor U5698 (N_5698,N_5187,N_5387);
xor U5699 (N_5699,N_5461,N_5132);
or U5700 (N_5700,N_5362,N_5233);
nor U5701 (N_5701,N_5228,N_5014);
xor U5702 (N_5702,N_5161,N_5190);
xor U5703 (N_5703,N_5006,N_5456);
and U5704 (N_5704,N_5250,N_5497);
nand U5705 (N_5705,N_5025,N_5338);
or U5706 (N_5706,N_5074,N_5449);
and U5707 (N_5707,N_5239,N_5098);
xor U5708 (N_5708,N_5087,N_5136);
nand U5709 (N_5709,N_5393,N_5378);
or U5710 (N_5710,N_5135,N_5254);
nor U5711 (N_5711,N_5226,N_5054);
xor U5712 (N_5712,N_5160,N_5438);
or U5713 (N_5713,N_5209,N_5062);
xnor U5714 (N_5714,N_5193,N_5292);
nand U5715 (N_5715,N_5475,N_5467);
or U5716 (N_5716,N_5336,N_5333);
and U5717 (N_5717,N_5222,N_5341);
and U5718 (N_5718,N_5163,N_5117);
nand U5719 (N_5719,N_5059,N_5118);
xnor U5720 (N_5720,N_5189,N_5353);
nand U5721 (N_5721,N_5125,N_5120);
xor U5722 (N_5722,N_5243,N_5263);
nor U5723 (N_5723,N_5354,N_5274);
and U5724 (N_5724,N_5088,N_5266);
and U5725 (N_5725,N_5477,N_5319);
and U5726 (N_5726,N_5144,N_5017);
and U5727 (N_5727,N_5440,N_5072);
xnor U5728 (N_5728,N_5173,N_5159);
nor U5729 (N_5729,N_5103,N_5302);
xnor U5730 (N_5730,N_5464,N_5439);
xor U5731 (N_5731,N_5443,N_5248);
nand U5732 (N_5732,N_5397,N_5177);
xnor U5733 (N_5733,N_5079,N_5342);
or U5734 (N_5734,N_5320,N_5337);
nor U5735 (N_5735,N_5184,N_5066);
nand U5736 (N_5736,N_5101,N_5468);
nand U5737 (N_5737,N_5422,N_5049);
or U5738 (N_5738,N_5472,N_5139);
or U5739 (N_5739,N_5416,N_5408);
xnor U5740 (N_5740,N_5427,N_5421);
nand U5741 (N_5741,N_5498,N_5123);
and U5742 (N_5742,N_5055,N_5238);
nand U5743 (N_5743,N_5077,N_5102);
nor U5744 (N_5744,N_5365,N_5316);
nand U5745 (N_5745,N_5081,N_5242);
xnor U5746 (N_5746,N_5020,N_5488);
and U5747 (N_5747,N_5058,N_5028);
nor U5748 (N_5748,N_5481,N_5301);
nor U5749 (N_5749,N_5108,N_5156);
xnor U5750 (N_5750,N_5468,N_5093);
and U5751 (N_5751,N_5140,N_5384);
or U5752 (N_5752,N_5270,N_5057);
nand U5753 (N_5753,N_5150,N_5018);
and U5754 (N_5754,N_5253,N_5200);
nand U5755 (N_5755,N_5297,N_5448);
nor U5756 (N_5756,N_5108,N_5097);
or U5757 (N_5757,N_5313,N_5120);
xor U5758 (N_5758,N_5198,N_5046);
or U5759 (N_5759,N_5322,N_5246);
and U5760 (N_5760,N_5057,N_5122);
xnor U5761 (N_5761,N_5460,N_5059);
and U5762 (N_5762,N_5232,N_5459);
xnor U5763 (N_5763,N_5378,N_5244);
and U5764 (N_5764,N_5165,N_5292);
and U5765 (N_5765,N_5336,N_5226);
nor U5766 (N_5766,N_5245,N_5382);
xor U5767 (N_5767,N_5289,N_5276);
and U5768 (N_5768,N_5195,N_5072);
xnor U5769 (N_5769,N_5206,N_5462);
or U5770 (N_5770,N_5076,N_5340);
nor U5771 (N_5771,N_5055,N_5224);
or U5772 (N_5772,N_5086,N_5475);
and U5773 (N_5773,N_5292,N_5204);
xnor U5774 (N_5774,N_5421,N_5479);
or U5775 (N_5775,N_5306,N_5456);
and U5776 (N_5776,N_5014,N_5270);
and U5777 (N_5777,N_5113,N_5064);
or U5778 (N_5778,N_5330,N_5375);
and U5779 (N_5779,N_5358,N_5147);
nor U5780 (N_5780,N_5249,N_5212);
nand U5781 (N_5781,N_5425,N_5063);
or U5782 (N_5782,N_5092,N_5269);
or U5783 (N_5783,N_5337,N_5141);
or U5784 (N_5784,N_5311,N_5147);
xnor U5785 (N_5785,N_5196,N_5457);
nor U5786 (N_5786,N_5449,N_5399);
nand U5787 (N_5787,N_5171,N_5015);
or U5788 (N_5788,N_5460,N_5071);
nand U5789 (N_5789,N_5285,N_5061);
xor U5790 (N_5790,N_5220,N_5149);
or U5791 (N_5791,N_5170,N_5216);
xor U5792 (N_5792,N_5498,N_5381);
nand U5793 (N_5793,N_5476,N_5061);
and U5794 (N_5794,N_5390,N_5476);
and U5795 (N_5795,N_5381,N_5265);
nand U5796 (N_5796,N_5395,N_5392);
and U5797 (N_5797,N_5110,N_5026);
nand U5798 (N_5798,N_5394,N_5170);
nor U5799 (N_5799,N_5198,N_5453);
and U5800 (N_5800,N_5371,N_5265);
or U5801 (N_5801,N_5249,N_5194);
nand U5802 (N_5802,N_5345,N_5179);
xnor U5803 (N_5803,N_5322,N_5347);
and U5804 (N_5804,N_5292,N_5441);
nor U5805 (N_5805,N_5104,N_5201);
and U5806 (N_5806,N_5161,N_5289);
nor U5807 (N_5807,N_5445,N_5277);
xnor U5808 (N_5808,N_5429,N_5100);
nor U5809 (N_5809,N_5273,N_5123);
or U5810 (N_5810,N_5418,N_5230);
nor U5811 (N_5811,N_5328,N_5110);
nor U5812 (N_5812,N_5042,N_5437);
and U5813 (N_5813,N_5007,N_5314);
xnor U5814 (N_5814,N_5141,N_5310);
or U5815 (N_5815,N_5051,N_5054);
nand U5816 (N_5816,N_5486,N_5272);
or U5817 (N_5817,N_5052,N_5353);
xor U5818 (N_5818,N_5062,N_5001);
xor U5819 (N_5819,N_5212,N_5307);
nand U5820 (N_5820,N_5282,N_5100);
and U5821 (N_5821,N_5195,N_5046);
or U5822 (N_5822,N_5077,N_5140);
nand U5823 (N_5823,N_5020,N_5409);
nor U5824 (N_5824,N_5280,N_5151);
or U5825 (N_5825,N_5048,N_5027);
nor U5826 (N_5826,N_5485,N_5135);
nor U5827 (N_5827,N_5009,N_5299);
and U5828 (N_5828,N_5158,N_5129);
xnor U5829 (N_5829,N_5284,N_5074);
nor U5830 (N_5830,N_5257,N_5136);
nand U5831 (N_5831,N_5100,N_5440);
xnor U5832 (N_5832,N_5342,N_5151);
or U5833 (N_5833,N_5050,N_5474);
nand U5834 (N_5834,N_5449,N_5185);
or U5835 (N_5835,N_5129,N_5184);
nand U5836 (N_5836,N_5313,N_5243);
or U5837 (N_5837,N_5370,N_5344);
or U5838 (N_5838,N_5129,N_5043);
nor U5839 (N_5839,N_5354,N_5065);
and U5840 (N_5840,N_5493,N_5078);
or U5841 (N_5841,N_5290,N_5088);
xor U5842 (N_5842,N_5477,N_5157);
nand U5843 (N_5843,N_5295,N_5401);
nand U5844 (N_5844,N_5125,N_5026);
or U5845 (N_5845,N_5253,N_5294);
and U5846 (N_5846,N_5227,N_5130);
nor U5847 (N_5847,N_5046,N_5410);
nor U5848 (N_5848,N_5164,N_5395);
xnor U5849 (N_5849,N_5241,N_5374);
or U5850 (N_5850,N_5423,N_5408);
or U5851 (N_5851,N_5416,N_5498);
nor U5852 (N_5852,N_5382,N_5432);
nand U5853 (N_5853,N_5487,N_5046);
or U5854 (N_5854,N_5484,N_5367);
or U5855 (N_5855,N_5127,N_5290);
xor U5856 (N_5856,N_5104,N_5067);
nor U5857 (N_5857,N_5046,N_5466);
nand U5858 (N_5858,N_5331,N_5459);
nand U5859 (N_5859,N_5288,N_5303);
xor U5860 (N_5860,N_5281,N_5272);
xor U5861 (N_5861,N_5406,N_5224);
nor U5862 (N_5862,N_5427,N_5409);
xnor U5863 (N_5863,N_5329,N_5163);
and U5864 (N_5864,N_5027,N_5227);
nand U5865 (N_5865,N_5111,N_5247);
and U5866 (N_5866,N_5061,N_5499);
nand U5867 (N_5867,N_5220,N_5255);
or U5868 (N_5868,N_5174,N_5238);
and U5869 (N_5869,N_5476,N_5488);
or U5870 (N_5870,N_5139,N_5475);
nor U5871 (N_5871,N_5010,N_5269);
xor U5872 (N_5872,N_5071,N_5486);
nor U5873 (N_5873,N_5232,N_5355);
nor U5874 (N_5874,N_5403,N_5158);
or U5875 (N_5875,N_5347,N_5122);
nand U5876 (N_5876,N_5002,N_5473);
nand U5877 (N_5877,N_5434,N_5311);
or U5878 (N_5878,N_5365,N_5272);
nor U5879 (N_5879,N_5184,N_5082);
xnor U5880 (N_5880,N_5199,N_5109);
or U5881 (N_5881,N_5238,N_5493);
or U5882 (N_5882,N_5020,N_5499);
nand U5883 (N_5883,N_5129,N_5297);
nor U5884 (N_5884,N_5020,N_5173);
or U5885 (N_5885,N_5393,N_5232);
nand U5886 (N_5886,N_5166,N_5111);
nand U5887 (N_5887,N_5305,N_5049);
nand U5888 (N_5888,N_5468,N_5221);
xnor U5889 (N_5889,N_5078,N_5081);
nor U5890 (N_5890,N_5395,N_5071);
and U5891 (N_5891,N_5140,N_5021);
xor U5892 (N_5892,N_5241,N_5176);
xnor U5893 (N_5893,N_5374,N_5279);
nor U5894 (N_5894,N_5218,N_5477);
nor U5895 (N_5895,N_5376,N_5275);
nor U5896 (N_5896,N_5038,N_5456);
nand U5897 (N_5897,N_5314,N_5381);
xnor U5898 (N_5898,N_5403,N_5476);
nand U5899 (N_5899,N_5418,N_5006);
nand U5900 (N_5900,N_5266,N_5379);
nand U5901 (N_5901,N_5118,N_5116);
and U5902 (N_5902,N_5258,N_5079);
and U5903 (N_5903,N_5373,N_5122);
xnor U5904 (N_5904,N_5370,N_5459);
or U5905 (N_5905,N_5353,N_5028);
and U5906 (N_5906,N_5100,N_5069);
and U5907 (N_5907,N_5429,N_5467);
nand U5908 (N_5908,N_5027,N_5120);
nand U5909 (N_5909,N_5392,N_5010);
and U5910 (N_5910,N_5092,N_5289);
nor U5911 (N_5911,N_5246,N_5478);
xnor U5912 (N_5912,N_5038,N_5208);
or U5913 (N_5913,N_5316,N_5099);
xor U5914 (N_5914,N_5050,N_5334);
nor U5915 (N_5915,N_5169,N_5181);
and U5916 (N_5916,N_5274,N_5471);
nand U5917 (N_5917,N_5343,N_5326);
or U5918 (N_5918,N_5180,N_5295);
and U5919 (N_5919,N_5434,N_5064);
or U5920 (N_5920,N_5448,N_5008);
or U5921 (N_5921,N_5032,N_5016);
and U5922 (N_5922,N_5161,N_5387);
nor U5923 (N_5923,N_5002,N_5253);
nand U5924 (N_5924,N_5455,N_5306);
and U5925 (N_5925,N_5233,N_5236);
xor U5926 (N_5926,N_5431,N_5002);
or U5927 (N_5927,N_5179,N_5101);
and U5928 (N_5928,N_5238,N_5029);
nand U5929 (N_5929,N_5057,N_5042);
nand U5930 (N_5930,N_5104,N_5054);
xnor U5931 (N_5931,N_5195,N_5439);
or U5932 (N_5932,N_5118,N_5114);
nor U5933 (N_5933,N_5484,N_5360);
and U5934 (N_5934,N_5352,N_5150);
xor U5935 (N_5935,N_5017,N_5364);
nor U5936 (N_5936,N_5244,N_5349);
or U5937 (N_5937,N_5331,N_5219);
xnor U5938 (N_5938,N_5205,N_5471);
nand U5939 (N_5939,N_5221,N_5489);
or U5940 (N_5940,N_5391,N_5433);
and U5941 (N_5941,N_5369,N_5433);
nor U5942 (N_5942,N_5146,N_5171);
nor U5943 (N_5943,N_5059,N_5179);
and U5944 (N_5944,N_5022,N_5002);
or U5945 (N_5945,N_5312,N_5077);
nor U5946 (N_5946,N_5017,N_5478);
nor U5947 (N_5947,N_5358,N_5392);
or U5948 (N_5948,N_5107,N_5366);
and U5949 (N_5949,N_5472,N_5268);
nand U5950 (N_5950,N_5481,N_5391);
and U5951 (N_5951,N_5390,N_5193);
nor U5952 (N_5952,N_5221,N_5127);
nand U5953 (N_5953,N_5286,N_5371);
nand U5954 (N_5954,N_5416,N_5467);
nand U5955 (N_5955,N_5315,N_5386);
or U5956 (N_5956,N_5381,N_5000);
nor U5957 (N_5957,N_5349,N_5182);
xor U5958 (N_5958,N_5303,N_5325);
xnor U5959 (N_5959,N_5210,N_5464);
xnor U5960 (N_5960,N_5035,N_5355);
or U5961 (N_5961,N_5159,N_5247);
nand U5962 (N_5962,N_5235,N_5405);
xor U5963 (N_5963,N_5298,N_5183);
xor U5964 (N_5964,N_5065,N_5279);
and U5965 (N_5965,N_5269,N_5455);
xnor U5966 (N_5966,N_5265,N_5341);
and U5967 (N_5967,N_5371,N_5030);
or U5968 (N_5968,N_5048,N_5254);
nor U5969 (N_5969,N_5369,N_5354);
xor U5970 (N_5970,N_5207,N_5201);
or U5971 (N_5971,N_5173,N_5272);
xor U5972 (N_5972,N_5424,N_5305);
or U5973 (N_5973,N_5195,N_5084);
nor U5974 (N_5974,N_5497,N_5373);
nor U5975 (N_5975,N_5407,N_5339);
nor U5976 (N_5976,N_5109,N_5412);
xnor U5977 (N_5977,N_5245,N_5293);
nand U5978 (N_5978,N_5340,N_5407);
xor U5979 (N_5979,N_5109,N_5449);
nor U5980 (N_5980,N_5169,N_5007);
nand U5981 (N_5981,N_5090,N_5491);
or U5982 (N_5982,N_5220,N_5114);
nand U5983 (N_5983,N_5072,N_5124);
xor U5984 (N_5984,N_5381,N_5232);
xnor U5985 (N_5985,N_5291,N_5217);
or U5986 (N_5986,N_5189,N_5301);
xor U5987 (N_5987,N_5456,N_5373);
nand U5988 (N_5988,N_5173,N_5028);
nor U5989 (N_5989,N_5458,N_5327);
and U5990 (N_5990,N_5417,N_5241);
or U5991 (N_5991,N_5079,N_5293);
and U5992 (N_5992,N_5175,N_5498);
xnor U5993 (N_5993,N_5086,N_5155);
xnor U5994 (N_5994,N_5355,N_5470);
nand U5995 (N_5995,N_5240,N_5018);
nor U5996 (N_5996,N_5455,N_5199);
nor U5997 (N_5997,N_5268,N_5042);
nor U5998 (N_5998,N_5454,N_5468);
xnor U5999 (N_5999,N_5459,N_5187);
xnor U6000 (N_6000,N_5845,N_5652);
xnor U6001 (N_6001,N_5911,N_5964);
nand U6002 (N_6002,N_5857,N_5963);
xor U6003 (N_6003,N_5751,N_5633);
nor U6004 (N_6004,N_5916,N_5691);
and U6005 (N_6005,N_5664,N_5820);
nand U6006 (N_6006,N_5680,N_5665);
nor U6007 (N_6007,N_5979,N_5807);
or U6008 (N_6008,N_5802,N_5954);
xor U6009 (N_6009,N_5611,N_5959);
xor U6010 (N_6010,N_5697,N_5658);
or U6011 (N_6011,N_5726,N_5672);
or U6012 (N_6012,N_5733,N_5705);
xor U6013 (N_6013,N_5772,N_5773);
nand U6014 (N_6014,N_5581,N_5529);
and U6015 (N_6015,N_5592,N_5923);
or U6016 (N_6016,N_5739,N_5595);
nor U6017 (N_6017,N_5904,N_5943);
nor U6018 (N_6018,N_5747,N_5885);
or U6019 (N_6019,N_5644,N_5789);
and U6020 (N_6020,N_5610,N_5525);
xnor U6021 (N_6021,N_5559,N_5537);
nor U6022 (N_6022,N_5850,N_5908);
nor U6023 (N_6023,N_5765,N_5735);
nor U6024 (N_6024,N_5939,N_5626);
nor U6025 (N_6025,N_5686,N_5915);
nand U6026 (N_6026,N_5841,N_5783);
or U6027 (N_6027,N_5758,N_5986);
nand U6028 (N_6028,N_5548,N_5565);
or U6029 (N_6029,N_5708,N_5724);
nor U6030 (N_6030,N_5641,N_5897);
and U6031 (N_6031,N_5893,N_5771);
and U6032 (N_6032,N_5585,N_5926);
or U6033 (N_6033,N_5945,N_5865);
and U6034 (N_6034,N_5669,N_5535);
xor U6035 (N_6035,N_5952,N_5949);
xor U6036 (N_6036,N_5696,N_5929);
nor U6037 (N_6037,N_5987,N_5609);
xor U6038 (N_6038,N_5598,N_5554);
xnor U6039 (N_6039,N_5822,N_5709);
nand U6040 (N_6040,N_5524,N_5511);
or U6041 (N_6041,N_5689,N_5608);
xnor U6042 (N_6042,N_5871,N_5973);
nand U6043 (N_6043,N_5536,N_5702);
nor U6044 (N_6044,N_5936,N_5994);
and U6045 (N_6045,N_5571,N_5797);
or U6046 (N_6046,N_5599,N_5970);
nand U6047 (N_6047,N_5553,N_5866);
nor U6048 (N_6048,N_5882,N_5587);
and U6049 (N_6049,N_5606,N_5942);
and U6050 (N_6050,N_5920,N_5740);
or U6051 (N_6051,N_5748,N_5806);
and U6052 (N_6052,N_5619,N_5519);
xnor U6053 (N_6053,N_5584,N_5918);
xnor U6054 (N_6054,N_5564,N_5552);
nand U6055 (N_6055,N_5960,N_5951);
and U6056 (N_6056,N_5907,N_5779);
nand U6057 (N_6057,N_5539,N_5812);
or U6058 (N_6058,N_5622,N_5925);
nand U6059 (N_6059,N_5732,N_5794);
and U6060 (N_6060,N_5900,N_5505);
or U6061 (N_6061,N_5870,N_5764);
nor U6062 (N_6062,N_5543,N_5744);
nand U6063 (N_6063,N_5905,N_5769);
xor U6064 (N_6064,N_5984,N_5588);
nor U6065 (N_6065,N_5755,N_5815);
nor U6066 (N_6066,N_5913,N_5808);
xor U6067 (N_6067,N_5766,N_5995);
nand U6068 (N_6068,N_5506,N_5837);
xnor U6069 (N_6069,N_5714,N_5736);
or U6070 (N_6070,N_5583,N_5607);
xor U6071 (N_6071,N_5863,N_5706);
xnor U6072 (N_6072,N_5650,N_5823);
and U6073 (N_6073,N_5924,N_5563);
xnor U6074 (N_6074,N_5731,N_5701);
and U6075 (N_6075,N_5629,N_5778);
and U6076 (N_6076,N_5813,N_5946);
nand U6077 (N_6077,N_5781,N_5886);
or U6078 (N_6078,N_5958,N_5544);
or U6079 (N_6079,N_5613,N_5874);
and U6080 (N_6080,N_5788,N_5528);
and U6081 (N_6081,N_5504,N_5522);
or U6082 (N_6082,N_5884,N_5551);
and U6083 (N_6083,N_5627,N_5657);
nand U6084 (N_6084,N_5903,N_5743);
or U6085 (N_6085,N_5558,N_5877);
or U6086 (N_6086,N_5694,N_5892);
or U6087 (N_6087,N_5785,N_5547);
nor U6088 (N_6088,N_5621,N_5967);
nand U6089 (N_6089,N_5719,N_5844);
nand U6090 (N_6090,N_5555,N_5809);
or U6091 (N_6091,N_5717,N_5759);
nand U6092 (N_6092,N_5966,N_5508);
and U6093 (N_6093,N_5947,N_5515);
or U6094 (N_6094,N_5600,N_5521);
or U6095 (N_6095,N_5612,N_5763);
nand U6096 (N_6096,N_5941,N_5533);
or U6097 (N_6097,N_5927,N_5725);
or U6098 (N_6098,N_5989,N_5974);
or U6099 (N_6099,N_5881,N_5721);
xnor U6100 (N_6100,N_5957,N_5562);
xnor U6101 (N_6101,N_5860,N_5596);
nand U6102 (N_6102,N_5969,N_5604);
nand U6103 (N_6103,N_5878,N_5898);
xnor U6104 (N_6104,N_5617,N_5512);
xnor U6105 (N_6105,N_5998,N_5623);
nand U6106 (N_6106,N_5741,N_5711);
xor U6107 (N_6107,N_5757,N_5560);
and U6108 (N_6108,N_5668,N_5527);
xor U6109 (N_6109,N_5990,N_5568);
nor U6110 (N_6110,N_5688,N_5876);
or U6111 (N_6111,N_5981,N_5654);
or U6112 (N_6112,N_5997,N_5780);
nand U6113 (N_6113,N_5513,N_5591);
nand U6114 (N_6114,N_5695,N_5909);
nand U6115 (N_6115,N_5687,N_5753);
nor U6116 (N_6116,N_5832,N_5645);
or U6117 (N_6117,N_5854,N_5602);
or U6118 (N_6118,N_5932,N_5566);
nor U6119 (N_6119,N_5700,N_5821);
and U6120 (N_6120,N_5526,N_5935);
nand U6121 (N_6121,N_5569,N_5578);
nor U6122 (N_6122,N_5514,N_5840);
nor U6123 (N_6123,N_5576,N_5985);
or U6124 (N_6124,N_5872,N_5727);
and U6125 (N_6125,N_5589,N_5638);
xnor U6126 (N_6126,N_5729,N_5518);
and U6127 (N_6127,N_5679,N_5503);
nand U6128 (N_6128,N_5805,N_5673);
nand U6129 (N_6129,N_5646,N_5856);
xor U6130 (N_6130,N_5698,N_5570);
and U6131 (N_6131,N_5710,N_5507);
nor U6132 (N_6132,N_5746,N_5824);
nor U6133 (N_6133,N_5800,N_5699);
nor U6134 (N_6134,N_5858,N_5894);
xnor U6135 (N_6135,N_5540,N_5676);
and U6136 (N_6136,N_5742,N_5752);
nand U6137 (N_6137,N_5520,N_5628);
xnor U6138 (N_6138,N_5501,N_5605);
nor U6139 (N_6139,N_5980,N_5715);
nor U6140 (N_6140,N_5816,N_5818);
or U6141 (N_6141,N_5579,N_5827);
nor U6142 (N_6142,N_5948,N_5692);
and U6143 (N_6143,N_5983,N_5712);
xnor U6144 (N_6144,N_5713,N_5671);
or U6145 (N_6145,N_5851,N_5685);
and U6146 (N_6146,N_5843,N_5546);
and U6147 (N_6147,N_5594,N_5636);
and U6148 (N_6148,N_5683,N_5879);
and U6149 (N_6149,N_5745,N_5653);
xnor U6150 (N_6150,N_5933,N_5848);
and U6151 (N_6151,N_5649,N_5760);
or U6152 (N_6152,N_5928,N_5775);
nor U6153 (N_6153,N_5573,N_5965);
and U6154 (N_6154,N_5756,N_5718);
xnor U6155 (N_6155,N_5834,N_5867);
and U6156 (N_6156,N_5722,N_5978);
nand U6157 (N_6157,N_5557,N_5703);
xnor U6158 (N_6158,N_5922,N_5919);
or U6159 (N_6159,N_5620,N_5762);
xnor U6160 (N_6160,N_5982,N_5639);
xnor U6161 (N_6161,N_5906,N_5864);
nand U6162 (N_6162,N_5890,N_5798);
nand U6163 (N_6163,N_5660,N_5853);
xnor U6164 (N_6164,N_5852,N_5632);
nand U6165 (N_6165,N_5791,N_5561);
nand U6166 (N_6166,N_5647,N_5795);
xor U6167 (N_6167,N_5869,N_5835);
xnor U6168 (N_6168,N_5681,N_5754);
and U6169 (N_6169,N_5517,N_5530);
and U6170 (N_6170,N_5531,N_5901);
xnor U6171 (N_6171,N_5817,N_5782);
xnor U6172 (N_6172,N_5663,N_5784);
and U6173 (N_6173,N_5545,N_5804);
or U6174 (N_6174,N_5938,N_5801);
and U6175 (N_6175,N_5770,N_5899);
nor U6176 (N_6176,N_5937,N_5625);
or U6177 (N_6177,N_5593,N_5955);
or U6178 (N_6178,N_5988,N_5829);
xor U6179 (N_6179,N_5643,N_5577);
or U6180 (N_6180,N_5953,N_5761);
xor U6181 (N_6181,N_5793,N_5950);
xnor U6182 (N_6182,N_5931,N_5614);
nor U6183 (N_6183,N_5895,N_5693);
nor U6184 (N_6184,N_5831,N_5883);
or U6185 (N_6185,N_5523,N_5634);
nand U6186 (N_6186,N_5737,N_5930);
nor U6187 (N_6187,N_5637,N_5640);
or U6188 (N_6188,N_5532,N_5912);
or U6189 (N_6189,N_5534,N_5855);
nor U6190 (N_6190,N_5655,N_5842);
xor U6191 (N_6191,N_5846,N_5509);
nor U6192 (N_6192,N_5549,N_5723);
nor U6193 (N_6193,N_5580,N_5999);
nand U6194 (N_6194,N_5738,N_5968);
and U6195 (N_6195,N_5648,N_5510);
or U6196 (N_6196,N_5572,N_5861);
nor U6197 (N_6197,N_5944,N_5830);
nor U6198 (N_6198,N_5992,N_5811);
xnor U6199 (N_6199,N_5796,N_5684);
nor U6200 (N_6200,N_5790,N_5888);
xnor U6201 (N_6201,N_5889,N_5616);
xor U6202 (N_6202,N_5838,N_5993);
or U6203 (N_6203,N_5961,N_5603);
and U6204 (N_6204,N_5971,N_5690);
and U6205 (N_6205,N_5662,N_5792);
and U6206 (N_6206,N_5873,N_5996);
nor U6207 (N_6207,N_5656,N_5975);
nor U6208 (N_6208,N_5910,N_5902);
and U6209 (N_6209,N_5674,N_5538);
nor U6210 (N_6210,N_5749,N_5777);
nor U6211 (N_6211,N_5836,N_5720);
or U6212 (N_6212,N_5839,N_5618);
nand U6213 (N_6213,N_5972,N_5887);
nand U6214 (N_6214,N_5768,N_5917);
nor U6215 (N_6215,N_5776,N_5819);
xor U6216 (N_6216,N_5875,N_5859);
xor U6217 (N_6217,N_5976,N_5601);
nor U6218 (N_6218,N_5849,N_5635);
or U6219 (N_6219,N_5582,N_5574);
and U6220 (N_6220,N_5586,N_5728);
or U6221 (N_6221,N_5734,N_5707);
nand U6222 (N_6222,N_5541,N_5624);
nand U6223 (N_6223,N_5550,N_5934);
xnor U6224 (N_6224,N_5730,N_5940);
and U6225 (N_6225,N_5651,N_5991);
nand U6226 (N_6226,N_5828,N_5677);
and U6227 (N_6227,N_5962,N_5921);
nand U6228 (N_6228,N_5704,N_5787);
and U6229 (N_6229,N_5615,N_5659);
xor U6230 (N_6230,N_5678,N_5826);
nor U6231 (N_6231,N_5667,N_5767);
and U6232 (N_6232,N_5810,N_5750);
and U6233 (N_6233,N_5642,N_5880);
xor U6234 (N_6234,N_5575,N_5670);
nor U6235 (N_6235,N_5891,N_5774);
or U6236 (N_6236,N_5661,N_5847);
and U6237 (N_6237,N_5799,N_5825);
xor U6238 (N_6238,N_5500,N_5786);
nand U6239 (N_6239,N_5956,N_5675);
and U6240 (N_6240,N_5630,N_5716);
nor U6241 (N_6241,N_5682,N_5833);
and U6242 (N_6242,N_5590,N_5862);
nor U6243 (N_6243,N_5914,N_5516);
nand U6244 (N_6244,N_5803,N_5814);
or U6245 (N_6245,N_5542,N_5567);
nor U6246 (N_6246,N_5597,N_5977);
xor U6247 (N_6247,N_5868,N_5666);
xnor U6248 (N_6248,N_5631,N_5896);
or U6249 (N_6249,N_5556,N_5502);
or U6250 (N_6250,N_5918,N_5925);
nand U6251 (N_6251,N_5595,N_5668);
nor U6252 (N_6252,N_5919,N_5807);
xor U6253 (N_6253,N_5905,N_5988);
nor U6254 (N_6254,N_5936,N_5963);
nand U6255 (N_6255,N_5748,N_5885);
nand U6256 (N_6256,N_5922,N_5657);
nand U6257 (N_6257,N_5699,N_5665);
nor U6258 (N_6258,N_5941,N_5834);
nand U6259 (N_6259,N_5639,N_5905);
or U6260 (N_6260,N_5636,N_5697);
nor U6261 (N_6261,N_5603,N_5746);
and U6262 (N_6262,N_5685,N_5649);
or U6263 (N_6263,N_5515,N_5942);
nand U6264 (N_6264,N_5671,N_5796);
nand U6265 (N_6265,N_5982,N_5917);
nor U6266 (N_6266,N_5806,N_5721);
nand U6267 (N_6267,N_5947,N_5802);
nor U6268 (N_6268,N_5554,N_5868);
nor U6269 (N_6269,N_5753,N_5870);
nand U6270 (N_6270,N_5920,N_5652);
and U6271 (N_6271,N_5501,N_5875);
nand U6272 (N_6272,N_5572,N_5868);
nor U6273 (N_6273,N_5642,N_5631);
and U6274 (N_6274,N_5732,N_5932);
xor U6275 (N_6275,N_5556,N_5805);
and U6276 (N_6276,N_5752,N_5976);
or U6277 (N_6277,N_5992,N_5876);
nor U6278 (N_6278,N_5647,N_5823);
nand U6279 (N_6279,N_5594,N_5743);
or U6280 (N_6280,N_5865,N_5981);
or U6281 (N_6281,N_5619,N_5755);
nand U6282 (N_6282,N_5680,N_5841);
nand U6283 (N_6283,N_5687,N_5706);
nor U6284 (N_6284,N_5847,N_5675);
or U6285 (N_6285,N_5898,N_5755);
nor U6286 (N_6286,N_5525,N_5869);
xnor U6287 (N_6287,N_5850,N_5985);
nor U6288 (N_6288,N_5668,N_5902);
nor U6289 (N_6289,N_5982,N_5790);
nand U6290 (N_6290,N_5593,N_5963);
nor U6291 (N_6291,N_5724,N_5742);
xor U6292 (N_6292,N_5659,N_5939);
and U6293 (N_6293,N_5565,N_5594);
and U6294 (N_6294,N_5516,N_5570);
or U6295 (N_6295,N_5684,N_5801);
nand U6296 (N_6296,N_5961,N_5827);
xnor U6297 (N_6297,N_5670,N_5508);
and U6298 (N_6298,N_5805,N_5953);
or U6299 (N_6299,N_5543,N_5848);
nand U6300 (N_6300,N_5756,N_5592);
or U6301 (N_6301,N_5658,N_5728);
nand U6302 (N_6302,N_5618,N_5979);
xor U6303 (N_6303,N_5841,N_5960);
or U6304 (N_6304,N_5702,N_5616);
or U6305 (N_6305,N_5608,N_5856);
nor U6306 (N_6306,N_5572,N_5574);
xor U6307 (N_6307,N_5919,N_5525);
xnor U6308 (N_6308,N_5934,N_5743);
nor U6309 (N_6309,N_5858,N_5972);
xnor U6310 (N_6310,N_5868,N_5899);
nand U6311 (N_6311,N_5687,N_5540);
and U6312 (N_6312,N_5655,N_5893);
xor U6313 (N_6313,N_5791,N_5721);
xor U6314 (N_6314,N_5734,N_5747);
xnor U6315 (N_6315,N_5500,N_5584);
nor U6316 (N_6316,N_5780,N_5869);
and U6317 (N_6317,N_5670,N_5553);
nor U6318 (N_6318,N_5874,N_5718);
xnor U6319 (N_6319,N_5771,N_5665);
and U6320 (N_6320,N_5936,N_5688);
nand U6321 (N_6321,N_5620,N_5696);
or U6322 (N_6322,N_5753,N_5598);
nor U6323 (N_6323,N_5855,N_5705);
nand U6324 (N_6324,N_5720,N_5675);
xnor U6325 (N_6325,N_5966,N_5983);
or U6326 (N_6326,N_5685,N_5869);
nand U6327 (N_6327,N_5613,N_5816);
nand U6328 (N_6328,N_5915,N_5522);
or U6329 (N_6329,N_5882,N_5890);
nor U6330 (N_6330,N_5884,N_5645);
and U6331 (N_6331,N_5707,N_5731);
xnor U6332 (N_6332,N_5687,N_5996);
nand U6333 (N_6333,N_5639,N_5868);
nand U6334 (N_6334,N_5802,N_5818);
nand U6335 (N_6335,N_5706,N_5882);
xnor U6336 (N_6336,N_5535,N_5987);
xor U6337 (N_6337,N_5868,N_5892);
xnor U6338 (N_6338,N_5521,N_5982);
and U6339 (N_6339,N_5816,N_5840);
and U6340 (N_6340,N_5828,N_5918);
or U6341 (N_6341,N_5583,N_5762);
nand U6342 (N_6342,N_5818,N_5734);
nand U6343 (N_6343,N_5555,N_5949);
xor U6344 (N_6344,N_5898,N_5529);
nand U6345 (N_6345,N_5544,N_5943);
xnor U6346 (N_6346,N_5522,N_5802);
or U6347 (N_6347,N_5709,N_5510);
nor U6348 (N_6348,N_5699,N_5957);
nor U6349 (N_6349,N_5894,N_5826);
nand U6350 (N_6350,N_5945,N_5544);
or U6351 (N_6351,N_5686,N_5731);
or U6352 (N_6352,N_5889,N_5981);
nand U6353 (N_6353,N_5508,N_5748);
nor U6354 (N_6354,N_5591,N_5784);
nor U6355 (N_6355,N_5819,N_5667);
nor U6356 (N_6356,N_5851,N_5582);
nor U6357 (N_6357,N_5710,N_5601);
nor U6358 (N_6358,N_5806,N_5589);
nor U6359 (N_6359,N_5879,N_5894);
nor U6360 (N_6360,N_5918,N_5950);
nand U6361 (N_6361,N_5923,N_5685);
nor U6362 (N_6362,N_5874,N_5755);
nor U6363 (N_6363,N_5739,N_5533);
and U6364 (N_6364,N_5528,N_5632);
or U6365 (N_6365,N_5932,N_5558);
xnor U6366 (N_6366,N_5714,N_5589);
or U6367 (N_6367,N_5915,N_5753);
or U6368 (N_6368,N_5716,N_5951);
nand U6369 (N_6369,N_5863,N_5776);
xor U6370 (N_6370,N_5611,N_5989);
nand U6371 (N_6371,N_5938,N_5985);
nand U6372 (N_6372,N_5801,N_5515);
xnor U6373 (N_6373,N_5522,N_5948);
xor U6374 (N_6374,N_5634,N_5552);
nand U6375 (N_6375,N_5969,N_5887);
and U6376 (N_6376,N_5734,N_5530);
nand U6377 (N_6377,N_5587,N_5758);
nor U6378 (N_6378,N_5648,N_5574);
and U6379 (N_6379,N_5632,N_5782);
nand U6380 (N_6380,N_5675,N_5610);
xnor U6381 (N_6381,N_5634,N_5525);
or U6382 (N_6382,N_5831,N_5818);
or U6383 (N_6383,N_5971,N_5949);
nor U6384 (N_6384,N_5646,N_5870);
nor U6385 (N_6385,N_5558,N_5632);
or U6386 (N_6386,N_5983,N_5943);
nor U6387 (N_6387,N_5951,N_5617);
and U6388 (N_6388,N_5806,N_5764);
or U6389 (N_6389,N_5694,N_5804);
nand U6390 (N_6390,N_5521,N_5867);
and U6391 (N_6391,N_5967,N_5564);
nor U6392 (N_6392,N_5594,N_5912);
or U6393 (N_6393,N_5542,N_5504);
xor U6394 (N_6394,N_5726,N_5615);
nor U6395 (N_6395,N_5879,N_5636);
nor U6396 (N_6396,N_5883,N_5752);
nor U6397 (N_6397,N_5878,N_5751);
nor U6398 (N_6398,N_5571,N_5746);
nor U6399 (N_6399,N_5912,N_5609);
nand U6400 (N_6400,N_5556,N_5667);
or U6401 (N_6401,N_5857,N_5979);
nand U6402 (N_6402,N_5514,N_5543);
and U6403 (N_6403,N_5782,N_5556);
and U6404 (N_6404,N_5773,N_5661);
xor U6405 (N_6405,N_5737,N_5613);
or U6406 (N_6406,N_5680,N_5700);
and U6407 (N_6407,N_5717,N_5747);
nor U6408 (N_6408,N_5878,N_5993);
or U6409 (N_6409,N_5968,N_5649);
nand U6410 (N_6410,N_5653,N_5500);
nor U6411 (N_6411,N_5514,N_5541);
and U6412 (N_6412,N_5723,N_5711);
and U6413 (N_6413,N_5944,N_5533);
xor U6414 (N_6414,N_5906,N_5603);
and U6415 (N_6415,N_5756,N_5608);
nand U6416 (N_6416,N_5702,N_5810);
and U6417 (N_6417,N_5527,N_5888);
xor U6418 (N_6418,N_5616,N_5874);
nand U6419 (N_6419,N_5817,N_5524);
nor U6420 (N_6420,N_5571,N_5951);
xnor U6421 (N_6421,N_5556,N_5959);
and U6422 (N_6422,N_5947,N_5984);
xor U6423 (N_6423,N_5811,N_5529);
nor U6424 (N_6424,N_5954,N_5758);
and U6425 (N_6425,N_5955,N_5887);
or U6426 (N_6426,N_5935,N_5864);
or U6427 (N_6427,N_5522,N_5955);
or U6428 (N_6428,N_5524,N_5665);
xor U6429 (N_6429,N_5570,N_5627);
nor U6430 (N_6430,N_5621,N_5728);
and U6431 (N_6431,N_5835,N_5744);
nor U6432 (N_6432,N_5588,N_5760);
and U6433 (N_6433,N_5960,N_5948);
nor U6434 (N_6434,N_5881,N_5573);
xor U6435 (N_6435,N_5778,N_5576);
and U6436 (N_6436,N_5653,N_5808);
or U6437 (N_6437,N_5577,N_5584);
or U6438 (N_6438,N_5649,N_5686);
and U6439 (N_6439,N_5749,N_5844);
nor U6440 (N_6440,N_5669,N_5883);
xor U6441 (N_6441,N_5812,N_5577);
xnor U6442 (N_6442,N_5797,N_5885);
xor U6443 (N_6443,N_5641,N_5729);
or U6444 (N_6444,N_5981,N_5554);
nand U6445 (N_6445,N_5830,N_5715);
and U6446 (N_6446,N_5765,N_5978);
xnor U6447 (N_6447,N_5619,N_5661);
nor U6448 (N_6448,N_5897,N_5757);
nand U6449 (N_6449,N_5522,N_5604);
nor U6450 (N_6450,N_5605,N_5732);
nand U6451 (N_6451,N_5579,N_5823);
nand U6452 (N_6452,N_5991,N_5938);
nor U6453 (N_6453,N_5691,N_5996);
xor U6454 (N_6454,N_5710,N_5970);
and U6455 (N_6455,N_5982,N_5601);
or U6456 (N_6456,N_5715,N_5891);
nor U6457 (N_6457,N_5939,N_5703);
nor U6458 (N_6458,N_5664,N_5665);
and U6459 (N_6459,N_5510,N_5827);
or U6460 (N_6460,N_5669,N_5728);
and U6461 (N_6461,N_5719,N_5509);
nand U6462 (N_6462,N_5643,N_5922);
and U6463 (N_6463,N_5862,N_5735);
nand U6464 (N_6464,N_5947,N_5523);
and U6465 (N_6465,N_5857,N_5897);
or U6466 (N_6466,N_5731,N_5533);
nand U6467 (N_6467,N_5544,N_5922);
nor U6468 (N_6468,N_5956,N_5963);
nand U6469 (N_6469,N_5662,N_5826);
xor U6470 (N_6470,N_5938,N_5545);
or U6471 (N_6471,N_5989,N_5622);
xnor U6472 (N_6472,N_5927,N_5674);
or U6473 (N_6473,N_5891,N_5853);
and U6474 (N_6474,N_5737,N_5543);
and U6475 (N_6475,N_5998,N_5506);
nor U6476 (N_6476,N_5504,N_5730);
and U6477 (N_6477,N_5510,N_5693);
or U6478 (N_6478,N_5546,N_5704);
nor U6479 (N_6479,N_5609,N_5986);
xor U6480 (N_6480,N_5839,N_5940);
and U6481 (N_6481,N_5616,N_5800);
or U6482 (N_6482,N_5871,N_5929);
and U6483 (N_6483,N_5785,N_5813);
and U6484 (N_6484,N_5994,N_5864);
xor U6485 (N_6485,N_5878,N_5874);
nor U6486 (N_6486,N_5854,N_5663);
nor U6487 (N_6487,N_5595,N_5978);
nor U6488 (N_6488,N_5524,N_5923);
or U6489 (N_6489,N_5887,N_5662);
xnor U6490 (N_6490,N_5777,N_5545);
or U6491 (N_6491,N_5998,N_5713);
xnor U6492 (N_6492,N_5512,N_5660);
nor U6493 (N_6493,N_5689,N_5917);
xor U6494 (N_6494,N_5540,N_5899);
and U6495 (N_6495,N_5755,N_5509);
and U6496 (N_6496,N_5955,N_5765);
nor U6497 (N_6497,N_5672,N_5997);
nand U6498 (N_6498,N_5905,N_5959);
or U6499 (N_6499,N_5520,N_5651);
and U6500 (N_6500,N_6051,N_6269);
or U6501 (N_6501,N_6274,N_6050);
nor U6502 (N_6502,N_6008,N_6130);
nand U6503 (N_6503,N_6141,N_6182);
xnor U6504 (N_6504,N_6053,N_6242);
and U6505 (N_6505,N_6097,N_6123);
and U6506 (N_6506,N_6469,N_6065);
xnor U6507 (N_6507,N_6232,N_6104);
nor U6508 (N_6508,N_6064,N_6186);
or U6509 (N_6509,N_6367,N_6244);
and U6510 (N_6510,N_6328,N_6144);
nand U6511 (N_6511,N_6233,N_6372);
nand U6512 (N_6512,N_6313,N_6149);
xor U6513 (N_6513,N_6259,N_6408);
nand U6514 (N_6514,N_6423,N_6380);
xor U6515 (N_6515,N_6049,N_6194);
xor U6516 (N_6516,N_6025,N_6337);
or U6517 (N_6517,N_6292,N_6207);
xnor U6518 (N_6518,N_6320,N_6377);
and U6519 (N_6519,N_6222,N_6121);
xor U6520 (N_6520,N_6155,N_6430);
or U6521 (N_6521,N_6005,N_6268);
and U6522 (N_6522,N_6083,N_6322);
or U6523 (N_6523,N_6001,N_6303);
xor U6524 (N_6524,N_6418,N_6312);
nor U6525 (N_6525,N_6206,N_6192);
nand U6526 (N_6526,N_6283,N_6470);
nand U6527 (N_6527,N_6093,N_6341);
xor U6528 (N_6528,N_6007,N_6483);
nor U6529 (N_6529,N_6250,N_6387);
nand U6530 (N_6530,N_6247,N_6090);
or U6531 (N_6531,N_6276,N_6358);
or U6532 (N_6532,N_6038,N_6397);
and U6533 (N_6533,N_6111,N_6286);
or U6534 (N_6534,N_6138,N_6249);
nor U6535 (N_6535,N_6096,N_6431);
and U6536 (N_6536,N_6238,N_6463);
nand U6537 (N_6537,N_6044,N_6391);
and U6538 (N_6538,N_6438,N_6285);
and U6539 (N_6539,N_6231,N_6190);
nor U6540 (N_6540,N_6376,N_6109);
and U6541 (N_6541,N_6160,N_6340);
nor U6542 (N_6542,N_6492,N_6355);
or U6543 (N_6543,N_6311,N_6471);
nor U6544 (N_6544,N_6494,N_6068);
xor U6545 (N_6545,N_6241,N_6421);
or U6546 (N_6546,N_6415,N_6026);
nand U6547 (N_6547,N_6239,N_6077);
and U6548 (N_6548,N_6115,N_6200);
nand U6549 (N_6549,N_6054,N_6331);
xnor U6550 (N_6550,N_6425,N_6344);
or U6551 (N_6551,N_6066,N_6323);
and U6552 (N_6552,N_6087,N_6099);
xnor U6553 (N_6553,N_6256,N_6079);
nand U6554 (N_6554,N_6092,N_6393);
nand U6555 (N_6555,N_6432,N_6378);
and U6556 (N_6556,N_6481,N_6027);
nand U6557 (N_6557,N_6370,N_6422);
or U6558 (N_6558,N_6437,N_6354);
nand U6559 (N_6559,N_6384,N_6227);
nor U6560 (N_6560,N_6347,N_6414);
xnor U6561 (N_6561,N_6113,N_6143);
or U6562 (N_6562,N_6265,N_6228);
nand U6563 (N_6563,N_6462,N_6018);
xnor U6564 (N_6564,N_6289,N_6124);
and U6565 (N_6565,N_6282,N_6279);
or U6566 (N_6566,N_6031,N_6270);
and U6567 (N_6567,N_6335,N_6224);
xor U6568 (N_6568,N_6448,N_6290);
and U6569 (N_6569,N_6450,N_6114);
and U6570 (N_6570,N_6205,N_6459);
nand U6571 (N_6571,N_6284,N_6366);
nand U6572 (N_6572,N_6125,N_6277);
or U6573 (N_6573,N_6017,N_6348);
nand U6574 (N_6574,N_6254,N_6101);
or U6575 (N_6575,N_6253,N_6310);
nand U6576 (N_6576,N_6363,N_6041);
nor U6577 (N_6577,N_6305,N_6489);
nand U6578 (N_6578,N_6266,N_6142);
and U6579 (N_6579,N_6103,N_6166);
xnor U6580 (N_6580,N_6074,N_6364);
or U6581 (N_6581,N_6082,N_6009);
xnor U6582 (N_6582,N_6043,N_6412);
nor U6583 (N_6583,N_6139,N_6336);
nor U6584 (N_6584,N_6003,N_6442);
nor U6585 (N_6585,N_6497,N_6296);
nand U6586 (N_6586,N_6201,N_6407);
nor U6587 (N_6587,N_6126,N_6246);
nor U6588 (N_6588,N_6342,N_6309);
or U6589 (N_6589,N_6151,N_6162);
xor U6590 (N_6590,N_6168,N_6332);
nor U6591 (N_6591,N_6175,N_6440);
nand U6592 (N_6592,N_6482,N_6374);
nor U6593 (N_6593,N_6157,N_6167);
nand U6594 (N_6594,N_6444,N_6002);
and U6595 (N_6595,N_6080,N_6076);
and U6596 (N_6596,N_6356,N_6392);
nor U6597 (N_6597,N_6446,N_6346);
or U6598 (N_6598,N_6004,N_6496);
and U6599 (N_6599,N_6034,N_6449);
and U6600 (N_6600,N_6088,N_6251);
nor U6601 (N_6601,N_6291,N_6174);
xor U6602 (N_6602,N_6181,N_6488);
xnor U6603 (N_6603,N_6381,N_6278);
xor U6604 (N_6604,N_6189,N_6297);
and U6605 (N_6605,N_6248,N_6135);
xnor U6606 (N_6606,N_6120,N_6447);
or U6607 (N_6607,N_6402,N_6211);
and U6608 (N_6608,N_6011,N_6304);
nand U6609 (N_6609,N_6028,N_6406);
nor U6610 (N_6610,N_6413,N_6287);
and U6611 (N_6611,N_6330,N_6257);
xor U6612 (N_6612,N_6013,N_6486);
xor U6613 (N_6613,N_6016,N_6417);
or U6614 (N_6614,N_6161,N_6229);
or U6615 (N_6615,N_6495,N_6436);
nand U6616 (N_6616,N_6301,N_6019);
and U6617 (N_6617,N_6493,N_6209);
xor U6618 (N_6618,N_6416,N_6293);
or U6619 (N_6619,N_6199,N_6343);
nand U6620 (N_6620,N_6014,N_6140);
xor U6621 (N_6621,N_6389,N_6221);
and U6622 (N_6622,N_6171,N_6237);
nand U6623 (N_6623,N_6198,N_6318);
nand U6624 (N_6624,N_6261,N_6006);
nand U6625 (N_6625,N_6308,N_6036);
xor U6626 (N_6626,N_6275,N_6294);
or U6627 (N_6627,N_6410,N_6477);
and U6628 (N_6628,N_6345,N_6434);
nor U6629 (N_6629,N_6105,N_6267);
nor U6630 (N_6630,N_6152,N_6165);
nor U6631 (N_6631,N_6339,N_6073);
xnor U6632 (N_6632,N_6252,N_6122);
nand U6633 (N_6633,N_6445,N_6490);
and U6634 (N_6634,N_6298,N_6060);
and U6635 (N_6635,N_6403,N_6146);
and U6636 (N_6636,N_6116,N_6176);
nor U6637 (N_6637,N_6147,N_6000);
xnor U6638 (N_6638,N_6480,N_6401);
or U6639 (N_6639,N_6321,N_6169);
xnor U6640 (N_6640,N_6178,N_6362);
nor U6641 (N_6641,N_6095,N_6338);
and U6642 (N_6642,N_6258,N_6193);
nor U6643 (N_6643,N_6315,N_6295);
and U6644 (N_6644,N_6170,N_6020);
nor U6645 (N_6645,N_6173,N_6390);
xor U6646 (N_6646,N_6059,N_6230);
nor U6647 (N_6647,N_6235,N_6150);
and U6648 (N_6648,N_6187,N_6210);
or U6649 (N_6649,N_6204,N_6273);
or U6650 (N_6650,N_6317,N_6188);
and U6651 (N_6651,N_6063,N_6131);
and U6652 (N_6652,N_6196,N_6365);
nand U6653 (N_6653,N_6467,N_6386);
and U6654 (N_6654,N_6236,N_6314);
nor U6655 (N_6655,N_6262,N_6098);
nor U6656 (N_6656,N_6375,N_6089);
or U6657 (N_6657,N_6172,N_6263);
nand U6658 (N_6658,N_6214,N_6491);
xor U6659 (N_6659,N_6145,N_6443);
or U6660 (N_6660,N_6136,N_6465);
and U6661 (N_6661,N_6218,N_6404);
nand U6662 (N_6662,N_6156,N_6048);
nor U6663 (N_6663,N_6225,N_6455);
or U6664 (N_6664,N_6302,N_6349);
and U6665 (N_6665,N_6454,N_6466);
nand U6666 (N_6666,N_6361,N_6106);
nor U6667 (N_6667,N_6394,N_6243);
xor U6668 (N_6668,N_6484,N_6058);
nand U6669 (N_6669,N_6351,N_6091);
nor U6670 (N_6670,N_6102,N_6062);
xor U6671 (N_6671,N_6220,N_6042);
xnor U6672 (N_6672,N_6353,N_6326);
nor U6673 (N_6673,N_6129,N_6396);
nand U6674 (N_6674,N_6385,N_6153);
xor U6675 (N_6675,N_6215,N_6468);
nor U6676 (N_6676,N_6179,N_6395);
nand U6677 (N_6677,N_6281,N_6216);
xnor U6678 (N_6678,N_6306,N_6219);
xor U6679 (N_6679,N_6071,N_6067);
nor U6680 (N_6680,N_6280,N_6223);
nor U6681 (N_6681,N_6100,N_6226);
and U6682 (N_6682,N_6327,N_6324);
nor U6683 (N_6683,N_6400,N_6203);
and U6684 (N_6684,N_6388,N_6056);
and U6685 (N_6685,N_6420,N_6197);
or U6686 (N_6686,N_6158,N_6072);
xnor U6687 (N_6687,N_6030,N_6163);
and U6688 (N_6688,N_6118,N_6154);
nand U6689 (N_6689,N_6010,N_6319);
or U6690 (N_6690,N_6498,N_6107);
and U6691 (N_6691,N_6035,N_6360);
or U6692 (N_6692,N_6428,N_6047);
nor U6693 (N_6693,N_6399,N_6382);
xor U6694 (N_6694,N_6039,N_6405);
nand U6695 (N_6695,N_6180,N_6451);
or U6696 (N_6696,N_6078,N_6456);
or U6697 (N_6697,N_6127,N_6055);
xor U6698 (N_6698,N_6255,N_6046);
or U6699 (N_6699,N_6094,N_6022);
nor U6700 (N_6700,N_6184,N_6373);
nor U6701 (N_6701,N_6137,N_6021);
nand U6702 (N_6702,N_6134,N_6040);
or U6703 (N_6703,N_6473,N_6409);
or U6704 (N_6704,N_6457,N_6108);
and U6705 (N_6705,N_6128,N_6212);
and U6706 (N_6706,N_6119,N_6075);
xnor U6707 (N_6707,N_6368,N_6427);
nand U6708 (N_6708,N_6217,N_6369);
nor U6709 (N_6709,N_6350,N_6271);
or U6710 (N_6710,N_6429,N_6177);
and U6711 (N_6711,N_6419,N_6029);
nor U6712 (N_6712,N_6478,N_6245);
and U6713 (N_6713,N_6061,N_6359);
nand U6714 (N_6714,N_6475,N_6299);
nor U6715 (N_6715,N_6325,N_6133);
nand U6716 (N_6716,N_6479,N_6272);
and U6717 (N_6717,N_6015,N_6460);
xnor U6718 (N_6718,N_6045,N_6458);
and U6719 (N_6719,N_6260,N_6439);
nor U6720 (N_6720,N_6398,N_6300);
nand U6721 (N_6721,N_6112,N_6464);
xor U6722 (N_6722,N_6316,N_6307);
and U6723 (N_6723,N_6461,N_6452);
and U6724 (N_6724,N_6499,N_6012);
nor U6725 (N_6725,N_6069,N_6476);
nand U6726 (N_6726,N_6033,N_6333);
nand U6727 (N_6727,N_6084,N_6191);
nand U6728 (N_6728,N_6487,N_6213);
or U6729 (N_6729,N_6234,N_6183);
or U6730 (N_6730,N_6159,N_6023);
xnor U6731 (N_6731,N_6195,N_6383);
nand U6732 (N_6732,N_6329,N_6379);
or U6733 (N_6733,N_6357,N_6202);
nor U6734 (N_6734,N_6164,N_6024);
nor U6735 (N_6735,N_6264,N_6110);
or U6736 (N_6736,N_6352,N_6441);
nor U6737 (N_6737,N_6148,N_6070);
nand U6738 (N_6738,N_6208,N_6334);
xor U6739 (N_6739,N_6426,N_6433);
nor U6740 (N_6740,N_6132,N_6474);
xor U6741 (N_6741,N_6032,N_6424);
nor U6742 (N_6742,N_6086,N_6052);
xor U6743 (N_6743,N_6085,N_6057);
nand U6744 (N_6744,N_6411,N_6117);
xor U6745 (N_6745,N_6435,N_6081);
xnor U6746 (N_6746,N_6472,N_6485);
or U6747 (N_6747,N_6288,N_6371);
and U6748 (N_6748,N_6185,N_6453);
and U6749 (N_6749,N_6037,N_6240);
nor U6750 (N_6750,N_6094,N_6268);
xor U6751 (N_6751,N_6143,N_6345);
or U6752 (N_6752,N_6005,N_6076);
nand U6753 (N_6753,N_6288,N_6216);
nand U6754 (N_6754,N_6136,N_6354);
and U6755 (N_6755,N_6084,N_6291);
xnor U6756 (N_6756,N_6378,N_6347);
nor U6757 (N_6757,N_6459,N_6361);
nand U6758 (N_6758,N_6189,N_6427);
or U6759 (N_6759,N_6055,N_6311);
and U6760 (N_6760,N_6079,N_6092);
nor U6761 (N_6761,N_6004,N_6242);
nor U6762 (N_6762,N_6341,N_6103);
nor U6763 (N_6763,N_6496,N_6283);
nand U6764 (N_6764,N_6245,N_6178);
and U6765 (N_6765,N_6135,N_6260);
or U6766 (N_6766,N_6355,N_6182);
xnor U6767 (N_6767,N_6040,N_6156);
xnor U6768 (N_6768,N_6132,N_6407);
nand U6769 (N_6769,N_6114,N_6481);
xor U6770 (N_6770,N_6229,N_6196);
and U6771 (N_6771,N_6308,N_6206);
nand U6772 (N_6772,N_6027,N_6018);
or U6773 (N_6773,N_6095,N_6140);
nand U6774 (N_6774,N_6071,N_6370);
nor U6775 (N_6775,N_6213,N_6003);
nor U6776 (N_6776,N_6434,N_6374);
or U6777 (N_6777,N_6473,N_6484);
nand U6778 (N_6778,N_6482,N_6303);
nand U6779 (N_6779,N_6306,N_6468);
and U6780 (N_6780,N_6417,N_6179);
nand U6781 (N_6781,N_6238,N_6455);
or U6782 (N_6782,N_6357,N_6275);
or U6783 (N_6783,N_6452,N_6327);
nor U6784 (N_6784,N_6038,N_6146);
nor U6785 (N_6785,N_6295,N_6201);
nor U6786 (N_6786,N_6286,N_6146);
xor U6787 (N_6787,N_6292,N_6199);
and U6788 (N_6788,N_6268,N_6259);
xor U6789 (N_6789,N_6008,N_6090);
and U6790 (N_6790,N_6254,N_6463);
nor U6791 (N_6791,N_6279,N_6423);
or U6792 (N_6792,N_6342,N_6181);
nand U6793 (N_6793,N_6461,N_6146);
nor U6794 (N_6794,N_6110,N_6309);
nor U6795 (N_6795,N_6079,N_6189);
nor U6796 (N_6796,N_6352,N_6329);
and U6797 (N_6797,N_6056,N_6146);
and U6798 (N_6798,N_6446,N_6359);
nand U6799 (N_6799,N_6063,N_6186);
or U6800 (N_6800,N_6454,N_6323);
and U6801 (N_6801,N_6199,N_6470);
nor U6802 (N_6802,N_6301,N_6015);
nor U6803 (N_6803,N_6204,N_6005);
xnor U6804 (N_6804,N_6373,N_6347);
or U6805 (N_6805,N_6068,N_6359);
xor U6806 (N_6806,N_6138,N_6352);
or U6807 (N_6807,N_6017,N_6402);
or U6808 (N_6808,N_6030,N_6089);
or U6809 (N_6809,N_6172,N_6484);
nor U6810 (N_6810,N_6008,N_6248);
nand U6811 (N_6811,N_6022,N_6130);
or U6812 (N_6812,N_6284,N_6470);
or U6813 (N_6813,N_6144,N_6057);
xnor U6814 (N_6814,N_6094,N_6462);
or U6815 (N_6815,N_6247,N_6398);
nor U6816 (N_6816,N_6273,N_6339);
nor U6817 (N_6817,N_6217,N_6387);
xnor U6818 (N_6818,N_6180,N_6256);
nor U6819 (N_6819,N_6052,N_6072);
xnor U6820 (N_6820,N_6021,N_6306);
nor U6821 (N_6821,N_6270,N_6126);
nand U6822 (N_6822,N_6193,N_6050);
xnor U6823 (N_6823,N_6305,N_6391);
or U6824 (N_6824,N_6409,N_6221);
nor U6825 (N_6825,N_6139,N_6112);
nand U6826 (N_6826,N_6296,N_6302);
xor U6827 (N_6827,N_6213,N_6132);
or U6828 (N_6828,N_6287,N_6383);
nor U6829 (N_6829,N_6353,N_6105);
nor U6830 (N_6830,N_6031,N_6355);
and U6831 (N_6831,N_6419,N_6027);
nand U6832 (N_6832,N_6084,N_6391);
nor U6833 (N_6833,N_6434,N_6158);
nand U6834 (N_6834,N_6406,N_6096);
xnor U6835 (N_6835,N_6233,N_6451);
or U6836 (N_6836,N_6480,N_6077);
and U6837 (N_6837,N_6384,N_6038);
nor U6838 (N_6838,N_6344,N_6113);
xnor U6839 (N_6839,N_6472,N_6052);
and U6840 (N_6840,N_6407,N_6408);
or U6841 (N_6841,N_6403,N_6231);
or U6842 (N_6842,N_6412,N_6377);
xor U6843 (N_6843,N_6059,N_6225);
or U6844 (N_6844,N_6136,N_6303);
nor U6845 (N_6845,N_6388,N_6486);
nand U6846 (N_6846,N_6445,N_6469);
xnor U6847 (N_6847,N_6453,N_6486);
nand U6848 (N_6848,N_6168,N_6041);
nor U6849 (N_6849,N_6405,N_6148);
xnor U6850 (N_6850,N_6185,N_6458);
nand U6851 (N_6851,N_6135,N_6207);
and U6852 (N_6852,N_6168,N_6211);
and U6853 (N_6853,N_6152,N_6369);
or U6854 (N_6854,N_6057,N_6293);
nor U6855 (N_6855,N_6023,N_6421);
xor U6856 (N_6856,N_6390,N_6425);
nand U6857 (N_6857,N_6209,N_6167);
nor U6858 (N_6858,N_6460,N_6268);
and U6859 (N_6859,N_6246,N_6356);
xnor U6860 (N_6860,N_6188,N_6112);
xnor U6861 (N_6861,N_6467,N_6488);
xnor U6862 (N_6862,N_6118,N_6205);
and U6863 (N_6863,N_6051,N_6207);
or U6864 (N_6864,N_6449,N_6129);
nand U6865 (N_6865,N_6040,N_6305);
nand U6866 (N_6866,N_6356,N_6132);
and U6867 (N_6867,N_6332,N_6262);
nand U6868 (N_6868,N_6457,N_6237);
nand U6869 (N_6869,N_6411,N_6034);
nor U6870 (N_6870,N_6361,N_6453);
nand U6871 (N_6871,N_6109,N_6067);
nor U6872 (N_6872,N_6420,N_6005);
and U6873 (N_6873,N_6238,N_6488);
xor U6874 (N_6874,N_6462,N_6371);
or U6875 (N_6875,N_6072,N_6177);
xnor U6876 (N_6876,N_6297,N_6214);
xor U6877 (N_6877,N_6076,N_6471);
and U6878 (N_6878,N_6397,N_6279);
nand U6879 (N_6879,N_6303,N_6313);
nand U6880 (N_6880,N_6454,N_6441);
nand U6881 (N_6881,N_6344,N_6343);
or U6882 (N_6882,N_6194,N_6242);
nor U6883 (N_6883,N_6464,N_6137);
and U6884 (N_6884,N_6319,N_6288);
nor U6885 (N_6885,N_6087,N_6241);
or U6886 (N_6886,N_6155,N_6311);
or U6887 (N_6887,N_6210,N_6167);
xnor U6888 (N_6888,N_6208,N_6402);
and U6889 (N_6889,N_6421,N_6043);
or U6890 (N_6890,N_6339,N_6214);
xor U6891 (N_6891,N_6136,N_6225);
or U6892 (N_6892,N_6138,N_6121);
or U6893 (N_6893,N_6304,N_6271);
nand U6894 (N_6894,N_6248,N_6072);
nand U6895 (N_6895,N_6132,N_6263);
xnor U6896 (N_6896,N_6435,N_6138);
or U6897 (N_6897,N_6156,N_6467);
nand U6898 (N_6898,N_6258,N_6248);
and U6899 (N_6899,N_6088,N_6271);
and U6900 (N_6900,N_6147,N_6447);
nand U6901 (N_6901,N_6260,N_6275);
nor U6902 (N_6902,N_6181,N_6199);
xor U6903 (N_6903,N_6296,N_6471);
nor U6904 (N_6904,N_6137,N_6120);
or U6905 (N_6905,N_6413,N_6097);
or U6906 (N_6906,N_6283,N_6197);
xor U6907 (N_6907,N_6163,N_6406);
or U6908 (N_6908,N_6086,N_6031);
nand U6909 (N_6909,N_6448,N_6015);
xor U6910 (N_6910,N_6243,N_6166);
xor U6911 (N_6911,N_6134,N_6299);
nand U6912 (N_6912,N_6478,N_6399);
xnor U6913 (N_6913,N_6019,N_6294);
nand U6914 (N_6914,N_6124,N_6103);
xor U6915 (N_6915,N_6342,N_6453);
nor U6916 (N_6916,N_6414,N_6166);
xor U6917 (N_6917,N_6245,N_6405);
nand U6918 (N_6918,N_6467,N_6335);
nand U6919 (N_6919,N_6039,N_6021);
nor U6920 (N_6920,N_6442,N_6248);
nor U6921 (N_6921,N_6026,N_6323);
xor U6922 (N_6922,N_6026,N_6206);
or U6923 (N_6923,N_6405,N_6308);
nand U6924 (N_6924,N_6310,N_6362);
or U6925 (N_6925,N_6427,N_6311);
nor U6926 (N_6926,N_6296,N_6210);
or U6927 (N_6927,N_6220,N_6108);
nor U6928 (N_6928,N_6151,N_6197);
nor U6929 (N_6929,N_6425,N_6000);
nand U6930 (N_6930,N_6091,N_6159);
and U6931 (N_6931,N_6409,N_6035);
nor U6932 (N_6932,N_6250,N_6367);
nor U6933 (N_6933,N_6337,N_6017);
xnor U6934 (N_6934,N_6198,N_6270);
nor U6935 (N_6935,N_6084,N_6277);
nand U6936 (N_6936,N_6116,N_6225);
nor U6937 (N_6937,N_6010,N_6463);
and U6938 (N_6938,N_6450,N_6072);
and U6939 (N_6939,N_6074,N_6439);
nand U6940 (N_6940,N_6024,N_6109);
nor U6941 (N_6941,N_6466,N_6115);
xnor U6942 (N_6942,N_6131,N_6380);
nand U6943 (N_6943,N_6025,N_6332);
or U6944 (N_6944,N_6405,N_6201);
nor U6945 (N_6945,N_6104,N_6170);
nor U6946 (N_6946,N_6176,N_6052);
nor U6947 (N_6947,N_6056,N_6218);
nor U6948 (N_6948,N_6259,N_6266);
xnor U6949 (N_6949,N_6057,N_6401);
nor U6950 (N_6950,N_6069,N_6028);
or U6951 (N_6951,N_6483,N_6260);
nor U6952 (N_6952,N_6052,N_6006);
nand U6953 (N_6953,N_6223,N_6048);
and U6954 (N_6954,N_6151,N_6057);
nand U6955 (N_6955,N_6448,N_6264);
or U6956 (N_6956,N_6490,N_6422);
xor U6957 (N_6957,N_6303,N_6416);
nand U6958 (N_6958,N_6299,N_6235);
nand U6959 (N_6959,N_6052,N_6361);
or U6960 (N_6960,N_6472,N_6131);
nand U6961 (N_6961,N_6238,N_6487);
nand U6962 (N_6962,N_6295,N_6318);
nor U6963 (N_6963,N_6360,N_6298);
and U6964 (N_6964,N_6260,N_6385);
nand U6965 (N_6965,N_6394,N_6228);
nand U6966 (N_6966,N_6480,N_6249);
nand U6967 (N_6967,N_6475,N_6241);
or U6968 (N_6968,N_6017,N_6291);
xor U6969 (N_6969,N_6319,N_6116);
and U6970 (N_6970,N_6361,N_6437);
xor U6971 (N_6971,N_6261,N_6463);
nand U6972 (N_6972,N_6140,N_6407);
nand U6973 (N_6973,N_6303,N_6369);
xnor U6974 (N_6974,N_6206,N_6369);
or U6975 (N_6975,N_6335,N_6244);
xnor U6976 (N_6976,N_6251,N_6358);
and U6977 (N_6977,N_6331,N_6198);
or U6978 (N_6978,N_6286,N_6302);
nor U6979 (N_6979,N_6072,N_6304);
or U6980 (N_6980,N_6242,N_6477);
nor U6981 (N_6981,N_6110,N_6340);
or U6982 (N_6982,N_6432,N_6223);
and U6983 (N_6983,N_6310,N_6316);
and U6984 (N_6984,N_6263,N_6214);
nand U6985 (N_6985,N_6233,N_6073);
xnor U6986 (N_6986,N_6344,N_6463);
nor U6987 (N_6987,N_6105,N_6047);
or U6988 (N_6988,N_6011,N_6381);
or U6989 (N_6989,N_6494,N_6251);
or U6990 (N_6990,N_6437,N_6443);
or U6991 (N_6991,N_6253,N_6364);
nand U6992 (N_6992,N_6412,N_6367);
nand U6993 (N_6993,N_6140,N_6152);
and U6994 (N_6994,N_6250,N_6203);
or U6995 (N_6995,N_6243,N_6175);
xor U6996 (N_6996,N_6380,N_6369);
xor U6997 (N_6997,N_6401,N_6335);
and U6998 (N_6998,N_6485,N_6287);
and U6999 (N_6999,N_6388,N_6395);
nand U7000 (N_7000,N_6845,N_6704);
nor U7001 (N_7001,N_6767,N_6913);
nand U7002 (N_7002,N_6677,N_6896);
xnor U7003 (N_7003,N_6951,N_6539);
or U7004 (N_7004,N_6738,N_6734);
xnor U7005 (N_7005,N_6865,N_6795);
xor U7006 (N_7006,N_6668,N_6524);
nor U7007 (N_7007,N_6639,N_6712);
nand U7008 (N_7008,N_6983,N_6915);
and U7009 (N_7009,N_6556,N_6519);
xor U7010 (N_7010,N_6981,N_6755);
nor U7011 (N_7011,N_6581,N_6813);
nand U7012 (N_7012,N_6529,N_6846);
nor U7013 (N_7013,N_6544,N_6957);
and U7014 (N_7014,N_6949,N_6579);
nand U7015 (N_7015,N_6572,N_6779);
nand U7016 (N_7016,N_6920,N_6891);
and U7017 (N_7017,N_6757,N_6526);
nand U7018 (N_7018,N_6614,N_6771);
or U7019 (N_7019,N_6561,N_6597);
nor U7020 (N_7020,N_6724,N_6793);
nor U7021 (N_7021,N_6853,N_6875);
and U7022 (N_7022,N_6855,N_6772);
nand U7023 (N_7023,N_6617,N_6815);
xor U7024 (N_7024,N_6641,N_6858);
or U7025 (N_7025,N_6825,N_6551);
and U7026 (N_7026,N_6821,N_6986);
or U7027 (N_7027,N_6722,N_6732);
or U7028 (N_7028,N_6792,N_6765);
or U7029 (N_7029,N_6691,N_6850);
nand U7030 (N_7030,N_6895,N_6522);
or U7031 (N_7031,N_6726,N_6884);
nand U7032 (N_7032,N_6684,N_6801);
or U7033 (N_7033,N_6616,N_6747);
nand U7034 (N_7034,N_6952,N_6856);
or U7035 (N_7035,N_6973,N_6511);
xnor U7036 (N_7036,N_6545,N_6903);
xnor U7037 (N_7037,N_6535,N_6809);
nor U7038 (N_7038,N_6723,N_6701);
and U7039 (N_7039,N_6532,N_6506);
or U7040 (N_7040,N_6642,N_6688);
nor U7041 (N_7041,N_6708,N_6868);
and U7042 (N_7042,N_6750,N_6509);
and U7043 (N_7043,N_6596,N_6580);
and U7044 (N_7044,N_6512,N_6749);
nand U7045 (N_7045,N_6721,N_6907);
and U7046 (N_7046,N_6810,N_6824);
and U7047 (N_7047,N_6897,N_6840);
xnor U7048 (N_7048,N_6626,N_6842);
nor U7049 (N_7049,N_6553,N_6823);
nand U7050 (N_7050,N_6909,N_6656);
nand U7051 (N_7051,N_6740,N_6817);
or U7052 (N_7052,N_6621,N_6925);
or U7053 (N_7053,N_6820,N_6569);
or U7054 (N_7054,N_6518,N_6733);
and U7055 (N_7055,N_6504,N_6816);
nand U7056 (N_7056,N_6961,N_6864);
nor U7057 (N_7057,N_6716,N_6727);
and U7058 (N_7058,N_6784,N_6670);
xor U7059 (N_7059,N_6835,N_6690);
xnor U7060 (N_7060,N_6568,N_6660);
nand U7061 (N_7061,N_6782,N_6759);
xnor U7062 (N_7062,N_6559,N_6904);
xnor U7063 (N_7063,N_6631,N_6698);
or U7064 (N_7064,N_6836,N_6542);
nor U7065 (N_7065,N_6586,N_6911);
or U7066 (N_7066,N_6847,N_6681);
or U7067 (N_7067,N_6968,N_6826);
and U7068 (N_7068,N_6959,N_6988);
xnor U7069 (N_7069,N_6797,N_6878);
or U7070 (N_7070,N_6989,N_6618);
xor U7071 (N_7071,N_6935,N_6877);
nand U7072 (N_7072,N_6623,N_6540);
nand U7073 (N_7073,N_6859,N_6997);
nor U7074 (N_7074,N_6994,N_6502);
and U7075 (N_7075,N_6743,N_6564);
or U7076 (N_7076,N_6565,N_6972);
nor U7077 (N_7077,N_6598,N_6888);
xnor U7078 (N_7078,N_6803,N_6978);
and U7079 (N_7079,N_6653,N_6683);
nand U7080 (N_7080,N_6508,N_6971);
and U7081 (N_7081,N_6881,N_6744);
or U7082 (N_7082,N_6672,N_6876);
nor U7083 (N_7083,N_6692,N_6657);
nor U7084 (N_7084,N_6894,N_6600);
nor U7085 (N_7085,N_6916,N_6886);
and U7086 (N_7086,N_6520,N_6808);
nand U7087 (N_7087,N_6606,N_6848);
or U7088 (N_7088,N_6742,N_6887);
or U7089 (N_7089,N_6662,N_6863);
nand U7090 (N_7090,N_6777,N_6576);
nand U7091 (N_7091,N_6831,N_6599);
nand U7092 (N_7092,N_6638,N_6584);
nor U7093 (N_7093,N_6912,N_6667);
nor U7094 (N_7094,N_6676,N_6958);
nand U7095 (N_7095,N_6892,N_6788);
and U7096 (N_7096,N_6900,N_6658);
or U7097 (N_7097,N_6607,N_6866);
or U7098 (N_7098,N_6622,N_6562);
and U7099 (N_7099,N_6729,N_6645);
xnor U7100 (N_7100,N_6785,N_6929);
and U7101 (N_7101,N_6828,N_6554);
nand U7102 (N_7102,N_6939,N_6787);
nor U7103 (N_7103,N_6905,N_6937);
xnor U7104 (N_7104,N_6583,N_6770);
and U7105 (N_7105,N_6790,N_6609);
nand U7106 (N_7106,N_6711,N_6654);
or U7107 (N_7107,N_6985,N_6830);
nor U7108 (N_7108,N_6906,N_6893);
nor U7109 (N_7109,N_6902,N_6608);
or U7110 (N_7110,N_6928,N_6758);
xnor U7111 (N_7111,N_6873,N_6604);
nand U7112 (N_7112,N_6574,N_6625);
and U7113 (N_7113,N_6687,N_6955);
or U7114 (N_7114,N_6773,N_6992);
and U7115 (N_7115,N_6976,N_6548);
nor U7116 (N_7116,N_6694,N_6812);
and U7117 (N_7117,N_6999,N_6860);
nand U7118 (N_7118,N_6550,N_6696);
xnor U7119 (N_7119,N_6500,N_6965);
and U7120 (N_7120,N_6854,N_6523);
nor U7121 (N_7121,N_6590,N_6947);
nand U7122 (N_7122,N_6567,N_6807);
or U7123 (N_7123,N_6970,N_6924);
xnor U7124 (N_7124,N_6932,N_6753);
and U7125 (N_7125,N_6852,N_6635);
nor U7126 (N_7126,N_6751,N_6980);
xor U7127 (N_7127,N_6543,N_6769);
nand U7128 (N_7128,N_6552,N_6710);
or U7129 (N_7129,N_6977,N_6630);
xnor U7130 (N_7130,N_6686,N_6882);
nand U7131 (N_7131,N_6774,N_6620);
nor U7132 (N_7132,N_6998,N_6762);
xnor U7133 (N_7133,N_6885,N_6501);
nor U7134 (N_7134,N_6601,N_6814);
and U7135 (N_7135,N_6967,N_6781);
nand U7136 (N_7136,N_6778,N_6528);
or U7137 (N_7137,N_6592,N_6637);
nand U7138 (N_7138,N_6533,N_6948);
or U7139 (N_7139,N_6923,N_6697);
nand U7140 (N_7140,N_6546,N_6934);
nor U7141 (N_7141,N_6640,N_6754);
nor U7142 (N_7142,N_6731,N_6883);
nor U7143 (N_7143,N_6615,N_6619);
nor U7144 (N_7144,N_6736,N_6776);
and U7145 (N_7145,N_6841,N_6521);
nand U7146 (N_7146,N_6987,N_6602);
xnor U7147 (N_7147,N_6818,N_6730);
and U7148 (N_7148,N_6946,N_6570);
and U7149 (N_7149,N_6950,N_6857);
xnor U7150 (N_7150,N_6990,N_6764);
nor U7151 (N_7151,N_6761,N_6833);
nand U7152 (N_7152,N_6557,N_6707);
nand U7153 (N_7153,N_6647,N_6588);
or U7154 (N_7154,N_6666,N_6555);
and U7155 (N_7155,N_6851,N_6627);
nand U7156 (N_7156,N_6665,N_6589);
nand U7157 (N_7157,N_6943,N_6699);
nand U7158 (N_7158,N_6908,N_6664);
xnor U7159 (N_7159,N_6862,N_6735);
or U7160 (N_7160,N_6984,N_6838);
or U7161 (N_7161,N_6587,N_6563);
and U7162 (N_7162,N_6930,N_6582);
nor U7163 (N_7163,N_6652,N_6964);
or U7164 (N_7164,N_6700,N_6629);
xnor U7165 (N_7165,N_6940,N_6786);
and U7166 (N_7166,N_6648,N_6577);
xor U7167 (N_7167,N_6944,N_6603);
xor U7168 (N_7168,N_6613,N_6612);
nand U7169 (N_7169,N_6991,N_6796);
or U7170 (N_7170,N_6673,N_6513);
nor U7171 (N_7171,N_6760,N_6956);
and U7172 (N_7172,N_6671,N_6936);
xor U7173 (N_7173,N_6960,N_6517);
xnor U7174 (N_7174,N_6921,N_6610);
nor U7175 (N_7175,N_6679,N_6982);
and U7176 (N_7176,N_6611,N_6516);
nand U7177 (N_7177,N_6541,N_6922);
or U7178 (N_7178,N_6595,N_6822);
nand U7179 (N_7179,N_6689,N_6725);
xor U7180 (N_7180,N_6644,N_6867);
nand U7181 (N_7181,N_6558,N_6593);
or U7182 (N_7182,N_6507,N_6879);
or U7183 (N_7183,N_6632,N_6942);
and U7184 (N_7184,N_6663,N_6996);
nor U7185 (N_7185,N_6746,N_6702);
nand U7186 (N_7186,N_6514,N_6919);
nand U7187 (N_7187,N_6861,N_6962);
or U7188 (N_7188,N_6804,N_6931);
or U7189 (N_7189,N_6674,N_6693);
or U7190 (N_7190,N_6872,N_6870);
and U7191 (N_7191,N_6536,N_6655);
nand U7192 (N_7192,N_6510,N_6910);
nor U7193 (N_7193,N_6926,N_6719);
nor U7194 (N_7194,N_6800,N_6953);
nand U7195 (N_7195,N_6829,N_6703);
nor U7196 (N_7196,N_6917,N_6874);
and U7197 (N_7197,N_6775,N_6525);
or U7198 (N_7198,N_6680,N_6537);
xor U7199 (N_7199,N_6748,N_6571);
or U7200 (N_7200,N_6649,N_6752);
nor U7201 (N_7201,N_6993,N_6651);
nand U7202 (N_7202,N_6954,N_6745);
xor U7203 (N_7203,N_6505,N_6695);
nor U7204 (N_7204,N_6871,N_6768);
and U7205 (N_7205,N_6901,N_6578);
xor U7206 (N_7206,N_6780,N_6685);
nand U7207 (N_7207,N_6643,N_6975);
nand U7208 (N_7208,N_6789,N_6869);
nor U7209 (N_7209,N_6628,N_6566);
xor U7210 (N_7210,N_6933,N_6794);
or U7211 (N_7211,N_6624,N_6515);
and U7212 (N_7212,N_6591,N_6979);
and U7213 (N_7213,N_6718,N_6669);
or U7214 (N_7214,N_6927,N_6941);
and U7215 (N_7215,N_6741,N_6791);
xor U7216 (N_7216,N_6898,N_6739);
nor U7217 (N_7217,N_6560,N_6715);
or U7218 (N_7218,N_6633,N_6661);
or U7219 (N_7219,N_6918,N_6575);
nor U7220 (N_7220,N_6995,N_6547);
nor U7221 (N_7221,N_6811,N_6837);
nor U7222 (N_7222,N_6880,N_6705);
and U7223 (N_7223,N_6714,N_6527);
nand U7224 (N_7224,N_6538,N_6717);
or U7225 (N_7225,N_6675,N_6737);
xnor U7226 (N_7226,N_6573,N_6728);
or U7227 (N_7227,N_6849,N_6819);
nand U7228 (N_7228,N_6963,N_6890);
nor U7229 (N_7229,N_6720,N_6969);
xnor U7230 (N_7230,N_6914,N_6889);
xnor U7231 (N_7231,N_6605,N_6938);
nand U7232 (N_7232,N_6594,N_6636);
or U7233 (N_7233,N_6678,N_6799);
nand U7234 (N_7234,N_6798,N_6709);
nand U7235 (N_7235,N_6530,N_6549);
or U7236 (N_7236,N_6706,N_6805);
xnor U7237 (N_7237,N_6650,N_6844);
xnor U7238 (N_7238,N_6839,N_6899);
nor U7239 (N_7239,N_6783,N_6974);
and U7240 (N_7240,N_6682,N_6834);
nand U7241 (N_7241,N_6531,N_6646);
or U7242 (N_7242,N_6832,N_6802);
and U7243 (N_7243,N_6945,N_6966);
and U7244 (N_7244,N_6766,N_6503);
nand U7245 (N_7245,N_6756,N_6534);
nor U7246 (N_7246,N_6806,N_6843);
nor U7247 (N_7247,N_6827,N_6634);
xor U7248 (N_7248,N_6763,N_6713);
nor U7249 (N_7249,N_6585,N_6659);
nand U7250 (N_7250,N_6914,N_6844);
and U7251 (N_7251,N_6508,N_6776);
or U7252 (N_7252,N_6753,N_6935);
nor U7253 (N_7253,N_6647,N_6689);
nor U7254 (N_7254,N_6681,N_6530);
nand U7255 (N_7255,N_6927,N_6682);
nor U7256 (N_7256,N_6831,N_6683);
xnor U7257 (N_7257,N_6670,N_6964);
nand U7258 (N_7258,N_6735,N_6613);
xor U7259 (N_7259,N_6796,N_6815);
or U7260 (N_7260,N_6663,N_6501);
nor U7261 (N_7261,N_6841,N_6813);
xnor U7262 (N_7262,N_6741,N_6828);
xor U7263 (N_7263,N_6769,N_6737);
and U7264 (N_7264,N_6542,N_6828);
nor U7265 (N_7265,N_6641,N_6789);
nand U7266 (N_7266,N_6846,N_6668);
nor U7267 (N_7267,N_6969,N_6644);
nand U7268 (N_7268,N_6812,N_6965);
nor U7269 (N_7269,N_6589,N_6563);
nor U7270 (N_7270,N_6956,N_6721);
nand U7271 (N_7271,N_6764,N_6689);
xor U7272 (N_7272,N_6956,N_6868);
and U7273 (N_7273,N_6944,N_6795);
nand U7274 (N_7274,N_6898,N_6712);
nor U7275 (N_7275,N_6956,N_6510);
nor U7276 (N_7276,N_6774,N_6816);
or U7277 (N_7277,N_6539,N_6656);
nor U7278 (N_7278,N_6771,N_6994);
nand U7279 (N_7279,N_6587,N_6580);
or U7280 (N_7280,N_6685,N_6919);
nand U7281 (N_7281,N_6650,N_6786);
nor U7282 (N_7282,N_6630,N_6784);
or U7283 (N_7283,N_6828,N_6599);
or U7284 (N_7284,N_6738,N_6500);
or U7285 (N_7285,N_6874,N_6576);
nand U7286 (N_7286,N_6558,N_6683);
nor U7287 (N_7287,N_6748,N_6533);
nand U7288 (N_7288,N_6612,N_6546);
nor U7289 (N_7289,N_6962,N_6676);
xnor U7290 (N_7290,N_6612,N_6920);
nor U7291 (N_7291,N_6564,N_6509);
nor U7292 (N_7292,N_6789,N_6818);
and U7293 (N_7293,N_6773,N_6706);
xor U7294 (N_7294,N_6987,N_6932);
nand U7295 (N_7295,N_6868,N_6569);
and U7296 (N_7296,N_6937,N_6837);
nand U7297 (N_7297,N_6848,N_6883);
nor U7298 (N_7298,N_6763,N_6790);
or U7299 (N_7299,N_6564,N_6537);
and U7300 (N_7300,N_6591,N_6835);
and U7301 (N_7301,N_6820,N_6983);
xnor U7302 (N_7302,N_6561,N_6686);
or U7303 (N_7303,N_6591,N_6729);
xnor U7304 (N_7304,N_6901,N_6894);
or U7305 (N_7305,N_6684,N_6746);
nand U7306 (N_7306,N_6563,N_6746);
xor U7307 (N_7307,N_6727,N_6685);
nor U7308 (N_7308,N_6613,N_6843);
and U7309 (N_7309,N_6705,N_6513);
nand U7310 (N_7310,N_6654,N_6633);
nor U7311 (N_7311,N_6744,N_6871);
or U7312 (N_7312,N_6863,N_6933);
xor U7313 (N_7313,N_6980,N_6817);
or U7314 (N_7314,N_6943,N_6971);
nand U7315 (N_7315,N_6548,N_6514);
xnor U7316 (N_7316,N_6848,N_6530);
and U7317 (N_7317,N_6723,N_6873);
nand U7318 (N_7318,N_6937,N_6948);
and U7319 (N_7319,N_6911,N_6996);
and U7320 (N_7320,N_6812,N_6696);
nand U7321 (N_7321,N_6513,N_6957);
nand U7322 (N_7322,N_6817,N_6779);
and U7323 (N_7323,N_6972,N_6934);
xor U7324 (N_7324,N_6967,N_6880);
xor U7325 (N_7325,N_6782,N_6825);
and U7326 (N_7326,N_6585,N_6710);
and U7327 (N_7327,N_6594,N_6748);
xnor U7328 (N_7328,N_6891,N_6857);
and U7329 (N_7329,N_6547,N_6883);
nand U7330 (N_7330,N_6735,N_6839);
nor U7331 (N_7331,N_6519,N_6724);
nor U7332 (N_7332,N_6901,N_6652);
nor U7333 (N_7333,N_6541,N_6774);
or U7334 (N_7334,N_6638,N_6924);
xor U7335 (N_7335,N_6639,N_6873);
nand U7336 (N_7336,N_6712,N_6648);
nand U7337 (N_7337,N_6884,N_6637);
nor U7338 (N_7338,N_6942,N_6884);
nand U7339 (N_7339,N_6915,N_6533);
or U7340 (N_7340,N_6918,N_6585);
and U7341 (N_7341,N_6547,N_6661);
and U7342 (N_7342,N_6593,N_6527);
and U7343 (N_7343,N_6574,N_6715);
nor U7344 (N_7344,N_6636,N_6503);
or U7345 (N_7345,N_6903,N_6555);
xnor U7346 (N_7346,N_6700,N_6932);
nor U7347 (N_7347,N_6841,N_6704);
xor U7348 (N_7348,N_6740,N_6928);
or U7349 (N_7349,N_6706,N_6807);
xor U7350 (N_7350,N_6548,N_6849);
xnor U7351 (N_7351,N_6759,N_6944);
xor U7352 (N_7352,N_6772,N_6632);
or U7353 (N_7353,N_6919,N_6535);
and U7354 (N_7354,N_6841,N_6900);
nand U7355 (N_7355,N_6918,N_6516);
or U7356 (N_7356,N_6699,N_6565);
and U7357 (N_7357,N_6901,N_6681);
nor U7358 (N_7358,N_6824,N_6551);
nand U7359 (N_7359,N_6517,N_6978);
xor U7360 (N_7360,N_6591,N_6758);
nand U7361 (N_7361,N_6746,N_6892);
and U7362 (N_7362,N_6518,N_6792);
nor U7363 (N_7363,N_6931,N_6756);
nor U7364 (N_7364,N_6519,N_6707);
and U7365 (N_7365,N_6677,N_6731);
and U7366 (N_7366,N_6610,N_6689);
xor U7367 (N_7367,N_6828,N_6714);
nor U7368 (N_7368,N_6919,N_6538);
or U7369 (N_7369,N_6504,N_6773);
or U7370 (N_7370,N_6878,N_6963);
nand U7371 (N_7371,N_6941,N_6942);
or U7372 (N_7372,N_6957,N_6767);
nor U7373 (N_7373,N_6802,N_6769);
nor U7374 (N_7374,N_6986,N_6657);
nor U7375 (N_7375,N_6844,N_6736);
nand U7376 (N_7376,N_6908,N_6826);
nand U7377 (N_7377,N_6713,N_6575);
or U7378 (N_7378,N_6827,N_6718);
and U7379 (N_7379,N_6923,N_6893);
nand U7380 (N_7380,N_6618,N_6883);
nand U7381 (N_7381,N_6724,N_6688);
xnor U7382 (N_7382,N_6559,N_6750);
or U7383 (N_7383,N_6529,N_6964);
or U7384 (N_7384,N_6770,N_6621);
xor U7385 (N_7385,N_6537,N_6507);
or U7386 (N_7386,N_6658,N_6617);
nand U7387 (N_7387,N_6586,N_6948);
nor U7388 (N_7388,N_6888,N_6595);
nand U7389 (N_7389,N_6803,N_6747);
xnor U7390 (N_7390,N_6699,N_6736);
xnor U7391 (N_7391,N_6966,N_6862);
or U7392 (N_7392,N_6581,N_6793);
and U7393 (N_7393,N_6615,N_6832);
or U7394 (N_7394,N_6867,N_6933);
xor U7395 (N_7395,N_6695,N_6623);
nor U7396 (N_7396,N_6631,N_6892);
and U7397 (N_7397,N_6867,N_6563);
or U7398 (N_7398,N_6884,N_6856);
nor U7399 (N_7399,N_6988,N_6862);
nor U7400 (N_7400,N_6527,N_6666);
nand U7401 (N_7401,N_6744,N_6570);
nor U7402 (N_7402,N_6924,N_6706);
nor U7403 (N_7403,N_6748,N_6825);
or U7404 (N_7404,N_6742,N_6688);
xnor U7405 (N_7405,N_6829,N_6925);
xor U7406 (N_7406,N_6794,N_6989);
nand U7407 (N_7407,N_6845,N_6781);
xor U7408 (N_7408,N_6741,N_6667);
or U7409 (N_7409,N_6963,N_6694);
xor U7410 (N_7410,N_6676,N_6585);
or U7411 (N_7411,N_6610,N_6892);
and U7412 (N_7412,N_6668,N_6853);
or U7413 (N_7413,N_6967,N_6974);
nor U7414 (N_7414,N_6854,N_6972);
xnor U7415 (N_7415,N_6808,N_6716);
nand U7416 (N_7416,N_6710,N_6650);
nand U7417 (N_7417,N_6855,N_6989);
xnor U7418 (N_7418,N_6804,N_6612);
nor U7419 (N_7419,N_6567,N_6598);
xor U7420 (N_7420,N_6741,N_6654);
or U7421 (N_7421,N_6796,N_6642);
xnor U7422 (N_7422,N_6650,N_6966);
nor U7423 (N_7423,N_6856,N_6528);
nand U7424 (N_7424,N_6988,N_6851);
or U7425 (N_7425,N_6554,N_6544);
xnor U7426 (N_7426,N_6601,N_6779);
xor U7427 (N_7427,N_6845,N_6562);
nor U7428 (N_7428,N_6912,N_6801);
xnor U7429 (N_7429,N_6862,N_6858);
nor U7430 (N_7430,N_6572,N_6521);
and U7431 (N_7431,N_6630,N_6891);
nand U7432 (N_7432,N_6670,N_6659);
or U7433 (N_7433,N_6614,N_6620);
or U7434 (N_7434,N_6933,N_6629);
nor U7435 (N_7435,N_6792,N_6587);
nand U7436 (N_7436,N_6652,N_6949);
nor U7437 (N_7437,N_6683,N_6633);
nor U7438 (N_7438,N_6841,N_6593);
and U7439 (N_7439,N_6918,N_6695);
nand U7440 (N_7440,N_6986,N_6597);
xnor U7441 (N_7441,N_6616,N_6926);
xor U7442 (N_7442,N_6708,N_6728);
nor U7443 (N_7443,N_6641,N_6921);
nor U7444 (N_7444,N_6815,N_6615);
nor U7445 (N_7445,N_6719,N_6735);
nand U7446 (N_7446,N_6710,N_6887);
xor U7447 (N_7447,N_6875,N_6698);
or U7448 (N_7448,N_6739,N_6756);
nor U7449 (N_7449,N_6811,N_6596);
nor U7450 (N_7450,N_6852,N_6874);
and U7451 (N_7451,N_6865,N_6973);
nor U7452 (N_7452,N_6728,N_6601);
nor U7453 (N_7453,N_6890,N_6998);
or U7454 (N_7454,N_6596,N_6633);
or U7455 (N_7455,N_6932,N_6948);
nand U7456 (N_7456,N_6656,N_6586);
or U7457 (N_7457,N_6804,N_6569);
nand U7458 (N_7458,N_6956,N_6506);
nand U7459 (N_7459,N_6683,N_6669);
xor U7460 (N_7460,N_6924,N_6942);
xnor U7461 (N_7461,N_6872,N_6838);
xor U7462 (N_7462,N_6696,N_6751);
and U7463 (N_7463,N_6825,N_6916);
and U7464 (N_7464,N_6994,N_6938);
or U7465 (N_7465,N_6541,N_6880);
or U7466 (N_7466,N_6824,N_6569);
nand U7467 (N_7467,N_6897,N_6855);
or U7468 (N_7468,N_6631,N_6732);
or U7469 (N_7469,N_6810,N_6571);
nand U7470 (N_7470,N_6539,N_6820);
or U7471 (N_7471,N_6530,N_6795);
nand U7472 (N_7472,N_6561,N_6650);
nand U7473 (N_7473,N_6690,N_6921);
and U7474 (N_7474,N_6677,N_6642);
xor U7475 (N_7475,N_6624,N_6628);
nor U7476 (N_7476,N_6640,N_6516);
nor U7477 (N_7477,N_6905,N_6664);
or U7478 (N_7478,N_6775,N_6872);
nand U7479 (N_7479,N_6806,N_6643);
nor U7480 (N_7480,N_6509,N_6827);
nand U7481 (N_7481,N_6524,N_6658);
nand U7482 (N_7482,N_6837,N_6558);
and U7483 (N_7483,N_6945,N_6630);
xor U7484 (N_7484,N_6587,N_6678);
nor U7485 (N_7485,N_6855,N_6589);
and U7486 (N_7486,N_6738,N_6994);
or U7487 (N_7487,N_6924,N_6605);
xor U7488 (N_7488,N_6944,N_6679);
or U7489 (N_7489,N_6983,N_6566);
or U7490 (N_7490,N_6830,N_6952);
nor U7491 (N_7491,N_6747,N_6549);
nor U7492 (N_7492,N_6577,N_6651);
nor U7493 (N_7493,N_6736,N_6995);
nor U7494 (N_7494,N_6705,N_6807);
or U7495 (N_7495,N_6840,N_6557);
nor U7496 (N_7496,N_6912,N_6763);
nor U7497 (N_7497,N_6871,N_6852);
xnor U7498 (N_7498,N_6774,N_6855);
nand U7499 (N_7499,N_6805,N_6642);
nor U7500 (N_7500,N_7150,N_7065);
or U7501 (N_7501,N_7446,N_7130);
nor U7502 (N_7502,N_7124,N_7141);
nor U7503 (N_7503,N_7139,N_7306);
nor U7504 (N_7504,N_7222,N_7485);
or U7505 (N_7505,N_7027,N_7015);
nor U7506 (N_7506,N_7285,N_7350);
and U7507 (N_7507,N_7283,N_7380);
nor U7508 (N_7508,N_7120,N_7125);
xor U7509 (N_7509,N_7046,N_7236);
xnor U7510 (N_7510,N_7345,N_7189);
nor U7511 (N_7511,N_7491,N_7068);
or U7512 (N_7512,N_7374,N_7220);
nand U7513 (N_7513,N_7296,N_7223);
or U7514 (N_7514,N_7021,N_7392);
nand U7515 (N_7515,N_7096,N_7209);
and U7516 (N_7516,N_7472,N_7231);
nor U7517 (N_7517,N_7254,N_7430);
nor U7518 (N_7518,N_7421,N_7369);
nor U7519 (N_7519,N_7084,N_7034);
or U7520 (N_7520,N_7171,N_7023);
and U7521 (N_7521,N_7388,N_7211);
and U7522 (N_7522,N_7303,N_7198);
nor U7523 (N_7523,N_7357,N_7429);
and U7524 (N_7524,N_7230,N_7183);
nand U7525 (N_7525,N_7343,N_7473);
nand U7526 (N_7526,N_7381,N_7165);
nor U7527 (N_7527,N_7269,N_7062);
xor U7528 (N_7528,N_7090,N_7455);
and U7529 (N_7529,N_7358,N_7266);
nand U7530 (N_7530,N_7241,N_7174);
or U7531 (N_7531,N_7496,N_7397);
nand U7532 (N_7532,N_7178,N_7041);
nor U7533 (N_7533,N_7323,N_7272);
nand U7534 (N_7534,N_7190,N_7099);
or U7535 (N_7535,N_7408,N_7404);
or U7536 (N_7536,N_7252,N_7024);
or U7537 (N_7537,N_7103,N_7310);
and U7538 (N_7538,N_7137,N_7438);
nand U7539 (N_7539,N_7471,N_7295);
nor U7540 (N_7540,N_7132,N_7032);
nand U7541 (N_7541,N_7423,N_7131);
nor U7542 (N_7542,N_7251,N_7179);
or U7543 (N_7543,N_7436,N_7441);
nand U7544 (N_7544,N_7087,N_7080);
or U7545 (N_7545,N_7426,N_7164);
and U7546 (N_7546,N_7460,N_7278);
xnor U7547 (N_7547,N_7177,N_7005);
nor U7548 (N_7548,N_7000,N_7051);
nor U7549 (N_7549,N_7271,N_7093);
nor U7550 (N_7550,N_7454,N_7347);
and U7551 (N_7551,N_7203,N_7311);
xor U7552 (N_7552,N_7001,N_7199);
xnor U7553 (N_7553,N_7086,N_7258);
nand U7554 (N_7554,N_7243,N_7493);
and U7555 (N_7555,N_7273,N_7147);
and U7556 (N_7556,N_7242,N_7465);
nor U7557 (N_7557,N_7308,N_7486);
or U7558 (N_7558,N_7011,N_7144);
or U7559 (N_7559,N_7387,N_7229);
xor U7560 (N_7560,N_7158,N_7031);
nand U7561 (N_7561,N_7324,N_7365);
xor U7562 (N_7562,N_7316,N_7201);
or U7563 (N_7563,N_7420,N_7386);
or U7564 (N_7564,N_7287,N_7302);
nor U7565 (N_7565,N_7235,N_7371);
xnor U7566 (N_7566,N_7204,N_7444);
nor U7567 (N_7567,N_7116,N_7325);
and U7568 (N_7568,N_7006,N_7044);
nand U7569 (N_7569,N_7063,N_7092);
and U7570 (N_7570,N_7342,N_7362);
nor U7571 (N_7571,N_7028,N_7425);
nor U7572 (N_7572,N_7340,N_7136);
nor U7573 (N_7573,N_7114,N_7205);
and U7574 (N_7574,N_7334,N_7361);
or U7575 (N_7575,N_7246,N_7354);
and U7576 (N_7576,N_7176,N_7383);
or U7577 (N_7577,N_7240,N_7359);
nor U7578 (N_7578,N_7221,N_7284);
nand U7579 (N_7579,N_7403,N_7385);
nand U7580 (N_7580,N_7257,N_7428);
and U7581 (N_7581,N_7298,N_7218);
or U7582 (N_7582,N_7217,N_7344);
nor U7583 (N_7583,N_7082,N_7382);
xnor U7584 (N_7584,N_7039,N_7250);
xnor U7585 (N_7585,N_7304,N_7160);
nor U7586 (N_7586,N_7346,N_7315);
and U7587 (N_7587,N_7094,N_7356);
nor U7588 (N_7588,N_7477,N_7076);
nand U7589 (N_7589,N_7053,N_7018);
nand U7590 (N_7590,N_7212,N_7047);
nand U7591 (N_7591,N_7059,N_7305);
nor U7592 (N_7592,N_7100,N_7012);
and U7593 (N_7593,N_7464,N_7475);
and U7594 (N_7594,N_7140,N_7108);
nand U7595 (N_7595,N_7153,N_7418);
xor U7596 (N_7596,N_7476,N_7291);
nor U7597 (N_7597,N_7327,N_7301);
or U7598 (N_7598,N_7413,N_7233);
nor U7599 (N_7599,N_7279,N_7170);
and U7600 (N_7600,N_7196,N_7148);
or U7601 (N_7601,N_7417,N_7469);
nand U7602 (N_7602,N_7280,N_7339);
xor U7603 (N_7603,N_7110,N_7091);
and U7604 (N_7604,N_7297,N_7121);
xor U7605 (N_7605,N_7187,N_7307);
and U7606 (N_7606,N_7260,N_7489);
nor U7607 (N_7607,N_7262,N_7329);
xor U7608 (N_7608,N_7411,N_7225);
or U7609 (N_7609,N_7452,N_7433);
nand U7610 (N_7610,N_7073,N_7451);
xor U7611 (N_7611,N_7427,N_7497);
or U7612 (N_7612,N_7450,N_7267);
nor U7613 (N_7613,N_7331,N_7159);
and U7614 (N_7614,N_7249,N_7293);
nand U7615 (N_7615,N_7321,N_7461);
and U7616 (N_7616,N_7393,N_7234);
nor U7617 (N_7617,N_7195,N_7069);
or U7618 (N_7618,N_7363,N_7341);
nand U7619 (N_7619,N_7416,N_7332);
and U7620 (N_7620,N_7134,N_7168);
and U7621 (N_7621,N_7226,N_7399);
nor U7622 (N_7622,N_7088,N_7289);
nor U7623 (N_7623,N_7457,N_7415);
nor U7624 (N_7624,N_7122,N_7490);
nand U7625 (N_7625,N_7017,N_7435);
and U7626 (N_7626,N_7364,N_7057);
or U7627 (N_7627,N_7202,N_7412);
nor U7628 (N_7628,N_7245,N_7424);
nor U7629 (N_7629,N_7194,N_7419);
and U7630 (N_7630,N_7377,N_7089);
nor U7631 (N_7631,N_7247,N_7228);
nand U7632 (N_7632,N_7030,N_7155);
nor U7633 (N_7633,N_7142,N_7055);
or U7634 (N_7634,N_7318,N_7468);
or U7635 (N_7635,N_7276,N_7462);
and U7636 (N_7636,N_7210,N_7395);
or U7637 (N_7637,N_7330,N_7098);
or U7638 (N_7638,N_7216,N_7402);
or U7639 (N_7639,N_7050,N_7135);
or U7640 (N_7640,N_7264,N_7227);
xnor U7641 (N_7641,N_7104,N_7274);
or U7642 (N_7642,N_7186,N_7107);
and U7643 (N_7643,N_7035,N_7238);
xnor U7644 (N_7644,N_7167,N_7169);
xnor U7645 (N_7645,N_7482,N_7478);
and U7646 (N_7646,N_7463,N_7379);
or U7647 (N_7647,N_7275,N_7317);
or U7648 (N_7648,N_7193,N_7109);
xnor U7649 (N_7649,N_7097,N_7045);
xor U7650 (N_7650,N_7064,N_7237);
and U7651 (N_7651,N_7286,N_7398);
xnor U7652 (N_7652,N_7367,N_7085);
or U7653 (N_7653,N_7111,N_7002);
nor U7654 (N_7654,N_7129,N_7467);
nor U7655 (N_7655,N_7326,N_7095);
and U7656 (N_7656,N_7390,N_7070);
xnor U7657 (N_7657,N_7016,N_7410);
xor U7658 (N_7658,N_7447,N_7375);
nand U7659 (N_7659,N_7391,N_7355);
and U7660 (N_7660,N_7470,N_7256);
xnor U7661 (N_7661,N_7014,N_7396);
and U7662 (N_7662,N_7060,N_7054);
xor U7663 (N_7663,N_7352,N_7061);
nor U7664 (N_7664,N_7113,N_7081);
xnor U7665 (N_7665,N_7128,N_7040);
nand U7666 (N_7666,N_7299,N_7029);
xor U7667 (N_7667,N_7019,N_7349);
xor U7668 (N_7668,N_7025,N_7072);
nor U7669 (N_7669,N_7488,N_7052);
or U7670 (N_7670,N_7338,N_7495);
or U7671 (N_7671,N_7138,N_7492);
nor U7672 (N_7672,N_7115,N_7117);
or U7673 (N_7673,N_7077,N_7145);
nor U7674 (N_7674,N_7290,N_7154);
xnor U7675 (N_7675,N_7105,N_7008);
and U7676 (N_7676,N_7373,N_7337);
nor U7677 (N_7677,N_7048,N_7414);
nor U7678 (N_7678,N_7182,N_7188);
or U7679 (N_7679,N_7214,N_7009);
xor U7680 (N_7680,N_7172,N_7185);
or U7681 (N_7681,N_7456,N_7127);
nor U7682 (N_7682,N_7206,N_7437);
and U7683 (N_7683,N_7022,N_7376);
and U7684 (N_7684,N_7314,N_7253);
nor U7685 (N_7685,N_7149,N_7288);
xnor U7686 (N_7686,N_7440,N_7036);
xnor U7687 (N_7687,N_7434,N_7366);
nand U7688 (N_7688,N_7265,N_7431);
xnor U7689 (N_7689,N_7261,N_7038);
nand U7690 (N_7690,N_7268,N_7207);
xnor U7691 (N_7691,N_7056,N_7432);
xnor U7692 (N_7692,N_7439,N_7333);
or U7693 (N_7693,N_7370,N_7405);
or U7694 (N_7694,N_7156,N_7479);
nor U7695 (N_7695,N_7407,N_7033);
or U7696 (N_7696,N_7078,N_7200);
xor U7697 (N_7697,N_7152,N_7058);
nand U7698 (N_7698,N_7320,N_7010);
and U7699 (N_7699,N_7197,N_7083);
nand U7700 (N_7700,N_7215,N_7409);
and U7701 (N_7701,N_7401,N_7074);
and U7702 (N_7702,N_7394,N_7255);
or U7703 (N_7703,N_7348,N_7020);
and U7704 (N_7704,N_7213,N_7270);
or U7705 (N_7705,N_7474,N_7184);
and U7706 (N_7706,N_7281,N_7162);
or U7707 (N_7707,N_7498,N_7157);
or U7708 (N_7708,N_7487,N_7384);
nor U7709 (N_7709,N_7481,N_7119);
nand U7710 (N_7710,N_7353,N_7312);
xnor U7711 (N_7711,N_7466,N_7004);
and U7712 (N_7712,N_7300,N_7313);
xor U7713 (N_7713,N_7143,N_7037);
and U7714 (N_7714,N_7049,N_7224);
xor U7715 (N_7715,N_7239,N_7494);
nand U7716 (N_7716,N_7043,N_7079);
or U7717 (N_7717,N_7118,N_7003);
xnor U7718 (N_7718,N_7232,N_7335);
nand U7719 (N_7719,N_7042,N_7181);
or U7720 (N_7720,N_7101,N_7442);
xor U7721 (N_7721,N_7173,N_7459);
xnor U7722 (N_7722,N_7309,N_7453);
nand U7723 (N_7723,N_7259,N_7483);
or U7724 (N_7724,N_7484,N_7406);
nor U7725 (N_7725,N_7071,N_7146);
nor U7726 (N_7726,N_7123,N_7208);
or U7727 (N_7727,N_7126,N_7328);
xnor U7728 (N_7728,N_7106,N_7219);
nand U7729 (N_7729,N_7422,N_7389);
and U7730 (N_7730,N_7351,N_7448);
nor U7731 (N_7731,N_7248,N_7180);
and U7732 (N_7732,N_7458,N_7166);
nand U7733 (N_7733,N_7322,N_7066);
nand U7734 (N_7734,N_7112,N_7360);
and U7735 (N_7735,N_7192,N_7244);
or U7736 (N_7736,N_7151,N_7319);
xnor U7737 (N_7737,N_7102,N_7191);
nor U7738 (N_7738,N_7292,N_7443);
xnor U7739 (N_7739,N_7445,N_7449);
nor U7740 (N_7740,N_7075,N_7480);
or U7741 (N_7741,N_7007,N_7161);
nand U7742 (N_7742,N_7372,N_7282);
nor U7743 (N_7743,N_7163,N_7026);
nor U7744 (N_7744,N_7499,N_7400);
or U7745 (N_7745,N_7013,N_7378);
nor U7746 (N_7746,N_7263,N_7368);
nand U7747 (N_7747,N_7336,N_7175);
nor U7748 (N_7748,N_7133,N_7277);
nand U7749 (N_7749,N_7067,N_7294);
or U7750 (N_7750,N_7316,N_7233);
nor U7751 (N_7751,N_7269,N_7271);
and U7752 (N_7752,N_7297,N_7123);
or U7753 (N_7753,N_7463,N_7357);
and U7754 (N_7754,N_7437,N_7040);
nor U7755 (N_7755,N_7391,N_7020);
or U7756 (N_7756,N_7193,N_7310);
and U7757 (N_7757,N_7210,N_7473);
nand U7758 (N_7758,N_7313,N_7070);
nand U7759 (N_7759,N_7282,N_7054);
and U7760 (N_7760,N_7291,N_7255);
xor U7761 (N_7761,N_7346,N_7017);
and U7762 (N_7762,N_7334,N_7012);
and U7763 (N_7763,N_7229,N_7415);
nor U7764 (N_7764,N_7086,N_7425);
nor U7765 (N_7765,N_7087,N_7411);
xnor U7766 (N_7766,N_7055,N_7399);
nand U7767 (N_7767,N_7150,N_7199);
and U7768 (N_7768,N_7392,N_7029);
nor U7769 (N_7769,N_7436,N_7102);
nand U7770 (N_7770,N_7034,N_7229);
or U7771 (N_7771,N_7098,N_7351);
xor U7772 (N_7772,N_7419,N_7172);
xor U7773 (N_7773,N_7347,N_7036);
nor U7774 (N_7774,N_7196,N_7338);
xnor U7775 (N_7775,N_7347,N_7403);
and U7776 (N_7776,N_7085,N_7282);
or U7777 (N_7777,N_7003,N_7077);
or U7778 (N_7778,N_7239,N_7008);
and U7779 (N_7779,N_7044,N_7262);
nor U7780 (N_7780,N_7352,N_7429);
and U7781 (N_7781,N_7086,N_7000);
xnor U7782 (N_7782,N_7433,N_7076);
nor U7783 (N_7783,N_7153,N_7242);
nand U7784 (N_7784,N_7077,N_7356);
nor U7785 (N_7785,N_7151,N_7347);
nor U7786 (N_7786,N_7176,N_7245);
xor U7787 (N_7787,N_7250,N_7267);
nand U7788 (N_7788,N_7211,N_7025);
nand U7789 (N_7789,N_7415,N_7408);
and U7790 (N_7790,N_7168,N_7268);
and U7791 (N_7791,N_7300,N_7074);
nor U7792 (N_7792,N_7055,N_7353);
nand U7793 (N_7793,N_7328,N_7043);
or U7794 (N_7794,N_7290,N_7081);
nor U7795 (N_7795,N_7399,N_7242);
nand U7796 (N_7796,N_7281,N_7468);
nor U7797 (N_7797,N_7170,N_7208);
or U7798 (N_7798,N_7365,N_7348);
and U7799 (N_7799,N_7405,N_7051);
xnor U7800 (N_7800,N_7152,N_7134);
nor U7801 (N_7801,N_7353,N_7346);
and U7802 (N_7802,N_7274,N_7440);
nand U7803 (N_7803,N_7316,N_7133);
and U7804 (N_7804,N_7106,N_7273);
nand U7805 (N_7805,N_7132,N_7405);
nor U7806 (N_7806,N_7189,N_7097);
xnor U7807 (N_7807,N_7298,N_7163);
xnor U7808 (N_7808,N_7308,N_7056);
or U7809 (N_7809,N_7339,N_7254);
nor U7810 (N_7810,N_7273,N_7242);
nand U7811 (N_7811,N_7236,N_7047);
xor U7812 (N_7812,N_7096,N_7166);
and U7813 (N_7813,N_7360,N_7008);
xor U7814 (N_7814,N_7070,N_7449);
and U7815 (N_7815,N_7039,N_7482);
nor U7816 (N_7816,N_7344,N_7222);
nor U7817 (N_7817,N_7211,N_7401);
or U7818 (N_7818,N_7161,N_7044);
or U7819 (N_7819,N_7198,N_7246);
and U7820 (N_7820,N_7446,N_7266);
xnor U7821 (N_7821,N_7323,N_7237);
nand U7822 (N_7822,N_7479,N_7491);
nand U7823 (N_7823,N_7409,N_7169);
or U7824 (N_7824,N_7011,N_7041);
or U7825 (N_7825,N_7080,N_7106);
and U7826 (N_7826,N_7034,N_7099);
nand U7827 (N_7827,N_7030,N_7224);
nand U7828 (N_7828,N_7101,N_7240);
or U7829 (N_7829,N_7281,N_7280);
or U7830 (N_7830,N_7107,N_7329);
xor U7831 (N_7831,N_7015,N_7192);
xor U7832 (N_7832,N_7233,N_7240);
and U7833 (N_7833,N_7262,N_7479);
xor U7834 (N_7834,N_7194,N_7004);
or U7835 (N_7835,N_7204,N_7240);
and U7836 (N_7836,N_7235,N_7049);
xor U7837 (N_7837,N_7449,N_7035);
or U7838 (N_7838,N_7108,N_7253);
and U7839 (N_7839,N_7399,N_7488);
xnor U7840 (N_7840,N_7182,N_7276);
nor U7841 (N_7841,N_7030,N_7126);
xnor U7842 (N_7842,N_7424,N_7296);
nand U7843 (N_7843,N_7087,N_7237);
and U7844 (N_7844,N_7193,N_7298);
xnor U7845 (N_7845,N_7236,N_7224);
xnor U7846 (N_7846,N_7337,N_7124);
or U7847 (N_7847,N_7095,N_7215);
and U7848 (N_7848,N_7372,N_7244);
or U7849 (N_7849,N_7479,N_7399);
nor U7850 (N_7850,N_7094,N_7147);
or U7851 (N_7851,N_7060,N_7207);
nand U7852 (N_7852,N_7236,N_7012);
and U7853 (N_7853,N_7026,N_7299);
or U7854 (N_7854,N_7117,N_7113);
nor U7855 (N_7855,N_7089,N_7497);
xor U7856 (N_7856,N_7113,N_7090);
and U7857 (N_7857,N_7361,N_7368);
or U7858 (N_7858,N_7106,N_7130);
nor U7859 (N_7859,N_7461,N_7347);
xor U7860 (N_7860,N_7360,N_7240);
or U7861 (N_7861,N_7372,N_7182);
and U7862 (N_7862,N_7274,N_7304);
nand U7863 (N_7863,N_7474,N_7189);
and U7864 (N_7864,N_7204,N_7248);
nand U7865 (N_7865,N_7328,N_7318);
or U7866 (N_7866,N_7361,N_7483);
nand U7867 (N_7867,N_7238,N_7422);
and U7868 (N_7868,N_7337,N_7324);
nor U7869 (N_7869,N_7081,N_7457);
nor U7870 (N_7870,N_7389,N_7223);
or U7871 (N_7871,N_7141,N_7454);
or U7872 (N_7872,N_7176,N_7112);
nor U7873 (N_7873,N_7166,N_7198);
xnor U7874 (N_7874,N_7141,N_7191);
nor U7875 (N_7875,N_7298,N_7321);
and U7876 (N_7876,N_7415,N_7157);
and U7877 (N_7877,N_7221,N_7098);
nand U7878 (N_7878,N_7307,N_7283);
xnor U7879 (N_7879,N_7363,N_7184);
nor U7880 (N_7880,N_7089,N_7468);
and U7881 (N_7881,N_7328,N_7154);
or U7882 (N_7882,N_7091,N_7190);
or U7883 (N_7883,N_7103,N_7174);
nor U7884 (N_7884,N_7076,N_7086);
xnor U7885 (N_7885,N_7083,N_7069);
xnor U7886 (N_7886,N_7070,N_7366);
nand U7887 (N_7887,N_7058,N_7249);
nor U7888 (N_7888,N_7351,N_7420);
and U7889 (N_7889,N_7215,N_7255);
and U7890 (N_7890,N_7491,N_7332);
and U7891 (N_7891,N_7059,N_7290);
xnor U7892 (N_7892,N_7245,N_7487);
or U7893 (N_7893,N_7373,N_7473);
nand U7894 (N_7894,N_7462,N_7367);
xor U7895 (N_7895,N_7255,N_7194);
or U7896 (N_7896,N_7117,N_7074);
nor U7897 (N_7897,N_7286,N_7468);
xnor U7898 (N_7898,N_7035,N_7236);
nand U7899 (N_7899,N_7117,N_7324);
xnor U7900 (N_7900,N_7088,N_7402);
nor U7901 (N_7901,N_7116,N_7191);
and U7902 (N_7902,N_7441,N_7337);
and U7903 (N_7903,N_7075,N_7083);
nor U7904 (N_7904,N_7469,N_7002);
nor U7905 (N_7905,N_7484,N_7140);
xnor U7906 (N_7906,N_7293,N_7443);
nor U7907 (N_7907,N_7258,N_7336);
nand U7908 (N_7908,N_7113,N_7453);
or U7909 (N_7909,N_7289,N_7150);
and U7910 (N_7910,N_7471,N_7106);
nor U7911 (N_7911,N_7338,N_7328);
nand U7912 (N_7912,N_7243,N_7050);
and U7913 (N_7913,N_7049,N_7473);
and U7914 (N_7914,N_7262,N_7182);
and U7915 (N_7915,N_7063,N_7388);
nand U7916 (N_7916,N_7491,N_7212);
or U7917 (N_7917,N_7435,N_7342);
or U7918 (N_7918,N_7194,N_7238);
nor U7919 (N_7919,N_7230,N_7062);
xor U7920 (N_7920,N_7032,N_7428);
nand U7921 (N_7921,N_7455,N_7473);
and U7922 (N_7922,N_7197,N_7127);
and U7923 (N_7923,N_7364,N_7004);
nor U7924 (N_7924,N_7370,N_7066);
and U7925 (N_7925,N_7293,N_7340);
nand U7926 (N_7926,N_7120,N_7424);
and U7927 (N_7927,N_7412,N_7400);
xnor U7928 (N_7928,N_7163,N_7434);
or U7929 (N_7929,N_7170,N_7354);
nand U7930 (N_7930,N_7065,N_7062);
and U7931 (N_7931,N_7175,N_7450);
nor U7932 (N_7932,N_7154,N_7291);
and U7933 (N_7933,N_7497,N_7083);
and U7934 (N_7934,N_7252,N_7137);
xor U7935 (N_7935,N_7469,N_7444);
nor U7936 (N_7936,N_7031,N_7397);
nor U7937 (N_7937,N_7199,N_7086);
or U7938 (N_7938,N_7127,N_7382);
nor U7939 (N_7939,N_7096,N_7017);
and U7940 (N_7940,N_7284,N_7040);
xnor U7941 (N_7941,N_7301,N_7483);
or U7942 (N_7942,N_7029,N_7169);
xnor U7943 (N_7943,N_7116,N_7345);
nand U7944 (N_7944,N_7371,N_7449);
xor U7945 (N_7945,N_7008,N_7162);
nor U7946 (N_7946,N_7466,N_7187);
and U7947 (N_7947,N_7473,N_7015);
and U7948 (N_7948,N_7397,N_7431);
or U7949 (N_7949,N_7385,N_7137);
xnor U7950 (N_7950,N_7252,N_7131);
nand U7951 (N_7951,N_7217,N_7260);
nand U7952 (N_7952,N_7016,N_7146);
and U7953 (N_7953,N_7411,N_7421);
nand U7954 (N_7954,N_7057,N_7395);
xor U7955 (N_7955,N_7297,N_7097);
xnor U7956 (N_7956,N_7370,N_7442);
xor U7957 (N_7957,N_7461,N_7445);
nand U7958 (N_7958,N_7154,N_7343);
nor U7959 (N_7959,N_7049,N_7182);
or U7960 (N_7960,N_7266,N_7119);
or U7961 (N_7961,N_7326,N_7080);
and U7962 (N_7962,N_7337,N_7315);
or U7963 (N_7963,N_7162,N_7473);
xor U7964 (N_7964,N_7482,N_7006);
nand U7965 (N_7965,N_7422,N_7365);
xnor U7966 (N_7966,N_7416,N_7255);
nand U7967 (N_7967,N_7210,N_7378);
nand U7968 (N_7968,N_7138,N_7481);
xor U7969 (N_7969,N_7399,N_7215);
nand U7970 (N_7970,N_7123,N_7321);
xor U7971 (N_7971,N_7307,N_7409);
xor U7972 (N_7972,N_7064,N_7013);
nand U7973 (N_7973,N_7375,N_7253);
nand U7974 (N_7974,N_7161,N_7367);
nand U7975 (N_7975,N_7120,N_7081);
xor U7976 (N_7976,N_7028,N_7128);
xnor U7977 (N_7977,N_7329,N_7270);
xnor U7978 (N_7978,N_7388,N_7146);
xor U7979 (N_7979,N_7070,N_7003);
nand U7980 (N_7980,N_7418,N_7257);
xnor U7981 (N_7981,N_7429,N_7192);
and U7982 (N_7982,N_7444,N_7452);
nor U7983 (N_7983,N_7198,N_7025);
and U7984 (N_7984,N_7366,N_7285);
nor U7985 (N_7985,N_7438,N_7429);
nand U7986 (N_7986,N_7498,N_7338);
or U7987 (N_7987,N_7337,N_7103);
or U7988 (N_7988,N_7443,N_7294);
or U7989 (N_7989,N_7096,N_7221);
or U7990 (N_7990,N_7453,N_7196);
xnor U7991 (N_7991,N_7051,N_7347);
xnor U7992 (N_7992,N_7349,N_7038);
nor U7993 (N_7993,N_7451,N_7106);
xnor U7994 (N_7994,N_7442,N_7105);
or U7995 (N_7995,N_7254,N_7139);
or U7996 (N_7996,N_7405,N_7087);
nor U7997 (N_7997,N_7362,N_7377);
and U7998 (N_7998,N_7364,N_7433);
xor U7999 (N_7999,N_7308,N_7038);
nor U8000 (N_8000,N_7755,N_7523);
nand U8001 (N_8001,N_7695,N_7752);
nor U8002 (N_8002,N_7834,N_7561);
nor U8003 (N_8003,N_7587,N_7871);
xor U8004 (N_8004,N_7851,N_7746);
xnor U8005 (N_8005,N_7771,N_7933);
or U8006 (N_8006,N_7715,N_7744);
nand U8007 (N_8007,N_7585,N_7685);
and U8008 (N_8008,N_7699,N_7790);
or U8009 (N_8009,N_7538,N_7892);
nand U8010 (N_8010,N_7612,N_7841);
nand U8011 (N_8011,N_7954,N_7897);
or U8012 (N_8012,N_7916,N_7516);
and U8013 (N_8013,N_7729,N_7743);
nor U8014 (N_8014,N_7658,N_7889);
nand U8015 (N_8015,N_7529,N_7815);
nor U8016 (N_8016,N_7631,N_7659);
or U8017 (N_8017,N_7964,N_7522);
nor U8018 (N_8018,N_7803,N_7642);
nand U8019 (N_8019,N_7598,N_7694);
nand U8020 (N_8020,N_7608,N_7630);
xor U8021 (N_8021,N_7848,N_7722);
nor U8022 (N_8022,N_7850,N_7976);
and U8023 (N_8023,N_7718,N_7800);
xnor U8024 (N_8024,N_7861,N_7874);
or U8025 (N_8025,N_7860,N_7619);
and U8026 (N_8026,N_7993,N_7568);
nor U8027 (N_8027,N_7886,N_7578);
or U8028 (N_8028,N_7610,N_7702);
xnor U8029 (N_8029,N_7651,N_7502);
nor U8030 (N_8030,N_7534,N_7667);
xor U8031 (N_8031,N_7939,N_7925);
nor U8032 (N_8032,N_7589,N_7931);
and U8033 (N_8033,N_7799,N_7688);
or U8034 (N_8034,N_7710,N_7643);
nand U8035 (N_8035,N_7543,N_7704);
xor U8036 (N_8036,N_7927,N_7641);
and U8037 (N_8037,N_7547,N_7508);
nand U8038 (N_8038,N_7811,N_7842);
nor U8039 (N_8039,N_7994,N_7652);
or U8040 (N_8040,N_7967,N_7614);
xnor U8041 (N_8041,N_7678,N_7726);
or U8042 (N_8042,N_7539,N_7697);
nand U8043 (N_8043,N_7930,N_7596);
and U8044 (N_8044,N_7607,N_7914);
and U8045 (N_8045,N_7648,N_7951);
or U8046 (N_8046,N_7572,N_7501);
and U8047 (N_8047,N_7582,N_7550);
nor U8048 (N_8048,N_7968,N_7580);
and U8049 (N_8049,N_7809,N_7801);
and U8050 (N_8050,N_7932,N_7858);
xnor U8051 (N_8051,N_7990,N_7626);
nand U8052 (N_8052,N_7813,N_7512);
xnor U8053 (N_8053,N_7756,N_7765);
or U8054 (N_8054,N_7884,N_7936);
nor U8055 (N_8055,N_7958,N_7613);
nor U8056 (N_8056,N_7804,N_7881);
or U8057 (N_8057,N_7785,N_7594);
xor U8058 (N_8058,N_7928,N_7778);
and U8059 (N_8059,N_7987,N_7693);
xor U8060 (N_8060,N_7513,N_7821);
xnor U8061 (N_8061,N_7818,N_7581);
xnor U8062 (N_8062,N_7888,N_7959);
xnor U8063 (N_8063,N_7797,N_7611);
nor U8064 (N_8064,N_7966,N_7773);
xnor U8065 (N_8065,N_7961,N_7989);
xnor U8066 (N_8066,N_7977,N_7946);
and U8067 (N_8067,N_7776,N_7998);
xnor U8068 (N_8068,N_7747,N_7524);
xor U8069 (N_8069,N_7810,N_7711);
or U8070 (N_8070,N_7760,N_7542);
or U8071 (N_8071,N_7759,N_7733);
xor U8072 (N_8072,N_7908,N_7527);
and U8073 (N_8073,N_7983,N_7774);
and U8074 (N_8074,N_7671,N_7792);
xnor U8075 (N_8075,N_7504,N_7978);
or U8076 (N_8076,N_7896,N_7764);
or U8077 (N_8077,N_7681,N_7979);
nand U8078 (N_8078,N_7955,N_7661);
and U8079 (N_8079,N_7570,N_7625);
xor U8080 (N_8080,N_7532,N_7721);
and U8081 (N_8081,N_7690,N_7624);
xnor U8082 (N_8082,N_7505,N_7766);
nand U8083 (N_8083,N_7736,N_7653);
or U8084 (N_8084,N_7664,N_7814);
xor U8085 (N_8085,N_7817,N_7565);
or U8086 (N_8086,N_7745,N_7638);
or U8087 (N_8087,N_7775,N_7899);
or U8088 (N_8088,N_7795,N_7960);
and U8089 (N_8089,N_7825,N_7944);
nand U8090 (N_8090,N_7541,N_7635);
or U8091 (N_8091,N_7526,N_7629);
or U8092 (N_8092,N_7820,N_7903);
nor U8093 (N_8093,N_7616,N_7838);
or U8094 (N_8094,N_7560,N_7957);
and U8095 (N_8095,N_7772,N_7969);
xor U8096 (N_8096,N_7984,N_7556);
and U8097 (N_8097,N_7684,N_7657);
xor U8098 (N_8098,N_7591,N_7862);
or U8099 (N_8099,N_7731,N_7869);
xor U8100 (N_8100,N_7844,N_7943);
or U8101 (N_8101,N_7950,N_7751);
and U8102 (N_8102,N_7615,N_7533);
nor U8103 (N_8103,N_7822,N_7605);
nor U8104 (N_8104,N_7609,N_7761);
nor U8105 (N_8105,N_7794,N_7975);
or U8106 (N_8106,N_7714,N_7637);
nand U8107 (N_8107,N_7553,N_7885);
xnor U8108 (N_8108,N_7528,N_7901);
nor U8109 (N_8109,N_7839,N_7549);
xor U8110 (N_8110,N_7974,N_7555);
nand U8111 (N_8111,N_7852,N_7518);
nor U8112 (N_8112,N_7781,N_7677);
xnor U8113 (N_8113,N_7540,N_7971);
or U8114 (N_8114,N_7823,N_7995);
and U8115 (N_8115,N_7573,N_7606);
nand U8116 (N_8116,N_7949,N_7696);
nand U8117 (N_8117,N_7701,N_7511);
xnor U8118 (N_8118,N_7798,N_7698);
xor U8119 (N_8119,N_7712,N_7856);
nand U8120 (N_8120,N_7986,N_7926);
nand U8121 (N_8121,N_7590,N_7812);
nor U8122 (N_8122,N_7520,N_7544);
xnor U8123 (N_8123,N_7758,N_7668);
nor U8124 (N_8124,N_7855,N_7519);
or U8125 (N_8125,N_7947,N_7847);
nor U8126 (N_8126,N_7551,N_7909);
and U8127 (N_8127,N_7819,N_7618);
xnor U8128 (N_8128,N_7672,N_7674);
xor U8129 (N_8129,N_7600,N_7749);
or U8130 (N_8130,N_7724,N_7827);
and U8131 (N_8131,N_7537,N_7649);
or U8132 (N_8132,N_7929,N_7833);
and U8133 (N_8133,N_7962,N_7577);
nand U8134 (N_8134,N_7628,N_7786);
xnor U8135 (N_8135,N_7576,N_7700);
xnor U8136 (N_8136,N_7571,N_7632);
nor U8137 (N_8137,N_7999,N_7675);
nand U8138 (N_8138,N_7876,N_7782);
or U8139 (N_8139,N_7557,N_7627);
nor U8140 (N_8140,N_7521,N_7934);
nor U8141 (N_8141,N_7942,N_7554);
or U8142 (N_8142,N_7603,N_7676);
nand U8143 (N_8143,N_7566,N_7866);
nand U8144 (N_8144,N_7535,N_7592);
nand U8145 (N_8145,N_7666,N_7913);
nor U8146 (N_8146,N_7757,N_7748);
nor U8147 (N_8147,N_7621,N_7753);
or U8148 (N_8148,N_7859,N_7552);
or U8149 (N_8149,N_7895,N_7679);
or U8150 (N_8150,N_7669,N_7890);
xnor U8151 (N_8151,N_7686,N_7604);
or U8152 (N_8152,N_7910,N_7660);
or U8153 (N_8153,N_7770,N_7793);
and U8154 (N_8154,N_7846,N_7644);
nor U8155 (N_8155,N_7545,N_7938);
nand U8156 (N_8156,N_7691,N_7980);
and U8157 (N_8157,N_7683,N_7739);
and U8158 (N_8158,N_7530,N_7777);
nor U8159 (N_8159,N_7740,N_7824);
and U8160 (N_8160,N_7981,N_7991);
xor U8161 (N_8161,N_7918,N_7655);
and U8162 (N_8162,N_7720,N_7564);
nor U8163 (N_8163,N_7891,N_7647);
or U8164 (N_8164,N_7662,N_7569);
nand U8165 (N_8165,N_7732,N_7921);
xor U8166 (N_8166,N_7692,N_7830);
nor U8167 (N_8167,N_7937,N_7623);
nor U8168 (N_8168,N_7920,N_7972);
or U8169 (N_8169,N_7788,N_7900);
nor U8170 (N_8170,N_7670,N_7857);
or U8171 (N_8171,N_7832,N_7507);
or U8172 (N_8172,N_7730,N_7601);
xor U8173 (N_8173,N_7878,N_7898);
and U8174 (N_8174,N_7911,N_7597);
xor U8175 (N_8175,N_7880,N_7558);
nor U8176 (N_8176,N_7919,N_7877);
and U8177 (N_8177,N_7816,N_7735);
xor U8178 (N_8178,N_7510,N_7787);
and U8179 (N_8179,N_7645,N_7883);
or U8180 (N_8180,N_7707,N_7705);
nand U8181 (N_8181,N_7650,N_7808);
nor U8182 (N_8182,N_7840,N_7574);
or U8183 (N_8183,N_7728,N_7988);
and U8184 (N_8184,N_7762,N_7789);
or U8185 (N_8185,N_7639,N_7506);
nor U8186 (N_8186,N_7515,N_7873);
and U8187 (N_8187,N_7912,N_7734);
xor U8188 (N_8188,N_7970,N_7500);
or U8189 (N_8189,N_7828,N_7907);
or U8190 (N_8190,N_7768,N_7875);
and U8191 (N_8191,N_7738,N_7716);
nand U8192 (N_8192,N_7953,N_7656);
nor U8193 (N_8193,N_7708,N_7741);
nand U8194 (N_8194,N_7536,N_7985);
nor U8195 (N_8195,N_7941,N_7867);
nand U8196 (N_8196,N_7563,N_7807);
xnor U8197 (N_8197,N_7719,N_7654);
xnor U8198 (N_8198,N_7703,N_7997);
and U8199 (N_8199,N_7870,N_7562);
nor U8200 (N_8200,N_7948,N_7905);
and U8201 (N_8201,N_7887,N_7783);
nand U8202 (N_8202,N_7879,N_7706);
or U8203 (N_8203,N_7849,N_7796);
nand U8204 (N_8204,N_7663,N_7567);
xor U8205 (N_8205,N_7665,N_7593);
and U8206 (N_8206,N_7868,N_7713);
or U8207 (N_8207,N_7791,N_7617);
xor U8208 (N_8208,N_7682,N_7586);
nand U8209 (N_8209,N_7853,N_7935);
or U8210 (N_8210,N_7805,N_7784);
and U8211 (N_8211,N_7843,N_7525);
nand U8212 (N_8212,N_7917,N_7992);
xnor U8213 (N_8213,N_7906,N_7963);
and U8214 (N_8214,N_7845,N_7717);
or U8215 (N_8215,N_7894,N_7575);
xnor U8216 (N_8216,N_7872,N_7882);
nand U8217 (N_8217,N_7514,N_7588);
nor U8218 (N_8218,N_7973,N_7952);
or U8219 (N_8219,N_7826,N_7620);
nor U8220 (N_8220,N_7584,N_7965);
nand U8221 (N_8221,N_7503,N_7854);
nor U8222 (N_8222,N_7689,N_7633);
nor U8223 (N_8223,N_7559,N_7646);
and U8224 (N_8224,N_7673,N_7831);
or U8225 (N_8225,N_7982,N_7864);
nor U8226 (N_8226,N_7767,N_7802);
nand U8227 (N_8227,N_7915,N_7835);
nor U8228 (N_8228,N_7750,N_7602);
nor U8229 (N_8229,N_7924,N_7517);
nand U8230 (N_8230,N_7531,N_7622);
xnor U8231 (N_8231,N_7709,N_7595);
nor U8232 (N_8232,N_7829,N_7680);
and U8233 (N_8233,N_7737,N_7687);
xor U8234 (N_8234,N_7996,N_7904);
nor U8235 (N_8235,N_7863,N_7902);
xnor U8236 (N_8236,N_7754,N_7780);
xnor U8237 (N_8237,N_7865,N_7742);
xnor U8238 (N_8238,N_7945,N_7763);
xnor U8239 (N_8239,N_7806,N_7599);
and U8240 (N_8240,N_7727,N_7636);
xnor U8241 (N_8241,N_7548,N_7640);
xor U8242 (N_8242,N_7837,N_7723);
or U8243 (N_8243,N_7509,N_7769);
nand U8244 (N_8244,N_7923,N_7922);
nand U8245 (N_8245,N_7634,N_7583);
xnor U8246 (N_8246,N_7579,N_7725);
and U8247 (N_8247,N_7956,N_7546);
nor U8248 (N_8248,N_7779,N_7836);
nor U8249 (N_8249,N_7893,N_7940);
nand U8250 (N_8250,N_7665,N_7991);
xnor U8251 (N_8251,N_7767,N_7745);
or U8252 (N_8252,N_7500,N_7702);
or U8253 (N_8253,N_7883,N_7902);
xor U8254 (N_8254,N_7635,N_7945);
nor U8255 (N_8255,N_7912,N_7659);
and U8256 (N_8256,N_7804,N_7648);
nand U8257 (N_8257,N_7717,N_7874);
xnor U8258 (N_8258,N_7739,N_7686);
or U8259 (N_8259,N_7775,N_7526);
or U8260 (N_8260,N_7685,N_7692);
nor U8261 (N_8261,N_7554,N_7849);
xnor U8262 (N_8262,N_7954,N_7947);
and U8263 (N_8263,N_7662,N_7526);
or U8264 (N_8264,N_7581,N_7555);
and U8265 (N_8265,N_7960,N_7961);
nand U8266 (N_8266,N_7696,N_7507);
or U8267 (N_8267,N_7763,N_7837);
xor U8268 (N_8268,N_7502,N_7983);
and U8269 (N_8269,N_7636,N_7743);
and U8270 (N_8270,N_7830,N_7725);
nand U8271 (N_8271,N_7813,N_7627);
nor U8272 (N_8272,N_7884,N_7580);
and U8273 (N_8273,N_7975,N_7633);
xor U8274 (N_8274,N_7850,N_7893);
xor U8275 (N_8275,N_7526,N_7561);
xor U8276 (N_8276,N_7933,N_7874);
or U8277 (N_8277,N_7563,N_7822);
and U8278 (N_8278,N_7619,N_7799);
nor U8279 (N_8279,N_7907,N_7756);
xor U8280 (N_8280,N_7703,N_7518);
or U8281 (N_8281,N_7565,N_7824);
or U8282 (N_8282,N_7632,N_7862);
nand U8283 (N_8283,N_7697,N_7658);
nand U8284 (N_8284,N_7922,N_7958);
and U8285 (N_8285,N_7847,N_7568);
and U8286 (N_8286,N_7655,N_7721);
nand U8287 (N_8287,N_7672,N_7619);
or U8288 (N_8288,N_7521,N_7847);
nor U8289 (N_8289,N_7799,N_7901);
and U8290 (N_8290,N_7866,N_7827);
and U8291 (N_8291,N_7975,N_7965);
xnor U8292 (N_8292,N_7940,N_7916);
nor U8293 (N_8293,N_7978,N_7812);
nand U8294 (N_8294,N_7869,N_7738);
xnor U8295 (N_8295,N_7804,N_7749);
and U8296 (N_8296,N_7897,N_7560);
nor U8297 (N_8297,N_7656,N_7856);
nand U8298 (N_8298,N_7665,N_7619);
or U8299 (N_8299,N_7649,N_7830);
nand U8300 (N_8300,N_7627,N_7963);
nand U8301 (N_8301,N_7777,N_7997);
or U8302 (N_8302,N_7974,N_7817);
xor U8303 (N_8303,N_7746,N_7932);
xnor U8304 (N_8304,N_7564,N_7760);
and U8305 (N_8305,N_7540,N_7748);
nor U8306 (N_8306,N_7763,N_7894);
or U8307 (N_8307,N_7824,N_7628);
and U8308 (N_8308,N_7875,N_7727);
xnor U8309 (N_8309,N_7675,N_7726);
and U8310 (N_8310,N_7756,N_7768);
nand U8311 (N_8311,N_7878,N_7896);
xor U8312 (N_8312,N_7755,N_7605);
xor U8313 (N_8313,N_7720,N_7968);
or U8314 (N_8314,N_7784,N_7609);
nor U8315 (N_8315,N_7679,N_7598);
and U8316 (N_8316,N_7787,N_7676);
nand U8317 (N_8317,N_7595,N_7664);
xor U8318 (N_8318,N_7553,N_7878);
nor U8319 (N_8319,N_7816,N_7663);
xor U8320 (N_8320,N_7565,N_7811);
or U8321 (N_8321,N_7937,N_7907);
nor U8322 (N_8322,N_7567,N_7714);
xor U8323 (N_8323,N_7645,N_7865);
and U8324 (N_8324,N_7543,N_7738);
xnor U8325 (N_8325,N_7759,N_7548);
xnor U8326 (N_8326,N_7740,N_7880);
and U8327 (N_8327,N_7870,N_7677);
or U8328 (N_8328,N_7926,N_7579);
xnor U8329 (N_8329,N_7966,N_7829);
or U8330 (N_8330,N_7831,N_7783);
and U8331 (N_8331,N_7527,N_7582);
or U8332 (N_8332,N_7852,N_7740);
nand U8333 (N_8333,N_7692,N_7826);
xnor U8334 (N_8334,N_7938,N_7836);
xor U8335 (N_8335,N_7772,N_7866);
nor U8336 (N_8336,N_7904,N_7760);
or U8337 (N_8337,N_7725,N_7508);
or U8338 (N_8338,N_7763,N_7898);
nand U8339 (N_8339,N_7836,N_7586);
xnor U8340 (N_8340,N_7683,N_7501);
xnor U8341 (N_8341,N_7611,N_7631);
nor U8342 (N_8342,N_7987,N_7721);
nand U8343 (N_8343,N_7550,N_7579);
nor U8344 (N_8344,N_7645,N_7542);
and U8345 (N_8345,N_7974,N_7759);
nor U8346 (N_8346,N_7639,N_7977);
xnor U8347 (N_8347,N_7796,N_7606);
nor U8348 (N_8348,N_7623,N_7658);
nand U8349 (N_8349,N_7734,N_7886);
or U8350 (N_8350,N_7588,N_7916);
nor U8351 (N_8351,N_7803,N_7729);
xor U8352 (N_8352,N_7614,N_7847);
xnor U8353 (N_8353,N_7772,N_7570);
and U8354 (N_8354,N_7838,N_7721);
nand U8355 (N_8355,N_7555,N_7506);
or U8356 (N_8356,N_7503,N_7707);
nand U8357 (N_8357,N_7780,N_7949);
nand U8358 (N_8358,N_7667,N_7573);
nand U8359 (N_8359,N_7881,N_7606);
and U8360 (N_8360,N_7772,N_7945);
nor U8361 (N_8361,N_7984,N_7645);
nor U8362 (N_8362,N_7933,N_7948);
or U8363 (N_8363,N_7975,N_7686);
and U8364 (N_8364,N_7782,N_7705);
and U8365 (N_8365,N_7581,N_7569);
nor U8366 (N_8366,N_7934,N_7694);
nor U8367 (N_8367,N_7938,N_7802);
nor U8368 (N_8368,N_7920,N_7591);
nor U8369 (N_8369,N_7726,N_7610);
xnor U8370 (N_8370,N_7819,N_7722);
nor U8371 (N_8371,N_7973,N_7536);
nand U8372 (N_8372,N_7569,N_7758);
xor U8373 (N_8373,N_7622,N_7956);
xnor U8374 (N_8374,N_7987,N_7545);
and U8375 (N_8375,N_7752,N_7852);
nand U8376 (N_8376,N_7726,N_7887);
or U8377 (N_8377,N_7915,N_7723);
nor U8378 (N_8378,N_7920,N_7907);
xor U8379 (N_8379,N_7872,N_7601);
and U8380 (N_8380,N_7659,N_7909);
and U8381 (N_8381,N_7741,N_7558);
xor U8382 (N_8382,N_7759,N_7725);
nor U8383 (N_8383,N_7501,N_7999);
or U8384 (N_8384,N_7519,N_7726);
nand U8385 (N_8385,N_7734,N_7924);
and U8386 (N_8386,N_7541,N_7971);
or U8387 (N_8387,N_7643,N_7995);
and U8388 (N_8388,N_7674,N_7627);
nand U8389 (N_8389,N_7989,N_7553);
nor U8390 (N_8390,N_7624,N_7655);
xnor U8391 (N_8391,N_7860,N_7989);
and U8392 (N_8392,N_7853,N_7934);
xnor U8393 (N_8393,N_7941,N_7685);
xor U8394 (N_8394,N_7668,N_7905);
or U8395 (N_8395,N_7613,N_7984);
and U8396 (N_8396,N_7640,N_7633);
or U8397 (N_8397,N_7893,N_7660);
and U8398 (N_8398,N_7728,N_7640);
xor U8399 (N_8399,N_7665,N_7517);
nand U8400 (N_8400,N_7602,N_7713);
or U8401 (N_8401,N_7922,N_7514);
nor U8402 (N_8402,N_7551,N_7630);
nor U8403 (N_8403,N_7794,N_7789);
nor U8404 (N_8404,N_7632,N_7537);
or U8405 (N_8405,N_7689,N_7897);
xnor U8406 (N_8406,N_7839,N_7941);
xnor U8407 (N_8407,N_7981,N_7587);
xor U8408 (N_8408,N_7945,N_7877);
nor U8409 (N_8409,N_7646,N_7769);
nand U8410 (N_8410,N_7880,N_7613);
and U8411 (N_8411,N_7977,N_7984);
xor U8412 (N_8412,N_7877,N_7567);
and U8413 (N_8413,N_7613,N_7826);
xor U8414 (N_8414,N_7898,N_7537);
or U8415 (N_8415,N_7935,N_7816);
nor U8416 (N_8416,N_7774,N_7908);
or U8417 (N_8417,N_7924,N_7728);
nor U8418 (N_8418,N_7789,N_7746);
xnor U8419 (N_8419,N_7839,N_7693);
nand U8420 (N_8420,N_7587,N_7798);
and U8421 (N_8421,N_7744,N_7986);
nand U8422 (N_8422,N_7839,N_7621);
and U8423 (N_8423,N_7870,N_7952);
xor U8424 (N_8424,N_7696,N_7750);
and U8425 (N_8425,N_7906,N_7726);
nand U8426 (N_8426,N_7728,N_7669);
xor U8427 (N_8427,N_7879,N_7655);
or U8428 (N_8428,N_7618,N_7770);
and U8429 (N_8429,N_7726,N_7776);
or U8430 (N_8430,N_7909,N_7574);
and U8431 (N_8431,N_7685,N_7990);
xor U8432 (N_8432,N_7913,N_7880);
xor U8433 (N_8433,N_7969,N_7608);
nor U8434 (N_8434,N_7661,N_7974);
nand U8435 (N_8435,N_7846,N_7913);
nor U8436 (N_8436,N_7551,N_7900);
xnor U8437 (N_8437,N_7552,N_7875);
nor U8438 (N_8438,N_7760,N_7861);
xnor U8439 (N_8439,N_7518,N_7955);
or U8440 (N_8440,N_7703,N_7972);
and U8441 (N_8441,N_7889,N_7870);
nand U8442 (N_8442,N_7827,N_7834);
or U8443 (N_8443,N_7592,N_7625);
and U8444 (N_8444,N_7780,N_7619);
nor U8445 (N_8445,N_7927,N_7885);
nand U8446 (N_8446,N_7738,N_7878);
xor U8447 (N_8447,N_7737,N_7515);
and U8448 (N_8448,N_7609,N_7899);
or U8449 (N_8449,N_7952,N_7889);
xnor U8450 (N_8450,N_7831,N_7734);
nor U8451 (N_8451,N_7893,N_7713);
nor U8452 (N_8452,N_7800,N_7882);
and U8453 (N_8453,N_7752,N_7995);
xnor U8454 (N_8454,N_7725,N_7766);
nor U8455 (N_8455,N_7603,N_7692);
nor U8456 (N_8456,N_7847,N_7618);
or U8457 (N_8457,N_7833,N_7529);
nand U8458 (N_8458,N_7750,N_7894);
nand U8459 (N_8459,N_7668,N_7943);
nand U8460 (N_8460,N_7588,N_7819);
and U8461 (N_8461,N_7795,N_7993);
xor U8462 (N_8462,N_7998,N_7783);
nand U8463 (N_8463,N_7795,N_7598);
xor U8464 (N_8464,N_7728,N_7778);
xnor U8465 (N_8465,N_7916,N_7994);
nor U8466 (N_8466,N_7925,N_7610);
xnor U8467 (N_8467,N_7593,N_7536);
nand U8468 (N_8468,N_7552,N_7502);
or U8469 (N_8469,N_7777,N_7834);
nand U8470 (N_8470,N_7916,N_7625);
or U8471 (N_8471,N_7610,N_7753);
nand U8472 (N_8472,N_7803,N_7837);
nand U8473 (N_8473,N_7882,N_7829);
and U8474 (N_8474,N_7699,N_7994);
and U8475 (N_8475,N_7760,N_7621);
or U8476 (N_8476,N_7763,N_7579);
or U8477 (N_8477,N_7792,N_7961);
xor U8478 (N_8478,N_7952,N_7800);
or U8479 (N_8479,N_7969,N_7749);
or U8480 (N_8480,N_7668,N_7723);
nor U8481 (N_8481,N_7545,N_7788);
nand U8482 (N_8482,N_7953,N_7721);
and U8483 (N_8483,N_7645,N_7719);
and U8484 (N_8484,N_7640,N_7564);
xnor U8485 (N_8485,N_7681,N_7799);
xnor U8486 (N_8486,N_7624,N_7766);
nand U8487 (N_8487,N_7590,N_7762);
and U8488 (N_8488,N_7882,N_7659);
and U8489 (N_8489,N_7756,N_7673);
and U8490 (N_8490,N_7574,N_7665);
or U8491 (N_8491,N_7825,N_7518);
nand U8492 (N_8492,N_7906,N_7575);
and U8493 (N_8493,N_7828,N_7810);
or U8494 (N_8494,N_7695,N_7753);
nand U8495 (N_8495,N_7902,N_7846);
nand U8496 (N_8496,N_7793,N_7775);
xor U8497 (N_8497,N_7548,N_7922);
xor U8498 (N_8498,N_7573,N_7815);
and U8499 (N_8499,N_7600,N_7905);
or U8500 (N_8500,N_8090,N_8172);
nand U8501 (N_8501,N_8005,N_8118);
nand U8502 (N_8502,N_8196,N_8021);
nand U8503 (N_8503,N_8470,N_8405);
nand U8504 (N_8504,N_8261,N_8302);
nand U8505 (N_8505,N_8378,N_8154);
nor U8506 (N_8506,N_8436,N_8145);
and U8507 (N_8507,N_8432,N_8173);
and U8508 (N_8508,N_8252,N_8075);
and U8509 (N_8509,N_8494,N_8319);
nor U8510 (N_8510,N_8217,N_8002);
and U8511 (N_8511,N_8025,N_8257);
nand U8512 (N_8512,N_8422,N_8143);
nand U8513 (N_8513,N_8496,N_8469);
nand U8514 (N_8514,N_8442,N_8138);
nor U8515 (N_8515,N_8310,N_8419);
nor U8516 (N_8516,N_8408,N_8165);
xor U8517 (N_8517,N_8328,N_8079);
and U8518 (N_8518,N_8158,N_8339);
nor U8519 (N_8519,N_8170,N_8398);
xnor U8520 (N_8520,N_8092,N_8293);
xnor U8521 (N_8521,N_8239,N_8355);
or U8522 (N_8522,N_8268,N_8135);
nand U8523 (N_8523,N_8406,N_8198);
nor U8524 (N_8524,N_8255,N_8142);
nand U8525 (N_8525,N_8070,N_8280);
and U8526 (N_8526,N_8010,N_8474);
and U8527 (N_8527,N_8253,N_8227);
xor U8528 (N_8528,N_8472,N_8338);
xnor U8529 (N_8529,N_8367,N_8159);
and U8530 (N_8530,N_8362,N_8059);
or U8531 (N_8531,N_8213,N_8073);
nand U8532 (N_8532,N_8490,N_8038);
nor U8533 (N_8533,N_8134,N_8177);
or U8534 (N_8534,N_8153,N_8131);
nand U8535 (N_8535,N_8308,N_8036);
xor U8536 (N_8536,N_8449,N_8195);
and U8537 (N_8537,N_8381,N_8263);
and U8538 (N_8538,N_8150,N_8063);
xor U8539 (N_8539,N_8477,N_8218);
nand U8540 (N_8540,N_8467,N_8087);
nand U8541 (N_8541,N_8215,N_8459);
or U8542 (N_8542,N_8137,N_8330);
or U8543 (N_8543,N_8337,N_8234);
xnor U8544 (N_8544,N_8363,N_8298);
or U8545 (N_8545,N_8418,N_8274);
nand U8546 (N_8546,N_8169,N_8123);
and U8547 (N_8547,N_8081,N_8240);
or U8548 (N_8548,N_8389,N_8236);
or U8549 (N_8549,N_8178,N_8219);
and U8550 (N_8550,N_8006,N_8383);
nor U8551 (N_8551,N_8311,N_8284);
and U8552 (N_8552,N_8190,N_8281);
nor U8553 (N_8553,N_8214,N_8283);
nand U8554 (N_8554,N_8035,N_8113);
and U8555 (N_8555,N_8409,N_8428);
nor U8556 (N_8556,N_8372,N_8313);
nor U8557 (N_8557,N_8163,N_8478);
nor U8558 (N_8558,N_8421,N_8392);
nor U8559 (N_8559,N_8466,N_8486);
or U8560 (N_8560,N_8033,N_8034);
xor U8561 (N_8561,N_8146,N_8055);
nand U8562 (N_8562,N_8402,N_8208);
xnor U8563 (N_8563,N_8191,N_8031);
and U8564 (N_8564,N_8384,N_8228);
and U8565 (N_8565,N_8209,N_8288);
nor U8566 (N_8566,N_8220,N_8291);
and U8567 (N_8567,N_8399,N_8183);
xor U8568 (N_8568,N_8053,N_8394);
and U8569 (N_8569,N_8229,N_8451);
nor U8570 (N_8570,N_8426,N_8304);
nor U8571 (N_8571,N_8047,N_8111);
xor U8572 (N_8572,N_8060,N_8414);
xor U8573 (N_8573,N_8011,N_8185);
nand U8574 (N_8574,N_8433,N_8050);
and U8575 (N_8575,N_8270,N_8062);
or U8576 (N_8576,N_8357,N_8175);
nand U8577 (N_8577,N_8093,N_8224);
nand U8578 (N_8578,N_8144,N_8462);
or U8579 (N_8579,N_8015,N_8151);
and U8580 (N_8580,N_8120,N_8251);
xor U8581 (N_8581,N_8121,N_8187);
and U8582 (N_8582,N_8373,N_8119);
or U8583 (N_8583,N_8309,N_8277);
nand U8584 (N_8584,N_8285,N_8094);
or U8585 (N_8585,N_8267,N_8057);
and U8586 (N_8586,N_8431,N_8312);
xor U8587 (N_8587,N_8456,N_8305);
and U8588 (N_8588,N_8371,N_8122);
and U8589 (N_8589,N_8030,N_8226);
xor U8590 (N_8590,N_8260,N_8282);
nand U8591 (N_8591,N_8171,N_8333);
xor U8592 (N_8592,N_8325,N_8349);
nand U8593 (N_8593,N_8231,N_8071);
xor U8594 (N_8594,N_8056,N_8427);
nor U8595 (N_8595,N_8259,N_8105);
nor U8596 (N_8596,N_8447,N_8415);
nor U8597 (N_8597,N_8039,N_8463);
and U8598 (N_8598,N_8242,N_8160);
and U8599 (N_8599,N_8300,N_8279);
xor U8600 (N_8600,N_8335,N_8243);
xnor U8601 (N_8601,N_8124,N_8222);
xor U8602 (N_8602,N_8434,N_8126);
or U8603 (N_8603,N_8018,N_8082);
nor U8604 (N_8604,N_8179,N_8404);
xnor U8605 (N_8605,N_8497,N_8495);
nor U8606 (N_8606,N_8321,N_8139);
or U8607 (N_8607,N_8230,N_8080);
or U8608 (N_8608,N_8382,N_8106);
or U8609 (N_8609,N_8471,N_8186);
nor U8610 (N_8610,N_8238,N_8387);
nand U8611 (N_8611,N_8391,N_8200);
nand U8612 (N_8612,N_8483,N_8117);
and U8613 (N_8613,N_8316,N_8354);
and U8614 (N_8614,N_8072,N_8343);
xnor U8615 (N_8615,N_8232,N_8003);
xor U8616 (N_8616,N_8443,N_8019);
and U8617 (N_8617,N_8029,N_8104);
and U8618 (N_8618,N_8395,N_8058);
or U8619 (N_8619,N_8249,N_8350);
and U8620 (N_8620,N_8344,N_8484);
and U8621 (N_8621,N_8364,N_8237);
xor U8622 (N_8622,N_8379,N_8192);
and U8623 (N_8623,N_8370,N_8199);
or U8624 (N_8624,N_8247,N_8439);
xnor U8625 (N_8625,N_8413,N_8101);
or U8626 (N_8626,N_8017,N_8425);
or U8627 (N_8627,N_8109,N_8098);
and U8628 (N_8628,N_8448,N_8468);
or U8629 (N_8629,N_8008,N_8386);
or U8630 (N_8630,N_8007,N_8041);
xor U8631 (N_8631,N_8161,N_8390);
and U8632 (N_8632,N_8128,N_8489);
and U8633 (N_8633,N_8303,N_8326);
nor U8634 (N_8634,N_8223,N_8435);
nor U8635 (N_8635,N_8216,N_8086);
and U8636 (N_8636,N_8482,N_8046);
and U8637 (N_8637,N_8174,N_8444);
and U8638 (N_8638,N_8180,N_8042);
and U8639 (N_8639,N_8088,N_8317);
nor U8640 (N_8640,N_8149,N_8084);
and U8641 (N_8641,N_8287,N_8068);
nor U8642 (N_8642,N_8385,N_8301);
nor U8643 (N_8643,N_8076,N_8193);
or U8644 (N_8644,N_8182,N_8125);
or U8645 (N_8645,N_8417,N_8012);
nand U8646 (N_8646,N_8108,N_8194);
and U8647 (N_8647,N_8212,N_8157);
and U8648 (N_8648,N_8491,N_8412);
xnor U8649 (N_8649,N_8396,N_8167);
and U8650 (N_8650,N_8393,N_8152);
nor U8651 (N_8651,N_8318,N_8295);
and U8652 (N_8652,N_8256,N_8254);
or U8653 (N_8653,N_8248,N_8027);
nand U8654 (N_8654,N_8074,N_8410);
and U8655 (N_8655,N_8001,N_8473);
nor U8656 (N_8656,N_8233,N_8361);
nand U8657 (N_8657,N_8114,N_8376);
or U8658 (N_8658,N_8156,N_8351);
xor U8659 (N_8659,N_8023,N_8380);
xnor U8660 (N_8660,N_8347,N_8440);
and U8661 (N_8661,N_8329,N_8014);
nand U8662 (N_8662,N_8374,N_8264);
xnor U8663 (N_8663,N_8272,N_8365);
nand U8664 (N_8664,N_8102,N_8097);
and U8665 (N_8665,N_8162,N_8481);
and U8666 (N_8666,N_8258,N_8375);
xor U8667 (N_8667,N_8132,N_8327);
or U8668 (N_8668,N_8437,N_8420);
and U8669 (N_8669,N_8429,N_8441);
and U8670 (N_8670,N_8341,N_8176);
nand U8671 (N_8671,N_8089,N_8324);
and U8672 (N_8672,N_8269,N_8052);
or U8673 (N_8673,N_8278,N_8368);
xnor U8674 (N_8674,N_8452,N_8078);
or U8675 (N_8675,N_8026,N_8077);
or U8676 (N_8676,N_8028,N_8207);
xnor U8677 (N_8677,N_8266,N_8352);
xnor U8678 (N_8678,N_8290,N_8377);
nand U8679 (N_8679,N_8356,N_8403);
nand U8680 (N_8680,N_8022,N_8453);
nand U8681 (N_8681,N_8485,N_8292);
nor U8682 (N_8682,N_8276,N_8099);
xnor U8683 (N_8683,N_8184,N_8205);
or U8684 (N_8684,N_8069,N_8043);
or U8685 (N_8685,N_8457,N_8211);
nand U8686 (N_8686,N_8155,N_8455);
and U8687 (N_8687,N_8320,N_8342);
nand U8688 (N_8688,N_8446,N_8112);
nor U8689 (N_8689,N_8107,N_8140);
and U8690 (N_8690,N_8438,N_8476);
nand U8691 (N_8691,N_8133,N_8488);
and U8692 (N_8692,N_8464,N_8009);
nor U8693 (N_8693,N_8265,N_8130);
nor U8694 (N_8694,N_8366,N_8083);
nor U8695 (N_8695,N_8091,N_8400);
nand U8696 (N_8696,N_8294,N_8407);
and U8697 (N_8697,N_8299,N_8044);
and U8698 (N_8698,N_8061,N_8181);
or U8699 (N_8699,N_8246,N_8332);
or U8700 (N_8700,N_8315,N_8066);
or U8701 (N_8701,N_8450,N_8024);
nand U8702 (N_8702,N_8067,N_8037);
or U8703 (N_8703,N_8336,N_8168);
xnor U8704 (N_8704,N_8100,N_8314);
xor U8705 (N_8705,N_8323,N_8250);
nor U8706 (N_8706,N_8095,N_8388);
and U8707 (N_8707,N_8141,N_8460);
or U8708 (N_8708,N_8454,N_8235);
nor U8709 (N_8709,N_8210,N_8147);
nor U8710 (N_8710,N_8116,N_8480);
xor U8711 (N_8711,N_8397,N_8166);
xnor U8712 (N_8712,N_8051,N_8423);
nor U8713 (N_8713,N_8129,N_8334);
xnor U8714 (N_8714,N_8085,N_8359);
or U8715 (N_8715,N_8475,N_8498);
or U8716 (N_8716,N_8241,N_8103);
nor U8717 (N_8717,N_8458,N_8164);
or U8718 (N_8718,N_8189,N_8348);
and U8719 (N_8719,N_8040,N_8204);
nor U8720 (N_8720,N_8045,N_8271);
and U8721 (N_8721,N_8273,N_8244);
xnor U8722 (N_8722,N_8020,N_8297);
or U8723 (N_8723,N_8358,N_8401);
or U8724 (N_8724,N_8096,N_8322);
nor U8725 (N_8725,N_8346,N_8445);
and U8726 (N_8726,N_8127,N_8000);
nand U8727 (N_8727,N_8340,N_8360);
xor U8728 (N_8728,N_8197,N_8487);
nor U8729 (N_8729,N_8245,N_8499);
and U8730 (N_8730,N_8203,N_8064);
and U8731 (N_8731,N_8289,N_8188);
nand U8732 (N_8732,N_8206,N_8411);
nand U8733 (N_8733,N_8221,N_8430);
nor U8734 (N_8734,N_8492,N_8369);
nand U8735 (N_8735,N_8013,N_8353);
and U8736 (N_8736,N_8065,N_8286);
and U8737 (N_8737,N_8296,N_8110);
nor U8738 (N_8738,N_8465,N_8416);
or U8739 (N_8739,N_8262,N_8424);
nor U8740 (N_8740,N_8201,N_8054);
nor U8741 (N_8741,N_8461,N_8136);
nand U8742 (N_8742,N_8016,N_8049);
nand U8743 (N_8743,N_8331,N_8275);
xor U8744 (N_8744,N_8493,N_8479);
xnor U8745 (N_8745,N_8115,N_8048);
xor U8746 (N_8746,N_8307,N_8345);
nor U8747 (N_8747,N_8148,N_8306);
and U8748 (N_8748,N_8032,N_8004);
and U8749 (N_8749,N_8225,N_8202);
nand U8750 (N_8750,N_8241,N_8164);
nor U8751 (N_8751,N_8116,N_8005);
and U8752 (N_8752,N_8097,N_8082);
or U8753 (N_8753,N_8499,N_8138);
nand U8754 (N_8754,N_8388,N_8324);
xor U8755 (N_8755,N_8402,N_8410);
or U8756 (N_8756,N_8162,N_8380);
or U8757 (N_8757,N_8188,N_8153);
nor U8758 (N_8758,N_8467,N_8335);
and U8759 (N_8759,N_8398,N_8465);
and U8760 (N_8760,N_8419,N_8071);
nor U8761 (N_8761,N_8195,N_8396);
nor U8762 (N_8762,N_8034,N_8060);
nor U8763 (N_8763,N_8151,N_8309);
nor U8764 (N_8764,N_8229,N_8467);
nand U8765 (N_8765,N_8489,N_8486);
nor U8766 (N_8766,N_8332,N_8354);
nor U8767 (N_8767,N_8380,N_8155);
nor U8768 (N_8768,N_8217,N_8346);
xor U8769 (N_8769,N_8468,N_8415);
xor U8770 (N_8770,N_8037,N_8147);
or U8771 (N_8771,N_8128,N_8136);
nor U8772 (N_8772,N_8281,N_8223);
and U8773 (N_8773,N_8109,N_8155);
nand U8774 (N_8774,N_8276,N_8426);
nor U8775 (N_8775,N_8202,N_8331);
and U8776 (N_8776,N_8039,N_8217);
nor U8777 (N_8777,N_8045,N_8343);
nor U8778 (N_8778,N_8107,N_8287);
or U8779 (N_8779,N_8098,N_8112);
or U8780 (N_8780,N_8226,N_8198);
and U8781 (N_8781,N_8006,N_8426);
and U8782 (N_8782,N_8102,N_8308);
and U8783 (N_8783,N_8382,N_8129);
nand U8784 (N_8784,N_8426,N_8383);
nor U8785 (N_8785,N_8466,N_8338);
xor U8786 (N_8786,N_8032,N_8158);
nand U8787 (N_8787,N_8062,N_8242);
and U8788 (N_8788,N_8200,N_8463);
nand U8789 (N_8789,N_8174,N_8004);
nand U8790 (N_8790,N_8088,N_8008);
xor U8791 (N_8791,N_8435,N_8351);
or U8792 (N_8792,N_8117,N_8237);
xnor U8793 (N_8793,N_8065,N_8318);
and U8794 (N_8794,N_8369,N_8128);
xor U8795 (N_8795,N_8198,N_8047);
and U8796 (N_8796,N_8120,N_8157);
xnor U8797 (N_8797,N_8330,N_8100);
and U8798 (N_8798,N_8267,N_8124);
xnor U8799 (N_8799,N_8017,N_8441);
nand U8800 (N_8800,N_8311,N_8156);
nor U8801 (N_8801,N_8202,N_8055);
nand U8802 (N_8802,N_8309,N_8049);
and U8803 (N_8803,N_8425,N_8009);
nand U8804 (N_8804,N_8248,N_8029);
or U8805 (N_8805,N_8398,N_8337);
nand U8806 (N_8806,N_8037,N_8476);
or U8807 (N_8807,N_8117,N_8297);
and U8808 (N_8808,N_8392,N_8045);
xor U8809 (N_8809,N_8265,N_8258);
nand U8810 (N_8810,N_8317,N_8263);
nand U8811 (N_8811,N_8053,N_8319);
xor U8812 (N_8812,N_8093,N_8011);
or U8813 (N_8813,N_8205,N_8006);
nand U8814 (N_8814,N_8450,N_8094);
and U8815 (N_8815,N_8006,N_8318);
nand U8816 (N_8816,N_8232,N_8412);
nand U8817 (N_8817,N_8083,N_8220);
nand U8818 (N_8818,N_8257,N_8485);
nor U8819 (N_8819,N_8460,N_8458);
and U8820 (N_8820,N_8013,N_8020);
nand U8821 (N_8821,N_8190,N_8299);
xnor U8822 (N_8822,N_8257,N_8171);
nand U8823 (N_8823,N_8145,N_8238);
xnor U8824 (N_8824,N_8411,N_8249);
and U8825 (N_8825,N_8331,N_8362);
xnor U8826 (N_8826,N_8030,N_8467);
and U8827 (N_8827,N_8165,N_8208);
xor U8828 (N_8828,N_8334,N_8499);
xor U8829 (N_8829,N_8470,N_8232);
and U8830 (N_8830,N_8246,N_8221);
nor U8831 (N_8831,N_8244,N_8176);
nand U8832 (N_8832,N_8150,N_8378);
and U8833 (N_8833,N_8096,N_8418);
nor U8834 (N_8834,N_8276,N_8302);
or U8835 (N_8835,N_8146,N_8250);
or U8836 (N_8836,N_8375,N_8002);
nor U8837 (N_8837,N_8086,N_8010);
or U8838 (N_8838,N_8180,N_8333);
xor U8839 (N_8839,N_8205,N_8016);
nand U8840 (N_8840,N_8371,N_8111);
nor U8841 (N_8841,N_8174,N_8136);
xnor U8842 (N_8842,N_8313,N_8016);
nand U8843 (N_8843,N_8261,N_8368);
nand U8844 (N_8844,N_8087,N_8453);
xnor U8845 (N_8845,N_8416,N_8498);
and U8846 (N_8846,N_8243,N_8190);
nor U8847 (N_8847,N_8490,N_8190);
and U8848 (N_8848,N_8006,N_8480);
xnor U8849 (N_8849,N_8037,N_8259);
or U8850 (N_8850,N_8283,N_8303);
nand U8851 (N_8851,N_8349,N_8002);
or U8852 (N_8852,N_8256,N_8113);
or U8853 (N_8853,N_8121,N_8267);
or U8854 (N_8854,N_8309,N_8160);
xor U8855 (N_8855,N_8039,N_8444);
or U8856 (N_8856,N_8346,N_8240);
nand U8857 (N_8857,N_8315,N_8086);
nand U8858 (N_8858,N_8238,N_8071);
nand U8859 (N_8859,N_8064,N_8209);
or U8860 (N_8860,N_8005,N_8071);
or U8861 (N_8861,N_8071,N_8178);
or U8862 (N_8862,N_8306,N_8105);
and U8863 (N_8863,N_8488,N_8057);
nor U8864 (N_8864,N_8056,N_8446);
nand U8865 (N_8865,N_8177,N_8222);
and U8866 (N_8866,N_8067,N_8358);
or U8867 (N_8867,N_8047,N_8362);
and U8868 (N_8868,N_8109,N_8396);
xnor U8869 (N_8869,N_8001,N_8295);
nand U8870 (N_8870,N_8257,N_8292);
xor U8871 (N_8871,N_8429,N_8110);
and U8872 (N_8872,N_8113,N_8107);
xor U8873 (N_8873,N_8001,N_8172);
and U8874 (N_8874,N_8023,N_8393);
xor U8875 (N_8875,N_8484,N_8399);
nand U8876 (N_8876,N_8106,N_8295);
nand U8877 (N_8877,N_8411,N_8194);
and U8878 (N_8878,N_8487,N_8104);
nand U8879 (N_8879,N_8155,N_8369);
nand U8880 (N_8880,N_8094,N_8308);
nor U8881 (N_8881,N_8324,N_8408);
and U8882 (N_8882,N_8439,N_8069);
and U8883 (N_8883,N_8316,N_8060);
and U8884 (N_8884,N_8496,N_8144);
nand U8885 (N_8885,N_8137,N_8172);
and U8886 (N_8886,N_8195,N_8143);
or U8887 (N_8887,N_8342,N_8000);
and U8888 (N_8888,N_8359,N_8391);
nand U8889 (N_8889,N_8009,N_8042);
nand U8890 (N_8890,N_8338,N_8256);
or U8891 (N_8891,N_8224,N_8161);
or U8892 (N_8892,N_8229,N_8202);
xor U8893 (N_8893,N_8170,N_8091);
nor U8894 (N_8894,N_8112,N_8001);
nor U8895 (N_8895,N_8192,N_8213);
and U8896 (N_8896,N_8029,N_8187);
nand U8897 (N_8897,N_8326,N_8319);
nand U8898 (N_8898,N_8386,N_8233);
nand U8899 (N_8899,N_8454,N_8277);
and U8900 (N_8900,N_8019,N_8351);
and U8901 (N_8901,N_8387,N_8041);
xnor U8902 (N_8902,N_8397,N_8161);
nor U8903 (N_8903,N_8204,N_8476);
nor U8904 (N_8904,N_8403,N_8140);
nor U8905 (N_8905,N_8035,N_8022);
or U8906 (N_8906,N_8445,N_8472);
nand U8907 (N_8907,N_8184,N_8073);
and U8908 (N_8908,N_8233,N_8195);
nand U8909 (N_8909,N_8406,N_8446);
nor U8910 (N_8910,N_8067,N_8164);
or U8911 (N_8911,N_8024,N_8406);
nand U8912 (N_8912,N_8013,N_8499);
xor U8913 (N_8913,N_8430,N_8148);
nand U8914 (N_8914,N_8428,N_8106);
or U8915 (N_8915,N_8164,N_8072);
nor U8916 (N_8916,N_8079,N_8165);
nand U8917 (N_8917,N_8299,N_8267);
or U8918 (N_8918,N_8159,N_8458);
xor U8919 (N_8919,N_8413,N_8475);
xnor U8920 (N_8920,N_8097,N_8186);
nand U8921 (N_8921,N_8086,N_8099);
nand U8922 (N_8922,N_8093,N_8253);
and U8923 (N_8923,N_8387,N_8010);
or U8924 (N_8924,N_8015,N_8327);
nand U8925 (N_8925,N_8204,N_8477);
and U8926 (N_8926,N_8139,N_8047);
xor U8927 (N_8927,N_8219,N_8152);
xor U8928 (N_8928,N_8443,N_8277);
xor U8929 (N_8929,N_8066,N_8344);
or U8930 (N_8930,N_8417,N_8324);
or U8931 (N_8931,N_8118,N_8416);
xnor U8932 (N_8932,N_8165,N_8139);
nor U8933 (N_8933,N_8300,N_8151);
nor U8934 (N_8934,N_8168,N_8224);
and U8935 (N_8935,N_8069,N_8247);
or U8936 (N_8936,N_8256,N_8321);
xnor U8937 (N_8937,N_8244,N_8028);
nor U8938 (N_8938,N_8042,N_8157);
nand U8939 (N_8939,N_8040,N_8379);
or U8940 (N_8940,N_8015,N_8082);
xor U8941 (N_8941,N_8295,N_8417);
xnor U8942 (N_8942,N_8344,N_8225);
and U8943 (N_8943,N_8466,N_8255);
and U8944 (N_8944,N_8003,N_8483);
nand U8945 (N_8945,N_8373,N_8374);
nand U8946 (N_8946,N_8398,N_8143);
xnor U8947 (N_8947,N_8428,N_8272);
nand U8948 (N_8948,N_8143,N_8460);
or U8949 (N_8949,N_8062,N_8159);
nor U8950 (N_8950,N_8463,N_8094);
and U8951 (N_8951,N_8381,N_8032);
xor U8952 (N_8952,N_8102,N_8319);
or U8953 (N_8953,N_8274,N_8280);
or U8954 (N_8954,N_8143,N_8217);
nand U8955 (N_8955,N_8308,N_8330);
xor U8956 (N_8956,N_8354,N_8483);
nand U8957 (N_8957,N_8009,N_8027);
nor U8958 (N_8958,N_8300,N_8456);
nand U8959 (N_8959,N_8153,N_8365);
and U8960 (N_8960,N_8063,N_8083);
nand U8961 (N_8961,N_8287,N_8164);
and U8962 (N_8962,N_8197,N_8386);
or U8963 (N_8963,N_8169,N_8032);
xnor U8964 (N_8964,N_8312,N_8354);
nand U8965 (N_8965,N_8424,N_8053);
nor U8966 (N_8966,N_8448,N_8423);
nor U8967 (N_8967,N_8430,N_8067);
nand U8968 (N_8968,N_8394,N_8002);
and U8969 (N_8969,N_8445,N_8381);
nand U8970 (N_8970,N_8078,N_8250);
xor U8971 (N_8971,N_8237,N_8357);
nor U8972 (N_8972,N_8296,N_8081);
and U8973 (N_8973,N_8219,N_8109);
and U8974 (N_8974,N_8471,N_8288);
nand U8975 (N_8975,N_8107,N_8324);
nand U8976 (N_8976,N_8009,N_8276);
nor U8977 (N_8977,N_8254,N_8150);
xor U8978 (N_8978,N_8489,N_8370);
and U8979 (N_8979,N_8027,N_8049);
and U8980 (N_8980,N_8253,N_8033);
or U8981 (N_8981,N_8382,N_8071);
xnor U8982 (N_8982,N_8397,N_8089);
and U8983 (N_8983,N_8226,N_8467);
and U8984 (N_8984,N_8278,N_8433);
or U8985 (N_8985,N_8361,N_8229);
xnor U8986 (N_8986,N_8170,N_8027);
and U8987 (N_8987,N_8166,N_8335);
and U8988 (N_8988,N_8206,N_8133);
xor U8989 (N_8989,N_8089,N_8385);
nand U8990 (N_8990,N_8025,N_8136);
xor U8991 (N_8991,N_8156,N_8315);
xnor U8992 (N_8992,N_8268,N_8179);
and U8993 (N_8993,N_8337,N_8205);
and U8994 (N_8994,N_8237,N_8287);
nand U8995 (N_8995,N_8317,N_8104);
or U8996 (N_8996,N_8283,N_8332);
nor U8997 (N_8997,N_8063,N_8363);
and U8998 (N_8998,N_8361,N_8489);
or U8999 (N_8999,N_8412,N_8101);
nand U9000 (N_9000,N_8845,N_8979);
and U9001 (N_9001,N_8988,N_8698);
nand U9002 (N_9002,N_8636,N_8831);
and U9003 (N_9003,N_8873,N_8977);
and U9004 (N_9004,N_8826,N_8927);
xnor U9005 (N_9005,N_8651,N_8877);
and U9006 (N_9006,N_8894,N_8849);
and U9007 (N_9007,N_8930,N_8991);
nand U9008 (N_9008,N_8607,N_8596);
xnor U9009 (N_9009,N_8934,N_8707);
nand U9010 (N_9010,N_8601,N_8806);
nor U9011 (N_9011,N_8741,N_8678);
or U9012 (N_9012,N_8560,N_8994);
nand U9013 (N_9013,N_8783,N_8896);
or U9014 (N_9014,N_8549,N_8591);
and U9015 (N_9015,N_8587,N_8650);
and U9016 (N_9016,N_8617,N_8971);
nor U9017 (N_9017,N_8833,N_8964);
nor U9018 (N_9018,N_8682,N_8703);
xnor U9019 (N_9019,N_8611,N_8565);
nor U9020 (N_9020,N_8909,N_8809);
xnor U9021 (N_9021,N_8816,N_8693);
nor U9022 (N_9022,N_8840,N_8538);
and U9023 (N_9023,N_8956,N_8644);
nor U9024 (N_9024,N_8668,N_8759);
nor U9025 (N_9025,N_8985,N_8555);
nand U9026 (N_9026,N_8861,N_8666);
nand U9027 (N_9027,N_8615,N_8737);
or U9028 (N_9028,N_8540,N_8745);
nor U9029 (N_9029,N_8616,N_8773);
and U9030 (N_9030,N_8603,N_8642);
nand U9031 (N_9031,N_8545,N_8959);
nor U9032 (N_9032,N_8825,N_8670);
or U9033 (N_9033,N_8695,N_8900);
or U9034 (N_9034,N_8676,N_8802);
xor U9035 (N_9035,N_8867,N_8641);
and U9036 (N_9036,N_8890,N_8761);
nand U9037 (N_9037,N_8594,N_8880);
nor U9038 (N_9038,N_8680,N_8599);
nand U9039 (N_9039,N_8659,N_8697);
and U9040 (N_9040,N_8704,N_8799);
nand U9041 (N_9041,N_8618,N_8700);
nor U9042 (N_9042,N_8923,N_8740);
or U9043 (N_9043,N_8928,N_8951);
nand U9044 (N_9044,N_8683,N_8812);
nor U9045 (N_9045,N_8602,N_8577);
nand U9046 (N_9046,N_8576,N_8583);
nor U9047 (N_9047,N_8661,N_8897);
nand U9048 (N_9048,N_8790,N_8581);
nor U9049 (N_9049,N_8613,N_8818);
xnor U9050 (N_9050,N_8715,N_8733);
and U9051 (N_9051,N_8535,N_8515);
or U9052 (N_9052,N_8557,N_8968);
xnor U9053 (N_9053,N_8620,N_8584);
xnor U9054 (N_9054,N_8905,N_8797);
nand U9055 (N_9055,N_8552,N_8984);
and U9056 (N_9056,N_8972,N_8739);
nand U9057 (N_9057,N_8946,N_8776);
nor U9058 (N_9058,N_8610,N_8958);
nor U9059 (N_9059,N_8888,N_8742);
xnor U9060 (N_9060,N_8865,N_8672);
or U9061 (N_9061,N_8949,N_8820);
and U9062 (N_9062,N_8643,N_8710);
or U9063 (N_9063,N_8689,N_8544);
or U9064 (N_9064,N_8539,N_8992);
nor U9065 (N_9065,N_8690,N_8970);
nand U9066 (N_9066,N_8735,N_8981);
nand U9067 (N_9067,N_8714,N_8886);
nand U9068 (N_9068,N_8559,N_8932);
or U9069 (N_9069,N_8782,N_8630);
and U9070 (N_9070,N_8669,N_8772);
nand U9071 (N_9071,N_8838,N_8609);
nand U9072 (N_9072,N_8671,N_8537);
nor U9073 (N_9073,N_8685,N_8862);
nor U9074 (N_9074,N_8852,N_8796);
and U9075 (N_9075,N_8996,N_8652);
and U9076 (N_9076,N_8542,N_8954);
and U9077 (N_9077,N_8738,N_8995);
and U9078 (N_9078,N_8974,N_8990);
xnor U9079 (N_9079,N_8960,N_8815);
xnor U9080 (N_9080,N_8748,N_8883);
or U9081 (N_9081,N_8983,N_8887);
and U9082 (N_9082,N_8572,N_8752);
and U9083 (N_9083,N_8943,N_8973);
or U9084 (N_9084,N_8645,N_8548);
nor U9085 (N_9085,N_8933,N_8876);
nand U9086 (N_9086,N_8595,N_8784);
or U9087 (N_9087,N_8777,N_8866);
nor U9088 (N_9088,N_8585,N_8863);
and U9089 (N_9089,N_8571,N_8763);
nand U9090 (N_9090,N_8966,N_8639);
nand U9091 (N_9091,N_8899,N_8513);
nand U9092 (N_9092,N_8870,N_8551);
nand U9093 (N_9093,N_8649,N_8526);
or U9094 (N_9094,N_8766,N_8721);
or U9095 (N_9095,N_8502,N_8800);
xnor U9096 (N_9096,N_8658,N_8647);
xor U9097 (N_9097,N_8916,N_8699);
nor U9098 (N_9098,N_8623,N_8924);
nand U9099 (N_9099,N_8997,N_8857);
xor U9100 (N_9100,N_8936,N_8885);
xor U9101 (N_9101,N_8534,N_8921);
or U9102 (N_9102,N_8504,N_8533);
and U9103 (N_9103,N_8638,N_8525);
xor U9104 (N_9104,N_8906,N_8575);
xnor U9105 (N_9105,N_8846,N_8579);
or U9106 (N_9106,N_8633,N_8634);
nand U9107 (N_9107,N_8662,N_8589);
xnor U9108 (N_9108,N_8744,N_8566);
nor U9109 (N_9109,N_8787,N_8901);
or U9110 (N_9110,N_8569,N_8986);
xnor U9111 (N_9111,N_8586,N_8653);
nand U9112 (N_9112,N_8687,N_8881);
and U9113 (N_9113,N_8543,N_8821);
nand U9114 (N_9114,N_8874,N_8531);
xnor U9115 (N_9115,N_8998,N_8774);
and U9116 (N_9116,N_8859,N_8719);
nand U9117 (N_9117,N_8509,N_8764);
xor U9118 (N_9118,N_8528,N_8889);
or U9119 (N_9119,N_8872,N_8965);
nor U9120 (N_9120,N_8629,N_8891);
xor U9121 (N_9121,N_8904,N_8913);
nand U9122 (N_9122,N_8530,N_8953);
or U9123 (N_9123,N_8523,N_8729);
or U9124 (N_9124,N_8590,N_8593);
and U9125 (N_9125,N_8805,N_8788);
nand U9126 (N_9126,N_8856,N_8828);
nor U9127 (N_9127,N_8597,N_8546);
and U9128 (N_9128,N_8918,N_8898);
xnor U9129 (N_9129,N_8541,N_8500);
nand U9130 (N_9130,N_8696,N_8747);
and U9131 (N_9131,N_8632,N_8520);
and U9132 (N_9132,N_8558,N_8875);
nor U9133 (N_9133,N_8789,N_8604);
and U9134 (N_9134,N_8722,N_8762);
and U9135 (N_9135,N_8684,N_8702);
or U9136 (N_9136,N_8769,N_8841);
nor U9137 (N_9137,N_8713,N_8770);
xnor U9138 (N_9138,N_8836,N_8524);
nand U9139 (N_9139,N_8945,N_8824);
nor U9140 (N_9140,N_8794,N_8834);
and U9141 (N_9141,N_8771,N_8963);
xnor U9142 (N_9142,N_8832,N_8758);
and U9143 (N_9143,N_8518,N_8795);
nor U9144 (N_9144,N_8731,N_8780);
xnor U9145 (N_9145,N_8993,N_8847);
nand U9146 (N_9146,N_8674,N_8754);
and U9147 (N_9147,N_8765,N_8786);
nand U9148 (N_9148,N_8871,N_8907);
nor U9149 (N_9149,N_8948,N_8570);
nand U9150 (N_9150,N_8734,N_8708);
xor U9151 (N_9151,N_8660,N_8844);
nor U9152 (N_9152,N_8627,N_8574);
or U9153 (N_9153,N_8978,N_8550);
nor U9154 (N_9154,N_8562,N_8868);
and U9155 (N_9155,N_8519,N_8961);
or U9156 (N_9156,N_8701,N_8506);
or U9157 (N_9157,N_8510,N_8726);
xor U9158 (N_9158,N_8514,N_8681);
nor U9159 (N_9159,N_8631,N_8512);
and U9160 (N_9160,N_8819,N_8622);
xnor U9161 (N_9161,N_8665,N_8655);
or U9162 (N_9162,N_8706,N_8711);
and U9163 (N_9163,N_8619,N_8508);
and U9164 (N_9164,N_8529,N_8792);
or U9165 (N_9165,N_8567,N_8736);
nand U9166 (N_9166,N_8950,N_8839);
and U9167 (N_9167,N_8929,N_8751);
xor U9168 (N_9168,N_8768,N_8612);
nor U9169 (N_9169,N_8635,N_8716);
or U9170 (N_9170,N_8801,N_8648);
and U9171 (N_9171,N_8851,N_8720);
and U9172 (N_9172,N_8536,N_8582);
and U9173 (N_9173,N_8803,N_8743);
or U9174 (N_9174,N_8804,N_8937);
or U9175 (N_9175,N_8848,N_8691);
nand U9176 (N_9176,N_8675,N_8884);
nand U9177 (N_9177,N_8568,N_8791);
nor U9178 (N_9178,N_8882,N_8673);
or U9179 (N_9179,N_8902,N_8982);
xor U9180 (N_9180,N_8915,N_8664);
nor U9181 (N_9181,N_8608,N_8573);
or U9182 (N_9182,N_8592,N_8600);
xnor U9183 (N_9183,N_8753,N_8517);
nor U9184 (N_9184,N_8511,N_8941);
and U9185 (N_9185,N_8922,N_8892);
xor U9186 (N_9186,N_8778,N_8793);
xor U9187 (N_9187,N_8830,N_8926);
or U9188 (N_9188,N_8750,N_8709);
nand U9189 (N_9189,N_8823,N_8903);
or U9190 (N_9190,N_8781,N_8969);
xnor U9191 (N_9191,N_8853,N_8858);
nand U9192 (N_9192,N_8705,N_8999);
and U9193 (N_9193,N_8692,N_8501);
nand U9194 (N_9194,N_8938,N_8925);
nand U9195 (N_9195,N_8967,N_8580);
and U9196 (N_9196,N_8855,N_8654);
and U9197 (N_9197,N_8756,N_8561);
or U9198 (N_9198,N_8908,N_8944);
nor U9199 (N_9199,N_8939,N_8718);
or U9200 (N_9200,N_8606,N_8808);
xor U9201 (N_9201,N_8628,N_8746);
nand U9202 (N_9202,N_8717,N_8728);
nor U9203 (N_9203,N_8869,N_8779);
nand U9204 (N_9204,N_8621,N_8657);
and U9205 (N_9205,N_8980,N_8686);
or U9206 (N_9206,N_8640,N_8864);
and U9207 (N_9207,N_8955,N_8931);
nor U9208 (N_9208,N_8814,N_8843);
and U9209 (N_9209,N_8757,N_8516);
and U9210 (N_9210,N_8521,N_8775);
xnor U9211 (N_9211,N_8588,N_8910);
xor U9212 (N_9212,N_8755,N_8637);
xnor U9213 (N_9213,N_8785,N_8942);
nand U9214 (N_9214,N_8663,N_8811);
nor U9215 (N_9215,N_8625,N_8813);
nor U9216 (N_9216,N_8503,N_8679);
xnor U9217 (N_9217,N_8952,N_8940);
nor U9218 (N_9218,N_8624,N_8614);
xnor U9219 (N_9219,N_8976,N_8626);
nor U9220 (N_9220,N_8646,N_8712);
and U9221 (N_9221,N_8798,N_8760);
xor U9222 (N_9222,N_8829,N_8947);
nor U9223 (N_9223,N_8554,N_8817);
and U9224 (N_9224,N_8919,N_8522);
nand U9225 (N_9225,N_8987,N_8553);
nand U9226 (N_9226,N_8605,N_8732);
nor U9227 (N_9227,N_8912,N_8917);
nor U9228 (N_9228,N_8879,N_8837);
nor U9229 (N_9229,N_8564,N_8957);
xor U9230 (N_9230,N_8920,N_8878);
or U9231 (N_9231,N_8730,N_8827);
nor U9232 (N_9232,N_8807,N_8724);
nor U9233 (N_9233,N_8749,N_8723);
and U9234 (N_9234,N_8822,N_8767);
nor U9235 (N_9235,N_8854,N_8505);
nor U9236 (N_9236,N_8532,N_8893);
nor U9237 (N_9237,N_8563,N_8694);
or U9238 (N_9238,N_8895,N_8667);
xor U9239 (N_9239,N_8962,N_8850);
and U9240 (N_9240,N_8727,N_8547);
or U9241 (N_9241,N_8527,N_8842);
or U9242 (N_9242,N_8688,N_8556);
xnor U9243 (N_9243,N_8935,N_8911);
or U9244 (N_9244,N_8835,N_8860);
nand U9245 (N_9245,N_8810,N_8975);
xor U9246 (N_9246,N_8989,N_8725);
nand U9247 (N_9247,N_8578,N_8507);
and U9248 (N_9248,N_8914,N_8677);
and U9249 (N_9249,N_8656,N_8598);
and U9250 (N_9250,N_8851,N_8958);
xnor U9251 (N_9251,N_8630,N_8719);
nor U9252 (N_9252,N_8648,N_8645);
nor U9253 (N_9253,N_8633,N_8563);
nor U9254 (N_9254,N_8883,N_8888);
nand U9255 (N_9255,N_8759,N_8608);
xnor U9256 (N_9256,N_8809,N_8752);
or U9257 (N_9257,N_8843,N_8759);
and U9258 (N_9258,N_8825,N_8721);
or U9259 (N_9259,N_8815,N_8538);
nor U9260 (N_9260,N_8894,N_8653);
xor U9261 (N_9261,N_8577,N_8536);
nor U9262 (N_9262,N_8718,N_8920);
nand U9263 (N_9263,N_8505,N_8809);
or U9264 (N_9264,N_8775,N_8774);
nand U9265 (N_9265,N_8540,N_8817);
and U9266 (N_9266,N_8940,N_8657);
nand U9267 (N_9267,N_8744,N_8696);
nor U9268 (N_9268,N_8902,N_8918);
nand U9269 (N_9269,N_8882,N_8700);
or U9270 (N_9270,N_8682,N_8679);
nor U9271 (N_9271,N_8728,N_8667);
and U9272 (N_9272,N_8960,N_8564);
xnor U9273 (N_9273,N_8786,N_8528);
nand U9274 (N_9274,N_8634,N_8693);
and U9275 (N_9275,N_8916,N_8751);
xor U9276 (N_9276,N_8831,N_8776);
or U9277 (N_9277,N_8746,N_8768);
nor U9278 (N_9278,N_8627,N_8809);
or U9279 (N_9279,N_8953,N_8929);
and U9280 (N_9280,N_8694,N_8618);
nor U9281 (N_9281,N_8868,N_8812);
or U9282 (N_9282,N_8545,N_8795);
nor U9283 (N_9283,N_8772,N_8990);
nand U9284 (N_9284,N_8600,N_8981);
nand U9285 (N_9285,N_8737,N_8512);
or U9286 (N_9286,N_8624,N_8606);
nand U9287 (N_9287,N_8875,N_8682);
and U9288 (N_9288,N_8660,N_8980);
nand U9289 (N_9289,N_8686,N_8934);
nor U9290 (N_9290,N_8864,N_8688);
and U9291 (N_9291,N_8523,N_8928);
xor U9292 (N_9292,N_8713,N_8818);
nand U9293 (N_9293,N_8873,N_8509);
and U9294 (N_9294,N_8598,N_8770);
nand U9295 (N_9295,N_8980,N_8936);
nand U9296 (N_9296,N_8579,N_8810);
nand U9297 (N_9297,N_8647,N_8556);
nand U9298 (N_9298,N_8991,N_8521);
or U9299 (N_9299,N_8529,N_8801);
and U9300 (N_9300,N_8664,N_8643);
nor U9301 (N_9301,N_8623,N_8713);
nor U9302 (N_9302,N_8544,N_8581);
or U9303 (N_9303,N_8652,N_8974);
nand U9304 (N_9304,N_8874,N_8589);
nand U9305 (N_9305,N_8634,N_8817);
and U9306 (N_9306,N_8617,N_8950);
nor U9307 (N_9307,N_8662,N_8564);
or U9308 (N_9308,N_8946,N_8713);
or U9309 (N_9309,N_8523,N_8683);
or U9310 (N_9310,N_8882,N_8729);
or U9311 (N_9311,N_8889,N_8729);
nand U9312 (N_9312,N_8758,N_8943);
and U9313 (N_9313,N_8634,N_8918);
xnor U9314 (N_9314,N_8647,N_8997);
or U9315 (N_9315,N_8966,N_8693);
nor U9316 (N_9316,N_8778,N_8849);
and U9317 (N_9317,N_8642,N_8725);
nand U9318 (N_9318,N_8786,N_8752);
nand U9319 (N_9319,N_8994,N_8893);
and U9320 (N_9320,N_8783,N_8964);
nor U9321 (N_9321,N_8513,N_8942);
xnor U9322 (N_9322,N_8735,N_8746);
and U9323 (N_9323,N_8766,N_8902);
or U9324 (N_9324,N_8977,N_8950);
and U9325 (N_9325,N_8585,N_8704);
nand U9326 (N_9326,N_8630,N_8897);
and U9327 (N_9327,N_8525,N_8624);
or U9328 (N_9328,N_8716,N_8564);
and U9329 (N_9329,N_8625,N_8743);
and U9330 (N_9330,N_8956,N_8519);
xnor U9331 (N_9331,N_8962,N_8719);
nand U9332 (N_9332,N_8594,N_8885);
nand U9333 (N_9333,N_8880,N_8605);
and U9334 (N_9334,N_8556,N_8769);
nor U9335 (N_9335,N_8542,N_8632);
nand U9336 (N_9336,N_8566,N_8543);
nand U9337 (N_9337,N_8810,N_8698);
nor U9338 (N_9338,N_8831,N_8699);
nor U9339 (N_9339,N_8641,N_8512);
xnor U9340 (N_9340,N_8957,N_8544);
xor U9341 (N_9341,N_8770,N_8969);
nand U9342 (N_9342,N_8567,N_8962);
nor U9343 (N_9343,N_8717,N_8865);
xnor U9344 (N_9344,N_8919,N_8780);
nand U9345 (N_9345,N_8728,N_8705);
nor U9346 (N_9346,N_8669,N_8917);
xnor U9347 (N_9347,N_8709,N_8646);
or U9348 (N_9348,N_8825,N_8515);
and U9349 (N_9349,N_8527,N_8942);
or U9350 (N_9350,N_8680,N_8617);
nor U9351 (N_9351,N_8925,N_8836);
nand U9352 (N_9352,N_8604,N_8872);
nand U9353 (N_9353,N_8980,N_8917);
xnor U9354 (N_9354,N_8756,N_8942);
nor U9355 (N_9355,N_8697,N_8507);
xnor U9356 (N_9356,N_8518,N_8689);
xnor U9357 (N_9357,N_8872,N_8583);
or U9358 (N_9358,N_8592,N_8674);
or U9359 (N_9359,N_8747,N_8904);
xnor U9360 (N_9360,N_8505,N_8785);
nor U9361 (N_9361,N_8741,N_8975);
nand U9362 (N_9362,N_8612,N_8568);
nand U9363 (N_9363,N_8514,N_8544);
nor U9364 (N_9364,N_8996,N_8648);
or U9365 (N_9365,N_8769,N_8669);
nand U9366 (N_9366,N_8865,N_8737);
nor U9367 (N_9367,N_8869,N_8893);
nor U9368 (N_9368,N_8890,N_8551);
nand U9369 (N_9369,N_8597,N_8791);
and U9370 (N_9370,N_8552,N_8633);
nor U9371 (N_9371,N_8573,N_8519);
nand U9372 (N_9372,N_8766,N_8716);
and U9373 (N_9373,N_8666,N_8562);
xnor U9374 (N_9374,N_8626,N_8832);
xnor U9375 (N_9375,N_8571,N_8989);
and U9376 (N_9376,N_8590,N_8890);
nor U9377 (N_9377,N_8781,N_8664);
nor U9378 (N_9378,N_8877,N_8934);
or U9379 (N_9379,N_8891,N_8582);
and U9380 (N_9380,N_8510,N_8522);
nor U9381 (N_9381,N_8978,N_8506);
and U9382 (N_9382,N_8896,N_8707);
and U9383 (N_9383,N_8961,N_8900);
nand U9384 (N_9384,N_8966,N_8698);
and U9385 (N_9385,N_8596,N_8546);
xor U9386 (N_9386,N_8577,N_8752);
xnor U9387 (N_9387,N_8724,N_8924);
xor U9388 (N_9388,N_8599,N_8989);
and U9389 (N_9389,N_8647,N_8749);
nor U9390 (N_9390,N_8666,N_8941);
nor U9391 (N_9391,N_8967,N_8791);
and U9392 (N_9392,N_8833,N_8871);
nor U9393 (N_9393,N_8624,N_8701);
or U9394 (N_9394,N_8968,N_8695);
nor U9395 (N_9395,N_8556,N_8727);
xor U9396 (N_9396,N_8612,N_8800);
and U9397 (N_9397,N_8947,N_8520);
and U9398 (N_9398,N_8846,N_8512);
and U9399 (N_9399,N_8958,N_8766);
nand U9400 (N_9400,N_8826,N_8679);
nand U9401 (N_9401,N_8566,N_8524);
xor U9402 (N_9402,N_8910,N_8581);
and U9403 (N_9403,N_8812,N_8839);
and U9404 (N_9404,N_8622,N_8607);
nor U9405 (N_9405,N_8726,N_8944);
xnor U9406 (N_9406,N_8938,N_8726);
and U9407 (N_9407,N_8824,N_8865);
and U9408 (N_9408,N_8804,N_8897);
nand U9409 (N_9409,N_8992,N_8796);
and U9410 (N_9410,N_8877,N_8843);
or U9411 (N_9411,N_8603,N_8548);
xnor U9412 (N_9412,N_8978,N_8555);
xnor U9413 (N_9413,N_8822,N_8704);
and U9414 (N_9414,N_8885,N_8727);
nor U9415 (N_9415,N_8657,N_8672);
nand U9416 (N_9416,N_8500,N_8620);
nor U9417 (N_9417,N_8533,N_8980);
and U9418 (N_9418,N_8782,N_8697);
or U9419 (N_9419,N_8511,N_8645);
nand U9420 (N_9420,N_8809,N_8855);
or U9421 (N_9421,N_8796,N_8862);
or U9422 (N_9422,N_8973,N_8800);
nor U9423 (N_9423,N_8617,N_8787);
nor U9424 (N_9424,N_8564,N_8527);
xnor U9425 (N_9425,N_8909,N_8767);
nor U9426 (N_9426,N_8908,N_8678);
or U9427 (N_9427,N_8655,N_8885);
or U9428 (N_9428,N_8865,N_8964);
xnor U9429 (N_9429,N_8647,N_8775);
nand U9430 (N_9430,N_8802,N_8823);
nand U9431 (N_9431,N_8531,N_8963);
or U9432 (N_9432,N_8848,N_8550);
nor U9433 (N_9433,N_8881,N_8939);
xnor U9434 (N_9434,N_8962,N_8846);
nor U9435 (N_9435,N_8575,N_8590);
nor U9436 (N_9436,N_8845,N_8629);
and U9437 (N_9437,N_8975,N_8606);
or U9438 (N_9438,N_8874,N_8805);
and U9439 (N_9439,N_8975,N_8573);
and U9440 (N_9440,N_8503,N_8788);
nor U9441 (N_9441,N_8836,N_8674);
or U9442 (N_9442,N_8500,N_8501);
and U9443 (N_9443,N_8603,N_8508);
nor U9444 (N_9444,N_8699,N_8962);
xnor U9445 (N_9445,N_8905,N_8675);
and U9446 (N_9446,N_8972,N_8783);
nand U9447 (N_9447,N_8857,N_8622);
or U9448 (N_9448,N_8931,N_8541);
xor U9449 (N_9449,N_8619,N_8823);
nand U9450 (N_9450,N_8537,N_8526);
nand U9451 (N_9451,N_8812,N_8892);
nor U9452 (N_9452,N_8740,N_8682);
or U9453 (N_9453,N_8863,N_8980);
nand U9454 (N_9454,N_8800,N_8897);
and U9455 (N_9455,N_8800,N_8866);
or U9456 (N_9456,N_8625,N_8668);
xor U9457 (N_9457,N_8726,N_8703);
nand U9458 (N_9458,N_8844,N_8867);
nor U9459 (N_9459,N_8862,N_8841);
xnor U9460 (N_9460,N_8611,N_8956);
or U9461 (N_9461,N_8765,N_8936);
or U9462 (N_9462,N_8571,N_8576);
xnor U9463 (N_9463,N_8711,N_8515);
nand U9464 (N_9464,N_8661,N_8641);
nand U9465 (N_9465,N_8771,N_8797);
and U9466 (N_9466,N_8768,N_8556);
and U9467 (N_9467,N_8854,N_8651);
xor U9468 (N_9468,N_8983,N_8547);
or U9469 (N_9469,N_8654,N_8974);
and U9470 (N_9470,N_8832,N_8564);
and U9471 (N_9471,N_8846,N_8854);
nor U9472 (N_9472,N_8592,N_8851);
or U9473 (N_9473,N_8707,N_8663);
nand U9474 (N_9474,N_8658,N_8826);
or U9475 (N_9475,N_8751,N_8718);
nand U9476 (N_9476,N_8633,N_8512);
nor U9477 (N_9477,N_8975,N_8852);
nor U9478 (N_9478,N_8670,N_8550);
nand U9479 (N_9479,N_8603,N_8856);
and U9480 (N_9480,N_8921,N_8886);
nand U9481 (N_9481,N_8626,N_8544);
nor U9482 (N_9482,N_8562,N_8955);
nor U9483 (N_9483,N_8691,N_8963);
xnor U9484 (N_9484,N_8677,N_8840);
and U9485 (N_9485,N_8647,N_8535);
or U9486 (N_9486,N_8683,N_8831);
nor U9487 (N_9487,N_8780,N_8862);
nor U9488 (N_9488,N_8701,N_8823);
or U9489 (N_9489,N_8644,N_8676);
nand U9490 (N_9490,N_8728,N_8962);
nor U9491 (N_9491,N_8626,N_8986);
nor U9492 (N_9492,N_8539,N_8925);
nor U9493 (N_9493,N_8585,N_8643);
nor U9494 (N_9494,N_8662,N_8548);
nand U9495 (N_9495,N_8718,N_8897);
nand U9496 (N_9496,N_8544,N_8844);
and U9497 (N_9497,N_8996,N_8874);
and U9498 (N_9498,N_8972,N_8651);
xor U9499 (N_9499,N_8603,N_8868);
and U9500 (N_9500,N_9468,N_9305);
or U9501 (N_9501,N_9013,N_9362);
and U9502 (N_9502,N_9392,N_9303);
nor U9503 (N_9503,N_9434,N_9312);
nor U9504 (N_9504,N_9272,N_9058);
nand U9505 (N_9505,N_9306,N_9060);
nor U9506 (N_9506,N_9154,N_9337);
or U9507 (N_9507,N_9111,N_9228);
nand U9508 (N_9508,N_9093,N_9103);
and U9509 (N_9509,N_9250,N_9295);
nand U9510 (N_9510,N_9176,N_9321);
and U9511 (N_9511,N_9401,N_9268);
xor U9512 (N_9512,N_9419,N_9325);
or U9513 (N_9513,N_9023,N_9221);
or U9514 (N_9514,N_9429,N_9424);
or U9515 (N_9515,N_9369,N_9115);
xor U9516 (N_9516,N_9237,N_9456);
nor U9517 (N_9517,N_9192,N_9018);
and U9518 (N_9518,N_9191,N_9219);
and U9519 (N_9519,N_9229,N_9186);
or U9520 (N_9520,N_9375,N_9099);
nor U9521 (N_9521,N_9061,N_9179);
nor U9522 (N_9522,N_9200,N_9175);
nand U9523 (N_9523,N_9478,N_9049);
and U9524 (N_9524,N_9247,N_9129);
or U9525 (N_9525,N_9435,N_9162);
nand U9526 (N_9526,N_9274,N_9213);
nand U9527 (N_9527,N_9291,N_9211);
nor U9528 (N_9528,N_9113,N_9085);
and U9529 (N_9529,N_9430,N_9395);
nor U9530 (N_9530,N_9479,N_9293);
nand U9531 (N_9531,N_9070,N_9351);
nand U9532 (N_9532,N_9064,N_9254);
nand U9533 (N_9533,N_9102,N_9195);
nand U9534 (N_9534,N_9095,N_9109);
or U9535 (N_9535,N_9040,N_9354);
nand U9536 (N_9536,N_9053,N_9051);
or U9537 (N_9537,N_9091,N_9065);
nor U9538 (N_9538,N_9164,N_9133);
nor U9539 (N_9539,N_9309,N_9017);
nor U9540 (N_9540,N_9160,N_9216);
nor U9541 (N_9541,N_9277,N_9033);
and U9542 (N_9542,N_9495,N_9346);
and U9543 (N_9543,N_9173,N_9433);
and U9544 (N_9544,N_9112,N_9097);
xor U9545 (N_9545,N_9364,N_9082);
xor U9546 (N_9546,N_9130,N_9232);
xnor U9547 (N_9547,N_9482,N_9038);
nand U9548 (N_9548,N_9122,N_9035);
xnor U9549 (N_9549,N_9452,N_9444);
nor U9550 (N_9550,N_9246,N_9220);
nor U9551 (N_9551,N_9454,N_9032);
and U9552 (N_9552,N_9014,N_9402);
nand U9553 (N_9553,N_9279,N_9118);
or U9554 (N_9554,N_9207,N_9174);
xor U9555 (N_9555,N_9413,N_9438);
nand U9556 (N_9556,N_9043,N_9374);
nor U9557 (N_9557,N_9345,N_9157);
or U9558 (N_9558,N_9496,N_9031);
or U9559 (N_9559,N_9236,N_9089);
or U9560 (N_9560,N_9336,N_9359);
and U9561 (N_9561,N_9125,N_9094);
and U9562 (N_9562,N_9466,N_9259);
or U9563 (N_9563,N_9255,N_9080);
nor U9564 (N_9564,N_9432,N_9230);
nand U9565 (N_9565,N_9441,N_9439);
nor U9566 (N_9566,N_9172,N_9187);
or U9567 (N_9567,N_9296,N_9119);
and U9568 (N_9568,N_9077,N_9282);
and U9569 (N_9569,N_9404,N_9161);
nand U9570 (N_9570,N_9283,N_9223);
nand U9571 (N_9571,N_9238,N_9193);
nor U9572 (N_9572,N_9455,N_9492);
xnor U9573 (N_9573,N_9298,N_9066);
nor U9574 (N_9574,N_9458,N_9069);
nand U9575 (N_9575,N_9499,N_9147);
nor U9576 (N_9576,N_9227,N_9015);
nor U9577 (N_9577,N_9090,N_9009);
or U9578 (N_9578,N_9156,N_9101);
nand U9579 (N_9579,N_9280,N_9206);
and U9580 (N_9580,N_9394,N_9356);
xnor U9581 (N_9581,N_9029,N_9287);
nand U9582 (N_9582,N_9411,N_9343);
xnor U9583 (N_9583,N_9096,N_9241);
nor U9584 (N_9584,N_9263,N_9275);
nor U9585 (N_9585,N_9169,N_9436);
and U9586 (N_9586,N_9471,N_9467);
nor U9587 (N_9587,N_9235,N_9063);
and U9588 (N_9588,N_9039,N_9218);
xor U9589 (N_9589,N_9453,N_9002);
nor U9590 (N_9590,N_9257,N_9037);
nor U9591 (N_9591,N_9300,N_9184);
nor U9592 (N_9592,N_9322,N_9056);
nand U9593 (N_9593,N_9417,N_9067);
nand U9594 (N_9594,N_9363,N_9188);
or U9595 (N_9595,N_9477,N_9057);
nand U9596 (N_9596,N_9062,N_9408);
xnor U9597 (N_9597,N_9016,N_9372);
or U9598 (N_9598,N_9311,N_9365);
nor U9599 (N_9599,N_9198,N_9106);
or U9600 (N_9600,N_9290,N_9324);
and U9601 (N_9601,N_9258,N_9025);
and U9602 (N_9602,N_9072,N_9476);
xnor U9603 (N_9603,N_9138,N_9110);
and U9604 (N_9604,N_9137,N_9407);
xnor U9605 (N_9605,N_9001,N_9423);
nor U9606 (N_9606,N_9486,N_9197);
xnor U9607 (N_9607,N_9339,N_9338);
xor U9608 (N_9608,N_9000,N_9403);
xor U9609 (N_9609,N_9472,N_9483);
and U9610 (N_9610,N_9368,N_9445);
nand U9611 (N_9611,N_9044,N_9024);
or U9612 (N_9612,N_9448,N_9212);
nand U9613 (N_9613,N_9159,N_9415);
and U9614 (N_9614,N_9320,N_9270);
or U9615 (N_9615,N_9030,N_9326);
and U9616 (N_9616,N_9028,N_9204);
or U9617 (N_9617,N_9127,N_9301);
nor U9618 (N_9618,N_9412,N_9047);
xnor U9619 (N_9619,N_9202,N_9331);
nand U9620 (N_9620,N_9196,N_9153);
or U9621 (N_9621,N_9449,N_9469);
and U9622 (N_9622,N_9075,N_9285);
and U9623 (N_9623,N_9457,N_9328);
and U9624 (N_9624,N_9352,N_9052);
and U9625 (N_9625,N_9481,N_9034);
nor U9626 (N_9626,N_9450,N_9386);
nor U9627 (N_9627,N_9086,N_9353);
and U9628 (N_9628,N_9234,N_9209);
and U9629 (N_9629,N_9284,N_9107);
xor U9630 (N_9630,N_9244,N_9414);
and U9631 (N_9631,N_9281,N_9006);
nor U9632 (N_9632,N_9494,N_9489);
or U9633 (N_9633,N_9189,N_9149);
and U9634 (N_9634,N_9260,N_9177);
nand U9635 (N_9635,N_9005,N_9132);
nor U9636 (N_9636,N_9140,N_9488);
nor U9637 (N_9637,N_9048,N_9314);
xor U9638 (N_9638,N_9418,N_9431);
xor U9639 (N_9639,N_9021,N_9400);
nand U9640 (N_9640,N_9329,N_9340);
xor U9641 (N_9641,N_9010,N_9335);
and U9642 (N_9642,N_9498,N_9054);
or U9643 (N_9643,N_9273,N_9083);
and U9644 (N_9644,N_9341,N_9243);
nand U9645 (N_9645,N_9461,N_9170);
or U9646 (N_9646,N_9366,N_9276);
xnor U9647 (N_9647,N_9380,N_9022);
or U9648 (N_9648,N_9383,N_9078);
and U9649 (N_9649,N_9373,N_9165);
and U9650 (N_9650,N_9146,N_9425);
or U9651 (N_9651,N_9242,N_9464);
or U9652 (N_9652,N_9185,N_9484);
and U9653 (N_9653,N_9194,N_9168);
xnor U9654 (N_9654,N_9388,N_9092);
or U9655 (N_9655,N_9117,N_9289);
nand U9656 (N_9656,N_9098,N_9249);
nor U9657 (N_9657,N_9490,N_9178);
and U9658 (N_9658,N_9286,N_9307);
nand U9659 (N_9659,N_9349,N_9355);
xnor U9660 (N_9660,N_9139,N_9134);
or U9661 (N_9661,N_9152,N_9084);
or U9662 (N_9662,N_9074,N_9378);
and U9663 (N_9663,N_9406,N_9382);
or U9664 (N_9664,N_9334,N_9473);
nor U9665 (N_9665,N_9155,N_9357);
nor U9666 (N_9666,N_9203,N_9076);
or U9667 (N_9667,N_9264,N_9042);
nor U9668 (N_9668,N_9302,N_9148);
or U9669 (N_9669,N_9465,N_9451);
and U9670 (N_9670,N_9447,N_9123);
nand U9671 (N_9671,N_9391,N_9226);
or U9672 (N_9672,N_9233,N_9493);
and U9673 (N_9673,N_9003,N_9261);
or U9674 (N_9674,N_9371,N_9377);
nor U9675 (N_9675,N_9208,N_9027);
nand U9676 (N_9676,N_9379,N_9294);
and U9677 (N_9677,N_9239,N_9318);
nor U9678 (N_9678,N_9055,N_9304);
or U9679 (N_9679,N_9087,N_9114);
nor U9680 (N_9680,N_9396,N_9428);
or U9681 (N_9681,N_9019,N_9350);
nand U9682 (N_9682,N_9361,N_9399);
or U9683 (N_9683,N_9292,N_9358);
nor U9684 (N_9684,N_9491,N_9248);
nor U9685 (N_9685,N_9384,N_9166);
and U9686 (N_9686,N_9121,N_9141);
nor U9687 (N_9687,N_9059,N_9143);
nand U9688 (N_9688,N_9385,N_9442);
nand U9689 (N_9689,N_9199,N_9462);
or U9690 (N_9690,N_9167,N_9446);
nand U9691 (N_9691,N_9079,N_9262);
and U9692 (N_9692,N_9007,N_9460);
or U9693 (N_9693,N_9136,N_9108);
or U9694 (N_9694,N_9316,N_9151);
nand U9695 (N_9695,N_9426,N_9330);
and U9696 (N_9696,N_9381,N_9308);
nor U9697 (N_9697,N_9011,N_9267);
nor U9698 (N_9698,N_9313,N_9265);
and U9699 (N_9699,N_9182,N_9266);
xnor U9700 (N_9700,N_9183,N_9397);
and U9701 (N_9701,N_9104,N_9142);
or U9702 (N_9702,N_9120,N_9474);
and U9703 (N_9703,N_9041,N_9145);
or U9704 (N_9704,N_9463,N_9323);
and U9705 (N_9705,N_9440,N_9297);
xnor U9706 (N_9706,N_9071,N_9150);
xor U9707 (N_9707,N_9475,N_9420);
nor U9708 (N_9708,N_9171,N_9215);
nor U9709 (N_9709,N_9100,N_9004);
and U9710 (N_9710,N_9008,N_9126);
nor U9711 (N_9711,N_9427,N_9144);
or U9712 (N_9712,N_9214,N_9181);
or U9713 (N_9713,N_9333,N_9421);
nor U9714 (N_9714,N_9158,N_9327);
or U9715 (N_9715,N_9470,N_9240);
and U9716 (N_9716,N_9315,N_9344);
nand U9717 (N_9717,N_9342,N_9347);
nand U9718 (N_9718,N_9487,N_9116);
or U9719 (N_9719,N_9348,N_9251);
or U9720 (N_9720,N_9256,N_9269);
or U9721 (N_9721,N_9081,N_9319);
and U9722 (N_9722,N_9073,N_9278);
nand U9723 (N_9723,N_9317,N_9480);
nor U9724 (N_9724,N_9046,N_9390);
nand U9725 (N_9725,N_9231,N_9245);
and U9726 (N_9726,N_9405,N_9485);
nor U9727 (N_9727,N_9367,N_9105);
nand U9728 (N_9728,N_9224,N_9497);
nor U9729 (N_9729,N_9217,N_9332);
and U9730 (N_9730,N_9201,N_9310);
and U9731 (N_9731,N_9370,N_9422);
or U9732 (N_9732,N_9180,N_9036);
nor U9733 (N_9733,N_9190,N_9387);
nand U9734 (N_9734,N_9135,N_9026);
xor U9735 (N_9735,N_9210,N_9271);
xor U9736 (N_9736,N_9252,N_9068);
nand U9737 (N_9737,N_9459,N_9299);
xor U9738 (N_9738,N_9050,N_9409);
and U9739 (N_9739,N_9389,N_9131);
xor U9740 (N_9740,N_9410,N_9360);
and U9741 (N_9741,N_9045,N_9225);
and U9742 (N_9742,N_9253,N_9437);
nor U9743 (N_9743,N_9124,N_9163);
xnor U9744 (N_9744,N_9288,N_9416);
nor U9745 (N_9745,N_9398,N_9012);
and U9746 (N_9746,N_9376,N_9128);
nor U9747 (N_9747,N_9088,N_9443);
nor U9748 (N_9748,N_9205,N_9222);
and U9749 (N_9749,N_9393,N_9020);
and U9750 (N_9750,N_9165,N_9009);
and U9751 (N_9751,N_9167,N_9017);
nand U9752 (N_9752,N_9221,N_9101);
and U9753 (N_9753,N_9458,N_9377);
and U9754 (N_9754,N_9495,N_9261);
xnor U9755 (N_9755,N_9159,N_9320);
nand U9756 (N_9756,N_9026,N_9235);
nand U9757 (N_9757,N_9012,N_9344);
or U9758 (N_9758,N_9294,N_9464);
nand U9759 (N_9759,N_9225,N_9006);
and U9760 (N_9760,N_9136,N_9167);
and U9761 (N_9761,N_9336,N_9282);
nor U9762 (N_9762,N_9312,N_9208);
nand U9763 (N_9763,N_9424,N_9255);
or U9764 (N_9764,N_9462,N_9185);
and U9765 (N_9765,N_9119,N_9238);
xnor U9766 (N_9766,N_9090,N_9041);
and U9767 (N_9767,N_9352,N_9324);
and U9768 (N_9768,N_9100,N_9190);
and U9769 (N_9769,N_9017,N_9320);
nand U9770 (N_9770,N_9216,N_9314);
or U9771 (N_9771,N_9065,N_9000);
xor U9772 (N_9772,N_9378,N_9056);
and U9773 (N_9773,N_9298,N_9096);
and U9774 (N_9774,N_9164,N_9070);
and U9775 (N_9775,N_9232,N_9114);
xor U9776 (N_9776,N_9051,N_9229);
and U9777 (N_9777,N_9302,N_9255);
nand U9778 (N_9778,N_9308,N_9151);
xnor U9779 (N_9779,N_9424,N_9022);
xnor U9780 (N_9780,N_9256,N_9108);
nor U9781 (N_9781,N_9463,N_9410);
and U9782 (N_9782,N_9112,N_9265);
nor U9783 (N_9783,N_9399,N_9175);
or U9784 (N_9784,N_9223,N_9048);
nand U9785 (N_9785,N_9085,N_9136);
xnor U9786 (N_9786,N_9240,N_9169);
or U9787 (N_9787,N_9126,N_9412);
and U9788 (N_9788,N_9141,N_9480);
xor U9789 (N_9789,N_9032,N_9152);
xnor U9790 (N_9790,N_9378,N_9008);
or U9791 (N_9791,N_9031,N_9229);
nand U9792 (N_9792,N_9093,N_9052);
or U9793 (N_9793,N_9097,N_9246);
and U9794 (N_9794,N_9260,N_9081);
xor U9795 (N_9795,N_9380,N_9476);
or U9796 (N_9796,N_9361,N_9223);
nand U9797 (N_9797,N_9294,N_9390);
and U9798 (N_9798,N_9005,N_9486);
and U9799 (N_9799,N_9021,N_9338);
or U9800 (N_9800,N_9250,N_9467);
nor U9801 (N_9801,N_9373,N_9009);
and U9802 (N_9802,N_9172,N_9314);
xnor U9803 (N_9803,N_9442,N_9217);
nand U9804 (N_9804,N_9336,N_9416);
xor U9805 (N_9805,N_9338,N_9461);
nand U9806 (N_9806,N_9256,N_9409);
nor U9807 (N_9807,N_9279,N_9352);
and U9808 (N_9808,N_9141,N_9166);
and U9809 (N_9809,N_9422,N_9467);
nand U9810 (N_9810,N_9091,N_9220);
or U9811 (N_9811,N_9395,N_9118);
nor U9812 (N_9812,N_9440,N_9049);
and U9813 (N_9813,N_9052,N_9280);
or U9814 (N_9814,N_9216,N_9199);
or U9815 (N_9815,N_9045,N_9049);
or U9816 (N_9816,N_9457,N_9375);
or U9817 (N_9817,N_9284,N_9124);
xor U9818 (N_9818,N_9352,N_9321);
or U9819 (N_9819,N_9351,N_9251);
nand U9820 (N_9820,N_9294,N_9337);
nor U9821 (N_9821,N_9117,N_9371);
nand U9822 (N_9822,N_9036,N_9261);
or U9823 (N_9823,N_9314,N_9296);
and U9824 (N_9824,N_9345,N_9274);
xnor U9825 (N_9825,N_9029,N_9100);
nand U9826 (N_9826,N_9145,N_9425);
nand U9827 (N_9827,N_9427,N_9290);
nand U9828 (N_9828,N_9373,N_9163);
and U9829 (N_9829,N_9076,N_9440);
nand U9830 (N_9830,N_9277,N_9015);
nand U9831 (N_9831,N_9178,N_9085);
nand U9832 (N_9832,N_9118,N_9335);
xor U9833 (N_9833,N_9283,N_9305);
and U9834 (N_9834,N_9022,N_9404);
nor U9835 (N_9835,N_9166,N_9365);
nor U9836 (N_9836,N_9062,N_9061);
nor U9837 (N_9837,N_9271,N_9314);
or U9838 (N_9838,N_9103,N_9169);
nor U9839 (N_9839,N_9254,N_9374);
and U9840 (N_9840,N_9000,N_9438);
or U9841 (N_9841,N_9284,N_9122);
and U9842 (N_9842,N_9454,N_9450);
xor U9843 (N_9843,N_9009,N_9208);
nor U9844 (N_9844,N_9260,N_9224);
nand U9845 (N_9845,N_9186,N_9049);
nand U9846 (N_9846,N_9463,N_9060);
nor U9847 (N_9847,N_9113,N_9173);
nor U9848 (N_9848,N_9265,N_9162);
xnor U9849 (N_9849,N_9050,N_9025);
nor U9850 (N_9850,N_9494,N_9034);
or U9851 (N_9851,N_9025,N_9082);
and U9852 (N_9852,N_9047,N_9049);
xor U9853 (N_9853,N_9141,N_9325);
xnor U9854 (N_9854,N_9395,N_9123);
or U9855 (N_9855,N_9064,N_9185);
and U9856 (N_9856,N_9414,N_9321);
xor U9857 (N_9857,N_9423,N_9368);
or U9858 (N_9858,N_9484,N_9025);
xnor U9859 (N_9859,N_9450,N_9176);
or U9860 (N_9860,N_9156,N_9124);
nand U9861 (N_9861,N_9273,N_9194);
nand U9862 (N_9862,N_9454,N_9017);
nand U9863 (N_9863,N_9402,N_9080);
nand U9864 (N_9864,N_9290,N_9114);
nor U9865 (N_9865,N_9113,N_9349);
xor U9866 (N_9866,N_9243,N_9364);
xor U9867 (N_9867,N_9447,N_9207);
nor U9868 (N_9868,N_9004,N_9306);
or U9869 (N_9869,N_9202,N_9375);
xor U9870 (N_9870,N_9129,N_9366);
nand U9871 (N_9871,N_9225,N_9063);
nand U9872 (N_9872,N_9014,N_9419);
xor U9873 (N_9873,N_9084,N_9410);
xor U9874 (N_9874,N_9310,N_9174);
xnor U9875 (N_9875,N_9428,N_9251);
and U9876 (N_9876,N_9302,N_9064);
xor U9877 (N_9877,N_9394,N_9370);
nand U9878 (N_9878,N_9483,N_9200);
xnor U9879 (N_9879,N_9366,N_9428);
nor U9880 (N_9880,N_9122,N_9010);
and U9881 (N_9881,N_9043,N_9337);
nor U9882 (N_9882,N_9110,N_9072);
nor U9883 (N_9883,N_9115,N_9451);
xor U9884 (N_9884,N_9157,N_9406);
and U9885 (N_9885,N_9201,N_9228);
xor U9886 (N_9886,N_9358,N_9401);
and U9887 (N_9887,N_9141,N_9147);
and U9888 (N_9888,N_9429,N_9498);
and U9889 (N_9889,N_9087,N_9231);
nand U9890 (N_9890,N_9080,N_9264);
xnor U9891 (N_9891,N_9223,N_9459);
nor U9892 (N_9892,N_9466,N_9309);
xnor U9893 (N_9893,N_9420,N_9331);
nor U9894 (N_9894,N_9467,N_9227);
nand U9895 (N_9895,N_9217,N_9431);
and U9896 (N_9896,N_9229,N_9391);
and U9897 (N_9897,N_9142,N_9300);
nor U9898 (N_9898,N_9366,N_9261);
or U9899 (N_9899,N_9350,N_9154);
or U9900 (N_9900,N_9294,N_9229);
xnor U9901 (N_9901,N_9341,N_9482);
nand U9902 (N_9902,N_9298,N_9424);
nor U9903 (N_9903,N_9223,N_9084);
and U9904 (N_9904,N_9259,N_9060);
and U9905 (N_9905,N_9101,N_9445);
xnor U9906 (N_9906,N_9136,N_9068);
or U9907 (N_9907,N_9039,N_9192);
nor U9908 (N_9908,N_9304,N_9143);
and U9909 (N_9909,N_9364,N_9148);
or U9910 (N_9910,N_9337,N_9357);
or U9911 (N_9911,N_9151,N_9207);
nor U9912 (N_9912,N_9363,N_9155);
xnor U9913 (N_9913,N_9026,N_9001);
nand U9914 (N_9914,N_9486,N_9351);
nand U9915 (N_9915,N_9229,N_9332);
nor U9916 (N_9916,N_9093,N_9331);
xor U9917 (N_9917,N_9117,N_9482);
nor U9918 (N_9918,N_9448,N_9230);
and U9919 (N_9919,N_9107,N_9451);
nor U9920 (N_9920,N_9301,N_9156);
or U9921 (N_9921,N_9473,N_9153);
xnor U9922 (N_9922,N_9284,N_9116);
and U9923 (N_9923,N_9240,N_9247);
or U9924 (N_9924,N_9181,N_9434);
nor U9925 (N_9925,N_9122,N_9220);
nand U9926 (N_9926,N_9026,N_9040);
nand U9927 (N_9927,N_9360,N_9109);
nor U9928 (N_9928,N_9334,N_9210);
xnor U9929 (N_9929,N_9040,N_9024);
nor U9930 (N_9930,N_9052,N_9180);
or U9931 (N_9931,N_9059,N_9047);
nand U9932 (N_9932,N_9073,N_9198);
nand U9933 (N_9933,N_9086,N_9489);
xnor U9934 (N_9934,N_9048,N_9272);
nand U9935 (N_9935,N_9140,N_9201);
and U9936 (N_9936,N_9118,N_9242);
or U9937 (N_9937,N_9010,N_9341);
and U9938 (N_9938,N_9284,N_9017);
nand U9939 (N_9939,N_9157,N_9212);
xnor U9940 (N_9940,N_9222,N_9435);
nand U9941 (N_9941,N_9368,N_9211);
xnor U9942 (N_9942,N_9378,N_9202);
xor U9943 (N_9943,N_9158,N_9160);
nand U9944 (N_9944,N_9100,N_9201);
nand U9945 (N_9945,N_9372,N_9453);
and U9946 (N_9946,N_9389,N_9106);
nand U9947 (N_9947,N_9154,N_9045);
nor U9948 (N_9948,N_9265,N_9246);
nor U9949 (N_9949,N_9387,N_9441);
and U9950 (N_9950,N_9164,N_9214);
and U9951 (N_9951,N_9015,N_9092);
xor U9952 (N_9952,N_9046,N_9020);
and U9953 (N_9953,N_9068,N_9345);
xor U9954 (N_9954,N_9332,N_9379);
xor U9955 (N_9955,N_9196,N_9078);
nand U9956 (N_9956,N_9101,N_9357);
nand U9957 (N_9957,N_9028,N_9453);
or U9958 (N_9958,N_9241,N_9253);
nor U9959 (N_9959,N_9382,N_9197);
or U9960 (N_9960,N_9315,N_9003);
nor U9961 (N_9961,N_9229,N_9035);
and U9962 (N_9962,N_9125,N_9278);
and U9963 (N_9963,N_9405,N_9369);
nor U9964 (N_9964,N_9384,N_9272);
or U9965 (N_9965,N_9181,N_9261);
xnor U9966 (N_9966,N_9298,N_9315);
nor U9967 (N_9967,N_9347,N_9333);
nor U9968 (N_9968,N_9471,N_9097);
nor U9969 (N_9969,N_9394,N_9431);
nor U9970 (N_9970,N_9332,N_9178);
nand U9971 (N_9971,N_9248,N_9189);
or U9972 (N_9972,N_9290,N_9081);
xor U9973 (N_9973,N_9302,N_9040);
xnor U9974 (N_9974,N_9335,N_9231);
xnor U9975 (N_9975,N_9339,N_9251);
nand U9976 (N_9976,N_9124,N_9248);
xor U9977 (N_9977,N_9047,N_9214);
nor U9978 (N_9978,N_9453,N_9370);
xor U9979 (N_9979,N_9139,N_9199);
nor U9980 (N_9980,N_9081,N_9372);
nand U9981 (N_9981,N_9246,N_9191);
xnor U9982 (N_9982,N_9108,N_9057);
or U9983 (N_9983,N_9495,N_9412);
nor U9984 (N_9984,N_9273,N_9239);
and U9985 (N_9985,N_9414,N_9139);
nor U9986 (N_9986,N_9065,N_9349);
xnor U9987 (N_9987,N_9245,N_9454);
and U9988 (N_9988,N_9114,N_9302);
or U9989 (N_9989,N_9473,N_9295);
and U9990 (N_9990,N_9251,N_9199);
nor U9991 (N_9991,N_9207,N_9180);
and U9992 (N_9992,N_9331,N_9401);
xor U9993 (N_9993,N_9396,N_9146);
or U9994 (N_9994,N_9318,N_9116);
nand U9995 (N_9995,N_9311,N_9212);
nor U9996 (N_9996,N_9342,N_9249);
or U9997 (N_9997,N_9124,N_9233);
or U9998 (N_9998,N_9046,N_9214);
and U9999 (N_9999,N_9258,N_9320);
nor U10000 (N_10000,N_9897,N_9607);
nand U10001 (N_10001,N_9919,N_9899);
or U10002 (N_10002,N_9650,N_9742);
nand U10003 (N_10003,N_9905,N_9608);
or U10004 (N_10004,N_9846,N_9610);
nand U10005 (N_10005,N_9616,N_9868);
nand U10006 (N_10006,N_9848,N_9936);
or U10007 (N_10007,N_9702,N_9827);
nand U10008 (N_10008,N_9867,N_9979);
and U10009 (N_10009,N_9681,N_9554);
nand U10010 (N_10010,N_9631,N_9830);
or U10011 (N_10011,N_9926,N_9525);
xnor U10012 (N_10012,N_9747,N_9706);
nor U10013 (N_10013,N_9965,N_9611);
and U10014 (N_10014,N_9595,N_9874);
nand U10015 (N_10015,N_9977,N_9673);
xnor U10016 (N_10016,N_9590,N_9816);
or U10017 (N_10017,N_9916,N_9589);
nand U10018 (N_10018,N_9643,N_9885);
nor U10019 (N_10019,N_9800,N_9748);
or U10020 (N_10020,N_9869,N_9508);
or U10021 (N_10021,N_9985,N_9888);
nand U10022 (N_10022,N_9907,N_9829);
xor U10023 (N_10023,N_9939,N_9909);
and U10024 (N_10024,N_9606,N_9730);
and U10025 (N_10025,N_9638,N_9957);
and U10026 (N_10026,N_9860,N_9657);
nand U10027 (N_10027,N_9944,N_9810);
nand U10028 (N_10028,N_9592,N_9720);
or U10029 (N_10029,N_9775,N_9719);
and U10030 (N_10030,N_9959,N_9697);
and U10031 (N_10031,N_9922,N_9973);
and U10032 (N_10032,N_9883,N_9565);
nor U10033 (N_10033,N_9685,N_9954);
xor U10034 (N_10034,N_9645,N_9893);
xnor U10035 (N_10035,N_9620,N_9815);
nor U10036 (N_10036,N_9577,N_9951);
xnor U10037 (N_10037,N_9512,N_9859);
or U10038 (N_10038,N_9735,N_9511);
nand U10039 (N_10039,N_9597,N_9786);
nor U10040 (N_10040,N_9805,N_9779);
or U10041 (N_10041,N_9535,N_9982);
nand U10042 (N_10042,N_9516,N_9528);
or U10043 (N_10043,N_9534,N_9801);
and U10044 (N_10044,N_9552,N_9793);
nand U10045 (N_10045,N_9857,N_9763);
or U10046 (N_10046,N_9622,N_9837);
nand U10047 (N_10047,N_9776,N_9875);
or U10048 (N_10048,N_9828,N_9601);
or U10049 (N_10049,N_9822,N_9953);
or U10050 (N_10050,N_9966,N_9819);
or U10051 (N_10051,N_9896,N_9632);
nand U10052 (N_10052,N_9698,N_9785);
and U10053 (N_10053,N_9787,N_9940);
xor U10054 (N_10054,N_9509,N_9696);
xor U10055 (N_10055,N_9757,N_9758);
xor U10056 (N_10056,N_9553,N_9618);
xor U10057 (N_10057,N_9671,N_9501);
and U10058 (N_10058,N_9559,N_9996);
nand U10059 (N_10059,N_9835,N_9813);
xor U10060 (N_10060,N_9823,N_9574);
nand U10061 (N_10061,N_9617,N_9962);
nor U10062 (N_10062,N_9773,N_9906);
and U10063 (N_10063,N_9680,N_9731);
and U10064 (N_10064,N_9510,N_9566);
xnor U10065 (N_10065,N_9579,N_9584);
xnor U10066 (N_10066,N_9881,N_9960);
xor U10067 (N_10067,N_9599,N_9911);
and U10068 (N_10068,N_9556,N_9955);
or U10069 (N_10069,N_9563,N_9678);
or U10070 (N_10070,N_9935,N_9715);
nand U10071 (N_10071,N_9729,N_9796);
nor U10072 (N_10072,N_9961,N_9852);
nand U10073 (N_10073,N_9933,N_9652);
nor U10074 (N_10074,N_9604,N_9997);
and U10075 (N_10075,N_9877,N_9900);
nand U10076 (N_10076,N_9653,N_9783);
or U10077 (N_10077,N_9746,N_9537);
nor U10078 (N_10078,N_9658,N_9981);
or U10079 (N_10079,N_9513,N_9704);
nor U10080 (N_10080,N_9821,N_9505);
nor U10081 (N_10081,N_9798,N_9844);
nor U10082 (N_10082,N_9695,N_9865);
xnor U10083 (N_10083,N_9969,N_9915);
xor U10084 (N_10084,N_9555,N_9947);
and U10085 (N_10085,N_9762,N_9726);
and U10086 (N_10086,N_9521,N_9789);
nor U10087 (N_10087,N_9891,N_9856);
xnor U10088 (N_10088,N_9581,N_9722);
nand U10089 (N_10089,N_9612,N_9992);
xnor U10090 (N_10090,N_9629,N_9750);
xor U10091 (N_10091,N_9724,N_9721);
xor U10092 (N_10092,N_9921,N_9895);
xnor U10093 (N_10093,N_9864,N_9526);
nor U10094 (N_10094,N_9711,N_9790);
nand U10095 (N_10095,N_9978,N_9500);
nor U10096 (N_10096,N_9630,N_9792);
nand U10097 (N_10097,N_9656,N_9700);
and U10098 (N_10098,N_9541,N_9561);
nand U10099 (N_10099,N_9683,N_9761);
nand U10100 (N_10100,N_9917,N_9976);
nor U10101 (N_10101,N_9692,N_9707);
xor U10102 (N_10102,N_9972,N_9932);
and U10103 (N_10103,N_9841,N_9633);
nor U10104 (N_10104,N_9937,N_9910);
nor U10105 (N_10105,N_9585,N_9994);
or U10106 (N_10106,N_9980,N_9738);
or U10107 (N_10107,N_9826,N_9832);
nor U10108 (N_10108,N_9648,N_9672);
or U10109 (N_10109,N_9862,N_9654);
and U10110 (N_10110,N_9788,N_9710);
nand U10111 (N_10111,N_9502,N_9587);
nand U10112 (N_10112,N_9743,N_9703);
nand U10113 (N_10113,N_9941,N_9912);
or U10114 (N_10114,N_9839,N_9766);
nand U10115 (N_10115,N_9536,N_9918);
nand U10116 (N_10116,N_9811,N_9873);
or U10117 (N_10117,N_9755,N_9791);
nand U10118 (N_10118,N_9717,N_9665);
nand U10119 (N_10119,N_9963,N_9894);
and U10120 (N_10120,N_9855,N_9814);
or U10121 (N_10121,N_9770,N_9804);
and U10122 (N_10122,N_9540,N_9642);
and U10123 (N_10123,N_9795,N_9767);
nand U10124 (N_10124,N_9503,N_9999);
nand U10125 (N_10125,N_9754,N_9740);
and U10126 (N_10126,N_9799,N_9991);
nor U10127 (N_10127,N_9544,N_9908);
nor U10128 (N_10128,N_9573,N_9531);
and U10129 (N_10129,N_9925,N_9676);
nor U10130 (N_10130,N_9545,N_9718);
and U10131 (N_10131,N_9725,N_9551);
nand U10132 (N_10132,N_9903,N_9504);
nand U10133 (N_10133,N_9902,N_9733);
or U10134 (N_10134,N_9898,N_9807);
nor U10135 (N_10135,N_9651,N_9781);
and U10136 (N_10136,N_9570,N_9686);
xnor U10137 (N_10137,N_9831,N_9533);
xor U10138 (N_10138,N_9970,N_9675);
xnor U10139 (N_10139,N_9693,N_9634);
nand U10140 (N_10140,N_9927,N_9974);
nor U10141 (N_10141,N_9639,N_9749);
or U10142 (N_10142,N_9866,N_9560);
and U10143 (N_10143,N_9929,N_9986);
xnor U10144 (N_10144,N_9923,N_9655);
and U10145 (N_10145,N_9532,N_9641);
and U10146 (N_10146,N_9971,N_9548);
nand U10147 (N_10147,N_9774,N_9572);
and U10148 (N_10148,N_9514,N_9594);
or U10149 (N_10149,N_9674,N_9884);
or U10150 (N_10150,N_9945,N_9557);
xnor U10151 (N_10151,N_9694,N_9716);
xor U10152 (N_10152,N_9809,N_9619);
and U10153 (N_10153,N_9851,N_9708);
nand U10154 (N_10154,N_9625,N_9518);
nand U10155 (N_10155,N_9660,N_9878);
or U10156 (N_10156,N_9803,N_9712);
nor U10157 (N_10157,N_9946,N_9772);
nand U10158 (N_10158,N_9613,N_9863);
and U10159 (N_10159,N_9628,N_9664);
nor U10160 (N_10160,N_9580,N_9778);
xor U10161 (N_10161,N_9538,N_9668);
nand U10162 (N_10162,N_9930,N_9659);
xor U10163 (N_10163,N_9627,N_9993);
or U10164 (N_10164,N_9546,N_9600);
nor U10165 (N_10165,N_9956,N_9777);
xnor U10166 (N_10166,N_9598,N_9820);
and U10167 (N_10167,N_9780,N_9667);
xnor U10168 (N_10168,N_9596,N_9812);
and U10169 (N_10169,N_9568,N_9669);
nor U10170 (N_10170,N_9522,N_9964);
nand U10171 (N_10171,N_9760,N_9886);
and U10172 (N_10172,N_9666,N_9771);
nand U10173 (N_10173,N_9687,N_9952);
or U10174 (N_10174,N_9825,N_9769);
nand U10175 (N_10175,N_9913,N_9797);
xor U10176 (N_10176,N_9871,N_9690);
nand U10177 (N_10177,N_9723,N_9904);
xnor U10178 (N_10178,N_9759,N_9728);
or U10179 (N_10179,N_9752,N_9876);
nor U10180 (N_10180,N_9679,N_9934);
nand U10181 (N_10181,N_9924,N_9853);
and U10182 (N_10182,N_9849,N_9817);
xnor U10183 (N_10183,N_9987,N_9621);
nand U10184 (N_10184,N_9609,N_9764);
or U10185 (N_10185,N_9988,N_9836);
or U10186 (N_10186,N_9880,N_9990);
and U10187 (N_10187,N_9824,N_9688);
xnor U10188 (N_10188,N_9768,N_9879);
nor U10189 (N_10189,N_9586,N_9920);
and U10190 (N_10190,N_9644,N_9756);
nor U10191 (N_10191,N_9870,N_9564);
nand U10192 (N_10192,N_9714,N_9808);
nand U10193 (N_10193,N_9833,N_9529);
nand U10194 (N_10194,N_9968,N_9578);
xnor U10195 (N_10195,N_9948,N_9689);
and U10196 (N_10196,N_9858,N_9684);
xnor U10197 (N_10197,N_9614,N_9571);
and U10198 (N_10198,N_9701,N_9998);
and U10199 (N_10199,N_9591,N_9989);
or U10200 (N_10200,N_9637,N_9569);
xor U10201 (N_10201,N_9539,N_9682);
nand U10202 (N_10202,N_9842,N_9765);
or U10203 (N_10203,N_9975,N_9739);
nor U10204 (N_10204,N_9802,N_9887);
or U10205 (N_10205,N_9662,N_9649);
nor U10206 (N_10206,N_9736,N_9709);
xor U10207 (N_10207,N_9699,N_9984);
or U10208 (N_10208,N_9931,N_9753);
or U10209 (N_10209,N_9872,N_9995);
xor U10210 (N_10210,N_9562,N_9588);
xnor U10211 (N_10211,N_9806,N_9943);
xor U10212 (N_10212,N_9737,N_9890);
and U10213 (N_10213,N_9751,N_9602);
nor U10214 (N_10214,N_9914,N_9889);
nand U10215 (N_10215,N_9567,N_9661);
xnor U10216 (N_10216,N_9593,N_9515);
nor U10217 (N_10217,N_9530,N_9575);
xor U10218 (N_10218,N_9547,N_9519);
or U10219 (N_10219,N_9507,N_9727);
or U10220 (N_10220,N_9558,N_9734);
nand U10221 (N_10221,N_9623,N_9517);
nor U10222 (N_10222,N_9670,N_9646);
xnor U10223 (N_10223,N_9605,N_9663);
and U10224 (N_10224,N_9861,N_9845);
nor U10225 (N_10225,N_9967,N_9854);
or U10226 (N_10226,N_9834,N_9741);
nor U10227 (N_10227,N_9543,N_9784);
xnor U10228 (N_10228,N_9626,N_9691);
xnor U10229 (N_10229,N_9847,N_9949);
xnor U10230 (N_10230,N_9840,N_9782);
nor U10231 (N_10231,N_9950,N_9524);
nor U10232 (N_10232,N_9603,N_9983);
or U10233 (N_10233,N_9744,N_9647);
nor U10234 (N_10234,N_9542,N_9850);
and U10235 (N_10235,N_9705,N_9942);
or U10236 (N_10236,N_9576,N_9549);
nor U10237 (N_10237,N_9582,N_9794);
or U10238 (N_10238,N_9958,N_9938);
and U10239 (N_10239,N_9882,N_9677);
xnor U10240 (N_10240,N_9928,N_9520);
nand U10241 (N_10241,N_9640,N_9732);
xnor U10242 (N_10242,N_9818,N_9624);
xnor U10243 (N_10243,N_9713,N_9745);
or U10244 (N_10244,N_9901,N_9506);
nor U10245 (N_10245,N_9636,N_9843);
nor U10246 (N_10246,N_9838,N_9635);
xor U10247 (N_10247,N_9892,N_9615);
or U10248 (N_10248,N_9550,N_9523);
nor U10249 (N_10249,N_9583,N_9527);
and U10250 (N_10250,N_9689,N_9900);
nand U10251 (N_10251,N_9677,N_9647);
or U10252 (N_10252,N_9881,N_9599);
nand U10253 (N_10253,N_9778,N_9822);
xor U10254 (N_10254,N_9773,N_9673);
or U10255 (N_10255,N_9667,N_9714);
or U10256 (N_10256,N_9762,N_9535);
or U10257 (N_10257,N_9957,N_9559);
and U10258 (N_10258,N_9599,N_9507);
xor U10259 (N_10259,N_9774,N_9738);
xor U10260 (N_10260,N_9960,N_9540);
or U10261 (N_10261,N_9650,N_9869);
xnor U10262 (N_10262,N_9704,N_9947);
xor U10263 (N_10263,N_9958,N_9892);
xor U10264 (N_10264,N_9899,N_9961);
nor U10265 (N_10265,N_9899,N_9648);
nor U10266 (N_10266,N_9724,N_9594);
nor U10267 (N_10267,N_9976,N_9641);
xor U10268 (N_10268,N_9794,N_9619);
nand U10269 (N_10269,N_9857,N_9647);
or U10270 (N_10270,N_9547,N_9959);
or U10271 (N_10271,N_9822,N_9782);
nand U10272 (N_10272,N_9948,N_9744);
and U10273 (N_10273,N_9942,N_9982);
or U10274 (N_10274,N_9755,N_9565);
nand U10275 (N_10275,N_9959,N_9694);
and U10276 (N_10276,N_9851,N_9642);
nor U10277 (N_10277,N_9611,N_9958);
or U10278 (N_10278,N_9523,N_9694);
or U10279 (N_10279,N_9857,N_9943);
xor U10280 (N_10280,N_9504,N_9837);
xnor U10281 (N_10281,N_9666,N_9760);
or U10282 (N_10282,N_9517,N_9949);
nand U10283 (N_10283,N_9737,N_9986);
nor U10284 (N_10284,N_9904,N_9501);
nand U10285 (N_10285,N_9882,N_9904);
and U10286 (N_10286,N_9884,N_9772);
nand U10287 (N_10287,N_9583,N_9915);
xnor U10288 (N_10288,N_9505,N_9794);
nand U10289 (N_10289,N_9940,N_9741);
and U10290 (N_10290,N_9667,N_9817);
nand U10291 (N_10291,N_9810,N_9954);
nor U10292 (N_10292,N_9826,N_9891);
or U10293 (N_10293,N_9837,N_9712);
nor U10294 (N_10294,N_9744,N_9881);
and U10295 (N_10295,N_9671,N_9888);
or U10296 (N_10296,N_9553,N_9798);
nand U10297 (N_10297,N_9612,N_9924);
nor U10298 (N_10298,N_9639,N_9740);
or U10299 (N_10299,N_9561,N_9562);
nand U10300 (N_10300,N_9600,N_9758);
and U10301 (N_10301,N_9895,N_9938);
and U10302 (N_10302,N_9680,N_9663);
nor U10303 (N_10303,N_9765,N_9837);
nor U10304 (N_10304,N_9561,N_9522);
and U10305 (N_10305,N_9577,N_9700);
nor U10306 (N_10306,N_9575,N_9705);
nor U10307 (N_10307,N_9792,N_9526);
nor U10308 (N_10308,N_9606,N_9553);
nor U10309 (N_10309,N_9812,N_9963);
or U10310 (N_10310,N_9772,N_9660);
and U10311 (N_10311,N_9548,N_9536);
nand U10312 (N_10312,N_9541,N_9693);
nand U10313 (N_10313,N_9666,N_9673);
or U10314 (N_10314,N_9785,N_9700);
xor U10315 (N_10315,N_9524,N_9653);
xnor U10316 (N_10316,N_9756,N_9742);
or U10317 (N_10317,N_9996,N_9525);
and U10318 (N_10318,N_9984,N_9538);
nand U10319 (N_10319,N_9831,N_9701);
nand U10320 (N_10320,N_9887,N_9799);
or U10321 (N_10321,N_9584,N_9958);
nand U10322 (N_10322,N_9974,N_9816);
and U10323 (N_10323,N_9504,N_9802);
or U10324 (N_10324,N_9944,N_9885);
nor U10325 (N_10325,N_9738,N_9849);
or U10326 (N_10326,N_9519,N_9505);
xnor U10327 (N_10327,N_9879,N_9626);
and U10328 (N_10328,N_9658,N_9640);
nand U10329 (N_10329,N_9696,N_9949);
or U10330 (N_10330,N_9860,N_9809);
nor U10331 (N_10331,N_9938,N_9623);
or U10332 (N_10332,N_9864,N_9940);
nand U10333 (N_10333,N_9831,N_9708);
or U10334 (N_10334,N_9804,N_9936);
xnor U10335 (N_10335,N_9867,N_9973);
nor U10336 (N_10336,N_9926,N_9564);
or U10337 (N_10337,N_9589,N_9660);
xor U10338 (N_10338,N_9766,N_9593);
and U10339 (N_10339,N_9763,N_9621);
or U10340 (N_10340,N_9851,N_9586);
nor U10341 (N_10341,N_9527,N_9941);
xor U10342 (N_10342,N_9916,N_9662);
nor U10343 (N_10343,N_9634,N_9531);
xnor U10344 (N_10344,N_9938,N_9905);
nor U10345 (N_10345,N_9710,N_9523);
or U10346 (N_10346,N_9823,N_9757);
or U10347 (N_10347,N_9876,N_9516);
nand U10348 (N_10348,N_9671,N_9573);
xnor U10349 (N_10349,N_9946,N_9691);
or U10350 (N_10350,N_9574,N_9783);
nand U10351 (N_10351,N_9533,N_9791);
nand U10352 (N_10352,N_9555,N_9739);
nand U10353 (N_10353,N_9759,N_9791);
nand U10354 (N_10354,N_9682,N_9665);
xor U10355 (N_10355,N_9791,N_9722);
or U10356 (N_10356,N_9998,N_9518);
xnor U10357 (N_10357,N_9983,N_9856);
and U10358 (N_10358,N_9876,N_9732);
xor U10359 (N_10359,N_9791,N_9972);
nor U10360 (N_10360,N_9752,N_9672);
nor U10361 (N_10361,N_9677,N_9874);
xnor U10362 (N_10362,N_9741,N_9794);
xor U10363 (N_10363,N_9755,N_9745);
and U10364 (N_10364,N_9519,N_9869);
and U10365 (N_10365,N_9756,N_9734);
nor U10366 (N_10366,N_9579,N_9799);
nand U10367 (N_10367,N_9808,N_9648);
xor U10368 (N_10368,N_9959,N_9704);
and U10369 (N_10369,N_9699,N_9760);
and U10370 (N_10370,N_9873,N_9985);
or U10371 (N_10371,N_9633,N_9815);
and U10372 (N_10372,N_9801,N_9935);
or U10373 (N_10373,N_9727,N_9900);
xor U10374 (N_10374,N_9805,N_9981);
nand U10375 (N_10375,N_9600,N_9537);
xor U10376 (N_10376,N_9501,N_9787);
or U10377 (N_10377,N_9882,N_9694);
xnor U10378 (N_10378,N_9950,N_9912);
and U10379 (N_10379,N_9994,N_9815);
xor U10380 (N_10380,N_9949,N_9931);
nand U10381 (N_10381,N_9872,N_9867);
or U10382 (N_10382,N_9693,N_9758);
and U10383 (N_10383,N_9506,N_9803);
and U10384 (N_10384,N_9518,N_9720);
xor U10385 (N_10385,N_9926,N_9825);
and U10386 (N_10386,N_9549,N_9638);
nor U10387 (N_10387,N_9508,N_9806);
nand U10388 (N_10388,N_9653,N_9687);
nor U10389 (N_10389,N_9910,N_9891);
xnor U10390 (N_10390,N_9657,N_9501);
xnor U10391 (N_10391,N_9635,N_9802);
and U10392 (N_10392,N_9790,N_9510);
nand U10393 (N_10393,N_9988,N_9705);
and U10394 (N_10394,N_9506,N_9637);
xnor U10395 (N_10395,N_9806,N_9642);
nand U10396 (N_10396,N_9660,N_9627);
xnor U10397 (N_10397,N_9771,N_9531);
xnor U10398 (N_10398,N_9604,N_9686);
nor U10399 (N_10399,N_9818,N_9844);
and U10400 (N_10400,N_9811,N_9769);
nand U10401 (N_10401,N_9553,N_9772);
nand U10402 (N_10402,N_9632,N_9563);
or U10403 (N_10403,N_9527,N_9968);
xnor U10404 (N_10404,N_9779,N_9968);
nand U10405 (N_10405,N_9817,N_9758);
or U10406 (N_10406,N_9888,N_9803);
xor U10407 (N_10407,N_9591,N_9823);
nand U10408 (N_10408,N_9749,N_9556);
nand U10409 (N_10409,N_9861,N_9739);
nor U10410 (N_10410,N_9927,N_9651);
nand U10411 (N_10411,N_9996,N_9781);
nor U10412 (N_10412,N_9668,N_9523);
xnor U10413 (N_10413,N_9944,N_9844);
nand U10414 (N_10414,N_9941,N_9891);
nor U10415 (N_10415,N_9500,N_9633);
nor U10416 (N_10416,N_9748,N_9902);
nor U10417 (N_10417,N_9678,N_9714);
or U10418 (N_10418,N_9688,N_9793);
or U10419 (N_10419,N_9686,N_9872);
xnor U10420 (N_10420,N_9956,N_9609);
xor U10421 (N_10421,N_9976,N_9566);
and U10422 (N_10422,N_9659,N_9708);
nor U10423 (N_10423,N_9614,N_9641);
xor U10424 (N_10424,N_9853,N_9724);
xnor U10425 (N_10425,N_9846,N_9590);
nor U10426 (N_10426,N_9768,N_9554);
nand U10427 (N_10427,N_9632,N_9653);
and U10428 (N_10428,N_9644,N_9696);
nor U10429 (N_10429,N_9953,N_9760);
nand U10430 (N_10430,N_9712,N_9844);
or U10431 (N_10431,N_9510,N_9679);
or U10432 (N_10432,N_9989,N_9832);
or U10433 (N_10433,N_9795,N_9566);
nor U10434 (N_10434,N_9517,N_9595);
xnor U10435 (N_10435,N_9776,N_9695);
nor U10436 (N_10436,N_9745,N_9565);
nor U10437 (N_10437,N_9541,N_9883);
nand U10438 (N_10438,N_9845,N_9700);
xnor U10439 (N_10439,N_9701,N_9922);
xnor U10440 (N_10440,N_9923,N_9922);
nand U10441 (N_10441,N_9649,N_9781);
nand U10442 (N_10442,N_9852,N_9672);
or U10443 (N_10443,N_9578,N_9774);
nand U10444 (N_10444,N_9893,N_9825);
and U10445 (N_10445,N_9542,N_9780);
or U10446 (N_10446,N_9737,N_9535);
xnor U10447 (N_10447,N_9761,N_9691);
xnor U10448 (N_10448,N_9833,N_9697);
xor U10449 (N_10449,N_9780,N_9682);
nand U10450 (N_10450,N_9611,N_9749);
and U10451 (N_10451,N_9632,N_9959);
xor U10452 (N_10452,N_9533,N_9977);
nand U10453 (N_10453,N_9792,N_9840);
and U10454 (N_10454,N_9846,N_9528);
nor U10455 (N_10455,N_9582,N_9886);
nand U10456 (N_10456,N_9682,N_9853);
xor U10457 (N_10457,N_9954,N_9990);
nand U10458 (N_10458,N_9639,N_9686);
nand U10459 (N_10459,N_9666,N_9639);
nor U10460 (N_10460,N_9760,N_9752);
xnor U10461 (N_10461,N_9905,N_9573);
nor U10462 (N_10462,N_9534,N_9827);
nor U10463 (N_10463,N_9829,N_9986);
or U10464 (N_10464,N_9861,N_9791);
nor U10465 (N_10465,N_9523,N_9530);
and U10466 (N_10466,N_9583,N_9872);
and U10467 (N_10467,N_9810,N_9526);
or U10468 (N_10468,N_9641,N_9543);
nand U10469 (N_10469,N_9716,N_9772);
or U10470 (N_10470,N_9743,N_9820);
and U10471 (N_10471,N_9823,N_9588);
nor U10472 (N_10472,N_9765,N_9809);
xnor U10473 (N_10473,N_9890,N_9758);
or U10474 (N_10474,N_9976,N_9956);
nor U10475 (N_10475,N_9738,N_9792);
nand U10476 (N_10476,N_9606,N_9978);
nand U10477 (N_10477,N_9850,N_9711);
nor U10478 (N_10478,N_9511,N_9784);
and U10479 (N_10479,N_9901,N_9950);
nor U10480 (N_10480,N_9607,N_9977);
nand U10481 (N_10481,N_9683,N_9876);
xnor U10482 (N_10482,N_9914,N_9794);
nor U10483 (N_10483,N_9712,N_9648);
and U10484 (N_10484,N_9851,N_9687);
or U10485 (N_10485,N_9941,N_9740);
and U10486 (N_10486,N_9952,N_9590);
nand U10487 (N_10487,N_9998,N_9779);
xor U10488 (N_10488,N_9568,N_9896);
and U10489 (N_10489,N_9877,N_9883);
and U10490 (N_10490,N_9905,N_9720);
and U10491 (N_10491,N_9978,N_9758);
nor U10492 (N_10492,N_9801,N_9578);
nand U10493 (N_10493,N_9612,N_9622);
nor U10494 (N_10494,N_9844,N_9830);
nor U10495 (N_10495,N_9724,N_9733);
xnor U10496 (N_10496,N_9529,N_9839);
nor U10497 (N_10497,N_9553,N_9610);
or U10498 (N_10498,N_9934,N_9613);
nand U10499 (N_10499,N_9970,N_9661);
xor U10500 (N_10500,N_10417,N_10271);
or U10501 (N_10501,N_10085,N_10088);
nand U10502 (N_10502,N_10148,N_10495);
nand U10503 (N_10503,N_10469,N_10489);
and U10504 (N_10504,N_10346,N_10114);
xor U10505 (N_10505,N_10118,N_10139);
nor U10506 (N_10506,N_10215,N_10020);
or U10507 (N_10507,N_10479,N_10392);
xnor U10508 (N_10508,N_10269,N_10299);
nor U10509 (N_10509,N_10437,N_10099);
nor U10510 (N_10510,N_10446,N_10157);
and U10511 (N_10511,N_10044,N_10352);
xnor U10512 (N_10512,N_10096,N_10001);
and U10513 (N_10513,N_10339,N_10310);
or U10514 (N_10514,N_10292,N_10401);
xnor U10515 (N_10515,N_10094,N_10104);
nor U10516 (N_10516,N_10187,N_10427);
nor U10517 (N_10517,N_10337,N_10270);
nand U10518 (N_10518,N_10325,N_10230);
nor U10519 (N_10519,N_10426,N_10361);
and U10520 (N_10520,N_10138,N_10472);
nand U10521 (N_10521,N_10209,N_10405);
nor U10522 (N_10522,N_10009,N_10467);
or U10523 (N_10523,N_10212,N_10123);
nor U10524 (N_10524,N_10057,N_10155);
and U10525 (N_10525,N_10025,N_10314);
xor U10526 (N_10526,N_10394,N_10181);
xor U10527 (N_10527,N_10254,N_10186);
or U10528 (N_10528,N_10082,N_10222);
nand U10529 (N_10529,N_10399,N_10201);
nor U10530 (N_10530,N_10093,N_10216);
nand U10531 (N_10531,N_10203,N_10326);
nor U10532 (N_10532,N_10443,N_10423);
nor U10533 (N_10533,N_10047,N_10288);
and U10534 (N_10534,N_10317,N_10006);
nand U10535 (N_10535,N_10459,N_10294);
nand U10536 (N_10536,N_10413,N_10162);
nor U10537 (N_10537,N_10341,N_10109);
xor U10538 (N_10538,N_10493,N_10452);
xnor U10539 (N_10539,N_10062,N_10355);
or U10540 (N_10540,N_10046,N_10349);
nor U10541 (N_10541,N_10257,N_10244);
xor U10542 (N_10542,N_10362,N_10435);
nand U10543 (N_10543,N_10280,N_10211);
or U10544 (N_10544,N_10455,N_10131);
xor U10545 (N_10545,N_10466,N_10195);
nand U10546 (N_10546,N_10327,N_10028);
nand U10547 (N_10547,N_10272,N_10053);
xor U10548 (N_10548,N_10330,N_10070);
and U10549 (N_10549,N_10385,N_10408);
or U10550 (N_10550,N_10185,N_10389);
and U10551 (N_10551,N_10482,N_10438);
nand U10552 (N_10552,N_10322,N_10285);
nand U10553 (N_10553,N_10376,N_10007);
nand U10554 (N_10554,N_10125,N_10273);
xnor U10555 (N_10555,N_10089,N_10372);
xor U10556 (N_10556,N_10188,N_10253);
and U10557 (N_10557,N_10412,N_10226);
xnor U10558 (N_10558,N_10112,N_10370);
xnor U10559 (N_10559,N_10040,N_10160);
nor U10560 (N_10560,N_10237,N_10180);
and U10561 (N_10561,N_10431,N_10301);
nand U10562 (N_10562,N_10205,N_10276);
and U10563 (N_10563,N_10079,N_10225);
nand U10564 (N_10564,N_10286,N_10266);
or U10565 (N_10565,N_10054,N_10419);
and U10566 (N_10566,N_10060,N_10086);
nor U10567 (N_10567,N_10458,N_10202);
or U10568 (N_10568,N_10154,N_10039);
nand U10569 (N_10569,N_10245,N_10307);
xnor U10570 (N_10570,N_10281,N_10196);
nor U10571 (N_10571,N_10116,N_10277);
nand U10572 (N_10572,N_10061,N_10134);
nand U10573 (N_10573,N_10439,N_10456);
nand U10574 (N_10574,N_10013,N_10130);
and U10575 (N_10575,N_10179,N_10045);
nor U10576 (N_10576,N_10393,N_10476);
or U10577 (N_10577,N_10074,N_10477);
or U10578 (N_10578,N_10016,N_10219);
xor U10579 (N_10579,N_10305,N_10197);
xnor U10580 (N_10580,N_10316,N_10142);
nand U10581 (N_10581,N_10059,N_10350);
xnor U10582 (N_10582,N_10158,N_10071);
or U10583 (N_10583,N_10019,N_10003);
xor U10584 (N_10584,N_10300,N_10256);
nand U10585 (N_10585,N_10425,N_10066);
and U10586 (N_10586,N_10144,N_10081);
nand U10587 (N_10587,N_10106,N_10296);
nand U10588 (N_10588,N_10255,N_10461);
xor U10589 (N_10589,N_10097,N_10382);
and U10590 (N_10590,N_10000,N_10008);
nor U10591 (N_10591,N_10132,N_10429);
xnor U10592 (N_10592,N_10369,N_10119);
nand U10593 (N_10593,N_10463,N_10208);
nor U10594 (N_10594,N_10191,N_10032);
or U10595 (N_10595,N_10448,N_10491);
xor U10596 (N_10596,N_10166,N_10036);
nand U10597 (N_10597,N_10414,N_10178);
nor U10598 (N_10598,N_10051,N_10150);
nand U10599 (N_10599,N_10430,N_10284);
nand U10600 (N_10600,N_10340,N_10497);
or U10601 (N_10601,N_10387,N_10147);
nand U10602 (N_10602,N_10121,N_10395);
xnor U10603 (N_10603,N_10090,N_10034);
nand U10604 (N_10604,N_10368,N_10083);
xor U10605 (N_10605,N_10265,N_10453);
nand U10606 (N_10606,N_10484,N_10258);
nor U10607 (N_10607,N_10014,N_10236);
or U10608 (N_10608,N_10231,N_10092);
nor U10609 (N_10609,N_10274,N_10328);
and U10610 (N_10610,N_10353,N_10383);
nand U10611 (N_10611,N_10320,N_10210);
nand U10612 (N_10612,N_10037,N_10363);
nand U10613 (N_10613,N_10329,N_10483);
or U10614 (N_10614,N_10168,N_10367);
nand U10615 (N_10615,N_10137,N_10073);
nor U10616 (N_10616,N_10403,N_10335);
and U10617 (N_10617,N_10105,N_10224);
nor U10618 (N_10618,N_10026,N_10315);
or U10619 (N_10619,N_10145,N_10240);
xnor U10620 (N_10620,N_10379,N_10342);
xor U10621 (N_10621,N_10289,N_10029);
and U10622 (N_10622,N_10441,N_10371);
and U10623 (N_10623,N_10422,N_10141);
nor U10624 (N_10624,N_10420,N_10193);
nor U10625 (N_10625,N_10323,N_10129);
nor U10626 (N_10626,N_10103,N_10449);
nand U10627 (N_10627,N_10149,N_10033);
nand U10628 (N_10628,N_10424,N_10217);
and U10629 (N_10629,N_10264,N_10474);
xnor U10630 (N_10630,N_10357,N_10199);
xnor U10631 (N_10631,N_10220,N_10331);
or U10632 (N_10632,N_10391,N_10133);
or U10633 (N_10633,N_10221,N_10100);
nand U10634 (N_10634,N_10238,N_10189);
xor U10635 (N_10635,N_10135,N_10293);
or U10636 (N_10636,N_10072,N_10041);
nand U10637 (N_10637,N_10485,N_10080);
nor U10638 (N_10638,N_10246,N_10251);
nor U10639 (N_10639,N_10428,N_10445);
and U10640 (N_10640,N_10462,N_10023);
and U10641 (N_10641,N_10140,N_10295);
and U10642 (N_10642,N_10063,N_10283);
and U10643 (N_10643,N_10214,N_10321);
nand U10644 (N_10644,N_10468,N_10067);
xnor U10645 (N_10645,N_10113,N_10184);
or U10646 (N_10646,N_10402,N_10465);
xnor U10647 (N_10647,N_10303,N_10398);
and U10648 (N_10648,N_10291,N_10318);
nand U10649 (N_10649,N_10262,N_10388);
and U10650 (N_10650,N_10290,N_10332);
or U10651 (N_10651,N_10002,N_10374);
nor U10652 (N_10652,N_10111,N_10043);
nand U10653 (N_10653,N_10030,N_10260);
nor U10654 (N_10654,N_10267,N_10304);
nand U10655 (N_10655,N_10249,N_10409);
nor U10656 (N_10656,N_10364,N_10415);
nor U10657 (N_10657,N_10015,N_10234);
or U10658 (N_10658,N_10297,N_10171);
nor U10659 (N_10659,N_10464,N_10451);
nand U10660 (N_10660,N_10263,N_10200);
nor U10661 (N_10661,N_10242,N_10207);
nor U10662 (N_10662,N_10194,N_10259);
nor U10663 (N_10663,N_10319,N_10174);
xnor U10664 (N_10664,N_10136,N_10351);
and U10665 (N_10665,N_10470,N_10400);
xor U10666 (N_10666,N_10486,N_10488);
nand U10667 (N_10667,N_10377,N_10359);
xor U10668 (N_10668,N_10024,N_10365);
nor U10669 (N_10669,N_10078,N_10334);
nor U10670 (N_10670,N_10475,N_10473);
nor U10671 (N_10671,N_10213,N_10324);
or U10672 (N_10672,N_10447,N_10027);
and U10673 (N_10673,N_10165,N_10192);
or U10674 (N_10674,N_10248,N_10287);
and U10675 (N_10675,N_10042,N_10161);
nor U10676 (N_10676,N_10065,N_10252);
nor U10677 (N_10677,N_10011,N_10309);
xor U10678 (N_10678,N_10356,N_10115);
nand U10679 (N_10679,N_10152,N_10373);
and U10680 (N_10680,N_10153,N_10480);
and U10681 (N_10681,N_10492,N_10250);
and U10682 (N_10682,N_10124,N_10035);
nor U10683 (N_10683,N_10390,N_10436);
nand U10684 (N_10684,N_10095,N_10416);
and U10685 (N_10685,N_10375,N_10360);
nor U10686 (N_10686,N_10167,N_10010);
or U10687 (N_10687,N_10075,N_10204);
xnor U10688 (N_10688,N_10418,N_10017);
nor U10689 (N_10689,N_10345,N_10055);
nand U10690 (N_10690,N_10173,N_10247);
nand U10691 (N_10691,N_10396,N_10235);
and U10692 (N_10692,N_10454,N_10440);
and U10693 (N_10693,N_10022,N_10442);
xor U10694 (N_10694,N_10498,N_10170);
nand U10695 (N_10695,N_10198,N_10049);
and U10696 (N_10696,N_10050,N_10223);
and U10697 (N_10697,N_10313,N_10278);
xor U10698 (N_10698,N_10261,N_10084);
nor U10699 (N_10699,N_10176,N_10146);
or U10700 (N_10700,N_10478,N_10298);
nor U10701 (N_10701,N_10433,N_10312);
and U10702 (N_10702,N_10005,N_10122);
xor U10703 (N_10703,N_10243,N_10381);
nand U10704 (N_10704,N_10183,N_10336);
xor U10705 (N_10705,N_10275,N_10333);
xnor U10706 (N_10706,N_10126,N_10499);
xor U10707 (N_10707,N_10064,N_10163);
nand U10708 (N_10708,N_10076,N_10120);
or U10709 (N_10709,N_10233,N_10172);
xnor U10710 (N_10710,N_10229,N_10159);
nor U10711 (N_10711,N_10338,N_10175);
nand U10712 (N_10712,N_10117,N_10102);
nand U10713 (N_10713,N_10490,N_10241);
and U10714 (N_10714,N_10177,N_10282);
and U10715 (N_10715,N_10411,N_10206);
nand U10716 (N_10716,N_10487,N_10457);
and U10717 (N_10717,N_10410,N_10471);
or U10718 (N_10718,N_10306,N_10496);
and U10719 (N_10719,N_10107,N_10004);
nand U10720 (N_10720,N_10308,N_10397);
nor U10721 (N_10721,N_10380,N_10384);
nor U10722 (N_10722,N_10151,N_10021);
nand U10723 (N_10723,N_10077,N_10228);
xnor U10724 (N_10724,N_10378,N_10421);
or U10725 (N_10725,N_10038,N_10108);
nand U10726 (N_10726,N_10347,N_10450);
nor U10727 (N_10727,N_10087,N_10012);
nor U10728 (N_10728,N_10460,N_10343);
nor U10729 (N_10729,N_10358,N_10406);
nand U10730 (N_10730,N_10190,N_10127);
nor U10731 (N_10731,N_10018,N_10348);
nand U10732 (N_10732,N_10386,N_10239);
or U10733 (N_10733,N_10068,N_10366);
nor U10734 (N_10734,N_10101,N_10279);
and U10735 (N_10735,N_10218,N_10494);
xnor U10736 (N_10736,N_10354,N_10434);
nand U10737 (N_10737,N_10232,N_10481);
and U10738 (N_10738,N_10091,N_10227);
nand U10739 (N_10739,N_10069,N_10031);
or U10740 (N_10740,N_10169,N_10128);
and U10741 (N_10741,N_10268,N_10056);
nor U10742 (N_10742,N_10110,N_10182);
and U10743 (N_10743,N_10098,N_10407);
xnor U10744 (N_10744,N_10143,N_10444);
nand U10745 (N_10745,N_10344,N_10048);
nand U10746 (N_10746,N_10432,N_10164);
and U10747 (N_10747,N_10311,N_10156);
nand U10748 (N_10748,N_10404,N_10058);
nand U10749 (N_10749,N_10052,N_10302);
or U10750 (N_10750,N_10480,N_10414);
nand U10751 (N_10751,N_10005,N_10095);
xor U10752 (N_10752,N_10371,N_10295);
or U10753 (N_10753,N_10304,N_10234);
or U10754 (N_10754,N_10414,N_10202);
or U10755 (N_10755,N_10116,N_10359);
or U10756 (N_10756,N_10146,N_10024);
or U10757 (N_10757,N_10222,N_10306);
nand U10758 (N_10758,N_10468,N_10338);
or U10759 (N_10759,N_10237,N_10326);
nor U10760 (N_10760,N_10165,N_10155);
xor U10761 (N_10761,N_10495,N_10196);
xor U10762 (N_10762,N_10451,N_10273);
or U10763 (N_10763,N_10323,N_10459);
nand U10764 (N_10764,N_10425,N_10453);
and U10765 (N_10765,N_10406,N_10465);
xor U10766 (N_10766,N_10130,N_10270);
or U10767 (N_10767,N_10005,N_10039);
xor U10768 (N_10768,N_10275,N_10140);
nand U10769 (N_10769,N_10209,N_10439);
nand U10770 (N_10770,N_10388,N_10258);
or U10771 (N_10771,N_10278,N_10460);
or U10772 (N_10772,N_10128,N_10478);
nor U10773 (N_10773,N_10307,N_10152);
nor U10774 (N_10774,N_10240,N_10348);
nand U10775 (N_10775,N_10472,N_10289);
and U10776 (N_10776,N_10265,N_10474);
nor U10777 (N_10777,N_10281,N_10356);
and U10778 (N_10778,N_10059,N_10459);
or U10779 (N_10779,N_10019,N_10481);
xnor U10780 (N_10780,N_10249,N_10049);
xor U10781 (N_10781,N_10182,N_10267);
or U10782 (N_10782,N_10150,N_10011);
nand U10783 (N_10783,N_10026,N_10348);
and U10784 (N_10784,N_10191,N_10259);
nor U10785 (N_10785,N_10089,N_10071);
or U10786 (N_10786,N_10122,N_10195);
and U10787 (N_10787,N_10231,N_10222);
nor U10788 (N_10788,N_10017,N_10279);
or U10789 (N_10789,N_10108,N_10327);
xnor U10790 (N_10790,N_10286,N_10243);
nor U10791 (N_10791,N_10244,N_10446);
xor U10792 (N_10792,N_10154,N_10099);
xnor U10793 (N_10793,N_10358,N_10464);
and U10794 (N_10794,N_10012,N_10367);
nor U10795 (N_10795,N_10427,N_10460);
and U10796 (N_10796,N_10365,N_10401);
or U10797 (N_10797,N_10432,N_10348);
nand U10798 (N_10798,N_10421,N_10064);
xnor U10799 (N_10799,N_10165,N_10326);
xor U10800 (N_10800,N_10056,N_10179);
xor U10801 (N_10801,N_10206,N_10216);
or U10802 (N_10802,N_10102,N_10126);
nand U10803 (N_10803,N_10494,N_10035);
xor U10804 (N_10804,N_10120,N_10469);
xnor U10805 (N_10805,N_10318,N_10269);
and U10806 (N_10806,N_10307,N_10368);
and U10807 (N_10807,N_10396,N_10085);
and U10808 (N_10808,N_10104,N_10343);
and U10809 (N_10809,N_10092,N_10181);
nor U10810 (N_10810,N_10143,N_10419);
or U10811 (N_10811,N_10412,N_10403);
or U10812 (N_10812,N_10339,N_10093);
and U10813 (N_10813,N_10152,N_10167);
nand U10814 (N_10814,N_10401,N_10273);
nand U10815 (N_10815,N_10200,N_10264);
xnor U10816 (N_10816,N_10375,N_10192);
xnor U10817 (N_10817,N_10240,N_10080);
nand U10818 (N_10818,N_10032,N_10198);
and U10819 (N_10819,N_10257,N_10234);
or U10820 (N_10820,N_10209,N_10397);
xor U10821 (N_10821,N_10070,N_10014);
nand U10822 (N_10822,N_10045,N_10296);
and U10823 (N_10823,N_10411,N_10310);
and U10824 (N_10824,N_10254,N_10041);
or U10825 (N_10825,N_10221,N_10177);
xnor U10826 (N_10826,N_10029,N_10372);
xnor U10827 (N_10827,N_10434,N_10085);
and U10828 (N_10828,N_10437,N_10445);
nand U10829 (N_10829,N_10463,N_10405);
and U10830 (N_10830,N_10145,N_10071);
xnor U10831 (N_10831,N_10447,N_10300);
nor U10832 (N_10832,N_10371,N_10123);
xnor U10833 (N_10833,N_10429,N_10322);
xnor U10834 (N_10834,N_10306,N_10157);
xor U10835 (N_10835,N_10364,N_10351);
and U10836 (N_10836,N_10367,N_10094);
nor U10837 (N_10837,N_10201,N_10117);
or U10838 (N_10838,N_10499,N_10304);
or U10839 (N_10839,N_10170,N_10294);
xor U10840 (N_10840,N_10189,N_10217);
and U10841 (N_10841,N_10217,N_10264);
xnor U10842 (N_10842,N_10437,N_10134);
and U10843 (N_10843,N_10284,N_10446);
nand U10844 (N_10844,N_10023,N_10435);
xnor U10845 (N_10845,N_10348,N_10032);
or U10846 (N_10846,N_10122,N_10497);
or U10847 (N_10847,N_10212,N_10204);
or U10848 (N_10848,N_10273,N_10082);
nor U10849 (N_10849,N_10476,N_10316);
and U10850 (N_10850,N_10226,N_10161);
xor U10851 (N_10851,N_10441,N_10339);
nand U10852 (N_10852,N_10298,N_10442);
and U10853 (N_10853,N_10405,N_10205);
nor U10854 (N_10854,N_10486,N_10091);
and U10855 (N_10855,N_10466,N_10125);
xnor U10856 (N_10856,N_10204,N_10264);
and U10857 (N_10857,N_10319,N_10150);
xor U10858 (N_10858,N_10460,N_10231);
nand U10859 (N_10859,N_10442,N_10219);
or U10860 (N_10860,N_10124,N_10377);
or U10861 (N_10861,N_10364,N_10329);
or U10862 (N_10862,N_10396,N_10354);
nor U10863 (N_10863,N_10221,N_10363);
or U10864 (N_10864,N_10071,N_10189);
or U10865 (N_10865,N_10097,N_10381);
nand U10866 (N_10866,N_10320,N_10163);
and U10867 (N_10867,N_10090,N_10392);
xnor U10868 (N_10868,N_10293,N_10123);
nand U10869 (N_10869,N_10029,N_10165);
nand U10870 (N_10870,N_10233,N_10132);
or U10871 (N_10871,N_10355,N_10016);
nor U10872 (N_10872,N_10378,N_10454);
or U10873 (N_10873,N_10008,N_10046);
nand U10874 (N_10874,N_10348,N_10224);
nand U10875 (N_10875,N_10239,N_10260);
xnor U10876 (N_10876,N_10346,N_10187);
and U10877 (N_10877,N_10009,N_10369);
and U10878 (N_10878,N_10432,N_10201);
nor U10879 (N_10879,N_10263,N_10431);
nor U10880 (N_10880,N_10452,N_10471);
or U10881 (N_10881,N_10341,N_10027);
and U10882 (N_10882,N_10167,N_10029);
and U10883 (N_10883,N_10010,N_10434);
nor U10884 (N_10884,N_10113,N_10194);
and U10885 (N_10885,N_10104,N_10444);
and U10886 (N_10886,N_10429,N_10308);
nor U10887 (N_10887,N_10144,N_10487);
nand U10888 (N_10888,N_10364,N_10035);
xor U10889 (N_10889,N_10182,N_10424);
nand U10890 (N_10890,N_10371,N_10160);
or U10891 (N_10891,N_10131,N_10098);
nor U10892 (N_10892,N_10084,N_10071);
or U10893 (N_10893,N_10117,N_10227);
and U10894 (N_10894,N_10272,N_10159);
xor U10895 (N_10895,N_10347,N_10344);
nor U10896 (N_10896,N_10323,N_10208);
and U10897 (N_10897,N_10414,N_10411);
or U10898 (N_10898,N_10465,N_10044);
xor U10899 (N_10899,N_10454,N_10463);
nand U10900 (N_10900,N_10368,N_10249);
nor U10901 (N_10901,N_10009,N_10111);
nand U10902 (N_10902,N_10214,N_10397);
xnor U10903 (N_10903,N_10063,N_10149);
nor U10904 (N_10904,N_10009,N_10165);
xnor U10905 (N_10905,N_10387,N_10299);
nor U10906 (N_10906,N_10026,N_10228);
or U10907 (N_10907,N_10004,N_10340);
nor U10908 (N_10908,N_10083,N_10434);
xor U10909 (N_10909,N_10273,N_10480);
nor U10910 (N_10910,N_10274,N_10087);
and U10911 (N_10911,N_10048,N_10091);
or U10912 (N_10912,N_10146,N_10350);
nand U10913 (N_10913,N_10097,N_10261);
and U10914 (N_10914,N_10483,N_10492);
nand U10915 (N_10915,N_10328,N_10127);
nor U10916 (N_10916,N_10377,N_10429);
nor U10917 (N_10917,N_10244,N_10015);
nor U10918 (N_10918,N_10153,N_10092);
or U10919 (N_10919,N_10252,N_10133);
and U10920 (N_10920,N_10272,N_10313);
xnor U10921 (N_10921,N_10483,N_10142);
nand U10922 (N_10922,N_10147,N_10360);
nor U10923 (N_10923,N_10297,N_10411);
or U10924 (N_10924,N_10205,N_10196);
or U10925 (N_10925,N_10440,N_10398);
xnor U10926 (N_10926,N_10164,N_10470);
or U10927 (N_10927,N_10227,N_10328);
nor U10928 (N_10928,N_10117,N_10467);
nand U10929 (N_10929,N_10188,N_10332);
nor U10930 (N_10930,N_10287,N_10110);
or U10931 (N_10931,N_10115,N_10460);
xnor U10932 (N_10932,N_10263,N_10110);
nor U10933 (N_10933,N_10163,N_10246);
and U10934 (N_10934,N_10106,N_10186);
nor U10935 (N_10935,N_10343,N_10434);
or U10936 (N_10936,N_10350,N_10128);
xnor U10937 (N_10937,N_10252,N_10413);
nor U10938 (N_10938,N_10097,N_10423);
or U10939 (N_10939,N_10084,N_10065);
nor U10940 (N_10940,N_10306,N_10247);
or U10941 (N_10941,N_10075,N_10303);
and U10942 (N_10942,N_10199,N_10035);
nand U10943 (N_10943,N_10386,N_10275);
nand U10944 (N_10944,N_10045,N_10155);
nand U10945 (N_10945,N_10221,N_10059);
nor U10946 (N_10946,N_10418,N_10411);
or U10947 (N_10947,N_10148,N_10449);
and U10948 (N_10948,N_10223,N_10212);
or U10949 (N_10949,N_10497,N_10284);
and U10950 (N_10950,N_10070,N_10155);
nor U10951 (N_10951,N_10239,N_10428);
nand U10952 (N_10952,N_10068,N_10415);
xor U10953 (N_10953,N_10308,N_10326);
and U10954 (N_10954,N_10002,N_10413);
and U10955 (N_10955,N_10033,N_10326);
or U10956 (N_10956,N_10316,N_10393);
and U10957 (N_10957,N_10203,N_10452);
xor U10958 (N_10958,N_10288,N_10090);
and U10959 (N_10959,N_10106,N_10200);
nand U10960 (N_10960,N_10307,N_10008);
xor U10961 (N_10961,N_10334,N_10470);
and U10962 (N_10962,N_10430,N_10415);
xor U10963 (N_10963,N_10124,N_10328);
nand U10964 (N_10964,N_10237,N_10471);
or U10965 (N_10965,N_10453,N_10187);
nand U10966 (N_10966,N_10485,N_10136);
and U10967 (N_10967,N_10126,N_10370);
xor U10968 (N_10968,N_10478,N_10299);
nor U10969 (N_10969,N_10187,N_10116);
or U10970 (N_10970,N_10282,N_10084);
or U10971 (N_10971,N_10477,N_10348);
xnor U10972 (N_10972,N_10004,N_10297);
or U10973 (N_10973,N_10393,N_10265);
or U10974 (N_10974,N_10471,N_10372);
nand U10975 (N_10975,N_10381,N_10092);
nand U10976 (N_10976,N_10339,N_10013);
nand U10977 (N_10977,N_10445,N_10363);
xor U10978 (N_10978,N_10215,N_10311);
and U10979 (N_10979,N_10129,N_10078);
and U10980 (N_10980,N_10491,N_10307);
nand U10981 (N_10981,N_10406,N_10417);
or U10982 (N_10982,N_10209,N_10308);
or U10983 (N_10983,N_10054,N_10468);
nor U10984 (N_10984,N_10459,N_10214);
xor U10985 (N_10985,N_10128,N_10122);
xnor U10986 (N_10986,N_10437,N_10325);
nand U10987 (N_10987,N_10438,N_10132);
and U10988 (N_10988,N_10057,N_10206);
xnor U10989 (N_10989,N_10229,N_10447);
and U10990 (N_10990,N_10010,N_10149);
or U10991 (N_10991,N_10379,N_10079);
and U10992 (N_10992,N_10391,N_10053);
and U10993 (N_10993,N_10480,N_10038);
nor U10994 (N_10994,N_10008,N_10119);
or U10995 (N_10995,N_10013,N_10126);
xnor U10996 (N_10996,N_10446,N_10076);
xnor U10997 (N_10997,N_10318,N_10338);
or U10998 (N_10998,N_10055,N_10459);
xor U10999 (N_10999,N_10167,N_10108);
or U11000 (N_11000,N_10804,N_10905);
or U11001 (N_11001,N_10711,N_10811);
nand U11002 (N_11002,N_10938,N_10575);
or U11003 (N_11003,N_10697,N_10590);
nor U11004 (N_11004,N_10599,N_10844);
xor U11005 (N_11005,N_10556,N_10629);
xnor U11006 (N_11006,N_10975,N_10836);
xor U11007 (N_11007,N_10601,N_10799);
or U11008 (N_11008,N_10684,N_10837);
or U11009 (N_11009,N_10874,N_10501);
or U11010 (N_11010,N_10890,N_10536);
xnor U11011 (N_11011,N_10880,N_10869);
xor U11012 (N_11012,N_10524,N_10542);
or U11013 (N_11013,N_10682,N_10506);
or U11014 (N_11014,N_10879,N_10801);
nor U11015 (N_11015,N_10663,N_10841);
and U11016 (N_11016,N_10757,N_10912);
xnor U11017 (N_11017,N_10987,N_10835);
and U11018 (N_11018,N_10892,N_10510);
or U11019 (N_11019,N_10883,N_10725);
nand U11020 (N_11020,N_10852,N_10698);
nand U11021 (N_11021,N_10878,N_10621);
nor U11022 (N_11022,N_10974,N_10894);
xor U11023 (N_11023,N_10911,N_10768);
or U11024 (N_11024,N_10956,N_10834);
nor U11025 (N_11025,N_10661,N_10942);
nand U11026 (N_11026,N_10659,N_10752);
xor U11027 (N_11027,N_10808,N_10960);
xnor U11028 (N_11028,N_10641,N_10703);
nand U11029 (N_11029,N_10673,N_10988);
nand U11030 (N_11030,N_10769,N_10753);
or U11031 (N_11031,N_10791,N_10613);
nand U11032 (N_11032,N_10903,N_10782);
nand U11033 (N_11033,N_10785,N_10686);
nor U11034 (N_11034,N_10679,N_10587);
nand U11035 (N_11035,N_10802,N_10593);
or U11036 (N_11036,N_10934,N_10657);
nor U11037 (N_11037,N_10548,N_10794);
or U11038 (N_11038,N_10625,N_10868);
and U11039 (N_11039,N_10756,N_10718);
or U11040 (N_11040,N_10717,N_10652);
and U11041 (N_11041,N_10516,N_10821);
and U11042 (N_11042,N_10700,N_10944);
xnor U11043 (N_11043,N_10685,N_10680);
nand U11044 (N_11044,N_10677,N_10538);
nor U11045 (N_11045,N_10866,N_10990);
nand U11046 (N_11046,N_10598,N_10906);
and U11047 (N_11047,N_10527,N_10747);
nand U11048 (N_11048,N_10740,N_10992);
and U11049 (N_11049,N_10568,N_10676);
and U11050 (N_11050,N_10929,N_10735);
and U11051 (N_11051,N_10732,N_10644);
nand U11052 (N_11052,N_10724,N_10889);
nor U11053 (N_11053,N_10594,N_10646);
nand U11054 (N_11054,N_10543,N_10754);
nand U11055 (N_11055,N_10643,N_10925);
nand U11056 (N_11056,N_10557,N_10876);
nand U11057 (N_11057,N_10867,N_10623);
nor U11058 (N_11058,N_10777,N_10537);
nand U11059 (N_11059,N_10519,N_10504);
and U11060 (N_11060,N_10591,N_10639);
nand U11061 (N_11061,N_10694,N_10742);
nand U11062 (N_11062,N_10619,N_10508);
nand U11063 (N_11063,N_10775,N_10710);
nor U11064 (N_11064,N_10743,N_10529);
xnor U11065 (N_11065,N_10983,N_10668);
or U11066 (N_11066,N_10976,N_10952);
or U11067 (N_11067,N_10848,N_10946);
nand U11068 (N_11068,N_10585,N_10935);
and U11069 (N_11069,N_10721,N_10931);
nand U11070 (N_11070,N_10574,N_10603);
or U11071 (N_11071,N_10991,N_10970);
and U11072 (N_11072,N_10772,N_10515);
or U11073 (N_11073,N_10546,N_10569);
or U11074 (N_11074,N_10793,N_10616);
xnor U11075 (N_11075,N_10653,N_10761);
xor U11076 (N_11076,N_10887,N_10885);
and U11077 (N_11077,N_10654,N_10505);
or U11078 (N_11078,N_10691,N_10640);
or U11079 (N_11079,N_10534,N_10770);
xnor U11080 (N_11080,N_10642,N_10749);
xnor U11081 (N_11081,N_10798,N_10994);
nor U11082 (N_11082,N_10588,N_10859);
and U11083 (N_11083,N_10738,N_10986);
and U11084 (N_11084,N_10972,N_10949);
and U11085 (N_11085,N_10571,N_10672);
nand U11086 (N_11086,N_10541,N_10719);
nand U11087 (N_11087,N_10726,N_10513);
nand U11088 (N_11088,N_10873,N_10830);
or U11089 (N_11089,N_10933,N_10555);
nor U11090 (N_11090,N_10628,N_10815);
xnor U11091 (N_11091,N_10984,N_10609);
and U11092 (N_11092,N_10670,N_10843);
nand U11093 (N_11093,N_10778,N_10796);
or U11094 (N_11094,N_10688,N_10664);
nand U11095 (N_11095,N_10893,N_10671);
and U11096 (N_11096,N_10577,N_10759);
and U11097 (N_11097,N_10832,N_10792);
nor U11098 (N_11098,N_10596,N_10918);
or U11099 (N_11099,N_10667,N_10825);
and U11100 (N_11100,N_10560,N_10714);
nand U11101 (N_11101,N_10838,N_10611);
and U11102 (N_11102,N_10958,N_10583);
or U11103 (N_11103,N_10584,N_10532);
nor U11104 (N_11104,N_10520,N_10985);
and U11105 (N_11105,N_10552,N_10689);
and U11106 (N_11106,N_10922,N_10900);
nand U11107 (N_11107,N_10779,N_10813);
nor U11108 (N_11108,N_10981,N_10712);
xnor U11109 (N_11109,N_10612,N_10713);
or U11110 (N_11110,N_10540,N_10803);
nor U11111 (N_11111,N_10518,N_10982);
nor U11112 (N_11112,N_10699,N_10839);
nor U11113 (N_11113,N_10704,N_10898);
nand U11114 (N_11114,N_10955,N_10943);
and U11115 (N_11115,N_10678,N_10891);
xnor U11116 (N_11116,N_10845,N_10549);
nor U11117 (N_11117,N_10610,N_10503);
nor U11118 (N_11118,N_10702,N_10851);
xnor U11119 (N_11119,N_10608,N_10683);
nor U11120 (N_11120,N_10731,N_10969);
xnor U11121 (N_11121,N_10705,N_10865);
or U11122 (N_11122,N_10822,N_10805);
or U11123 (N_11123,N_10924,N_10957);
nand U11124 (N_11124,N_10927,N_10744);
xor U11125 (N_11125,N_10675,N_10662);
nand U11126 (N_11126,N_10788,N_10860);
or U11127 (N_11127,N_10758,N_10950);
nand U11128 (N_11128,N_10962,N_10923);
or U11129 (N_11129,N_10530,N_10550);
nand U11130 (N_11130,N_10771,N_10833);
or U11131 (N_11131,N_10736,N_10895);
nand U11132 (N_11132,N_10635,N_10637);
nor U11133 (N_11133,N_10763,N_10511);
or U11134 (N_11134,N_10904,N_10787);
or U11135 (N_11135,N_10539,N_10553);
and U11136 (N_11136,N_10881,N_10776);
nand U11137 (N_11137,N_10709,N_10854);
xor U11138 (N_11138,N_10762,N_10930);
nor U11139 (N_11139,N_10998,N_10597);
xnor U11140 (N_11140,N_10996,N_10914);
xnor U11141 (N_11141,N_10669,N_10936);
or U11142 (N_11142,N_10857,N_10795);
or U11143 (N_11143,N_10812,N_10526);
xor U11144 (N_11144,N_10966,N_10733);
xor U11145 (N_11145,N_10600,N_10720);
nor U11146 (N_11146,N_10727,N_10514);
xor U11147 (N_11147,N_10863,N_10502);
or U11148 (N_11148,N_10809,N_10897);
or U11149 (N_11149,N_10564,N_10765);
xor U11150 (N_11150,N_10707,N_10977);
or U11151 (N_11151,N_10917,N_10989);
and U11152 (N_11152,N_10947,N_10919);
xnor U11153 (N_11153,N_10728,N_10622);
nor U11154 (N_11154,N_10693,N_10937);
nand U11155 (N_11155,N_10655,N_10806);
nor U11156 (N_11156,N_10995,N_10921);
or U11157 (N_11157,N_10522,N_10861);
and U11158 (N_11158,N_10630,N_10939);
nor U11159 (N_11159,N_10884,N_10696);
xnor U11160 (N_11160,N_10722,N_10886);
nor U11161 (N_11161,N_10558,N_10807);
and U11162 (N_11162,N_10824,N_10650);
xnor U11163 (N_11163,N_10716,N_10820);
nor U11164 (N_11164,N_10627,N_10606);
nor U11165 (N_11165,N_10547,N_10945);
xor U11166 (N_11166,N_10647,N_10563);
or U11167 (N_11167,N_10739,N_10614);
and U11168 (N_11168,N_10823,N_10831);
nor U11169 (N_11169,N_10959,N_10875);
xor U11170 (N_11170,N_10973,N_10554);
xnor U11171 (N_11171,N_10666,N_10658);
nor U11172 (N_11172,N_10559,N_10500);
and U11173 (N_11173,N_10797,N_10764);
or U11174 (N_11174,N_10523,N_10853);
and U11175 (N_11175,N_10638,N_10544);
nand U11176 (N_11176,N_10877,N_10636);
xnor U11177 (N_11177,N_10858,N_10649);
nor U11178 (N_11178,N_10872,N_10971);
nand U11179 (N_11179,N_10800,N_10734);
or U11180 (N_11180,N_10856,N_10509);
or U11181 (N_11181,N_10964,N_10978);
xor U11182 (N_11182,N_10748,N_10774);
nor U11183 (N_11183,N_10902,N_10790);
or U11184 (N_11184,N_10737,N_10531);
or U11185 (N_11185,N_10783,N_10656);
or U11186 (N_11186,N_10741,N_10589);
nor U11187 (N_11187,N_10660,N_10701);
and U11188 (N_11188,N_10545,N_10827);
nand U11189 (N_11189,N_10690,N_10850);
nand U11190 (N_11190,N_10915,N_10789);
or U11191 (N_11191,N_10784,N_10648);
nand U11192 (N_11192,N_10521,N_10665);
nand U11193 (N_11193,N_10525,N_10751);
nor U11194 (N_11194,N_10692,N_10602);
nor U11195 (N_11195,N_10979,N_10512);
nor U11196 (N_11196,N_10948,N_10913);
xor U11197 (N_11197,N_10968,N_10864);
and U11198 (N_11198,N_10870,N_10965);
xor U11199 (N_11199,N_10829,N_10633);
or U11200 (N_11200,N_10626,N_10745);
or U11201 (N_11201,N_10535,N_10573);
nand U11202 (N_11202,N_10579,N_10615);
xnor U11203 (N_11203,N_10817,N_10561);
nor U11204 (N_11204,N_10816,N_10826);
nor U11205 (N_11205,N_10941,N_10729);
and U11206 (N_11206,N_10961,N_10708);
nand U11207 (N_11207,N_10617,N_10760);
nand U11208 (N_11208,N_10651,N_10624);
nand U11209 (N_11209,N_10818,N_10755);
and U11210 (N_11210,N_10862,N_10730);
xnor U11211 (N_11211,N_10828,N_10967);
and U11212 (N_11212,N_10871,N_10576);
xor U11213 (N_11213,N_10681,N_10715);
nor U11214 (N_11214,N_10780,N_10706);
and U11215 (N_11215,N_10562,N_10814);
or U11216 (N_11216,N_10842,N_10882);
xnor U11217 (N_11217,N_10566,N_10582);
or U11218 (N_11218,N_10773,N_10580);
nand U11219 (N_11219,N_10618,N_10632);
nand U11220 (N_11220,N_10951,N_10819);
and U11221 (N_11221,N_10781,N_10551);
nor U11222 (N_11222,N_10908,N_10810);
nor U11223 (N_11223,N_10631,N_10855);
or U11224 (N_11224,N_10901,N_10953);
nand U11225 (N_11225,N_10786,N_10963);
and U11226 (N_11226,N_10645,N_10767);
and U11227 (N_11227,N_10907,N_10533);
xnor U11228 (N_11228,N_10940,N_10849);
nor U11229 (N_11229,N_10840,N_10565);
and U11230 (N_11230,N_10567,N_10604);
nor U11231 (N_11231,N_10634,N_10746);
nand U11232 (N_11232,N_10750,N_10980);
xor U11233 (N_11233,N_10954,N_10620);
and U11234 (N_11234,N_10920,N_10607);
or U11235 (N_11235,N_10687,N_10993);
nor U11236 (N_11236,N_10605,N_10570);
or U11237 (N_11237,N_10928,N_10932);
nor U11238 (N_11238,N_10723,N_10766);
xor U11239 (N_11239,N_10586,N_10846);
nor U11240 (N_11240,N_10926,N_10595);
or U11241 (N_11241,N_10916,N_10572);
xnor U11242 (N_11242,N_10997,N_10999);
xor U11243 (N_11243,N_10528,N_10910);
nor U11244 (N_11244,N_10847,N_10899);
xor U11245 (N_11245,N_10507,N_10896);
nor U11246 (N_11246,N_10909,N_10578);
or U11247 (N_11247,N_10695,N_10674);
xnor U11248 (N_11248,N_10888,N_10581);
and U11249 (N_11249,N_10517,N_10592);
or U11250 (N_11250,N_10794,N_10829);
xor U11251 (N_11251,N_10577,N_10524);
and U11252 (N_11252,N_10778,N_10568);
and U11253 (N_11253,N_10625,N_10732);
xnor U11254 (N_11254,N_10719,N_10957);
nand U11255 (N_11255,N_10786,N_10788);
nor U11256 (N_11256,N_10515,N_10560);
and U11257 (N_11257,N_10858,N_10843);
or U11258 (N_11258,N_10891,N_10877);
nor U11259 (N_11259,N_10501,N_10616);
or U11260 (N_11260,N_10682,N_10898);
xor U11261 (N_11261,N_10618,N_10805);
and U11262 (N_11262,N_10916,N_10607);
xnor U11263 (N_11263,N_10507,N_10641);
and U11264 (N_11264,N_10990,N_10812);
nand U11265 (N_11265,N_10780,N_10748);
or U11266 (N_11266,N_10759,N_10596);
nand U11267 (N_11267,N_10737,N_10664);
xnor U11268 (N_11268,N_10696,N_10843);
and U11269 (N_11269,N_10898,N_10883);
and U11270 (N_11270,N_10664,N_10624);
xor U11271 (N_11271,N_10828,N_10806);
nor U11272 (N_11272,N_10984,N_10778);
and U11273 (N_11273,N_10831,N_10687);
and U11274 (N_11274,N_10709,N_10944);
xnor U11275 (N_11275,N_10721,N_10990);
xor U11276 (N_11276,N_10709,N_10548);
nand U11277 (N_11277,N_10817,N_10614);
nand U11278 (N_11278,N_10905,N_10968);
or U11279 (N_11279,N_10985,N_10888);
xnor U11280 (N_11280,N_10568,N_10593);
xnor U11281 (N_11281,N_10675,N_10572);
nand U11282 (N_11282,N_10603,N_10662);
and U11283 (N_11283,N_10864,N_10724);
xnor U11284 (N_11284,N_10920,N_10995);
nor U11285 (N_11285,N_10604,N_10580);
nand U11286 (N_11286,N_10576,N_10924);
and U11287 (N_11287,N_10904,N_10682);
or U11288 (N_11288,N_10644,N_10838);
or U11289 (N_11289,N_10583,N_10647);
nand U11290 (N_11290,N_10556,N_10637);
or U11291 (N_11291,N_10971,N_10952);
xor U11292 (N_11292,N_10582,N_10752);
xor U11293 (N_11293,N_10746,N_10968);
or U11294 (N_11294,N_10801,N_10809);
nor U11295 (N_11295,N_10645,N_10835);
and U11296 (N_11296,N_10598,N_10612);
xor U11297 (N_11297,N_10843,N_10531);
and U11298 (N_11298,N_10962,N_10972);
nand U11299 (N_11299,N_10826,N_10766);
nor U11300 (N_11300,N_10601,N_10740);
nor U11301 (N_11301,N_10886,N_10649);
xor U11302 (N_11302,N_10928,N_10567);
xnor U11303 (N_11303,N_10788,N_10805);
or U11304 (N_11304,N_10615,N_10971);
nor U11305 (N_11305,N_10898,N_10644);
nand U11306 (N_11306,N_10845,N_10923);
or U11307 (N_11307,N_10695,N_10551);
xor U11308 (N_11308,N_10646,N_10787);
nand U11309 (N_11309,N_10659,N_10885);
or U11310 (N_11310,N_10887,N_10604);
xnor U11311 (N_11311,N_10957,N_10705);
and U11312 (N_11312,N_10977,N_10603);
or U11313 (N_11313,N_10727,N_10833);
and U11314 (N_11314,N_10771,N_10683);
or U11315 (N_11315,N_10526,N_10845);
nor U11316 (N_11316,N_10974,N_10917);
nor U11317 (N_11317,N_10876,N_10712);
nor U11318 (N_11318,N_10699,N_10509);
and U11319 (N_11319,N_10937,N_10667);
nand U11320 (N_11320,N_10618,N_10981);
or U11321 (N_11321,N_10877,N_10512);
nand U11322 (N_11322,N_10631,N_10721);
or U11323 (N_11323,N_10978,N_10946);
nor U11324 (N_11324,N_10518,N_10562);
nor U11325 (N_11325,N_10513,N_10799);
nor U11326 (N_11326,N_10895,N_10784);
nor U11327 (N_11327,N_10880,N_10916);
and U11328 (N_11328,N_10697,N_10952);
nor U11329 (N_11329,N_10732,N_10500);
nand U11330 (N_11330,N_10849,N_10854);
and U11331 (N_11331,N_10853,N_10554);
nor U11332 (N_11332,N_10605,N_10852);
or U11333 (N_11333,N_10666,N_10737);
and U11334 (N_11334,N_10538,N_10925);
nand U11335 (N_11335,N_10625,N_10892);
nand U11336 (N_11336,N_10993,N_10924);
nand U11337 (N_11337,N_10994,N_10593);
xnor U11338 (N_11338,N_10868,N_10841);
nor U11339 (N_11339,N_10669,N_10759);
and U11340 (N_11340,N_10904,N_10581);
and U11341 (N_11341,N_10686,N_10939);
xor U11342 (N_11342,N_10656,N_10557);
and U11343 (N_11343,N_10703,N_10738);
nand U11344 (N_11344,N_10852,N_10516);
xnor U11345 (N_11345,N_10675,N_10691);
xor U11346 (N_11346,N_10997,N_10726);
nor U11347 (N_11347,N_10569,N_10864);
or U11348 (N_11348,N_10945,N_10822);
nand U11349 (N_11349,N_10814,N_10685);
and U11350 (N_11350,N_10943,N_10880);
or U11351 (N_11351,N_10740,N_10960);
xnor U11352 (N_11352,N_10808,N_10669);
and U11353 (N_11353,N_10734,N_10825);
nand U11354 (N_11354,N_10903,N_10864);
or U11355 (N_11355,N_10897,N_10563);
nand U11356 (N_11356,N_10625,N_10619);
and U11357 (N_11357,N_10949,N_10862);
nand U11358 (N_11358,N_10904,N_10917);
nand U11359 (N_11359,N_10643,N_10939);
nor U11360 (N_11360,N_10898,N_10658);
nand U11361 (N_11361,N_10936,N_10909);
nand U11362 (N_11362,N_10872,N_10697);
nor U11363 (N_11363,N_10664,N_10775);
xor U11364 (N_11364,N_10781,N_10893);
or U11365 (N_11365,N_10983,N_10998);
xor U11366 (N_11366,N_10545,N_10717);
nor U11367 (N_11367,N_10562,N_10530);
xor U11368 (N_11368,N_10540,N_10568);
nor U11369 (N_11369,N_10619,N_10861);
xor U11370 (N_11370,N_10957,N_10891);
xnor U11371 (N_11371,N_10561,N_10933);
nor U11372 (N_11372,N_10614,N_10647);
xnor U11373 (N_11373,N_10736,N_10585);
and U11374 (N_11374,N_10864,N_10714);
xor U11375 (N_11375,N_10828,N_10717);
or U11376 (N_11376,N_10595,N_10691);
xnor U11377 (N_11377,N_10557,N_10776);
nor U11378 (N_11378,N_10533,N_10874);
or U11379 (N_11379,N_10667,N_10990);
and U11380 (N_11380,N_10855,N_10988);
nand U11381 (N_11381,N_10683,N_10975);
and U11382 (N_11382,N_10862,N_10905);
and U11383 (N_11383,N_10847,N_10836);
xor U11384 (N_11384,N_10816,N_10519);
xnor U11385 (N_11385,N_10681,N_10693);
xor U11386 (N_11386,N_10691,N_10859);
and U11387 (N_11387,N_10561,N_10765);
nand U11388 (N_11388,N_10983,N_10521);
nor U11389 (N_11389,N_10936,N_10528);
xor U11390 (N_11390,N_10992,N_10938);
nand U11391 (N_11391,N_10851,N_10751);
and U11392 (N_11392,N_10729,N_10902);
nor U11393 (N_11393,N_10848,N_10637);
nor U11394 (N_11394,N_10500,N_10541);
nand U11395 (N_11395,N_10828,N_10733);
and U11396 (N_11396,N_10536,N_10619);
nand U11397 (N_11397,N_10878,N_10535);
xor U11398 (N_11398,N_10853,N_10684);
and U11399 (N_11399,N_10505,N_10511);
nor U11400 (N_11400,N_10745,N_10527);
nand U11401 (N_11401,N_10872,N_10838);
and U11402 (N_11402,N_10996,N_10708);
nand U11403 (N_11403,N_10528,N_10660);
nor U11404 (N_11404,N_10815,N_10546);
nor U11405 (N_11405,N_10699,N_10849);
xor U11406 (N_11406,N_10669,N_10731);
nand U11407 (N_11407,N_10994,N_10544);
xor U11408 (N_11408,N_10862,N_10508);
or U11409 (N_11409,N_10626,N_10871);
or U11410 (N_11410,N_10704,N_10938);
xor U11411 (N_11411,N_10858,N_10621);
and U11412 (N_11412,N_10941,N_10551);
nand U11413 (N_11413,N_10619,N_10569);
nor U11414 (N_11414,N_10773,N_10665);
or U11415 (N_11415,N_10809,N_10818);
or U11416 (N_11416,N_10822,N_10987);
nand U11417 (N_11417,N_10679,N_10906);
xor U11418 (N_11418,N_10705,N_10570);
nand U11419 (N_11419,N_10596,N_10702);
xor U11420 (N_11420,N_10902,N_10823);
xor U11421 (N_11421,N_10558,N_10533);
or U11422 (N_11422,N_10946,N_10895);
and U11423 (N_11423,N_10780,N_10637);
and U11424 (N_11424,N_10621,N_10733);
xor U11425 (N_11425,N_10633,N_10867);
or U11426 (N_11426,N_10943,N_10665);
and U11427 (N_11427,N_10699,N_10714);
nand U11428 (N_11428,N_10834,N_10914);
and U11429 (N_11429,N_10807,N_10748);
or U11430 (N_11430,N_10866,N_10552);
or U11431 (N_11431,N_10913,N_10708);
nand U11432 (N_11432,N_10884,N_10974);
nor U11433 (N_11433,N_10669,N_10525);
nand U11434 (N_11434,N_10952,N_10782);
nand U11435 (N_11435,N_10916,N_10967);
xor U11436 (N_11436,N_10812,N_10519);
nand U11437 (N_11437,N_10653,N_10855);
and U11438 (N_11438,N_10569,N_10999);
or U11439 (N_11439,N_10591,N_10660);
xor U11440 (N_11440,N_10977,N_10921);
xnor U11441 (N_11441,N_10838,N_10502);
and U11442 (N_11442,N_10820,N_10563);
or U11443 (N_11443,N_10674,N_10686);
and U11444 (N_11444,N_10545,N_10562);
or U11445 (N_11445,N_10974,N_10636);
or U11446 (N_11446,N_10603,N_10763);
or U11447 (N_11447,N_10819,N_10975);
xor U11448 (N_11448,N_10608,N_10613);
or U11449 (N_11449,N_10935,N_10700);
and U11450 (N_11450,N_10600,N_10838);
or U11451 (N_11451,N_10835,N_10710);
xor U11452 (N_11452,N_10516,N_10553);
xor U11453 (N_11453,N_10974,N_10714);
and U11454 (N_11454,N_10854,N_10572);
nand U11455 (N_11455,N_10984,N_10843);
nor U11456 (N_11456,N_10889,N_10720);
or U11457 (N_11457,N_10600,N_10915);
nor U11458 (N_11458,N_10949,N_10849);
or U11459 (N_11459,N_10924,N_10682);
and U11460 (N_11460,N_10896,N_10959);
xnor U11461 (N_11461,N_10857,N_10601);
nand U11462 (N_11462,N_10806,N_10562);
nand U11463 (N_11463,N_10970,N_10692);
or U11464 (N_11464,N_10808,N_10950);
or U11465 (N_11465,N_10754,N_10827);
nor U11466 (N_11466,N_10753,N_10926);
nand U11467 (N_11467,N_10573,N_10826);
or U11468 (N_11468,N_10914,N_10565);
nand U11469 (N_11469,N_10943,N_10957);
nand U11470 (N_11470,N_10651,N_10722);
xor U11471 (N_11471,N_10520,N_10941);
and U11472 (N_11472,N_10745,N_10633);
nand U11473 (N_11473,N_10806,N_10650);
or U11474 (N_11474,N_10636,N_10887);
or U11475 (N_11475,N_10588,N_10589);
or U11476 (N_11476,N_10657,N_10552);
nand U11477 (N_11477,N_10536,N_10506);
or U11478 (N_11478,N_10856,N_10576);
xor U11479 (N_11479,N_10968,N_10874);
xor U11480 (N_11480,N_10896,N_10549);
and U11481 (N_11481,N_10636,N_10862);
or U11482 (N_11482,N_10827,N_10981);
or U11483 (N_11483,N_10558,N_10909);
nand U11484 (N_11484,N_10680,N_10838);
and U11485 (N_11485,N_10698,N_10931);
and U11486 (N_11486,N_10983,N_10928);
and U11487 (N_11487,N_10809,N_10549);
nor U11488 (N_11488,N_10613,N_10551);
and U11489 (N_11489,N_10707,N_10549);
or U11490 (N_11490,N_10959,N_10818);
and U11491 (N_11491,N_10752,N_10506);
and U11492 (N_11492,N_10716,N_10773);
xnor U11493 (N_11493,N_10576,N_10870);
and U11494 (N_11494,N_10667,N_10987);
nand U11495 (N_11495,N_10717,N_10669);
nor U11496 (N_11496,N_10641,N_10743);
nor U11497 (N_11497,N_10906,N_10557);
or U11498 (N_11498,N_10791,N_10897);
or U11499 (N_11499,N_10617,N_10974);
nand U11500 (N_11500,N_11241,N_11077);
xnor U11501 (N_11501,N_11229,N_11366);
or U11502 (N_11502,N_11365,N_11245);
nand U11503 (N_11503,N_11086,N_11412);
and U11504 (N_11504,N_11251,N_11113);
nand U11505 (N_11505,N_11421,N_11068);
and U11506 (N_11506,N_11410,N_11160);
nor U11507 (N_11507,N_11411,N_11362);
or U11508 (N_11508,N_11234,N_11022);
xor U11509 (N_11509,N_11282,N_11424);
xnor U11510 (N_11510,N_11111,N_11479);
nand U11511 (N_11511,N_11401,N_11448);
nand U11512 (N_11512,N_11019,N_11271);
xor U11513 (N_11513,N_11453,N_11011);
nor U11514 (N_11514,N_11480,N_11288);
nor U11515 (N_11515,N_11198,N_11031);
and U11516 (N_11516,N_11335,N_11294);
xor U11517 (N_11517,N_11139,N_11498);
nor U11518 (N_11518,N_11418,N_11233);
nor U11519 (N_11519,N_11308,N_11432);
or U11520 (N_11520,N_11322,N_11004);
nor U11521 (N_11521,N_11191,N_11240);
nand U11522 (N_11522,N_11426,N_11003);
nand U11523 (N_11523,N_11008,N_11005);
nand U11524 (N_11524,N_11243,N_11330);
or U11525 (N_11525,N_11007,N_11168);
xor U11526 (N_11526,N_11326,N_11306);
nand U11527 (N_11527,N_11056,N_11201);
or U11528 (N_11528,N_11457,N_11475);
nand U11529 (N_11529,N_11493,N_11205);
nand U11530 (N_11530,N_11211,N_11488);
or U11531 (N_11531,N_11334,N_11486);
nor U11532 (N_11532,N_11473,N_11038);
nand U11533 (N_11533,N_11236,N_11069);
nor U11534 (N_11534,N_11222,N_11394);
xnor U11535 (N_11535,N_11329,N_11262);
nor U11536 (N_11536,N_11070,N_11268);
or U11537 (N_11537,N_11417,N_11055);
and U11538 (N_11538,N_11231,N_11438);
nor U11539 (N_11539,N_11097,N_11199);
xnor U11540 (N_11540,N_11416,N_11336);
nand U11541 (N_11541,N_11396,N_11147);
xor U11542 (N_11542,N_11140,N_11254);
nor U11543 (N_11543,N_11067,N_11152);
or U11544 (N_11544,N_11323,N_11000);
or U11545 (N_11545,N_11403,N_11181);
xnor U11546 (N_11546,N_11024,N_11006);
and U11547 (N_11547,N_11103,N_11481);
nor U11548 (N_11548,N_11376,N_11230);
nand U11549 (N_11549,N_11435,N_11300);
xor U11550 (N_11550,N_11149,N_11409);
and U11551 (N_11551,N_11018,N_11387);
xnor U11552 (N_11552,N_11227,N_11203);
nand U11553 (N_11553,N_11183,N_11184);
nand U11554 (N_11554,N_11249,N_11182);
or U11555 (N_11555,N_11001,N_11291);
and U11556 (N_11556,N_11063,N_11154);
and U11557 (N_11557,N_11050,N_11261);
and U11558 (N_11558,N_11355,N_11253);
xor U11559 (N_11559,N_11162,N_11075);
xor U11560 (N_11560,N_11037,N_11039);
and U11561 (N_11561,N_11247,N_11419);
xnor U11562 (N_11562,N_11360,N_11277);
xnor U11563 (N_11563,N_11440,N_11290);
nor U11564 (N_11564,N_11248,N_11172);
and U11565 (N_11565,N_11451,N_11225);
or U11566 (N_11566,N_11458,N_11136);
nand U11567 (N_11567,N_11084,N_11476);
and U11568 (N_11568,N_11081,N_11073);
nor U11569 (N_11569,N_11372,N_11027);
nor U11570 (N_11570,N_11302,N_11014);
and U11571 (N_11571,N_11361,N_11464);
or U11572 (N_11572,N_11337,N_11135);
and U11573 (N_11573,N_11094,N_11218);
nand U11574 (N_11574,N_11100,N_11487);
or U11575 (N_11575,N_11058,N_11207);
or U11576 (N_11576,N_11364,N_11491);
and U11577 (N_11577,N_11275,N_11313);
xor U11578 (N_11578,N_11144,N_11485);
nor U11579 (N_11579,N_11499,N_11118);
nor U11580 (N_11580,N_11307,N_11404);
xnor U11581 (N_11581,N_11369,N_11321);
nor U11582 (N_11582,N_11434,N_11345);
and U11583 (N_11583,N_11331,N_11352);
xor U11584 (N_11584,N_11133,N_11375);
or U11585 (N_11585,N_11319,N_11289);
nor U11586 (N_11586,N_11353,N_11456);
or U11587 (N_11587,N_11310,N_11129);
xor U11588 (N_11588,N_11472,N_11455);
or U11589 (N_11589,N_11064,N_11042);
and U11590 (N_11590,N_11017,N_11060);
nor U11591 (N_11591,N_11425,N_11420);
xnor U11592 (N_11592,N_11287,N_11213);
or U11593 (N_11593,N_11119,N_11284);
nand U11594 (N_11594,N_11212,N_11358);
and U11595 (N_11595,N_11188,N_11130);
or U11596 (N_11596,N_11304,N_11303);
nand U11597 (N_11597,N_11382,N_11301);
nand U11598 (N_11598,N_11398,N_11093);
and U11599 (N_11599,N_11413,N_11071);
nand U11600 (N_11600,N_11428,N_11347);
xnor U11601 (N_11601,N_11433,N_11167);
xor U11602 (N_11602,N_11020,N_11354);
nor U11603 (N_11603,N_11047,N_11496);
nand U11604 (N_11604,N_11048,N_11083);
nand U11605 (N_11605,N_11328,N_11185);
or U11606 (N_11606,N_11250,N_11497);
and U11607 (N_11607,N_11286,N_11105);
or U11608 (N_11608,N_11223,N_11034);
and U11609 (N_11609,N_11078,N_11214);
xnor U11610 (N_11610,N_11276,N_11080);
or U11611 (N_11611,N_11040,N_11053);
xnor U11612 (N_11612,N_11390,N_11357);
or U11613 (N_11613,N_11195,N_11171);
and U11614 (N_11614,N_11257,N_11327);
and U11615 (N_11615,N_11052,N_11033);
xor U11616 (N_11616,N_11489,N_11112);
xnor U11617 (N_11617,N_11346,N_11132);
nor U11618 (N_11618,N_11108,N_11494);
nand U11619 (N_11619,N_11383,N_11091);
or U11620 (N_11620,N_11082,N_11166);
and U11621 (N_11621,N_11274,N_11454);
nor U11622 (N_11622,N_11415,N_11441);
and U11623 (N_11623,N_11202,N_11102);
xnor U11624 (N_11624,N_11309,N_11232);
xor U11625 (N_11625,N_11459,N_11386);
nor U11626 (N_11626,N_11397,N_11175);
nor U11627 (N_11627,N_11127,N_11079);
and U11628 (N_11628,N_11338,N_11384);
nand U11629 (N_11629,N_11228,N_11340);
nand U11630 (N_11630,N_11490,N_11076);
or U11631 (N_11631,N_11393,N_11348);
and U11632 (N_11632,N_11148,N_11349);
nand U11633 (N_11633,N_11279,N_11278);
and U11634 (N_11634,N_11002,N_11138);
xor U11635 (N_11635,N_11155,N_11466);
nor U11636 (N_11636,N_11315,N_11442);
or U11637 (N_11637,N_11283,N_11312);
nand U11638 (N_11638,N_11344,N_11235);
xnor U11639 (N_11639,N_11204,N_11012);
nand U11640 (N_11640,N_11074,N_11174);
and U11641 (N_11641,N_11450,N_11297);
and U11642 (N_11642,N_11314,N_11395);
nor U11643 (N_11643,N_11117,N_11392);
or U11644 (N_11644,N_11427,N_11122);
or U11645 (N_11645,N_11495,N_11317);
and U11646 (N_11646,N_11374,N_11324);
or U11647 (N_11647,N_11165,N_11281);
and U11648 (N_11648,N_11263,N_11096);
or U11649 (N_11649,N_11028,N_11359);
xor U11650 (N_11650,N_11484,N_11462);
or U11651 (N_11651,N_11131,N_11126);
nor U11652 (N_11652,N_11046,N_11157);
nor U11653 (N_11653,N_11025,N_11380);
or U11654 (N_11654,N_11368,N_11371);
nor U11655 (N_11655,N_11273,N_11333);
nand U11656 (N_11656,N_11461,N_11035);
nor U11657 (N_11657,N_11242,N_11176);
or U11658 (N_11658,N_11219,N_11153);
nand U11659 (N_11659,N_11180,N_11021);
or U11660 (N_11660,N_11095,N_11173);
nand U11661 (N_11661,N_11187,N_11054);
nor U11662 (N_11662,N_11363,N_11237);
and U11663 (N_11663,N_11085,N_11471);
and U11664 (N_11664,N_11252,N_11146);
or U11665 (N_11665,N_11087,N_11446);
or U11666 (N_11666,N_11305,N_11292);
nor U11667 (N_11667,N_11143,N_11266);
xor U11668 (N_11668,N_11381,N_11036);
and U11669 (N_11669,N_11178,N_11158);
xnor U11670 (N_11670,N_11217,N_11116);
xor U11671 (N_11671,N_11057,N_11460);
nand U11672 (N_11672,N_11032,N_11164);
and U11673 (N_11673,N_11110,N_11325);
xor U11674 (N_11674,N_11269,N_11389);
and U11675 (N_11675,N_11430,N_11370);
or U11676 (N_11676,N_11339,N_11142);
or U11677 (N_11677,N_11316,N_11373);
nand U11678 (N_11678,N_11391,N_11469);
xor U11679 (N_11679,N_11089,N_11467);
and U11680 (N_11680,N_11114,N_11026);
nand U11681 (N_11681,N_11436,N_11123);
xnor U11682 (N_11682,N_11072,N_11090);
nand U11683 (N_11683,N_11452,N_11221);
nor U11684 (N_11684,N_11402,N_11244);
nand U11685 (N_11685,N_11260,N_11216);
xor U11686 (N_11686,N_11378,N_11134);
nand U11687 (N_11687,N_11265,N_11196);
nor U11688 (N_11688,N_11351,N_11049);
nor U11689 (N_11689,N_11407,N_11170);
nor U11690 (N_11690,N_11156,N_11179);
xnor U11691 (N_11691,N_11189,N_11379);
and U11692 (N_11692,N_11474,N_11255);
nor U11693 (N_11693,N_11177,N_11399);
nor U11694 (N_11694,N_11051,N_11492);
nand U11695 (N_11695,N_11408,N_11088);
nor U11696 (N_11696,N_11041,N_11258);
and U11697 (N_11697,N_11200,N_11013);
nand U11698 (N_11698,N_11465,N_11120);
or U11699 (N_11699,N_11208,N_11197);
xor U11700 (N_11700,N_11377,N_11099);
or U11701 (N_11701,N_11029,N_11206);
xnor U11702 (N_11702,N_11104,N_11121);
xnor U11703 (N_11703,N_11066,N_11264);
nand U11704 (N_11704,N_11311,N_11341);
or U11705 (N_11705,N_11141,N_11044);
and U11706 (N_11706,N_11385,N_11367);
and U11707 (N_11707,N_11065,N_11043);
nand U11708 (N_11708,N_11423,N_11023);
nor U11709 (N_11709,N_11280,N_11125);
nor U11710 (N_11710,N_11115,N_11159);
nor U11711 (N_11711,N_11414,N_11016);
nor U11712 (N_11712,N_11470,N_11030);
nor U11713 (N_11713,N_11443,N_11342);
nand U11714 (N_11714,N_11293,N_11009);
nor U11715 (N_11715,N_11145,N_11406);
nor U11716 (N_11716,N_11210,N_11190);
nand U11717 (N_11717,N_11192,N_11098);
nor U11718 (N_11718,N_11238,N_11437);
nor U11719 (N_11719,N_11444,N_11463);
xor U11720 (N_11720,N_11062,N_11296);
and U11721 (N_11721,N_11356,N_11483);
or U11722 (N_11722,N_11137,N_11124);
or U11723 (N_11723,N_11477,N_11109);
or U11724 (N_11724,N_11194,N_11285);
nand U11725 (N_11725,N_11163,N_11332);
nand U11726 (N_11726,N_11439,N_11468);
xnor U11727 (N_11727,N_11295,N_11299);
xnor U11728 (N_11728,N_11061,N_11405);
nand U11729 (N_11729,N_11318,N_11422);
nor U11730 (N_11730,N_11400,N_11246);
and U11731 (N_11731,N_11267,N_11045);
xor U11732 (N_11732,N_11447,N_11010);
or U11733 (N_11733,N_11220,N_11015);
nand U11734 (N_11734,N_11106,N_11107);
or U11735 (N_11735,N_11343,N_11259);
nor U11736 (N_11736,N_11272,N_11226);
or U11737 (N_11737,N_11350,N_11161);
or U11738 (N_11738,N_11059,N_11298);
and U11739 (N_11739,N_11209,N_11151);
nor U11740 (N_11740,N_11431,N_11150);
or U11741 (N_11741,N_11445,N_11388);
nand U11742 (N_11742,N_11224,N_11256);
nand U11743 (N_11743,N_11215,N_11429);
and U11744 (N_11744,N_11193,N_11482);
and U11745 (N_11745,N_11478,N_11320);
or U11746 (N_11746,N_11092,N_11239);
nand U11747 (N_11747,N_11101,N_11128);
nand U11748 (N_11748,N_11186,N_11169);
nor U11749 (N_11749,N_11270,N_11449);
nor U11750 (N_11750,N_11075,N_11298);
xor U11751 (N_11751,N_11115,N_11435);
or U11752 (N_11752,N_11073,N_11344);
xnor U11753 (N_11753,N_11321,N_11000);
nor U11754 (N_11754,N_11047,N_11209);
xor U11755 (N_11755,N_11014,N_11456);
nor U11756 (N_11756,N_11453,N_11053);
or U11757 (N_11757,N_11238,N_11110);
or U11758 (N_11758,N_11456,N_11131);
and U11759 (N_11759,N_11420,N_11318);
and U11760 (N_11760,N_11073,N_11088);
xor U11761 (N_11761,N_11170,N_11209);
or U11762 (N_11762,N_11214,N_11147);
or U11763 (N_11763,N_11333,N_11269);
and U11764 (N_11764,N_11078,N_11199);
nand U11765 (N_11765,N_11492,N_11073);
xor U11766 (N_11766,N_11052,N_11071);
xor U11767 (N_11767,N_11055,N_11223);
xor U11768 (N_11768,N_11448,N_11116);
nor U11769 (N_11769,N_11097,N_11358);
xnor U11770 (N_11770,N_11463,N_11308);
nor U11771 (N_11771,N_11040,N_11169);
and U11772 (N_11772,N_11115,N_11117);
and U11773 (N_11773,N_11103,N_11045);
or U11774 (N_11774,N_11360,N_11448);
nand U11775 (N_11775,N_11186,N_11373);
xnor U11776 (N_11776,N_11099,N_11488);
or U11777 (N_11777,N_11294,N_11174);
and U11778 (N_11778,N_11243,N_11346);
xor U11779 (N_11779,N_11184,N_11470);
nand U11780 (N_11780,N_11388,N_11413);
xnor U11781 (N_11781,N_11029,N_11447);
and U11782 (N_11782,N_11068,N_11412);
and U11783 (N_11783,N_11446,N_11128);
nand U11784 (N_11784,N_11452,N_11105);
nand U11785 (N_11785,N_11322,N_11446);
nand U11786 (N_11786,N_11263,N_11150);
and U11787 (N_11787,N_11285,N_11007);
xor U11788 (N_11788,N_11327,N_11136);
or U11789 (N_11789,N_11068,N_11004);
nor U11790 (N_11790,N_11463,N_11335);
nor U11791 (N_11791,N_11084,N_11385);
and U11792 (N_11792,N_11346,N_11394);
nand U11793 (N_11793,N_11155,N_11490);
nand U11794 (N_11794,N_11082,N_11018);
or U11795 (N_11795,N_11391,N_11372);
nor U11796 (N_11796,N_11212,N_11221);
xor U11797 (N_11797,N_11216,N_11486);
xnor U11798 (N_11798,N_11338,N_11206);
nor U11799 (N_11799,N_11179,N_11432);
xor U11800 (N_11800,N_11143,N_11359);
and U11801 (N_11801,N_11007,N_11485);
and U11802 (N_11802,N_11201,N_11494);
and U11803 (N_11803,N_11031,N_11291);
nand U11804 (N_11804,N_11324,N_11412);
nor U11805 (N_11805,N_11229,N_11178);
or U11806 (N_11806,N_11092,N_11468);
or U11807 (N_11807,N_11365,N_11032);
or U11808 (N_11808,N_11435,N_11143);
and U11809 (N_11809,N_11024,N_11373);
or U11810 (N_11810,N_11009,N_11241);
or U11811 (N_11811,N_11266,N_11134);
or U11812 (N_11812,N_11186,N_11196);
nand U11813 (N_11813,N_11493,N_11150);
xor U11814 (N_11814,N_11190,N_11221);
xor U11815 (N_11815,N_11041,N_11008);
and U11816 (N_11816,N_11419,N_11403);
nor U11817 (N_11817,N_11154,N_11048);
or U11818 (N_11818,N_11408,N_11013);
nor U11819 (N_11819,N_11271,N_11297);
nor U11820 (N_11820,N_11166,N_11134);
nand U11821 (N_11821,N_11226,N_11310);
nand U11822 (N_11822,N_11212,N_11357);
nor U11823 (N_11823,N_11345,N_11231);
xor U11824 (N_11824,N_11034,N_11289);
nor U11825 (N_11825,N_11247,N_11447);
or U11826 (N_11826,N_11435,N_11464);
nand U11827 (N_11827,N_11280,N_11156);
nand U11828 (N_11828,N_11315,N_11458);
nor U11829 (N_11829,N_11156,N_11035);
xor U11830 (N_11830,N_11189,N_11180);
nand U11831 (N_11831,N_11273,N_11431);
nand U11832 (N_11832,N_11284,N_11164);
or U11833 (N_11833,N_11256,N_11113);
nand U11834 (N_11834,N_11442,N_11263);
and U11835 (N_11835,N_11258,N_11194);
and U11836 (N_11836,N_11287,N_11070);
and U11837 (N_11837,N_11019,N_11185);
or U11838 (N_11838,N_11236,N_11039);
nand U11839 (N_11839,N_11245,N_11089);
and U11840 (N_11840,N_11050,N_11454);
or U11841 (N_11841,N_11152,N_11028);
xor U11842 (N_11842,N_11429,N_11005);
or U11843 (N_11843,N_11454,N_11366);
nand U11844 (N_11844,N_11480,N_11261);
nor U11845 (N_11845,N_11482,N_11452);
nand U11846 (N_11846,N_11476,N_11216);
xnor U11847 (N_11847,N_11018,N_11140);
and U11848 (N_11848,N_11046,N_11431);
or U11849 (N_11849,N_11096,N_11293);
and U11850 (N_11850,N_11070,N_11143);
nor U11851 (N_11851,N_11333,N_11145);
and U11852 (N_11852,N_11082,N_11370);
and U11853 (N_11853,N_11062,N_11324);
xnor U11854 (N_11854,N_11414,N_11385);
and U11855 (N_11855,N_11019,N_11133);
nor U11856 (N_11856,N_11056,N_11202);
or U11857 (N_11857,N_11223,N_11476);
nand U11858 (N_11858,N_11219,N_11339);
nand U11859 (N_11859,N_11080,N_11253);
nor U11860 (N_11860,N_11204,N_11355);
nor U11861 (N_11861,N_11494,N_11175);
nor U11862 (N_11862,N_11039,N_11320);
xor U11863 (N_11863,N_11217,N_11473);
nor U11864 (N_11864,N_11203,N_11476);
nor U11865 (N_11865,N_11170,N_11174);
or U11866 (N_11866,N_11487,N_11455);
nand U11867 (N_11867,N_11472,N_11261);
nand U11868 (N_11868,N_11215,N_11014);
xnor U11869 (N_11869,N_11343,N_11193);
nor U11870 (N_11870,N_11021,N_11072);
nand U11871 (N_11871,N_11248,N_11149);
or U11872 (N_11872,N_11176,N_11167);
nand U11873 (N_11873,N_11096,N_11308);
and U11874 (N_11874,N_11172,N_11135);
nor U11875 (N_11875,N_11411,N_11239);
nand U11876 (N_11876,N_11149,N_11454);
xor U11877 (N_11877,N_11200,N_11416);
and U11878 (N_11878,N_11341,N_11361);
nand U11879 (N_11879,N_11433,N_11261);
or U11880 (N_11880,N_11484,N_11363);
xor U11881 (N_11881,N_11309,N_11276);
or U11882 (N_11882,N_11267,N_11041);
or U11883 (N_11883,N_11393,N_11131);
nand U11884 (N_11884,N_11352,N_11160);
nor U11885 (N_11885,N_11028,N_11005);
and U11886 (N_11886,N_11356,N_11349);
nand U11887 (N_11887,N_11265,N_11038);
nor U11888 (N_11888,N_11455,N_11052);
nor U11889 (N_11889,N_11485,N_11424);
xnor U11890 (N_11890,N_11481,N_11248);
and U11891 (N_11891,N_11114,N_11139);
xnor U11892 (N_11892,N_11117,N_11324);
xnor U11893 (N_11893,N_11404,N_11435);
nand U11894 (N_11894,N_11369,N_11081);
xor U11895 (N_11895,N_11415,N_11256);
nand U11896 (N_11896,N_11009,N_11351);
nand U11897 (N_11897,N_11125,N_11055);
or U11898 (N_11898,N_11193,N_11249);
nand U11899 (N_11899,N_11420,N_11131);
xnor U11900 (N_11900,N_11452,N_11182);
nand U11901 (N_11901,N_11137,N_11387);
or U11902 (N_11902,N_11384,N_11203);
and U11903 (N_11903,N_11251,N_11063);
nand U11904 (N_11904,N_11082,N_11286);
and U11905 (N_11905,N_11235,N_11487);
or U11906 (N_11906,N_11327,N_11428);
nand U11907 (N_11907,N_11477,N_11277);
and U11908 (N_11908,N_11396,N_11179);
xnor U11909 (N_11909,N_11064,N_11097);
or U11910 (N_11910,N_11049,N_11250);
xor U11911 (N_11911,N_11051,N_11324);
or U11912 (N_11912,N_11453,N_11164);
xnor U11913 (N_11913,N_11135,N_11091);
nor U11914 (N_11914,N_11130,N_11370);
or U11915 (N_11915,N_11235,N_11480);
nor U11916 (N_11916,N_11405,N_11244);
xor U11917 (N_11917,N_11077,N_11028);
nor U11918 (N_11918,N_11491,N_11391);
and U11919 (N_11919,N_11388,N_11371);
or U11920 (N_11920,N_11284,N_11036);
or U11921 (N_11921,N_11179,N_11144);
xnor U11922 (N_11922,N_11099,N_11402);
xnor U11923 (N_11923,N_11122,N_11105);
nand U11924 (N_11924,N_11489,N_11290);
nor U11925 (N_11925,N_11182,N_11200);
xor U11926 (N_11926,N_11413,N_11079);
and U11927 (N_11927,N_11051,N_11323);
xor U11928 (N_11928,N_11156,N_11314);
nor U11929 (N_11929,N_11498,N_11423);
and U11930 (N_11930,N_11014,N_11405);
and U11931 (N_11931,N_11237,N_11487);
xnor U11932 (N_11932,N_11102,N_11394);
nor U11933 (N_11933,N_11117,N_11230);
and U11934 (N_11934,N_11460,N_11400);
xnor U11935 (N_11935,N_11037,N_11093);
xnor U11936 (N_11936,N_11201,N_11370);
nand U11937 (N_11937,N_11363,N_11469);
nand U11938 (N_11938,N_11308,N_11085);
and U11939 (N_11939,N_11071,N_11056);
nand U11940 (N_11940,N_11467,N_11197);
nand U11941 (N_11941,N_11246,N_11116);
nand U11942 (N_11942,N_11403,N_11277);
xnor U11943 (N_11943,N_11007,N_11411);
nand U11944 (N_11944,N_11248,N_11406);
xnor U11945 (N_11945,N_11216,N_11073);
or U11946 (N_11946,N_11249,N_11367);
xnor U11947 (N_11947,N_11169,N_11445);
nand U11948 (N_11948,N_11176,N_11442);
or U11949 (N_11949,N_11281,N_11080);
xnor U11950 (N_11950,N_11388,N_11135);
xor U11951 (N_11951,N_11127,N_11169);
nand U11952 (N_11952,N_11498,N_11079);
nand U11953 (N_11953,N_11212,N_11133);
or U11954 (N_11954,N_11497,N_11014);
nand U11955 (N_11955,N_11044,N_11339);
or U11956 (N_11956,N_11035,N_11217);
nor U11957 (N_11957,N_11061,N_11278);
xor U11958 (N_11958,N_11462,N_11145);
xnor U11959 (N_11959,N_11391,N_11138);
xnor U11960 (N_11960,N_11024,N_11173);
or U11961 (N_11961,N_11360,N_11498);
xor U11962 (N_11962,N_11194,N_11025);
nor U11963 (N_11963,N_11076,N_11193);
xor U11964 (N_11964,N_11080,N_11003);
xor U11965 (N_11965,N_11137,N_11030);
nor U11966 (N_11966,N_11104,N_11250);
xor U11967 (N_11967,N_11319,N_11406);
and U11968 (N_11968,N_11303,N_11007);
or U11969 (N_11969,N_11359,N_11144);
or U11970 (N_11970,N_11056,N_11313);
xnor U11971 (N_11971,N_11015,N_11032);
nand U11972 (N_11972,N_11095,N_11156);
or U11973 (N_11973,N_11428,N_11278);
xnor U11974 (N_11974,N_11092,N_11395);
nand U11975 (N_11975,N_11268,N_11404);
xor U11976 (N_11976,N_11029,N_11376);
and U11977 (N_11977,N_11336,N_11471);
nand U11978 (N_11978,N_11018,N_11239);
nor U11979 (N_11979,N_11049,N_11493);
or U11980 (N_11980,N_11289,N_11023);
nor U11981 (N_11981,N_11429,N_11148);
or U11982 (N_11982,N_11184,N_11301);
or U11983 (N_11983,N_11189,N_11218);
nand U11984 (N_11984,N_11148,N_11267);
and U11985 (N_11985,N_11000,N_11487);
nor U11986 (N_11986,N_11038,N_11169);
xor U11987 (N_11987,N_11380,N_11215);
nand U11988 (N_11988,N_11110,N_11072);
and U11989 (N_11989,N_11437,N_11341);
nand U11990 (N_11990,N_11280,N_11410);
or U11991 (N_11991,N_11222,N_11465);
and U11992 (N_11992,N_11008,N_11421);
nand U11993 (N_11993,N_11315,N_11014);
nor U11994 (N_11994,N_11180,N_11351);
xor U11995 (N_11995,N_11456,N_11470);
and U11996 (N_11996,N_11413,N_11178);
nor U11997 (N_11997,N_11343,N_11330);
and U11998 (N_11998,N_11030,N_11052);
xor U11999 (N_11999,N_11459,N_11221);
xor U12000 (N_12000,N_11618,N_11791);
nand U12001 (N_12001,N_11823,N_11611);
xnor U12002 (N_12002,N_11686,N_11723);
or U12003 (N_12003,N_11673,N_11911);
nand U12004 (N_12004,N_11832,N_11716);
nor U12005 (N_12005,N_11822,N_11523);
or U12006 (N_12006,N_11806,N_11601);
or U12007 (N_12007,N_11691,N_11811);
nand U12008 (N_12008,N_11758,N_11631);
xnor U12009 (N_12009,N_11545,N_11574);
nand U12010 (N_12010,N_11831,N_11995);
xnor U12011 (N_12011,N_11794,N_11533);
nand U12012 (N_12012,N_11827,N_11935);
and U12013 (N_12013,N_11527,N_11625);
nor U12014 (N_12014,N_11514,N_11848);
nand U12015 (N_12015,N_11540,N_11513);
and U12016 (N_12016,N_11619,N_11666);
xnor U12017 (N_12017,N_11500,N_11539);
or U12018 (N_12018,N_11706,N_11603);
nand U12019 (N_12019,N_11924,N_11787);
nand U12020 (N_12020,N_11947,N_11524);
or U12021 (N_12021,N_11685,N_11897);
nand U12022 (N_12022,N_11595,N_11970);
nor U12023 (N_12023,N_11896,N_11607);
nor U12024 (N_12024,N_11663,N_11845);
nor U12025 (N_12025,N_11857,N_11866);
and U12026 (N_12026,N_11665,N_11775);
nand U12027 (N_12027,N_11708,N_11839);
or U12028 (N_12028,N_11739,N_11677);
and U12029 (N_12029,N_11749,N_11735);
and U12030 (N_12030,N_11833,N_11696);
nand U12031 (N_12031,N_11629,N_11988);
nand U12032 (N_12032,N_11541,N_11772);
nand U12033 (N_12033,N_11846,N_11905);
xnor U12034 (N_12034,N_11626,N_11765);
xnor U12035 (N_12035,N_11678,N_11843);
xnor U12036 (N_12036,N_11732,N_11519);
or U12037 (N_12037,N_11713,N_11585);
nor U12038 (N_12038,N_11930,N_11768);
or U12039 (N_12039,N_11759,N_11565);
and U12040 (N_12040,N_11805,N_11676);
xnor U12041 (N_12041,N_11633,N_11801);
xor U12042 (N_12042,N_11987,N_11655);
nor U12043 (N_12043,N_11920,N_11694);
or U12044 (N_12044,N_11721,N_11756);
nor U12045 (N_12045,N_11570,N_11720);
xor U12046 (N_12046,N_11628,N_11544);
nor U12047 (N_12047,N_11581,N_11999);
or U12048 (N_12048,N_11737,N_11647);
nand U12049 (N_12049,N_11571,N_11838);
and U12050 (N_12050,N_11926,N_11908);
and U12051 (N_12051,N_11914,N_11651);
nor U12052 (N_12052,N_11815,N_11637);
or U12053 (N_12053,N_11669,N_11909);
nor U12054 (N_12054,N_11847,N_11824);
or U12055 (N_12055,N_11931,N_11900);
or U12056 (N_12056,N_11818,N_11979);
nor U12057 (N_12057,N_11622,N_11837);
and U12058 (N_12058,N_11809,N_11980);
or U12059 (N_12059,N_11736,N_11933);
xnor U12060 (N_12060,N_11521,N_11813);
xor U12061 (N_12061,N_11958,N_11741);
or U12062 (N_12062,N_11657,N_11556);
or U12063 (N_12063,N_11899,N_11877);
and U12064 (N_12064,N_11512,N_11971);
xor U12065 (N_12065,N_11841,N_11821);
or U12066 (N_12066,N_11653,N_11638);
and U12067 (N_12067,N_11798,N_11714);
xnor U12068 (N_12068,N_11754,N_11826);
nor U12069 (N_12069,N_11510,N_11985);
or U12070 (N_12070,N_11589,N_11766);
and U12071 (N_12071,N_11921,N_11803);
xnor U12072 (N_12072,N_11812,N_11779);
and U12073 (N_12073,N_11748,N_11690);
and U12074 (N_12074,N_11733,N_11855);
and U12075 (N_12075,N_11851,N_11769);
or U12076 (N_12076,N_11623,N_11726);
xnor U12077 (N_12077,N_11904,N_11817);
nand U12078 (N_12078,N_11644,N_11557);
and U12079 (N_12079,N_11796,N_11982);
xnor U12080 (N_12080,N_11918,N_11760);
xnor U12081 (N_12081,N_11927,N_11871);
xor U12082 (N_12082,N_11828,N_11861);
xnor U12083 (N_12083,N_11661,N_11802);
and U12084 (N_12084,N_11808,N_11517);
and U12085 (N_12085,N_11879,N_11569);
xnor U12086 (N_12086,N_11604,N_11542);
and U12087 (N_12087,N_11525,N_11778);
and U12088 (N_12088,N_11800,N_11887);
and U12089 (N_12089,N_11888,N_11953);
nand U12090 (N_12090,N_11964,N_11627);
nor U12091 (N_12091,N_11770,N_11998);
or U12092 (N_12092,N_11789,N_11782);
xor U12093 (N_12093,N_11816,N_11873);
xnor U12094 (N_12094,N_11608,N_11575);
nand U12095 (N_12095,N_11950,N_11865);
xor U12096 (N_12096,N_11504,N_11858);
nand U12097 (N_12097,N_11693,N_11698);
or U12098 (N_12098,N_11610,N_11767);
xor U12099 (N_12099,N_11674,N_11515);
nand U12100 (N_12100,N_11591,N_11670);
xnor U12101 (N_12101,N_11790,N_11548);
nor U12102 (N_12102,N_11849,N_11606);
xnor U12103 (N_12103,N_11901,N_11695);
or U12104 (N_12104,N_11856,N_11639);
nor U12105 (N_12105,N_11593,N_11543);
nand U12106 (N_12106,N_11889,N_11939);
xnor U12107 (N_12107,N_11773,N_11505);
and U12108 (N_12108,N_11878,N_11859);
nor U12109 (N_12109,N_11885,N_11867);
nor U12110 (N_12110,N_11614,N_11617);
and U12111 (N_12111,N_11654,N_11916);
or U12112 (N_12112,N_11938,N_11600);
xor U12113 (N_12113,N_11943,N_11783);
xor U12114 (N_12114,N_11962,N_11937);
nor U12115 (N_12115,N_11854,N_11531);
xnor U12116 (N_12116,N_11605,N_11876);
xnor U12117 (N_12117,N_11940,N_11649);
nor U12118 (N_12118,N_11648,N_11566);
xor U12119 (N_12119,N_11738,N_11990);
xor U12120 (N_12120,N_11560,N_11704);
or U12121 (N_12121,N_11630,N_11946);
and U12122 (N_12122,N_11799,N_11751);
nand U12123 (N_12123,N_11573,N_11744);
nand U12124 (N_12124,N_11536,N_11810);
nand U12125 (N_12125,N_11797,N_11983);
and U12126 (N_12126,N_11786,N_11973);
nor U12127 (N_12127,N_11898,N_11840);
and U12128 (N_12128,N_11688,N_11780);
nand U12129 (N_12129,N_11547,N_11699);
and U12130 (N_12130,N_11596,N_11507);
xnor U12131 (N_12131,N_11715,N_11534);
or U12132 (N_12132,N_11740,N_11532);
nand U12133 (N_12133,N_11568,N_11894);
or U12134 (N_12134,N_11961,N_11893);
and U12135 (N_12135,N_11597,N_11615);
nor U12136 (N_12136,N_11850,N_11977);
nor U12137 (N_12137,N_11872,N_11522);
nor U12138 (N_12138,N_11520,N_11928);
nor U12139 (N_12139,N_11718,N_11612);
nor U12140 (N_12140,N_11529,N_11771);
or U12141 (N_12141,N_11645,N_11819);
nor U12142 (N_12142,N_11884,N_11701);
or U12143 (N_12143,N_11755,N_11503);
nand U12144 (N_12144,N_11717,N_11853);
nand U12145 (N_12145,N_11672,N_11886);
nor U12146 (N_12146,N_11864,N_11616);
and U12147 (N_12147,N_11729,N_11577);
nand U12148 (N_12148,N_11588,N_11746);
nand U12149 (N_12149,N_11852,N_11662);
or U12150 (N_12150,N_11963,N_11640);
nor U12151 (N_12151,N_11907,N_11558);
and U12152 (N_12152,N_11697,N_11793);
nand U12153 (N_12153,N_11679,N_11609);
nor U12154 (N_12154,N_11700,N_11820);
or U12155 (N_12155,N_11795,N_11981);
nor U12156 (N_12156,N_11883,N_11863);
or U12157 (N_12157,N_11646,N_11579);
xor U12158 (N_12158,N_11881,N_11763);
or U12159 (N_12159,N_11702,N_11842);
nand U12160 (N_12160,N_11643,N_11502);
and U12161 (N_12161,N_11613,N_11922);
nand U12162 (N_12162,N_11870,N_11632);
or U12163 (N_12163,N_11967,N_11890);
and U12164 (N_12164,N_11621,N_11976);
xor U12165 (N_12165,N_11902,N_11882);
or U12166 (N_12166,N_11903,N_11705);
nand U12167 (N_12167,N_11572,N_11978);
nand U12168 (N_12168,N_11844,N_11682);
xor U12169 (N_12169,N_11551,N_11762);
nand U12170 (N_12170,N_11975,N_11664);
and U12171 (N_12171,N_11993,N_11804);
nand U12172 (N_12172,N_11750,N_11835);
xnor U12173 (N_12173,N_11582,N_11658);
and U12174 (N_12174,N_11745,N_11917);
and U12175 (N_12175,N_11722,N_11761);
xnor U12176 (N_12176,N_11683,N_11776);
xor U12177 (N_12177,N_11501,N_11731);
and U12178 (N_12178,N_11511,N_11537);
nand U12179 (N_12179,N_11635,N_11952);
and U12180 (N_12180,N_11587,N_11956);
xnor U12181 (N_12181,N_11709,N_11836);
xnor U12182 (N_12182,N_11586,N_11969);
or U12183 (N_12183,N_11730,N_11652);
nor U12184 (N_12184,N_11974,N_11727);
nor U12185 (N_12185,N_11968,N_11792);
and U12186 (N_12186,N_11689,N_11668);
nor U12187 (N_12187,N_11594,N_11526);
or U12188 (N_12188,N_11659,N_11561);
or U12189 (N_12189,N_11874,N_11546);
xnor U12190 (N_12190,N_11925,N_11602);
and U12191 (N_12191,N_11530,N_11707);
and U12192 (N_12192,N_11675,N_11862);
or U12193 (N_12193,N_11860,N_11687);
nand U12194 (N_12194,N_11583,N_11642);
xor U12195 (N_12195,N_11554,N_11915);
and U12196 (N_12196,N_11564,N_11936);
and U12197 (N_12197,N_11660,N_11681);
and U12198 (N_12198,N_11991,N_11725);
or U12199 (N_12199,N_11757,N_11892);
xor U12200 (N_12200,N_11984,N_11559);
nor U12201 (N_12201,N_11923,N_11788);
nand U12202 (N_12202,N_11951,N_11567);
xnor U12203 (N_12203,N_11948,N_11552);
and U12204 (N_12204,N_11747,N_11580);
xnor U12205 (N_12205,N_11880,N_11562);
and U12206 (N_12206,N_11703,N_11919);
xnor U12207 (N_12207,N_11590,N_11667);
xor U12208 (N_12208,N_11986,N_11641);
nand U12209 (N_12209,N_11549,N_11868);
xor U12210 (N_12210,N_11781,N_11656);
nand U12211 (N_12211,N_11620,N_11734);
nand U12212 (N_12212,N_11728,N_11997);
or U12213 (N_12213,N_11711,N_11650);
nor U12214 (N_12214,N_11960,N_11784);
nor U12215 (N_12215,N_11509,N_11671);
nor U12216 (N_12216,N_11989,N_11825);
or U12217 (N_12217,N_11774,N_11829);
nor U12218 (N_12218,N_11814,N_11941);
xor U12219 (N_12219,N_11949,N_11834);
xor U12220 (N_12220,N_11553,N_11724);
nand U12221 (N_12221,N_11555,N_11891);
and U12222 (N_12222,N_11910,N_11680);
nand U12223 (N_12223,N_11996,N_11692);
and U12224 (N_12224,N_11752,N_11636);
or U12225 (N_12225,N_11753,N_11584);
or U12226 (N_12226,N_11785,N_11966);
or U12227 (N_12227,N_11550,N_11875);
nand U12228 (N_12228,N_11576,N_11895);
or U12229 (N_12229,N_11506,N_11592);
nor U12230 (N_12230,N_11598,N_11972);
xor U12231 (N_12231,N_11710,N_11764);
nand U12232 (N_12232,N_11807,N_11992);
and U12233 (N_12233,N_11955,N_11954);
nand U12234 (N_12234,N_11912,N_11624);
xnor U12235 (N_12235,N_11934,N_11959);
nor U12236 (N_12236,N_11777,N_11944);
and U12237 (N_12237,N_11719,N_11913);
xnor U12238 (N_12238,N_11528,N_11538);
nand U12239 (N_12239,N_11942,N_11563);
nand U12240 (N_12240,N_11965,N_11957);
nand U12241 (N_12241,N_11712,N_11599);
nand U12242 (N_12242,N_11906,N_11932);
xnor U12243 (N_12243,N_11518,N_11634);
xor U12244 (N_12244,N_11994,N_11945);
and U12245 (N_12245,N_11535,N_11929);
nor U12246 (N_12246,N_11742,N_11516);
nand U12247 (N_12247,N_11869,N_11743);
nor U12248 (N_12248,N_11684,N_11508);
xor U12249 (N_12249,N_11578,N_11830);
nand U12250 (N_12250,N_11725,N_11866);
nor U12251 (N_12251,N_11542,N_11830);
and U12252 (N_12252,N_11912,N_11844);
nor U12253 (N_12253,N_11954,N_11626);
and U12254 (N_12254,N_11749,N_11565);
nor U12255 (N_12255,N_11534,N_11526);
xor U12256 (N_12256,N_11604,N_11737);
xor U12257 (N_12257,N_11500,N_11894);
nand U12258 (N_12258,N_11817,N_11905);
and U12259 (N_12259,N_11738,N_11924);
and U12260 (N_12260,N_11554,N_11727);
nand U12261 (N_12261,N_11936,N_11935);
nand U12262 (N_12262,N_11867,N_11512);
nand U12263 (N_12263,N_11549,N_11853);
nor U12264 (N_12264,N_11667,N_11947);
nand U12265 (N_12265,N_11745,N_11596);
or U12266 (N_12266,N_11772,N_11911);
nand U12267 (N_12267,N_11698,N_11733);
nand U12268 (N_12268,N_11670,N_11683);
and U12269 (N_12269,N_11838,N_11979);
or U12270 (N_12270,N_11825,N_11631);
nand U12271 (N_12271,N_11746,N_11994);
nand U12272 (N_12272,N_11682,N_11836);
nor U12273 (N_12273,N_11966,N_11849);
or U12274 (N_12274,N_11774,N_11979);
or U12275 (N_12275,N_11763,N_11686);
and U12276 (N_12276,N_11508,N_11647);
nor U12277 (N_12277,N_11921,N_11900);
nor U12278 (N_12278,N_11818,N_11753);
nor U12279 (N_12279,N_11659,N_11746);
or U12280 (N_12280,N_11786,N_11948);
and U12281 (N_12281,N_11716,N_11534);
nand U12282 (N_12282,N_11620,N_11559);
nor U12283 (N_12283,N_11806,N_11598);
or U12284 (N_12284,N_11934,N_11915);
nand U12285 (N_12285,N_11980,N_11534);
xor U12286 (N_12286,N_11798,N_11732);
nand U12287 (N_12287,N_11556,N_11983);
xor U12288 (N_12288,N_11618,N_11654);
nor U12289 (N_12289,N_11789,N_11778);
and U12290 (N_12290,N_11835,N_11575);
nand U12291 (N_12291,N_11640,N_11574);
and U12292 (N_12292,N_11712,N_11519);
nand U12293 (N_12293,N_11569,N_11578);
and U12294 (N_12294,N_11893,N_11737);
and U12295 (N_12295,N_11819,N_11657);
nor U12296 (N_12296,N_11803,N_11537);
nand U12297 (N_12297,N_11827,N_11565);
and U12298 (N_12298,N_11899,N_11984);
nand U12299 (N_12299,N_11579,N_11703);
and U12300 (N_12300,N_11613,N_11527);
and U12301 (N_12301,N_11868,N_11615);
or U12302 (N_12302,N_11896,N_11602);
xnor U12303 (N_12303,N_11633,N_11942);
nand U12304 (N_12304,N_11602,N_11754);
xor U12305 (N_12305,N_11675,N_11512);
nor U12306 (N_12306,N_11548,N_11742);
or U12307 (N_12307,N_11854,N_11935);
and U12308 (N_12308,N_11579,N_11707);
nor U12309 (N_12309,N_11612,N_11972);
nand U12310 (N_12310,N_11669,N_11546);
nand U12311 (N_12311,N_11927,N_11888);
xnor U12312 (N_12312,N_11594,N_11602);
nand U12313 (N_12313,N_11640,N_11711);
nand U12314 (N_12314,N_11825,N_11914);
nand U12315 (N_12315,N_11985,N_11516);
xnor U12316 (N_12316,N_11822,N_11600);
nor U12317 (N_12317,N_11733,N_11511);
or U12318 (N_12318,N_11843,N_11735);
and U12319 (N_12319,N_11877,N_11638);
xor U12320 (N_12320,N_11983,N_11922);
xnor U12321 (N_12321,N_11899,N_11665);
or U12322 (N_12322,N_11559,N_11610);
nand U12323 (N_12323,N_11520,N_11999);
xor U12324 (N_12324,N_11855,N_11555);
or U12325 (N_12325,N_11625,N_11532);
nor U12326 (N_12326,N_11783,N_11562);
xnor U12327 (N_12327,N_11704,N_11510);
and U12328 (N_12328,N_11602,N_11800);
xor U12329 (N_12329,N_11919,N_11982);
or U12330 (N_12330,N_11781,N_11583);
nor U12331 (N_12331,N_11783,N_11518);
xnor U12332 (N_12332,N_11686,N_11792);
nor U12333 (N_12333,N_11903,N_11622);
nand U12334 (N_12334,N_11867,N_11870);
xor U12335 (N_12335,N_11753,N_11721);
or U12336 (N_12336,N_11789,N_11619);
or U12337 (N_12337,N_11669,N_11626);
or U12338 (N_12338,N_11987,N_11760);
xor U12339 (N_12339,N_11977,N_11570);
or U12340 (N_12340,N_11871,N_11945);
xor U12341 (N_12341,N_11508,N_11968);
nand U12342 (N_12342,N_11729,N_11908);
nor U12343 (N_12343,N_11775,N_11703);
and U12344 (N_12344,N_11988,N_11868);
xor U12345 (N_12345,N_11940,N_11563);
nor U12346 (N_12346,N_11826,N_11670);
or U12347 (N_12347,N_11568,N_11773);
and U12348 (N_12348,N_11996,N_11556);
nor U12349 (N_12349,N_11787,N_11755);
nand U12350 (N_12350,N_11611,N_11797);
or U12351 (N_12351,N_11747,N_11663);
nand U12352 (N_12352,N_11867,N_11614);
nand U12353 (N_12353,N_11637,N_11534);
nor U12354 (N_12354,N_11756,N_11969);
nor U12355 (N_12355,N_11562,N_11844);
and U12356 (N_12356,N_11562,N_11652);
nor U12357 (N_12357,N_11583,N_11975);
nand U12358 (N_12358,N_11677,N_11941);
xor U12359 (N_12359,N_11893,N_11936);
nand U12360 (N_12360,N_11742,N_11833);
or U12361 (N_12361,N_11800,N_11959);
xor U12362 (N_12362,N_11506,N_11750);
nor U12363 (N_12363,N_11633,N_11957);
or U12364 (N_12364,N_11906,N_11664);
nor U12365 (N_12365,N_11938,N_11768);
or U12366 (N_12366,N_11777,N_11955);
xnor U12367 (N_12367,N_11939,N_11866);
nand U12368 (N_12368,N_11739,N_11710);
nand U12369 (N_12369,N_11683,N_11613);
and U12370 (N_12370,N_11684,N_11871);
or U12371 (N_12371,N_11710,N_11695);
or U12372 (N_12372,N_11610,N_11561);
and U12373 (N_12373,N_11767,N_11678);
nand U12374 (N_12374,N_11707,N_11735);
xnor U12375 (N_12375,N_11914,N_11922);
or U12376 (N_12376,N_11753,N_11904);
xor U12377 (N_12377,N_11772,N_11548);
xnor U12378 (N_12378,N_11832,N_11539);
xnor U12379 (N_12379,N_11941,N_11994);
xnor U12380 (N_12380,N_11537,N_11798);
and U12381 (N_12381,N_11511,N_11702);
and U12382 (N_12382,N_11547,N_11857);
and U12383 (N_12383,N_11569,N_11720);
nor U12384 (N_12384,N_11543,N_11856);
and U12385 (N_12385,N_11576,N_11667);
nand U12386 (N_12386,N_11741,N_11606);
and U12387 (N_12387,N_11718,N_11735);
or U12388 (N_12388,N_11873,N_11844);
xnor U12389 (N_12389,N_11596,N_11865);
nor U12390 (N_12390,N_11530,N_11669);
xnor U12391 (N_12391,N_11741,N_11645);
nor U12392 (N_12392,N_11695,N_11921);
nand U12393 (N_12393,N_11915,N_11955);
nand U12394 (N_12394,N_11908,N_11648);
xnor U12395 (N_12395,N_11854,N_11791);
and U12396 (N_12396,N_11940,N_11696);
nor U12397 (N_12397,N_11835,N_11565);
and U12398 (N_12398,N_11939,N_11673);
nor U12399 (N_12399,N_11593,N_11781);
nand U12400 (N_12400,N_11727,N_11562);
or U12401 (N_12401,N_11532,N_11676);
nand U12402 (N_12402,N_11717,N_11671);
xnor U12403 (N_12403,N_11976,N_11872);
and U12404 (N_12404,N_11564,N_11921);
nor U12405 (N_12405,N_11810,N_11900);
and U12406 (N_12406,N_11503,N_11913);
xnor U12407 (N_12407,N_11604,N_11721);
and U12408 (N_12408,N_11536,N_11668);
nand U12409 (N_12409,N_11960,N_11855);
and U12410 (N_12410,N_11820,N_11585);
and U12411 (N_12411,N_11998,N_11663);
nor U12412 (N_12412,N_11908,N_11886);
or U12413 (N_12413,N_11628,N_11820);
and U12414 (N_12414,N_11968,N_11908);
nor U12415 (N_12415,N_11535,N_11848);
nor U12416 (N_12416,N_11742,N_11827);
nand U12417 (N_12417,N_11977,N_11623);
and U12418 (N_12418,N_11968,N_11754);
nor U12419 (N_12419,N_11824,N_11926);
and U12420 (N_12420,N_11983,N_11638);
and U12421 (N_12421,N_11713,N_11529);
and U12422 (N_12422,N_11737,N_11628);
and U12423 (N_12423,N_11554,N_11728);
nand U12424 (N_12424,N_11721,N_11922);
xor U12425 (N_12425,N_11809,N_11586);
or U12426 (N_12426,N_11585,N_11901);
or U12427 (N_12427,N_11899,N_11736);
or U12428 (N_12428,N_11806,N_11667);
nor U12429 (N_12429,N_11641,N_11981);
xor U12430 (N_12430,N_11607,N_11511);
or U12431 (N_12431,N_11874,N_11730);
xnor U12432 (N_12432,N_11697,N_11594);
nor U12433 (N_12433,N_11672,N_11846);
xnor U12434 (N_12434,N_11756,N_11906);
or U12435 (N_12435,N_11647,N_11517);
nor U12436 (N_12436,N_11890,N_11753);
nor U12437 (N_12437,N_11715,N_11812);
nor U12438 (N_12438,N_11970,N_11628);
xnor U12439 (N_12439,N_11722,N_11833);
nor U12440 (N_12440,N_11646,N_11614);
xor U12441 (N_12441,N_11717,N_11774);
nand U12442 (N_12442,N_11676,N_11951);
xor U12443 (N_12443,N_11839,N_11802);
nand U12444 (N_12444,N_11509,N_11534);
or U12445 (N_12445,N_11925,N_11541);
xor U12446 (N_12446,N_11586,N_11580);
and U12447 (N_12447,N_11639,N_11530);
or U12448 (N_12448,N_11939,N_11804);
or U12449 (N_12449,N_11856,N_11981);
or U12450 (N_12450,N_11799,N_11742);
or U12451 (N_12451,N_11872,N_11627);
and U12452 (N_12452,N_11867,N_11703);
nor U12453 (N_12453,N_11758,N_11509);
or U12454 (N_12454,N_11583,N_11541);
nand U12455 (N_12455,N_11839,N_11901);
xor U12456 (N_12456,N_11771,N_11945);
nand U12457 (N_12457,N_11900,N_11880);
nor U12458 (N_12458,N_11962,N_11880);
nand U12459 (N_12459,N_11869,N_11962);
or U12460 (N_12460,N_11788,N_11999);
xor U12461 (N_12461,N_11714,N_11634);
xnor U12462 (N_12462,N_11807,N_11842);
nor U12463 (N_12463,N_11841,N_11592);
nor U12464 (N_12464,N_11830,N_11548);
nor U12465 (N_12465,N_11792,N_11755);
nor U12466 (N_12466,N_11770,N_11559);
and U12467 (N_12467,N_11947,N_11669);
nand U12468 (N_12468,N_11947,N_11869);
nand U12469 (N_12469,N_11922,N_11985);
nor U12470 (N_12470,N_11940,N_11566);
and U12471 (N_12471,N_11926,N_11910);
or U12472 (N_12472,N_11805,N_11553);
nand U12473 (N_12473,N_11501,N_11653);
nor U12474 (N_12474,N_11876,N_11987);
and U12475 (N_12475,N_11850,N_11821);
xnor U12476 (N_12476,N_11582,N_11510);
nor U12477 (N_12477,N_11689,N_11605);
nand U12478 (N_12478,N_11858,N_11935);
and U12479 (N_12479,N_11905,N_11781);
or U12480 (N_12480,N_11782,N_11742);
or U12481 (N_12481,N_11918,N_11555);
and U12482 (N_12482,N_11701,N_11896);
or U12483 (N_12483,N_11917,N_11502);
and U12484 (N_12484,N_11950,N_11560);
nor U12485 (N_12485,N_11930,N_11651);
and U12486 (N_12486,N_11656,N_11705);
nor U12487 (N_12487,N_11961,N_11635);
or U12488 (N_12488,N_11879,N_11896);
nor U12489 (N_12489,N_11822,N_11869);
xnor U12490 (N_12490,N_11662,N_11715);
or U12491 (N_12491,N_11634,N_11748);
and U12492 (N_12492,N_11811,N_11692);
nand U12493 (N_12493,N_11922,N_11882);
nand U12494 (N_12494,N_11709,N_11547);
or U12495 (N_12495,N_11659,N_11694);
and U12496 (N_12496,N_11787,N_11728);
or U12497 (N_12497,N_11939,N_11698);
and U12498 (N_12498,N_11771,N_11577);
xor U12499 (N_12499,N_11524,N_11552);
nor U12500 (N_12500,N_12155,N_12245);
or U12501 (N_12501,N_12394,N_12139);
or U12502 (N_12502,N_12439,N_12246);
xnor U12503 (N_12503,N_12190,N_12038);
nand U12504 (N_12504,N_12170,N_12168);
xnor U12505 (N_12505,N_12127,N_12290);
or U12506 (N_12506,N_12288,N_12000);
nor U12507 (N_12507,N_12276,N_12418);
nand U12508 (N_12508,N_12129,N_12470);
nand U12509 (N_12509,N_12485,N_12272);
nor U12510 (N_12510,N_12396,N_12091);
xnor U12511 (N_12511,N_12344,N_12187);
nand U12512 (N_12512,N_12199,N_12298);
xnor U12513 (N_12513,N_12277,N_12071);
nand U12514 (N_12514,N_12269,N_12119);
nand U12515 (N_12515,N_12350,N_12032);
and U12516 (N_12516,N_12186,N_12236);
nand U12517 (N_12517,N_12058,N_12002);
or U12518 (N_12518,N_12413,N_12135);
nand U12519 (N_12519,N_12082,N_12251);
and U12520 (N_12520,N_12178,N_12469);
nor U12521 (N_12521,N_12339,N_12005);
nand U12522 (N_12522,N_12393,N_12435);
or U12523 (N_12523,N_12432,N_12254);
nor U12524 (N_12524,N_12315,N_12067);
and U12525 (N_12525,N_12208,N_12025);
nor U12526 (N_12526,N_12030,N_12084);
or U12527 (N_12527,N_12447,N_12281);
or U12528 (N_12528,N_12222,N_12039);
xnor U12529 (N_12529,N_12337,N_12090);
nor U12530 (N_12530,N_12059,N_12402);
nor U12531 (N_12531,N_12473,N_12318);
and U12532 (N_12532,N_12335,N_12361);
nor U12533 (N_12533,N_12427,N_12358);
or U12534 (N_12534,N_12471,N_12107);
nor U12535 (N_12535,N_12184,N_12438);
and U12536 (N_12536,N_12087,N_12064);
nor U12537 (N_12537,N_12003,N_12467);
or U12538 (N_12538,N_12089,N_12121);
and U12539 (N_12539,N_12468,N_12444);
nor U12540 (N_12540,N_12264,N_12301);
or U12541 (N_12541,N_12144,N_12492);
or U12542 (N_12542,N_12282,N_12386);
xor U12543 (N_12543,N_12412,N_12248);
and U12544 (N_12544,N_12179,N_12283);
xnor U12545 (N_12545,N_12211,N_12227);
or U12546 (N_12546,N_12011,N_12406);
and U12547 (N_12547,N_12371,N_12325);
xnor U12548 (N_12548,N_12451,N_12268);
nor U12549 (N_12549,N_12183,N_12150);
or U12550 (N_12550,N_12065,N_12161);
and U12551 (N_12551,N_12314,N_12271);
and U12552 (N_12552,N_12052,N_12378);
and U12553 (N_12553,N_12247,N_12464);
and U12554 (N_12554,N_12196,N_12200);
or U12555 (N_12555,N_12345,N_12053);
and U12556 (N_12556,N_12327,N_12321);
and U12557 (N_12557,N_12255,N_12369);
nor U12558 (N_12558,N_12173,N_12426);
or U12559 (N_12559,N_12416,N_12115);
and U12560 (N_12560,N_12037,N_12031);
or U12561 (N_12561,N_12049,N_12017);
xor U12562 (N_12562,N_12098,N_12220);
and U12563 (N_12563,N_12232,N_12195);
and U12564 (N_12564,N_12312,N_12258);
and U12565 (N_12565,N_12384,N_12275);
xor U12566 (N_12566,N_12180,N_12128);
nor U12567 (N_12567,N_12273,N_12289);
or U12568 (N_12568,N_12287,N_12141);
nor U12569 (N_12569,N_12233,N_12134);
nand U12570 (N_12570,N_12160,N_12478);
and U12571 (N_12571,N_12352,N_12353);
or U12572 (N_12572,N_12302,N_12081);
xnor U12573 (N_12573,N_12270,N_12142);
nor U12574 (N_12574,N_12061,N_12400);
and U12575 (N_12575,N_12218,N_12235);
nor U12576 (N_12576,N_12365,N_12363);
nand U12577 (N_12577,N_12320,N_12423);
xor U12578 (N_12578,N_12182,N_12442);
or U12579 (N_12579,N_12420,N_12216);
and U12580 (N_12580,N_12201,N_12307);
nor U12581 (N_12581,N_12021,N_12349);
nand U12582 (N_12582,N_12231,N_12185);
and U12583 (N_12583,N_12020,N_12055);
xnor U12584 (N_12584,N_12382,N_12136);
nor U12585 (N_12585,N_12040,N_12433);
nand U12586 (N_12586,N_12051,N_12441);
nand U12587 (N_12587,N_12007,N_12351);
xor U12588 (N_12588,N_12070,N_12153);
nor U12589 (N_12589,N_12425,N_12257);
xnor U12590 (N_12590,N_12319,N_12079);
nor U12591 (N_12591,N_12300,N_12445);
nor U12592 (N_12592,N_12226,N_12225);
xor U12593 (N_12593,N_12401,N_12151);
nor U12594 (N_12594,N_12198,N_12080);
and U12595 (N_12595,N_12095,N_12377);
nand U12596 (N_12596,N_12172,N_12143);
xnor U12597 (N_12597,N_12243,N_12106);
xor U12598 (N_12598,N_12175,N_12110);
or U12599 (N_12599,N_12176,N_12159);
or U12600 (N_12600,N_12317,N_12297);
nor U12601 (N_12601,N_12075,N_12117);
nand U12602 (N_12602,N_12260,N_12023);
or U12603 (N_12603,N_12304,N_12299);
xnor U12604 (N_12604,N_12165,N_12486);
and U12605 (N_12605,N_12440,N_12463);
nor U12606 (N_12606,N_12250,N_12221);
nand U12607 (N_12607,N_12375,N_12072);
or U12608 (N_12608,N_12336,N_12417);
nor U12609 (N_12609,N_12322,N_12157);
or U12610 (N_12610,N_12193,N_12097);
xor U12611 (N_12611,N_12408,N_12376);
nand U12612 (N_12612,N_12404,N_12126);
nand U12613 (N_12613,N_12379,N_12383);
nor U12614 (N_12614,N_12364,N_12224);
and U12615 (N_12615,N_12405,N_12476);
nor U12616 (N_12616,N_12140,N_12120);
or U12617 (N_12617,N_12449,N_12101);
and U12618 (N_12618,N_12448,N_12309);
or U12619 (N_12619,N_12356,N_12498);
xnor U12620 (N_12620,N_12118,N_12256);
or U12621 (N_12621,N_12239,N_12050);
or U12622 (N_12622,N_12398,N_12411);
xnor U12623 (N_12623,N_12306,N_12284);
or U12624 (N_12624,N_12388,N_12459);
xnor U12625 (N_12625,N_12152,N_12028);
nor U12626 (N_12626,N_12483,N_12206);
nand U12627 (N_12627,N_12105,N_12391);
nor U12628 (N_12628,N_12062,N_12456);
or U12629 (N_12629,N_12421,N_12036);
or U12630 (N_12630,N_12415,N_12063);
or U12631 (N_12631,N_12296,N_12026);
and U12632 (N_12632,N_12347,N_12035);
or U12633 (N_12633,N_12261,N_12373);
and U12634 (N_12634,N_12454,N_12479);
xor U12635 (N_12635,N_12455,N_12214);
nand U12636 (N_12636,N_12112,N_12450);
nand U12637 (N_12637,N_12278,N_12437);
or U12638 (N_12638,N_12313,N_12100);
or U12639 (N_12639,N_12043,N_12217);
and U12640 (N_12640,N_12409,N_12331);
nor U12641 (N_12641,N_12474,N_12237);
or U12642 (N_12642,N_12054,N_12279);
and U12643 (N_12643,N_12267,N_12446);
and U12644 (N_12644,N_12001,N_12203);
or U12645 (N_12645,N_12209,N_12457);
and U12646 (N_12646,N_12368,N_12076);
nand U12647 (N_12647,N_12181,N_12499);
and U12648 (N_12648,N_12234,N_12443);
and U12649 (N_12649,N_12330,N_12374);
nor U12650 (N_12650,N_12019,N_12164);
xor U12651 (N_12651,N_12362,N_12004);
and U12652 (N_12652,N_12066,N_12453);
nor U12653 (N_12653,N_12125,N_12108);
xor U12654 (N_12654,N_12163,N_12013);
nand U12655 (N_12655,N_12360,N_12434);
nand U12656 (N_12656,N_12266,N_12009);
and U12657 (N_12657,N_12311,N_12329);
nand U12658 (N_12658,N_12274,N_12088);
and U12659 (N_12659,N_12074,N_12018);
or U12660 (N_12660,N_12060,N_12166);
xor U12661 (N_12661,N_12240,N_12219);
or U12662 (N_12662,N_12008,N_12249);
xnor U12663 (N_12663,N_12242,N_12328);
nand U12664 (N_12664,N_12042,N_12099);
nor U12665 (N_12665,N_12215,N_12047);
nor U12666 (N_12666,N_12194,N_12428);
nand U12667 (N_12667,N_12029,N_12292);
and U12668 (N_12668,N_12122,N_12103);
or U12669 (N_12669,N_12452,N_12280);
and U12670 (N_12670,N_12124,N_12348);
and U12671 (N_12671,N_12487,N_12431);
and U12672 (N_12672,N_12016,N_12238);
nand U12673 (N_12673,N_12202,N_12424);
or U12674 (N_12674,N_12244,N_12094);
and U12675 (N_12675,N_12346,N_12109);
nand U12676 (N_12676,N_12410,N_12354);
nor U12677 (N_12677,N_12359,N_12380);
xnor U12678 (N_12678,N_12489,N_12162);
or U12679 (N_12679,N_12147,N_12068);
or U12680 (N_12680,N_12169,N_12044);
or U12681 (N_12681,N_12262,N_12482);
and U12682 (N_12682,N_12460,N_12156);
nand U12683 (N_12683,N_12495,N_12148);
or U12684 (N_12684,N_12387,N_12341);
nor U12685 (N_12685,N_12041,N_12293);
xnor U12686 (N_12686,N_12138,N_12015);
nor U12687 (N_12687,N_12343,N_12114);
nor U12688 (N_12688,N_12263,N_12012);
xor U12689 (N_12689,N_12332,N_12113);
nor U12690 (N_12690,N_12370,N_12305);
or U12691 (N_12691,N_12265,N_12092);
nor U12692 (N_12692,N_12291,N_12392);
and U12693 (N_12693,N_12048,N_12207);
nor U12694 (N_12694,N_12310,N_12340);
nor U12695 (N_12695,N_12116,N_12395);
or U12696 (N_12696,N_12057,N_12197);
nor U12697 (N_12697,N_12381,N_12259);
or U12698 (N_12698,N_12131,N_12034);
xor U12699 (N_12699,N_12073,N_12472);
and U12700 (N_12700,N_12462,N_12223);
or U12701 (N_12701,N_12083,N_12085);
xnor U12702 (N_12702,N_12390,N_12188);
nand U12703 (N_12703,N_12422,N_12496);
nor U12704 (N_12704,N_12294,N_12093);
or U12705 (N_12705,N_12130,N_12286);
nand U12706 (N_12706,N_12481,N_12484);
or U12707 (N_12707,N_12465,N_12355);
nor U12708 (N_12708,N_12334,N_12132);
xor U12709 (N_12709,N_12022,N_12407);
and U12710 (N_12710,N_12006,N_12477);
or U12711 (N_12711,N_12494,N_12230);
nor U12712 (N_12712,N_12078,N_12493);
and U12713 (N_12713,N_12191,N_12146);
xnor U12714 (N_12714,N_12177,N_12324);
nand U12715 (N_12715,N_12295,N_12046);
nor U12716 (N_12716,N_12205,N_12326);
nor U12717 (N_12717,N_12241,N_12123);
nand U12718 (N_12718,N_12096,N_12167);
xor U12719 (N_12719,N_12228,N_12414);
xor U12720 (N_12720,N_12491,N_12010);
xor U12721 (N_12721,N_12308,N_12212);
and U12722 (N_12722,N_12104,N_12385);
nand U12723 (N_12723,N_12253,N_12342);
xor U12724 (N_12724,N_12213,N_12174);
nor U12725 (N_12725,N_12171,N_12077);
xnor U12726 (N_12726,N_12316,N_12333);
and U12727 (N_12727,N_12497,N_12086);
or U12728 (N_12728,N_12189,N_12069);
xnor U12729 (N_12729,N_12488,N_12338);
xor U12730 (N_12730,N_12192,N_12367);
or U12731 (N_12731,N_12490,N_12475);
or U12732 (N_12732,N_12366,N_12145);
nor U12733 (N_12733,N_12458,N_12033);
xor U12734 (N_12734,N_12403,N_12204);
nor U12735 (N_12735,N_12429,N_12461);
and U12736 (N_12736,N_12045,N_12133);
and U12737 (N_12737,N_12102,N_12372);
nand U12738 (N_12738,N_12056,N_12111);
or U12739 (N_12739,N_12303,N_12480);
and U12740 (N_12740,N_12436,N_12397);
nand U12741 (N_12741,N_12357,N_12210);
and U12742 (N_12742,N_12027,N_12252);
xor U12743 (N_12743,N_12154,N_12024);
or U12744 (N_12744,N_12285,N_12014);
nand U12745 (N_12745,N_12149,N_12430);
nand U12746 (N_12746,N_12399,N_12323);
nand U12747 (N_12747,N_12229,N_12137);
nand U12748 (N_12748,N_12419,N_12466);
xnor U12749 (N_12749,N_12158,N_12389);
and U12750 (N_12750,N_12403,N_12244);
or U12751 (N_12751,N_12083,N_12330);
or U12752 (N_12752,N_12322,N_12235);
nor U12753 (N_12753,N_12216,N_12138);
nor U12754 (N_12754,N_12258,N_12011);
nor U12755 (N_12755,N_12004,N_12379);
nor U12756 (N_12756,N_12177,N_12329);
or U12757 (N_12757,N_12277,N_12335);
xor U12758 (N_12758,N_12228,N_12070);
xnor U12759 (N_12759,N_12179,N_12471);
nand U12760 (N_12760,N_12295,N_12326);
nand U12761 (N_12761,N_12069,N_12090);
nor U12762 (N_12762,N_12485,N_12173);
and U12763 (N_12763,N_12492,N_12105);
nand U12764 (N_12764,N_12320,N_12483);
nor U12765 (N_12765,N_12480,N_12144);
nor U12766 (N_12766,N_12141,N_12481);
nor U12767 (N_12767,N_12179,N_12142);
and U12768 (N_12768,N_12117,N_12378);
xor U12769 (N_12769,N_12183,N_12251);
xor U12770 (N_12770,N_12499,N_12461);
and U12771 (N_12771,N_12150,N_12157);
nand U12772 (N_12772,N_12185,N_12046);
xnor U12773 (N_12773,N_12286,N_12294);
and U12774 (N_12774,N_12006,N_12300);
nor U12775 (N_12775,N_12374,N_12059);
or U12776 (N_12776,N_12471,N_12239);
nor U12777 (N_12777,N_12401,N_12044);
xnor U12778 (N_12778,N_12286,N_12278);
and U12779 (N_12779,N_12234,N_12046);
nor U12780 (N_12780,N_12092,N_12391);
nand U12781 (N_12781,N_12104,N_12204);
xnor U12782 (N_12782,N_12096,N_12168);
nand U12783 (N_12783,N_12112,N_12040);
xnor U12784 (N_12784,N_12225,N_12114);
or U12785 (N_12785,N_12387,N_12323);
or U12786 (N_12786,N_12173,N_12151);
or U12787 (N_12787,N_12398,N_12187);
xnor U12788 (N_12788,N_12234,N_12131);
xor U12789 (N_12789,N_12240,N_12078);
xor U12790 (N_12790,N_12192,N_12394);
nor U12791 (N_12791,N_12064,N_12120);
or U12792 (N_12792,N_12183,N_12296);
and U12793 (N_12793,N_12076,N_12297);
or U12794 (N_12794,N_12208,N_12050);
or U12795 (N_12795,N_12014,N_12442);
and U12796 (N_12796,N_12019,N_12468);
nor U12797 (N_12797,N_12424,N_12069);
nand U12798 (N_12798,N_12365,N_12161);
nand U12799 (N_12799,N_12492,N_12030);
and U12800 (N_12800,N_12403,N_12367);
xor U12801 (N_12801,N_12182,N_12414);
nor U12802 (N_12802,N_12451,N_12229);
nor U12803 (N_12803,N_12495,N_12087);
nand U12804 (N_12804,N_12029,N_12422);
and U12805 (N_12805,N_12300,N_12007);
or U12806 (N_12806,N_12405,N_12288);
nor U12807 (N_12807,N_12349,N_12298);
nor U12808 (N_12808,N_12324,N_12181);
nand U12809 (N_12809,N_12293,N_12007);
or U12810 (N_12810,N_12345,N_12484);
and U12811 (N_12811,N_12070,N_12069);
nor U12812 (N_12812,N_12498,N_12303);
xnor U12813 (N_12813,N_12033,N_12217);
xnor U12814 (N_12814,N_12218,N_12184);
nor U12815 (N_12815,N_12031,N_12258);
and U12816 (N_12816,N_12342,N_12169);
nand U12817 (N_12817,N_12004,N_12048);
or U12818 (N_12818,N_12316,N_12075);
or U12819 (N_12819,N_12224,N_12324);
nor U12820 (N_12820,N_12208,N_12023);
or U12821 (N_12821,N_12123,N_12292);
nand U12822 (N_12822,N_12143,N_12375);
nor U12823 (N_12823,N_12390,N_12122);
xor U12824 (N_12824,N_12377,N_12375);
nor U12825 (N_12825,N_12435,N_12297);
or U12826 (N_12826,N_12106,N_12198);
nand U12827 (N_12827,N_12491,N_12433);
or U12828 (N_12828,N_12414,N_12037);
and U12829 (N_12829,N_12336,N_12326);
nor U12830 (N_12830,N_12457,N_12033);
xnor U12831 (N_12831,N_12465,N_12360);
nand U12832 (N_12832,N_12071,N_12161);
or U12833 (N_12833,N_12212,N_12332);
nor U12834 (N_12834,N_12340,N_12116);
or U12835 (N_12835,N_12315,N_12114);
xor U12836 (N_12836,N_12471,N_12150);
or U12837 (N_12837,N_12073,N_12140);
nand U12838 (N_12838,N_12149,N_12337);
nor U12839 (N_12839,N_12218,N_12329);
and U12840 (N_12840,N_12186,N_12333);
and U12841 (N_12841,N_12216,N_12295);
nand U12842 (N_12842,N_12215,N_12141);
nor U12843 (N_12843,N_12068,N_12432);
xor U12844 (N_12844,N_12408,N_12045);
nand U12845 (N_12845,N_12499,N_12028);
nand U12846 (N_12846,N_12268,N_12004);
nand U12847 (N_12847,N_12359,N_12450);
nor U12848 (N_12848,N_12172,N_12348);
nor U12849 (N_12849,N_12461,N_12276);
and U12850 (N_12850,N_12131,N_12143);
and U12851 (N_12851,N_12467,N_12353);
xor U12852 (N_12852,N_12029,N_12304);
or U12853 (N_12853,N_12127,N_12068);
and U12854 (N_12854,N_12274,N_12256);
nor U12855 (N_12855,N_12174,N_12128);
xor U12856 (N_12856,N_12429,N_12423);
nor U12857 (N_12857,N_12489,N_12016);
and U12858 (N_12858,N_12305,N_12055);
xor U12859 (N_12859,N_12225,N_12190);
and U12860 (N_12860,N_12078,N_12417);
xor U12861 (N_12861,N_12252,N_12359);
and U12862 (N_12862,N_12079,N_12265);
xnor U12863 (N_12863,N_12129,N_12184);
or U12864 (N_12864,N_12321,N_12337);
nor U12865 (N_12865,N_12226,N_12268);
and U12866 (N_12866,N_12176,N_12332);
or U12867 (N_12867,N_12342,N_12194);
or U12868 (N_12868,N_12116,N_12109);
xnor U12869 (N_12869,N_12269,N_12005);
and U12870 (N_12870,N_12094,N_12253);
or U12871 (N_12871,N_12117,N_12485);
and U12872 (N_12872,N_12226,N_12287);
nand U12873 (N_12873,N_12144,N_12449);
nor U12874 (N_12874,N_12280,N_12040);
or U12875 (N_12875,N_12423,N_12127);
nand U12876 (N_12876,N_12473,N_12469);
and U12877 (N_12877,N_12171,N_12001);
or U12878 (N_12878,N_12159,N_12042);
xor U12879 (N_12879,N_12219,N_12407);
xnor U12880 (N_12880,N_12473,N_12065);
and U12881 (N_12881,N_12079,N_12029);
nor U12882 (N_12882,N_12358,N_12471);
xor U12883 (N_12883,N_12435,N_12128);
xor U12884 (N_12884,N_12456,N_12267);
nand U12885 (N_12885,N_12054,N_12394);
nand U12886 (N_12886,N_12258,N_12105);
or U12887 (N_12887,N_12156,N_12223);
and U12888 (N_12888,N_12301,N_12097);
or U12889 (N_12889,N_12434,N_12039);
nand U12890 (N_12890,N_12097,N_12285);
xor U12891 (N_12891,N_12278,N_12465);
nor U12892 (N_12892,N_12479,N_12039);
nand U12893 (N_12893,N_12113,N_12282);
nor U12894 (N_12894,N_12451,N_12165);
and U12895 (N_12895,N_12043,N_12301);
nor U12896 (N_12896,N_12286,N_12381);
nand U12897 (N_12897,N_12218,N_12125);
or U12898 (N_12898,N_12053,N_12072);
and U12899 (N_12899,N_12032,N_12104);
or U12900 (N_12900,N_12202,N_12099);
and U12901 (N_12901,N_12081,N_12146);
or U12902 (N_12902,N_12026,N_12042);
xnor U12903 (N_12903,N_12458,N_12280);
nand U12904 (N_12904,N_12016,N_12069);
nor U12905 (N_12905,N_12050,N_12491);
and U12906 (N_12906,N_12309,N_12273);
or U12907 (N_12907,N_12456,N_12219);
nand U12908 (N_12908,N_12337,N_12246);
and U12909 (N_12909,N_12116,N_12029);
xor U12910 (N_12910,N_12041,N_12196);
and U12911 (N_12911,N_12047,N_12360);
nand U12912 (N_12912,N_12279,N_12378);
or U12913 (N_12913,N_12189,N_12044);
nand U12914 (N_12914,N_12163,N_12335);
xor U12915 (N_12915,N_12092,N_12001);
or U12916 (N_12916,N_12030,N_12136);
nand U12917 (N_12917,N_12399,N_12366);
nand U12918 (N_12918,N_12288,N_12120);
nor U12919 (N_12919,N_12130,N_12195);
and U12920 (N_12920,N_12406,N_12495);
nand U12921 (N_12921,N_12445,N_12029);
xnor U12922 (N_12922,N_12439,N_12333);
nor U12923 (N_12923,N_12412,N_12240);
nor U12924 (N_12924,N_12077,N_12268);
or U12925 (N_12925,N_12034,N_12161);
xnor U12926 (N_12926,N_12095,N_12198);
xnor U12927 (N_12927,N_12256,N_12257);
xor U12928 (N_12928,N_12404,N_12484);
or U12929 (N_12929,N_12137,N_12425);
or U12930 (N_12930,N_12037,N_12067);
nand U12931 (N_12931,N_12416,N_12468);
nor U12932 (N_12932,N_12067,N_12493);
and U12933 (N_12933,N_12373,N_12198);
xnor U12934 (N_12934,N_12261,N_12394);
xnor U12935 (N_12935,N_12143,N_12325);
or U12936 (N_12936,N_12088,N_12050);
nand U12937 (N_12937,N_12028,N_12493);
nand U12938 (N_12938,N_12088,N_12323);
nand U12939 (N_12939,N_12049,N_12246);
and U12940 (N_12940,N_12289,N_12382);
nor U12941 (N_12941,N_12450,N_12019);
and U12942 (N_12942,N_12347,N_12245);
nand U12943 (N_12943,N_12126,N_12295);
xnor U12944 (N_12944,N_12362,N_12340);
xor U12945 (N_12945,N_12257,N_12176);
nand U12946 (N_12946,N_12121,N_12498);
xnor U12947 (N_12947,N_12133,N_12069);
nor U12948 (N_12948,N_12331,N_12121);
nand U12949 (N_12949,N_12140,N_12006);
or U12950 (N_12950,N_12303,N_12164);
nor U12951 (N_12951,N_12260,N_12300);
and U12952 (N_12952,N_12457,N_12150);
xor U12953 (N_12953,N_12151,N_12403);
nand U12954 (N_12954,N_12239,N_12266);
nor U12955 (N_12955,N_12220,N_12080);
nand U12956 (N_12956,N_12103,N_12496);
nand U12957 (N_12957,N_12013,N_12280);
nor U12958 (N_12958,N_12466,N_12037);
nand U12959 (N_12959,N_12161,N_12355);
nor U12960 (N_12960,N_12174,N_12460);
and U12961 (N_12961,N_12339,N_12225);
nor U12962 (N_12962,N_12107,N_12306);
nor U12963 (N_12963,N_12179,N_12192);
nor U12964 (N_12964,N_12451,N_12463);
or U12965 (N_12965,N_12248,N_12336);
or U12966 (N_12966,N_12273,N_12170);
nand U12967 (N_12967,N_12245,N_12387);
nand U12968 (N_12968,N_12487,N_12078);
or U12969 (N_12969,N_12062,N_12029);
or U12970 (N_12970,N_12243,N_12221);
and U12971 (N_12971,N_12109,N_12391);
and U12972 (N_12972,N_12234,N_12486);
nand U12973 (N_12973,N_12334,N_12029);
nand U12974 (N_12974,N_12043,N_12408);
and U12975 (N_12975,N_12148,N_12439);
and U12976 (N_12976,N_12024,N_12240);
and U12977 (N_12977,N_12226,N_12492);
and U12978 (N_12978,N_12418,N_12318);
nand U12979 (N_12979,N_12433,N_12099);
and U12980 (N_12980,N_12495,N_12031);
xnor U12981 (N_12981,N_12065,N_12208);
nor U12982 (N_12982,N_12162,N_12211);
or U12983 (N_12983,N_12441,N_12139);
nand U12984 (N_12984,N_12344,N_12078);
and U12985 (N_12985,N_12344,N_12452);
and U12986 (N_12986,N_12141,N_12127);
xnor U12987 (N_12987,N_12141,N_12193);
and U12988 (N_12988,N_12412,N_12094);
xor U12989 (N_12989,N_12221,N_12331);
nand U12990 (N_12990,N_12496,N_12143);
nor U12991 (N_12991,N_12310,N_12164);
nand U12992 (N_12992,N_12300,N_12167);
nor U12993 (N_12993,N_12187,N_12292);
nor U12994 (N_12994,N_12192,N_12312);
nor U12995 (N_12995,N_12222,N_12098);
or U12996 (N_12996,N_12496,N_12276);
xor U12997 (N_12997,N_12122,N_12378);
or U12998 (N_12998,N_12327,N_12251);
xor U12999 (N_12999,N_12149,N_12194);
nor U13000 (N_13000,N_12632,N_12710);
nor U13001 (N_13001,N_12860,N_12976);
or U13002 (N_13002,N_12914,N_12761);
xnor U13003 (N_13003,N_12576,N_12959);
nor U13004 (N_13004,N_12921,N_12788);
nor U13005 (N_13005,N_12563,N_12748);
or U13006 (N_13006,N_12801,N_12852);
or U13007 (N_13007,N_12782,N_12695);
or U13008 (N_13008,N_12538,N_12677);
or U13009 (N_13009,N_12739,N_12835);
and U13010 (N_13010,N_12689,N_12787);
xor U13011 (N_13011,N_12947,N_12807);
nand U13012 (N_13012,N_12719,N_12679);
or U13013 (N_13013,N_12631,N_12968);
or U13014 (N_13014,N_12507,N_12777);
nor U13015 (N_13015,N_12556,N_12714);
nand U13016 (N_13016,N_12757,N_12519);
xor U13017 (N_13017,N_12655,N_12809);
nor U13018 (N_13018,N_12609,N_12585);
xor U13019 (N_13019,N_12523,N_12876);
nor U13020 (N_13020,N_12767,N_12928);
nand U13021 (N_13021,N_12681,N_12682);
and U13022 (N_13022,N_12615,N_12721);
nor U13023 (N_13023,N_12736,N_12918);
xor U13024 (N_13024,N_12709,N_12793);
nand U13025 (N_13025,N_12636,N_12840);
nand U13026 (N_13026,N_12561,N_12865);
and U13027 (N_13027,N_12587,N_12594);
nor U13028 (N_13028,N_12597,N_12554);
xor U13029 (N_13029,N_12885,N_12588);
xor U13030 (N_13030,N_12954,N_12572);
or U13031 (N_13031,N_12846,N_12937);
nor U13032 (N_13032,N_12766,N_12528);
xnor U13033 (N_13033,N_12649,N_12798);
or U13034 (N_13034,N_12532,N_12771);
nor U13035 (N_13035,N_12505,N_12931);
nand U13036 (N_13036,N_12905,N_12794);
nor U13037 (N_13037,N_12863,N_12772);
nand U13038 (N_13038,N_12715,N_12819);
nor U13039 (N_13039,N_12664,N_12527);
and U13040 (N_13040,N_12596,N_12702);
xor U13041 (N_13041,N_12734,N_12502);
nor U13042 (N_13042,N_12984,N_12708);
or U13043 (N_13043,N_12616,N_12866);
xor U13044 (N_13044,N_12637,N_12839);
and U13045 (N_13045,N_12907,N_12613);
and U13046 (N_13046,N_12699,N_12762);
nor U13047 (N_13047,N_12768,N_12864);
nor U13048 (N_13048,N_12514,N_12555);
and U13049 (N_13049,N_12672,N_12660);
nand U13050 (N_13050,N_12844,N_12881);
nand U13051 (N_13051,N_12601,N_12706);
and U13052 (N_13052,N_12756,N_12849);
or U13053 (N_13053,N_12818,N_12848);
nand U13054 (N_13054,N_12593,N_12758);
and U13055 (N_13055,N_12770,N_12912);
nand U13056 (N_13056,N_12573,N_12648);
nand U13057 (N_13057,N_12871,N_12557);
xnor U13058 (N_13058,N_12967,N_12598);
and U13059 (N_13059,N_12898,N_12744);
nor U13060 (N_13060,N_12753,N_12607);
nand U13061 (N_13061,N_12583,N_12738);
nand U13062 (N_13062,N_12579,N_12539);
xnor U13063 (N_13063,N_12675,N_12624);
or U13064 (N_13064,N_12558,N_12717);
nor U13065 (N_13065,N_12570,N_12812);
xnor U13066 (N_13066,N_12994,N_12985);
and U13067 (N_13067,N_12800,N_12590);
and U13068 (N_13068,N_12535,N_12831);
xnor U13069 (N_13069,N_12680,N_12843);
nor U13070 (N_13070,N_12541,N_12902);
nand U13071 (N_13071,N_12763,N_12741);
nor U13072 (N_13072,N_12640,N_12617);
nor U13073 (N_13073,N_12652,N_12900);
or U13074 (N_13074,N_12608,N_12773);
xor U13075 (N_13075,N_12740,N_12981);
nor U13076 (N_13076,N_12603,N_12989);
or U13077 (N_13077,N_12543,N_12893);
nand U13078 (N_13078,N_12999,N_12656);
and U13079 (N_13079,N_12635,N_12899);
xnor U13080 (N_13080,N_12694,N_12990);
or U13081 (N_13081,N_12678,N_12837);
nor U13082 (N_13082,N_12829,N_12906);
nor U13083 (N_13083,N_12992,N_12980);
nor U13084 (N_13084,N_12877,N_12669);
xnor U13085 (N_13085,N_12910,N_12786);
and U13086 (N_13086,N_12641,N_12929);
and U13087 (N_13087,N_12661,N_12857);
and U13088 (N_13088,N_12537,N_12913);
xor U13089 (N_13089,N_12972,N_12611);
xnor U13090 (N_13090,N_12964,N_12803);
and U13091 (N_13091,N_12759,N_12657);
nor U13092 (N_13092,N_12911,N_12614);
xor U13093 (N_13093,N_12956,N_12546);
or U13094 (N_13094,N_12855,N_12925);
nor U13095 (N_13095,N_12955,N_12935);
xor U13096 (N_13096,N_12540,N_12693);
nand U13097 (N_13097,N_12700,N_12804);
nand U13098 (N_13098,N_12671,N_12960);
xor U13099 (N_13099,N_12799,N_12854);
or U13100 (N_13100,N_12979,N_12834);
xnor U13101 (N_13101,N_12703,N_12904);
nor U13102 (N_13102,N_12534,N_12723);
and U13103 (N_13103,N_12692,N_12567);
xnor U13104 (N_13104,N_12683,N_12595);
nand U13105 (N_13105,N_12847,N_12524);
or U13106 (N_13106,N_12936,N_12975);
xor U13107 (N_13107,N_12665,N_12642);
and U13108 (N_13108,N_12584,N_12821);
or U13109 (N_13109,N_12784,N_12944);
nor U13110 (N_13110,N_12684,N_12581);
or U13111 (N_13111,N_12605,N_12512);
and U13112 (N_13112,N_12606,N_12765);
or U13113 (N_13113,N_12932,N_12789);
nand U13114 (N_13114,N_12988,N_12745);
and U13115 (N_13115,N_12589,N_12806);
and U13116 (N_13116,N_12506,N_12903);
xor U13117 (N_13117,N_12653,N_12971);
xnor U13118 (N_13118,N_12752,N_12500);
nor U13119 (N_13119,N_12861,N_12574);
xnor U13120 (N_13120,N_12737,N_12895);
and U13121 (N_13121,N_12577,N_12892);
nand U13122 (N_13122,N_12965,N_12628);
or U13123 (N_13123,N_12663,N_12850);
and U13124 (N_13124,N_12630,N_12888);
or U13125 (N_13125,N_12633,N_12897);
nand U13126 (N_13126,N_12549,N_12511);
xor U13127 (N_13127,N_12610,N_12529);
nand U13128 (N_13128,N_12559,N_12544);
xor U13129 (N_13129,N_12645,N_12517);
and U13130 (N_13130,N_12670,N_12949);
nor U13131 (N_13131,N_12668,N_12817);
nor U13132 (N_13132,N_12824,N_12940);
nor U13133 (N_13133,N_12580,N_12868);
and U13134 (N_13134,N_12676,N_12845);
xnor U13135 (N_13135,N_12566,N_12531);
nor U13136 (N_13136,N_12711,N_12571);
nand U13137 (N_13137,N_12720,N_12697);
nand U13138 (N_13138,N_12815,N_12504);
and U13139 (N_13139,N_12982,N_12909);
and U13140 (N_13140,N_12878,N_12934);
xor U13141 (N_13141,N_12733,N_12930);
nand U13142 (N_13142,N_12802,N_12643);
or U13143 (N_13143,N_12945,N_12578);
and U13144 (N_13144,N_12942,N_12569);
nand U13145 (N_13145,N_12521,N_12662);
nand U13146 (N_13146,N_12747,N_12833);
nand U13147 (N_13147,N_12810,N_12729);
and U13148 (N_13148,N_12701,N_12751);
xor U13149 (N_13149,N_12634,N_12749);
and U13150 (N_13150,N_12627,N_12939);
or U13151 (N_13151,N_12779,N_12969);
nand U13152 (N_13152,N_12639,N_12966);
nor U13153 (N_13153,N_12755,N_12704);
or U13154 (N_13154,N_12508,N_12530);
nor U13155 (N_13155,N_12862,N_12908);
nor U13156 (N_13156,N_12974,N_12823);
xor U13157 (N_13157,N_12725,N_12983);
xor U13158 (N_13158,N_12896,N_12644);
and U13159 (N_13159,N_12783,N_12727);
nor U13160 (N_13160,N_12948,N_12775);
xnor U13161 (N_13161,N_12933,N_12894);
xor U13162 (N_13162,N_12814,N_12873);
nand U13163 (N_13163,N_12619,N_12686);
nor U13164 (N_13164,N_12638,N_12551);
and U13165 (N_13165,N_12575,N_12826);
and U13166 (N_13166,N_12875,N_12732);
and U13167 (N_13167,N_12998,N_12986);
nor U13168 (N_13168,N_12722,N_12991);
nand U13169 (N_13169,N_12997,N_12618);
nor U13170 (N_13170,N_12816,N_12522);
or U13171 (N_13171,N_12957,N_12962);
xor U13172 (N_13172,N_12769,N_12625);
xnor U13173 (N_13173,N_12901,N_12586);
nor U13174 (N_13174,N_12730,N_12889);
nor U13175 (N_13175,N_12778,N_12890);
or U13176 (N_13176,N_12958,N_12518);
nand U13177 (N_13177,N_12688,N_12869);
and U13178 (N_13178,N_12716,N_12724);
nand U13179 (N_13179,N_12516,N_12674);
xnor U13180 (N_13180,N_12510,N_12883);
nor U13181 (N_13181,N_12827,N_12764);
nand U13182 (N_13182,N_12743,N_12841);
xnor U13183 (N_13183,N_12728,N_12951);
or U13184 (N_13184,N_12791,N_12503);
nand U13185 (N_13185,N_12880,N_12659);
and U13186 (N_13186,N_12884,N_12582);
xor U13187 (N_13187,N_12562,N_12667);
nand U13188 (N_13188,N_12978,N_12602);
xor U13189 (N_13189,N_12629,N_12795);
or U13190 (N_13190,N_12856,N_12828);
nor U13191 (N_13191,N_12977,N_12654);
nand U13192 (N_13192,N_12533,N_12851);
nand U13193 (N_13193,N_12926,N_12525);
and U13194 (N_13194,N_12970,N_12760);
and U13195 (N_13195,N_12646,N_12565);
and U13196 (N_13196,N_12825,N_12647);
nand U13197 (N_13197,N_12797,N_12886);
xor U13198 (N_13198,N_12993,N_12754);
and U13199 (N_13199,N_12600,N_12650);
and U13200 (N_13200,N_12927,N_12950);
nor U13201 (N_13201,N_12790,N_12938);
xnor U13202 (N_13202,N_12859,N_12995);
nand U13203 (N_13203,N_12891,N_12685);
or U13204 (N_13204,N_12526,N_12917);
nand U13205 (N_13205,N_12776,N_12987);
or U13206 (N_13206,N_12658,N_12879);
nand U13207 (N_13207,N_12696,N_12592);
xor U13208 (N_13208,N_12698,N_12515);
nor U13209 (N_13209,N_12712,N_12996);
or U13210 (N_13210,N_12564,N_12780);
or U13211 (N_13211,N_12853,N_12626);
or U13212 (N_13212,N_12520,N_12501);
nand U13213 (N_13213,N_12742,N_12805);
nor U13214 (N_13214,N_12735,N_12872);
nand U13215 (N_13215,N_12820,N_12621);
nor U13216 (N_13216,N_12811,N_12666);
xnor U13217 (N_13217,N_12553,N_12604);
nand U13218 (N_13218,N_12545,N_12838);
or U13219 (N_13219,N_12882,N_12963);
and U13220 (N_13220,N_12513,N_12915);
nor U13221 (N_13221,N_12691,N_12796);
nor U13222 (N_13222,N_12785,N_12750);
nor U13223 (N_13223,N_12687,N_12705);
xnor U13224 (N_13224,N_12746,N_12874);
or U13225 (N_13225,N_12887,N_12924);
nor U13226 (N_13226,N_12690,N_12953);
or U13227 (N_13227,N_12622,N_12612);
and U13228 (N_13228,N_12870,N_12599);
or U13229 (N_13229,N_12973,N_12836);
xor U13230 (N_13230,N_12920,N_12916);
or U13231 (N_13231,N_12832,N_12792);
xnor U13232 (N_13232,N_12552,N_12673);
xor U13233 (N_13233,N_12591,N_12707);
xnor U13234 (N_13234,N_12943,N_12731);
nor U13235 (N_13235,N_12542,N_12813);
or U13236 (N_13236,N_12923,N_12774);
nand U13237 (N_13237,N_12548,N_12961);
nor U13238 (N_13238,N_12858,N_12808);
nor U13239 (N_13239,N_12946,N_12919);
nand U13240 (N_13240,N_12536,N_12842);
nand U13241 (N_13241,N_12781,N_12822);
xnor U13242 (N_13242,N_12651,N_12941);
and U13243 (N_13243,N_12550,N_12623);
nand U13244 (N_13244,N_12726,N_12867);
xnor U13245 (N_13245,N_12718,N_12560);
nand U13246 (N_13246,N_12713,N_12547);
and U13247 (N_13247,N_12620,N_12922);
xnor U13248 (N_13248,N_12509,N_12830);
nand U13249 (N_13249,N_12952,N_12568);
nand U13250 (N_13250,N_12874,N_12693);
nor U13251 (N_13251,N_12515,N_12531);
and U13252 (N_13252,N_12724,N_12838);
nor U13253 (N_13253,N_12784,N_12733);
nor U13254 (N_13254,N_12706,N_12593);
or U13255 (N_13255,N_12955,N_12590);
or U13256 (N_13256,N_12564,N_12976);
nand U13257 (N_13257,N_12611,N_12737);
and U13258 (N_13258,N_12681,N_12740);
nand U13259 (N_13259,N_12859,N_12711);
xnor U13260 (N_13260,N_12855,N_12710);
nor U13261 (N_13261,N_12836,N_12948);
and U13262 (N_13262,N_12911,N_12615);
or U13263 (N_13263,N_12875,N_12669);
or U13264 (N_13264,N_12871,N_12500);
xnor U13265 (N_13265,N_12790,N_12640);
nand U13266 (N_13266,N_12707,N_12901);
or U13267 (N_13267,N_12833,N_12745);
nand U13268 (N_13268,N_12528,N_12954);
nor U13269 (N_13269,N_12858,N_12756);
xor U13270 (N_13270,N_12981,N_12758);
nand U13271 (N_13271,N_12507,N_12648);
and U13272 (N_13272,N_12732,N_12519);
xor U13273 (N_13273,N_12627,N_12538);
and U13274 (N_13274,N_12907,N_12834);
nor U13275 (N_13275,N_12952,N_12723);
nor U13276 (N_13276,N_12938,N_12519);
and U13277 (N_13277,N_12527,N_12736);
nor U13278 (N_13278,N_12667,N_12617);
nand U13279 (N_13279,N_12594,N_12931);
nand U13280 (N_13280,N_12965,N_12940);
nand U13281 (N_13281,N_12659,N_12913);
nor U13282 (N_13282,N_12560,N_12970);
or U13283 (N_13283,N_12668,N_12687);
and U13284 (N_13284,N_12828,N_12936);
or U13285 (N_13285,N_12747,N_12756);
and U13286 (N_13286,N_12775,N_12629);
or U13287 (N_13287,N_12758,N_12654);
and U13288 (N_13288,N_12960,N_12781);
or U13289 (N_13289,N_12987,N_12851);
nor U13290 (N_13290,N_12936,N_12883);
nand U13291 (N_13291,N_12519,N_12849);
xor U13292 (N_13292,N_12601,N_12741);
nor U13293 (N_13293,N_12732,N_12651);
nand U13294 (N_13294,N_12712,N_12624);
nor U13295 (N_13295,N_12619,N_12819);
nor U13296 (N_13296,N_12728,N_12583);
nor U13297 (N_13297,N_12851,N_12813);
xor U13298 (N_13298,N_12821,N_12870);
nand U13299 (N_13299,N_12754,N_12762);
nand U13300 (N_13300,N_12723,N_12684);
nor U13301 (N_13301,N_12511,N_12877);
or U13302 (N_13302,N_12625,N_12605);
nor U13303 (N_13303,N_12862,N_12696);
nor U13304 (N_13304,N_12936,N_12983);
and U13305 (N_13305,N_12898,N_12847);
nor U13306 (N_13306,N_12841,N_12733);
nand U13307 (N_13307,N_12787,N_12588);
xor U13308 (N_13308,N_12927,N_12549);
nand U13309 (N_13309,N_12743,N_12785);
nor U13310 (N_13310,N_12600,N_12950);
nor U13311 (N_13311,N_12686,N_12740);
xnor U13312 (N_13312,N_12994,N_12820);
and U13313 (N_13313,N_12643,N_12634);
nand U13314 (N_13314,N_12917,N_12811);
xor U13315 (N_13315,N_12955,N_12554);
or U13316 (N_13316,N_12840,N_12868);
and U13317 (N_13317,N_12518,N_12936);
nor U13318 (N_13318,N_12943,N_12855);
nor U13319 (N_13319,N_12838,N_12827);
nor U13320 (N_13320,N_12568,N_12919);
nor U13321 (N_13321,N_12892,N_12868);
xor U13322 (N_13322,N_12893,N_12968);
nor U13323 (N_13323,N_12943,N_12770);
nor U13324 (N_13324,N_12618,N_12501);
nor U13325 (N_13325,N_12551,N_12907);
nand U13326 (N_13326,N_12967,N_12526);
nor U13327 (N_13327,N_12899,N_12508);
xnor U13328 (N_13328,N_12652,N_12843);
or U13329 (N_13329,N_12966,N_12517);
xor U13330 (N_13330,N_12660,N_12597);
or U13331 (N_13331,N_12916,N_12610);
nor U13332 (N_13332,N_12924,N_12801);
or U13333 (N_13333,N_12751,N_12998);
xor U13334 (N_13334,N_12948,N_12574);
nor U13335 (N_13335,N_12816,N_12620);
and U13336 (N_13336,N_12821,N_12970);
or U13337 (N_13337,N_12896,N_12826);
or U13338 (N_13338,N_12570,N_12979);
nor U13339 (N_13339,N_12926,N_12855);
nor U13340 (N_13340,N_12638,N_12904);
xnor U13341 (N_13341,N_12550,N_12996);
nor U13342 (N_13342,N_12676,N_12907);
xnor U13343 (N_13343,N_12895,N_12576);
nor U13344 (N_13344,N_12813,N_12707);
nand U13345 (N_13345,N_12818,N_12840);
nor U13346 (N_13346,N_12582,N_12777);
xnor U13347 (N_13347,N_12958,N_12778);
xor U13348 (N_13348,N_12752,N_12755);
nand U13349 (N_13349,N_12937,N_12665);
xor U13350 (N_13350,N_12560,N_12726);
or U13351 (N_13351,N_12928,N_12722);
or U13352 (N_13352,N_12519,N_12552);
nand U13353 (N_13353,N_12991,N_12900);
nand U13354 (N_13354,N_12749,N_12941);
nand U13355 (N_13355,N_12795,N_12737);
xnor U13356 (N_13356,N_12608,N_12690);
xnor U13357 (N_13357,N_12688,N_12661);
xor U13358 (N_13358,N_12558,N_12851);
and U13359 (N_13359,N_12739,N_12539);
or U13360 (N_13360,N_12788,N_12684);
and U13361 (N_13361,N_12725,N_12756);
nor U13362 (N_13362,N_12980,N_12815);
and U13363 (N_13363,N_12743,N_12548);
nor U13364 (N_13364,N_12942,N_12580);
nand U13365 (N_13365,N_12916,N_12712);
or U13366 (N_13366,N_12612,N_12752);
nand U13367 (N_13367,N_12841,N_12719);
nand U13368 (N_13368,N_12780,N_12654);
nand U13369 (N_13369,N_12676,N_12685);
or U13370 (N_13370,N_12591,N_12931);
or U13371 (N_13371,N_12531,N_12780);
xor U13372 (N_13372,N_12705,N_12545);
nor U13373 (N_13373,N_12950,N_12548);
or U13374 (N_13374,N_12847,N_12605);
nor U13375 (N_13375,N_12714,N_12599);
nand U13376 (N_13376,N_12945,N_12959);
nor U13377 (N_13377,N_12524,N_12756);
xnor U13378 (N_13378,N_12545,N_12845);
nand U13379 (N_13379,N_12906,N_12816);
nand U13380 (N_13380,N_12741,N_12607);
or U13381 (N_13381,N_12886,N_12829);
nor U13382 (N_13382,N_12520,N_12907);
nor U13383 (N_13383,N_12850,N_12716);
or U13384 (N_13384,N_12872,N_12898);
nor U13385 (N_13385,N_12915,N_12688);
nand U13386 (N_13386,N_12684,N_12531);
and U13387 (N_13387,N_12559,N_12874);
xnor U13388 (N_13388,N_12573,N_12744);
nand U13389 (N_13389,N_12786,N_12516);
nor U13390 (N_13390,N_12697,N_12635);
xnor U13391 (N_13391,N_12705,N_12532);
and U13392 (N_13392,N_12601,N_12974);
nand U13393 (N_13393,N_12609,N_12576);
or U13394 (N_13394,N_12547,N_12902);
and U13395 (N_13395,N_12922,N_12573);
or U13396 (N_13396,N_12904,N_12682);
nor U13397 (N_13397,N_12638,N_12920);
nor U13398 (N_13398,N_12617,N_12933);
and U13399 (N_13399,N_12946,N_12658);
nand U13400 (N_13400,N_12854,N_12646);
and U13401 (N_13401,N_12844,N_12803);
nor U13402 (N_13402,N_12739,N_12611);
and U13403 (N_13403,N_12527,N_12755);
or U13404 (N_13404,N_12629,N_12696);
nand U13405 (N_13405,N_12757,N_12758);
or U13406 (N_13406,N_12604,N_12953);
nand U13407 (N_13407,N_12823,N_12948);
nand U13408 (N_13408,N_12536,N_12551);
xor U13409 (N_13409,N_12706,N_12634);
nor U13410 (N_13410,N_12943,N_12773);
and U13411 (N_13411,N_12765,N_12921);
xor U13412 (N_13412,N_12704,N_12649);
nand U13413 (N_13413,N_12837,N_12985);
xnor U13414 (N_13414,N_12568,N_12559);
xnor U13415 (N_13415,N_12665,N_12817);
or U13416 (N_13416,N_12753,N_12505);
nand U13417 (N_13417,N_12744,N_12758);
xor U13418 (N_13418,N_12975,N_12917);
and U13419 (N_13419,N_12675,N_12994);
or U13420 (N_13420,N_12520,N_12968);
or U13421 (N_13421,N_12839,N_12524);
nand U13422 (N_13422,N_12889,N_12558);
nand U13423 (N_13423,N_12987,N_12755);
or U13424 (N_13424,N_12605,N_12553);
and U13425 (N_13425,N_12992,N_12621);
nand U13426 (N_13426,N_12981,N_12913);
or U13427 (N_13427,N_12707,N_12890);
nand U13428 (N_13428,N_12723,N_12903);
xor U13429 (N_13429,N_12739,N_12740);
nor U13430 (N_13430,N_12514,N_12619);
or U13431 (N_13431,N_12563,N_12628);
nor U13432 (N_13432,N_12832,N_12565);
nor U13433 (N_13433,N_12802,N_12591);
xor U13434 (N_13434,N_12754,N_12731);
or U13435 (N_13435,N_12503,N_12653);
and U13436 (N_13436,N_12652,N_12708);
and U13437 (N_13437,N_12650,N_12837);
xor U13438 (N_13438,N_12749,N_12684);
and U13439 (N_13439,N_12500,N_12929);
xnor U13440 (N_13440,N_12669,N_12560);
xnor U13441 (N_13441,N_12737,N_12558);
or U13442 (N_13442,N_12679,N_12756);
and U13443 (N_13443,N_12723,N_12963);
nand U13444 (N_13444,N_12687,N_12714);
nor U13445 (N_13445,N_12871,N_12504);
or U13446 (N_13446,N_12843,N_12612);
nand U13447 (N_13447,N_12987,N_12685);
nand U13448 (N_13448,N_12974,N_12813);
nand U13449 (N_13449,N_12561,N_12769);
nand U13450 (N_13450,N_12731,N_12787);
nand U13451 (N_13451,N_12843,N_12918);
nor U13452 (N_13452,N_12633,N_12648);
and U13453 (N_13453,N_12688,N_12645);
xor U13454 (N_13454,N_12572,N_12603);
nor U13455 (N_13455,N_12936,N_12679);
and U13456 (N_13456,N_12668,N_12964);
xnor U13457 (N_13457,N_12998,N_12861);
nand U13458 (N_13458,N_12749,N_12766);
nand U13459 (N_13459,N_12657,N_12740);
nand U13460 (N_13460,N_12774,N_12712);
or U13461 (N_13461,N_12970,N_12881);
and U13462 (N_13462,N_12707,N_12910);
and U13463 (N_13463,N_12537,N_12914);
or U13464 (N_13464,N_12974,N_12801);
xor U13465 (N_13465,N_12531,N_12553);
nor U13466 (N_13466,N_12964,N_12671);
nand U13467 (N_13467,N_12596,N_12866);
or U13468 (N_13468,N_12643,N_12827);
or U13469 (N_13469,N_12741,N_12542);
nor U13470 (N_13470,N_12586,N_12542);
nand U13471 (N_13471,N_12541,N_12732);
xnor U13472 (N_13472,N_12760,N_12561);
xnor U13473 (N_13473,N_12991,N_12562);
or U13474 (N_13474,N_12638,N_12985);
or U13475 (N_13475,N_12917,N_12551);
or U13476 (N_13476,N_12695,N_12775);
and U13477 (N_13477,N_12670,N_12538);
or U13478 (N_13478,N_12604,N_12853);
nand U13479 (N_13479,N_12857,N_12864);
nand U13480 (N_13480,N_12894,N_12743);
or U13481 (N_13481,N_12937,N_12527);
nand U13482 (N_13482,N_12973,N_12738);
nand U13483 (N_13483,N_12843,N_12974);
xnor U13484 (N_13484,N_12778,N_12713);
or U13485 (N_13485,N_12886,N_12732);
nor U13486 (N_13486,N_12525,N_12720);
nand U13487 (N_13487,N_12593,N_12729);
nor U13488 (N_13488,N_12515,N_12880);
nor U13489 (N_13489,N_12585,N_12640);
or U13490 (N_13490,N_12655,N_12533);
nor U13491 (N_13491,N_12713,N_12741);
nand U13492 (N_13492,N_12942,N_12543);
and U13493 (N_13493,N_12583,N_12946);
xor U13494 (N_13494,N_12610,N_12566);
nand U13495 (N_13495,N_12748,N_12768);
xor U13496 (N_13496,N_12773,N_12951);
and U13497 (N_13497,N_12966,N_12511);
or U13498 (N_13498,N_12868,N_12513);
nand U13499 (N_13499,N_12963,N_12964);
and U13500 (N_13500,N_13230,N_13098);
and U13501 (N_13501,N_13185,N_13199);
or U13502 (N_13502,N_13457,N_13276);
nor U13503 (N_13503,N_13122,N_13130);
xnor U13504 (N_13504,N_13260,N_13488);
nor U13505 (N_13505,N_13176,N_13269);
nor U13506 (N_13506,N_13053,N_13338);
nand U13507 (N_13507,N_13479,N_13118);
nor U13508 (N_13508,N_13080,N_13412);
xnor U13509 (N_13509,N_13375,N_13351);
or U13510 (N_13510,N_13154,N_13440);
or U13511 (N_13511,N_13366,N_13107);
nand U13512 (N_13512,N_13277,N_13064);
xnor U13513 (N_13513,N_13310,N_13234);
xor U13514 (N_13514,N_13026,N_13158);
nor U13515 (N_13515,N_13293,N_13051);
xor U13516 (N_13516,N_13301,N_13240);
xnor U13517 (N_13517,N_13494,N_13490);
and U13518 (N_13518,N_13177,N_13091);
and U13519 (N_13519,N_13078,N_13453);
xor U13520 (N_13520,N_13447,N_13413);
and U13521 (N_13521,N_13133,N_13034);
nor U13522 (N_13522,N_13170,N_13493);
nand U13523 (N_13523,N_13065,N_13250);
xor U13524 (N_13524,N_13278,N_13031);
or U13525 (N_13525,N_13332,N_13265);
nand U13526 (N_13526,N_13329,N_13465);
xor U13527 (N_13527,N_13152,N_13414);
or U13528 (N_13528,N_13268,N_13295);
nand U13529 (N_13529,N_13280,N_13448);
nand U13530 (N_13530,N_13027,N_13491);
xnor U13531 (N_13531,N_13073,N_13344);
nand U13532 (N_13532,N_13151,N_13178);
and U13533 (N_13533,N_13258,N_13405);
nor U13534 (N_13534,N_13229,N_13473);
nor U13535 (N_13535,N_13458,N_13009);
or U13536 (N_13536,N_13474,N_13377);
nand U13537 (N_13537,N_13323,N_13367);
or U13538 (N_13538,N_13285,N_13005);
nor U13539 (N_13539,N_13215,N_13043);
xnor U13540 (N_13540,N_13181,N_13341);
or U13541 (N_13541,N_13320,N_13114);
or U13542 (N_13542,N_13356,N_13401);
nor U13543 (N_13543,N_13291,N_13217);
and U13544 (N_13544,N_13220,N_13451);
xor U13545 (N_13545,N_13007,N_13013);
nor U13546 (N_13546,N_13456,N_13049);
and U13547 (N_13547,N_13436,N_13101);
and U13548 (N_13548,N_13339,N_13120);
and U13549 (N_13549,N_13259,N_13106);
xor U13550 (N_13550,N_13183,N_13407);
or U13551 (N_13551,N_13316,N_13334);
nand U13552 (N_13552,N_13076,N_13104);
nor U13553 (N_13553,N_13109,N_13205);
nand U13554 (N_13554,N_13161,N_13153);
nand U13555 (N_13555,N_13175,N_13000);
or U13556 (N_13556,N_13214,N_13206);
and U13557 (N_13557,N_13054,N_13201);
nor U13558 (N_13558,N_13068,N_13385);
and U13559 (N_13559,N_13040,N_13237);
and U13560 (N_13560,N_13195,N_13135);
or U13561 (N_13561,N_13357,N_13388);
xor U13562 (N_13562,N_13470,N_13372);
nand U13563 (N_13563,N_13108,N_13184);
or U13564 (N_13564,N_13012,N_13055);
xor U13565 (N_13565,N_13204,N_13390);
and U13566 (N_13566,N_13402,N_13305);
xnor U13567 (N_13567,N_13330,N_13431);
and U13568 (N_13568,N_13089,N_13452);
and U13569 (N_13569,N_13428,N_13358);
xnor U13570 (N_13570,N_13125,N_13062);
or U13571 (N_13571,N_13123,N_13324);
xnor U13572 (N_13572,N_13492,N_13124);
nor U13573 (N_13573,N_13117,N_13315);
nand U13574 (N_13574,N_13166,N_13111);
nor U13575 (N_13575,N_13126,N_13409);
xnor U13576 (N_13576,N_13360,N_13266);
nand U13577 (N_13577,N_13001,N_13248);
xor U13578 (N_13578,N_13231,N_13219);
nand U13579 (N_13579,N_13383,N_13096);
or U13580 (N_13580,N_13198,N_13264);
xnor U13581 (N_13581,N_13289,N_13081);
and U13582 (N_13582,N_13174,N_13016);
nand U13583 (N_13583,N_13397,N_13059);
or U13584 (N_13584,N_13032,N_13483);
nand U13585 (N_13585,N_13411,N_13300);
nor U13586 (N_13586,N_13050,N_13380);
or U13587 (N_13587,N_13480,N_13399);
nor U13588 (N_13588,N_13134,N_13398);
xor U13589 (N_13589,N_13283,N_13066);
and U13590 (N_13590,N_13203,N_13128);
nand U13591 (N_13591,N_13381,N_13193);
nand U13592 (N_13592,N_13370,N_13481);
or U13593 (N_13593,N_13311,N_13461);
nor U13594 (N_13594,N_13086,N_13349);
nand U13595 (N_13595,N_13226,N_13342);
nand U13596 (N_13596,N_13189,N_13247);
xor U13597 (N_13597,N_13365,N_13438);
xnor U13598 (N_13598,N_13468,N_13200);
or U13599 (N_13599,N_13030,N_13450);
nor U13600 (N_13600,N_13218,N_13420);
or U13601 (N_13601,N_13004,N_13477);
xnor U13602 (N_13602,N_13116,N_13037);
nor U13603 (N_13603,N_13466,N_13057);
xor U13604 (N_13604,N_13426,N_13395);
or U13605 (N_13605,N_13225,N_13352);
nor U13606 (N_13606,N_13322,N_13239);
nand U13607 (N_13607,N_13441,N_13262);
and U13608 (N_13608,N_13484,N_13121);
nor U13609 (N_13609,N_13303,N_13029);
and U13610 (N_13610,N_13169,N_13403);
nor U13611 (N_13611,N_13139,N_13256);
nor U13612 (N_13612,N_13254,N_13298);
nand U13613 (N_13613,N_13343,N_13495);
nand U13614 (N_13614,N_13286,N_13314);
nand U13615 (N_13615,N_13228,N_13171);
xor U13616 (N_13616,N_13213,N_13319);
nand U13617 (N_13617,N_13362,N_13485);
or U13618 (N_13618,N_13039,N_13434);
xnor U13619 (N_13619,N_13296,N_13389);
xor U13620 (N_13620,N_13449,N_13041);
nand U13621 (N_13621,N_13318,N_13163);
or U13622 (N_13622,N_13140,N_13425);
nor U13623 (N_13623,N_13348,N_13267);
nand U13624 (N_13624,N_13088,N_13423);
xor U13625 (N_13625,N_13359,N_13432);
xnor U13626 (N_13626,N_13421,N_13384);
and U13627 (N_13627,N_13025,N_13442);
or U13628 (N_13628,N_13036,N_13061);
xor U13629 (N_13629,N_13033,N_13083);
nand U13630 (N_13630,N_13015,N_13261);
nor U13631 (N_13631,N_13306,N_13345);
nor U13632 (N_13632,N_13075,N_13227);
nand U13633 (N_13633,N_13246,N_13454);
nand U13634 (N_13634,N_13326,N_13327);
nand U13635 (N_13635,N_13340,N_13090);
and U13636 (N_13636,N_13287,N_13424);
and U13637 (N_13637,N_13044,N_13475);
xnor U13638 (N_13638,N_13263,N_13003);
or U13639 (N_13639,N_13346,N_13058);
nor U13640 (N_13640,N_13202,N_13238);
and U13641 (N_13641,N_13071,N_13018);
or U13642 (N_13642,N_13404,N_13060);
nand U13643 (N_13643,N_13476,N_13355);
nor U13644 (N_13644,N_13353,N_13144);
and U13645 (N_13645,N_13222,N_13212);
xor U13646 (N_13646,N_13284,N_13095);
and U13647 (N_13647,N_13325,N_13241);
nand U13648 (N_13648,N_13006,N_13435);
xnor U13649 (N_13649,N_13354,N_13087);
or U13650 (N_13650,N_13136,N_13471);
xnor U13651 (N_13651,N_13371,N_13188);
nand U13652 (N_13652,N_13197,N_13145);
and U13653 (N_13653,N_13167,N_13072);
nand U13654 (N_13654,N_13251,N_13244);
or U13655 (N_13655,N_13499,N_13186);
nor U13656 (N_13656,N_13379,N_13419);
nand U13657 (N_13657,N_13321,N_13085);
or U13658 (N_13658,N_13410,N_13460);
xor U13659 (N_13659,N_13275,N_13069);
nand U13660 (N_13660,N_13022,N_13270);
or U13661 (N_13661,N_13308,N_13331);
xnor U13662 (N_13662,N_13047,N_13444);
nand U13663 (N_13663,N_13496,N_13363);
nor U13664 (N_13664,N_13211,N_13093);
nor U13665 (N_13665,N_13112,N_13313);
nor U13666 (N_13666,N_13232,N_13074);
or U13667 (N_13667,N_13079,N_13021);
or U13668 (N_13668,N_13035,N_13459);
nand U13669 (N_13669,N_13317,N_13307);
or U13670 (N_13670,N_13223,N_13048);
xor U13671 (N_13671,N_13019,N_13290);
nand U13672 (N_13672,N_13418,N_13427);
xor U13673 (N_13673,N_13209,N_13417);
nor U13674 (N_13674,N_13462,N_13196);
or U13675 (N_13675,N_13067,N_13100);
or U13676 (N_13676,N_13392,N_13486);
and U13677 (N_13677,N_13002,N_13023);
and U13678 (N_13678,N_13180,N_13156);
and U13679 (N_13679,N_13252,N_13396);
nor U13680 (N_13680,N_13257,N_13393);
nand U13681 (N_13681,N_13155,N_13302);
nor U13682 (N_13682,N_13309,N_13092);
nand U13683 (N_13683,N_13373,N_13221);
nor U13684 (N_13684,N_13210,N_13110);
xnor U13685 (N_13685,N_13235,N_13439);
xnor U13686 (N_13686,N_13113,N_13017);
nor U13687 (N_13687,N_13386,N_13445);
and U13688 (N_13688,N_13281,N_13347);
and U13689 (N_13689,N_13408,N_13129);
xnor U13690 (N_13690,N_13143,N_13378);
nor U13691 (N_13691,N_13008,N_13160);
nand U13692 (N_13692,N_13224,N_13253);
nand U13693 (N_13693,N_13020,N_13288);
or U13694 (N_13694,N_13046,N_13446);
xnor U13695 (N_13695,N_13333,N_13159);
nand U13696 (N_13696,N_13455,N_13255);
nand U13697 (N_13697,N_13374,N_13187);
xnor U13698 (N_13698,N_13115,N_13028);
or U13699 (N_13699,N_13131,N_13472);
or U13700 (N_13700,N_13245,N_13437);
and U13701 (N_13701,N_13103,N_13394);
nor U13702 (N_13702,N_13304,N_13147);
or U13703 (N_13703,N_13146,N_13097);
nand U13704 (N_13704,N_13182,N_13282);
or U13705 (N_13705,N_13045,N_13038);
xor U13706 (N_13706,N_13070,N_13132);
nand U13707 (N_13707,N_13119,N_13024);
xor U13708 (N_13708,N_13207,N_13216);
and U13709 (N_13709,N_13084,N_13142);
and U13710 (N_13710,N_13272,N_13094);
nor U13711 (N_13711,N_13063,N_13497);
xor U13712 (N_13712,N_13077,N_13279);
xnor U13713 (N_13713,N_13082,N_13292);
or U13714 (N_13714,N_13336,N_13489);
and U13715 (N_13715,N_13328,N_13312);
nand U13716 (N_13716,N_13137,N_13478);
and U13717 (N_13717,N_13376,N_13274);
and U13718 (N_13718,N_13194,N_13463);
xnor U13719 (N_13719,N_13191,N_13249);
or U13720 (N_13720,N_13387,N_13297);
or U13721 (N_13721,N_13422,N_13138);
and U13722 (N_13722,N_13369,N_13148);
nor U13723 (N_13723,N_13102,N_13105);
nor U13724 (N_13724,N_13416,N_13391);
nand U13725 (N_13725,N_13406,N_13052);
xnor U13726 (N_13726,N_13192,N_13242);
or U13727 (N_13727,N_13236,N_13173);
xnor U13728 (N_13728,N_13168,N_13299);
or U13729 (N_13729,N_13350,N_13010);
nand U13730 (N_13730,N_13482,N_13400);
xnor U13731 (N_13731,N_13150,N_13487);
xor U13732 (N_13732,N_13208,N_13172);
xor U13733 (N_13733,N_13056,N_13271);
and U13734 (N_13734,N_13233,N_13364);
and U13735 (N_13735,N_13179,N_13433);
or U13736 (N_13736,N_13368,N_13157);
xnor U13737 (N_13737,N_13165,N_13011);
xnor U13738 (N_13738,N_13149,N_13294);
nor U13739 (N_13739,N_13430,N_13361);
and U13740 (N_13740,N_13127,N_13469);
or U13741 (N_13741,N_13382,N_13464);
nor U13742 (N_13742,N_13415,N_13014);
and U13743 (N_13743,N_13099,N_13243);
or U13744 (N_13744,N_13498,N_13273);
nor U13745 (N_13745,N_13335,N_13164);
xnor U13746 (N_13746,N_13443,N_13141);
or U13747 (N_13747,N_13042,N_13190);
xnor U13748 (N_13748,N_13337,N_13162);
nor U13749 (N_13749,N_13429,N_13467);
nand U13750 (N_13750,N_13317,N_13239);
or U13751 (N_13751,N_13169,N_13359);
or U13752 (N_13752,N_13273,N_13390);
and U13753 (N_13753,N_13090,N_13164);
and U13754 (N_13754,N_13464,N_13431);
nor U13755 (N_13755,N_13367,N_13115);
and U13756 (N_13756,N_13184,N_13219);
or U13757 (N_13757,N_13314,N_13148);
nand U13758 (N_13758,N_13067,N_13473);
nand U13759 (N_13759,N_13185,N_13181);
nand U13760 (N_13760,N_13398,N_13124);
nand U13761 (N_13761,N_13379,N_13001);
xor U13762 (N_13762,N_13399,N_13366);
or U13763 (N_13763,N_13145,N_13475);
and U13764 (N_13764,N_13270,N_13146);
or U13765 (N_13765,N_13019,N_13241);
and U13766 (N_13766,N_13451,N_13180);
nor U13767 (N_13767,N_13382,N_13353);
xnor U13768 (N_13768,N_13113,N_13485);
nand U13769 (N_13769,N_13200,N_13393);
nand U13770 (N_13770,N_13129,N_13402);
nand U13771 (N_13771,N_13308,N_13133);
xor U13772 (N_13772,N_13176,N_13405);
nor U13773 (N_13773,N_13292,N_13488);
or U13774 (N_13774,N_13008,N_13212);
xor U13775 (N_13775,N_13193,N_13283);
or U13776 (N_13776,N_13393,N_13072);
nand U13777 (N_13777,N_13270,N_13370);
nand U13778 (N_13778,N_13026,N_13491);
or U13779 (N_13779,N_13374,N_13348);
nand U13780 (N_13780,N_13111,N_13114);
and U13781 (N_13781,N_13111,N_13374);
or U13782 (N_13782,N_13456,N_13438);
or U13783 (N_13783,N_13005,N_13106);
or U13784 (N_13784,N_13116,N_13258);
xor U13785 (N_13785,N_13455,N_13121);
xor U13786 (N_13786,N_13078,N_13291);
and U13787 (N_13787,N_13399,N_13467);
nor U13788 (N_13788,N_13257,N_13010);
nor U13789 (N_13789,N_13192,N_13022);
and U13790 (N_13790,N_13012,N_13196);
nand U13791 (N_13791,N_13032,N_13315);
or U13792 (N_13792,N_13257,N_13269);
xnor U13793 (N_13793,N_13273,N_13267);
xor U13794 (N_13794,N_13249,N_13396);
and U13795 (N_13795,N_13123,N_13242);
or U13796 (N_13796,N_13214,N_13466);
nor U13797 (N_13797,N_13213,N_13468);
nor U13798 (N_13798,N_13187,N_13015);
or U13799 (N_13799,N_13060,N_13280);
nand U13800 (N_13800,N_13338,N_13194);
xnor U13801 (N_13801,N_13000,N_13382);
or U13802 (N_13802,N_13481,N_13145);
xnor U13803 (N_13803,N_13428,N_13093);
nor U13804 (N_13804,N_13375,N_13067);
or U13805 (N_13805,N_13138,N_13293);
or U13806 (N_13806,N_13004,N_13492);
and U13807 (N_13807,N_13308,N_13009);
and U13808 (N_13808,N_13271,N_13320);
or U13809 (N_13809,N_13435,N_13493);
nand U13810 (N_13810,N_13245,N_13216);
xnor U13811 (N_13811,N_13031,N_13252);
xnor U13812 (N_13812,N_13271,N_13018);
or U13813 (N_13813,N_13344,N_13430);
nand U13814 (N_13814,N_13449,N_13269);
nand U13815 (N_13815,N_13328,N_13497);
or U13816 (N_13816,N_13302,N_13475);
or U13817 (N_13817,N_13216,N_13302);
or U13818 (N_13818,N_13384,N_13276);
and U13819 (N_13819,N_13204,N_13087);
nor U13820 (N_13820,N_13261,N_13307);
nand U13821 (N_13821,N_13452,N_13497);
nor U13822 (N_13822,N_13086,N_13499);
or U13823 (N_13823,N_13110,N_13141);
xnor U13824 (N_13824,N_13086,N_13032);
nor U13825 (N_13825,N_13012,N_13000);
xnor U13826 (N_13826,N_13251,N_13449);
xnor U13827 (N_13827,N_13143,N_13258);
or U13828 (N_13828,N_13338,N_13496);
nand U13829 (N_13829,N_13194,N_13072);
nor U13830 (N_13830,N_13161,N_13487);
nand U13831 (N_13831,N_13013,N_13063);
or U13832 (N_13832,N_13457,N_13001);
or U13833 (N_13833,N_13491,N_13401);
and U13834 (N_13834,N_13426,N_13142);
nand U13835 (N_13835,N_13027,N_13001);
and U13836 (N_13836,N_13162,N_13358);
or U13837 (N_13837,N_13172,N_13002);
or U13838 (N_13838,N_13137,N_13366);
nand U13839 (N_13839,N_13416,N_13358);
nor U13840 (N_13840,N_13014,N_13344);
nand U13841 (N_13841,N_13196,N_13430);
nand U13842 (N_13842,N_13429,N_13280);
xnor U13843 (N_13843,N_13312,N_13178);
nor U13844 (N_13844,N_13069,N_13141);
nand U13845 (N_13845,N_13200,N_13452);
and U13846 (N_13846,N_13315,N_13041);
and U13847 (N_13847,N_13134,N_13297);
or U13848 (N_13848,N_13388,N_13184);
or U13849 (N_13849,N_13310,N_13145);
and U13850 (N_13850,N_13289,N_13467);
xor U13851 (N_13851,N_13422,N_13151);
or U13852 (N_13852,N_13228,N_13204);
nand U13853 (N_13853,N_13050,N_13156);
nor U13854 (N_13854,N_13056,N_13046);
nand U13855 (N_13855,N_13454,N_13326);
and U13856 (N_13856,N_13054,N_13374);
nor U13857 (N_13857,N_13145,N_13170);
nand U13858 (N_13858,N_13327,N_13033);
nand U13859 (N_13859,N_13300,N_13284);
or U13860 (N_13860,N_13125,N_13354);
xnor U13861 (N_13861,N_13259,N_13454);
or U13862 (N_13862,N_13048,N_13016);
nor U13863 (N_13863,N_13110,N_13243);
xnor U13864 (N_13864,N_13430,N_13279);
nor U13865 (N_13865,N_13385,N_13393);
or U13866 (N_13866,N_13016,N_13152);
and U13867 (N_13867,N_13189,N_13369);
nor U13868 (N_13868,N_13488,N_13101);
xnor U13869 (N_13869,N_13195,N_13276);
nor U13870 (N_13870,N_13033,N_13146);
or U13871 (N_13871,N_13487,N_13106);
nor U13872 (N_13872,N_13076,N_13251);
nand U13873 (N_13873,N_13031,N_13080);
and U13874 (N_13874,N_13156,N_13308);
nor U13875 (N_13875,N_13327,N_13179);
xor U13876 (N_13876,N_13020,N_13075);
or U13877 (N_13877,N_13470,N_13163);
nand U13878 (N_13878,N_13374,N_13071);
xnor U13879 (N_13879,N_13447,N_13446);
nand U13880 (N_13880,N_13164,N_13248);
nor U13881 (N_13881,N_13174,N_13275);
and U13882 (N_13882,N_13224,N_13182);
nand U13883 (N_13883,N_13496,N_13336);
xor U13884 (N_13884,N_13473,N_13351);
and U13885 (N_13885,N_13384,N_13464);
xor U13886 (N_13886,N_13309,N_13182);
nor U13887 (N_13887,N_13467,N_13344);
nand U13888 (N_13888,N_13454,N_13173);
nor U13889 (N_13889,N_13262,N_13471);
nor U13890 (N_13890,N_13110,N_13367);
or U13891 (N_13891,N_13320,N_13411);
xor U13892 (N_13892,N_13313,N_13361);
or U13893 (N_13893,N_13188,N_13372);
or U13894 (N_13894,N_13238,N_13444);
or U13895 (N_13895,N_13325,N_13031);
or U13896 (N_13896,N_13280,N_13251);
and U13897 (N_13897,N_13135,N_13086);
xor U13898 (N_13898,N_13351,N_13426);
and U13899 (N_13899,N_13200,N_13029);
or U13900 (N_13900,N_13102,N_13096);
or U13901 (N_13901,N_13135,N_13083);
xnor U13902 (N_13902,N_13454,N_13398);
nor U13903 (N_13903,N_13469,N_13060);
and U13904 (N_13904,N_13290,N_13393);
and U13905 (N_13905,N_13008,N_13307);
and U13906 (N_13906,N_13493,N_13343);
or U13907 (N_13907,N_13267,N_13423);
xor U13908 (N_13908,N_13342,N_13043);
and U13909 (N_13909,N_13473,N_13187);
nand U13910 (N_13910,N_13089,N_13140);
or U13911 (N_13911,N_13483,N_13361);
nand U13912 (N_13912,N_13388,N_13390);
nand U13913 (N_13913,N_13383,N_13079);
xnor U13914 (N_13914,N_13163,N_13092);
xor U13915 (N_13915,N_13195,N_13157);
and U13916 (N_13916,N_13384,N_13105);
and U13917 (N_13917,N_13076,N_13445);
nand U13918 (N_13918,N_13296,N_13103);
xor U13919 (N_13919,N_13478,N_13088);
xor U13920 (N_13920,N_13036,N_13147);
nor U13921 (N_13921,N_13095,N_13333);
or U13922 (N_13922,N_13318,N_13162);
nand U13923 (N_13923,N_13326,N_13317);
nand U13924 (N_13924,N_13143,N_13137);
or U13925 (N_13925,N_13499,N_13496);
or U13926 (N_13926,N_13273,N_13113);
xnor U13927 (N_13927,N_13059,N_13071);
xnor U13928 (N_13928,N_13340,N_13349);
nand U13929 (N_13929,N_13362,N_13276);
and U13930 (N_13930,N_13003,N_13364);
xnor U13931 (N_13931,N_13187,N_13429);
nor U13932 (N_13932,N_13089,N_13429);
nand U13933 (N_13933,N_13191,N_13316);
nand U13934 (N_13934,N_13199,N_13457);
nand U13935 (N_13935,N_13001,N_13393);
and U13936 (N_13936,N_13208,N_13027);
nor U13937 (N_13937,N_13442,N_13308);
or U13938 (N_13938,N_13451,N_13313);
xnor U13939 (N_13939,N_13221,N_13054);
nor U13940 (N_13940,N_13322,N_13213);
or U13941 (N_13941,N_13066,N_13185);
nor U13942 (N_13942,N_13160,N_13173);
and U13943 (N_13943,N_13127,N_13296);
and U13944 (N_13944,N_13452,N_13290);
and U13945 (N_13945,N_13036,N_13183);
or U13946 (N_13946,N_13244,N_13330);
and U13947 (N_13947,N_13477,N_13402);
and U13948 (N_13948,N_13126,N_13111);
nor U13949 (N_13949,N_13407,N_13070);
and U13950 (N_13950,N_13204,N_13338);
and U13951 (N_13951,N_13419,N_13341);
or U13952 (N_13952,N_13380,N_13251);
or U13953 (N_13953,N_13431,N_13300);
or U13954 (N_13954,N_13088,N_13105);
and U13955 (N_13955,N_13205,N_13093);
and U13956 (N_13956,N_13416,N_13291);
and U13957 (N_13957,N_13382,N_13478);
or U13958 (N_13958,N_13245,N_13299);
xor U13959 (N_13959,N_13434,N_13142);
nand U13960 (N_13960,N_13150,N_13097);
nor U13961 (N_13961,N_13149,N_13398);
or U13962 (N_13962,N_13367,N_13012);
and U13963 (N_13963,N_13434,N_13125);
nor U13964 (N_13964,N_13174,N_13144);
and U13965 (N_13965,N_13493,N_13217);
or U13966 (N_13966,N_13088,N_13282);
nor U13967 (N_13967,N_13499,N_13282);
nand U13968 (N_13968,N_13162,N_13296);
or U13969 (N_13969,N_13270,N_13494);
nand U13970 (N_13970,N_13250,N_13210);
nand U13971 (N_13971,N_13022,N_13495);
nand U13972 (N_13972,N_13076,N_13147);
and U13973 (N_13973,N_13246,N_13170);
nand U13974 (N_13974,N_13304,N_13296);
nor U13975 (N_13975,N_13279,N_13122);
or U13976 (N_13976,N_13426,N_13400);
xor U13977 (N_13977,N_13018,N_13421);
or U13978 (N_13978,N_13494,N_13473);
or U13979 (N_13979,N_13357,N_13043);
and U13980 (N_13980,N_13432,N_13472);
and U13981 (N_13981,N_13375,N_13161);
nor U13982 (N_13982,N_13122,N_13213);
nor U13983 (N_13983,N_13032,N_13054);
nor U13984 (N_13984,N_13483,N_13038);
nand U13985 (N_13985,N_13239,N_13343);
nor U13986 (N_13986,N_13021,N_13461);
xor U13987 (N_13987,N_13104,N_13343);
xnor U13988 (N_13988,N_13186,N_13347);
and U13989 (N_13989,N_13049,N_13297);
and U13990 (N_13990,N_13170,N_13152);
xnor U13991 (N_13991,N_13356,N_13044);
and U13992 (N_13992,N_13327,N_13092);
nand U13993 (N_13993,N_13400,N_13243);
xnor U13994 (N_13994,N_13051,N_13314);
nand U13995 (N_13995,N_13336,N_13093);
nor U13996 (N_13996,N_13220,N_13333);
nand U13997 (N_13997,N_13012,N_13477);
xor U13998 (N_13998,N_13106,N_13140);
nor U13999 (N_13999,N_13014,N_13225);
and U14000 (N_14000,N_13748,N_13918);
or U14001 (N_14001,N_13515,N_13761);
or U14002 (N_14002,N_13544,N_13874);
or U14003 (N_14003,N_13832,N_13583);
nand U14004 (N_14004,N_13581,N_13893);
and U14005 (N_14005,N_13501,N_13891);
and U14006 (N_14006,N_13680,N_13785);
nand U14007 (N_14007,N_13890,N_13804);
xnor U14008 (N_14008,N_13984,N_13957);
or U14009 (N_14009,N_13749,N_13702);
or U14010 (N_14010,N_13968,N_13799);
and U14011 (N_14011,N_13575,N_13936);
and U14012 (N_14012,N_13925,N_13860);
nand U14013 (N_14013,N_13552,N_13563);
xor U14014 (N_14014,N_13590,N_13762);
xor U14015 (N_14015,N_13753,N_13756);
nand U14016 (N_14016,N_13695,N_13899);
nor U14017 (N_14017,N_13989,N_13873);
or U14018 (N_14018,N_13657,N_13861);
or U14019 (N_14019,N_13933,N_13942);
nor U14020 (N_14020,N_13634,N_13813);
or U14021 (N_14021,N_13580,N_13611);
or U14022 (N_14022,N_13865,N_13682);
xor U14023 (N_14023,N_13676,N_13765);
xnor U14024 (N_14024,N_13913,N_13779);
and U14025 (N_14025,N_13617,N_13642);
nor U14026 (N_14026,N_13632,N_13825);
nand U14027 (N_14027,N_13994,N_13721);
nor U14028 (N_14028,N_13605,N_13710);
nand U14029 (N_14029,N_13754,N_13567);
or U14030 (N_14030,N_13996,N_13606);
xor U14031 (N_14031,N_13621,N_13803);
xnor U14032 (N_14032,N_13595,N_13896);
or U14033 (N_14033,N_13910,N_13693);
nor U14034 (N_14034,N_13908,N_13856);
or U14035 (N_14035,N_13953,N_13921);
nor U14036 (N_14036,N_13585,N_13817);
and U14037 (N_14037,N_13539,N_13673);
or U14038 (N_14038,N_13938,N_13919);
and U14039 (N_14039,N_13979,N_13841);
or U14040 (N_14040,N_13559,N_13698);
or U14041 (N_14041,N_13780,N_13558);
and U14042 (N_14042,N_13616,N_13724);
nand U14043 (N_14043,N_13985,N_13823);
nor U14044 (N_14044,N_13986,N_13534);
xnor U14045 (N_14045,N_13728,N_13808);
xnor U14046 (N_14046,N_13707,N_13742);
and U14047 (N_14047,N_13751,N_13527);
nand U14048 (N_14048,N_13647,N_13653);
and U14049 (N_14049,N_13871,N_13665);
nor U14050 (N_14050,N_13814,N_13509);
nor U14051 (N_14051,N_13589,N_13988);
or U14052 (N_14052,N_13939,N_13935);
nor U14053 (N_14053,N_13648,N_13758);
and U14054 (N_14054,N_13679,N_13579);
and U14055 (N_14055,N_13533,N_13556);
and U14056 (N_14056,N_13858,N_13535);
xnor U14057 (N_14057,N_13626,N_13880);
and U14058 (N_14058,N_13675,N_13674);
xnor U14059 (N_14059,N_13637,N_13571);
and U14060 (N_14060,N_13798,N_13564);
and U14061 (N_14061,N_13949,N_13592);
xnor U14062 (N_14062,N_13655,N_13965);
or U14063 (N_14063,N_13517,N_13900);
and U14064 (N_14064,N_13594,N_13663);
and U14065 (N_14065,N_13809,N_13875);
nand U14066 (N_14066,N_13639,N_13864);
nand U14067 (N_14067,N_13969,N_13999);
or U14068 (N_14068,N_13706,N_13725);
nor U14069 (N_14069,N_13755,N_13739);
nand U14070 (N_14070,N_13981,N_13694);
nand U14071 (N_14071,N_13628,N_13831);
and U14072 (N_14072,N_13568,N_13777);
nand U14073 (N_14073,N_13894,N_13800);
xor U14074 (N_14074,N_13738,N_13726);
and U14075 (N_14075,N_13962,N_13767);
or U14076 (N_14076,N_13670,N_13811);
nand U14077 (N_14077,N_13541,N_13772);
xor U14078 (N_14078,N_13623,N_13946);
xor U14079 (N_14079,N_13795,N_13652);
xor U14080 (N_14080,N_13818,N_13542);
or U14081 (N_14081,N_13960,N_13995);
and U14082 (N_14082,N_13505,N_13796);
and U14083 (N_14083,N_13862,N_13669);
and U14084 (N_14084,N_13712,N_13897);
nand U14085 (N_14085,N_13993,N_13783);
xnor U14086 (N_14086,N_13692,N_13743);
or U14087 (N_14087,N_13850,N_13930);
xnor U14088 (N_14088,N_13516,N_13781);
nor U14089 (N_14089,N_13826,N_13704);
xor U14090 (N_14090,N_13855,N_13554);
or U14091 (N_14091,N_13760,N_13645);
nor U14092 (N_14092,N_13500,N_13685);
nand U14093 (N_14093,N_13906,N_13833);
and U14094 (N_14094,N_13598,N_13518);
xnor U14095 (N_14095,N_13502,N_13883);
xor U14096 (N_14096,N_13603,N_13786);
xnor U14097 (N_14097,N_13869,N_13846);
nor U14098 (N_14098,N_13536,N_13876);
or U14099 (N_14099,N_13610,N_13773);
nor U14100 (N_14100,N_13717,N_13895);
xnor U14101 (N_14101,N_13591,N_13976);
nor U14102 (N_14102,N_13940,N_13952);
or U14103 (N_14103,N_13577,N_13911);
or U14104 (N_14104,N_13678,N_13904);
xnor U14105 (N_14105,N_13565,N_13889);
nor U14106 (N_14106,N_13791,N_13683);
and U14107 (N_14107,N_13787,N_13790);
nand U14108 (N_14108,N_13863,N_13792);
nand U14109 (N_14109,N_13914,N_13966);
xnor U14110 (N_14110,N_13766,N_13715);
xor U14111 (N_14111,N_13703,N_13625);
or U14112 (N_14112,N_13691,N_13820);
and U14113 (N_14113,N_13987,N_13569);
xor U14114 (N_14114,N_13633,N_13711);
nand U14115 (N_14115,N_13593,N_13572);
or U14116 (N_14116,N_13801,N_13584);
nand U14117 (N_14117,N_13723,N_13805);
nand U14118 (N_14118,N_13506,N_13708);
or U14119 (N_14119,N_13822,N_13700);
nor U14120 (N_14120,N_13638,N_13955);
nand U14121 (N_14121,N_13870,N_13614);
nand U14122 (N_14122,N_13838,N_13526);
or U14123 (N_14123,N_13696,N_13973);
nor U14124 (N_14124,N_13643,N_13608);
xor U14125 (N_14125,N_13847,N_13757);
nand U14126 (N_14126,N_13654,N_13510);
xor U14127 (N_14127,N_13943,N_13701);
or U14128 (N_14128,N_13980,N_13576);
or U14129 (N_14129,N_13888,N_13821);
nor U14130 (N_14130,N_13884,N_13937);
nor U14131 (N_14131,N_13546,N_13523);
nor U14132 (N_14132,N_13731,N_13551);
xnor U14133 (N_14133,N_13834,N_13956);
and U14134 (N_14134,N_13521,N_13615);
and U14135 (N_14135,N_13970,N_13944);
nand U14136 (N_14136,N_13882,N_13793);
xor U14137 (N_14137,N_13902,N_13845);
and U14138 (N_14138,N_13774,N_13529);
and U14139 (N_14139,N_13802,N_13531);
nand U14140 (N_14140,N_13901,N_13684);
xor U14141 (N_14141,N_13978,N_13797);
or U14142 (N_14142,N_13836,N_13961);
nand U14143 (N_14143,N_13532,N_13636);
nor U14144 (N_14144,N_13697,N_13954);
nor U14145 (N_14145,N_13649,N_13794);
and U14146 (N_14146,N_13658,N_13829);
or U14147 (N_14147,N_13714,N_13624);
xnor U14148 (N_14148,N_13664,N_13807);
xor U14149 (N_14149,N_13746,N_13612);
or U14150 (N_14150,N_13540,N_13926);
xnor U14151 (N_14151,N_13932,N_13646);
and U14152 (N_14152,N_13892,N_13732);
or U14153 (N_14153,N_13844,N_13992);
nor U14154 (N_14154,N_13827,N_13602);
nor U14155 (N_14155,N_13548,N_13514);
nand U14156 (N_14156,N_13771,N_13690);
xnor U14157 (N_14157,N_13924,N_13828);
and U14158 (N_14158,N_13503,N_13709);
xor U14159 (N_14159,N_13991,N_13644);
nor U14160 (N_14160,N_13600,N_13784);
nand U14161 (N_14161,N_13782,N_13830);
or U14162 (N_14162,N_13736,N_13549);
nor U14163 (N_14163,N_13522,N_13843);
or U14164 (N_14164,N_13586,N_13607);
nor U14165 (N_14165,N_13635,N_13705);
and U14166 (N_14166,N_13916,N_13967);
nor U14167 (N_14167,N_13768,N_13618);
or U14168 (N_14168,N_13997,N_13839);
nand U14169 (N_14169,N_13713,N_13689);
nor U14170 (N_14170,N_13806,N_13513);
or U14171 (N_14171,N_13859,N_13974);
xor U14172 (N_14172,N_13641,N_13963);
and U14173 (N_14173,N_13912,N_13759);
or U14174 (N_14174,N_13789,N_13866);
and U14175 (N_14175,N_13613,N_13666);
or U14176 (N_14176,N_13920,N_13842);
nor U14177 (N_14177,N_13819,N_13630);
and U14178 (N_14178,N_13629,N_13719);
nor U14179 (N_14179,N_13877,N_13915);
and U14180 (N_14180,N_13735,N_13851);
nor U14181 (N_14181,N_13941,N_13776);
or U14182 (N_14182,N_13778,N_13927);
nand U14183 (N_14183,N_13835,N_13727);
or U14184 (N_14184,N_13878,N_13972);
nand U14185 (N_14185,N_13744,N_13601);
xor U14186 (N_14186,N_13686,N_13868);
and U14187 (N_14187,N_13651,N_13917);
or U14188 (N_14188,N_13752,N_13545);
nand U14189 (N_14189,N_13929,N_13729);
and U14190 (N_14190,N_13543,N_13507);
and U14191 (N_14191,N_13677,N_13672);
and U14192 (N_14192,N_13812,N_13547);
nor U14193 (N_14193,N_13815,N_13853);
xnor U14194 (N_14194,N_13597,N_13631);
xnor U14195 (N_14195,N_13504,N_13619);
or U14196 (N_14196,N_13661,N_13627);
or U14197 (N_14197,N_13537,N_13945);
xnor U14198 (N_14198,N_13750,N_13720);
nand U14199 (N_14199,N_13886,N_13971);
xor U14200 (N_14200,N_13668,N_13560);
or U14201 (N_14201,N_13508,N_13857);
or U14202 (N_14202,N_13609,N_13769);
nand U14203 (N_14203,N_13587,N_13745);
xnor U14204 (N_14204,N_13730,N_13553);
or U14205 (N_14205,N_13650,N_13562);
or U14206 (N_14206,N_13722,N_13733);
nor U14207 (N_14207,N_13747,N_13948);
or U14208 (N_14208,N_13950,N_13764);
or U14209 (N_14209,N_13983,N_13982);
or U14210 (N_14210,N_13879,N_13975);
nor U14211 (N_14211,N_13931,N_13620);
or U14212 (N_14212,N_13872,N_13898);
nor U14213 (N_14213,N_13770,N_13582);
xor U14214 (N_14214,N_13604,N_13959);
or U14215 (N_14215,N_13511,N_13566);
or U14216 (N_14216,N_13907,N_13824);
nand U14217 (N_14217,N_13763,N_13775);
xnor U14218 (N_14218,N_13699,N_13848);
or U14219 (N_14219,N_13538,N_13816);
or U14220 (N_14220,N_13687,N_13990);
nor U14221 (N_14221,N_13656,N_13958);
xnor U14222 (N_14222,N_13903,N_13737);
nor U14223 (N_14223,N_13574,N_13561);
xnor U14224 (N_14224,N_13810,N_13688);
or U14225 (N_14225,N_13640,N_13881);
nand U14226 (N_14226,N_13512,N_13928);
nor U14227 (N_14227,N_13977,N_13867);
nand U14228 (N_14228,N_13837,N_13555);
or U14229 (N_14229,N_13530,N_13909);
xor U14230 (N_14230,N_13923,N_13741);
nand U14231 (N_14231,N_13887,N_13599);
nor U14232 (N_14232,N_13525,N_13519);
xor U14233 (N_14233,N_13716,N_13596);
nand U14234 (N_14234,N_13934,N_13788);
and U14235 (N_14235,N_13681,N_13718);
nor U14236 (N_14236,N_13849,N_13667);
nor U14237 (N_14237,N_13922,N_13854);
nor U14238 (N_14238,N_13622,N_13570);
nand U14239 (N_14239,N_13840,N_13524);
nor U14240 (N_14240,N_13520,N_13557);
xnor U14241 (N_14241,N_13852,N_13528);
nor U14242 (N_14242,N_13659,N_13588);
nor U14243 (N_14243,N_13740,N_13905);
nand U14244 (N_14244,N_13998,N_13578);
nand U14245 (N_14245,N_13660,N_13951);
nor U14246 (N_14246,N_13885,N_13734);
xor U14247 (N_14247,N_13671,N_13550);
xnor U14248 (N_14248,N_13947,N_13964);
and U14249 (N_14249,N_13662,N_13573);
or U14250 (N_14250,N_13950,N_13581);
nor U14251 (N_14251,N_13900,N_13764);
and U14252 (N_14252,N_13708,N_13580);
and U14253 (N_14253,N_13626,N_13755);
nand U14254 (N_14254,N_13993,N_13695);
xor U14255 (N_14255,N_13720,N_13978);
nor U14256 (N_14256,N_13523,N_13741);
nand U14257 (N_14257,N_13968,N_13535);
and U14258 (N_14258,N_13751,N_13772);
nand U14259 (N_14259,N_13561,N_13879);
or U14260 (N_14260,N_13631,N_13849);
xnor U14261 (N_14261,N_13628,N_13547);
or U14262 (N_14262,N_13827,N_13619);
nand U14263 (N_14263,N_13755,N_13587);
nand U14264 (N_14264,N_13977,N_13783);
xnor U14265 (N_14265,N_13650,N_13556);
nand U14266 (N_14266,N_13827,N_13677);
or U14267 (N_14267,N_13505,N_13921);
nor U14268 (N_14268,N_13830,N_13940);
and U14269 (N_14269,N_13925,N_13895);
nor U14270 (N_14270,N_13741,N_13673);
nor U14271 (N_14271,N_13819,N_13516);
and U14272 (N_14272,N_13680,N_13613);
and U14273 (N_14273,N_13829,N_13888);
xor U14274 (N_14274,N_13568,N_13705);
nand U14275 (N_14275,N_13807,N_13630);
xor U14276 (N_14276,N_13912,N_13702);
xor U14277 (N_14277,N_13933,N_13592);
nand U14278 (N_14278,N_13758,N_13507);
and U14279 (N_14279,N_13524,N_13565);
or U14280 (N_14280,N_13819,N_13945);
and U14281 (N_14281,N_13844,N_13620);
nand U14282 (N_14282,N_13736,N_13944);
and U14283 (N_14283,N_13704,N_13685);
and U14284 (N_14284,N_13780,N_13717);
xnor U14285 (N_14285,N_13992,N_13913);
or U14286 (N_14286,N_13634,N_13617);
and U14287 (N_14287,N_13747,N_13835);
xor U14288 (N_14288,N_13515,N_13541);
nor U14289 (N_14289,N_13694,N_13946);
xor U14290 (N_14290,N_13944,N_13924);
nor U14291 (N_14291,N_13675,N_13612);
or U14292 (N_14292,N_13739,N_13989);
and U14293 (N_14293,N_13838,N_13743);
and U14294 (N_14294,N_13643,N_13765);
nand U14295 (N_14295,N_13978,N_13734);
nand U14296 (N_14296,N_13842,N_13766);
xor U14297 (N_14297,N_13852,N_13954);
nand U14298 (N_14298,N_13909,N_13504);
and U14299 (N_14299,N_13759,N_13523);
nand U14300 (N_14300,N_13807,N_13934);
and U14301 (N_14301,N_13825,N_13641);
nand U14302 (N_14302,N_13853,N_13522);
nand U14303 (N_14303,N_13664,N_13539);
xor U14304 (N_14304,N_13744,N_13914);
and U14305 (N_14305,N_13700,N_13814);
xor U14306 (N_14306,N_13664,N_13792);
and U14307 (N_14307,N_13799,N_13595);
xnor U14308 (N_14308,N_13672,N_13592);
and U14309 (N_14309,N_13928,N_13767);
xor U14310 (N_14310,N_13897,N_13732);
xor U14311 (N_14311,N_13824,N_13913);
and U14312 (N_14312,N_13908,N_13591);
or U14313 (N_14313,N_13715,N_13867);
xor U14314 (N_14314,N_13709,N_13854);
nor U14315 (N_14315,N_13517,N_13709);
nor U14316 (N_14316,N_13789,N_13764);
or U14317 (N_14317,N_13796,N_13727);
or U14318 (N_14318,N_13659,N_13692);
nor U14319 (N_14319,N_13842,N_13874);
and U14320 (N_14320,N_13708,N_13691);
xnor U14321 (N_14321,N_13795,N_13600);
xor U14322 (N_14322,N_13995,N_13998);
or U14323 (N_14323,N_13769,N_13553);
nor U14324 (N_14324,N_13777,N_13846);
and U14325 (N_14325,N_13683,N_13632);
or U14326 (N_14326,N_13844,N_13733);
xor U14327 (N_14327,N_13633,N_13613);
nor U14328 (N_14328,N_13687,N_13783);
nand U14329 (N_14329,N_13845,N_13677);
and U14330 (N_14330,N_13871,N_13652);
nand U14331 (N_14331,N_13993,N_13503);
xor U14332 (N_14332,N_13775,N_13636);
nor U14333 (N_14333,N_13745,N_13810);
xor U14334 (N_14334,N_13598,N_13597);
or U14335 (N_14335,N_13943,N_13632);
and U14336 (N_14336,N_13561,N_13839);
nand U14337 (N_14337,N_13759,N_13654);
nand U14338 (N_14338,N_13941,N_13597);
xor U14339 (N_14339,N_13935,N_13937);
nand U14340 (N_14340,N_13774,N_13965);
nor U14341 (N_14341,N_13992,N_13662);
xnor U14342 (N_14342,N_13962,N_13765);
or U14343 (N_14343,N_13974,N_13708);
xnor U14344 (N_14344,N_13542,N_13582);
xnor U14345 (N_14345,N_13781,N_13627);
nor U14346 (N_14346,N_13864,N_13676);
nand U14347 (N_14347,N_13724,N_13862);
or U14348 (N_14348,N_13517,N_13688);
or U14349 (N_14349,N_13606,N_13520);
nor U14350 (N_14350,N_13594,N_13990);
xor U14351 (N_14351,N_13757,N_13649);
or U14352 (N_14352,N_13713,N_13665);
and U14353 (N_14353,N_13822,N_13962);
nor U14354 (N_14354,N_13548,N_13551);
and U14355 (N_14355,N_13523,N_13514);
nor U14356 (N_14356,N_13656,N_13505);
xnor U14357 (N_14357,N_13896,N_13573);
or U14358 (N_14358,N_13521,N_13863);
and U14359 (N_14359,N_13518,N_13859);
and U14360 (N_14360,N_13594,N_13715);
nor U14361 (N_14361,N_13794,N_13895);
nor U14362 (N_14362,N_13759,N_13704);
nand U14363 (N_14363,N_13570,N_13609);
and U14364 (N_14364,N_13744,N_13540);
and U14365 (N_14365,N_13556,N_13926);
and U14366 (N_14366,N_13793,N_13992);
nand U14367 (N_14367,N_13685,N_13912);
and U14368 (N_14368,N_13821,N_13670);
or U14369 (N_14369,N_13517,N_13648);
or U14370 (N_14370,N_13548,N_13561);
nor U14371 (N_14371,N_13982,N_13871);
and U14372 (N_14372,N_13969,N_13555);
nor U14373 (N_14373,N_13848,N_13932);
nand U14374 (N_14374,N_13553,N_13677);
nand U14375 (N_14375,N_13712,N_13805);
nand U14376 (N_14376,N_13812,N_13818);
or U14377 (N_14377,N_13860,N_13554);
nor U14378 (N_14378,N_13756,N_13960);
or U14379 (N_14379,N_13663,N_13995);
nand U14380 (N_14380,N_13658,N_13530);
and U14381 (N_14381,N_13641,N_13610);
and U14382 (N_14382,N_13634,N_13711);
or U14383 (N_14383,N_13911,N_13975);
nor U14384 (N_14384,N_13770,N_13860);
nor U14385 (N_14385,N_13640,N_13729);
and U14386 (N_14386,N_13893,N_13807);
and U14387 (N_14387,N_13895,N_13926);
or U14388 (N_14388,N_13607,N_13902);
nand U14389 (N_14389,N_13595,N_13528);
nor U14390 (N_14390,N_13573,N_13663);
nor U14391 (N_14391,N_13599,N_13767);
and U14392 (N_14392,N_13752,N_13536);
or U14393 (N_14393,N_13646,N_13915);
nand U14394 (N_14394,N_13956,N_13590);
xor U14395 (N_14395,N_13633,N_13770);
and U14396 (N_14396,N_13694,N_13609);
xor U14397 (N_14397,N_13926,N_13560);
nand U14398 (N_14398,N_13872,N_13666);
or U14399 (N_14399,N_13666,N_13938);
and U14400 (N_14400,N_13579,N_13591);
and U14401 (N_14401,N_13628,N_13551);
nor U14402 (N_14402,N_13558,N_13942);
and U14403 (N_14403,N_13800,N_13947);
or U14404 (N_14404,N_13692,N_13538);
and U14405 (N_14405,N_13846,N_13812);
or U14406 (N_14406,N_13991,N_13597);
nand U14407 (N_14407,N_13752,N_13920);
nand U14408 (N_14408,N_13844,N_13924);
nor U14409 (N_14409,N_13660,N_13600);
nand U14410 (N_14410,N_13882,N_13708);
nand U14411 (N_14411,N_13775,N_13871);
or U14412 (N_14412,N_13962,N_13613);
nand U14413 (N_14413,N_13630,N_13673);
nand U14414 (N_14414,N_13965,N_13973);
nor U14415 (N_14415,N_13827,N_13545);
or U14416 (N_14416,N_13773,N_13847);
and U14417 (N_14417,N_13531,N_13998);
nor U14418 (N_14418,N_13774,N_13520);
or U14419 (N_14419,N_13533,N_13578);
nor U14420 (N_14420,N_13552,N_13522);
or U14421 (N_14421,N_13553,N_13898);
and U14422 (N_14422,N_13736,N_13621);
and U14423 (N_14423,N_13688,N_13942);
nand U14424 (N_14424,N_13749,N_13689);
xnor U14425 (N_14425,N_13963,N_13973);
or U14426 (N_14426,N_13680,N_13656);
and U14427 (N_14427,N_13592,N_13750);
nand U14428 (N_14428,N_13835,N_13843);
or U14429 (N_14429,N_13925,N_13972);
nand U14430 (N_14430,N_13605,N_13737);
nand U14431 (N_14431,N_13866,N_13762);
xnor U14432 (N_14432,N_13955,N_13818);
and U14433 (N_14433,N_13817,N_13658);
nor U14434 (N_14434,N_13801,N_13596);
or U14435 (N_14435,N_13656,N_13688);
nand U14436 (N_14436,N_13727,N_13833);
and U14437 (N_14437,N_13578,N_13736);
nor U14438 (N_14438,N_13944,N_13696);
nor U14439 (N_14439,N_13959,N_13774);
and U14440 (N_14440,N_13797,N_13596);
nor U14441 (N_14441,N_13786,N_13500);
xor U14442 (N_14442,N_13852,N_13749);
nor U14443 (N_14443,N_13725,N_13703);
nor U14444 (N_14444,N_13641,N_13939);
nor U14445 (N_14445,N_13630,N_13706);
and U14446 (N_14446,N_13520,N_13618);
or U14447 (N_14447,N_13833,N_13510);
and U14448 (N_14448,N_13796,N_13704);
nand U14449 (N_14449,N_13637,N_13725);
xnor U14450 (N_14450,N_13997,N_13952);
or U14451 (N_14451,N_13724,N_13579);
nor U14452 (N_14452,N_13587,N_13736);
nand U14453 (N_14453,N_13781,N_13929);
nor U14454 (N_14454,N_13600,N_13793);
nand U14455 (N_14455,N_13983,N_13814);
nand U14456 (N_14456,N_13831,N_13593);
and U14457 (N_14457,N_13511,N_13946);
or U14458 (N_14458,N_13984,N_13972);
or U14459 (N_14459,N_13945,N_13533);
xor U14460 (N_14460,N_13638,N_13910);
and U14461 (N_14461,N_13769,N_13710);
or U14462 (N_14462,N_13955,N_13849);
nand U14463 (N_14463,N_13798,N_13923);
or U14464 (N_14464,N_13653,N_13866);
and U14465 (N_14465,N_13997,N_13880);
or U14466 (N_14466,N_13993,N_13752);
xor U14467 (N_14467,N_13597,N_13837);
and U14468 (N_14468,N_13922,N_13960);
nor U14469 (N_14469,N_13830,N_13796);
and U14470 (N_14470,N_13834,N_13977);
or U14471 (N_14471,N_13851,N_13882);
xor U14472 (N_14472,N_13860,N_13841);
xnor U14473 (N_14473,N_13939,N_13949);
nor U14474 (N_14474,N_13732,N_13871);
and U14475 (N_14475,N_13960,N_13965);
nand U14476 (N_14476,N_13715,N_13559);
nor U14477 (N_14477,N_13535,N_13541);
nor U14478 (N_14478,N_13897,N_13969);
nand U14479 (N_14479,N_13915,N_13739);
or U14480 (N_14480,N_13687,N_13881);
xnor U14481 (N_14481,N_13500,N_13798);
nand U14482 (N_14482,N_13748,N_13830);
nand U14483 (N_14483,N_13564,N_13757);
xnor U14484 (N_14484,N_13798,N_13824);
nor U14485 (N_14485,N_13531,N_13826);
nand U14486 (N_14486,N_13599,N_13557);
and U14487 (N_14487,N_13509,N_13992);
and U14488 (N_14488,N_13967,N_13767);
nand U14489 (N_14489,N_13600,N_13980);
and U14490 (N_14490,N_13874,N_13838);
nor U14491 (N_14491,N_13893,N_13856);
or U14492 (N_14492,N_13655,N_13879);
and U14493 (N_14493,N_13973,N_13909);
xnor U14494 (N_14494,N_13702,N_13836);
or U14495 (N_14495,N_13776,N_13649);
nand U14496 (N_14496,N_13708,N_13697);
nand U14497 (N_14497,N_13994,N_13869);
nor U14498 (N_14498,N_13958,N_13503);
nand U14499 (N_14499,N_13841,N_13685);
nand U14500 (N_14500,N_14191,N_14012);
and U14501 (N_14501,N_14437,N_14404);
xnor U14502 (N_14502,N_14489,N_14438);
nand U14503 (N_14503,N_14253,N_14001);
xor U14504 (N_14504,N_14213,N_14259);
nand U14505 (N_14505,N_14076,N_14083);
and U14506 (N_14506,N_14323,N_14379);
or U14507 (N_14507,N_14337,N_14449);
nand U14508 (N_14508,N_14137,N_14156);
xor U14509 (N_14509,N_14212,N_14096);
xnor U14510 (N_14510,N_14490,N_14055);
or U14511 (N_14511,N_14401,N_14045);
nand U14512 (N_14512,N_14269,N_14183);
or U14513 (N_14513,N_14487,N_14053);
and U14514 (N_14514,N_14427,N_14483);
or U14515 (N_14515,N_14425,N_14226);
nand U14516 (N_14516,N_14312,N_14287);
nor U14517 (N_14517,N_14331,N_14235);
and U14518 (N_14518,N_14221,N_14171);
or U14519 (N_14519,N_14015,N_14162);
xnor U14520 (N_14520,N_14362,N_14336);
and U14521 (N_14521,N_14376,N_14266);
nor U14522 (N_14522,N_14227,N_14219);
or U14523 (N_14523,N_14245,N_14407);
nand U14524 (N_14524,N_14155,N_14298);
nand U14525 (N_14525,N_14163,N_14468);
or U14526 (N_14526,N_14103,N_14014);
or U14527 (N_14527,N_14192,N_14218);
or U14528 (N_14528,N_14327,N_14410);
or U14529 (N_14529,N_14320,N_14193);
and U14530 (N_14530,N_14148,N_14047);
xor U14531 (N_14531,N_14054,N_14088);
nor U14532 (N_14532,N_14247,N_14277);
nand U14533 (N_14533,N_14321,N_14005);
or U14534 (N_14534,N_14081,N_14369);
nand U14535 (N_14535,N_14041,N_14339);
and U14536 (N_14536,N_14236,N_14002);
xnor U14537 (N_14537,N_14290,N_14216);
and U14538 (N_14538,N_14030,N_14286);
xor U14539 (N_14539,N_14318,N_14090);
or U14540 (N_14540,N_14089,N_14328);
and U14541 (N_14541,N_14164,N_14330);
or U14542 (N_14542,N_14201,N_14185);
nand U14543 (N_14543,N_14058,N_14107);
xnor U14544 (N_14544,N_14241,N_14256);
nor U14545 (N_14545,N_14264,N_14310);
nor U14546 (N_14546,N_14324,N_14099);
or U14547 (N_14547,N_14040,N_14249);
or U14548 (N_14548,N_14434,N_14451);
and U14549 (N_14549,N_14319,N_14342);
or U14550 (N_14550,N_14347,N_14203);
and U14551 (N_14551,N_14303,N_14305);
xor U14552 (N_14552,N_14311,N_14016);
or U14553 (N_14553,N_14460,N_14222);
nand U14554 (N_14554,N_14072,N_14220);
nand U14555 (N_14555,N_14032,N_14409);
nor U14556 (N_14556,N_14051,N_14050);
or U14557 (N_14557,N_14144,N_14364);
or U14558 (N_14558,N_14093,N_14413);
xor U14559 (N_14559,N_14448,N_14059);
nand U14560 (N_14560,N_14215,N_14372);
nor U14561 (N_14561,N_14146,N_14273);
xor U14562 (N_14562,N_14013,N_14140);
nand U14563 (N_14563,N_14112,N_14181);
nor U14564 (N_14564,N_14289,N_14262);
nand U14565 (N_14565,N_14452,N_14282);
and U14566 (N_14566,N_14242,N_14458);
or U14567 (N_14567,N_14399,N_14348);
nor U14568 (N_14568,N_14010,N_14354);
nand U14569 (N_14569,N_14422,N_14027);
and U14570 (N_14570,N_14066,N_14465);
nor U14571 (N_14571,N_14154,N_14217);
or U14572 (N_14572,N_14157,N_14393);
xnor U14573 (N_14573,N_14223,N_14430);
and U14574 (N_14574,N_14017,N_14341);
nand U14575 (N_14575,N_14044,N_14447);
nor U14576 (N_14576,N_14145,N_14190);
and U14577 (N_14577,N_14435,N_14138);
and U14578 (N_14578,N_14123,N_14308);
or U14579 (N_14579,N_14060,N_14113);
and U14580 (N_14580,N_14159,N_14023);
nor U14581 (N_14581,N_14075,N_14382);
xnor U14582 (N_14582,N_14065,N_14326);
xor U14583 (N_14583,N_14477,N_14349);
and U14584 (N_14584,N_14120,N_14199);
and U14585 (N_14585,N_14248,N_14028);
or U14586 (N_14586,N_14283,N_14254);
xnor U14587 (N_14587,N_14469,N_14378);
or U14588 (N_14588,N_14400,N_14414);
xor U14589 (N_14589,N_14357,N_14478);
or U14590 (N_14590,N_14296,N_14432);
and U14591 (N_14591,N_14069,N_14431);
nand U14592 (N_14592,N_14472,N_14237);
xnor U14593 (N_14593,N_14428,N_14003);
or U14594 (N_14594,N_14007,N_14068);
nand U14595 (N_14595,N_14109,N_14322);
xor U14596 (N_14596,N_14251,N_14125);
and U14597 (N_14597,N_14272,N_14009);
nand U14598 (N_14598,N_14476,N_14367);
nor U14599 (N_14599,N_14333,N_14474);
xor U14600 (N_14600,N_14317,N_14111);
or U14601 (N_14601,N_14355,N_14240);
xnor U14602 (N_14602,N_14149,N_14124);
nand U14603 (N_14603,N_14134,N_14441);
or U14604 (N_14604,N_14229,N_14356);
and U14605 (N_14605,N_14481,N_14383);
nand U14606 (N_14606,N_14151,N_14482);
nor U14607 (N_14607,N_14291,N_14270);
nand U14608 (N_14608,N_14231,N_14423);
or U14609 (N_14609,N_14126,N_14417);
nor U14610 (N_14610,N_14178,N_14386);
and U14611 (N_14611,N_14029,N_14384);
nand U14612 (N_14612,N_14129,N_14358);
nor U14613 (N_14613,N_14209,N_14280);
or U14614 (N_14614,N_14394,N_14067);
and U14615 (N_14615,N_14132,N_14142);
and U14616 (N_14616,N_14471,N_14117);
nand U14617 (N_14617,N_14118,N_14091);
xor U14618 (N_14618,N_14301,N_14025);
xnor U14619 (N_14619,N_14039,N_14133);
or U14620 (N_14620,N_14211,N_14371);
xnor U14621 (N_14621,N_14411,N_14436);
xor U14622 (N_14622,N_14167,N_14456);
and U14623 (N_14623,N_14388,N_14198);
nor U14624 (N_14624,N_14257,N_14176);
nand U14625 (N_14625,N_14115,N_14492);
xnor U14626 (N_14626,N_14078,N_14292);
nand U14627 (N_14627,N_14228,N_14197);
nand U14628 (N_14628,N_14353,N_14043);
xor U14629 (N_14629,N_14061,N_14244);
nor U14630 (N_14630,N_14480,N_14080);
nor U14631 (N_14631,N_14000,N_14498);
xor U14632 (N_14632,N_14136,N_14499);
nand U14633 (N_14633,N_14359,N_14034);
and U14634 (N_14634,N_14454,N_14079);
or U14635 (N_14635,N_14127,N_14252);
xnor U14636 (N_14636,N_14175,N_14405);
nand U14637 (N_14637,N_14325,N_14275);
nor U14638 (N_14638,N_14214,N_14020);
xnor U14639 (N_14639,N_14035,N_14467);
xor U14640 (N_14640,N_14122,N_14462);
or U14641 (N_14641,N_14334,N_14152);
or U14642 (N_14642,N_14415,N_14189);
and U14643 (N_14643,N_14166,N_14139);
nand U14644 (N_14644,N_14461,N_14094);
and U14645 (N_14645,N_14085,N_14365);
nand U14646 (N_14646,N_14445,N_14375);
and U14647 (N_14647,N_14338,N_14052);
or U14648 (N_14648,N_14457,N_14443);
and U14649 (N_14649,N_14486,N_14316);
nor U14650 (N_14650,N_14306,N_14466);
nor U14651 (N_14651,N_14426,N_14293);
or U14652 (N_14652,N_14300,N_14455);
nor U14653 (N_14653,N_14173,N_14370);
and U14654 (N_14654,N_14108,N_14104);
or U14655 (N_14655,N_14082,N_14150);
nor U14656 (N_14656,N_14281,N_14470);
or U14657 (N_14657,N_14402,N_14497);
nand U14658 (N_14658,N_14390,N_14473);
xor U14659 (N_14659,N_14086,N_14442);
nand U14660 (N_14660,N_14267,N_14019);
and U14661 (N_14661,N_14479,N_14391);
and U14662 (N_14662,N_14011,N_14395);
nand U14663 (N_14663,N_14366,N_14006);
nor U14664 (N_14664,N_14194,N_14130);
xnor U14665 (N_14665,N_14314,N_14179);
xnor U14666 (N_14666,N_14206,N_14440);
xor U14667 (N_14667,N_14098,N_14343);
and U14668 (N_14668,N_14250,N_14377);
or U14669 (N_14669,N_14315,N_14444);
and U14670 (N_14670,N_14351,N_14260);
nand U14671 (N_14671,N_14463,N_14459);
xor U14672 (N_14672,N_14268,N_14346);
and U14673 (N_14673,N_14294,N_14288);
and U14674 (N_14674,N_14380,N_14488);
or U14675 (N_14675,N_14121,N_14381);
or U14676 (N_14676,N_14169,N_14070);
xnor U14677 (N_14677,N_14284,N_14225);
and U14678 (N_14678,N_14429,N_14398);
xnor U14679 (N_14679,N_14036,N_14485);
and U14680 (N_14680,N_14018,N_14106);
and U14681 (N_14681,N_14309,N_14446);
nand U14682 (N_14682,N_14038,N_14397);
and U14683 (N_14683,N_14453,N_14238);
nor U14684 (N_14684,N_14495,N_14184);
nor U14685 (N_14685,N_14101,N_14265);
nor U14686 (N_14686,N_14464,N_14233);
nor U14687 (N_14687,N_14373,N_14484);
or U14688 (N_14688,N_14494,N_14307);
and U14689 (N_14689,N_14196,N_14403);
nand U14690 (N_14690,N_14056,N_14165);
or U14691 (N_14691,N_14433,N_14074);
xnor U14692 (N_14692,N_14439,N_14182);
and U14693 (N_14693,N_14204,N_14493);
nand U14694 (N_14694,N_14285,N_14042);
nand U14695 (N_14695,N_14361,N_14340);
and U14696 (N_14696,N_14412,N_14246);
nand U14697 (N_14697,N_14186,N_14297);
or U14698 (N_14698,N_14232,N_14363);
xor U14699 (N_14699,N_14119,N_14385);
nor U14700 (N_14700,N_14295,N_14202);
and U14701 (N_14701,N_14424,N_14160);
xnor U14702 (N_14702,N_14224,N_14174);
nor U14703 (N_14703,N_14491,N_14350);
nor U14704 (N_14704,N_14057,N_14168);
and U14705 (N_14705,N_14374,N_14332);
or U14706 (N_14706,N_14304,N_14102);
nand U14707 (N_14707,N_14177,N_14063);
and U14708 (N_14708,N_14161,N_14406);
and U14709 (N_14709,N_14004,N_14274);
or U14710 (N_14710,N_14263,N_14026);
nand U14711 (N_14711,N_14210,N_14450);
xor U14712 (N_14712,N_14077,N_14258);
and U14713 (N_14713,N_14131,N_14008);
or U14714 (N_14714,N_14170,N_14416);
nand U14715 (N_14715,N_14147,N_14408);
and U14716 (N_14716,N_14031,N_14116);
and U14717 (N_14717,N_14135,N_14352);
nor U14718 (N_14718,N_14114,N_14392);
nor U14719 (N_14719,N_14087,N_14188);
xnor U14720 (N_14720,N_14313,N_14208);
nor U14721 (N_14721,N_14048,N_14143);
nand U14722 (N_14722,N_14345,N_14128);
nor U14723 (N_14723,N_14421,N_14100);
and U14724 (N_14724,N_14071,N_14299);
and U14725 (N_14725,N_14475,N_14097);
nand U14726 (N_14726,N_14368,N_14046);
nor U14727 (N_14727,N_14024,N_14239);
or U14728 (N_14728,N_14073,N_14092);
and U14729 (N_14729,N_14195,N_14271);
nand U14730 (N_14730,N_14105,N_14172);
nand U14731 (N_14731,N_14255,N_14084);
nor U14732 (N_14732,N_14180,N_14279);
nor U14733 (N_14733,N_14153,N_14064);
or U14734 (N_14734,N_14207,N_14496);
or U14735 (N_14735,N_14062,N_14389);
nor U14736 (N_14736,N_14335,N_14095);
or U14737 (N_14737,N_14200,N_14205);
nand U14738 (N_14738,N_14243,N_14033);
nand U14739 (N_14739,N_14110,N_14037);
and U14740 (N_14740,N_14187,N_14396);
nor U14741 (N_14741,N_14344,N_14158);
nand U14742 (N_14742,N_14419,N_14141);
nand U14743 (N_14743,N_14234,N_14230);
and U14744 (N_14744,N_14302,N_14021);
nand U14745 (N_14745,N_14276,N_14049);
xor U14746 (N_14746,N_14360,N_14022);
nor U14747 (N_14747,N_14420,N_14387);
and U14748 (N_14748,N_14418,N_14278);
nor U14749 (N_14749,N_14261,N_14329);
and U14750 (N_14750,N_14287,N_14460);
xor U14751 (N_14751,N_14267,N_14031);
nand U14752 (N_14752,N_14096,N_14377);
nor U14753 (N_14753,N_14062,N_14006);
nand U14754 (N_14754,N_14396,N_14181);
nand U14755 (N_14755,N_14249,N_14306);
nor U14756 (N_14756,N_14047,N_14471);
and U14757 (N_14757,N_14491,N_14098);
nor U14758 (N_14758,N_14037,N_14050);
nand U14759 (N_14759,N_14427,N_14317);
xnor U14760 (N_14760,N_14051,N_14092);
nand U14761 (N_14761,N_14375,N_14065);
or U14762 (N_14762,N_14356,N_14313);
or U14763 (N_14763,N_14308,N_14327);
nor U14764 (N_14764,N_14307,N_14139);
and U14765 (N_14765,N_14180,N_14338);
xor U14766 (N_14766,N_14150,N_14384);
nor U14767 (N_14767,N_14252,N_14394);
nor U14768 (N_14768,N_14093,N_14454);
nor U14769 (N_14769,N_14253,N_14189);
xor U14770 (N_14770,N_14253,N_14225);
nor U14771 (N_14771,N_14412,N_14041);
nor U14772 (N_14772,N_14300,N_14433);
xnor U14773 (N_14773,N_14097,N_14238);
and U14774 (N_14774,N_14143,N_14137);
or U14775 (N_14775,N_14036,N_14467);
nand U14776 (N_14776,N_14318,N_14093);
xnor U14777 (N_14777,N_14393,N_14458);
nand U14778 (N_14778,N_14226,N_14170);
nor U14779 (N_14779,N_14129,N_14222);
nor U14780 (N_14780,N_14030,N_14363);
nand U14781 (N_14781,N_14220,N_14199);
nor U14782 (N_14782,N_14138,N_14465);
xor U14783 (N_14783,N_14234,N_14324);
or U14784 (N_14784,N_14034,N_14479);
xnor U14785 (N_14785,N_14244,N_14421);
and U14786 (N_14786,N_14483,N_14224);
nor U14787 (N_14787,N_14103,N_14224);
and U14788 (N_14788,N_14089,N_14209);
and U14789 (N_14789,N_14486,N_14032);
and U14790 (N_14790,N_14072,N_14122);
nor U14791 (N_14791,N_14258,N_14030);
xnor U14792 (N_14792,N_14133,N_14119);
and U14793 (N_14793,N_14238,N_14062);
and U14794 (N_14794,N_14295,N_14319);
nor U14795 (N_14795,N_14002,N_14305);
or U14796 (N_14796,N_14196,N_14238);
nor U14797 (N_14797,N_14376,N_14148);
and U14798 (N_14798,N_14383,N_14399);
or U14799 (N_14799,N_14188,N_14015);
nor U14800 (N_14800,N_14391,N_14154);
and U14801 (N_14801,N_14482,N_14181);
and U14802 (N_14802,N_14225,N_14450);
nand U14803 (N_14803,N_14125,N_14262);
or U14804 (N_14804,N_14496,N_14348);
nor U14805 (N_14805,N_14345,N_14354);
and U14806 (N_14806,N_14452,N_14279);
or U14807 (N_14807,N_14010,N_14272);
nand U14808 (N_14808,N_14014,N_14027);
or U14809 (N_14809,N_14498,N_14419);
or U14810 (N_14810,N_14017,N_14468);
and U14811 (N_14811,N_14331,N_14027);
xnor U14812 (N_14812,N_14101,N_14272);
or U14813 (N_14813,N_14049,N_14489);
nor U14814 (N_14814,N_14424,N_14292);
xnor U14815 (N_14815,N_14414,N_14433);
or U14816 (N_14816,N_14333,N_14003);
nand U14817 (N_14817,N_14471,N_14141);
or U14818 (N_14818,N_14275,N_14411);
or U14819 (N_14819,N_14286,N_14106);
nor U14820 (N_14820,N_14306,N_14027);
xnor U14821 (N_14821,N_14251,N_14014);
and U14822 (N_14822,N_14205,N_14105);
and U14823 (N_14823,N_14306,N_14317);
nor U14824 (N_14824,N_14008,N_14321);
xnor U14825 (N_14825,N_14105,N_14126);
xor U14826 (N_14826,N_14410,N_14243);
xnor U14827 (N_14827,N_14334,N_14109);
xor U14828 (N_14828,N_14115,N_14219);
or U14829 (N_14829,N_14299,N_14432);
and U14830 (N_14830,N_14270,N_14093);
or U14831 (N_14831,N_14219,N_14345);
and U14832 (N_14832,N_14494,N_14349);
nand U14833 (N_14833,N_14268,N_14020);
xnor U14834 (N_14834,N_14360,N_14183);
and U14835 (N_14835,N_14291,N_14170);
xnor U14836 (N_14836,N_14024,N_14470);
nor U14837 (N_14837,N_14231,N_14480);
nor U14838 (N_14838,N_14211,N_14357);
xor U14839 (N_14839,N_14259,N_14092);
nor U14840 (N_14840,N_14219,N_14425);
or U14841 (N_14841,N_14093,N_14259);
nand U14842 (N_14842,N_14036,N_14186);
xor U14843 (N_14843,N_14450,N_14424);
nor U14844 (N_14844,N_14379,N_14471);
or U14845 (N_14845,N_14088,N_14444);
or U14846 (N_14846,N_14174,N_14445);
xnor U14847 (N_14847,N_14261,N_14277);
or U14848 (N_14848,N_14033,N_14055);
nor U14849 (N_14849,N_14176,N_14086);
nand U14850 (N_14850,N_14056,N_14388);
or U14851 (N_14851,N_14487,N_14265);
nor U14852 (N_14852,N_14370,N_14211);
or U14853 (N_14853,N_14005,N_14334);
nand U14854 (N_14854,N_14256,N_14000);
or U14855 (N_14855,N_14346,N_14210);
nor U14856 (N_14856,N_14333,N_14117);
xnor U14857 (N_14857,N_14054,N_14399);
or U14858 (N_14858,N_14399,N_14019);
or U14859 (N_14859,N_14026,N_14482);
xor U14860 (N_14860,N_14096,N_14178);
and U14861 (N_14861,N_14100,N_14431);
xnor U14862 (N_14862,N_14045,N_14111);
nand U14863 (N_14863,N_14013,N_14463);
nor U14864 (N_14864,N_14018,N_14045);
nor U14865 (N_14865,N_14093,N_14103);
and U14866 (N_14866,N_14061,N_14199);
nor U14867 (N_14867,N_14370,N_14014);
nand U14868 (N_14868,N_14210,N_14165);
nand U14869 (N_14869,N_14037,N_14023);
or U14870 (N_14870,N_14320,N_14061);
or U14871 (N_14871,N_14022,N_14322);
nor U14872 (N_14872,N_14082,N_14157);
and U14873 (N_14873,N_14212,N_14451);
xnor U14874 (N_14874,N_14214,N_14287);
or U14875 (N_14875,N_14262,N_14467);
or U14876 (N_14876,N_14054,N_14368);
nand U14877 (N_14877,N_14126,N_14185);
nand U14878 (N_14878,N_14308,N_14105);
and U14879 (N_14879,N_14195,N_14404);
nor U14880 (N_14880,N_14076,N_14139);
nand U14881 (N_14881,N_14250,N_14314);
nor U14882 (N_14882,N_14335,N_14132);
nand U14883 (N_14883,N_14272,N_14241);
or U14884 (N_14884,N_14235,N_14212);
nand U14885 (N_14885,N_14277,N_14008);
nand U14886 (N_14886,N_14357,N_14041);
nor U14887 (N_14887,N_14446,N_14020);
nand U14888 (N_14888,N_14007,N_14423);
nand U14889 (N_14889,N_14498,N_14216);
nand U14890 (N_14890,N_14197,N_14246);
nor U14891 (N_14891,N_14416,N_14018);
nor U14892 (N_14892,N_14057,N_14439);
xor U14893 (N_14893,N_14222,N_14491);
and U14894 (N_14894,N_14133,N_14495);
nand U14895 (N_14895,N_14204,N_14194);
and U14896 (N_14896,N_14328,N_14447);
or U14897 (N_14897,N_14034,N_14074);
nor U14898 (N_14898,N_14147,N_14238);
and U14899 (N_14899,N_14280,N_14157);
xnor U14900 (N_14900,N_14126,N_14217);
or U14901 (N_14901,N_14241,N_14487);
and U14902 (N_14902,N_14426,N_14048);
xor U14903 (N_14903,N_14287,N_14151);
nand U14904 (N_14904,N_14065,N_14077);
xor U14905 (N_14905,N_14216,N_14052);
or U14906 (N_14906,N_14009,N_14042);
xnor U14907 (N_14907,N_14389,N_14473);
or U14908 (N_14908,N_14111,N_14007);
or U14909 (N_14909,N_14011,N_14251);
nor U14910 (N_14910,N_14358,N_14245);
nor U14911 (N_14911,N_14270,N_14280);
xnor U14912 (N_14912,N_14493,N_14213);
xnor U14913 (N_14913,N_14204,N_14403);
or U14914 (N_14914,N_14089,N_14466);
nor U14915 (N_14915,N_14387,N_14498);
nand U14916 (N_14916,N_14070,N_14459);
or U14917 (N_14917,N_14185,N_14211);
nor U14918 (N_14918,N_14192,N_14134);
xor U14919 (N_14919,N_14053,N_14438);
xnor U14920 (N_14920,N_14458,N_14499);
xor U14921 (N_14921,N_14465,N_14083);
and U14922 (N_14922,N_14036,N_14060);
xnor U14923 (N_14923,N_14196,N_14483);
or U14924 (N_14924,N_14056,N_14235);
or U14925 (N_14925,N_14266,N_14370);
nor U14926 (N_14926,N_14173,N_14413);
xor U14927 (N_14927,N_14176,N_14386);
nand U14928 (N_14928,N_14139,N_14083);
or U14929 (N_14929,N_14328,N_14472);
and U14930 (N_14930,N_14161,N_14003);
or U14931 (N_14931,N_14284,N_14280);
or U14932 (N_14932,N_14154,N_14411);
and U14933 (N_14933,N_14052,N_14483);
xnor U14934 (N_14934,N_14012,N_14408);
nor U14935 (N_14935,N_14252,N_14192);
nor U14936 (N_14936,N_14093,N_14417);
and U14937 (N_14937,N_14094,N_14151);
and U14938 (N_14938,N_14274,N_14418);
nor U14939 (N_14939,N_14003,N_14120);
nor U14940 (N_14940,N_14200,N_14040);
nand U14941 (N_14941,N_14012,N_14134);
xnor U14942 (N_14942,N_14428,N_14304);
and U14943 (N_14943,N_14267,N_14098);
and U14944 (N_14944,N_14035,N_14351);
nor U14945 (N_14945,N_14347,N_14496);
or U14946 (N_14946,N_14047,N_14063);
nand U14947 (N_14947,N_14374,N_14067);
nor U14948 (N_14948,N_14291,N_14383);
nor U14949 (N_14949,N_14387,N_14202);
nand U14950 (N_14950,N_14077,N_14234);
or U14951 (N_14951,N_14144,N_14150);
and U14952 (N_14952,N_14151,N_14000);
xor U14953 (N_14953,N_14444,N_14250);
xnor U14954 (N_14954,N_14272,N_14268);
and U14955 (N_14955,N_14230,N_14312);
nand U14956 (N_14956,N_14161,N_14239);
and U14957 (N_14957,N_14491,N_14252);
and U14958 (N_14958,N_14190,N_14034);
and U14959 (N_14959,N_14427,N_14444);
nand U14960 (N_14960,N_14051,N_14289);
or U14961 (N_14961,N_14315,N_14077);
xor U14962 (N_14962,N_14067,N_14312);
nand U14963 (N_14963,N_14111,N_14051);
xor U14964 (N_14964,N_14287,N_14163);
and U14965 (N_14965,N_14401,N_14003);
nor U14966 (N_14966,N_14210,N_14124);
nand U14967 (N_14967,N_14218,N_14361);
or U14968 (N_14968,N_14187,N_14094);
xnor U14969 (N_14969,N_14069,N_14338);
nor U14970 (N_14970,N_14236,N_14062);
nor U14971 (N_14971,N_14189,N_14029);
and U14972 (N_14972,N_14467,N_14248);
nand U14973 (N_14973,N_14352,N_14177);
nand U14974 (N_14974,N_14068,N_14061);
xor U14975 (N_14975,N_14118,N_14125);
nand U14976 (N_14976,N_14085,N_14473);
and U14977 (N_14977,N_14400,N_14218);
nand U14978 (N_14978,N_14027,N_14262);
xor U14979 (N_14979,N_14254,N_14440);
or U14980 (N_14980,N_14246,N_14364);
or U14981 (N_14981,N_14355,N_14310);
and U14982 (N_14982,N_14163,N_14153);
xnor U14983 (N_14983,N_14451,N_14175);
xor U14984 (N_14984,N_14111,N_14307);
and U14985 (N_14985,N_14389,N_14237);
and U14986 (N_14986,N_14348,N_14408);
nor U14987 (N_14987,N_14087,N_14297);
and U14988 (N_14988,N_14295,N_14149);
xnor U14989 (N_14989,N_14102,N_14429);
or U14990 (N_14990,N_14307,N_14154);
and U14991 (N_14991,N_14199,N_14126);
nand U14992 (N_14992,N_14109,N_14257);
nor U14993 (N_14993,N_14201,N_14486);
nor U14994 (N_14994,N_14219,N_14046);
nand U14995 (N_14995,N_14008,N_14211);
nor U14996 (N_14996,N_14134,N_14251);
xor U14997 (N_14997,N_14485,N_14117);
nor U14998 (N_14998,N_14057,N_14142);
nand U14999 (N_14999,N_14265,N_14112);
xnor UO_0 (O_0,N_14568,N_14978);
xor UO_1 (O_1,N_14667,N_14567);
nor UO_2 (O_2,N_14949,N_14767);
xor UO_3 (O_3,N_14985,N_14589);
xnor UO_4 (O_4,N_14757,N_14513);
nand UO_5 (O_5,N_14634,N_14947);
nor UO_6 (O_6,N_14695,N_14810);
and UO_7 (O_7,N_14710,N_14764);
xor UO_8 (O_8,N_14912,N_14822);
nor UO_9 (O_9,N_14701,N_14597);
xor UO_10 (O_10,N_14739,N_14966);
xor UO_11 (O_11,N_14833,N_14694);
nor UO_12 (O_12,N_14962,N_14829);
nor UO_13 (O_13,N_14877,N_14609);
and UO_14 (O_14,N_14522,N_14570);
xnor UO_15 (O_15,N_14948,N_14685);
or UO_16 (O_16,N_14569,N_14809);
xor UO_17 (O_17,N_14578,N_14774);
or UO_18 (O_18,N_14624,N_14780);
nand UO_19 (O_19,N_14890,N_14608);
or UO_20 (O_20,N_14705,N_14857);
xnor UO_21 (O_21,N_14687,N_14721);
nor UO_22 (O_22,N_14799,N_14737);
nand UO_23 (O_23,N_14808,N_14841);
or UO_24 (O_24,N_14756,N_14700);
nand UO_25 (O_25,N_14750,N_14885);
or UO_26 (O_26,N_14862,N_14738);
or UO_27 (O_27,N_14731,N_14903);
or UO_28 (O_28,N_14743,N_14664);
nor UO_29 (O_29,N_14753,N_14509);
xor UO_30 (O_30,N_14768,N_14538);
nand UO_31 (O_31,N_14963,N_14927);
or UO_32 (O_32,N_14717,N_14755);
and UO_33 (O_33,N_14916,N_14747);
or UO_34 (O_34,N_14576,N_14956);
xnor UO_35 (O_35,N_14742,N_14734);
nor UO_36 (O_36,N_14842,N_14791);
and UO_37 (O_37,N_14584,N_14587);
nor UO_38 (O_38,N_14713,N_14585);
or UO_39 (O_39,N_14543,N_14815);
or UO_40 (O_40,N_14817,N_14825);
or UO_41 (O_41,N_14663,N_14970);
xor UO_42 (O_42,N_14577,N_14586);
or UO_43 (O_43,N_14725,N_14816);
and UO_44 (O_44,N_14804,N_14910);
or UO_45 (O_45,N_14714,N_14891);
nor UO_46 (O_46,N_14630,N_14800);
or UO_47 (O_47,N_14836,N_14880);
and UO_48 (O_48,N_14666,N_14790);
or UO_49 (O_49,N_14937,N_14660);
nor UO_50 (O_50,N_14573,N_14803);
nor UO_51 (O_51,N_14698,N_14802);
nor UO_52 (O_52,N_14986,N_14989);
or UO_53 (O_53,N_14792,N_14559);
nand UO_54 (O_54,N_14508,N_14621);
or UO_55 (O_55,N_14794,N_14869);
xor UO_56 (O_56,N_14652,N_14548);
nor UO_57 (O_57,N_14574,N_14661);
xnor UO_58 (O_58,N_14872,N_14563);
nand UO_59 (O_59,N_14723,N_14798);
or UO_60 (O_60,N_14535,N_14580);
xor UO_61 (O_61,N_14888,N_14846);
nor UO_62 (O_62,N_14754,N_14752);
or UO_63 (O_63,N_14882,N_14680);
nor UO_64 (O_64,N_14840,N_14579);
and UO_65 (O_65,N_14997,N_14759);
or UO_66 (O_66,N_14517,N_14765);
nor UO_67 (O_67,N_14730,N_14635);
nor UO_68 (O_68,N_14532,N_14541);
nor UO_69 (O_69,N_14893,N_14636);
nand UO_70 (O_70,N_14950,N_14847);
xor UO_71 (O_71,N_14732,N_14902);
nor UO_72 (O_72,N_14940,N_14853);
nand UO_73 (O_73,N_14644,N_14684);
nand UO_74 (O_74,N_14672,N_14646);
xor UO_75 (O_75,N_14565,N_14600);
xor UO_76 (O_76,N_14631,N_14931);
nand UO_77 (O_77,N_14760,N_14834);
xor UO_78 (O_78,N_14605,N_14826);
xor UO_79 (O_79,N_14859,N_14995);
nand UO_80 (O_80,N_14536,N_14921);
and UO_81 (O_81,N_14554,N_14715);
or UO_82 (O_82,N_14861,N_14524);
nand UO_83 (O_83,N_14789,N_14654);
nand UO_84 (O_84,N_14828,N_14892);
xor UO_85 (O_85,N_14736,N_14958);
xor UO_86 (O_86,N_14788,N_14643);
nor UO_87 (O_87,N_14819,N_14926);
nor UO_88 (O_88,N_14674,N_14657);
nand UO_89 (O_89,N_14653,N_14607);
and UO_90 (O_90,N_14735,N_14914);
or UO_91 (O_91,N_14516,N_14545);
or UO_92 (O_92,N_14603,N_14992);
and UO_93 (O_93,N_14843,N_14782);
nand UO_94 (O_94,N_14557,N_14951);
and UO_95 (O_95,N_14677,N_14542);
xor UO_96 (O_96,N_14669,N_14974);
nor UO_97 (O_97,N_14683,N_14983);
nand UO_98 (O_98,N_14620,N_14855);
xnor UO_99 (O_99,N_14614,N_14924);
or UO_100 (O_100,N_14581,N_14839);
or UO_101 (O_101,N_14783,N_14566);
nand UO_102 (O_102,N_14886,N_14727);
nor UO_103 (O_103,N_14645,N_14813);
nor UO_104 (O_104,N_14728,N_14709);
or UO_105 (O_105,N_14628,N_14518);
and UO_106 (O_106,N_14604,N_14812);
nor UO_107 (O_107,N_14500,N_14741);
nor UO_108 (O_108,N_14900,N_14638);
or UO_109 (O_109,N_14823,N_14712);
or UO_110 (O_110,N_14529,N_14520);
nor UO_111 (O_111,N_14575,N_14606);
or UO_112 (O_112,N_14533,N_14611);
nor UO_113 (O_113,N_14501,N_14623);
nand UO_114 (O_114,N_14671,N_14719);
nor UO_115 (O_115,N_14686,N_14656);
xor UO_116 (O_116,N_14934,N_14873);
xnor UO_117 (O_117,N_14746,N_14758);
nor UO_118 (O_118,N_14771,N_14786);
xnor UO_119 (O_119,N_14688,N_14954);
xnor UO_120 (O_120,N_14655,N_14851);
nor UO_121 (O_121,N_14519,N_14773);
xnor UO_122 (O_122,N_14964,N_14689);
xnor UO_123 (O_123,N_14633,N_14864);
and UO_124 (O_124,N_14599,N_14503);
nand UO_125 (O_125,N_14530,N_14965);
and UO_126 (O_126,N_14512,N_14820);
xnor UO_127 (O_127,N_14668,N_14561);
or UO_128 (O_128,N_14918,N_14720);
nor UO_129 (O_129,N_14676,N_14592);
and UO_130 (O_130,N_14973,N_14593);
nor UO_131 (O_131,N_14544,N_14733);
nand UO_132 (O_132,N_14722,N_14955);
or UO_133 (O_133,N_14928,N_14960);
nand UO_134 (O_134,N_14762,N_14953);
and UO_135 (O_135,N_14572,N_14785);
nand UO_136 (O_136,N_14551,N_14944);
nand UO_137 (O_137,N_14935,N_14941);
nor UO_138 (O_138,N_14514,N_14506);
and UO_139 (O_139,N_14881,N_14675);
and UO_140 (O_140,N_14521,N_14899);
nand UO_141 (O_141,N_14933,N_14549);
or UO_142 (O_142,N_14547,N_14852);
xor UO_143 (O_143,N_14523,N_14854);
nor UO_144 (O_144,N_14740,N_14590);
nand UO_145 (O_145,N_14844,N_14837);
nor UO_146 (O_146,N_14612,N_14831);
nand UO_147 (O_147,N_14601,N_14795);
xnor UO_148 (O_148,N_14845,N_14784);
xor UO_149 (O_149,N_14699,N_14748);
nand UO_150 (O_150,N_14832,N_14778);
nor UO_151 (O_151,N_14678,N_14874);
nor UO_152 (O_152,N_14796,N_14534);
and UO_153 (O_153,N_14776,N_14648);
and UO_154 (O_154,N_14860,N_14507);
nor UO_155 (O_155,N_14595,N_14868);
xnor UO_156 (O_156,N_14887,N_14560);
or UO_157 (O_157,N_14856,N_14658);
and UO_158 (O_158,N_14979,N_14641);
xor UO_159 (O_159,N_14805,N_14649);
nand UO_160 (O_160,N_14904,N_14761);
nand UO_161 (O_161,N_14775,N_14811);
nor UO_162 (O_162,N_14878,N_14884);
and UO_163 (O_163,N_14537,N_14711);
xnor UO_164 (O_164,N_14702,N_14932);
nor UO_165 (O_165,N_14998,N_14591);
xnor UO_166 (O_166,N_14691,N_14894);
nand UO_167 (O_167,N_14703,N_14527);
and UO_168 (O_168,N_14779,N_14708);
and UO_169 (O_169,N_14824,N_14555);
nor UO_170 (O_170,N_14562,N_14911);
xor UO_171 (O_171,N_14629,N_14959);
or UO_172 (O_172,N_14982,N_14745);
and UO_173 (O_173,N_14632,N_14571);
nor UO_174 (O_174,N_14769,N_14618);
or UO_175 (O_175,N_14639,N_14787);
and UO_176 (O_176,N_14697,N_14777);
nor UO_177 (O_177,N_14984,N_14505);
nand UO_178 (O_178,N_14640,N_14670);
and UO_179 (O_179,N_14981,N_14602);
or UO_180 (O_180,N_14943,N_14692);
and UO_181 (O_181,N_14976,N_14550);
xnor UO_182 (O_182,N_14716,N_14946);
and UO_183 (O_183,N_14724,N_14619);
and UO_184 (O_184,N_14510,N_14922);
and UO_185 (O_185,N_14896,N_14617);
nand UO_186 (O_186,N_14763,N_14920);
nor UO_187 (O_187,N_14865,N_14801);
nor UO_188 (O_188,N_14991,N_14980);
xnor UO_189 (O_189,N_14988,N_14729);
xnor UO_190 (O_190,N_14969,N_14908);
nand UO_191 (O_191,N_14807,N_14511);
nand UO_192 (O_192,N_14679,N_14744);
xor UO_193 (O_193,N_14525,N_14594);
and UO_194 (O_194,N_14539,N_14961);
and UO_195 (O_195,N_14662,N_14936);
or UO_196 (O_196,N_14704,N_14673);
nand UO_197 (O_197,N_14564,N_14651);
xnor UO_198 (O_198,N_14830,N_14552);
nor UO_199 (O_199,N_14770,N_14863);
and UO_200 (O_200,N_14528,N_14693);
and UO_201 (O_201,N_14682,N_14526);
and UO_202 (O_202,N_14766,N_14626);
nor UO_203 (O_203,N_14919,N_14977);
nand UO_204 (O_204,N_14987,N_14850);
nand UO_205 (O_205,N_14647,N_14690);
and UO_206 (O_206,N_14866,N_14909);
and UO_207 (O_207,N_14913,N_14515);
nor UO_208 (O_208,N_14967,N_14616);
nand UO_209 (O_209,N_14917,N_14999);
or UO_210 (O_210,N_14504,N_14659);
and UO_211 (O_211,N_14625,N_14797);
and UO_212 (O_212,N_14994,N_14827);
nand UO_213 (O_213,N_14906,N_14696);
and UO_214 (O_214,N_14772,N_14793);
or UO_215 (O_215,N_14818,N_14583);
or UO_216 (O_216,N_14939,N_14971);
nor UO_217 (O_217,N_14706,N_14867);
xnor UO_218 (O_218,N_14895,N_14875);
nor UO_219 (O_219,N_14749,N_14613);
xor UO_220 (O_220,N_14883,N_14642);
and UO_221 (O_221,N_14622,N_14929);
xor UO_222 (O_222,N_14650,N_14938);
or UO_223 (O_223,N_14871,N_14821);
or UO_224 (O_224,N_14915,N_14540);
and UO_225 (O_225,N_14781,N_14901);
xnor UO_226 (O_226,N_14957,N_14870);
or UO_227 (O_227,N_14598,N_14972);
or UO_228 (O_228,N_14558,N_14996);
xnor UO_229 (O_229,N_14848,N_14907);
nand UO_230 (O_230,N_14993,N_14531);
xor UO_231 (O_231,N_14588,N_14968);
or UO_232 (O_232,N_14849,N_14546);
nand UO_233 (O_233,N_14814,N_14726);
and UO_234 (O_234,N_14751,N_14923);
or UO_235 (O_235,N_14707,N_14615);
or UO_236 (O_236,N_14665,N_14942);
nor UO_237 (O_237,N_14838,N_14553);
xnor UO_238 (O_238,N_14610,N_14627);
and UO_239 (O_239,N_14990,N_14502);
nand UO_240 (O_240,N_14898,N_14582);
or UO_241 (O_241,N_14681,N_14945);
nand UO_242 (O_242,N_14556,N_14718);
nand UO_243 (O_243,N_14975,N_14637);
or UO_244 (O_244,N_14876,N_14925);
nand UO_245 (O_245,N_14858,N_14905);
xnor UO_246 (O_246,N_14879,N_14897);
and UO_247 (O_247,N_14930,N_14952);
or UO_248 (O_248,N_14596,N_14889);
nor UO_249 (O_249,N_14835,N_14806);
xor UO_250 (O_250,N_14976,N_14500);
nor UO_251 (O_251,N_14769,N_14689);
and UO_252 (O_252,N_14718,N_14846);
and UO_253 (O_253,N_14939,N_14647);
nand UO_254 (O_254,N_14545,N_14933);
xor UO_255 (O_255,N_14755,N_14812);
xnor UO_256 (O_256,N_14708,N_14777);
or UO_257 (O_257,N_14801,N_14626);
nor UO_258 (O_258,N_14591,N_14912);
and UO_259 (O_259,N_14723,N_14827);
nand UO_260 (O_260,N_14860,N_14774);
or UO_261 (O_261,N_14846,N_14745);
nor UO_262 (O_262,N_14881,N_14548);
nand UO_263 (O_263,N_14966,N_14680);
or UO_264 (O_264,N_14834,N_14878);
xor UO_265 (O_265,N_14995,N_14886);
nand UO_266 (O_266,N_14591,N_14513);
xor UO_267 (O_267,N_14764,N_14910);
nand UO_268 (O_268,N_14889,N_14748);
xnor UO_269 (O_269,N_14775,N_14641);
nor UO_270 (O_270,N_14830,N_14844);
nand UO_271 (O_271,N_14594,N_14750);
or UO_272 (O_272,N_14802,N_14924);
xor UO_273 (O_273,N_14626,N_14687);
nor UO_274 (O_274,N_14740,N_14791);
and UO_275 (O_275,N_14886,N_14519);
nor UO_276 (O_276,N_14892,N_14781);
xor UO_277 (O_277,N_14681,N_14624);
nand UO_278 (O_278,N_14784,N_14774);
xor UO_279 (O_279,N_14964,N_14610);
nand UO_280 (O_280,N_14890,N_14875);
nand UO_281 (O_281,N_14625,N_14770);
nand UO_282 (O_282,N_14984,N_14780);
nand UO_283 (O_283,N_14938,N_14540);
or UO_284 (O_284,N_14681,N_14850);
nand UO_285 (O_285,N_14937,N_14850);
nand UO_286 (O_286,N_14841,N_14934);
and UO_287 (O_287,N_14778,N_14564);
xnor UO_288 (O_288,N_14792,N_14589);
or UO_289 (O_289,N_14749,N_14821);
xor UO_290 (O_290,N_14571,N_14970);
xnor UO_291 (O_291,N_14807,N_14660);
nand UO_292 (O_292,N_14524,N_14979);
and UO_293 (O_293,N_14670,N_14552);
nand UO_294 (O_294,N_14831,N_14783);
or UO_295 (O_295,N_14883,N_14765);
xnor UO_296 (O_296,N_14689,N_14615);
nor UO_297 (O_297,N_14795,N_14944);
nand UO_298 (O_298,N_14688,N_14836);
and UO_299 (O_299,N_14656,N_14615);
or UO_300 (O_300,N_14894,N_14576);
xor UO_301 (O_301,N_14900,N_14913);
and UO_302 (O_302,N_14977,N_14674);
or UO_303 (O_303,N_14764,N_14666);
nand UO_304 (O_304,N_14656,N_14985);
xnor UO_305 (O_305,N_14970,N_14965);
nor UO_306 (O_306,N_14909,N_14991);
nand UO_307 (O_307,N_14718,N_14611);
nand UO_308 (O_308,N_14701,N_14796);
or UO_309 (O_309,N_14908,N_14759);
nor UO_310 (O_310,N_14803,N_14558);
nand UO_311 (O_311,N_14625,N_14863);
nor UO_312 (O_312,N_14974,N_14757);
xnor UO_313 (O_313,N_14606,N_14833);
or UO_314 (O_314,N_14872,N_14553);
and UO_315 (O_315,N_14773,N_14899);
nand UO_316 (O_316,N_14597,N_14846);
xnor UO_317 (O_317,N_14659,N_14983);
and UO_318 (O_318,N_14501,N_14827);
nand UO_319 (O_319,N_14622,N_14714);
nor UO_320 (O_320,N_14705,N_14603);
xor UO_321 (O_321,N_14578,N_14541);
nor UO_322 (O_322,N_14633,N_14793);
or UO_323 (O_323,N_14529,N_14865);
nor UO_324 (O_324,N_14656,N_14886);
nand UO_325 (O_325,N_14541,N_14696);
nor UO_326 (O_326,N_14853,N_14627);
nor UO_327 (O_327,N_14595,N_14814);
nor UO_328 (O_328,N_14914,N_14923);
and UO_329 (O_329,N_14936,N_14949);
nor UO_330 (O_330,N_14820,N_14507);
and UO_331 (O_331,N_14651,N_14951);
nor UO_332 (O_332,N_14919,N_14933);
nand UO_333 (O_333,N_14637,N_14544);
xnor UO_334 (O_334,N_14663,N_14650);
and UO_335 (O_335,N_14849,N_14859);
or UO_336 (O_336,N_14779,N_14500);
nor UO_337 (O_337,N_14858,N_14619);
nand UO_338 (O_338,N_14908,N_14982);
nor UO_339 (O_339,N_14993,N_14661);
nand UO_340 (O_340,N_14723,N_14609);
or UO_341 (O_341,N_14804,N_14605);
or UO_342 (O_342,N_14741,N_14952);
nor UO_343 (O_343,N_14685,N_14719);
and UO_344 (O_344,N_14999,N_14691);
xor UO_345 (O_345,N_14738,N_14666);
xor UO_346 (O_346,N_14647,N_14531);
or UO_347 (O_347,N_14532,N_14663);
or UO_348 (O_348,N_14545,N_14800);
xnor UO_349 (O_349,N_14837,N_14546);
xor UO_350 (O_350,N_14609,N_14990);
nor UO_351 (O_351,N_14800,N_14942);
nand UO_352 (O_352,N_14768,N_14758);
nor UO_353 (O_353,N_14622,N_14793);
nand UO_354 (O_354,N_14671,N_14913);
nor UO_355 (O_355,N_14707,N_14745);
nor UO_356 (O_356,N_14622,N_14688);
and UO_357 (O_357,N_14882,N_14608);
nand UO_358 (O_358,N_14550,N_14757);
and UO_359 (O_359,N_14950,N_14707);
and UO_360 (O_360,N_14514,N_14739);
or UO_361 (O_361,N_14543,N_14872);
nand UO_362 (O_362,N_14818,N_14584);
xor UO_363 (O_363,N_14986,N_14688);
or UO_364 (O_364,N_14627,N_14794);
and UO_365 (O_365,N_14689,N_14555);
nor UO_366 (O_366,N_14561,N_14895);
nand UO_367 (O_367,N_14517,N_14629);
or UO_368 (O_368,N_14748,N_14936);
and UO_369 (O_369,N_14516,N_14699);
and UO_370 (O_370,N_14632,N_14746);
nand UO_371 (O_371,N_14751,N_14964);
nand UO_372 (O_372,N_14736,N_14988);
nand UO_373 (O_373,N_14547,N_14825);
nand UO_374 (O_374,N_14518,N_14772);
nor UO_375 (O_375,N_14959,N_14684);
xnor UO_376 (O_376,N_14922,N_14697);
xor UO_377 (O_377,N_14899,N_14945);
and UO_378 (O_378,N_14865,N_14779);
xor UO_379 (O_379,N_14632,N_14602);
nor UO_380 (O_380,N_14695,N_14710);
nand UO_381 (O_381,N_14855,N_14800);
or UO_382 (O_382,N_14978,N_14940);
xor UO_383 (O_383,N_14641,N_14556);
nor UO_384 (O_384,N_14985,N_14665);
or UO_385 (O_385,N_14808,N_14536);
xor UO_386 (O_386,N_14975,N_14802);
or UO_387 (O_387,N_14964,N_14793);
or UO_388 (O_388,N_14905,N_14755);
and UO_389 (O_389,N_14937,N_14970);
nand UO_390 (O_390,N_14625,N_14919);
and UO_391 (O_391,N_14638,N_14593);
or UO_392 (O_392,N_14818,N_14917);
nor UO_393 (O_393,N_14656,N_14811);
or UO_394 (O_394,N_14609,N_14645);
and UO_395 (O_395,N_14504,N_14891);
xnor UO_396 (O_396,N_14662,N_14618);
nand UO_397 (O_397,N_14561,N_14983);
and UO_398 (O_398,N_14890,N_14756);
nor UO_399 (O_399,N_14670,N_14571);
nand UO_400 (O_400,N_14567,N_14766);
and UO_401 (O_401,N_14791,N_14960);
xnor UO_402 (O_402,N_14973,N_14688);
nor UO_403 (O_403,N_14567,N_14982);
and UO_404 (O_404,N_14646,N_14518);
or UO_405 (O_405,N_14802,N_14621);
nand UO_406 (O_406,N_14698,N_14944);
nor UO_407 (O_407,N_14920,N_14850);
or UO_408 (O_408,N_14580,N_14865);
nor UO_409 (O_409,N_14991,N_14623);
or UO_410 (O_410,N_14799,N_14747);
xor UO_411 (O_411,N_14605,N_14731);
or UO_412 (O_412,N_14542,N_14686);
nor UO_413 (O_413,N_14556,N_14747);
or UO_414 (O_414,N_14566,N_14952);
nor UO_415 (O_415,N_14828,N_14516);
and UO_416 (O_416,N_14804,N_14524);
or UO_417 (O_417,N_14696,N_14941);
nand UO_418 (O_418,N_14651,N_14692);
xor UO_419 (O_419,N_14759,N_14928);
or UO_420 (O_420,N_14577,N_14969);
or UO_421 (O_421,N_14914,N_14801);
and UO_422 (O_422,N_14790,N_14679);
xor UO_423 (O_423,N_14561,N_14910);
and UO_424 (O_424,N_14682,N_14967);
nand UO_425 (O_425,N_14501,N_14539);
nand UO_426 (O_426,N_14507,N_14515);
or UO_427 (O_427,N_14789,N_14597);
and UO_428 (O_428,N_14516,N_14968);
nand UO_429 (O_429,N_14736,N_14878);
nand UO_430 (O_430,N_14976,N_14845);
nand UO_431 (O_431,N_14990,N_14604);
and UO_432 (O_432,N_14554,N_14829);
or UO_433 (O_433,N_14710,N_14757);
nand UO_434 (O_434,N_14513,N_14521);
xnor UO_435 (O_435,N_14639,N_14625);
xor UO_436 (O_436,N_14857,N_14593);
nor UO_437 (O_437,N_14537,N_14523);
nand UO_438 (O_438,N_14718,N_14980);
xor UO_439 (O_439,N_14686,N_14511);
and UO_440 (O_440,N_14625,N_14646);
and UO_441 (O_441,N_14608,N_14705);
or UO_442 (O_442,N_14987,N_14754);
nor UO_443 (O_443,N_14961,N_14951);
or UO_444 (O_444,N_14690,N_14774);
or UO_445 (O_445,N_14815,N_14645);
or UO_446 (O_446,N_14810,N_14645);
nand UO_447 (O_447,N_14512,N_14957);
or UO_448 (O_448,N_14874,N_14829);
and UO_449 (O_449,N_14778,N_14893);
and UO_450 (O_450,N_14923,N_14551);
nor UO_451 (O_451,N_14558,N_14711);
and UO_452 (O_452,N_14852,N_14693);
xnor UO_453 (O_453,N_14574,N_14874);
nor UO_454 (O_454,N_14713,N_14755);
and UO_455 (O_455,N_14762,N_14826);
xnor UO_456 (O_456,N_14661,N_14769);
nand UO_457 (O_457,N_14747,N_14769);
nand UO_458 (O_458,N_14642,N_14813);
xor UO_459 (O_459,N_14957,N_14500);
nand UO_460 (O_460,N_14731,N_14567);
xnor UO_461 (O_461,N_14781,N_14654);
nand UO_462 (O_462,N_14668,N_14677);
and UO_463 (O_463,N_14692,N_14814);
nor UO_464 (O_464,N_14717,N_14515);
and UO_465 (O_465,N_14984,N_14950);
and UO_466 (O_466,N_14701,N_14626);
nand UO_467 (O_467,N_14681,N_14778);
nor UO_468 (O_468,N_14919,N_14815);
or UO_469 (O_469,N_14855,N_14722);
nand UO_470 (O_470,N_14549,N_14930);
nand UO_471 (O_471,N_14935,N_14661);
or UO_472 (O_472,N_14601,N_14991);
nand UO_473 (O_473,N_14592,N_14737);
or UO_474 (O_474,N_14752,N_14706);
xor UO_475 (O_475,N_14944,N_14832);
xor UO_476 (O_476,N_14631,N_14938);
and UO_477 (O_477,N_14630,N_14755);
and UO_478 (O_478,N_14655,N_14637);
and UO_479 (O_479,N_14876,N_14856);
nand UO_480 (O_480,N_14869,N_14961);
or UO_481 (O_481,N_14576,N_14535);
nor UO_482 (O_482,N_14888,N_14500);
or UO_483 (O_483,N_14918,N_14669);
nand UO_484 (O_484,N_14948,N_14584);
xnor UO_485 (O_485,N_14709,N_14632);
nor UO_486 (O_486,N_14991,N_14863);
or UO_487 (O_487,N_14660,N_14593);
or UO_488 (O_488,N_14870,N_14688);
or UO_489 (O_489,N_14539,N_14586);
xor UO_490 (O_490,N_14809,N_14923);
and UO_491 (O_491,N_14645,N_14637);
and UO_492 (O_492,N_14567,N_14762);
xor UO_493 (O_493,N_14549,N_14632);
nor UO_494 (O_494,N_14921,N_14981);
nor UO_495 (O_495,N_14882,N_14551);
nor UO_496 (O_496,N_14610,N_14626);
nor UO_497 (O_497,N_14817,N_14744);
nand UO_498 (O_498,N_14517,N_14696);
or UO_499 (O_499,N_14874,N_14858);
and UO_500 (O_500,N_14782,N_14909);
nor UO_501 (O_501,N_14675,N_14600);
xor UO_502 (O_502,N_14524,N_14785);
and UO_503 (O_503,N_14655,N_14763);
and UO_504 (O_504,N_14946,N_14824);
nand UO_505 (O_505,N_14604,N_14904);
nand UO_506 (O_506,N_14937,N_14975);
nand UO_507 (O_507,N_14607,N_14534);
and UO_508 (O_508,N_14905,N_14586);
or UO_509 (O_509,N_14818,N_14737);
or UO_510 (O_510,N_14521,N_14788);
or UO_511 (O_511,N_14542,N_14837);
xnor UO_512 (O_512,N_14685,N_14829);
and UO_513 (O_513,N_14998,N_14761);
and UO_514 (O_514,N_14864,N_14511);
or UO_515 (O_515,N_14700,N_14875);
and UO_516 (O_516,N_14701,N_14860);
nor UO_517 (O_517,N_14651,N_14748);
nor UO_518 (O_518,N_14508,N_14933);
nor UO_519 (O_519,N_14749,N_14979);
xnor UO_520 (O_520,N_14790,N_14991);
nor UO_521 (O_521,N_14512,N_14740);
or UO_522 (O_522,N_14924,N_14948);
nand UO_523 (O_523,N_14710,N_14741);
nor UO_524 (O_524,N_14834,N_14610);
or UO_525 (O_525,N_14715,N_14935);
and UO_526 (O_526,N_14595,N_14881);
or UO_527 (O_527,N_14843,N_14973);
nor UO_528 (O_528,N_14612,N_14883);
nor UO_529 (O_529,N_14969,N_14892);
nor UO_530 (O_530,N_14619,N_14938);
or UO_531 (O_531,N_14814,N_14722);
and UO_532 (O_532,N_14622,N_14770);
and UO_533 (O_533,N_14634,N_14764);
xnor UO_534 (O_534,N_14909,N_14761);
or UO_535 (O_535,N_14645,N_14992);
xnor UO_536 (O_536,N_14945,N_14764);
or UO_537 (O_537,N_14908,N_14806);
or UO_538 (O_538,N_14833,N_14693);
or UO_539 (O_539,N_14712,N_14646);
nand UO_540 (O_540,N_14745,N_14544);
nor UO_541 (O_541,N_14989,N_14982);
nor UO_542 (O_542,N_14609,N_14655);
or UO_543 (O_543,N_14890,N_14538);
xnor UO_544 (O_544,N_14940,N_14682);
or UO_545 (O_545,N_14892,N_14991);
or UO_546 (O_546,N_14883,N_14877);
and UO_547 (O_547,N_14885,N_14782);
xor UO_548 (O_548,N_14978,N_14821);
nand UO_549 (O_549,N_14832,N_14781);
xor UO_550 (O_550,N_14702,N_14822);
nand UO_551 (O_551,N_14885,N_14802);
nand UO_552 (O_552,N_14840,N_14784);
xor UO_553 (O_553,N_14597,N_14750);
and UO_554 (O_554,N_14724,N_14813);
or UO_555 (O_555,N_14583,N_14765);
nand UO_556 (O_556,N_14962,N_14738);
nand UO_557 (O_557,N_14684,N_14682);
nand UO_558 (O_558,N_14732,N_14650);
or UO_559 (O_559,N_14815,N_14779);
and UO_560 (O_560,N_14536,N_14873);
or UO_561 (O_561,N_14787,N_14550);
nand UO_562 (O_562,N_14660,N_14648);
or UO_563 (O_563,N_14771,N_14922);
nor UO_564 (O_564,N_14505,N_14717);
xor UO_565 (O_565,N_14745,N_14815);
xnor UO_566 (O_566,N_14801,N_14787);
or UO_567 (O_567,N_14744,N_14802);
and UO_568 (O_568,N_14954,N_14725);
nor UO_569 (O_569,N_14553,N_14880);
nor UO_570 (O_570,N_14720,N_14685);
xor UO_571 (O_571,N_14610,N_14956);
or UO_572 (O_572,N_14895,N_14675);
or UO_573 (O_573,N_14781,N_14762);
nand UO_574 (O_574,N_14553,N_14977);
nor UO_575 (O_575,N_14559,N_14526);
or UO_576 (O_576,N_14765,N_14782);
or UO_577 (O_577,N_14579,N_14751);
nand UO_578 (O_578,N_14805,N_14724);
and UO_579 (O_579,N_14958,N_14808);
and UO_580 (O_580,N_14594,N_14511);
and UO_581 (O_581,N_14675,N_14571);
nor UO_582 (O_582,N_14891,N_14890);
nand UO_583 (O_583,N_14615,N_14895);
and UO_584 (O_584,N_14605,N_14653);
or UO_585 (O_585,N_14768,N_14531);
nand UO_586 (O_586,N_14882,N_14944);
xnor UO_587 (O_587,N_14851,N_14923);
nor UO_588 (O_588,N_14605,N_14848);
nand UO_589 (O_589,N_14609,N_14820);
nand UO_590 (O_590,N_14659,N_14676);
and UO_591 (O_591,N_14653,N_14919);
xnor UO_592 (O_592,N_14701,N_14523);
nand UO_593 (O_593,N_14606,N_14994);
xor UO_594 (O_594,N_14873,N_14985);
nor UO_595 (O_595,N_14794,N_14504);
nand UO_596 (O_596,N_14521,N_14576);
nand UO_597 (O_597,N_14779,N_14510);
or UO_598 (O_598,N_14873,N_14631);
nor UO_599 (O_599,N_14858,N_14824);
nand UO_600 (O_600,N_14790,N_14583);
nand UO_601 (O_601,N_14964,N_14501);
and UO_602 (O_602,N_14786,N_14602);
nor UO_603 (O_603,N_14925,N_14713);
or UO_604 (O_604,N_14765,N_14851);
and UO_605 (O_605,N_14876,N_14966);
and UO_606 (O_606,N_14521,N_14861);
xnor UO_607 (O_607,N_14803,N_14788);
and UO_608 (O_608,N_14815,N_14752);
nand UO_609 (O_609,N_14988,N_14685);
and UO_610 (O_610,N_14703,N_14636);
nor UO_611 (O_611,N_14981,N_14633);
and UO_612 (O_612,N_14882,N_14650);
nor UO_613 (O_613,N_14607,N_14955);
or UO_614 (O_614,N_14927,N_14990);
nor UO_615 (O_615,N_14931,N_14942);
xnor UO_616 (O_616,N_14505,N_14976);
and UO_617 (O_617,N_14972,N_14692);
xnor UO_618 (O_618,N_14921,N_14963);
and UO_619 (O_619,N_14958,N_14778);
nand UO_620 (O_620,N_14892,N_14806);
nor UO_621 (O_621,N_14830,N_14657);
or UO_622 (O_622,N_14673,N_14735);
and UO_623 (O_623,N_14659,N_14622);
or UO_624 (O_624,N_14762,N_14664);
xnor UO_625 (O_625,N_14791,N_14992);
nor UO_626 (O_626,N_14836,N_14749);
nor UO_627 (O_627,N_14565,N_14599);
nor UO_628 (O_628,N_14540,N_14974);
and UO_629 (O_629,N_14670,N_14568);
and UO_630 (O_630,N_14973,N_14937);
and UO_631 (O_631,N_14664,N_14781);
or UO_632 (O_632,N_14524,N_14662);
xnor UO_633 (O_633,N_14753,N_14777);
and UO_634 (O_634,N_14737,N_14712);
xnor UO_635 (O_635,N_14990,N_14532);
or UO_636 (O_636,N_14655,N_14671);
xnor UO_637 (O_637,N_14532,N_14915);
or UO_638 (O_638,N_14987,N_14724);
and UO_639 (O_639,N_14918,N_14868);
xnor UO_640 (O_640,N_14615,N_14889);
nor UO_641 (O_641,N_14616,N_14602);
or UO_642 (O_642,N_14631,N_14608);
nand UO_643 (O_643,N_14515,N_14881);
xnor UO_644 (O_644,N_14540,N_14804);
and UO_645 (O_645,N_14715,N_14890);
and UO_646 (O_646,N_14659,N_14883);
and UO_647 (O_647,N_14538,N_14927);
and UO_648 (O_648,N_14588,N_14574);
and UO_649 (O_649,N_14748,N_14981);
nand UO_650 (O_650,N_14872,N_14623);
and UO_651 (O_651,N_14541,N_14703);
nor UO_652 (O_652,N_14708,N_14635);
or UO_653 (O_653,N_14590,N_14728);
xnor UO_654 (O_654,N_14895,N_14527);
xor UO_655 (O_655,N_14735,N_14886);
nand UO_656 (O_656,N_14507,N_14933);
nor UO_657 (O_657,N_14831,N_14771);
nand UO_658 (O_658,N_14572,N_14709);
nand UO_659 (O_659,N_14506,N_14796);
nand UO_660 (O_660,N_14503,N_14610);
xor UO_661 (O_661,N_14726,N_14768);
and UO_662 (O_662,N_14787,N_14735);
nand UO_663 (O_663,N_14557,N_14756);
xor UO_664 (O_664,N_14651,N_14736);
nor UO_665 (O_665,N_14731,N_14610);
xnor UO_666 (O_666,N_14671,N_14500);
and UO_667 (O_667,N_14683,N_14616);
nand UO_668 (O_668,N_14567,N_14570);
or UO_669 (O_669,N_14843,N_14937);
nor UO_670 (O_670,N_14626,N_14987);
nor UO_671 (O_671,N_14771,N_14668);
nor UO_672 (O_672,N_14746,N_14846);
nor UO_673 (O_673,N_14800,N_14915);
nand UO_674 (O_674,N_14882,N_14822);
nand UO_675 (O_675,N_14689,N_14717);
nor UO_676 (O_676,N_14848,N_14713);
nor UO_677 (O_677,N_14915,N_14868);
nor UO_678 (O_678,N_14715,N_14722);
nor UO_679 (O_679,N_14854,N_14635);
nand UO_680 (O_680,N_14601,N_14520);
nand UO_681 (O_681,N_14512,N_14833);
xor UO_682 (O_682,N_14815,N_14798);
nor UO_683 (O_683,N_14902,N_14791);
and UO_684 (O_684,N_14811,N_14948);
xnor UO_685 (O_685,N_14646,N_14586);
and UO_686 (O_686,N_14824,N_14526);
nand UO_687 (O_687,N_14512,N_14745);
xor UO_688 (O_688,N_14799,N_14850);
nor UO_689 (O_689,N_14877,N_14880);
and UO_690 (O_690,N_14993,N_14769);
and UO_691 (O_691,N_14729,N_14612);
nand UO_692 (O_692,N_14856,N_14754);
nand UO_693 (O_693,N_14720,N_14871);
xor UO_694 (O_694,N_14570,N_14932);
and UO_695 (O_695,N_14884,N_14529);
or UO_696 (O_696,N_14640,N_14960);
nand UO_697 (O_697,N_14504,N_14992);
nor UO_698 (O_698,N_14826,N_14652);
and UO_699 (O_699,N_14539,N_14689);
or UO_700 (O_700,N_14793,N_14767);
xor UO_701 (O_701,N_14558,N_14995);
xor UO_702 (O_702,N_14661,N_14956);
and UO_703 (O_703,N_14548,N_14928);
nor UO_704 (O_704,N_14987,N_14917);
nor UO_705 (O_705,N_14692,N_14822);
nand UO_706 (O_706,N_14695,N_14752);
or UO_707 (O_707,N_14852,N_14788);
and UO_708 (O_708,N_14585,N_14695);
nand UO_709 (O_709,N_14578,N_14831);
or UO_710 (O_710,N_14847,N_14918);
nor UO_711 (O_711,N_14680,N_14897);
or UO_712 (O_712,N_14518,N_14589);
and UO_713 (O_713,N_14979,N_14528);
nand UO_714 (O_714,N_14792,N_14814);
nand UO_715 (O_715,N_14936,N_14754);
nand UO_716 (O_716,N_14738,N_14704);
or UO_717 (O_717,N_14992,N_14853);
xnor UO_718 (O_718,N_14602,N_14611);
and UO_719 (O_719,N_14687,N_14853);
nand UO_720 (O_720,N_14674,N_14985);
xor UO_721 (O_721,N_14656,N_14598);
nor UO_722 (O_722,N_14865,N_14881);
xnor UO_723 (O_723,N_14522,N_14515);
xor UO_724 (O_724,N_14646,N_14729);
nor UO_725 (O_725,N_14828,N_14781);
nand UO_726 (O_726,N_14578,N_14669);
or UO_727 (O_727,N_14615,N_14913);
xnor UO_728 (O_728,N_14510,N_14682);
xnor UO_729 (O_729,N_14992,N_14939);
or UO_730 (O_730,N_14575,N_14558);
nor UO_731 (O_731,N_14896,N_14841);
and UO_732 (O_732,N_14801,N_14597);
nand UO_733 (O_733,N_14772,N_14832);
xor UO_734 (O_734,N_14825,N_14964);
xnor UO_735 (O_735,N_14553,N_14790);
and UO_736 (O_736,N_14551,N_14825);
and UO_737 (O_737,N_14518,N_14630);
or UO_738 (O_738,N_14904,N_14978);
xor UO_739 (O_739,N_14982,N_14947);
or UO_740 (O_740,N_14531,N_14991);
nor UO_741 (O_741,N_14787,N_14813);
xor UO_742 (O_742,N_14571,N_14870);
or UO_743 (O_743,N_14890,N_14914);
and UO_744 (O_744,N_14961,N_14548);
nor UO_745 (O_745,N_14679,N_14716);
nor UO_746 (O_746,N_14840,N_14794);
xor UO_747 (O_747,N_14769,N_14756);
xor UO_748 (O_748,N_14822,N_14872);
or UO_749 (O_749,N_14904,N_14787);
nand UO_750 (O_750,N_14600,N_14774);
or UO_751 (O_751,N_14844,N_14749);
or UO_752 (O_752,N_14553,N_14771);
and UO_753 (O_753,N_14939,N_14605);
xor UO_754 (O_754,N_14612,N_14689);
nor UO_755 (O_755,N_14889,N_14664);
xnor UO_756 (O_756,N_14504,N_14942);
nor UO_757 (O_757,N_14995,N_14537);
xnor UO_758 (O_758,N_14678,N_14973);
nor UO_759 (O_759,N_14608,N_14975);
or UO_760 (O_760,N_14575,N_14705);
nand UO_761 (O_761,N_14916,N_14711);
nand UO_762 (O_762,N_14769,N_14789);
nand UO_763 (O_763,N_14889,N_14525);
xor UO_764 (O_764,N_14879,N_14633);
nand UO_765 (O_765,N_14716,N_14900);
nor UO_766 (O_766,N_14623,N_14714);
and UO_767 (O_767,N_14819,N_14911);
or UO_768 (O_768,N_14765,N_14649);
xor UO_769 (O_769,N_14705,N_14923);
or UO_770 (O_770,N_14649,N_14921);
and UO_771 (O_771,N_14886,N_14647);
and UO_772 (O_772,N_14578,N_14958);
nand UO_773 (O_773,N_14990,N_14781);
and UO_774 (O_774,N_14643,N_14541);
nor UO_775 (O_775,N_14521,N_14966);
nor UO_776 (O_776,N_14695,N_14582);
and UO_777 (O_777,N_14980,N_14817);
and UO_778 (O_778,N_14771,N_14972);
nor UO_779 (O_779,N_14743,N_14999);
xor UO_780 (O_780,N_14620,N_14693);
and UO_781 (O_781,N_14797,N_14915);
nor UO_782 (O_782,N_14779,N_14773);
nor UO_783 (O_783,N_14819,N_14857);
nor UO_784 (O_784,N_14924,N_14684);
nor UO_785 (O_785,N_14759,N_14823);
nand UO_786 (O_786,N_14873,N_14803);
or UO_787 (O_787,N_14638,N_14840);
nor UO_788 (O_788,N_14742,N_14754);
xor UO_789 (O_789,N_14738,N_14619);
nand UO_790 (O_790,N_14762,N_14663);
or UO_791 (O_791,N_14533,N_14965);
or UO_792 (O_792,N_14833,N_14930);
and UO_793 (O_793,N_14846,N_14931);
or UO_794 (O_794,N_14823,N_14866);
nor UO_795 (O_795,N_14840,N_14816);
or UO_796 (O_796,N_14935,N_14998);
xnor UO_797 (O_797,N_14665,N_14916);
nor UO_798 (O_798,N_14907,N_14738);
nor UO_799 (O_799,N_14553,N_14903);
xnor UO_800 (O_800,N_14841,N_14745);
nand UO_801 (O_801,N_14925,N_14542);
xor UO_802 (O_802,N_14571,N_14911);
nor UO_803 (O_803,N_14826,N_14638);
and UO_804 (O_804,N_14581,N_14935);
xnor UO_805 (O_805,N_14638,N_14891);
nor UO_806 (O_806,N_14744,N_14885);
nor UO_807 (O_807,N_14522,N_14930);
xnor UO_808 (O_808,N_14895,N_14588);
xnor UO_809 (O_809,N_14510,N_14826);
xor UO_810 (O_810,N_14688,N_14505);
and UO_811 (O_811,N_14903,N_14856);
and UO_812 (O_812,N_14804,N_14538);
and UO_813 (O_813,N_14837,N_14619);
nand UO_814 (O_814,N_14993,N_14798);
nand UO_815 (O_815,N_14569,N_14525);
xnor UO_816 (O_816,N_14771,N_14538);
and UO_817 (O_817,N_14634,N_14653);
nor UO_818 (O_818,N_14849,N_14931);
nand UO_819 (O_819,N_14649,N_14797);
and UO_820 (O_820,N_14987,N_14564);
or UO_821 (O_821,N_14867,N_14525);
and UO_822 (O_822,N_14858,N_14998);
and UO_823 (O_823,N_14519,N_14979);
nand UO_824 (O_824,N_14922,N_14647);
nor UO_825 (O_825,N_14575,N_14735);
nor UO_826 (O_826,N_14935,N_14872);
or UO_827 (O_827,N_14717,N_14911);
xnor UO_828 (O_828,N_14790,N_14631);
nand UO_829 (O_829,N_14518,N_14562);
xor UO_830 (O_830,N_14614,N_14928);
nor UO_831 (O_831,N_14853,N_14771);
nand UO_832 (O_832,N_14954,N_14659);
nand UO_833 (O_833,N_14760,N_14849);
nand UO_834 (O_834,N_14944,N_14839);
nor UO_835 (O_835,N_14544,N_14781);
nand UO_836 (O_836,N_14671,N_14561);
or UO_837 (O_837,N_14933,N_14546);
or UO_838 (O_838,N_14502,N_14501);
or UO_839 (O_839,N_14676,N_14651);
xnor UO_840 (O_840,N_14684,N_14587);
and UO_841 (O_841,N_14534,N_14710);
nor UO_842 (O_842,N_14873,N_14831);
or UO_843 (O_843,N_14953,N_14756);
nor UO_844 (O_844,N_14841,N_14713);
and UO_845 (O_845,N_14761,N_14669);
and UO_846 (O_846,N_14971,N_14976);
xor UO_847 (O_847,N_14914,N_14597);
nor UO_848 (O_848,N_14875,N_14511);
nand UO_849 (O_849,N_14897,N_14623);
and UO_850 (O_850,N_14773,N_14728);
nand UO_851 (O_851,N_14978,N_14606);
nor UO_852 (O_852,N_14769,N_14839);
or UO_853 (O_853,N_14552,N_14615);
and UO_854 (O_854,N_14985,N_14522);
nand UO_855 (O_855,N_14547,N_14714);
nor UO_856 (O_856,N_14752,N_14605);
xor UO_857 (O_857,N_14856,N_14544);
xor UO_858 (O_858,N_14774,N_14737);
nor UO_859 (O_859,N_14566,N_14517);
and UO_860 (O_860,N_14744,N_14762);
or UO_861 (O_861,N_14843,N_14643);
nand UO_862 (O_862,N_14573,N_14969);
and UO_863 (O_863,N_14999,N_14914);
xor UO_864 (O_864,N_14890,N_14931);
nand UO_865 (O_865,N_14960,N_14916);
or UO_866 (O_866,N_14544,N_14955);
nor UO_867 (O_867,N_14640,N_14602);
xnor UO_868 (O_868,N_14525,N_14759);
xnor UO_869 (O_869,N_14924,N_14954);
and UO_870 (O_870,N_14729,N_14551);
nand UO_871 (O_871,N_14511,N_14911);
nand UO_872 (O_872,N_14939,N_14811);
xor UO_873 (O_873,N_14920,N_14516);
nor UO_874 (O_874,N_14706,N_14847);
nand UO_875 (O_875,N_14883,N_14875);
nand UO_876 (O_876,N_14806,N_14564);
and UO_877 (O_877,N_14896,N_14867);
or UO_878 (O_878,N_14620,N_14719);
nor UO_879 (O_879,N_14567,N_14741);
nand UO_880 (O_880,N_14796,N_14651);
or UO_881 (O_881,N_14869,N_14531);
or UO_882 (O_882,N_14999,N_14614);
nor UO_883 (O_883,N_14631,N_14585);
or UO_884 (O_884,N_14596,N_14618);
nand UO_885 (O_885,N_14501,N_14580);
nand UO_886 (O_886,N_14922,N_14587);
nand UO_887 (O_887,N_14656,N_14659);
or UO_888 (O_888,N_14621,N_14591);
nor UO_889 (O_889,N_14533,N_14637);
xnor UO_890 (O_890,N_14983,N_14817);
or UO_891 (O_891,N_14955,N_14922);
xnor UO_892 (O_892,N_14653,N_14650);
xor UO_893 (O_893,N_14714,N_14940);
or UO_894 (O_894,N_14573,N_14851);
nand UO_895 (O_895,N_14902,N_14952);
xor UO_896 (O_896,N_14908,N_14910);
and UO_897 (O_897,N_14667,N_14913);
and UO_898 (O_898,N_14817,N_14691);
xnor UO_899 (O_899,N_14643,N_14609);
nor UO_900 (O_900,N_14818,N_14609);
xnor UO_901 (O_901,N_14766,N_14838);
and UO_902 (O_902,N_14868,N_14785);
or UO_903 (O_903,N_14588,N_14545);
or UO_904 (O_904,N_14813,N_14614);
or UO_905 (O_905,N_14929,N_14975);
or UO_906 (O_906,N_14666,N_14656);
xnor UO_907 (O_907,N_14605,N_14825);
or UO_908 (O_908,N_14781,N_14603);
xor UO_909 (O_909,N_14634,N_14794);
or UO_910 (O_910,N_14836,N_14685);
or UO_911 (O_911,N_14808,N_14834);
or UO_912 (O_912,N_14641,N_14763);
or UO_913 (O_913,N_14848,N_14804);
and UO_914 (O_914,N_14620,N_14765);
xnor UO_915 (O_915,N_14791,N_14789);
xor UO_916 (O_916,N_14619,N_14833);
nor UO_917 (O_917,N_14964,N_14943);
nand UO_918 (O_918,N_14845,N_14786);
xnor UO_919 (O_919,N_14568,N_14780);
or UO_920 (O_920,N_14667,N_14576);
xnor UO_921 (O_921,N_14936,N_14798);
nor UO_922 (O_922,N_14591,N_14596);
and UO_923 (O_923,N_14996,N_14800);
or UO_924 (O_924,N_14603,N_14950);
and UO_925 (O_925,N_14753,N_14556);
xor UO_926 (O_926,N_14911,N_14624);
or UO_927 (O_927,N_14940,N_14959);
nand UO_928 (O_928,N_14796,N_14630);
or UO_929 (O_929,N_14706,N_14504);
nand UO_930 (O_930,N_14843,N_14909);
nor UO_931 (O_931,N_14988,N_14821);
or UO_932 (O_932,N_14706,N_14843);
nor UO_933 (O_933,N_14560,N_14522);
or UO_934 (O_934,N_14686,N_14636);
nand UO_935 (O_935,N_14872,N_14656);
and UO_936 (O_936,N_14968,N_14754);
nand UO_937 (O_937,N_14974,N_14910);
nor UO_938 (O_938,N_14646,N_14958);
and UO_939 (O_939,N_14874,N_14713);
and UO_940 (O_940,N_14825,N_14740);
or UO_941 (O_941,N_14771,N_14796);
xor UO_942 (O_942,N_14820,N_14792);
nor UO_943 (O_943,N_14810,N_14520);
xor UO_944 (O_944,N_14596,N_14735);
xor UO_945 (O_945,N_14862,N_14849);
nor UO_946 (O_946,N_14930,N_14573);
xor UO_947 (O_947,N_14548,N_14714);
nand UO_948 (O_948,N_14855,N_14899);
or UO_949 (O_949,N_14758,N_14671);
and UO_950 (O_950,N_14836,N_14839);
or UO_951 (O_951,N_14958,N_14698);
nand UO_952 (O_952,N_14992,N_14865);
and UO_953 (O_953,N_14682,N_14855);
xor UO_954 (O_954,N_14611,N_14735);
xnor UO_955 (O_955,N_14649,N_14507);
xor UO_956 (O_956,N_14554,N_14701);
or UO_957 (O_957,N_14826,N_14772);
and UO_958 (O_958,N_14950,N_14786);
nor UO_959 (O_959,N_14615,N_14543);
xor UO_960 (O_960,N_14793,N_14856);
xnor UO_961 (O_961,N_14690,N_14839);
or UO_962 (O_962,N_14542,N_14581);
or UO_963 (O_963,N_14815,N_14825);
nand UO_964 (O_964,N_14741,N_14867);
nor UO_965 (O_965,N_14994,N_14814);
nor UO_966 (O_966,N_14920,N_14728);
or UO_967 (O_967,N_14731,N_14741);
xnor UO_968 (O_968,N_14658,N_14914);
or UO_969 (O_969,N_14852,N_14601);
xor UO_970 (O_970,N_14994,N_14516);
nor UO_971 (O_971,N_14948,N_14586);
xor UO_972 (O_972,N_14946,N_14894);
xnor UO_973 (O_973,N_14825,N_14882);
and UO_974 (O_974,N_14961,N_14643);
or UO_975 (O_975,N_14794,N_14883);
xnor UO_976 (O_976,N_14999,N_14607);
xor UO_977 (O_977,N_14811,N_14877);
or UO_978 (O_978,N_14708,N_14714);
nor UO_979 (O_979,N_14677,N_14806);
nand UO_980 (O_980,N_14892,N_14869);
or UO_981 (O_981,N_14933,N_14995);
or UO_982 (O_982,N_14931,N_14699);
xor UO_983 (O_983,N_14780,N_14980);
nand UO_984 (O_984,N_14948,N_14780);
nand UO_985 (O_985,N_14662,N_14728);
nand UO_986 (O_986,N_14778,N_14687);
and UO_987 (O_987,N_14982,N_14622);
xor UO_988 (O_988,N_14747,N_14841);
nand UO_989 (O_989,N_14708,N_14888);
xnor UO_990 (O_990,N_14617,N_14925);
nand UO_991 (O_991,N_14989,N_14541);
xnor UO_992 (O_992,N_14766,N_14599);
nand UO_993 (O_993,N_14967,N_14533);
nor UO_994 (O_994,N_14816,N_14598);
nor UO_995 (O_995,N_14670,N_14808);
or UO_996 (O_996,N_14743,N_14754);
or UO_997 (O_997,N_14586,N_14917);
and UO_998 (O_998,N_14623,N_14929);
nand UO_999 (O_999,N_14961,N_14559);
nor UO_1000 (O_1000,N_14879,N_14623);
and UO_1001 (O_1001,N_14550,N_14777);
or UO_1002 (O_1002,N_14731,N_14943);
xor UO_1003 (O_1003,N_14638,N_14903);
xnor UO_1004 (O_1004,N_14721,N_14992);
xnor UO_1005 (O_1005,N_14881,N_14610);
nand UO_1006 (O_1006,N_14776,N_14745);
and UO_1007 (O_1007,N_14700,N_14534);
xnor UO_1008 (O_1008,N_14776,N_14965);
and UO_1009 (O_1009,N_14564,N_14766);
and UO_1010 (O_1010,N_14973,N_14613);
or UO_1011 (O_1011,N_14689,N_14850);
nand UO_1012 (O_1012,N_14901,N_14517);
xnor UO_1013 (O_1013,N_14794,N_14811);
or UO_1014 (O_1014,N_14580,N_14733);
and UO_1015 (O_1015,N_14838,N_14639);
or UO_1016 (O_1016,N_14966,N_14621);
xor UO_1017 (O_1017,N_14657,N_14733);
nor UO_1018 (O_1018,N_14695,N_14758);
xnor UO_1019 (O_1019,N_14644,N_14695);
nand UO_1020 (O_1020,N_14533,N_14945);
nand UO_1021 (O_1021,N_14986,N_14910);
xnor UO_1022 (O_1022,N_14668,N_14983);
nand UO_1023 (O_1023,N_14977,N_14787);
xnor UO_1024 (O_1024,N_14864,N_14520);
or UO_1025 (O_1025,N_14579,N_14833);
xor UO_1026 (O_1026,N_14565,N_14798);
and UO_1027 (O_1027,N_14795,N_14563);
nor UO_1028 (O_1028,N_14733,N_14612);
or UO_1029 (O_1029,N_14832,N_14948);
or UO_1030 (O_1030,N_14953,N_14557);
nor UO_1031 (O_1031,N_14798,N_14948);
nor UO_1032 (O_1032,N_14741,N_14949);
nand UO_1033 (O_1033,N_14866,N_14773);
or UO_1034 (O_1034,N_14550,N_14927);
or UO_1035 (O_1035,N_14867,N_14639);
or UO_1036 (O_1036,N_14698,N_14877);
nor UO_1037 (O_1037,N_14633,N_14893);
nand UO_1038 (O_1038,N_14551,N_14844);
or UO_1039 (O_1039,N_14847,N_14698);
and UO_1040 (O_1040,N_14700,N_14750);
and UO_1041 (O_1041,N_14798,N_14695);
and UO_1042 (O_1042,N_14787,N_14820);
nor UO_1043 (O_1043,N_14924,N_14634);
and UO_1044 (O_1044,N_14819,N_14859);
xnor UO_1045 (O_1045,N_14551,N_14989);
nor UO_1046 (O_1046,N_14898,N_14512);
or UO_1047 (O_1047,N_14582,N_14931);
xor UO_1048 (O_1048,N_14786,N_14732);
and UO_1049 (O_1049,N_14956,N_14820);
xnor UO_1050 (O_1050,N_14513,N_14927);
nand UO_1051 (O_1051,N_14572,N_14616);
nor UO_1052 (O_1052,N_14704,N_14953);
xor UO_1053 (O_1053,N_14823,N_14598);
xor UO_1054 (O_1054,N_14989,N_14611);
nand UO_1055 (O_1055,N_14677,N_14843);
and UO_1056 (O_1056,N_14722,N_14523);
xnor UO_1057 (O_1057,N_14862,N_14740);
xor UO_1058 (O_1058,N_14780,N_14918);
and UO_1059 (O_1059,N_14999,N_14572);
nor UO_1060 (O_1060,N_14708,N_14855);
xor UO_1061 (O_1061,N_14926,N_14585);
or UO_1062 (O_1062,N_14718,N_14945);
or UO_1063 (O_1063,N_14923,N_14983);
or UO_1064 (O_1064,N_14799,N_14962);
and UO_1065 (O_1065,N_14793,N_14936);
and UO_1066 (O_1066,N_14873,N_14623);
or UO_1067 (O_1067,N_14962,N_14915);
nor UO_1068 (O_1068,N_14523,N_14663);
and UO_1069 (O_1069,N_14820,N_14883);
xnor UO_1070 (O_1070,N_14841,N_14818);
or UO_1071 (O_1071,N_14704,N_14575);
and UO_1072 (O_1072,N_14919,N_14817);
xnor UO_1073 (O_1073,N_14843,N_14925);
xor UO_1074 (O_1074,N_14785,N_14513);
nand UO_1075 (O_1075,N_14913,N_14768);
or UO_1076 (O_1076,N_14857,N_14848);
and UO_1077 (O_1077,N_14677,N_14645);
nand UO_1078 (O_1078,N_14723,N_14966);
xnor UO_1079 (O_1079,N_14933,N_14964);
nor UO_1080 (O_1080,N_14758,N_14931);
or UO_1081 (O_1081,N_14510,N_14708);
nand UO_1082 (O_1082,N_14996,N_14740);
or UO_1083 (O_1083,N_14626,N_14685);
nor UO_1084 (O_1084,N_14589,N_14871);
and UO_1085 (O_1085,N_14927,N_14802);
nand UO_1086 (O_1086,N_14762,N_14536);
xnor UO_1087 (O_1087,N_14973,N_14866);
nor UO_1088 (O_1088,N_14869,N_14524);
nand UO_1089 (O_1089,N_14822,N_14927);
or UO_1090 (O_1090,N_14883,N_14628);
xnor UO_1091 (O_1091,N_14547,N_14760);
xor UO_1092 (O_1092,N_14658,N_14821);
xor UO_1093 (O_1093,N_14540,N_14907);
nor UO_1094 (O_1094,N_14712,N_14764);
nand UO_1095 (O_1095,N_14616,N_14691);
xnor UO_1096 (O_1096,N_14635,N_14801);
nand UO_1097 (O_1097,N_14748,N_14620);
xor UO_1098 (O_1098,N_14828,N_14614);
and UO_1099 (O_1099,N_14886,N_14704);
and UO_1100 (O_1100,N_14519,N_14648);
xor UO_1101 (O_1101,N_14905,N_14719);
and UO_1102 (O_1102,N_14607,N_14894);
nor UO_1103 (O_1103,N_14980,N_14845);
or UO_1104 (O_1104,N_14571,N_14754);
nand UO_1105 (O_1105,N_14692,N_14888);
or UO_1106 (O_1106,N_14951,N_14528);
or UO_1107 (O_1107,N_14671,N_14512);
or UO_1108 (O_1108,N_14632,N_14970);
or UO_1109 (O_1109,N_14866,N_14669);
nand UO_1110 (O_1110,N_14896,N_14842);
xnor UO_1111 (O_1111,N_14940,N_14837);
nand UO_1112 (O_1112,N_14890,N_14717);
or UO_1113 (O_1113,N_14867,N_14758);
xnor UO_1114 (O_1114,N_14680,N_14533);
nand UO_1115 (O_1115,N_14906,N_14690);
nor UO_1116 (O_1116,N_14702,N_14622);
nand UO_1117 (O_1117,N_14971,N_14992);
or UO_1118 (O_1118,N_14585,N_14768);
and UO_1119 (O_1119,N_14550,N_14513);
or UO_1120 (O_1120,N_14555,N_14750);
nand UO_1121 (O_1121,N_14637,N_14993);
xnor UO_1122 (O_1122,N_14621,N_14521);
or UO_1123 (O_1123,N_14746,N_14709);
nand UO_1124 (O_1124,N_14934,N_14870);
or UO_1125 (O_1125,N_14831,N_14669);
and UO_1126 (O_1126,N_14613,N_14680);
nor UO_1127 (O_1127,N_14800,N_14913);
or UO_1128 (O_1128,N_14614,N_14759);
nor UO_1129 (O_1129,N_14814,N_14628);
and UO_1130 (O_1130,N_14936,N_14547);
nand UO_1131 (O_1131,N_14940,N_14963);
or UO_1132 (O_1132,N_14504,N_14960);
xnor UO_1133 (O_1133,N_14764,N_14706);
and UO_1134 (O_1134,N_14809,N_14950);
and UO_1135 (O_1135,N_14834,N_14503);
and UO_1136 (O_1136,N_14822,N_14574);
nand UO_1137 (O_1137,N_14657,N_14790);
nor UO_1138 (O_1138,N_14994,N_14628);
nor UO_1139 (O_1139,N_14666,N_14995);
and UO_1140 (O_1140,N_14820,N_14773);
nor UO_1141 (O_1141,N_14539,N_14671);
and UO_1142 (O_1142,N_14711,N_14512);
and UO_1143 (O_1143,N_14620,N_14894);
xor UO_1144 (O_1144,N_14696,N_14972);
and UO_1145 (O_1145,N_14877,N_14979);
or UO_1146 (O_1146,N_14599,N_14702);
nor UO_1147 (O_1147,N_14771,N_14760);
nand UO_1148 (O_1148,N_14781,N_14734);
nor UO_1149 (O_1149,N_14867,N_14535);
xor UO_1150 (O_1150,N_14619,N_14641);
and UO_1151 (O_1151,N_14970,N_14702);
xnor UO_1152 (O_1152,N_14823,N_14707);
and UO_1153 (O_1153,N_14663,N_14965);
or UO_1154 (O_1154,N_14683,N_14947);
nor UO_1155 (O_1155,N_14589,N_14785);
xnor UO_1156 (O_1156,N_14637,N_14794);
nand UO_1157 (O_1157,N_14960,N_14782);
and UO_1158 (O_1158,N_14943,N_14632);
and UO_1159 (O_1159,N_14959,N_14505);
or UO_1160 (O_1160,N_14716,N_14712);
and UO_1161 (O_1161,N_14650,N_14840);
nand UO_1162 (O_1162,N_14506,N_14930);
nor UO_1163 (O_1163,N_14600,N_14847);
or UO_1164 (O_1164,N_14832,N_14573);
nor UO_1165 (O_1165,N_14810,N_14668);
nor UO_1166 (O_1166,N_14629,N_14642);
nor UO_1167 (O_1167,N_14998,N_14910);
nor UO_1168 (O_1168,N_14918,N_14652);
nor UO_1169 (O_1169,N_14757,N_14724);
and UO_1170 (O_1170,N_14848,N_14579);
nand UO_1171 (O_1171,N_14577,N_14644);
or UO_1172 (O_1172,N_14788,N_14771);
and UO_1173 (O_1173,N_14572,N_14987);
or UO_1174 (O_1174,N_14656,N_14767);
nand UO_1175 (O_1175,N_14894,N_14571);
nor UO_1176 (O_1176,N_14611,N_14549);
or UO_1177 (O_1177,N_14906,N_14933);
and UO_1178 (O_1178,N_14520,N_14549);
nand UO_1179 (O_1179,N_14947,N_14713);
or UO_1180 (O_1180,N_14740,N_14734);
xnor UO_1181 (O_1181,N_14639,N_14836);
xnor UO_1182 (O_1182,N_14912,N_14577);
and UO_1183 (O_1183,N_14709,N_14987);
or UO_1184 (O_1184,N_14644,N_14848);
nor UO_1185 (O_1185,N_14937,N_14848);
nor UO_1186 (O_1186,N_14931,N_14805);
nand UO_1187 (O_1187,N_14650,N_14587);
xnor UO_1188 (O_1188,N_14697,N_14943);
and UO_1189 (O_1189,N_14787,N_14942);
and UO_1190 (O_1190,N_14818,N_14811);
and UO_1191 (O_1191,N_14650,N_14617);
or UO_1192 (O_1192,N_14669,N_14521);
xor UO_1193 (O_1193,N_14925,N_14687);
nor UO_1194 (O_1194,N_14712,N_14978);
and UO_1195 (O_1195,N_14967,N_14787);
nand UO_1196 (O_1196,N_14904,N_14913);
nand UO_1197 (O_1197,N_14644,N_14604);
nor UO_1198 (O_1198,N_14691,N_14644);
and UO_1199 (O_1199,N_14516,N_14935);
nand UO_1200 (O_1200,N_14567,N_14698);
or UO_1201 (O_1201,N_14853,N_14682);
and UO_1202 (O_1202,N_14927,N_14667);
nor UO_1203 (O_1203,N_14997,N_14754);
nor UO_1204 (O_1204,N_14572,N_14823);
xnor UO_1205 (O_1205,N_14564,N_14946);
and UO_1206 (O_1206,N_14666,N_14670);
nand UO_1207 (O_1207,N_14899,N_14844);
and UO_1208 (O_1208,N_14735,N_14978);
nor UO_1209 (O_1209,N_14711,N_14649);
nand UO_1210 (O_1210,N_14570,N_14902);
nand UO_1211 (O_1211,N_14927,N_14913);
nor UO_1212 (O_1212,N_14973,N_14987);
or UO_1213 (O_1213,N_14862,N_14596);
nor UO_1214 (O_1214,N_14703,N_14977);
or UO_1215 (O_1215,N_14830,N_14981);
xor UO_1216 (O_1216,N_14719,N_14961);
nand UO_1217 (O_1217,N_14633,N_14892);
nand UO_1218 (O_1218,N_14740,N_14904);
nand UO_1219 (O_1219,N_14577,N_14921);
or UO_1220 (O_1220,N_14627,N_14535);
nand UO_1221 (O_1221,N_14710,N_14912);
nand UO_1222 (O_1222,N_14730,N_14613);
xor UO_1223 (O_1223,N_14662,N_14801);
xor UO_1224 (O_1224,N_14910,N_14790);
xor UO_1225 (O_1225,N_14967,N_14632);
or UO_1226 (O_1226,N_14517,N_14732);
or UO_1227 (O_1227,N_14515,N_14826);
nand UO_1228 (O_1228,N_14771,N_14949);
or UO_1229 (O_1229,N_14811,N_14933);
and UO_1230 (O_1230,N_14831,N_14840);
xor UO_1231 (O_1231,N_14814,N_14578);
or UO_1232 (O_1232,N_14571,N_14719);
and UO_1233 (O_1233,N_14523,N_14560);
nand UO_1234 (O_1234,N_14610,N_14573);
or UO_1235 (O_1235,N_14968,N_14689);
nor UO_1236 (O_1236,N_14799,N_14512);
nand UO_1237 (O_1237,N_14781,N_14942);
nand UO_1238 (O_1238,N_14970,N_14885);
xnor UO_1239 (O_1239,N_14583,N_14543);
xnor UO_1240 (O_1240,N_14583,N_14619);
xor UO_1241 (O_1241,N_14539,N_14981);
nand UO_1242 (O_1242,N_14959,N_14799);
or UO_1243 (O_1243,N_14959,N_14661);
and UO_1244 (O_1244,N_14921,N_14663);
nand UO_1245 (O_1245,N_14640,N_14573);
nand UO_1246 (O_1246,N_14852,N_14619);
nor UO_1247 (O_1247,N_14648,N_14509);
nand UO_1248 (O_1248,N_14951,N_14618);
and UO_1249 (O_1249,N_14955,N_14849);
nand UO_1250 (O_1250,N_14600,N_14532);
xor UO_1251 (O_1251,N_14922,N_14556);
xnor UO_1252 (O_1252,N_14683,N_14785);
nor UO_1253 (O_1253,N_14741,N_14801);
and UO_1254 (O_1254,N_14581,N_14577);
or UO_1255 (O_1255,N_14582,N_14601);
or UO_1256 (O_1256,N_14996,N_14659);
and UO_1257 (O_1257,N_14804,N_14696);
or UO_1258 (O_1258,N_14804,N_14641);
and UO_1259 (O_1259,N_14701,N_14989);
nor UO_1260 (O_1260,N_14817,N_14890);
and UO_1261 (O_1261,N_14750,N_14934);
and UO_1262 (O_1262,N_14781,N_14936);
nor UO_1263 (O_1263,N_14888,N_14616);
and UO_1264 (O_1264,N_14805,N_14788);
xnor UO_1265 (O_1265,N_14623,N_14760);
and UO_1266 (O_1266,N_14608,N_14980);
and UO_1267 (O_1267,N_14993,N_14796);
xor UO_1268 (O_1268,N_14530,N_14621);
xnor UO_1269 (O_1269,N_14917,N_14574);
and UO_1270 (O_1270,N_14958,N_14774);
nand UO_1271 (O_1271,N_14629,N_14526);
xor UO_1272 (O_1272,N_14760,N_14770);
or UO_1273 (O_1273,N_14920,N_14984);
nor UO_1274 (O_1274,N_14898,N_14609);
and UO_1275 (O_1275,N_14543,N_14985);
xor UO_1276 (O_1276,N_14561,N_14821);
nor UO_1277 (O_1277,N_14744,N_14989);
nor UO_1278 (O_1278,N_14506,N_14760);
and UO_1279 (O_1279,N_14926,N_14730);
xor UO_1280 (O_1280,N_14682,N_14959);
or UO_1281 (O_1281,N_14812,N_14873);
and UO_1282 (O_1282,N_14973,N_14971);
or UO_1283 (O_1283,N_14759,N_14943);
nand UO_1284 (O_1284,N_14923,N_14684);
nor UO_1285 (O_1285,N_14517,N_14804);
xnor UO_1286 (O_1286,N_14922,N_14825);
nor UO_1287 (O_1287,N_14798,N_14551);
nand UO_1288 (O_1288,N_14508,N_14924);
nand UO_1289 (O_1289,N_14696,N_14761);
nor UO_1290 (O_1290,N_14586,N_14752);
or UO_1291 (O_1291,N_14629,N_14716);
nand UO_1292 (O_1292,N_14892,N_14651);
nor UO_1293 (O_1293,N_14688,N_14716);
nand UO_1294 (O_1294,N_14762,N_14897);
nand UO_1295 (O_1295,N_14621,N_14729);
and UO_1296 (O_1296,N_14542,N_14890);
or UO_1297 (O_1297,N_14896,N_14526);
xnor UO_1298 (O_1298,N_14725,N_14938);
xor UO_1299 (O_1299,N_14577,N_14729);
and UO_1300 (O_1300,N_14975,N_14932);
or UO_1301 (O_1301,N_14505,N_14767);
and UO_1302 (O_1302,N_14999,N_14588);
nor UO_1303 (O_1303,N_14732,N_14787);
and UO_1304 (O_1304,N_14576,N_14967);
and UO_1305 (O_1305,N_14538,N_14994);
xor UO_1306 (O_1306,N_14958,N_14723);
or UO_1307 (O_1307,N_14826,N_14973);
nand UO_1308 (O_1308,N_14520,N_14834);
nand UO_1309 (O_1309,N_14874,N_14737);
nand UO_1310 (O_1310,N_14896,N_14649);
nor UO_1311 (O_1311,N_14959,N_14983);
xor UO_1312 (O_1312,N_14619,N_14767);
or UO_1313 (O_1313,N_14590,N_14834);
or UO_1314 (O_1314,N_14780,N_14885);
or UO_1315 (O_1315,N_14971,N_14829);
xnor UO_1316 (O_1316,N_14670,N_14748);
xor UO_1317 (O_1317,N_14710,N_14572);
and UO_1318 (O_1318,N_14573,N_14515);
or UO_1319 (O_1319,N_14772,N_14573);
or UO_1320 (O_1320,N_14539,N_14515);
and UO_1321 (O_1321,N_14594,N_14804);
nand UO_1322 (O_1322,N_14522,N_14887);
xnor UO_1323 (O_1323,N_14787,N_14745);
nand UO_1324 (O_1324,N_14649,N_14902);
and UO_1325 (O_1325,N_14994,N_14880);
nor UO_1326 (O_1326,N_14588,N_14917);
or UO_1327 (O_1327,N_14578,N_14732);
nand UO_1328 (O_1328,N_14796,N_14954);
xor UO_1329 (O_1329,N_14734,N_14889);
or UO_1330 (O_1330,N_14980,N_14946);
nand UO_1331 (O_1331,N_14851,N_14754);
or UO_1332 (O_1332,N_14525,N_14740);
nand UO_1333 (O_1333,N_14757,N_14510);
nor UO_1334 (O_1334,N_14666,N_14910);
nand UO_1335 (O_1335,N_14919,N_14612);
and UO_1336 (O_1336,N_14884,N_14640);
and UO_1337 (O_1337,N_14732,N_14527);
nor UO_1338 (O_1338,N_14935,N_14721);
or UO_1339 (O_1339,N_14788,N_14861);
nor UO_1340 (O_1340,N_14637,N_14727);
and UO_1341 (O_1341,N_14799,N_14980);
and UO_1342 (O_1342,N_14891,N_14697);
or UO_1343 (O_1343,N_14561,N_14965);
nand UO_1344 (O_1344,N_14523,N_14977);
xnor UO_1345 (O_1345,N_14846,N_14532);
and UO_1346 (O_1346,N_14782,N_14630);
or UO_1347 (O_1347,N_14624,N_14684);
nor UO_1348 (O_1348,N_14609,N_14998);
nand UO_1349 (O_1349,N_14767,N_14943);
nor UO_1350 (O_1350,N_14915,N_14966);
or UO_1351 (O_1351,N_14808,N_14897);
or UO_1352 (O_1352,N_14685,N_14888);
and UO_1353 (O_1353,N_14642,N_14769);
xor UO_1354 (O_1354,N_14691,N_14561);
and UO_1355 (O_1355,N_14584,N_14689);
nor UO_1356 (O_1356,N_14832,N_14590);
nand UO_1357 (O_1357,N_14912,N_14971);
and UO_1358 (O_1358,N_14573,N_14826);
nor UO_1359 (O_1359,N_14750,N_14729);
or UO_1360 (O_1360,N_14820,N_14886);
xor UO_1361 (O_1361,N_14559,N_14809);
nand UO_1362 (O_1362,N_14736,N_14865);
xnor UO_1363 (O_1363,N_14810,N_14995);
or UO_1364 (O_1364,N_14718,N_14677);
xnor UO_1365 (O_1365,N_14913,N_14752);
nand UO_1366 (O_1366,N_14625,N_14623);
or UO_1367 (O_1367,N_14950,N_14850);
nand UO_1368 (O_1368,N_14965,N_14963);
nand UO_1369 (O_1369,N_14755,N_14706);
or UO_1370 (O_1370,N_14882,N_14850);
nor UO_1371 (O_1371,N_14569,N_14813);
and UO_1372 (O_1372,N_14824,N_14634);
xnor UO_1373 (O_1373,N_14635,N_14770);
nor UO_1374 (O_1374,N_14959,N_14817);
nand UO_1375 (O_1375,N_14884,N_14668);
or UO_1376 (O_1376,N_14725,N_14910);
or UO_1377 (O_1377,N_14596,N_14915);
nor UO_1378 (O_1378,N_14567,N_14968);
xnor UO_1379 (O_1379,N_14821,N_14673);
nor UO_1380 (O_1380,N_14722,N_14539);
nand UO_1381 (O_1381,N_14859,N_14761);
or UO_1382 (O_1382,N_14709,N_14504);
nand UO_1383 (O_1383,N_14650,N_14783);
and UO_1384 (O_1384,N_14723,N_14569);
xnor UO_1385 (O_1385,N_14905,N_14791);
or UO_1386 (O_1386,N_14782,N_14606);
nor UO_1387 (O_1387,N_14856,N_14710);
or UO_1388 (O_1388,N_14745,N_14728);
or UO_1389 (O_1389,N_14667,N_14642);
nor UO_1390 (O_1390,N_14539,N_14638);
and UO_1391 (O_1391,N_14532,N_14833);
and UO_1392 (O_1392,N_14518,N_14991);
nor UO_1393 (O_1393,N_14568,N_14986);
and UO_1394 (O_1394,N_14548,N_14878);
and UO_1395 (O_1395,N_14894,N_14747);
xor UO_1396 (O_1396,N_14831,N_14679);
xnor UO_1397 (O_1397,N_14791,N_14899);
and UO_1398 (O_1398,N_14593,N_14907);
or UO_1399 (O_1399,N_14754,N_14889);
or UO_1400 (O_1400,N_14856,N_14669);
nor UO_1401 (O_1401,N_14668,N_14743);
xnor UO_1402 (O_1402,N_14600,N_14666);
and UO_1403 (O_1403,N_14911,N_14936);
xor UO_1404 (O_1404,N_14611,N_14704);
xnor UO_1405 (O_1405,N_14502,N_14737);
nand UO_1406 (O_1406,N_14588,N_14577);
and UO_1407 (O_1407,N_14932,N_14752);
xor UO_1408 (O_1408,N_14514,N_14762);
xnor UO_1409 (O_1409,N_14560,N_14519);
nand UO_1410 (O_1410,N_14784,N_14938);
xor UO_1411 (O_1411,N_14772,N_14605);
nor UO_1412 (O_1412,N_14836,N_14832);
or UO_1413 (O_1413,N_14695,N_14789);
nand UO_1414 (O_1414,N_14821,N_14973);
or UO_1415 (O_1415,N_14637,N_14516);
nor UO_1416 (O_1416,N_14506,N_14649);
and UO_1417 (O_1417,N_14836,N_14867);
and UO_1418 (O_1418,N_14843,N_14554);
nor UO_1419 (O_1419,N_14848,N_14552);
nor UO_1420 (O_1420,N_14644,N_14687);
and UO_1421 (O_1421,N_14527,N_14885);
nor UO_1422 (O_1422,N_14775,N_14774);
or UO_1423 (O_1423,N_14527,N_14540);
or UO_1424 (O_1424,N_14603,N_14840);
nand UO_1425 (O_1425,N_14664,N_14540);
or UO_1426 (O_1426,N_14965,N_14680);
and UO_1427 (O_1427,N_14912,N_14595);
nand UO_1428 (O_1428,N_14923,N_14863);
or UO_1429 (O_1429,N_14976,N_14638);
and UO_1430 (O_1430,N_14812,N_14664);
nand UO_1431 (O_1431,N_14807,N_14626);
xor UO_1432 (O_1432,N_14664,N_14868);
and UO_1433 (O_1433,N_14917,N_14544);
nand UO_1434 (O_1434,N_14999,N_14893);
and UO_1435 (O_1435,N_14820,N_14930);
or UO_1436 (O_1436,N_14695,N_14723);
and UO_1437 (O_1437,N_14691,N_14828);
and UO_1438 (O_1438,N_14633,N_14556);
nor UO_1439 (O_1439,N_14527,N_14641);
or UO_1440 (O_1440,N_14953,N_14878);
xor UO_1441 (O_1441,N_14678,N_14739);
nand UO_1442 (O_1442,N_14983,N_14623);
and UO_1443 (O_1443,N_14922,N_14526);
or UO_1444 (O_1444,N_14569,N_14761);
or UO_1445 (O_1445,N_14831,N_14546);
nand UO_1446 (O_1446,N_14765,N_14945);
nor UO_1447 (O_1447,N_14578,N_14919);
nor UO_1448 (O_1448,N_14529,N_14993);
nand UO_1449 (O_1449,N_14577,N_14824);
and UO_1450 (O_1450,N_14732,N_14617);
or UO_1451 (O_1451,N_14694,N_14862);
or UO_1452 (O_1452,N_14543,N_14520);
xor UO_1453 (O_1453,N_14776,N_14667);
nor UO_1454 (O_1454,N_14861,N_14917);
nor UO_1455 (O_1455,N_14528,N_14833);
or UO_1456 (O_1456,N_14791,N_14665);
xor UO_1457 (O_1457,N_14729,N_14948);
nand UO_1458 (O_1458,N_14937,N_14506);
nand UO_1459 (O_1459,N_14785,N_14962);
nand UO_1460 (O_1460,N_14579,N_14924);
nand UO_1461 (O_1461,N_14746,N_14910);
nor UO_1462 (O_1462,N_14768,N_14579);
nor UO_1463 (O_1463,N_14710,N_14786);
nor UO_1464 (O_1464,N_14517,N_14974);
nor UO_1465 (O_1465,N_14811,N_14792);
and UO_1466 (O_1466,N_14644,N_14536);
xnor UO_1467 (O_1467,N_14965,N_14805);
or UO_1468 (O_1468,N_14807,N_14698);
xnor UO_1469 (O_1469,N_14911,N_14700);
or UO_1470 (O_1470,N_14875,N_14948);
and UO_1471 (O_1471,N_14637,N_14760);
nor UO_1472 (O_1472,N_14508,N_14560);
nand UO_1473 (O_1473,N_14829,N_14521);
and UO_1474 (O_1474,N_14833,N_14658);
and UO_1475 (O_1475,N_14540,N_14929);
or UO_1476 (O_1476,N_14893,N_14616);
and UO_1477 (O_1477,N_14770,N_14961);
and UO_1478 (O_1478,N_14879,N_14504);
or UO_1479 (O_1479,N_14799,N_14779);
nor UO_1480 (O_1480,N_14611,N_14913);
nand UO_1481 (O_1481,N_14579,N_14972);
nor UO_1482 (O_1482,N_14807,N_14866);
nand UO_1483 (O_1483,N_14511,N_14757);
or UO_1484 (O_1484,N_14636,N_14998);
or UO_1485 (O_1485,N_14968,N_14820);
nand UO_1486 (O_1486,N_14593,N_14587);
nand UO_1487 (O_1487,N_14835,N_14788);
or UO_1488 (O_1488,N_14726,N_14795);
nand UO_1489 (O_1489,N_14541,N_14844);
nand UO_1490 (O_1490,N_14852,N_14826);
nor UO_1491 (O_1491,N_14647,N_14756);
or UO_1492 (O_1492,N_14594,N_14526);
xnor UO_1493 (O_1493,N_14941,N_14810);
xor UO_1494 (O_1494,N_14938,N_14855);
nor UO_1495 (O_1495,N_14985,N_14762);
xnor UO_1496 (O_1496,N_14775,N_14789);
nand UO_1497 (O_1497,N_14615,N_14660);
or UO_1498 (O_1498,N_14716,N_14583);
nor UO_1499 (O_1499,N_14569,N_14589);
nor UO_1500 (O_1500,N_14636,N_14832);
or UO_1501 (O_1501,N_14784,N_14749);
nor UO_1502 (O_1502,N_14517,N_14947);
nand UO_1503 (O_1503,N_14859,N_14782);
and UO_1504 (O_1504,N_14735,N_14822);
nand UO_1505 (O_1505,N_14590,N_14732);
and UO_1506 (O_1506,N_14826,N_14745);
and UO_1507 (O_1507,N_14921,N_14688);
nor UO_1508 (O_1508,N_14704,N_14823);
nand UO_1509 (O_1509,N_14811,N_14660);
nor UO_1510 (O_1510,N_14660,N_14629);
xnor UO_1511 (O_1511,N_14850,N_14728);
nor UO_1512 (O_1512,N_14515,N_14743);
xor UO_1513 (O_1513,N_14681,N_14771);
and UO_1514 (O_1514,N_14724,N_14523);
xnor UO_1515 (O_1515,N_14803,N_14880);
nand UO_1516 (O_1516,N_14705,N_14858);
nand UO_1517 (O_1517,N_14902,N_14860);
or UO_1518 (O_1518,N_14640,N_14685);
xor UO_1519 (O_1519,N_14941,N_14522);
or UO_1520 (O_1520,N_14547,N_14534);
nand UO_1521 (O_1521,N_14567,N_14764);
and UO_1522 (O_1522,N_14828,N_14841);
and UO_1523 (O_1523,N_14574,N_14501);
nand UO_1524 (O_1524,N_14886,N_14878);
and UO_1525 (O_1525,N_14910,N_14903);
nor UO_1526 (O_1526,N_14573,N_14585);
nor UO_1527 (O_1527,N_14832,N_14964);
or UO_1528 (O_1528,N_14810,N_14660);
or UO_1529 (O_1529,N_14531,N_14666);
nor UO_1530 (O_1530,N_14905,N_14667);
and UO_1531 (O_1531,N_14731,N_14669);
xor UO_1532 (O_1532,N_14534,N_14655);
nor UO_1533 (O_1533,N_14834,N_14893);
nand UO_1534 (O_1534,N_14785,N_14889);
nor UO_1535 (O_1535,N_14777,N_14694);
nor UO_1536 (O_1536,N_14709,N_14737);
or UO_1537 (O_1537,N_14790,N_14550);
xnor UO_1538 (O_1538,N_14573,N_14690);
nor UO_1539 (O_1539,N_14899,N_14520);
nand UO_1540 (O_1540,N_14918,N_14551);
xor UO_1541 (O_1541,N_14990,N_14752);
xnor UO_1542 (O_1542,N_14855,N_14921);
xor UO_1543 (O_1543,N_14651,N_14980);
nor UO_1544 (O_1544,N_14538,N_14902);
and UO_1545 (O_1545,N_14780,N_14864);
xor UO_1546 (O_1546,N_14813,N_14591);
xor UO_1547 (O_1547,N_14707,N_14557);
and UO_1548 (O_1548,N_14512,N_14570);
and UO_1549 (O_1549,N_14786,N_14709);
nand UO_1550 (O_1550,N_14900,N_14916);
and UO_1551 (O_1551,N_14884,N_14617);
nor UO_1552 (O_1552,N_14771,N_14918);
and UO_1553 (O_1553,N_14795,N_14975);
or UO_1554 (O_1554,N_14874,N_14863);
and UO_1555 (O_1555,N_14785,N_14717);
nor UO_1556 (O_1556,N_14748,N_14880);
or UO_1557 (O_1557,N_14843,N_14571);
and UO_1558 (O_1558,N_14914,N_14730);
or UO_1559 (O_1559,N_14609,N_14560);
nand UO_1560 (O_1560,N_14845,N_14983);
nor UO_1561 (O_1561,N_14769,N_14615);
or UO_1562 (O_1562,N_14738,N_14544);
or UO_1563 (O_1563,N_14689,N_14796);
nor UO_1564 (O_1564,N_14571,N_14945);
xnor UO_1565 (O_1565,N_14928,N_14670);
nor UO_1566 (O_1566,N_14564,N_14566);
and UO_1567 (O_1567,N_14997,N_14736);
or UO_1568 (O_1568,N_14638,N_14691);
nand UO_1569 (O_1569,N_14571,N_14693);
or UO_1570 (O_1570,N_14843,N_14875);
and UO_1571 (O_1571,N_14836,N_14595);
nor UO_1572 (O_1572,N_14852,N_14775);
nand UO_1573 (O_1573,N_14656,N_14574);
nor UO_1574 (O_1574,N_14816,N_14524);
and UO_1575 (O_1575,N_14547,N_14715);
nand UO_1576 (O_1576,N_14736,N_14956);
nand UO_1577 (O_1577,N_14853,N_14964);
and UO_1578 (O_1578,N_14694,N_14721);
or UO_1579 (O_1579,N_14846,N_14966);
or UO_1580 (O_1580,N_14682,N_14945);
or UO_1581 (O_1581,N_14602,N_14764);
or UO_1582 (O_1582,N_14587,N_14864);
and UO_1583 (O_1583,N_14530,N_14862);
nand UO_1584 (O_1584,N_14597,N_14618);
and UO_1585 (O_1585,N_14783,N_14628);
nand UO_1586 (O_1586,N_14833,N_14594);
or UO_1587 (O_1587,N_14853,N_14938);
xor UO_1588 (O_1588,N_14619,N_14899);
nand UO_1589 (O_1589,N_14891,N_14519);
or UO_1590 (O_1590,N_14881,N_14599);
xor UO_1591 (O_1591,N_14656,N_14716);
nand UO_1592 (O_1592,N_14795,N_14800);
nand UO_1593 (O_1593,N_14740,N_14756);
nand UO_1594 (O_1594,N_14654,N_14898);
nor UO_1595 (O_1595,N_14856,N_14885);
nor UO_1596 (O_1596,N_14853,N_14573);
and UO_1597 (O_1597,N_14988,N_14604);
and UO_1598 (O_1598,N_14658,N_14923);
xnor UO_1599 (O_1599,N_14732,N_14564);
or UO_1600 (O_1600,N_14901,N_14777);
and UO_1601 (O_1601,N_14807,N_14697);
nand UO_1602 (O_1602,N_14922,N_14892);
nor UO_1603 (O_1603,N_14886,N_14893);
xor UO_1604 (O_1604,N_14989,N_14954);
xor UO_1605 (O_1605,N_14511,N_14521);
nand UO_1606 (O_1606,N_14974,N_14795);
nor UO_1607 (O_1607,N_14982,N_14693);
nor UO_1608 (O_1608,N_14932,N_14979);
nand UO_1609 (O_1609,N_14534,N_14981);
or UO_1610 (O_1610,N_14742,N_14850);
nand UO_1611 (O_1611,N_14958,N_14533);
or UO_1612 (O_1612,N_14901,N_14641);
nor UO_1613 (O_1613,N_14685,N_14610);
nor UO_1614 (O_1614,N_14996,N_14726);
nor UO_1615 (O_1615,N_14771,N_14839);
or UO_1616 (O_1616,N_14593,N_14688);
nor UO_1617 (O_1617,N_14551,N_14812);
nor UO_1618 (O_1618,N_14666,N_14707);
xor UO_1619 (O_1619,N_14523,N_14885);
or UO_1620 (O_1620,N_14772,N_14616);
or UO_1621 (O_1621,N_14992,N_14720);
xnor UO_1622 (O_1622,N_14884,N_14933);
or UO_1623 (O_1623,N_14886,N_14618);
xor UO_1624 (O_1624,N_14772,N_14691);
and UO_1625 (O_1625,N_14721,N_14645);
or UO_1626 (O_1626,N_14542,N_14757);
or UO_1627 (O_1627,N_14728,N_14787);
nand UO_1628 (O_1628,N_14952,N_14660);
nand UO_1629 (O_1629,N_14713,N_14796);
xnor UO_1630 (O_1630,N_14500,N_14670);
nor UO_1631 (O_1631,N_14972,N_14539);
xnor UO_1632 (O_1632,N_14824,N_14769);
xor UO_1633 (O_1633,N_14804,N_14814);
nor UO_1634 (O_1634,N_14927,N_14512);
and UO_1635 (O_1635,N_14510,N_14626);
or UO_1636 (O_1636,N_14596,N_14955);
and UO_1637 (O_1637,N_14522,N_14924);
and UO_1638 (O_1638,N_14663,N_14876);
nor UO_1639 (O_1639,N_14895,N_14644);
and UO_1640 (O_1640,N_14715,N_14563);
or UO_1641 (O_1641,N_14747,N_14651);
or UO_1642 (O_1642,N_14898,N_14689);
nand UO_1643 (O_1643,N_14996,N_14916);
or UO_1644 (O_1644,N_14882,N_14706);
nor UO_1645 (O_1645,N_14532,N_14743);
or UO_1646 (O_1646,N_14678,N_14953);
nor UO_1647 (O_1647,N_14823,N_14714);
or UO_1648 (O_1648,N_14712,N_14663);
or UO_1649 (O_1649,N_14770,N_14805);
nand UO_1650 (O_1650,N_14947,N_14937);
and UO_1651 (O_1651,N_14948,N_14525);
nor UO_1652 (O_1652,N_14903,N_14565);
nand UO_1653 (O_1653,N_14519,N_14879);
nor UO_1654 (O_1654,N_14971,N_14870);
and UO_1655 (O_1655,N_14808,N_14650);
nor UO_1656 (O_1656,N_14677,N_14981);
nand UO_1657 (O_1657,N_14940,N_14559);
xor UO_1658 (O_1658,N_14963,N_14697);
or UO_1659 (O_1659,N_14645,N_14710);
xor UO_1660 (O_1660,N_14941,N_14699);
xnor UO_1661 (O_1661,N_14593,N_14935);
and UO_1662 (O_1662,N_14959,N_14600);
nand UO_1663 (O_1663,N_14974,N_14965);
or UO_1664 (O_1664,N_14763,N_14580);
nor UO_1665 (O_1665,N_14754,N_14501);
or UO_1666 (O_1666,N_14903,N_14539);
xnor UO_1667 (O_1667,N_14528,N_14813);
xnor UO_1668 (O_1668,N_14862,N_14868);
and UO_1669 (O_1669,N_14826,N_14948);
xnor UO_1670 (O_1670,N_14543,N_14567);
or UO_1671 (O_1671,N_14804,N_14778);
and UO_1672 (O_1672,N_14863,N_14606);
and UO_1673 (O_1673,N_14649,N_14648);
and UO_1674 (O_1674,N_14508,N_14752);
and UO_1675 (O_1675,N_14572,N_14749);
nand UO_1676 (O_1676,N_14618,N_14907);
nor UO_1677 (O_1677,N_14984,N_14891);
xnor UO_1678 (O_1678,N_14535,N_14993);
nand UO_1679 (O_1679,N_14906,N_14522);
xnor UO_1680 (O_1680,N_14909,N_14667);
or UO_1681 (O_1681,N_14670,N_14919);
nand UO_1682 (O_1682,N_14998,N_14649);
nand UO_1683 (O_1683,N_14707,N_14723);
or UO_1684 (O_1684,N_14524,N_14696);
nor UO_1685 (O_1685,N_14663,N_14690);
and UO_1686 (O_1686,N_14860,N_14534);
nand UO_1687 (O_1687,N_14761,N_14503);
nor UO_1688 (O_1688,N_14780,N_14924);
and UO_1689 (O_1689,N_14856,N_14940);
xor UO_1690 (O_1690,N_14971,N_14948);
or UO_1691 (O_1691,N_14543,N_14864);
and UO_1692 (O_1692,N_14665,N_14982);
nand UO_1693 (O_1693,N_14787,N_14932);
nor UO_1694 (O_1694,N_14643,N_14720);
nand UO_1695 (O_1695,N_14725,N_14866);
and UO_1696 (O_1696,N_14973,N_14962);
and UO_1697 (O_1697,N_14871,N_14991);
nor UO_1698 (O_1698,N_14760,N_14810);
nand UO_1699 (O_1699,N_14628,N_14708);
nand UO_1700 (O_1700,N_14989,N_14788);
nand UO_1701 (O_1701,N_14744,N_14957);
or UO_1702 (O_1702,N_14716,N_14825);
or UO_1703 (O_1703,N_14892,N_14708);
nor UO_1704 (O_1704,N_14655,N_14501);
xor UO_1705 (O_1705,N_14873,N_14628);
nor UO_1706 (O_1706,N_14689,N_14916);
or UO_1707 (O_1707,N_14575,N_14845);
nor UO_1708 (O_1708,N_14539,N_14559);
or UO_1709 (O_1709,N_14799,N_14817);
or UO_1710 (O_1710,N_14542,N_14780);
and UO_1711 (O_1711,N_14852,N_14823);
and UO_1712 (O_1712,N_14790,N_14715);
or UO_1713 (O_1713,N_14512,N_14943);
and UO_1714 (O_1714,N_14647,N_14563);
or UO_1715 (O_1715,N_14537,N_14690);
xnor UO_1716 (O_1716,N_14875,N_14835);
nor UO_1717 (O_1717,N_14904,N_14684);
xnor UO_1718 (O_1718,N_14635,N_14518);
xnor UO_1719 (O_1719,N_14939,N_14953);
xor UO_1720 (O_1720,N_14568,N_14784);
nor UO_1721 (O_1721,N_14547,N_14907);
nor UO_1722 (O_1722,N_14500,N_14537);
nand UO_1723 (O_1723,N_14985,N_14987);
xnor UO_1724 (O_1724,N_14690,N_14832);
or UO_1725 (O_1725,N_14893,N_14829);
nand UO_1726 (O_1726,N_14857,N_14661);
nand UO_1727 (O_1727,N_14618,N_14650);
nor UO_1728 (O_1728,N_14978,N_14788);
nor UO_1729 (O_1729,N_14730,N_14678);
nor UO_1730 (O_1730,N_14707,N_14623);
nand UO_1731 (O_1731,N_14746,N_14659);
and UO_1732 (O_1732,N_14694,N_14555);
xor UO_1733 (O_1733,N_14868,N_14859);
nand UO_1734 (O_1734,N_14890,N_14633);
or UO_1735 (O_1735,N_14712,N_14583);
nand UO_1736 (O_1736,N_14585,N_14892);
or UO_1737 (O_1737,N_14894,N_14878);
or UO_1738 (O_1738,N_14564,N_14899);
or UO_1739 (O_1739,N_14559,N_14713);
nand UO_1740 (O_1740,N_14828,N_14997);
xor UO_1741 (O_1741,N_14863,N_14585);
or UO_1742 (O_1742,N_14736,N_14570);
and UO_1743 (O_1743,N_14832,N_14909);
nor UO_1744 (O_1744,N_14507,N_14736);
nor UO_1745 (O_1745,N_14700,N_14788);
nand UO_1746 (O_1746,N_14522,N_14730);
and UO_1747 (O_1747,N_14529,N_14876);
nor UO_1748 (O_1748,N_14661,N_14559);
nand UO_1749 (O_1749,N_14783,N_14594);
nor UO_1750 (O_1750,N_14611,N_14782);
xor UO_1751 (O_1751,N_14653,N_14710);
or UO_1752 (O_1752,N_14768,N_14959);
nand UO_1753 (O_1753,N_14893,N_14583);
xnor UO_1754 (O_1754,N_14662,N_14836);
xor UO_1755 (O_1755,N_14506,N_14927);
xor UO_1756 (O_1756,N_14549,N_14737);
xor UO_1757 (O_1757,N_14736,N_14610);
or UO_1758 (O_1758,N_14697,N_14844);
and UO_1759 (O_1759,N_14589,N_14738);
nand UO_1760 (O_1760,N_14862,N_14999);
and UO_1761 (O_1761,N_14847,N_14582);
or UO_1762 (O_1762,N_14797,N_14622);
and UO_1763 (O_1763,N_14859,N_14679);
and UO_1764 (O_1764,N_14613,N_14583);
and UO_1765 (O_1765,N_14963,N_14861);
and UO_1766 (O_1766,N_14502,N_14749);
nand UO_1767 (O_1767,N_14976,N_14567);
and UO_1768 (O_1768,N_14947,N_14806);
or UO_1769 (O_1769,N_14552,N_14791);
nor UO_1770 (O_1770,N_14938,N_14820);
nand UO_1771 (O_1771,N_14575,N_14535);
nand UO_1772 (O_1772,N_14967,N_14561);
xnor UO_1773 (O_1773,N_14671,N_14897);
or UO_1774 (O_1774,N_14953,N_14698);
nor UO_1775 (O_1775,N_14730,N_14547);
or UO_1776 (O_1776,N_14566,N_14626);
xnor UO_1777 (O_1777,N_14745,N_14914);
nor UO_1778 (O_1778,N_14737,N_14656);
and UO_1779 (O_1779,N_14774,N_14933);
nand UO_1780 (O_1780,N_14979,N_14540);
and UO_1781 (O_1781,N_14825,N_14640);
and UO_1782 (O_1782,N_14503,N_14714);
or UO_1783 (O_1783,N_14655,N_14697);
and UO_1784 (O_1784,N_14616,N_14959);
nor UO_1785 (O_1785,N_14978,N_14895);
nand UO_1786 (O_1786,N_14666,N_14735);
nand UO_1787 (O_1787,N_14821,N_14976);
nand UO_1788 (O_1788,N_14618,N_14976);
nand UO_1789 (O_1789,N_14589,N_14915);
or UO_1790 (O_1790,N_14580,N_14723);
nand UO_1791 (O_1791,N_14715,N_14501);
and UO_1792 (O_1792,N_14506,N_14939);
or UO_1793 (O_1793,N_14643,N_14821);
and UO_1794 (O_1794,N_14783,N_14604);
or UO_1795 (O_1795,N_14513,N_14680);
nor UO_1796 (O_1796,N_14858,N_14648);
nand UO_1797 (O_1797,N_14689,N_14743);
and UO_1798 (O_1798,N_14686,N_14551);
xor UO_1799 (O_1799,N_14992,N_14742);
or UO_1800 (O_1800,N_14836,N_14577);
or UO_1801 (O_1801,N_14716,N_14519);
or UO_1802 (O_1802,N_14912,N_14993);
nand UO_1803 (O_1803,N_14707,N_14559);
xor UO_1804 (O_1804,N_14919,N_14819);
nor UO_1805 (O_1805,N_14852,N_14605);
nand UO_1806 (O_1806,N_14677,N_14531);
and UO_1807 (O_1807,N_14980,N_14833);
and UO_1808 (O_1808,N_14801,N_14868);
nand UO_1809 (O_1809,N_14644,N_14917);
nand UO_1810 (O_1810,N_14684,N_14922);
nand UO_1811 (O_1811,N_14704,N_14600);
nand UO_1812 (O_1812,N_14708,N_14843);
nor UO_1813 (O_1813,N_14582,N_14964);
xor UO_1814 (O_1814,N_14561,N_14744);
or UO_1815 (O_1815,N_14835,N_14853);
and UO_1816 (O_1816,N_14823,N_14716);
nor UO_1817 (O_1817,N_14731,N_14989);
and UO_1818 (O_1818,N_14669,N_14514);
nand UO_1819 (O_1819,N_14874,N_14986);
xnor UO_1820 (O_1820,N_14939,N_14683);
and UO_1821 (O_1821,N_14897,N_14785);
or UO_1822 (O_1822,N_14930,N_14652);
xnor UO_1823 (O_1823,N_14878,N_14728);
or UO_1824 (O_1824,N_14553,N_14761);
nand UO_1825 (O_1825,N_14657,N_14534);
nand UO_1826 (O_1826,N_14900,N_14648);
nor UO_1827 (O_1827,N_14567,N_14861);
and UO_1828 (O_1828,N_14724,N_14891);
nand UO_1829 (O_1829,N_14683,N_14724);
xor UO_1830 (O_1830,N_14943,N_14750);
nand UO_1831 (O_1831,N_14771,N_14604);
or UO_1832 (O_1832,N_14684,N_14798);
and UO_1833 (O_1833,N_14772,N_14681);
xor UO_1834 (O_1834,N_14780,N_14903);
nor UO_1835 (O_1835,N_14716,N_14964);
nand UO_1836 (O_1836,N_14771,N_14818);
nor UO_1837 (O_1837,N_14837,N_14675);
nor UO_1838 (O_1838,N_14559,N_14902);
or UO_1839 (O_1839,N_14544,N_14649);
or UO_1840 (O_1840,N_14690,N_14903);
or UO_1841 (O_1841,N_14884,N_14921);
nor UO_1842 (O_1842,N_14685,N_14516);
and UO_1843 (O_1843,N_14677,N_14897);
nand UO_1844 (O_1844,N_14760,N_14574);
nor UO_1845 (O_1845,N_14687,N_14753);
nor UO_1846 (O_1846,N_14765,N_14730);
nand UO_1847 (O_1847,N_14571,N_14620);
and UO_1848 (O_1848,N_14989,N_14674);
and UO_1849 (O_1849,N_14613,N_14597);
xor UO_1850 (O_1850,N_14978,N_14956);
and UO_1851 (O_1851,N_14987,N_14903);
and UO_1852 (O_1852,N_14578,N_14674);
nand UO_1853 (O_1853,N_14964,N_14562);
xor UO_1854 (O_1854,N_14963,N_14884);
and UO_1855 (O_1855,N_14544,N_14560);
nor UO_1856 (O_1856,N_14989,N_14903);
or UO_1857 (O_1857,N_14577,N_14700);
or UO_1858 (O_1858,N_14865,N_14960);
xnor UO_1859 (O_1859,N_14600,N_14558);
nand UO_1860 (O_1860,N_14734,N_14881);
nor UO_1861 (O_1861,N_14720,N_14622);
and UO_1862 (O_1862,N_14991,N_14751);
or UO_1863 (O_1863,N_14811,N_14645);
xor UO_1864 (O_1864,N_14541,N_14852);
nand UO_1865 (O_1865,N_14540,N_14790);
xor UO_1866 (O_1866,N_14817,N_14823);
or UO_1867 (O_1867,N_14634,N_14605);
xor UO_1868 (O_1868,N_14811,N_14639);
xnor UO_1869 (O_1869,N_14753,N_14756);
nor UO_1870 (O_1870,N_14745,N_14626);
xnor UO_1871 (O_1871,N_14884,N_14931);
and UO_1872 (O_1872,N_14514,N_14924);
and UO_1873 (O_1873,N_14782,N_14873);
or UO_1874 (O_1874,N_14608,N_14594);
and UO_1875 (O_1875,N_14928,N_14827);
and UO_1876 (O_1876,N_14769,N_14927);
nand UO_1877 (O_1877,N_14672,N_14704);
or UO_1878 (O_1878,N_14801,N_14854);
or UO_1879 (O_1879,N_14714,N_14890);
nor UO_1880 (O_1880,N_14686,N_14641);
xor UO_1881 (O_1881,N_14916,N_14828);
nor UO_1882 (O_1882,N_14967,N_14666);
and UO_1883 (O_1883,N_14921,N_14961);
nor UO_1884 (O_1884,N_14901,N_14895);
xor UO_1885 (O_1885,N_14988,N_14735);
nor UO_1886 (O_1886,N_14571,N_14539);
nor UO_1887 (O_1887,N_14597,N_14834);
nor UO_1888 (O_1888,N_14880,N_14533);
or UO_1889 (O_1889,N_14508,N_14664);
or UO_1890 (O_1890,N_14827,N_14570);
and UO_1891 (O_1891,N_14967,N_14878);
xnor UO_1892 (O_1892,N_14554,N_14521);
or UO_1893 (O_1893,N_14983,N_14980);
nand UO_1894 (O_1894,N_14892,N_14972);
nor UO_1895 (O_1895,N_14597,N_14548);
nand UO_1896 (O_1896,N_14689,N_14713);
nand UO_1897 (O_1897,N_14962,N_14618);
and UO_1898 (O_1898,N_14547,N_14522);
nor UO_1899 (O_1899,N_14987,N_14868);
xnor UO_1900 (O_1900,N_14642,N_14712);
xnor UO_1901 (O_1901,N_14686,N_14500);
xor UO_1902 (O_1902,N_14793,N_14828);
and UO_1903 (O_1903,N_14524,N_14857);
xor UO_1904 (O_1904,N_14862,N_14909);
or UO_1905 (O_1905,N_14870,N_14896);
nand UO_1906 (O_1906,N_14988,N_14624);
nor UO_1907 (O_1907,N_14664,N_14580);
nand UO_1908 (O_1908,N_14952,N_14572);
xnor UO_1909 (O_1909,N_14988,N_14585);
nor UO_1910 (O_1910,N_14704,N_14536);
nand UO_1911 (O_1911,N_14773,N_14669);
and UO_1912 (O_1912,N_14719,N_14987);
and UO_1913 (O_1913,N_14820,N_14652);
or UO_1914 (O_1914,N_14546,N_14737);
and UO_1915 (O_1915,N_14722,N_14879);
nor UO_1916 (O_1916,N_14978,N_14719);
xor UO_1917 (O_1917,N_14596,N_14674);
nand UO_1918 (O_1918,N_14848,N_14822);
nor UO_1919 (O_1919,N_14846,N_14701);
or UO_1920 (O_1920,N_14615,N_14670);
xor UO_1921 (O_1921,N_14921,N_14863);
nand UO_1922 (O_1922,N_14829,N_14707);
nand UO_1923 (O_1923,N_14513,N_14856);
and UO_1924 (O_1924,N_14526,N_14784);
xor UO_1925 (O_1925,N_14929,N_14821);
xor UO_1926 (O_1926,N_14900,N_14806);
nand UO_1927 (O_1927,N_14786,N_14609);
or UO_1928 (O_1928,N_14505,N_14703);
or UO_1929 (O_1929,N_14623,N_14555);
and UO_1930 (O_1930,N_14673,N_14765);
nor UO_1931 (O_1931,N_14832,N_14841);
and UO_1932 (O_1932,N_14951,N_14863);
and UO_1933 (O_1933,N_14747,N_14681);
nor UO_1934 (O_1934,N_14615,N_14622);
nand UO_1935 (O_1935,N_14520,N_14713);
xor UO_1936 (O_1936,N_14576,N_14642);
nand UO_1937 (O_1937,N_14864,N_14575);
nor UO_1938 (O_1938,N_14717,N_14562);
nand UO_1939 (O_1939,N_14525,N_14603);
nor UO_1940 (O_1940,N_14773,N_14884);
and UO_1941 (O_1941,N_14842,N_14556);
or UO_1942 (O_1942,N_14788,N_14742);
nand UO_1943 (O_1943,N_14636,N_14837);
nor UO_1944 (O_1944,N_14774,N_14545);
or UO_1945 (O_1945,N_14848,N_14890);
nand UO_1946 (O_1946,N_14571,N_14701);
and UO_1947 (O_1947,N_14980,N_14577);
xor UO_1948 (O_1948,N_14725,N_14706);
and UO_1949 (O_1949,N_14644,N_14972);
nor UO_1950 (O_1950,N_14756,N_14689);
xor UO_1951 (O_1951,N_14894,N_14862);
nor UO_1952 (O_1952,N_14811,N_14534);
nand UO_1953 (O_1953,N_14949,N_14605);
or UO_1954 (O_1954,N_14608,N_14695);
and UO_1955 (O_1955,N_14837,N_14592);
xnor UO_1956 (O_1956,N_14655,N_14897);
xnor UO_1957 (O_1957,N_14616,N_14697);
xnor UO_1958 (O_1958,N_14592,N_14602);
and UO_1959 (O_1959,N_14529,N_14735);
xnor UO_1960 (O_1960,N_14530,N_14810);
nor UO_1961 (O_1961,N_14605,N_14514);
and UO_1962 (O_1962,N_14788,N_14527);
xor UO_1963 (O_1963,N_14657,N_14834);
or UO_1964 (O_1964,N_14795,N_14926);
xnor UO_1965 (O_1965,N_14736,N_14757);
xnor UO_1966 (O_1966,N_14900,N_14833);
or UO_1967 (O_1967,N_14566,N_14843);
and UO_1968 (O_1968,N_14716,N_14881);
xor UO_1969 (O_1969,N_14521,N_14831);
or UO_1970 (O_1970,N_14814,N_14616);
or UO_1971 (O_1971,N_14988,N_14646);
nor UO_1972 (O_1972,N_14525,N_14521);
nor UO_1973 (O_1973,N_14877,N_14601);
nor UO_1974 (O_1974,N_14670,N_14899);
or UO_1975 (O_1975,N_14977,N_14795);
and UO_1976 (O_1976,N_14980,N_14535);
or UO_1977 (O_1977,N_14783,N_14600);
and UO_1978 (O_1978,N_14610,N_14524);
or UO_1979 (O_1979,N_14511,N_14564);
and UO_1980 (O_1980,N_14961,N_14634);
and UO_1981 (O_1981,N_14723,N_14542);
nand UO_1982 (O_1982,N_14709,N_14858);
nor UO_1983 (O_1983,N_14623,N_14824);
and UO_1984 (O_1984,N_14596,N_14834);
nor UO_1985 (O_1985,N_14564,N_14922);
or UO_1986 (O_1986,N_14742,N_14818);
nor UO_1987 (O_1987,N_14787,N_14670);
nor UO_1988 (O_1988,N_14669,N_14925);
nor UO_1989 (O_1989,N_14861,N_14830);
xor UO_1990 (O_1990,N_14995,N_14683);
xnor UO_1991 (O_1991,N_14931,N_14919);
or UO_1992 (O_1992,N_14574,N_14560);
nand UO_1993 (O_1993,N_14690,N_14697);
or UO_1994 (O_1994,N_14600,N_14966);
xnor UO_1995 (O_1995,N_14659,N_14641);
nor UO_1996 (O_1996,N_14637,N_14902);
and UO_1997 (O_1997,N_14792,N_14887);
nand UO_1998 (O_1998,N_14675,N_14938);
nand UO_1999 (O_1999,N_14589,N_14951);
endmodule