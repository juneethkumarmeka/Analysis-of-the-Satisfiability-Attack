module basic_500_3000_500_40_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xnor U0 (N_0,In_128,In_373);
nand U1 (N_1,In_33,In_147);
xor U2 (N_2,In_87,In_228);
nand U3 (N_3,In_378,In_192);
nand U4 (N_4,In_264,In_369);
nand U5 (N_5,In_32,In_55);
nand U6 (N_6,In_148,In_296);
nor U7 (N_7,In_453,In_115);
nor U8 (N_8,In_72,In_411);
nor U9 (N_9,In_393,In_387);
xnor U10 (N_10,In_493,In_27);
nor U11 (N_11,In_259,In_97);
and U12 (N_12,In_391,In_90);
nor U13 (N_13,In_281,In_421);
xor U14 (N_14,In_237,In_120);
xor U15 (N_15,In_386,In_69);
nand U16 (N_16,In_63,In_133);
xnor U17 (N_17,In_137,In_64);
nor U18 (N_18,In_82,In_336);
nor U19 (N_19,In_68,In_436);
xor U20 (N_20,In_494,In_103);
or U21 (N_21,In_301,In_451);
nand U22 (N_22,In_257,In_440);
or U23 (N_23,In_230,In_92);
or U24 (N_24,In_350,In_116);
nor U25 (N_25,In_160,In_40);
xnor U26 (N_26,In_271,In_111);
nor U27 (N_27,In_498,In_225);
or U28 (N_28,In_142,In_42);
xor U29 (N_29,In_61,In_420);
nor U30 (N_30,In_96,In_323);
nand U31 (N_31,In_52,In_374);
or U32 (N_32,In_191,In_222);
xnor U33 (N_33,In_246,In_452);
or U34 (N_34,In_5,In_140);
or U35 (N_35,In_57,In_18);
xnor U36 (N_36,In_499,In_149);
xnor U37 (N_37,In_292,In_73);
or U38 (N_38,In_270,In_445);
nor U39 (N_39,In_408,In_180);
xnor U40 (N_40,In_241,In_477);
or U41 (N_41,In_242,In_278);
xnor U42 (N_42,In_331,In_168);
and U43 (N_43,In_200,In_125);
xor U44 (N_44,In_434,In_474);
nand U45 (N_45,In_287,In_211);
nor U46 (N_46,In_199,In_272);
and U47 (N_47,In_54,In_483);
nor U48 (N_48,In_173,In_299);
and U49 (N_49,In_330,In_233);
and U50 (N_50,In_41,In_256);
nand U51 (N_51,In_203,In_406);
or U52 (N_52,In_495,In_85);
nor U53 (N_53,In_457,In_24);
xor U54 (N_54,In_370,In_51);
or U55 (N_55,In_353,In_315);
and U56 (N_56,In_109,In_9);
xnor U57 (N_57,In_439,In_465);
xnor U58 (N_58,In_482,In_107);
or U59 (N_59,In_244,In_260);
nor U60 (N_60,In_213,In_23);
nor U61 (N_61,In_352,In_255);
nor U62 (N_62,In_60,In_108);
xor U63 (N_63,In_417,In_265);
xor U64 (N_64,In_295,In_380);
nor U65 (N_65,In_306,In_45);
and U66 (N_66,In_124,In_189);
or U67 (N_67,In_321,In_314);
or U68 (N_68,In_332,In_14);
and U69 (N_69,In_119,In_384);
nor U70 (N_70,In_470,In_223);
nand U71 (N_71,In_433,In_58);
xnor U72 (N_72,In_39,In_50);
xnor U73 (N_73,In_358,In_235);
or U74 (N_74,In_98,In_162);
nor U75 (N_75,In_139,In_8);
or U76 (N_76,In_74,In_206);
nor U77 (N_77,In_100,N_65);
nor U78 (N_78,In_201,In_95);
xor U79 (N_79,N_51,In_334);
nor U80 (N_80,N_11,In_151);
and U81 (N_81,N_21,In_153);
nor U82 (N_82,In_335,In_489);
xnor U83 (N_83,In_79,In_447);
or U84 (N_84,In_398,In_431);
or U85 (N_85,In_15,In_490);
xor U86 (N_86,In_428,In_280);
nand U87 (N_87,In_170,In_480);
and U88 (N_88,In_44,In_416);
nand U89 (N_89,In_460,In_266);
xnor U90 (N_90,In_413,In_132);
or U91 (N_91,N_2,N_26);
xnor U92 (N_92,In_34,In_469);
nand U93 (N_93,In_487,In_478);
nand U94 (N_94,N_31,In_214);
xnor U95 (N_95,N_57,In_123);
xor U96 (N_96,In_190,In_443);
or U97 (N_97,N_55,In_19);
and U98 (N_98,In_12,In_348);
and U99 (N_99,N_28,In_365);
nor U100 (N_100,In_67,In_224);
and U101 (N_101,In_106,N_14);
and U102 (N_102,In_193,In_276);
nand U103 (N_103,N_7,In_466);
nor U104 (N_104,N_29,In_438);
xnor U105 (N_105,N_6,In_59);
xnor U106 (N_106,In_36,In_158);
nand U107 (N_107,In_220,In_53);
xnor U108 (N_108,In_227,In_178);
and U109 (N_109,In_194,N_8);
xor U110 (N_110,In_360,In_426);
nor U111 (N_111,In_375,In_282);
nor U112 (N_112,In_368,N_50);
and U113 (N_113,In_185,N_13);
nor U114 (N_114,In_117,In_383);
or U115 (N_115,N_53,N_9);
nor U116 (N_116,In_243,In_319);
nor U117 (N_117,In_449,In_28);
xnor U118 (N_118,N_56,N_34);
nand U119 (N_119,N_35,In_273);
xor U120 (N_120,In_175,In_361);
nor U121 (N_121,In_435,In_268);
or U122 (N_122,In_134,In_46);
nor U123 (N_123,In_432,In_410);
xnor U124 (N_124,In_293,In_208);
or U125 (N_125,N_37,N_36);
and U126 (N_126,In_309,In_164);
or U127 (N_127,In_186,In_250);
or U128 (N_128,In_56,In_485);
and U129 (N_129,In_359,In_357);
nand U130 (N_130,In_113,In_71);
xnor U131 (N_131,In_157,In_1);
nand U132 (N_132,In_121,In_130);
or U133 (N_133,In_83,In_300);
nor U134 (N_134,N_47,N_33);
nand U135 (N_135,In_218,In_342);
and U136 (N_136,In_392,In_401);
xor U137 (N_137,In_379,In_89);
and U138 (N_138,In_204,In_135);
or U139 (N_139,N_59,In_349);
and U140 (N_140,In_471,N_68);
or U141 (N_141,N_15,N_58);
or U142 (N_142,In_283,N_19);
or U143 (N_143,N_67,In_333);
and U144 (N_144,In_455,In_364);
or U145 (N_145,In_422,In_475);
nor U146 (N_146,N_74,In_326);
nand U147 (N_147,In_88,In_345);
nor U148 (N_148,In_394,In_0);
or U149 (N_149,In_16,In_167);
nand U150 (N_150,In_254,N_122);
xor U151 (N_151,N_4,In_110);
or U152 (N_152,In_188,N_49);
nor U153 (N_153,N_38,N_78);
nor U154 (N_154,In_486,N_62);
or U155 (N_155,In_263,In_93);
nand U156 (N_156,In_169,In_207);
nor U157 (N_157,In_179,N_148);
or U158 (N_158,In_497,In_390);
and U159 (N_159,N_102,N_123);
nand U160 (N_160,In_86,N_119);
xnor U161 (N_161,N_121,In_341);
or U162 (N_162,N_147,In_138);
xor U163 (N_163,In_303,N_92);
nand U164 (N_164,N_133,N_125);
nor U165 (N_165,In_454,N_80);
nand U166 (N_166,N_120,N_142);
and U167 (N_167,N_100,N_5);
nand U168 (N_168,In_6,In_297);
xnor U169 (N_169,In_118,N_45);
xnor U170 (N_170,In_317,In_152);
nor U171 (N_171,In_7,In_318);
or U172 (N_172,N_22,N_61);
or U173 (N_173,N_1,N_24);
xor U174 (N_174,N_118,In_286);
and U175 (N_175,In_473,N_101);
nor U176 (N_176,N_73,In_363);
xnor U177 (N_177,N_71,In_253);
or U178 (N_178,In_320,In_31);
nor U179 (N_179,N_30,In_25);
nand U180 (N_180,In_4,In_404);
xnor U181 (N_181,In_251,N_104);
nor U182 (N_182,In_424,In_221);
nor U183 (N_183,In_366,In_462);
nor U184 (N_184,In_274,N_138);
and U185 (N_185,N_107,In_141);
and U186 (N_186,N_129,In_425);
or U187 (N_187,In_302,In_146);
and U188 (N_188,N_60,N_117);
xnor U189 (N_189,In_122,In_442);
nand U190 (N_190,In_182,In_418);
or U191 (N_191,N_109,In_187);
and U192 (N_192,In_381,In_239);
nor U193 (N_193,In_129,In_156);
and U194 (N_194,In_184,N_69);
nand U195 (N_195,In_104,In_430);
nand U196 (N_196,In_226,In_240);
nor U197 (N_197,In_150,In_62);
nand U198 (N_198,In_21,In_145);
xor U199 (N_199,In_84,In_252);
nand U200 (N_200,In_308,In_249);
and U201 (N_201,In_234,In_316);
and U202 (N_202,In_338,In_305);
xnor U203 (N_203,In_304,In_205);
or U204 (N_204,In_114,N_88);
and U205 (N_205,In_229,In_277);
and U206 (N_206,In_219,N_48);
or U207 (N_207,In_288,N_99);
or U208 (N_208,N_112,In_38);
or U209 (N_209,In_267,In_310);
nor U210 (N_210,In_144,N_110);
or U211 (N_211,In_126,N_135);
and U212 (N_212,In_202,In_80);
nand U213 (N_213,In_248,In_427);
and U214 (N_214,In_183,N_18);
and U215 (N_215,In_376,In_212);
and U216 (N_216,In_284,In_388);
xor U217 (N_217,N_105,N_63);
or U218 (N_218,N_97,In_399);
or U219 (N_219,In_351,N_39);
and U220 (N_220,N_41,N_96);
nand U221 (N_221,In_29,In_372);
and U222 (N_222,N_146,N_54);
and U223 (N_223,In_488,In_197);
nor U224 (N_224,In_367,N_81);
or U225 (N_225,N_166,N_159);
nand U226 (N_226,N_190,N_145);
nor U227 (N_227,In_395,N_215);
nor U228 (N_228,N_72,In_468);
nor U229 (N_229,N_152,In_419);
nand U230 (N_230,In_415,N_176);
nand U231 (N_231,In_101,In_481);
or U232 (N_232,In_347,N_77);
nor U233 (N_233,N_94,In_344);
nor U234 (N_234,In_414,In_231);
nand U235 (N_235,N_113,In_262);
nor U236 (N_236,N_179,In_195);
nand U237 (N_237,In_30,In_238);
xor U238 (N_238,In_405,In_312);
and U239 (N_239,N_207,In_20);
xnor U240 (N_240,In_423,N_126);
nor U241 (N_241,In_311,N_12);
nor U242 (N_242,N_43,In_491);
nand U243 (N_243,In_407,In_3);
nand U244 (N_244,N_134,N_20);
xor U245 (N_245,N_40,In_261);
nor U246 (N_246,N_75,In_385);
or U247 (N_247,In_81,N_17);
xnor U248 (N_248,In_397,N_211);
nor U249 (N_249,N_222,In_441);
nand U250 (N_250,N_116,N_66);
xnor U251 (N_251,In_328,In_294);
and U252 (N_252,N_91,In_371);
or U253 (N_253,In_289,N_206);
nor U254 (N_254,N_203,N_191);
and U255 (N_255,In_464,In_10);
xor U256 (N_256,In_216,N_204);
or U257 (N_257,N_124,N_175);
or U258 (N_258,In_26,In_143);
nor U259 (N_259,N_182,In_444);
nand U260 (N_260,In_131,In_76);
nand U261 (N_261,In_217,In_458);
xnor U262 (N_262,In_43,N_108);
xor U263 (N_263,N_177,In_35);
and U264 (N_264,N_184,N_136);
xnor U265 (N_265,N_141,In_389);
or U266 (N_266,N_87,In_13);
or U267 (N_267,In_11,N_76);
xnor U268 (N_268,N_115,In_496);
xor U269 (N_269,N_153,In_165);
xnor U270 (N_270,In_313,N_85);
and U271 (N_271,N_44,N_192);
nor U272 (N_272,In_461,N_188);
nand U273 (N_273,In_2,In_362);
and U274 (N_274,N_130,N_223);
xor U275 (N_275,In_91,In_409);
nand U276 (N_276,In_172,N_3);
and U277 (N_277,In_196,N_25);
xnor U278 (N_278,N_103,N_162);
nor U279 (N_279,In_154,In_322);
nand U280 (N_280,N_200,In_402);
xnor U281 (N_281,N_212,N_183);
nor U282 (N_282,N_155,In_339);
xor U283 (N_283,N_219,N_172);
or U284 (N_284,In_99,N_128);
xnor U285 (N_285,N_16,In_437);
nor U286 (N_286,N_178,In_479);
nor U287 (N_287,N_205,In_75);
or U288 (N_288,In_94,In_17);
or U289 (N_289,In_463,N_79);
nor U290 (N_290,In_177,N_165);
nor U291 (N_291,N_86,In_377);
nand U292 (N_292,In_400,N_98);
and U293 (N_293,N_82,N_195);
nand U294 (N_294,In_291,In_48);
nor U295 (N_295,N_185,N_27);
nand U296 (N_296,In_269,N_168);
or U297 (N_297,In_396,N_52);
nand U298 (N_298,N_89,N_171);
nor U299 (N_299,In_102,N_158);
or U300 (N_300,In_78,In_22);
nor U301 (N_301,N_298,N_280);
nor U302 (N_302,N_228,In_459);
nand U303 (N_303,In_198,N_278);
nand U304 (N_304,In_448,N_83);
nor U305 (N_305,In_181,In_476);
or U306 (N_306,In_472,N_248);
xnor U307 (N_307,N_231,N_95);
nor U308 (N_308,N_232,N_274);
and U309 (N_309,N_282,N_224);
xnor U310 (N_310,N_255,N_163);
nand U311 (N_311,N_229,N_169);
xnor U312 (N_312,N_249,N_244);
nor U313 (N_313,N_174,In_247);
nor U314 (N_314,N_139,N_10);
xor U315 (N_315,N_227,N_247);
and U316 (N_316,N_233,In_66);
nand U317 (N_317,N_281,N_289);
xnor U318 (N_318,N_199,N_268);
xor U319 (N_319,In_166,In_245);
nand U320 (N_320,In_285,N_217);
xnor U321 (N_321,N_149,N_161);
nand U322 (N_322,N_127,In_174);
or U323 (N_323,N_196,N_253);
or U324 (N_324,N_263,N_46);
nand U325 (N_325,N_32,In_467);
nor U326 (N_326,N_288,N_273);
and U327 (N_327,N_257,In_215);
or U328 (N_328,N_296,N_198);
nand U329 (N_329,N_234,N_201);
and U330 (N_330,N_164,In_65);
or U331 (N_331,N_271,N_210);
nor U332 (N_332,N_70,In_327);
nand U333 (N_333,In_446,In_232);
and U334 (N_334,In_429,N_230);
nand U335 (N_335,N_243,In_105);
nand U336 (N_336,N_214,N_180);
nor U337 (N_337,In_456,N_262);
nand U338 (N_338,N_154,In_37);
and U339 (N_339,N_173,In_275);
xnor U340 (N_340,In_403,N_221);
xor U341 (N_341,N_251,N_245);
nand U342 (N_342,N_237,N_239);
nand U343 (N_343,N_216,N_260);
nand U344 (N_344,In_324,N_167);
and U345 (N_345,N_272,In_112);
nor U346 (N_346,N_93,N_267);
and U347 (N_347,N_252,In_210);
nor U348 (N_348,In_159,In_279);
and U349 (N_349,In_176,N_235);
xor U350 (N_350,N_209,N_170);
or U351 (N_351,In_127,N_258);
or U352 (N_352,In_70,N_287);
or U353 (N_353,In_343,N_220);
and U354 (N_354,N_0,N_143);
nor U355 (N_355,N_140,N_84);
nor U356 (N_356,N_114,In_355);
or U357 (N_357,N_132,In_412);
xnor U358 (N_358,In_236,N_294);
xor U359 (N_359,N_156,N_160);
and U360 (N_360,N_279,N_186);
or U361 (N_361,In_163,In_258);
xor U362 (N_362,N_269,In_450);
or U363 (N_363,N_277,In_209);
nor U364 (N_364,In_346,N_266);
nor U365 (N_365,N_265,N_137);
xor U366 (N_366,N_90,N_261);
nor U367 (N_367,N_246,In_337);
xnor U368 (N_368,N_291,N_284);
nand U369 (N_369,N_240,N_187);
nand U370 (N_370,N_150,N_236);
or U371 (N_371,N_290,N_238);
xor U372 (N_372,N_275,In_49);
nor U373 (N_373,N_194,N_193);
nor U374 (N_374,N_286,N_197);
nand U375 (N_375,N_343,N_329);
nand U376 (N_376,In_171,N_335);
and U377 (N_377,In_382,N_361);
nor U378 (N_378,In_484,N_324);
or U379 (N_379,N_344,N_304);
nor U380 (N_380,In_307,N_226);
and U381 (N_381,N_320,N_42);
and U382 (N_382,N_208,N_131);
nor U383 (N_383,N_213,N_345);
and U384 (N_384,N_332,N_322);
nand U385 (N_385,N_301,N_317);
xnor U386 (N_386,N_225,N_357);
xnor U387 (N_387,N_305,N_370);
or U388 (N_388,N_325,N_347);
nor U389 (N_389,In_354,N_309);
xor U390 (N_390,N_368,N_339);
nor U391 (N_391,N_358,N_366);
xor U392 (N_392,N_365,N_372);
nor U393 (N_393,N_363,N_323);
nor U394 (N_394,N_356,N_374);
or U395 (N_395,N_315,N_106);
nor U396 (N_396,N_341,N_334);
and U397 (N_397,N_242,N_313);
xnor U398 (N_398,N_295,N_311);
xor U399 (N_399,N_337,N_349);
and U400 (N_400,N_264,N_111);
or U401 (N_401,N_151,N_285);
xnor U402 (N_402,N_328,N_307);
xnor U403 (N_403,N_23,N_299);
xor U404 (N_404,N_355,In_325);
or U405 (N_405,N_218,In_161);
nand U406 (N_406,N_189,N_327);
and U407 (N_407,N_292,N_373);
and U408 (N_408,N_318,In_356);
or U409 (N_409,N_293,In_77);
or U410 (N_410,N_371,In_492);
nor U411 (N_411,In_329,N_64);
xor U412 (N_412,In_155,N_310);
or U413 (N_413,In_290,N_353);
xnor U414 (N_414,N_340,N_316);
and U415 (N_415,N_348,N_256);
xor U416 (N_416,N_283,N_336);
nand U417 (N_417,N_331,N_302);
and U418 (N_418,N_351,N_359);
and U419 (N_419,N_326,N_202);
nand U420 (N_420,N_352,N_333);
xor U421 (N_421,In_340,N_276);
or U422 (N_422,N_354,N_300);
xnor U423 (N_423,N_350,N_250);
nor U424 (N_424,N_362,N_312);
nor U425 (N_425,N_338,N_330);
or U426 (N_426,N_254,N_319);
nand U427 (N_427,N_364,N_241);
or U428 (N_428,In_47,N_369);
and U429 (N_429,N_270,N_314);
and U430 (N_430,N_306,N_259);
xor U431 (N_431,N_308,N_157);
nor U432 (N_432,N_346,N_321);
xor U433 (N_433,N_181,N_144);
xnor U434 (N_434,N_367,N_342);
nand U435 (N_435,N_360,N_297);
nand U436 (N_436,N_303,In_136);
or U437 (N_437,In_298,In_47);
nand U438 (N_438,N_317,N_318);
xnor U439 (N_439,N_337,N_326);
nor U440 (N_440,N_313,N_361);
nor U441 (N_441,N_332,N_312);
nor U442 (N_442,In_155,N_350);
nor U443 (N_443,N_306,N_327);
or U444 (N_444,N_370,N_347);
nor U445 (N_445,N_270,N_302);
or U446 (N_446,N_213,N_374);
nor U447 (N_447,N_254,N_373);
nand U448 (N_448,In_484,N_352);
xnor U449 (N_449,N_344,N_360);
nor U450 (N_450,N_398,N_412);
xor U451 (N_451,N_409,N_406);
nand U452 (N_452,N_415,N_397);
and U453 (N_453,N_435,N_445);
nand U454 (N_454,N_441,N_416);
nor U455 (N_455,N_426,N_437);
and U456 (N_456,N_376,N_432);
and U457 (N_457,N_428,N_433);
nor U458 (N_458,N_417,N_449);
nor U459 (N_459,N_418,N_385);
xnor U460 (N_460,N_420,N_427);
and U461 (N_461,N_394,N_399);
and U462 (N_462,N_447,N_431);
nand U463 (N_463,N_422,N_379);
and U464 (N_464,N_381,N_410);
nor U465 (N_465,N_423,N_408);
xor U466 (N_466,N_442,N_434);
xor U467 (N_467,N_407,N_440);
or U468 (N_468,N_429,N_425);
xnor U469 (N_469,N_390,N_421);
nor U470 (N_470,N_401,N_382);
and U471 (N_471,N_391,N_395);
xnor U472 (N_472,N_419,N_377);
and U473 (N_473,N_400,N_443);
and U474 (N_474,N_413,N_446);
nand U475 (N_475,N_438,N_405);
nor U476 (N_476,N_430,N_388);
and U477 (N_477,N_448,N_411);
nor U478 (N_478,N_414,N_378);
nand U479 (N_479,N_436,N_380);
and U480 (N_480,N_383,N_375);
xor U481 (N_481,N_424,N_386);
xor U482 (N_482,N_403,N_444);
or U483 (N_483,N_392,N_393);
nand U484 (N_484,N_384,N_387);
or U485 (N_485,N_439,N_396);
nor U486 (N_486,N_389,N_402);
and U487 (N_487,N_404,N_440);
or U488 (N_488,N_381,N_398);
nand U489 (N_489,N_375,N_376);
and U490 (N_490,N_376,N_383);
xnor U491 (N_491,N_385,N_390);
nor U492 (N_492,N_431,N_410);
and U493 (N_493,N_409,N_423);
xor U494 (N_494,N_396,N_436);
xnor U495 (N_495,N_443,N_444);
nor U496 (N_496,N_384,N_411);
nor U497 (N_497,N_435,N_387);
and U498 (N_498,N_407,N_391);
or U499 (N_499,N_396,N_381);
xnor U500 (N_500,N_384,N_417);
nor U501 (N_501,N_421,N_402);
and U502 (N_502,N_397,N_391);
xnor U503 (N_503,N_406,N_408);
or U504 (N_504,N_403,N_424);
or U505 (N_505,N_424,N_430);
nor U506 (N_506,N_419,N_389);
xnor U507 (N_507,N_402,N_427);
or U508 (N_508,N_384,N_426);
nor U509 (N_509,N_438,N_385);
or U510 (N_510,N_415,N_404);
xor U511 (N_511,N_407,N_380);
nand U512 (N_512,N_383,N_413);
nand U513 (N_513,N_388,N_440);
xnor U514 (N_514,N_409,N_444);
xor U515 (N_515,N_440,N_394);
or U516 (N_516,N_379,N_380);
and U517 (N_517,N_401,N_444);
and U518 (N_518,N_440,N_424);
xnor U519 (N_519,N_383,N_389);
or U520 (N_520,N_418,N_381);
or U521 (N_521,N_441,N_445);
and U522 (N_522,N_404,N_375);
or U523 (N_523,N_394,N_442);
xor U524 (N_524,N_442,N_392);
and U525 (N_525,N_512,N_502);
and U526 (N_526,N_481,N_492);
nor U527 (N_527,N_511,N_467);
and U528 (N_528,N_454,N_465);
nor U529 (N_529,N_456,N_495);
and U530 (N_530,N_475,N_469);
nor U531 (N_531,N_509,N_516);
or U532 (N_532,N_472,N_484);
xor U533 (N_533,N_458,N_459);
and U534 (N_534,N_524,N_463);
nor U535 (N_535,N_471,N_500);
or U536 (N_536,N_494,N_470);
nand U537 (N_537,N_522,N_510);
and U538 (N_538,N_478,N_468);
or U539 (N_539,N_477,N_485);
nand U540 (N_540,N_473,N_480);
and U541 (N_541,N_507,N_457);
nor U542 (N_542,N_464,N_488);
xnor U543 (N_543,N_503,N_460);
or U544 (N_544,N_474,N_479);
nor U545 (N_545,N_519,N_493);
and U546 (N_546,N_515,N_499);
nand U547 (N_547,N_520,N_514);
nand U548 (N_548,N_498,N_486);
nor U549 (N_549,N_523,N_482);
and U550 (N_550,N_513,N_504);
nor U551 (N_551,N_476,N_450);
nand U552 (N_552,N_521,N_455);
xnor U553 (N_553,N_453,N_517);
and U554 (N_554,N_489,N_487);
nor U555 (N_555,N_491,N_461);
nand U556 (N_556,N_462,N_466);
and U557 (N_557,N_506,N_490);
or U558 (N_558,N_501,N_508);
and U559 (N_559,N_518,N_452);
nor U560 (N_560,N_483,N_505);
nand U561 (N_561,N_497,N_451);
xnor U562 (N_562,N_496,N_477);
nand U563 (N_563,N_484,N_489);
nor U564 (N_564,N_491,N_496);
xor U565 (N_565,N_480,N_482);
nor U566 (N_566,N_488,N_468);
or U567 (N_567,N_479,N_463);
xnor U568 (N_568,N_477,N_503);
nand U569 (N_569,N_520,N_495);
or U570 (N_570,N_515,N_477);
or U571 (N_571,N_493,N_516);
nor U572 (N_572,N_470,N_485);
and U573 (N_573,N_495,N_457);
xor U574 (N_574,N_454,N_522);
nand U575 (N_575,N_478,N_503);
xor U576 (N_576,N_502,N_505);
and U577 (N_577,N_458,N_490);
nand U578 (N_578,N_454,N_484);
and U579 (N_579,N_458,N_523);
or U580 (N_580,N_503,N_467);
nand U581 (N_581,N_454,N_475);
nor U582 (N_582,N_490,N_456);
nor U583 (N_583,N_474,N_482);
nor U584 (N_584,N_470,N_500);
and U585 (N_585,N_465,N_470);
nor U586 (N_586,N_458,N_491);
nand U587 (N_587,N_516,N_484);
and U588 (N_588,N_489,N_469);
or U589 (N_589,N_452,N_456);
nand U590 (N_590,N_460,N_510);
nand U591 (N_591,N_512,N_466);
or U592 (N_592,N_489,N_488);
nand U593 (N_593,N_464,N_469);
nand U594 (N_594,N_503,N_452);
xor U595 (N_595,N_500,N_518);
nand U596 (N_596,N_454,N_512);
and U597 (N_597,N_501,N_455);
and U598 (N_598,N_463,N_481);
or U599 (N_599,N_491,N_463);
or U600 (N_600,N_570,N_571);
nand U601 (N_601,N_527,N_582);
nor U602 (N_602,N_530,N_587);
or U603 (N_603,N_588,N_566);
xnor U604 (N_604,N_540,N_532);
nand U605 (N_605,N_565,N_558);
or U606 (N_606,N_564,N_529);
and U607 (N_607,N_591,N_545);
nand U608 (N_608,N_561,N_576);
nand U609 (N_609,N_555,N_551);
nand U610 (N_610,N_544,N_573);
nor U611 (N_611,N_554,N_550);
nor U612 (N_612,N_538,N_577);
and U613 (N_613,N_542,N_595);
xor U614 (N_614,N_539,N_560);
and U615 (N_615,N_528,N_568);
nor U616 (N_616,N_536,N_531);
and U617 (N_617,N_557,N_552);
and U618 (N_618,N_559,N_584);
nor U619 (N_619,N_526,N_567);
xnor U620 (N_620,N_543,N_574);
nor U621 (N_621,N_563,N_525);
or U622 (N_622,N_548,N_583);
and U623 (N_623,N_533,N_594);
nand U624 (N_624,N_589,N_586);
nand U625 (N_625,N_575,N_590);
or U626 (N_626,N_534,N_553);
and U627 (N_627,N_547,N_597);
or U628 (N_628,N_541,N_569);
nand U629 (N_629,N_549,N_578);
xnor U630 (N_630,N_580,N_599);
nand U631 (N_631,N_598,N_535);
nand U632 (N_632,N_596,N_556);
or U633 (N_633,N_593,N_562);
nand U634 (N_634,N_592,N_537);
xnor U635 (N_635,N_585,N_579);
nand U636 (N_636,N_572,N_546);
and U637 (N_637,N_581,N_572);
nand U638 (N_638,N_538,N_529);
or U639 (N_639,N_578,N_540);
xor U640 (N_640,N_579,N_567);
or U641 (N_641,N_534,N_583);
nor U642 (N_642,N_567,N_574);
xor U643 (N_643,N_568,N_592);
xor U644 (N_644,N_573,N_595);
or U645 (N_645,N_575,N_585);
or U646 (N_646,N_550,N_555);
nand U647 (N_647,N_587,N_533);
and U648 (N_648,N_586,N_578);
nand U649 (N_649,N_525,N_534);
or U650 (N_650,N_575,N_540);
and U651 (N_651,N_567,N_556);
xnor U652 (N_652,N_576,N_597);
or U653 (N_653,N_577,N_586);
nand U654 (N_654,N_548,N_590);
nand U655 (N_655,N_593,N_575);
or U656 (N_656,N_563,N_545);
or U657 (N_657,N_542,N_581);
nand U658 (N_658,N_577,N_539);
nand U659 (N_659,N_530,N_533);
and U660 (N_660,N_576,N_569);
or U661 (N_661,N_528,N_560);
nand U662 (N_662,N_558,N_586);
and U663 (N_663,N_543,N_562);
or U664 (N_664,N_566,N_592);
or U665 (N_665,N_537,N_554);
or U666 (N_666,N_540,N_549);
xnor U667 (N_667,N_596,N_553);
nor U668 (N_668,N_537,N_596);
nand U669 (N_669,N_556,N_554);
nor U670 (N_670,N_577,N_595);
or U671 (N_671,N_571,N_526);
or U672 (N_672,N_549,N_572);
or U673 (N_673,N_586,N_547);
xor U674 (N_674,N_565,N_569);
or U675 (N_675,N_633,N_671);
nand U676 (N_676,N_622,N_624);
and U677 (N_677,N_610,N_637);
and U678 (N_678,N_646,N_600);
nand U679 (N_679,N_657,N_616);
xor U680 (N_680,N_673,N_641);
and U681 (N_681,N_636,N_651);
nand U682 (N_682,N_644,N_647);
and U683 (N_683,N_652,N_669);
or U684 (N_684,N_623,N_649);
xnor U685 (N_685,N_629,N_605);
and U686 (N_686,N_620,N_604);
nor U687 (N_687,N_625,N_654);
nand U688 (N_688,N_602,N_603);
xnor U689 (N_689,N_614,N_662);
nand U690 (N_690,N_611,N_634);
nor U691 (N_691,N_631,N_635);
xnor U692 (N_692,N_656,N_667);
or U693 (N_693,N_648,N_612);
nor U694 (N_694,N_618,N_638);
nand U695 (N_695,N_645,N_672);
nor U696 (N_696,N_650,N_627);
xnor U697 (N_697,N_640,N_655);
and U698 (N_698,N_643,N_630);
or U699 (N_699,N_664,N_666);
nand U700 (N_700,N_661,N_617);
xnor U701 (N_701,N_608,N_653);
or U702 (N_702,N_619,N_660);
or U703 (N_703,N_639,N_665);
nand U704 (N_704,N_607,N_609);
nor U705 (N_705,N_642,N_626);
xnor U706 (N_706,N_621,N_663);
nand U707 (N_707,N_632,N_658);
or U708 (N_708,N_674,N_668);
nand U709 (N_709,N_628,N_659);
xor U710 (N_710,N_613,N_670);
xor U711 (N_711,N_615,N_606);
and U712 (N_712,N_601,N_613);
nor U713 (N_713,N_659,N_620);
nand U714 (N_714,N_603,N_614);
nor U715 (N_715,N_641,N_674);
nor U716 (N_716,N_668,N_605);
or U717 (N_717,N_651,N_604);
and U718 (N_718,N_660,N_636);
xnor U719 (N_719,N_602,N_634);
nand U720 (N_720,N_647,N_661);
nor U721 (N_721,N_628,N_645);
or U722 (N_722,N_638,N_665);
xnor U723 (N_723,N_670,N_641);
and U724 (N_724,N_628,N_614);
nor U725 (N_725,N_627,N_642);
and U726 (N_726,N_617,N_668);
xnor U727 (N_727,N_652,N_643);
nand U728 (N_728,N_635,N_626);
nor U729 (N_729,N_618,N_616);
nand U730 (N_730,N_613,N_654);
or U731 (N_731,N_661,N_637);
xnor U732 (N_732,N_632,N_616);
or U733 (N_733,N_600,N_616);
or U734 (N_734,N_655,N_631);
and U735 (N_735,N_668,N_645);
nor U736 (N_736,N_653,N_612);
nor U737 (N_737,N_602,N_648);
nor U738 (N_738,N_607,N_603);
and U739 (N_739,N_642,N_608);
and U740 (N_740,N_666,N_659);
or U741 (N_741,N_643,N_619);
nor U742 (N_742,N_664,N_663);
or U743 (N_743,N_614,N_640);
or U744 (N_744,N_668,N_649);
xnor U745 (N_745,N_629,N_614);
nand U746 (N_746,N_602,N_640);
xor U747 (N_747,N_660,N_634);
nor U748 (N_748,N_609,N_642);
xor U749 (N_749,N_650,N_662);
or U750 (N_750,N_736,N_722);
xnor U751 (N_751,N_706,N_745);
nand U752 (N_752,N_690,N_686);
nand U753 (N_753,N_708,N_675);
xnor U754 (N_754,N_696,N_732);
xor U755 (N_755,N_682,N_692);
nand U756 (N_756,N_725,N_695);
nand U757 (N_757,N_731,N_707);
nand U758 (N_758,N_704,N_710);
nor U759 (N_759,N_747,N_721);
xor U760 (N_760,N_713,N_699);
nand U761 (N_761,N_698,N_697);
nor U762 (N_762,N_687,N_703);
and U763 (N_763,N_720,N_742);
and U764 (N_764,N_693,N_744);
and U765 (N_765,N_711,N_702);
xnor U766 (N_766,N_718,N_689);
nand U767 (N_767,N_700,N_714);
and U768 (N_768,N_701,N_746);
or U769 (N_769,N_705,N_685);
nor U770 (N_770,N_712,N_743);
nand U771 (N_771,N_679,N_741);
or U772 (N_772,N_688,N_726);
nand U773 (N_773,N_730,N_734);
nand U774 (N_774,N_680,N_738);
nand U775 (N_775,N_729,N_709);
nor U776 (N_776,N_719,N_735);
xnor U777 (N_777,N_733,N_728);
or U778 (N_778,N_715,N_694);
xor U779 (N_779,N_678,N_676);
xnor U780 (N_780,N_681,N_737);
xnor U781 (N_781,N_739,N_727);
and U782 (N_782,N_716,N_748);
nand U783 (N_783,N_684,N_717);
or U784 (N_784,N_749,N_724);
nor U785 (N_785,N_723,N_683);
xor U786 (N_786,N_691,N_677);
or U787 (N_787,N_740,N_698);
or U788 (N_788,N_738,N_699);
and U789 (N_789,N_744,N_703);
or U790 (N_790,N_695,N_726);
nand U791 (N_791,N_697,N_700);
xnor U792 (N_792,N_734,N_714);
or U793 (N_793,N_744,N_724);
or U794 (N_794,N_745,N_699);
or U795 (N_795,N_729,N_690);
nand U796 (N_796,N_749,N_734);
nor U797 (N_797,N_738,N_733);
xnor U798 (N_798,N_748,N_722);
xor U799 (N_799,N_746,N_732);
xor U800 (N_800,N_710,N_706);
nor U801 (N_801,N_701,N_732);
and U802 (N_802,N_733,N_731);
or U803 (N_803,N_684,N_698);
nand U804 (N_804,N_711,N_747);
xor U805 (N_805,N_731,N_697);
xor U806 (N_806,N_686,N_738);
and U807 (N_807,N_685,N_741);
and U808 (N_808,N_716,N_731);
nor U809 (N_809,N_692,N_709);
and U810 (N_810,N_706,N_738);
xor U811 (N_811,N_692,N_710);
and U812 (N_812,N_682,N_694);
and U813 (N_813,N_718,N_712);
nand U814 (N_814,N_697,N_711);
and U815 (N_815,N_684,N_719);
nor U816 (N_816,N_683,N_676);
xnor U817 (N_817,N_713,N_733);
nand U818 (N_818,N_711,N_712);
or U819 (N_819,N_685,N_720);
xor U820 (N_820,N_684,N_743);
nor U821 (N_821,N_679,N_706);
xor U822 (N_822,N_713,N_735);
and U823 (N_823,N_718,N_740);
and U824 (N_824,N_679,N_733);
nor U825 (N_825,N_820,N_811);
nor U826 (N_826,N_779,N_770);
and U827 (N_827,N_803,N_813);
and U828 (N_828,N_757,N_817);
and U829 (N_829,N_800,N_766);
nor U830 (N_830,N_773,N_760);
or U831 (N_831,N_814,N_793);
nor U832 (N_832,N_756,N_778);
nor U833 (N_833,N_790,N_775);
nand U834 (N_834,N_796,N_809);
or U835 (N_835,N_789,N_764);
or U836 (N_836,N_788,N_769);
or U837 (N_837,N_765,N_784);
xor U838 (N_838,N_751,N_761);
nand U839 (N_839,N_812,N_808);
or U840 (N_840,N_776,N_824);
and U841 (N_841,N_777,N_754);
nor U842 (N_842,N_767,N_801);
nor U843 (N_843,N_786,N_758);
and U844 (N_844,N_819,N_780);
xor U845 (N_845,N_804,N_816);
nand U846 (N_846,N_821,N_755);
or U847 (N_847,N_753,N_818);
nor U848 (N_848,N_815,N_822);
nor U849 (N_849,N_762,N_771);
nor U850 (N_850,N_810,N_805);
or U851 (N_851,N_797,N_759);
nand U852 (N_852,N_807,N_781);
or U853 (N_853,N_792,N_806);
and U854 (N_854,N_752,N_783);
xor U855 (N_855,N_785,N_774);
or U856 (N_856,N_787,N_763);
nor U857 (N_857,N_795,N_798);
and U858 (N_858,N_799,N_768);
and U859 (N_859,N_782,N_750);
xnor U860 (N_860,N_794,N_791);
nand U861 (N_861,N_823,N_802);
and U862 (N_862,N_772,N_796);
nor U863 (N_863,N_765,N_754);
nand U864 (N_864,N_818,N_757);
and U865 (N_865,N_752,N_792);
or U866 (N_866,N_763,N_808);
nor U867 (N_867,N_801,N_777);
nand U868 (N_868,N_752,N_814);
xnor U869 (N_869,N_804,N_795);
or U870 (N_870,N_771,N_780);
xor U871 (N_871,N_774,N_813);
and U872 (N_872,N_770,N_791);
nor U873 (N_873,N_781,N_759);
and U874 (N_874,N_777,N_803);
and U875 (N_875,N_800,N_784);
and U876 (N_876,N_750,N_775);
or U877 (N_877,N_762,N_775);
and U878 (N_878,N_778,N_801);
nor U879 (N_879,N_755,N_757);
xor U880 (N_880,N_813,N_754);
or U881 (N_881,N_758,N_820);
nand U882 (N_882,N_785,N_761);
nor U883 (N_883,N_795,N_787);
and U884 (N_884,N_818,N_755);
nor U885 (N_885,N_814,N_768);
nor U886 (N_886,N_760,N_821);
nand U887 (N_887,N_751,N_775);
xnor U888 (N_888,N_780,N_808);
xor U889 (N_889,N_780,N_751);
nor U890 (N_890,N_784,N_751);
and U891 (N_891,N_812,N_750);
xor U892 (N_892,N_808,N_806);
nor U893 (N_893,N_817,N_814);
or U894 (N_894,N_820,N_756);
xnor U895 (N_895,N_762,N_774);
and U896 (N_896,N_812,N_817);
nor U897 (N_897,N_780,N_810);
or U898 (N_898,N_821,N_800);
xor U899 (N_899,N_770,N_754);
or U900 (N_900,N_876,N_879);
nor U901 (N_901,N_863,N_861);
or U902 (N_902,N_887,N_841);
xnor U903 (N_903,N_898,N_834);
and U904 (N_904,N_880,N_864);
or U905 (N_905,N_825,N_852);
nor U906 (N_906,N_889,N_886);
or U907 (N_907,N_853,N_831);
or U908 (N_908,N_827,N_833);
nor U909 (N_909,N_891,N_892);
or U910 (N_910,N_851,N_842);
or U911 (N_911,N_896,N_888);
and U912 (N_912,N_848,N_854);
and U913 (N_913,N_862,N_835);
nor U914 (N_914,N_873,N_868);
xnor U915 (N_915,N_883,N_839);
nor U916 (N_916,N_870,N_882);
and U917 (N_917,N_881,N_872);
and U918 (N_918,N_899,N_885);
or U919 (N_919,N_830,N_840);
or U920 (N_920,N_832,N_847);
or U921 (N_921,N_894,N_866);
or U922 (N_922,N_836,N_828);
or U923 (N_923,N_897,N_867);
and U924 (N_924,N_871,N_850);
nor U925 (N_925,N_895,N_859);
nand U926 (N_926,N_890,N_844);
xnor U927 (N_927,N_874,N_858);
nand U928 (N_928,N_845,N_826);
nor U929 (N_929,N_865,N_860);
xnor U930 (N_930,N_884,N_878);
nand U931 (N_931,N_857,N_838);
or U932 (N_932,N_843,N_877);
and U933 (N_933,N_837,N_855);
nor U934 (N_934,N_829,N_869);
and U935 (N_935,N_849,N_875);
xnor U936 (N_936,N_893,N_846);
nand U937 (N_937,N_856,N_886);
xnor U938 (N_938,N_853,N_855);
and U939 (N_939,N_865,N_882);
xor U940 (N_940,N_874,N_859);
or U941 (N_941,N_872,N_873);
xor U942 (N_942,N_830,N_837);
xor U943 (N_943,N_843,N_846);
xor U944 (N_944,N_838,N_825);
nand U945 (N_945,N_842,N_881);
nand U946 (N_946,N_884,N_833);
nor U947 (N_947,N_878,N_831);
and U948 (N_948,N_862,N_851);
xor U949 (N_949,N_850,N_826);
nand U950 (N_950,N_868,N_858);
nor U951 (N_951,N_890,N_854);
nor U952 (N_952,N_826,N_842);
nor U953 (N_953,N_840,N_890);
nand U954 (N_954,N_866,N_847);
nand U955 (N_955,N_854,N_883);
nand U956 (N_956,N_829,N_844);
xnor U957 (N_957,N_827,N_862);
nor U958 (N_958,N_893,N_843);
or U959 (N_959,N_888,N_844);
nand U960 (N_960,N_833,N_863);
and U961 (N_961,N_860,N_862);
or U962 (N_962,N_835,N_841);
nand U963 (N_963,N_848,N_831);
or U964 (N_964,N_831,N_826);
nor U965 (N_965,N_855,N_830);
nand U966 (N_966,N_849,N_844);
and U967 (N_967,N_861,N_855);
nor U968 (N_968,N_838,N_892);
and U969 (N_969,N_872,N_889);
and U970 (N_970,N_833,N_831);
xor U971 (N_971,N_873,N_837);
and U972 (N_972,N_887,N_828);
or U973 (N_973,N_886,N_876);
xor U974 (N_974,N_879,N_895);
nor U975 (N_975,N_900,N_956);
nand U976 (N_976,N_954,N_903);
nand U977 (N_977,N_939,N_902);
nor U978 (N_978,N_912,N_957);
nand U979 (N_979,N_928,N_953);
xor U980 (N_980,N_906,N_955);
or U981 (N_981,N_942,N_950);
and U982 (N_982,N_908,N_919);
nand U983 (N_983,N_945,N_930);
nor U984 (N_984,N_926,N_921);
xor U985 (N_985,N_901,N_960);
or U986 (N_986,N_914,N_916);
xnor U987 (N_987,N_965,N_925);
nor U988 (N_988,N_944,N_959);
nand U989 (N_989,N_936,N_958);
nand U990 (N_990,N_910,N_968);
nand U991 (N_991,N_937,N_973);
nand U992 (N_992,N_907,N_924);
and U993 (N_993,N_929,N_971);
nand U994 (N_994,N_949,N_918);
and U995 (N_995,N_963,N_969);
and U996 (N_996,N_972,N_917);
nand U997 (N_997,N_951,N_966);
xor U998 (N_998,N_940,N_935);
and U999 (N_999,N_948,N_927);
and U1000 (N_1000,N_941,N_946);
and U1001 (N_1001,N_933,N_904);
nand U1002 (N_1002,N_962,N_961);
nand U1003 (N_1003,N_915,N_947);
xnor U1004 (N_1004,N_964,N_934);
nand U1005 (N_1005,N_931,N_967);
nand U1006 (N_1006,N_913,N_938);
nand U1007 (N_1007,N_943,N_974);
nor U1008 (N_1008,N_970,N_922);
xor U1009 (N_1009,N_923,N_905);
nand U1010 (N_1010,N_952,N_911);
xor U1011 (N_1011,N_909,N_920);
nand U1012 (N_1012,N_932,N_944);
nor U1013 (N_1013,N_900,N_929);
nand U1014 (N_1014,N_954,N_944);
xor U1015 (N_1015,N_926,N_915);
nand U1016 (N_1016,N_938,N_969);
xor U1017 (N_1017,N_927,N_937);
or U1018 (N_1018,N_932,N_904);
nand U1019 (N_1019,N_962,N_926);
nand U1020 (N_1020,N_955,N_948);
xnor U1021 (N_1021,N_911,N_966);
and U1022 (N_1022,N_947,N_906);
nand U1023 (N_1023,N_950,N_969);
and U1024 (N_1024,N_936,N_901);
or U1025 (N_1025,N_972,N_971);
and U1026 (N_1026,N_964,N_926);
nor U1027 (N_1027,N_963,N_972);
or U1028 (N_1028,N_970,N_938);
and U1029 (N_1029,N_919,N_943);
and U1030 (N_1030,N_936,N_938);
nor U1031 (N_1031,N_907,N_947);
or U1032 (N_1032,N_932,N_956);
nor U1033 (N_1033,N_915,N_904);
nand U1034 (N_1034,N_948,N_972);
nor U1035 (N_1035,N_947,N_943);
and U1036 (N_1036,N_940,N_944);
and U1037 (N_1037,N_960,N_925);
nand U1038 (N_1038,N_970,N_940);
and U1039 (N_1039,N_910,N_967);
nor U1040 (N_1040,N_900,N_949);
nand U1041 (N_1041,N_959,N_956);
or U1042 (N_1042,N_971,N_969);
xor U1043 (N_1043,N_969,N_946);
xnor U1044 (N_1044,N_960,N_973);
nor U1045 (N_1045,N_944,N_952);
nand U1046 (N_1046,N_950,N_930);
xor U1047 (N_1047,N_952,N_904);
xor U1048 (N_1048,N_926,N_953);
and U1049 (N_1049,N_950,N_961);
and U1050 (N_1050,N_979,N_1048);
or U1051 (N_1051,N_1020,N_978);
xor U1052 (N_1052,N_1007,N_982);
and U1053 (N_1053,N_1040,N_984);
and U1054 (N_1054,N_1016,N_1038);
xor U1055 (N_1055,N_985,N_1034);
xnor U1056 (N_1056,N_1013,N_1035);
nand U1057 (N_1057,N_991,N_1025);
or U1058 (N_1058,N_1024,N_987);
xnor U1059 (N_1059,N_988,N_1043);
nor U1060 (N_1060,N_1046,N_1042);
and U1061 (N_1061,N_983,N_1030);
xnor U1062 (N_1062,N_1044,N_1023);
xnor U1063 (N_1063,N_997,N_1049);
and U1064 (N_1064,N_1018,N_1022);
nor U1065 (N_1065,N_1017,N_1019);
xnor U1066 (N_1066,N_999,N_986);
and U1067 (N_1067,N_998,N_1015);
nand U1068 (N_1068,N_1039,N_992);
or U1069 (N_1069,N_980,N_996);
or U1070 (N_1070,N_1002,N_993);
and U1071 (N_1071,N_1032,N_975);
xnor U1072 (N_1072,N_1011,N_1009);
xnor U1073 (N_1073,N_1031,N_977);
nor U1074 (N_1074,N_989,N_1026);
nor U1075 (N_1075,N_1000,N_1014);
and U1076 (N_1076,N_1008,N_1029);
nand U1077 (N_1077,N_1037,N_1021);
nor U1078 (N_1078,N_1027,N_994);
nor U1079 (N_1079,N_1010,N_1045);
nand U1080 (N_1080,N_981,N_1006);
or U1081 (N_1081,N_1004,N_995);
and U1082 (N_1082,N_1003,N_1033);
or U1083 (N_1083,N_990,N_1047);
nand U1084 (N_1084,N_1005,N_1036);
and U1085 (N_1085,N_1012,N_976);
xnor U1086 (N_1086,N_1041,N_1028);
xnor U1087 (N_1087,N_1001,N_996);
or U1088 (N_1088,N_976,N_1000);
nand U1089 (N_1089,N_1044,N_1049);
nand U1090 (N_1090,N_993,N_1049);
nand U1091 (N_1091,N_984,N_1013);
nand U1092 (N_1092,N_1033,N_1010);
nand U1093 (N_1093,N_1000,N_990);
xnor U1094 (N_1094,N_993,N_979);
and U1095 (N_1095,N_988,N_1027);
and U1096 (N_1096,N_998,N_1002);
xnor U1097 (N_1097,N_995,N_1046);
nand U1098 (N_1098,N_1034,N_1008);
xor U1099 (N_1099,N_1035,N_983);
or U1100 (N_1100,N_982,N_995);
or U1101 (N_1101,N_1006,N_1040);
and U1102 (N_1102,N_984,N_1004);
or U1103 (N_1103,N_991,N_981);
and U1104 (N_1104,N_993,N_1013);
xor U1105 (N_1105,N_1014,N_1002);
and U1106 (N_1106,N_1015,N_990);
xor U1107 (N_1107,N_984,N_1019);
nor U1108 (N_1108,N_983,N_1036);
xnor U1109 (N_1109,N_976,N_1020);
and U1110 (N_1110,N_995,N_979);
or U1111 (N_1111,N_1023,N_1009);
nor U1112 (N_1112,N_1045,N_1012);
or U1113 (N_1113,N_980,N_994);
and U1114 (N_1114,N_1041,N_1048);
or U1115 (N_1115,N_986,N_1037);
and U1116 (N_1116,N_1034,N_1023);
or U1117 (N_1117,N_985,N_1001);
or U1118 (N_1118,N_1016,N_1011);
nor U1119 (N_1119,N_993,N_999);
and U1120 (N_1120,N_996,N_1037);
and U1121 (N_1121,N_1013,N_1009);
nand U1122 (N_1122,N_1030,N_982);
nand U1123 (N_1123,N_1038,N_1024);
nand U1124 (N_1124,N_1008,N_1031);
and U1125 (N_1125,N_1062,N_1109);
and U1126 (N_1126,N_1083,N_1110);
or U1127 (N_1127,N_1096,N_1090);
nand U1128 (N_1128,N_1067,N_1075);
nand U1129 (N_1129,N_1060,N_1057);
or U1130 (N_1130,N_1116,N_1073);
and U1131 (N_1131,N_1072,N_1066);
or U1132 (N_1132,N_1102,N_1054);
nand U1133 (N_1133,N_1061,N_1082);
nand U1134 (N_1134,N_1092,N_1089);
nand U1135 (N_1135,N_1068,N_1053);
or U1136 (N_1136,N_1076,N_1094);
and U1137 (N_1137,N_1106,N_1051);
nor U1138 (N_1138,N_1084,N_1063);
and U1139 (N_1139,N_1052,N_1065);
or U1140 (N_1140,N_1122,N_1100);
nor U1141 (N_1141,N_1107,N_1050);
or U1142 (N_1142,N_1056,N_1079);
nor U1143 (N_1143,N_1087,N_1111);
or U1144 (N_1144,N_1112,N_1059);
xnor U1145 (N_1145,N_1064,N_1123);
xnor U1146 (N_1146,N_1093,N_1118);
and U1147 (N_1147,N_1058,N_1099);
xor U1148 (N_1148,N_1070,N_1108);
nor U1149 (N_1149,N_1117,N_1124);
and U1150 (N_1150,N_1071,N_1080);
xor U1151 (N_1151,N_1055,N_1077);
nor U1152 (N_1152,N_1097,N_1069);
or U1153 (N_1153,N_1098,N_1119);
nor U1154 (N_1154,N_1103,N_1091);
or U1155 (N_1155,N_1121,N_1086);
or U1156 (N_1156,N_1095,N_1085);
nand U1157 (N_1157,N_1074,N_1114);
and U1158 (N_1158,N_1088,N_1078);
nand U1159 (N_1159,N_1115,N_1113);
or U1160 (N_1160,N_1120,N_1081);
or U1161 (N_1161,N_1101,N_1104);
nor U1162 (N_1162,N_1105,N_1066);
nand U1163 (N_1163,N_1114,N_1050);
nand U1164 (N_1164,N_1061,N_1104);
or U1165 (N_1165,N_1090,N_1087);
and U1166 (N_1166,N_1062,N_1104);
nor U1167 (N_1167,N_1082,N_1068);
or U1168 (N_1168,N_1084,N_1103);
or U1169 (N_1169,N_1066,N_1064);
xnor U1170 (N_1170,N_1118,N_1085);
and U1171 (N_1171,N_1085,N_1106);
nand U1172 (N_1172,N_1050,N_1086);
or U1173 (N_1173,N_1077,N_1099);
and U1174 (N_1174,N_1057,N_1117);
or U1175 (N_1175,N_1057,N_1096);
xnor U1176 (N_1176,N_1097,N_1110);
or U1177 (N_1177,N_1071,N_1061);
nor U1178 (N_1178,N_1119,N_1076);
nor U1179 (N_1179,N_1113,N_1075);
or U1180 (N_1180,N_1108,N_1100);
or U1181 (N_1181,N_1095,N_1078);
nor U1182 (N_1182,N_1118,N_1083);
nor U1183 (N_1183,N_1056,N_1053);
nor U1184 (N_1184,N_1054,N_1123);
or U1185 (N_1185,N_1122,N_1124);
xnor U1186 (N_1186,N_1110,N_1121);
or U1187 (N_1187,N_1089,N_1071);
or U1188 (N_1188,N_1114,N_1106);
or U1189 (N_1189,N_1095,N_1100);
or U1190 (N_1190,N_1114,N_1076);
xnor U1191 (N_1191,N_1117,N_1096);
nand U1192 (N_1192,N_1065,N_1079);
and U1193 (N_1193,N_1123,N_1111);
xnor U1194 (N_1194,N_1094,N_1120);
and U1195 (N_1195,N_1052,N_1109);
xor U1196 (N_1196,N_1064,N_1085);
nor U1197 (N_1197,N_1108,N_1122);
and U1198 (N_1198,N_1100,N_1082);
nor U1199 (N_1199,N_1066,N_1096);
xnor U1200 (N_1200,N_1145,N_1191);
nand U1201 (N_1201,N_1154,N_1175);
or U1202 (N_1202,N_1146,N_1162);
nor U1203 (N_1203,N_1169,N_1142);
xor U1204 (N_1204,N_1172,N_1149);
nor U1205 (N_1205,N_1197,N_1196);
and U1206 (N_1206,N_1153,N_1130);
or U1207 (N_1207,N_1139,N_1167);
xnor U1208 (N_1208,N_1168,N_1188);
nor U1209 (N_1209,N_1144,N_1177);
or U1210 (N_1210,N_1127,N_1173);
nor U1211 (N_1211,N_1161,N_1199);
nor U1212 (N_1212,N_1148,N_1141);
or U1213 (N_1213,N_1135,N_1189);
nand U1214 (N_1214,N_1159,N_1158);
nand U1215 (N_1215,N_1176,N_1181);
xor U1216 (N_1216,N_1171,N_1131);
nor U1217 (N_1217,N_1165,N_1155);
nand U1218 (N_1218,N_1195,N_1179);
xnor U1219 (N_1219,N_1170,N_1178);
nand U1220 (N_1220,N_1137,N_1183);
xnor U1221 (N_1221,N_1128,N_1190);
and U1222 (N_1222,N_1132,N_1138);
nand U1223 (N_1223,N_1133,N_1147);
or U1224 (N_1224,N_1134,N_1198);
or U1225 (N_1225,N_1157,N_1187);
xnor U1226 (N_1226,N_1192,N_1140);
nand U1227 (N_1227,N_1174,N_1126);
and U1228 (N_1228,N_1160,N_1180);
xor U1229 (N_1229,N_1193,N_1182);
nor U1230 (N_1230,N_1163,N_1150);
or U1231 (N_1231,N_1129,N_1166);
or U1232 (N_1232,N_1143,N_1186);
nor U1233 (N_1233,N_1194,N_1185);
xor U1234 (N_1234,N_1164,N_1156);
nor U1235 (N_1235,N_1151,N_1136);
or U1236 (N_1236,N_1125,N_1184);
and U1237 (N_1237,N_1152,N_1199);
xor U1238 (N_1238,N_1186,N_1161);
or U1239 (N_1239,N_1148,N_1150);
or U1240 (N_1240,N_1137,N_1165);
nor U1241 (N_1241,N_1127,N_1190);
and U1242 (N_1242,N_1127,N_1156);
nand U1243 (N_1243,N_1178,N_1176);
or U1244 (N_1244,N_1181,N_1199);
nand U1245 (N_1245,N_1175,N_1130);
nand U1246 (N_1246,N_1143,N_1140);
and U1247 (N_1247,N_1139,N_1164);
xnor U1248 (N_1248,N_1127,N_1148);
or U1249 (N_1249,N_1175,N_1185);
or U1250 (N_1250,N_1169,N_1185);
and U1251 (N_1251,N_1156,N_1184);
or U1252 (N_1252,N_1171,N_1138);
nand U1253 (N_1253,N_1135,N_1148);
or U1254 (N_1254,N_1132,N_1157);
and U1255 (N_1255,N_1137,N_1130);
xnor U1256 (N_1256,N_1197,N_1186);
and U1257 (N_1257,N_1158,N_1198);
xor U1258 (N_1258,N_1156,N_1165);
nor U1259 (N_1259,N_1165,N_1169);
nor U1260 (N_1260,N_1190,N_1130);
and U1261 (N_1261,N_1193,N_1142);
nand U1262 (N_1262,N_1149,N_1168);
nor U1263 (N_1263,N_1169,N_1139);
or U1264 (N_1264,N_1138,N_1153);
xor U1265 (N_1265,N_1135,N_1131);
nand U1266 (N_1266,N_1131,N_1153);
xnor U1267 (N_1267,N_1172,N_1146);
and U1268 (N_1268,N_1155,N_1162);
and U1269 (N_1269,N_1130,N_1139);
and U1270 (N_1270,N_1163,N_1131);
nor U1271 (N_1271,N_1131,N_1194);
nand U1272 (N_1272,N_1182,N_1188);
nor U1273 (N_1273,N_1164,N_1168);
and U1274 (N_1274,N_1193,N_1194);
nor U1275 (N_1275,N_1221,N_1257);
nor U1276 (N_1276,N_1253,N_1224);
or U1277 (N_1277,N_1201,N_1200);
nor U1278 (N_1278,N_1240,N_1256);
xor U1279 (N_1279,N_1232,N_1216);
and U1280 (N_1280,N_1208,N_1203);
xnor U1281 (N_1281,N_1218,N_1243);
or U1282 (N_1282,N_1263,N_1217);
nand U1283 (N_1283,N_1246,N_1266);
xnor U1284 (N_1284,N_1250,N_1213);
xnor U1285 (N_1285,N_1264,N_1244);
and U1286 (N_1286,N_1258,N_1241);
nand U1287 (N_1287,N_1247,N_1274);
and U1288 (N_1288,N_1252,N_1211);
nor U1289 (N_1289,N_1235,N_1238);
xnor U1290 (N_1290,N_1242,N_1271);
xor U1291 (N_1291,N_1227,N_1207);
xnor U1292 (N_1292,N_1223,N_1259);
and U1293 (N_1293,N_1239,N_1214);
and U1294 (N_1294,N_1269,N_1225);
xor U1295 (N_1295,N_1205,N_1245);
nand U1296 (N_1296,N_1233,N_1272);
nor U1297 (N_1297,N_1268,N_1249);
xor U1298 (N_1298,N_1237,N_1230);
xor U1299 (N_1299,N_1248,N_1220);
nor U1300 (N_1300,N_1228,N_1255);
nand U1301 (N_1301,N_1206,N_1231);
xor U1302 (N_1302,N_1267,N_1202);
nand U1303 (N_1303,N_1254,N_1261);
nand U1304 (N_1304,N_1251,N_1226);
and U1305 (N_1305,N_1229,N_1270);
xor U1306 (N_1306,N_1260,N_1210);
nand U1307 (N_1307,N_1212,N_1222);
xnor U1308 (N_1308,N_1204,N_1262);
xnor U1309 (N_1309,N_1265,N_1209);
or U1310 (N_1310,N_1215,N_1219);
xor U1311 (N_1311,N_1234,N_1236);
xor U1312 (N_1312,N_1273,N_1224);
nor U1313 (N_1313,N_1216,N_1228);
nand U1314 (N_1314,N_1207,N_1252);
xnor U1315 (N_1315,N_1270,N_1258);
and U1316 (N_1316,N_1251,N_1210);
nand U1317 (N_1317,N_1232,N_1218);
nand U1318 (N_1318,N_1209,N_1255);
nand U1319 (N_1319,N_1270,N_1202);
nand U1320 (N_1320,N_1214,N_1255);
and U1321 (N_1321,N_1200,N_1240);
or U1322 (N_1322,N_1243,N_1226);
nor U1323 (N_1323,N_1254,N_1260);
nand U1324 (N_1324,N_1238,N_1226);
or U1325 (N_1325,N_1225,N_1272);
nor U1326 (N_1326,N_1238,N_1205);
and U1327 (N_1327,N_1211,N_1225);
and U1328 (N_1328,N_1233,N_1244);
xor U1329 (N_1329,N_1248,N_1227);
or U1330 (N_1330,N_1236,N_1211);
or U1331 (N_1331,N_1219,N_1210);
xor U1332 (N_1332,N_1214,N_1243);
nor U1333 (N_1333,N_1208,N_1270);
nor U1334 (N_1334,N_1248,N_1200);
and U1335 (N_1335,N_1202,N_1260);
nand U1336 (N_1336,N_1220,N_1243);
and U1337 (N_1337,N_1261,N_1248);
xor U1338 (N_1338,N_1209,N_1251);
nor U1339 (N_1339,N_1250,N_1265);
nor U1340 (N_1340,N_1259,N_1212);
or U1341 (N_1341,N_1245,N_1265);
nand U1342 (N_1342,N_1250,N_1219);
and U1343 (N_1343,N_1256,N_1214);
nand U1344 (N_1344,N_1258,N_1255);
and U1345 (N_1345,N_1236,N_1221);
xnor U1346 (N_1346,N_1253,N_1207);
or U1347 (N_1347,N_1205,N_1254);
xnor U1348 (N_1348,N_1241,N_1264);
or U1349 (N_1349,N_1234,N_1202);
xnor U1350 (N_1350,N_1275,N_1346);
or U1351 (N_1351,N_1296,N_1302);
nor U1352 (N_1352,N_1340,N_1291);
and U1353 (N_1353,N_1335,N_1323);
nor U1354 (N_1354,N_1289,N_1347);
or U1355 (N_1355,N_1337,N_1277);
and U1356 (N_1356,N_1278,N_1281);
xor U1357 (N_1357,N_1287,N_1334);
nand U1358 (N_1358,N_1325,N_1343);
nand U1359 (N_1359,N_1326,N_1341);
and U1360 (N_1360,N_1345,N_1286);
or U1361 (N_1361,N_1310,N_1333);
xor U1362 (N_1362,N_1290,N_1309);
or U1363 (N_1363,N_1297,N_1307);
and U1364 (N_1364,N_1331,N_1324);
and U1365 (N_1365,N_1305,N_1320);
nor U1366 (N_1366,N_1298,N_1292);
nor U1367 (N_1367,N_1317,N_1339);
nand U1368 (N_1368,N_1300,N_1327);
nor U1369 (N_1369,N_1279,N_1313);
nand U1370 (N_1370,N_1348,N_1306);
nand U1371 (N_1371,N_1304,N_1342);
nand U1372 (N_1372,N_1321,N_1284);
xor U1373 (N_1373,N_1314,N_1336);
nand U1374 (N_1374,N_1311,N_1312);
nor U1375 (N_1375,N_1276,N_1330);
nand U1376 (N_1376,N_1316,N_1328);
nand U1377 (N_1377,N_1282,N_1303);
nand U1378 (N_1378,N_1294,N_1322);
nand U1379 (N_1379,N_1295,N_1344);
nand U1380 (N_1380,N_1299,N_1293);
nor U1381 (N_1381,N_1285,N_1280);
nor U1382 (N_1382,N_1318,N_1308);
and U1383 (N_1383,N_1288,N_1338);
xor U1384 (N_1384,N_1283,N_1329);
and U1385 (N_1385,N_1349,N_1301);
xnor U1386 (N_1386,N_1319,N_1332);
nor U1387 (N_1387,N_1315,N_1284);
xnor U1388 (N_1388,N_1306,N_1283);
or U1389 (N_1389,N_1343,N_1308);
or U1390 (N_1390,N_1296,N_1276);
xnor U1391 (N_1391,N_1278,N_1327);
or U1392 (N_1392,N_1286,N_1292);
or U1393 (N_1393,N_1290,N_1332);
or U1394 (N_1394,N_1301,N_1296);
and U1395 (N_1395,N_1304,N_1285);
nand U1396 (N_1396,N_1311,N_1329);
xor U1397 (N_1397,N_1277,N_1296);
or U1398 (N_1398,N_1280,N_1330);
nor U1399 (N_1399,N_1330,N_1335);
xor U1400 (N_1400,N_1299,N_1300);
nand U1401 (N_1401,N_1305,N_1325);
xor U1402 (N_1402,N_1348,N_1292);
and U1403 (N_1403,N_1340,N_1293);
or U1404 (N_1404,N_1342,N_1298);
or U1405 (N_1405,N_1313,N_1343);
nor U1406 (N_1406,N_1344,N_1320);
or U1407 (N_1407,N_1325,N_1316);
or U1408 (N_1408,N_1301,N_1284);
and U1409 (N_1409,N_1338,N_1320);
xnor U1410 (N_1410,N_1297,N_1338);
and U1411 (N_1411,N_1315,N_1336);
xnor U1412 (N_1412,N_1324,N_1306);
and U1413 (N_1413,N_1308,N_1347);
or U1414 (N_1414,N_1298,N_1284);
nor U1415 (N_1415,N_1349,N_1332);
and U1416 (N_1416,N_1309,N_1322);
and U1417 (N_1417,N_1280,N_1295);
nand U1418 (N_1418,N_1297,N_1281);
xor U1419 (N_1419,N_1300,N_1331);
and U1420 (N_1420,N_1300,N_1318);
or U1421 (N_1421,N_1298,N_1318);
and U1422 (N_1422,N_1312,N_1305);
xnor U1423 (N_1423,N_1304,N_1311);
nor U1424 (N_1424,N_1330,N_1293);
and U1425 (N_1425,N_1407,N_1405);
nand U1426 (N_1426,N_1398,N_1420);
and U1427 (N_1427,N_1415,N_1410);
or U1428 (N_1428,N_1390,N_1373);
nor U1429 (N_1429,N_1383,N_1374);
and U1430 (N_1430,N_1409,N_1423);
nor U1431 (N_1431,N_1376,N_1419);
xor U1432 (N_1432,N_1350,N_1366);
xnor U1433 (N_1433,N_1372,N_1396);
nand U1434 (N_1434,N_1354,N_1365);
nor U1435 (N_1435,N_1411,N_1386);
and U1436 (N_1436,N_1401,N_1353);
nand U1437 (N_1437,N_1378,N_1388);
nor U1438 (N_1438,N_1387,N_1408);
or U1439 (N_1439,N_1367,N_1377);
and U1440 (N_1440,N_1380,N_1382);
nor U1441 (N_1441,N_1359,N_1369);
and U1442 (N_1442,N_1357,N_1418);
nand U1443 (N_1443,N_1352,N_1356);
xnor U1444 (N_1444,N_1360,N_1393);
or U1445 (N_1445,N_1375,N_1381);
nand U1446 (N_1446,N_1379,N_1402);
or U1447 (N_1447,N_1385,N_1421);
nand U1448 (N_1448,N_1406,N_1412);
xnor U1449 (N_1449,N_1417,N_1392);
and U1450 (N_1450,N_1364,N_1403);
xnor U1451 (N_1451,N_1397,N_1355);
nor U1452 (N_1452,N_1391,N_1371);
or U1453 (N_1453,N_1351,N_1394);
or U1454 (N_1454,N_1370,N_1358);
and U1455 (N_1455,N_1416,N_1395);
xor U1456 (N_1456,N_1404,N_1399);
or U1457 (N_1457,N_1424,N_1361);
and U1458 (N_1458,N_1389,N_1422);
xnor U1459 (N_1459,N_1414,N_1384);
nand U1460 (N_1460,N_1368,N_1413);
or U1461 (N_1461,N_1362,N_1363);
nor U1462 (N_1462,N_1400,N_1375);
or U1463 (N_1463,N_1362,N_1364);
nand U1464 (N_1464,N_1416,N_1390);
xor U1465 (N_1465,N_1350,N_1386);
or U1466 (N_1466,N_1405,N_1365);
and U1467 (N_1467,N_1355,N_1354);
and U1468 (N_1468,N_1370,N_1355);
nand U1469 (N_1469,N_1395,N_1386);
nand U1470 (N_1470,N_1380,N_1378);
nand U1471 (N_1471,N_1404,N_1390);
and U1472 (N_1472,N_1403,N_1363);
nor U1473 (N_1473,N_1399,N_1382);
nand U1474 (N_1474,N_1415,N_1375);
or U1475 (N_1475,N_1357,N_1358);
nor U1476 (N_1476,N_1398,N_1382);
and U1477 (N_1477,N_1418,N_1414);
nor U1478 (N_1478,N_1383,N_1354);
xnor U1479 (N_1479,N_1407,N_1381);
and U1480 (N_1480,N_1372,N_1398);
nor U1481 (N_1481,N_1381,N_1416);
or U1482 (N_1482,N_1401,N_1404);
xor U1483 (N_1483,N_1395,N_1411);
nand U1484 (N_1484,N_1418,N_1355);
nor U1485 (N_1485,N_1414,N_1407);
xnor U1486 (N_1486,N_1381,N_1358);
nand U1487 (N_1487,N_1368,N_1380);
nand U1488 (N_1488,N_1368,N_1407);
xor U1489 (N_1489,N_1405,N_1419);
nor U1490 (N_1490,N_1407,N_1379);
and U1491 (N_1491,N_1373,N_1409);
xor U1492 (N_1492,N_1362,N_1390);
and U1493 (N_1493,N_1423,N_1393);
nand U1494 (N_1494,N_1409,N_1353);
nand U1495 (N_1495,N_1423,N_1400);
nand U1496 (N_1496,N_1393,N_1394);
and U1497 (N_1497,N_1379,N_1360);
or U1498 (N_1498,N_1360,N_1362);
and U1499 (N_1499,N_1400,N_1409);
or U1500 (N_1500,N_1457,N_1432);
nor U1501 (N_1501,N_1495,N_1442);
xnor U1502 (N_1502,N_1464,N_1440);
xor U1503 (N_1503,N_1447,N_1469);
nand U1504 (N_1504,N_1437,N_1467);
and U1505 (N_1505,N_1480,N_1446);
nand U1506 (N_1506,N_1492,N_1450);
or U1507 (N_1507,N_1448,N_1452);
and U1508 (N_1508,N_1462,N_1438);
or U1509 (N_1509,N_1470,N_1455);
nand U1510 (N_1510,N_1451,N_1456);
nand U1511 (N_1511,N_1461,N_1441);
nand U1512 (N_1512,N_1490,N_1476);
xnor U1513 (N_1513,N_1485,N_1443);
nor U1514 (N_1514,N_1493,N_1425);
xor U1515 (N_1515,N_1444,N_1463);
nand U1516 (N_1516,N_1459,N_1478);
and U1517 (N_1517,N_1486,N_1445);
nand U1518 (N_1518,N_1481,N_1454);
nor U1519 (N_1519,N_1436,N_1497);
nand U1520 (N_1520,N_1471,N_1453);
xor U1521 (N_1521,N_1489,N_1477);
and U1522 (N_1522,N_1479,N_1458);
xnor U1523 (N_1523,N_1491,N_1496);
nor U1524 (N_1524,N_1474,N_1433);
nor U1525 (N_1525,N_1472,N_1426);
and U1526 (N_1526,N_1475,N_1431);
and U1527 (N_1527,N_1482,N_1499);
xnor U1528 (N_1528,N_1483,N_1488);
nand U1529 (N_1529,N_1487,N_1484);
xor U1530 (N_1530,N_1460,N_1473);
nand U1531 (N_1531,N_1429,N_1435);
and U1532 (N_1532,N_1439,N_1465);
nand U1533 (N_1533,N_1449,N_1430);
nand U1534 (N_1534,N_1494,N_1428);
xor U1535 (N_1535,N_1434,N_1427);
nand U1536 (N_1536,N_1498,N_1466);
and U1537 (N_1537,N_1468,N_1481);
xor U1538 (N_1538,N_1467,N_1474);
nand U1539 (N_1539,N_1437,N_1431);
and U1540 (N_1540,N_1454,N_1463);
nor U1541 (N_1541,N_1487,N_1492);
and U1542 (N_1542,N_1491,N_1485);
and U1543 (N_1543,N_1442,N_1445);
nand U1544 (N_1544,N_1497,N_1458);
or U1545 (N_1545,N_1452,N_1491);
nor U1546 (N_1546,N_1457,N_1494);
xor U1547 (N_1547,N_1496,N_1440);
or U1548 (N_1548,N_1445,N_1454);
and U1549 (N_1549,N_1472,N_1482);
nor U1550 (N_1550,N_1490,N_1444);
or U1551 (N_1551,N_1472,N_1425);
or U1552 (N_1552,N_1444,N_1456);
or U1553 (N_1553,N_1476,N_1474);
and U1554 (N_1554,N_1468,N_1432);
or U1555 (N_1555,N_1474,N_1489);
and U1556 (N_1556,N_1494,N_1450);
nand U1557 (N_1557,N_1455,N_1462);
nand U1558 (N_1558,N_1482,N_1436);
and U1559 (N_1559,N_1429,N_1430);
and U1560 (N_1560,N_1455,N_1474);
and U1561 (N_1561,N_1475,N_1425);
xnor U1562 (N_1562,N_1467,N_1472);
or U1563 (N_1563,N_1448,N_1447);
and U1564 (N_1564,N_1473,N_1440);
nor U1565 (N_1565,N_1467,N_1451);
nor U1566 (N_1566,N_1428,N_1479);
and U1567 (N_1567,N_1460,N_1467);
and U1568 (N_1568,N_1499,N_1498);
or U1569 (N_1569,N_1480,N_1461);
or U1570 (N_1570,N_1463,N_1478);
and U1571 (N_1571,N_1466,N_1436);
nand U1572 (N_1572,N_1428,N_1439);
and U1573 (N_1573,N_1441,N_1430);
nand U1574 (N_1574,N_1468,N_1459);
nor U1575 (N_1575,N_1546,N_1564);
or U1576 (N_1576,N_1558,N_1551);
and U1577 (N_1577,N_1528,N_1550);
nand U1578 (N_1578,N_1547,N_1568);
and U1579 (N_1579,N_1553,N_1534);
and U1580 (N_1580,N_1503,N_1570);
or U1581 (N_1581,N_1560,N_1507);
or U1582 (N_1582,N_1542,N_1514);
or U1583 (N_1583,N_1543,N_1527);
nand U1584 (N_1584,N_1502,N_1519);
or U1585 (N_1585,N_1525,N_1538);
xnor U1586 (N_1586,N_1504,N_1548);
nor U1587 (N_1587,N_1513,N_1539);
or U1588 (N_1588,N_1501,N_1520);
nor U1589 (N_1589,N_1508,N_1569);
xor U1590 (N_1590,N_1566,N_1511);
or U1591 (N_1591,N_1573,N_1556);
or U1592 (N_1592,N_1535,N_1572);
nor U1593 (N_1593,N_1500,N_1559);
and U1594 (N_1594,N_1567,N_1561);
or U1595 (N_1595,N_1552,N_1574);
nand U1596 (N_1596,N_1540,N_1512);
and U1597 (N_1597,N_1515,N_1562);
and U1598 (N_1598,N_1523,N_1557);
or U1599 (N_1599,N_1555,N_1505);
nand U1600 (N_1600,N_1509,N_1549);
nand U1601 (N_1601,N_1571,N_1541);
and U1602 (N_1602,N_1530,N_1554);
xor U1603 (N_1603,N_1510,N_1521);
nor U1604 (N_1604,N_1518,N_1506);
or U1605 (N_1605,N_1563,N_1544);
and U1606 (N_1606,N_1526,N_1522);
nand U1607 (N_1607,N_1545,N_1565);
nand U1608 (N_1608,N_1536,N_1532);
nand U1609 (N_1609,N_1533,N_1524);
xnor U1610 (N_1610,N_1529,N_1517);
nand U1611 (N_1611,N_1531,N_1516);
nor U1612 (N_1612,N_1537,N_1513);
and U1613 (N_1613,N_1511,N_1513);
xor U1614 (N_1614,N_1549,N_1572);
nand U1615 (N_1615,N_1502,N_1523);
xor U1616 (N_1616,N_1525,N_1507);
nand U1617 (N_1617,N_1539,N_1523);
nor U1618 (N_1618,N_1557,N_1570);
nor U1619 (N_1619,N_1508,N_1506);
nor U1620 (N_1620,N_1537,N_1565);
xnor U1621 (N_1621,N_1536,N_1506);
or U1622 (N_1622,N_1507,N_1514);
and U1623 (N_1623,N_1528,N_1522);
xnor U1624 (N_1624,N_1572,N_1522);
or U1625 (N_1625,N_1561,N_1555);
nor U1626 (N_1626,N_1525,N_1558);
nor U1627 (N_1627,N_1516,N_1549);
nand U1628 (N_1628,N_1518,N_1511);
nand U1629 (N_1629,N_1545,N_1520);
nand U1630 (N_1630,N_1507,N_1500);
nor U1631 (N_1631,N_1546,N_1570);
or U1632 (N_1632,N_1542,N_1540);
nor U1633 (N_1633,N_1525,N_1535);
nand U1634 (N_1634,N_1544,N_1534);
or U1635 (N_1635,N_1553,N_1569);
or U1636 (N_1636,N_1552,N_1510);
xor U1637 (N_1637,N_1570,N_1573);
or U1638 (N_1638,N_1538,N_1528);
nor U1639 (N_1639,N_1529,N_1514);
or U1640 (N_1640,N_1553,N_1518);
nand U1641 (N_1641,N_1572,N_1541);
xor U1642 (N_1642,N_1526,N_1574);
xor U1643 (N_1643,N_1521,N_1527);
nor U1644 (N_1644,N_1526,N_1562);
nand U1645 (N_1645,N_1509,N_1556);
and U1646 (N_1646,N_1524,N_1540);
nor U1647 (N_1647,N_1521,N_1522);
nor U1648 (N_1648,N_1536,N_1567);
nand U1649 (N_1649,N_1552,N_1514);
nand U1650 (N_1650,N_1613,N_1594);
xor U1651 (N_1651,N_1601,N_1623);
nand U1652 (N_1652,N_1590,N_1585);
nor U1653 (N_1653,N_1617,N_1635);
xnor U1654 (N_1654,N_1605,N_1614);
and U1655 (N_1655,N_1598,N_1588);
xnor U1656 (N_1656,N_1636,N_1589);
nor U1657 (N_1657,N_1584,N_1631);
and U1658 (N_1658,N_1633,N_1586);
or U1659 (N_1659,N_1608,N_1579);
nor U1660 (N_1660,N_1647,N_1610);
and U1661 (N_1661,N_1627,N_1646);
nand U1662 (N_1662,N_1612,N_1628);
or U1663 (N_1663,N_1602,N_1592);
nor U1664 (N_1664,N_1611,N_1643);
or U1665 (N_1665,N_1581,N_1587);
nor U1666 (N_1666,N_1620,N_1578);
nor U1667 (N_1667,N_1576,N_1626);
nor U1668 (N_1668,N_1618,N_1577);
nand U1669 (N_1669,N_1593,N_1591);
nand U1670 (N_1670,N_1645,N_1583);
or U1671 (N_1671,N_1604,N_1575);
and U1672 (N_1672,N_1615,N_1641);
or U1673 (N_1673,N_1595,N_1622);
xor U1674 (N_1674,N_1624,N_1603);
nor U1675 (N_1675,N_1630,N_1580);
nor U1676 (N_1676,N_1644,N_1640);
xor U1677 (N_1677,N_1648,N_1639);
or U1678 (N_1678,N_1621,N_1632);
and U1679 (N_1679,N_1619,N_1607);
nand U1680 (N_1680,N_1609,N_1582);
xor U1681 (N_1681,N_1599,N_1629);
nand U1682 (N_1682,N_1649,N_1606);
nor U1683 (N_1683,N_1600,N_1638);
nand U1684 (N_1684,N_1634,N_1642);
or U1685 (N_1685,N_1616,N_1625);
xor U1686 (N_1686,N_1637,N_1597);
and U1687 (N_1687,N_1596,N_1642);
xor U1688 (N_1688,N_1633,N_1605);
or U1689 (N_1689,N_1614,N_1618);
nor U1690 (N_1690,N_1575,N_1634);
xnor U1691 (N_1691,N_1637,N_1613);
nor U1692 (N_1692,N_1631,N_1637);
and U1693 (N_1693,N_1600,N_1595);
or U1694 (N_1694,N_1641,N_1619);
or U1695 (N_1695,N_1636,N_1639);
nor U1696 (N_1696,N_1588,N_1577);
xnor U1697 (N_1697,N_1622,N_1592);
and U1698 (N_1698,N_1578,N_1642);
and U1699 (N_1699,N_1581,N_1643);
or U1700 (N_1700,N_1584,N_1645);
or U1701 (N_1701,N_1645,N_1639);
and U1702 (N_1702,N_1577,N_1617);
nand U1703 (N_1703,N_1633,N_1597);
nand U1704 (N_1704,N_1617,N_1610);
or U1705 (N_1705,N_1614,N_1637);
or U1706 (N_1706,N_1623,N_1630);
and U1707 (N_1707,N_1637,N_1649);
xnor U1708 (N_1708,N_1595,N_1638);
or U1709 (N_1709,N_1648,N_1632);
xor U1710 (N_1710,N_1615,N_1599);
xnor U1711 (N_1711,N_1646,N_1601);
and U1712 (N_1712,N_1616,N_1600);
nor U1713 (N_1713,N_1591,N_1629);
or U1714 (N_1714,N_1610,N_1605);
nor U1715 (N_1715,N_1620,N_1584);
or U1716 (N_1716,N_1624,N_1586);
or U1717 (N_1717,N_1610,N_1616);
xor U1718 (N_1718,N_1625,N_1575);
or U1719 (N_1719,N_1612,N_1607);
xnor U1720 (N_1720,N_1620,N_1617);
nand U1721 (N_1721,N_1641,N_1582);
or U1722 (N_1722,N_1637,N_1610);
nor U1723 (N_1723,N_1578,N_1615);
nand U1724 (N_1724,N_1611,N_1617);
and U1725 (N_1725,N_1664,N_1714);
and U1726 (N_1726,N_1665,N_1670);
nand U1727 (N_1727,N_1663,N_1654);
and U1728 (N_1728,N_1662,N_1696);
nand U1729 (N_1729,N_1671,N_1653);
and U1730 (N_1730,N_1668,N_1701);
nor U1731 (N_1731,N_1716,N_1712);
nor U1732 (N_1732,N_1658,N_1697);
and U1733 (N_1733,N_1676,N_1723);
xnor U1734 (N_1734,N_1715,N_1678);
and U1735 (N_1735,N_1704,N_1722);
nor U1736 (N_1736,N_1667,N_1680);
or U1737 (N_1737,N_1705,N_1710);
nor U1738 (N_1738,N_1679,N_1657);
nand U1739 (N_1739,N_1675,N_1694);
or U1740 (N_1740,N_1700,N_1719);
or U1741 (N_1741,N_1699,N_1660);
nor U1742 (N_1742,N_1674,N_1703);
nand U1743 (N_1743,N_1688,N_1717);
xnor U1744 (N_1744,N_1709,N_1652);
or U1745 (N_1745,N_1708,N_1661);
nand U1746 (N_1746,N_1691,N_1650);
xnor U1747 (N_1747,N_1689,N_1693);
nor U1748 (N_1748,N_1672,N_1656);
and U1749 (N_1749,N_1666,N_1695);
nand U1750 (N_1750,N_1684,N_1651);
and U1751 (N_1751,N_1655,N_1724);
and U1752 (N_1752,N_1707,N_1686);
xor U1753 (N_1753,N_1659,N_1683);
nor U1754 (N_1754,N_1706,N_1677);
nand U1755 (N_1755,N_1702,N_1698);
nand U1756 (N_1756,N_1711,N_1673);
or U1757 (N_1757,N_1669,N_1685);
xnor U1758 (N_1758,N_1692,N_1720);
or U1759 (N_1759,N_1687,N_1713);
nor U1760 (N_1760,N_1681,N_1690);
or U1761 (N_1761,N_1682,N_1718);
or U1762 (N_1762,N_1721,N_1706);
nand U1763 (N_1763,N_1705,N_1692);
xnor U1764 (N_1764,N_1711,N_1719);
or U1765 (N_1765,N_1658,N_1724);
xor U1766 (N_1766,N_1655,N_1686);
or U1767 (N_1767,N_1668,N_1720);
and U1768 (N_1768,N_1657,N_1722);
or U1769 (N_1769,N_1678,N_1687);
and U1770 (N_1770,N_1702,N_1654);
and U1771 (N_1771,N_1652,N_1684);
nor U1772 (N_1772,N_1665,N_1660);
and U1773 (N_1773,N_1694,N_1692);
nor U1774 (N_1774,N_1721,N_1700);
or U1775 (N_1775,N_1666,N_1652);
and U1776 (N_1776,N_1708,N_1707);
or U1777 (N_1777,N_1669,N_1717);
nand U1778 (N_1778,N_1700,N_1681);
or U1779 (N_1779,N_1673,N_1684);
nor U1780 (N_1780,N_1691,N_1681);
xor U1781 (N_1781,N_1683,N_1681);
or U1782 (N_1782,N_1720,N_1670);
or U1783 (N_1783,N_1684,N_1716);
xnor U1784 (N_1784,N_1655,N_1709);
nand U1785 (N_1785,N_1699,N_1673);
nor U1786 (N_1786,N_1667,N_1692);
nor U1787 (N_1787,N_1660,N_1702);
nor U1788 (N_1788,N_1719,N_1658);
or U1789 (N_1789,N_1705,N_1695);
nor U1790 (N_1790,N_1718,N_1666);
nand U1791 (N_1791,N_1671,N_1722);
nor U1792 (N_1792,N_1664,N_1715);
or U1793 (N_1793,N_1708,N_1673);
nor U1794 (N_1794,N_1693,N_1672);
or U1795 (N_1795,N_1691,N_1713);
xnor U1796 (N_1796,N_1672,N_1674);
nand U1797 (N_1797,N_1717,N_1716);
and U1798 (N_1798,N_1658,N_1666);
or U1799 (N_1799,N_1709,N_1700);
nor U1800 (N_1800,N_1733,N_1759);
and U1801 (N_1801,N_1768,N_1786);
nor U1802 (N_1802,N_1792,N_1781);
xnor U1803 (N_1803,N_1742,N_1771);
xnor U1804 (N_1804,N_1785,N_1755);
and U1805 (N_1805,N_1761,N_1740);
nor U1806 (N_1806,N_1773,N_1763);
nand U1807 (N_1807,N_1789,N_1748);
nand U1808 (N_1808,N_1729,N_1762);
or U1809 (N_1809,N_1725,N_1797);
nand U1810 (N_1810,N_1776,N_1784);
and U1811 (N_1811,N_1752,N_1788);
or U1812 (N_1812,N_1764,N_1727);
nand U1813 (N_1813,N_1737,N_1799);
nand U1814 (N_1814,N_1757,N_1793);
xnor U1815 (N_1815,N_1741,N_1754);
nand U1816 (N_1816,N_1738,N_1790);
and U1817 (N_1817,N_1747,N_1730);
nor U1818 (N_1818,N_1734,N_1749);
and U1819 (N_1819,N_1728,N_1794);
and U1820 (N_1820,N_1743,N_1732);
nor U1821 (N_1821,N_1798,N_1778);
nor U1822 (N_1822,N_1787,N_1791);
and U1823 (N_1823,N_1731,N_1750);
xnor U1824 (N_1824,N_1775,N_1758);
nand U1825 (N_1825,N_1746,N_1756);
xor U1826 (N_1826,N_1783,N_1774);
and U1827 (N_1827,N_1745,N_1772);
nor U1828 (N_1828,N_1766,N_1767);
xor U1829 (N_1829,N_1779,N_1736);
xor U1830 (N_1830,N_1726,N_1770);
xnor U1831 (N_1831,N_1777,N_1739);
nor U1832 (N_1832,N_1795,N_1735);
nand U1833 (N_1833,N_1751,N_1796);
and U1834 (N_1834,N_1760,N_1780);
nand U1835 (N_1835,N_1782,N_1765);
xnor U1836 (N_1836,N_1744,N_1769);
nand U1837 (N_1837,N_1753,N_1773);
xnor U1838 (N_1838,N_1738,N_1753);
nor U1839 (N_1839,N_1791,N_1770);
nand U1840 (N_1840,N_1746,N_1744);
xor U1841 (N_1841,N_1774,N_1761);
and U1842 (N_1842,N_1740,N_1725);
xor U1843 (N_1843,N_1735,N_1740);
xnor U1844 (N_1844,N_1752,N_1750);
and U1845 (N_1845,N_1763,N_1729);
nor U1846 (N_1846,N_1791,N_1757);
xnor U1847 (N_1847,N_1766,N_1764);
and U1848 (N_1848,N_1787,N_1781);
or U1849 (N_1849,N_1748,N_1762);
or U1850 (N_1850,N_1770,N_1785);
xor U1851 (N_1851,N_1793,N_1765);
xor U1852 (N_1852,N_1757,N_1751);
xor U1853 (N_1853,N_1753,N_1789);
nand U1854 (N_1854,N_1755,N_1759);
nor U1855 (N_1855,N_1732,N_1744);
and U1856 (N_1856,N_1743,N_1760);
xnor U1857 (N_1857,N_1733,N_1739);
and U1858 (N_1858,N_1778,N_1738);
and U1859 (N_1859,N_1794,N_1762);
nand U1860 (N_1860,N_1741,N_1756);
or U1861 (N_1861,N_1798,N_1783);
nand U1862 (N_1862,N_1726,N_1773);
nand U1863 (N_1863,N_1785,N_1780);
nor U1864 (N_1864,N_1773,N_1756);
and U1865 (N_1865,N_1763,N_1725);
nor U1866 (N_1866,N_1744,N_1798);
or U1867 (N_1867,N_1734,N_1767);
nand U1868 (N_1868,N_1757,N_1788);
nand U1869 (N_1869,N_1759,N_1743);
nor U1870 (N_1870,N_1782,N_1781);
nand U1871 (N_1871,N_1741,N_1758);
nor U1872 (N_1872,N_1738,N_1775);
xor U1873 (N_1873,N_1727,N_1777);
and U1874 (N_1874,N_1744,N_1774);
nor U1875 (N_1875,N_1802,N_1841);
nand U1876 (N_1876,N_1808,N_1870);
xnor U1877 (N_1877,N_1805,N_1815);
nor U1878 (N_1878,N_1835,N_1864);
and U1879 (N_1879,N_1849,N_1853);
or U1880 (N_1880,N_1844,N_1809);
xnor U1881 (N_1881,N_1834,N_1813);
or U1882 (N_1882,N_1868,N_1843);
xor U1883 (N_1883,N_1816,N_1838);
and U1884 (N_1884,N_1845,N_1842);
or U1885 (N_1885,N_1803,N_1850);
or U1886 (N_1886,N_1867,N_1833);
xor U1887 (N_1887,N_1810,N_1837);
nor U1888 (N_1888,N_1873,N_1857);
or U1889 (N_1889,N_1851,N_1800);
or U1890 (N_1890,N_1861,N_1831);
nor U1891 (N_1891,N_1854,N_1847);
and U1892 (N_1892,N_1822,N_1807);
and U1893 (N_1893,N_1824,N_1866);
and U1894 (N_1894,N_1855,N_1830);
nor U1895 (N_1895,N_1801,N_1856);
or U1896 (N_1896,N_1817,N_1823);
or U1897 (N_1897,N_1806,N_1812);
nand U1898 (N_1898,N_1874,N_1828);
nand U1899 (N_1899,N_1839,N_1865);
and U1900 (N_1900,N_1814,N_1848);
nor U1901 (N_1901,N_1819,N_1862);
and U1902 (N_1902,N_1858,N_1818);
xnor U1903 (N_1903,N_1869,N_1820);
nor U1904 (N_1904,N_1840,N_1821);
nor U1905 (N_1905,N_1811,N_1832);
or U1906 (N_1906,N_1872,N_1859);
nor U1907 (N_1907,N_1804,N_1846);
and U1908 (N_1908,N_1826,N_1825);
and U1909 (N_1909,N_1863,N_1829);
xor U1910 (N_1910,N_1852,N_1871);
or U1911 (N_1911,N_1860,N_1836);
nor U1912 (N_1912,N_1827,N_1874);
or U1913 (N_1913,N_1831,N_1863);
xnor U1914 (N_1914,N_1860,N_1848);
xor U1915 (N_1915,N_1869,N_1801);
or U1916 (N_1916,N_1821,N_1858);
nor U1917 (N_1917,N_1866,N_1827);
nor U1918 (N_1918,N_1873,N_1827);
xor U1919 (N_1919,N_1853,N_1808);
and U1920 (N_1920,N_1835,N_1821);
nand U1921 (N_1921,N_1821,N_1851);
xor U1922 (N_1922,N_1867,N_1853);
xnor U1923 (N_1923,N_1809,N_1851);
nor U1924 (N_1924,N_1872,N_1845);
nor U1925 (N_1925,N_1858,N_1847);
nor U1926 (N_1926,N_1864,N_1844);
nand U1927 (N_1927,N_1809,N_1854);
or U1928 (N_1928,N_1842,N_1817);
nand U1929 (N_1929,N_1868,N_1856);
xor U1930 (N_1930,N_1856,N_1806);
nor U1931 (N_1931,N_1837,N_1816);
nor U1932 (N_1932,N_1869,N_1870);
or U1933 (N_1933,N_1850,N_1820);
xnor U1934 (N_1934,N_1853,N_1812);
nand U1935 (N_1935,N_1814,N_1832);
nor U1936 (N_1936,N_1806,N_1834);
nand U1937 (N_1937,N_1842,N_1810);
or U1938 (N_1938,N_1833,N_1803);
xor U1939 (N_1939,N_1853,N_1872);
and U1940 (N_1940,N_1848,N_1824);
xor U1941 (N_1941,N_1850,N_1832);
or U1942 (N_1942,N_1856,N_1847);
and U1943 (N_1943,N_1830,N_1850);
nand U1944 (N_1944,N_1811,N_1817);
nand U1945 (N_1945,N_1804,N_1814);
and U1946 (N_1946,N_1810,N_1852);
or U1947 (N_1947,N_1822,N_1814);
xor U1948 (N_1948,N_1827,N_1847);
and U1949 (N_1949,N_1807,N_1866);
nand U1950 (N_1950,N_1901,N_1922);
or U1951 (N_1951,N_1909,N_1908);
nand U1952 (N_1952,N_1875,N_1887);
nand U1953 (N_1953,N_1933,N_1943);
and U1954 (N_1954,N_1923,N_1898);
nand U1955 (N_1955,N_1902,N_1876);
and U1956 (N_1956,N_1883,N_1885);
or U1957 (N_1957,N_1888,N_1894);
and U1958 (N_1958,N_1937,N_1947);
nand U1959 (N_1959,N_1919,N_1895);
nor U1960 (N_1960,N_1897,N_1896);
nand U1961 (N_1961,N_1904,N_1926);
and U1962 (N_1962,N_1912,N_1930);
nand U1963 (N_1963,N_1893,N_1940);
nand U1964 (N_1964,N_1877,N_1892);
or U1965 (N_1965,N_1917,N_1927);
xor U1966 (N_1966,N_1915,N_1913);
or U1967 (N_1967,N_1889,N_1882);
and U1968 (N_1968,N_1949,N_1942);
and U1969 (N_1969,N_1928,N_1948);
and U1970 (N_1970,N_1939,N_1890);
or U1971 (N_1971,N_1946,N_1905);
and U1972 (N_1972,N_1881,N_1903);
or U1973 (N_1973,N_1945,N_1935);
nand U1974 (N_1974,N_1932,N_1916);
nor U1975 (N_1975,N_1891,N_1920);
xnor U1976 (N_1976,N_1936,N_1878);
and U1977 (N_1977,N_1934,N_1880);
nand U1978 (N_1978,N_1910,N_1944);
nor U1979 (N_1979,N_1899,N_1879);
nor U1980 (N_1980,N_1929,N_1918);
nor U1981 (N_1981,N_1911,N_1925);
nand U1982 (N_1982,N_1886,N_1906);
nor U1983 (N_1983,N_1884,N_1907);
nor U1984 (N_1984,N_1900,N_1914);
and U1985 (N_1985,N_1924,N_1931);
xnor U1986 (N_1986,N_1938,N_1941);
nor U1987 (N_1987,N_1921,N_1926);
and U1988 (N_1988,N_1885,N_1934);
and U1989 (N_1989,N_1899,N_1885);
nor U1990 (N_1990,N_1935,N_1899);
nor U1991 (N_1991,N_1884,N_1922);
or U1992 (N_1992,N_1919,N_1927);
xor U1993 (N_1993,N_1941,N_1894);
nand U1994 (N_1994,N_1931,N_1927);
and U1995 (N_1995,N_1943,N_1877);
nand U1996 (N_1996,N_1888,N_1903);
nor U1997 (N_1997,N_1937,N_1909);
or U1998 (N_1998,N_1948,N_1915);
and U1999 (N_1999,N_1926,N_1947);
nand U2000 (N_2000,N_1901,N_1936);
nand U2001 (N_2001,N_1900,N_1937);
nand U2002 (N_2002,N_1910,N_1893);
xnor U2003 (N_2003,N_1890,N_1892);
xnor U2004 (N_2004,N_1926,N_1875);
and U2005 (N_2005,N_1886,N_1875);
and U2006 (N_2006,N_1887,N_1885);
nor U2007 (N_2007,N_1884,N_1935);
and U2008 (N_2008,N_1921,N_1910);
xor U2009 (N_2009,N_1922,N_1887);
and U2010 (N_2010,N_1934,N_1922);
xor U2011 (N_2011,N_1913,N_1925);
xnor U2012 (N_2012,N_1891,N_1930);
and U2013 (N_2013,N_1933,N_1908);
or U2014 (N_2014,N_1876,N_1939);
nor U2015 (N_2015,N_1918,N_1924);
nand U2016 (N_2016,N_1943,N_1939);
nor U2017 (N_2017,N_1946,N_1896);
and U2018 (N_2018,N_1899,N_1930);
nand U2019 (N_2019,N_1949,N_1924);
xor U2020 (N_2020,N_1911,N_1895);
and U2021 (N_2021,N_1897,N_1930);
xnor U2022 (N_2022,N_1942,N_1913);
or U2023 (N_2023,N_1899,N_1918);
or U2024 (N_2024,N_1877,N_1932);
or U2025 (N_2025,N_1979,N_1970);
and U2026 (N_2026,N_2016,N_1958);
nor U2027 (N_2027,N_2020,N_1984);
nand U2028 (N_2028,N_1994,N_2005);
nand U2029 (N_2029,N_2007,N_1957);
xor U2030 (N_2030,N_2010,N_1978);
and U2031 (N_2031,N_2009,N_1998);
xnor U2032 (N_2032,N_1951,N_2012);
and U2033 (N_2033,N_1967,N_2023);
and U2034 (N_2034,N_2004,N_1991);
nand U2035 (N_2035,N_1961,N_2018);
nor U2036 (N_2036,N_2019,N_2001);
nand U2037 (N_2037,N_1976,N_1956);
nand U2038 (N_2038,N_1983,N_1975);
or U2039 (N_2039,N_1955,N_1971);
nand U2040 (N_2040,N_1950,N_1988);
xor U2041 (N_2041,N_2000,N_1966);
nand U2042 (N_2042,N_1993,N_2021);
nor U2043 (N_2043,N_1969,N_1973);
and U2044 (N_2044,N_1995,N_1972);
xnor U2045 (N_2045,N_1981,N_1996);
and U2046 (N_2046,N_2014,N_1964);
or U2047 (N_2047,N_1989,N_1982);
or U2048 (N_2048,N_1954,N_2017);
and U2049 (N_2049,N_1985,N_1992);
and U2050 (N_2050,N_1968,N_1965);
xnor U2051 (N_2051,N_2013,N_1959);
and U2052 (N_2052,N_1999,N_2024);
nor U2053 (N_2053,N_2008,N_1952);
or U2054 (N_2054,N_1986,N_1960);
nor U2055 (N_2055,N_1990,N_2015);
nor U2056 (N_2056,N_1980,N_1997);
nand U2057 (N_2057,N_2006,N_1962);
or U2058 (N_2058,N_2022,N_1953);
nand U2059 (N_2059,N_2011,N_2003);
nor U2060 (N_2060,N_1987,N_1963);
xnor U2061 (N_2061,N_1977,N_1974);
xor U2062 (N_2062,N_2002,N_2019);
xnor U2063 (N_2063,N_1997,N_1979);
and U2064 (N_2064,N_2010,N_1996);
nor U2065 (N_2065,N_1966,N_1962);
and U2066 (N_2066,N_1959,N_1966);
nand U2067 (N_2067,N_1994,N_1974);
xor U2068 (N_2068,N_2014,N_1996);
nor U2069 (N_2069,N_1996,N_2017);
and U2070 (N_2070,N_1990,N_2018);
nor U2071 (N_2071,N_1983,N_1952);
xor U2072 (N_2072,N_2002,N_2020);
nand U2073 (N_2073,N_2003,N_1967);
nand U2074 (N_2074,N_1996,N_1964);
nor U2075 (N_2075,N_2023,N_1982);
and U2076 (N_2076,N_1986,N_1984);
nand U2077 (N_2077,N_1953,N_1955);
or U2078 (N_2078,N_1968,N_1962);
nor U2079 (N_2079,N_2019,N_2010);
xnor U2080 (N_2080,N_1992,N_1970);
or U2081 (N_2081,N_2002,N_1997);
nor U2082 (N_2082,N_1973,N_1959);
xnor U2083 (N_2083,N_2016,N_1998);
nor U2084 (N_2084,N_2007,N_1971);
nor U2085 (N_2085,N_1999,N_1964);
nor U2086 (N_2086,N_1990,N_2023);
or U2087 (N_2087,N_1992,N_2018);
and U2088 (N_2088,N_1967,N_1959);
or U2089 (N_2089,N_2010,N_2008);
xor U2090 (N_2090,N_1979,N_2023);
and U2091 (N_2091,N_1988,N_2002);
nand U2092 (N_2092,N_1997,N_1969);
or U2093 (N_2093,N_2023,N_1977);
or U2094 (N_2094,N_1950,N_2006);
xnor U2095 (N_2095,N_1976,N_1962);
nand U2096 (N_2096,N_1997,N_2021);
or U2097 (N_2097,N_1983,N_2020);
or U2098 (N_2098,N_1983,N_1962);
nand U2099 (N_2099,N_2018,N_1982);
or U2100 (N_2100,N_2028,N_2045);
or U2101 (N_2101,N_2046,N_2093);
nand U2102 (N_2102,N_2084,N_2083);
xnor U2103 (N_2103,N_2079,N_2048);
and U2104 (N_2104,N_2034,N_2066);
nand U2105 (N_2105,N_2096,N_2080);
and U2106 (N_2106,N_2072,N_2067);
or U2107 (N_2107,N_2041,N_2065);
xnor U2108 (N_2108,N_2090,N_2095);
and U2109 (N_2109,N_2099,N_2087);
nor U2110 (N_2110,N_2085,N_2092);
and U2111 (N_2111,N_2058,N_2064);
xor U2112 (N_2112,N_2055,N_2073);
nor U2113 (N_2113,N_2053,N_2033);
or U2114 (N_2114,N_2071,N_2039);
nor U2115 (N_2115,N_2040,N_2070);
nand U2116 (N_2116,N_2057,N_2091);
xnor U2117 (N_2117,N_2075,N_2038);
and U2118 (N_2118,N_2059,N_2054);
nor U2119 (N_2119,N_2069,N_2030);
nor U2120 (N_2120,N_2051,N_2037);
or U2121 (N_2121,N_2089,N_2047);
nand U2122 (N_2122,N_2027,N_2078);
or U2123 (N_2123,N_2060,N_2077);
xor U2124 (N_2124,N_2076,N_2074);
and U2125 (N_2125,N_2068,N_2026);
nand U2126 (N_2126,N_2098,N_2063);
xor U2127 (N_2127,N_2035,N_2082);
or U2128 (N_2128,N_2081,N_2097);
xor U2129 (N_2129,N_2061,N_2050);
xnor U2130 (N_2130,N_2086,N_2025);
nor U2131 (N_2131,N_2049,N_2088);
or U2132 (N_2132,N_2043,N_2044);
and U2133 (N_2133,N_2056,N_2052);
xor U2134 (N_2134,N_2062,N_2094);
and U2135 (N_2135,N_2032,N_2029);
nand U2136 (N_2136,N_2031,N_2042);
nor U2137 (N_2137,N_2036,N_2090);
or U2138 (N_2138,N_2053,N_2027);
xor U2139 (N_2139,N_2084,N_2075);
or U2140 (N_2140,N_2078,N_2032);
nor U2141 (N_2141,N_2079,N_2061);
and U2142 (N_2142,N_2064,N_2037);
nand U2143 (N_2143,N_2037,N_2068);
and U2144 (N_2144,N_2091,N_2033);
xnor U2145 (N_2145,N_2095,N_2088);
xnor U2146 (N_2146,N_2030,N_2047);
nor U2147 (N_2147,N_2037,N_2085);
xnor U2148 (N_2148,N_2027,N_2086);
xor U2149 (N_2149,N_2071,N_2076);
nor U2150 (N_2150,N_2049,N_2047);
or U2151 (N_2151,N_2087,N_2078);
nor U2152 (N_2152,N_2034,N_2035);
and U2153 (N_2153,N_2089,N_2071);
and U2154 (N_2154,N_2059,N_2083);
and U2155 (N_2155,N_2032,N_2051);
and U2156 (N_2156,N_2073,N_2067);
xnor U2157 (N_2157,N_2079,N_2031);
or U2158 (N_2158,N_2027,N_2043);
or U2159 (N_2159,N_2075,N_2045);
nor U2160 (N_2160,N_2088,N_2072);
nand U2161 (N_2161,N_2066,N_2042);
xnor U2162 (N_2162,N_2092,N_2056);
xor U2163 (N_2163,N_2074,N_2064);
nand U2164 (N_2164,N_2088,N_2061);
or U2165 (N_2165,N_2082,N_2079);
nand U2166 (N_2166,N_2096,N_2063);
xor U2167 (N_2167,N_2072,N_2040);
or U2168 (N_2168,N_2040,N_2042);
xor U2169 (N_2169,N_2054,N_2032);
nor U2170 (N_2170,N_2077,N_2047);
or U2171 (N_2171,N_2058,N_2093);
xor U2172 (N_2172,N_2076,N_2031);
nor U2173 (N_2173,N_2092,N_2027);
nand U2174 (N_2174,N_2070,N_2079);
xnor U2175 (N_2175,N_2126,N_2147);
and U2176 (N_2176,N_2130,N_2163);
or U2177 (N_2177,N_2160,N_2113);
and U2178 (N_2178,N_2156,N_2139);
and U2179 (N_2179,N_2125,N_2134);
xor U2180 (N_2180,N_2157,N_2166);
nor U2181 (N_2181,N_2119,N_2124);
nand U2182 (N_2182,N_2109,N_2158);
nand U2183 (N_2183,N_2149,N_2116);
nor U2184 (N_2184,N_2105,N_2135);
xnor U2185 (N_2185,N_2172,N_2137);
xor U2186 (N_2186,N_2122,N_2114);
or U2187 (N_2187,N_2123,N_2118);
xor U2188 (N_2188,N_2167,N_2132);
and U2189 (N_2189,N_2111,N_2150);
xnor U2190 (N_2190,N_2169,N_2117);
xnor U2191 (N_2191,N_2141,N_2171);
and U2192 (N_2192,N_2108,N_2143);
xor U2193 (N_2193,N_2144,N_2153);
xor U2194 (N_2194,N_2129,N_2127);
and U2195 (N_2195,N_2110,N_2104);
and U2196 (N_2196,N_2148,N_2131);
nand U2197 (N_2197,N_2115,N_2112);
and U2198 (N_2198,N_2100,N_2121);
xnor U2199 (N_2199,N_2162,N_2106);
nand U2200 (N_2200,N_2174,N_2152);
nor U2201 (N_2201,N_2164,N_2146);
or U2202 (N_2202,N_2159,N_2142);
xnor U2203 (N_2203,N_2155,N_2154);
nor U2204 (N_2204,N_2138,N_2168);
nand U2205 (N_2205,N_2170,N_2133);
nand U2206 (N_2206,N_2145,N_2128);
xnor U2207 (N_2207,N_2151,N_2107);
xor U2208 (N_2208,N_2103,N_2136);
or U2209 (N_2209,N_2165,N_2173);
nor U2210 (N_2210,N_2161,N_2120);
nand U2211 (N_2211,N_2101,N_2140);
xnor U2212 (N_2212,N_2102,N_2132);
nor U2213 (N_2213,N_2126,N_2149);
or U2214 (N_2214,N_2117,N_2133);
xor U2215 (N_2215,N_2122,N_2124);
and U2216 (N_2216,N_2145,N_2137);
nand U2217 (N_2217,N_2121,N_2164);
nand U2218 (N_2218,N_2166,N_2120);
nor U2219 (N_2219,N_2121,N_2117);
or U2220 (N_2220,N_2138,N_2101);
nor U2221 (N_2221,N_2165,N_2129);
or U2222 (N_2222,N_2163,N_2129);
nor U2223 (N_2223,N_2153,N_2141);
nor U2224 (N_2224,N_2156,N_2132);
or U2225 (N_2225,N_2137,N_2154);
and U2226 (N_2226,N_2102,N_2107);
nor U2227 (N_2227,N_2142,N_2124);
or U2228 (N_2228,N_2131,N_2157);
xnor U2229 (N_2229,N_2159,N_2130);
or U2230 (N_2230,N_2110,N_2137);
xor U2231 (N_2231,N_2154,N_2162);
nand U2232 (N_2232,N_2115,N_2116);
or U2233 (N_2233,N_2138,N_2113);
xnor U2234 (N_2234,N_2114,N_2110);
xor U2235 (N_2235,N_2104,N_2137);
or U2236 (N_2236,N_2124,N_2108);
or U2237 (N_2237,N_2148,N_2159);
nand U2238 (N_2238,N_2162,N_2166);
and U2239 (N_2239,N_2131,N_2140);
or U2240 (N_2240,N_2149,N_2150);
nand U2241 (N_2241,N_2139,N_2114);
nand U2242 (N_2242,N_2108,N_2174);
nand U2243 (N_2243,N_2151,N_2135);
nor U2244 (N_2244,N_2140,N_2141);
nor U2245 (N_2245,N_2160,N_2102);
nor U2246 (N_2246,N_2115,N_2129);
and U2247 (N_2247,N_2128,N_2131);
nand U2248 (N_2248,N_2168,N_2152);
xor U2249 (N_2249,N_2118,N_2107);
nor U2250 (N_2250,N_2218,N_2215);
and U2251 (N_2251,N_2248,N_2237);
or U2252 (N_2252,N_2236,N_2221);
nor U2253 (N_2253,N_2180,N_2232);
or U2254 (N_2254,N_2207,N_2200);
xor U2255 (N_2255,N_2183,N_2220);
or U2256 (N_2256,N_2210,N_2204);
nor U2257 (N_2257,N_2192,N_2205);
nand U2258 (N_2258,N_2189,N_2198);
or U2259 (N_2259,N_2203,N_2178);
or U2260 (N_2260,N_2185,N_2222);
or U2261 (N_2261,N_2177,N_2249);
or U2262 (N_2262,N_2233,N_2219);
nor U2263 (N_2263,N_2216,N_2226);
nor U2264 (N_2264,N_2190,N_2196);
nor U2265 (N_2265,N_2175,N_2208);
or U2266 (N_2266,N_2212,N_2247);
or U2267 (N_2267,N_2201,N_2197);
or U2268 (N_2268,N_2195,N_2224);
nor U2269 (N_2269,N_2217,N_2223);
xnor U2270 (N_2270,N_2239,N_2244);
nand U2271 (N_2271,N_2238,N_2243);
xnor U2272 (N_2272,N_2246,N_2186);
or U2273 (N_2273,N_2191,N_2202);
nor U2274 (N_2274,N_2184,N_2245);
xnor U2275 (N_2275,N_2188,N_2179);
xnor U2276 (N_2276,N_2194,N_2242);
nand U2277 (N_2277,N_2231,N_2206);
or U2278 (N_2278,N_2229,N_2240);
or U2279 (N_2279,N_2193,N_2182);
and U2280 (N_2280,N_2209,N_2225);
nor U2281 (N_2281,N_2187,N_2214);
and U2282 (N_2282,N_2241,N_2228);
nor U2283 (N_2283,N_2213,N_2181);
nand U2284 (N_2284,N_2234,N_2230);
and U2285 (N_2285,N_2235,N_2199);
nand U2286 (N_2286,N_2176,N_2211);
or U2287 (N_2287,N_2227,N_2230);
and U2288 (N_2288,N_2186,N_2195);
or U2289 (N_2289,N_2175,N_2219);
nand U2290 (N_2290,N_2228,N_2236);
and U2291 (N_2291,N_2187,N_2212);
xnor U2292 (N_2292,N_2214,N_2222);
or U2293 (N_2293,N_2205,N_2249);
nand U2294 (N_2294,N_2176,N_2234);
nor U2295 (N_2295,N_2215,N_2222);
or U2296 (N_2296,N_2215,N_2214);
or U2297 (N_2297,N_2193,N_2185);
and U2298 (N_2298,N_2222,N_2183);
nor U2299 (N_2299,N_2211,N_2249);
or U2300 (N_2300,N_2181,N_2216);
and U2301 (N_2301,N_2248,N_2241);
nor U2302 (N_2302,N_2207,N_2239);
and U2303 (N_2303,N_2198,N_2204);
or U2304 (N_2304,N_2246,N_2183);
or U2305 (N_2305,N_2196,N_2231);
xor U2306 (N_2306,N_2178,N_2184);
and U2307 (N_2307,N_2190,N_2217);
nand U2308 (N_2308,N_2223,N_2226);
nor U2309 (N_2309,N_2188,N_2232);
and U2310 (N_2310,N_2235,N_2195);
nand U2311 (N_2311,N_2205,N_2225);
nor U2312 (N_2312,N_2216,N_2196);
and U2313 (N_2313,N_2188,N_2247);
or U2314 (N_2314,N_2203,N_2179);
xor U2315 (N_2315,N_2235,N_2229);
xnor U2316 (N_2316,N_2243,N_2217);
nor U2317 (N_2317,N_2183,N_2236);
or U2318 (N_2318,N_2223,N_2228);
xor U2319 (N_2319,N_2219,N_2216);
nand U2320 (N_2320,N_2205,N_2221);
and U2321 (N_2321,N_2233,N_2199);
or U2322 (N_2322,N_2202,N_2242);
nor U2323 (N_2323,N_2229,N_2239);
nand U2324 (N_2324,N_2185,N_2204);
and U2325 (N_2325,N_2302,N_2265);
nand U2326 (N_2326,N_2285,N_2316);
nor U2327 (N_2327,N_2277,N_2296);
xnor U2328 (N_2328,N_2255,N_2250);
nor U2329 (N_2329,N_2309,N_2297);
or U2330 (N_2330,N_2313,N_2260);
and U2331 (N_2331,N_2266,N_2315);
nor U2332 (N_2332,N_2291,N_2253);
nor U2333 (N_2333,N_2301,N_2270);
xnor U2334 (N_2334,N_2319,N_2308);
xor U2335 (N_2335,N_2281,N_2256);
xor U2336 (N_2336,N_2298,N_2286);
or U2337 (N_2337,N_2274,N_2310);
or U2338 (N_2338,N_2269,N_2263);
nor U2339 (N_2339,N_2320,N_2314);
xnor U2340 (N_2340,N_2311,N_2312);
and U2341 (N_2341,N_2307,N_2258);
or U2342 (N_2342,N_2271,N_2305);
or U2343 (N_2343,N_2304,N_2318);
and U2344 (N_2344,N_2321,N_2273);
nor U2345 (N_2345,N_2306,N_2292);
xor U2346 (N_2346,N_2279,N_2280);
and U2347 (N_2347,N_2283,N_2268);
xnor U2348 (N_2348,N_2252,N_2264);
nand U2349 (N_2349,N_2254,N_2278);
xor U2350 (N_2350,N_2276,N_2293);
nor U2351 (N_2351,N_2288,N_2272);
and U2352 (N_2352,N_2317,N_2299);
nand U2353 (N_2353,N_2262,N_2294);
and U2354 (N_2354,N_2261,N_2300);
xor U2355 (N_2355,N_2324,N_2290);
and U2356 (N_2356,N_2282,N_2259);
nand U2357 (N_2357,N_2322,N_2287);
xor U2358 (N_2358,N_2257,N_2275);
or U2359 (N_2359,N_2284,N_2323);
nor U2360 (N_2360,N_2295,N_2267);
nand U2361 (N_2361,N_2289,N_2303);
or U2362 (N_2362,N_2251,N_2300);
or U2363 (N_2363,N_2295,N_2269);
nand U2364 (N_2364,N_2304,N_2263);
xor U2365 (N_2365,N_2262,N_2320);
nand U2366 (N_2366,N_2301,N_2288);
nor U2367 (N_2367,N_2263,N_2318);
nor U2368 (N_2368,N_2254,N_2282);
nand U2369 (N_2369,N_2295,N_2263);
and U2370 (N_2370,N_2252,N_2272);
and U2371 (N_2371,N_2320,N_2305);
nor U2372 (N_2372,N_2277,N_2294);
and U2373 (N_2373,N_2263,N_2288);
nand U2374 (N_2374,N_2280,N_2315);
nand U2375 (N_2375,N_2253,N_2285);
nand U2376 (N_2376,N_2299,N_2324);
or U2377 (N_2377,N_2318,N_2279);
or U2378 (N_2378,N_2300,N_2287);
and U2379 (N_2379,N_2288,N_2292);
and U2380 (N_2380,N_2287,N_2296);
xor U2381 (N_2381,N_2291,N_2306);
xnor U2382 (N_2382,N_2313,N_2285);
nor U2383 (N_2383,N_2317,N_2315);
xor U2384 (N_2384,N_2308,N_2253);
nor U2385 (N_2385,N_2268,N_2255);
nor U2386 (N_2386,N_2316,N_2286);
and U2387 (N_2387,N_2317,N_2258);
and U2388 (N_2388,N_2302,N_2263);
nor U2389 (N_2389,N_2319,N_2324);
xor U2390 (N_2390,N_2257,N_2288);
and U2391 (N_2391,N_2270,N_2297);
nand U2392 (N_2392,N_2322,N_2317);
or U2393 (N_2393,N_2312,N_2283);
nand U2394 (N_2394,N_2313,N_2320);
nand U2395 (N_2395,N_2262,N_2317);
nand U2396 (N_2396,N_2296,N_2267);
nor U2397 (N_2397,N_2294,N_2279);
xnor U2398 (N_2398,N_2311,N_2297);
or U2399 (N_2399,N_2317,N_2298);
and U2400 (N_2400,N_2359,N_2375);
or U2401 (N_2401,N_2380,N_2395);
and U2402 (N_2402,N_2332,N_2360);
or U2403 (N_2403,N_2330,N_2376);
nor U2404 (N_2404,N_2329,N_2327);
nand U2405 (N_2405,N_2334,N_2393);
nand U2406 (N_2406,N_2388,N_2397);
nor U2407 (N_2407,N_2326,N_2355);
and U2408 (N_2408,N_2386,N_2382);
nand U2409 (N_2409,N_2371,N_2384);
nor U2410 (N_2410,N_2362,N_2361);
or U2411 (N_2411,N_2353,N_2348);
and U2412 (N_2412,N_2373,N_2356);
xnor U2413 (N_2413,N_2363,N_2339);
and U2414 (N_2414,N_2383,N_2340);
or U2415 (N_2415,N_2350,N_2344);
nor U2416 (N_2416,N_2367,N_2366);
xnor U2417 (N_2417,N_2372,N_2399);
nand U2418 (N_2418,N_2335,N_2392);
and U2419 (N_2419,N_2368,N_2378);
xnor U2420 (N_2420,N_2333,N_2396);
nand U2421 (N_2421,N_2351,N_2352);
xor U2422 (N_2422,N_2357,N_2387);
or U2423 (N_2423,N_2394,N_2342);
nand U2424 (N_2424,N_2379,N_2377);
xnor U2425 (N_2425,N_2325,N_2389);
nor U2426 (N_2426,N_2337,N_2328);
nor U2427 (N_2427,N_2369,N_2358);
or U2428 (N_2428,N_2341,N_2354);
and U2429 (N_2429,N_2336,N_2346);
and U2430 (N_2430,N_2364,N_2398);
xor U2431 (N_2431,N_2385,N_2331);
nor U2432 (N_2432,N_2365,N_2349);
and U2433 (N_2433,N_2390,N_2391);
nand U2434 (N_2434,N_2370,N_2381);
and U2435 (N_2435,N_2347,N_2338);
or U2436 (N_2436,N_2345,N_2343);
and U2437 (N_2437,N_2374,N_2353);
xnor U2438 (N_2438,N_2399,N_2373);
xor U2439 (N_2439,N_2357,N_2378);
and U2440 (N_2440,N_2392,N_2378);
nand U2441 (N_2441,N_2335,N_2339);
nor U2442 (N_2442,N_2362,N_2329);
xor U2443 (N_2443,N_2334,N_2374);
or U2444 (N_2444,N_2350,N_2325);
nand U2445 (N_2445,N_2351,N_2399);
xor U2446 (N_2446,N_2378,N_2374);
or U2447 (N_2447,N_2391,N_2327);
nand U2448 (N_2448,N_2356,N_2355);
nand U2449 (N_2449,N_2346,N_2371);
or U2450 (N_2450,N_2352,N_2364);
xnor U2451 (N_2451,N_2346,N_2351);
nor U2452 (N_2452,N_2362,N_2392);
and U2453 (N_2453,N_2340,N_2329);
xor U2454 (N_2454,N_2351,N_2392);
and U2455 (N_2455,N_2332,N_2362);
nand U2456 (N_2456,N_2367,N_2329);
nor U2457 (N_2457,N_2367,N_2378);
nor U2458 (N_2458,N_2379,N_2337);
or U2459 (N_2459,N_2339,N_2328);
nor U2460 (N_2460,N_2362,N_2395);
or U2461 (N_2461,N_2325,N_2347);
xnor U2462 (N_2462,N_2328,N_2353);
or U2463 (N_2463,N_2329,N_2379);
xnor U2464 (N_2464,N_2350,N_2373);
nand U2465 (N_2465,N_2361,N_2333);
nor U2466 (N_2466,N_2364,N_2363);
nand U2467 (N_2467,N_2389,N_2336);
xor U2468 (N_2468,N_2327,N_2360);
nand U2469 (N_2469,N_2368,N_2397);
and U2470 (N_2470,N_2366,N_2359);
xnor U2471 (N_2471,N_2387,N_2353);
nand U2472 (N_2472,N_2376,N_2383);
and U2473 (N_2473,N_2346,N_2352);
or U2474 (N_2474,N_2360,N_2361);
nor U2475 (N_2475,N_2472,N_2418);
xor U2476 (N_2476,N_2411,N_2406);
and U2477 (N_2477,N_2471,N_2458);
nor U2478 (N_2478,N_2473,N_2415);
and U2479 (N_2479,N_2456,N_2455);
xor U2480 (N_2480,N_2459,N_2463);
or U2481 (N_2481,N_2462,N_2461);
nand U2482 (N_2482,N_2443,N_2416);
xnor U2483 (N_2483,N_2470,N_2407);
xor U2484 (N_2484,N_2434,N_2445);
nor U2485 (N_2485,N_2431,N_2405);
or U2486 (N_2486,N_2450,N_2408);
xor U2487 (N_2487,N_2469,N_2444);
xor U2488 (N_2488,N_2464,N_2452);
or U2489 (N_2489,N_2446,N_2453);
xor U2490 (N_2490,N_2403,N_2467);
nor U2491 (N_2491,N_2441,N_2460);
nand U2492 (N_2492,N_2420,N_2413);
nor U2493 (N_2493,N_2448,N_2412);
and U2494 (N_2494,N_2465,N_2402);
and U2495 (N_2495,N_2410,N_2435);
nor U2496 (N_2496,N_2430,N_2424);
nand U2497 (N_2497,N_2400,N_2427);
or U2498 (N_2498,N_2423,N_2422);
xnor U2499 (N_2499,N_2437,N_2447);
or U2500 (N_2500,N_2401,N_2442);
and U2501 (N_2501,N_2417,N_2439);
xnor U2502 (N_2502,N_2404,N_2466);
nand U2503 (N_2503,N_2426,N_2451);
nor U2504 (N_2504,N_2438,N_2449);
nand U2505 (N_2505,N_2428,N_2474);
or U2506 (N_2506,N_2433,N_2419);
and U2507 (N_2507,N_2414,N_2457);
and U2508 (N_2508,N_2432,N_2409);
xor U2509 (N_2509,N_2425,N_2454);
and U2510 (N_2510,N_2440,N_2421);
xor U2511 (N_2511,N_2468,N_2436);
or U2512 (N_2512,N_2429,N_2465);
nand U2513 (N_2513,N_2453,N_2448);
nor U2514 (N_2514,N_2469,N_2463);
xor U2515 (N_2515,N_2407,N_2426);
nor U2516 (N_2516,N_2453,N_2464);
nor U2517 (N_2517,N_2456,N_2437);
nand U2518 (N_2518,N_2468,N_2403);
nor U2519 (N_2519,N_2421,N_2469);
and U2520 (N_2520,N_2431,N_2458);
or U2521 (N_2521,N_2461,N_2416);
or U2522 (N_2522,N_2403,N_2446);
nand U2523 (N_2523,N_2400,N_2432);
and U2524 (N_2524,N_2407,N_2462);
or U2525 (N_2525,N_2446,N_2456);
xor U2526 (N_2526,N_2467,N_2442);
xnor U2527 (N_2527,N_2439,N_2418);
nor U2528 (N_2528,N_2462,N_2409);
nand U2529 (N_2529,N_2435,N_2405);
nor U2530 (N_2530,N_2436,N_2448);
xnor U2531 (N_2531,N_2409,N_2456);
xor U2532 (N_2532,N_2421,N_2462);
or U2533 (N_2533,N_2439,N_2438);
nor U2534 (N_2534,N_2458,N_2405);
or U2535 (N_2535,N_2425,N_2462);
nand U2536 (N_2536,N_2452,N_2449);
xnor U2537 (N_2537,N_2447,N_2421);
and U2538 (N_2538,N_2466,N_2461);
or U2539 (N_2539,N_2424,N_2441);
nand U2540 (N_2540,N_2456,N_2425);
or U2541 (N_2541,N_2470,N_2465);
or U2542 (N_2542,N_2454,N_2435);
xnor U2543 (N_2543,N_2429,N_2471);
or U2544 (N_2544,N_2471,N_2427);
and U2545 (N_2545,N_2461,N_2438);
nor U2546 (N_2546,N_2435,N_2411);
nor U2547 (N_2547,N_2440,N_2402);
nor U2548 (N_2548,N_2412,N_2442);
nand U2549 (N_2549,N_2428,N_2429);
nand U2550 (N_2550,N_2537,N_2510);
or U2551 (N_2551,N_2482,N_2496);
or U2552 (N_2552,N_2475,N_2514);
and U2553 (N_2553,N_2546,N_2505);
or U2554 (N_2554,N_2536,N_2540);
nor U2555 (N_2555,N_2490,N_2521);
xor U2556 (N_2556,N_2549,N_2499);
nand U2557 (N_2557,N_2547,N_2544);
nand U2558 (N_2558,N_2479,N_2526);
or U2559 (N_2559,N_2507,N_2495);
nand U2560 (N_2560,N_2515,N_2511);
nor U2561 (N_2561,N_2532,N_2483);
xor U2562 (N_2562,N_2517,N_2486);
and U2563 (N_2563,N_2516,N_2485);
nor U2564 (N_2564,N_2502,N_2524);
and U2565 (N_2565,N_2477,N_2493);
nand U2566 (N_2566,N_2506,N_2520);
xor U2567 (N_2567,N_2518,N_2528);
nand U2568 (N_2568,N_2497,N_2545);
nor U2569 (N_2569,N_2478,N_2480);
or U2570 (N_2570,N_2503,N_2530);
or U2571 (N_2571,N_2500,N_2476);
or U2572 (N_2572,N_2535,N_2508);
and U2573 (N_2573,N_2491,N_2541);
xor U2574 (N_2574,N_2525,N_2513);
nor U2575 (N_2575,N_2542,N_2539);
nand U2576 (N_2576,N_2519,N_2501);
nand U2577 (N_2577,N_2512,N_2523);
nor U2578 (N_2578,N_2504,N_2492);
nand U2579 (N_2579,N_2543,N_2527);
and U2580 (N_2580,N_2498,N_2489);
or U2581 (N_2581,N_2487,N_2531);
or U2582 (N_2582,N_2529,N_2481);
nand U2583 (N_2583,N_2534,N_2548);
nand U2584 (N_2584,N_2484,N_2509);
xor U2585 (N_2585,N_2494,N_2533);
nand U2586 (N_2586,N_2538,N_2522);
and U2587 (N_2587,N_2488,N_2480);
nand U2588 (N_2588,N_2512,N_2476);
nand U2589 (N_2589,N_2540,N_2518);
nor U2590 (N_2590,N_2478,N_2486);
and U2591 (N_2591,N_2516,N_2518);
xnor U2592 (N_2592,N_2522,N_2528);
nor U2593 (N_2593,N_2540,N_2515);
nor U2594 (N_2594,N_2509,N_2511);
nor U2595 (N_2595,N_2541,N_2481);
or U2596 (N_2596,N_2489,N_2475);
and U2597 (N_2597,N_2486,N_2497);
nor U2598 (N_2598,N_2527,N_2482);
nor U2599 (N_2599,N_2515,N_2520);
nand U2600 (N_2600,N_2542,N_2475);
xnor U2601 (N_2601,N_2506,N_2482);
xor U2602 (N_2602,N_2538,N_2510);
xor U2603 (N_2603,N_2535,N_2477);
and U2604 (N_2604,N_2542,N_2507);
xor U2605 (N_2605,N_2521,N_2481);
xnor U2606 (N_2606,N_2503,N_2533);
or U2607 (N_2607,N_2489,N_2540);
or U2608 (N_2608,N_2535,N_2548);
xor U2609 (N_2609,N_2478,N_2548);
nand U2610 (N_2610,N_2480,N_2498);
and U2611 (N_2611,N_2519,N_2487);
xor U2612 (N_2612,N_2503,N_2509);
xnor U2613 (N_2613,N_2481,N_2495);
nand U2614 (N_2614,N_2530,N_2495);
or U2615 (N_2615,N_2485,N_2524);
xnor U2616 (N_2616,N_2494,N_2491);
or U2617 (N_2617,N_2488,N_2485);
and U2618 (N_2618,N_2509,N_2482);
nand U2619 (N_2619,N_2548,N_2514);
or U2620 (N_2620,N_2491,N_2535);
or U2621 (N_2621,N_2505,N_2502);
xor U2622 (N_2622,N_2518,N_2524);
xnor U2623 (N_2623,N_2483,N_2503);
nor U2624 (N_2624,N_2535,N_2481);
nor U2625 (N_2625,N_2563,N_2568);
and U2626 (N_2626,N_2586,N_2553);
or U2627 (N_2627,N_2616,N_2598);
xnor U2628 (N_2628,N_2591,N_2613);
or U2629 (N_2629,N_2567,N_2585);
and U2630 (N_2630,N_2601,N_2605);
xor U2631 (N_2631,N_2608,N_2570);
or U2632 (N_2632,N_2577,N_2581);
and U2633 (N_2633,N_2590,N_2603);
and U2634 (N_2634,N_2597,N_2596);
xnor U2635 (N_2635,N_2622,N_2587);
and U2636 (N_2636,N_2595,N_2610);
and U2637 (N_2637,N_2588,N_2579);
nand U2638 (N_2638,N_2594,N_2551);
and U2639 (N_2639,N_2600,N_2584);
and U2640 (N_2640,N_2578,N_2560);
xnor U2641 (N_2641,N_2556,N_2607);
nand U2642 (N_2642,N_2561,N_2604);
xor U2643 (N_2643,N_2559,N_2602);
and U2644 (N_2644,N_2623,N_2565);
nand U2645 (N_2645,N_2614,N_2620);
and U2646 (N_2646,N_2583,N_2624);
or U2647 (N_2647,N_2569,N_2606);
nor U2648 (N_2648,N_2599,N_2617);
xor U2649 (N_2649,N_2564,N_2582);
and U2650 (N_2650,N_2621,N_2571);
xor U2651 (N_2651,N_2618,N_2615);
or U2652 (N_2652,N_2566,N_2576);
or U2653 (N_2653,N_2558,N_2612);
or U2654 (N_2654,N_2550,N_2592);
nand U2655 (N_2655,N_2552,N_2574);
or U2656 (N_2656,N_2573,N_2562);
or U2657 (N_2657,N_2611,N_2619);
nor U2658 (N_2658,N_2572,N_2557);
nand U2659 (N_2659,N_2609,N_2580);
nand U2660 (N_2660,N_2593,N_2589);
or U2661 (N_2661,N_2555,N_2575);
nand U2662 (N_2662,N_2554,N_2556);
nor U2663 (N_2663,N_2582,N_2592);
nor U2664 (N_2664,N_2581,N_2564);
xnor U2665 (N_2665,N_2577,N_2612);
or U2666 (N_2666,N_2585,N_2584);
xnor U2667 (N_2667,N_2589,N_2573);
or U2668 (N_2668,N_2606,N_2573);
and U2669 (N_2669,N_2615,N_2599);
nand U2670 (N_2670,N_2621,N_2604);
and U2671 (N_2671,N_2554,N_2614);
nor U2672 (N_2672,N_2606,N_2603);
xnor U2673 (N_2673,N_2584,N_2568);
xor U2674 (N_2674,N_2607,N_2597);
nor U2675 (N_2675,N_2608,N_2578);
or U2676 (N_2676,N_2576,N_2592);
xor U2677 (N_2677,N_2562,N_2616);
nor U2678 (N_2678,N_2568,N_2599);
xor U2679 (N_2679,N_2624,N_2603);
nand U2680 (N_2680,N_2577,N_2613);
xnor U2681 (N_2681,N_2569,N_2609);
nor U2682 (N_2682,N_2622,N_2612);
xor U2683 (N_2683,N_2557,N_2617);
or U2684 (N_2684,N_2582,N_2600);
nand U2685 (N_2685,N_2582,N_2559);
nand U2686 (N_2686,N_2597,N_2603);
and U2687 (N_2687,N_2599,N_2576);
xnor U2688 (N_2688,N_2624,N_2580);
nand U2689 (N_2689,N_2601,N_2580);
and U2690 (N_2690,N_2616,N_2580);
nor U2691 (N_2691,N_2578,N_2617);
or U2692 (N_2692,N_2593,N_2591);
nand U2693 (N_2693,N_2623,N_2576);
nor U2694 (N_2694,N_2573,N_2623);
and U2695 (N_2695,N_2559,N_2576);
and U2696 (N_2696,N_2584,N_2596);
nand U2697 (N_2697,N_2562,N_2613);
xnor U2698 (N_2698,N_2578,N_2616);
and U2699 (N_2699,N_2575,N_2594);
nand U2700 (N_2700,N_2650,N_2651);
nand U2701 (N_2701,N_2640,N_2688);
nand U2702 (N_2702,N_2625,N_2632);
nand U2703 (N_2703,N_2673,N_2665);
and U2704 (N_2704,N_2686,N_2695);
nand U2705 (N_2705,N_2644,N_2676);
nor U2706 (N_2706,N_2663,N_2694);
and U2707 (N_2707,N_2653,N_2637);
xor U2708 (N_2708,N_2677,N_2684);
nand U2709 (N_2709,N_2666,N_2698);
and U2710 (N_2710,N_2647,N_2639);
or U2711 (N_2711,N_2657,N_2661);
xnor U2712 (N_2712,N_2678,N_2654);
or U2713 (N_2713,N_2652,N_2696);
xnor U2714 (N_2714,N_2683,N_2628);
xor U2715 (N_2715,N_2691,N_2655);
or U2716 (N_2716,N_2646,N_2649);
xor U2717 (N_2717,N_2680,N_2697);
nor U2718 (N_2718,N_2660,N_2693);
or U2719 (N_2719,N_2645,N_2682);
or U2720 (N_2720,N_2689,N_2629);
xor U2721 (N_2721,N_2668,N_2634);
nand U2722 (N_2722,N_2692,N_2630);
xor U2723 (N_2723,N_2685,N_2658);
nand U2724 (N_2724,N_2669,N_2675);
nand U2725 (N_2725,N_2638,N_2681);
and U2726 (N_2726,N_2664,N_2659);
xnor U2727 (N_2727,N_2667,N_2648);
nand U2728 (N_2728,N_2662,N_2690);
nand U2729 (N_2729,N_2687,N_2679);
nand U2730 (N_2730,N_2642,N_2631);
xor U2731 (N_2731,N_2643,N_2656);
xnor U2732 (N_2732,N_2633,N_2672);
xor U2733 (N_2733,N_2636,N_2635);
xnor U2734 (N_2734,N_2641,N_2670);
nor U2735 (N_2735,N_2626,N_2699);
and U2736 (N_2736,N_2674,N_2671);
nand U2737 (N_2737,N_2627,N_2668);
nand U2738 (N_2738,N_2686,N_2644);
nand U2739 (N_2739,N_2687,N_2646);
or U2740 (N_2740,N_2642,N_2662);
and U2741 (N_2741,N_2647,N_2625);
or U2742 (N_2742,N_2627,N_2690);
or U2743 (N_2743,N_2626,N_2692);
nor U2744 (N_2744,N_2661,N_2687);
and U2745 (N_2745,N_2692,N_2640);
and U2746 (N_2746,N_2645,N_2636);
nor U2747 (N_2747,N_2644,N_2628);
xnor U2748 (N_2748,N_2648,N_2685);
xor U2749 (N_2749,N_2675,N_2699);
nor U2750 (N_2750,N_2660,N_2629);
nor U2751 (N_2751,N_2669,N_2645);
nand U2752 (N_2752,N_2685,N_2625);
nand U2753 (N_2753,N_2689,N_2670);
xnor U2754 (N_2754,N_2691,N_2678);
nand U2755 (N_2755,N_2686,N_2682);
and U2756 (N_2756,N_2678,N_2627);
xor U2757 (N_2757,N_2646,N_2661);
nor U2758 (N_2758,N_2654,N_2651);
nand U2759 (N_2759,N_2678,N_2689);
xor U2760 (N_2760,N_2698,N_2674);
or U2761 (N_2761,N_2664,N_2692);
nand U2762 (N_2762,N_2657,N_2630);
and U2763 (N_2763,N_2670,N_2643);
nor U2764 (N_2764,N_2682,N_2692);
and U2765 (N_2765,N_2691,N_2687);
nand U2766 (N_2766,N_2679,N_2668);
nand U2767 (N_2767,N_2693,N_2649);
and U2768 (N_2768,N_2629,N_2638);
nand U2769 (N_2769,N_2625,N_2667);
xor U2770 (N_2770,N_2646,N_2647);
or U2771 (N_2771,N_2678,N_2693);
xor U2772 (N_2772,N_2655,N_2633);
nand U2773 (N_2773,N_2666,N_2685);
and U2774 (N_2774,N_2672,N_2687);
and U2775 (N_2775,N_2725,N_2773);
nand U2776 (N_2776,N_2733,N_2744);
nand U2777 (N_2777,N_2738,N_2715);
nand U2778 (N_2778,N_2707,N_2705);
or U2779 (N_2779,N_2717,N_2768);
nand U2780 (N_2780,N_2748,N_2702);
and U2781 (N_2781,N_2752,N_2735);
nand U2782 (N_2782,N_2720,N_2710);
nor U2783 (N_2783,N_2741,N_2745);
nand U2784 (N_2784,N_2743,N_2724);
nor U2785 (N_2785,N_2711,N_2730);
or U2786 (N_2786,N_2746,N_2764);
xor U2787 (N_2787,N_2714,N_2771);
nand U2788 (N_2788,N_2753,N_2770);
and U2789 (N_2789,N_2713,N_2701);
xor U2790 (N_2790,N_2723,N_2736);
and U2791 (N_2791,N_2762,N_2765);
nor U2792 (N_2792,N_2718,N_2728);
nor U2793 (N_2793,N_2722,N_2704);
or U2794 (N_2794,N_2756,N_2740);
or U2795 (N_2795,N_2747,N_2755);
or U2796 (N_2796,N_2706,N_2766);
xor U2797 (N_2797,N_2731,N_2750);
nand U2798 (N_2798,N_2761,N_2760);
or U2799 (N_2799,N_2751,N_2742);
nand U2800 (N_2800,N_2769,N_2763);
or U2801 (N_2801,N_2716,N_2757);
xnor U2802 (N_2802,N_2726,N_2772);
xor U2803 (N_2803,N_2700,N_2737);
nand U2804 (N_2804,N_2754,N_2739);
nand U2805 (N_2805,N_2712,N_2721);
xnor U2806 (N_2806,N_2732,N_2749);
nand U2807 (N_2807,N_2708,N_2767);
nand U2808 (N_2808,N_2729,N_2774);
xnor U2809 (N_2809,N_2703,N_2719);
xnor U2810 (N_2810,N_2759,N_2709);
xnor U2811 (N_2811,N_2727,N_2758);
xor U2812 (N_2812,N_2734,N_2712);
or U2813 (N_2813,N_2703,N_2758);
and U2814 (N_2814,N_2737,N_2747);
nand U2815 (N_2815,N_2758,N_2728);
and U2816 (N_2816,N_2722,N_2768);
or U2817 (N_2817,N_2731,N_2764);
nand U2818 (N_2818,N_2708,N_2765);
or U2819 (N_2819,N_2739,N_2768);
xor U2820 (N_2820,N_2750,N_2727);
nor U2821 (N_2821,N_2774,N_2763);
and U2822 (N_2822,N_2743,N_2760);
and U2823 (N_2823,N_2732,N_2754);
and U2824 (N_2824,N_2765,N_2724);
xnor U2825 (N_2825,N_2725,N_2750);
and U2826 (N_2826,N_2755,N_2719);
xor U2827 (N_2827,N_2762,N_2753);
or U2828 (N_2828,N_2726,N_2725);
xor U2829 (N_2829,N_2705,N_2750);
nand U2830 (N_2830,N_2758,N_2755);
xnor U2831 (N_2831,N_2700,N_2770);
xnor U2832 (N_2832,N_2754,N_2773);
nor U2833 (N_2833,N_2755,N_2742);
nand U2834 (N_2834,N_2737,N_2733);
and U2835 (N_2835,N_2768,N_2754);
nor U2836 (N_2836,N_2751,N_2724);
or U2837 (N_2837,N_2759,N_2721);
nand U2838 (N_2838,N_2715,N_2751);
xnor U2839 (N_2839,N_2708,N_2772);
nand U2840 (N_2840,N_2767,N_2701);
xor U2841 (N_2841,N_2732,N_2743);
or U2842 (N_2842,N_2722,N_2751);
nor U2843 (N_2843,N_2724,N_2708);
nand U2844 (N_2844,N_2768,N_2710);
nand U2845 (N_2845,N_2707,N_2750);
nor U2846 (N_2846,N_2703,N_2744);
or U2847 (N_2847,N_2732,N_2724);
nand U2848 (N_2848,N_2706,N_2725);
and U2849 (N_2849,N_2743,N_2766);
nand U2850 (N_2850,N_2846,N_2819);
or U2851 (N_2851,N_2805,N_2784);
or U2852 (N_2852,N_2845,N_2849);
and U2853 (N_2853,N_2810,N_2787);
or U2854 (N_2854,N_2802,N_2780);
or U2855 (N_2855,N_2775,N_2794);
and U2856 (N_2856,N_2809,N_2823);
xor U2857 (N_2857,N_2778,N_2833);
and U2858 (N_2858,N_2788,N_2826);
and U2859 (N_2859,N_2801,N_2806);
nand U2860 (N_2860,N_2832,N_2785);
and U2861 (N_2861,N_2811,N_2821);
nor U2862 (N_2862,N_2796,N_2818);
xnor U2863 (N_2863,N_2779,N_2836);
nand U2864 (N_2864,N_2841,N_2807);
nor U2865 (N_2865,N_2830,N_2848);
nand U2866 (N_2866,N_2838,N_2790);
xnor U2867 (N_2867,N_2804,N_2812);
xor U2868 (N_2868,N_2827,N_2808);
nand U2869 (N_2869,N_2800,N_2803);
xor U2870 (N_2870,N_2783,N_2776);
xnor U2871 (N_2871,N_2840,N_2814);
and U2872 (N_2872,N_2777,N_2837);
xnor U2873 (N_2873,N_2834,N_2815);
or U2874 (N_2874,N_2799,N_2835);
or U2875 (N_2875,N_2797,N_2798);
and U2876 (N_2876,N_2817,N_2822);
and U2877 (N_2877,N_2789,N_2839);
or U2878 (N_2878,N_2842,N_2782);
and U2879 (N_2879,N_2831,N_2792);
and U2880 (N_2880,N_2843,N_2844);
and U2881 (N_2881,N_2813,N_2828);
xnor U2882 (N_2882,N_2825,N_2786);
or U2883 (N_2883,N_2793,N_2795);
nand U2884 (N_2884,N_2824,N_2829);
xor U2885 (N_2885,N_2816,N_2847);
or U2886 (N_2886,N_2781,N_2820);
and U2887 (N_2887,N_2791,N_2795);
nor U2888 (N_2888,N_2844,N_2795);
nand U2889 (N_2889,N_2835,N_2824);
and U2890 (N_2890,N_2776,N_2819);
xnor U2891 (N_2891,N_2823,N_2818);
nor U2892 (N_2892,N_2841,N_2791);
nand U2893 (N_2893,N_2840,N_2798);
nor U2894 (N_2894,N_2813,N_2848);
xor U2895 (N_2895,N_2821,N_2781);
nor U2896 (N_2896,N_2841,N_2816);
or U2897 (N_2897,N_2790,N_2846);
and U2898 (N_2898,N_2801,N_2815);
and U2899 (N_2899,N_2786,N_2781);
nor U2900 (N_2900,N_2796,N_2787);
nand U2901 (N_2901,N_2780,N_2790);
nand U2902 (N_2902,N_2839,N_2826);
and U2903 (N_2903,N_2818,N_2789);
or U2904 (N_2904,N_2847,N_2818);
nand U2905 (N_2905,N_2818,N_2825);
or U2906 (N_2906,N_2799,N_2790);
xnor U2907 (N_2907,N_2775,N_2813);
xor U2908 (N_2908,N_2826,N_2793);
nor U2909 (N_2909,N_2821,N_2834);
nor U2910 (N_2910,N_2834,N_2837);
and U2911 (N_2911,N_2780,N_2844);
nand U2912 (N_2912,N_2829,N_2795);
nand U2913 (N_2913,N_2833,N_2805);
and U2914 (N_2914,N_2789,N_2814);
and U2915 (N_2915,N_2797,N_2777);
or U2916 (N_2916,N_2785,N_2824);
xnor U2917 (N_2917,N_2799,N_2784);
and U2918 (N_2918,N_2793,N_2831);
or U2919 (N_2919,N_2797,N_2836);
or U2920 (N_2920,N_2823,N_2800);
or U2921 (N_2921,N_2839,N_2807);
nor U2922 (N_2922,N_2837,N_2830);
nand U2923 (N_2923,N_2790,N_2815);
and U2924 (N_2924,N_2805,N_2802);
or U2925 (N_2925,N_2871,N_2889);
nand U2926 (N_2926,N_2913,N_2898);
xnor U2927 (N_2927,N_2872,N_2893);
and U2928 (N_2928,N_2905,N_2902);
nor U2929 (N_2929,N_2903,N_2920);
and U2930 (N_2930,N_2882,N_2868);
and U2931 (N_2931,N_2896,N_2917);
nand U2932 (N_2932,N_2876,N_2918);
nand U2933 (N_2933,N_2892,N_2884);
and U2934 (N_2934,N_2873,N_2911);
xor U2935 (N_2935,N_2852,N_2904);
or U2936 (N_2936,N_2879,N_2885);
and U2937 (N_2937,N_2887,N_2863);
and U2938 (N_2938,N_2877,N_2921);
nor U2939 (N_2939,N_2907,N_2894);
nand U2940 (N_2940,N_2900,N_2857);
xnor U2941 (N_2941,N_2864,N_2909);
nand U2942 (N_2942,N_2858,N_2865);
and U2943 (N_2943,N_2880,N_2862);
xnor U2944 (N_2944,N_2881,N_2869);
xnor U2945 (N_2945,N_2851,N_2891);
nand U2946 (N_2946,N_2870,N_2850);
or U2947 (N_2947,N_2923,N_2883);
xnor U2948 (N_2948,N_2916,N_2924);
xor U2949 (N_2949,N_2908,N_2878);
nor U2950 (N_2950,N_2895,N_2859);
and U2951 (N_2951,N_2897,N_2853);
and U2952 (N_2952,N_2855,N_2899);
or U2953 (N_2953,N_2861,N_2919);
or U2954 (N_2954,N_2888,N_2875);
nand U2955 (N_2955,N_2901,N_2854);
nand U2956 (N_2956,N_2874,N_2886);
xnor U2957 (N_2957,N_2867,N_2856);
nor U2958 (N_2958,N_2860,N_2915);
nand U2959 (N_2959,N_2914,N_2922);
nand U2960 (N_2960,N_2912,N_2890);
or U2961 (N_2961,N_2866,N_2906);
and U2962 (N_2962,N_2910,N_2872);
nand U2963 (N_2963,N_2870,N_2851);
xnor U2964 (N_2964,N_2903,N_2918);
nor U2965 (N_2965,N_2862,N_2867);
xor U2966 (N_2966,N_2871,N_2872);
xor U2967 (N_2967,N_2911,N_2854);
nand U2968 (N_2968,N_2862,N_2883);
nor U2969 (N_2969,N_2880,N_2878);
nor U2970 (N_2970,N_2873,N_2918);
nor U2971 (N_2971,N_2902,N_2896);
and U2972 (N_2972,N_2916,N_2877);
nand U2973 (N_2973,N_2871,N_2875);
or U2974 (N_2974,N_2897,N_2888);
or U2975 (N_2975,N_2863,N_2878);
xor U2976 (N_2976,N_2894,N_2909);
xor U2977 (N_2977,N_2852,N_2900);
nor U2978 (N_2978,N_2920,N_2921);
nand U2979 (N_2979,N_2884,N_2888);
nand U2980 (N_2980,N_2886,N_2910);
or U2981 (N_2981,N_2895,N_2908);
nor U2982 (N_2982,N_2907,N_2922);
nand U2983 (N_2983,N_2869,N_2875);
nand U2984 (N_2984,N_2885,N_2855);
or U2985 (N_2985,N_2889,N_2902);
and U2986 (N_2986,N_2868,N_2880);
nor U2987 (N_2987,N_2918,N_2859);
or U2988 (N_2988,N_2874,N_2851);
nor U2989 (N_2989,N_2870,N_2895);
and U2990 (N_2990,N_2902,N_2872);
or U2991 (N_2991,N_2920,N_2872);
nor U2992 (N_2992,N_2860,N_2894);
and U2993 (N_2993,N_2895,N_2869);
nor U2994 (N_2994,N_2913,N_2875);
and U2995 (N_2995,N_2850,N_2902);
nand U2996 (N_2996,N_2875,N_2852);
and U2997 (N_2997,N_2911,N_2885);
nor U2998 (N_2998,N_2852,N_2898);
nor U2999 (N_2999,N_2921,N_2923);
or UO_0 (O_0,N_2935,N_2946);
nand UO_1 (O_1,N_2945,N_2975);
and UO_2 (O_2,N_2970,N_2966);
and UO_3 (O_3,N_2984,N_2978);
nor UO_4 (O_4,N_2983,N_2951);
nor UO_5 (O_5,N_2948,N_2931);
or UO_6 (O_6,N_2979,N_2961);
or UO_7 (O_7,N_2930,N_2958);
xnor UO_8 (O_8,N_2943,N_2953);
nand UO_9 (O_9,N_2938,N_2952);
nor UO_10 (O_10,N_2942,N_2980);
or UO_11 (O_11,N_2934,N_2986);
or UO_12 (O_12,N_2988,N_2995);
xor UO_13 (O_13,N_2976,N_2997);
xor UO_14 (O_14,N_2956,N_2973);
or UO_15 (O_15,N_2947,N_2964);
and UO_16 (O_16,N_2944,N_2972);
and UO_17 (O_17,N_2937,N_2941);
and UO_18 (O_18,N_2928,N_2940);
and UO_19 (O_19,N_2990,N_2949);
nand UO_20 (O_20,N_2999,N_2925);
nand UO_21 (O_21,N_2974,N_2982);
nor UO_22 (O_22,N_2959,N_2963);
xor UO_23 (O_23,N_2993,N_2977);
nor UO_24 (O_24,N_2929,N_2991);
nor UO_25 (O_25,N_2992,N_2955);
xor UO_26 (O_26,N_2981,N_2932);
xor UO_27 (O_27,N_2971,N_2998);
nand UO_28 (O_28,N_2985,N_2994);
or UO_29 (O_29,N_2965,N_2968);
xor UO_30 (O_30,N_2969,N_2967);
or UO_31 (O_31,N_2927,N_2954);
nand UO_32 (O_32,N_2939,N_2996);
nand UO_33 (O_33,N_2987,N_2960);
nand UO_34 (O_34,N_2989,N_2926);
xor UO_35 (O_35,N_2933,N_2936);
xnor UO_36 (O_36,N_2957,N_2962);
nand UO_37 (O_37,N_2950,N_2939);
nand UO_38 (O_38,N_2926,N_2946);
nand UO_39 (O_39,N_2998,N_2952);
nand UO_40 (O_40,N_2992,N_2968);
nand UO_41 (O_41,N_2993,N_2930);
and UO_42 (O_42,N_2981,N_2979);
nand UO_43 (O_43,N_2985,N_2986);
nand UO_44 (O_44,N_2964,N_2948);
or UO_45 (O_45,N_2965,N_2961);
xnor UO_46 (O_46,N_2961,N_2971);
nand UO_47 (O_47,N_2962,N_2966);
xnor UO_48 (O_48,N_2948,N_2943);
and UO_49 (O_49,N_2988,N_2987);
and UO_50 (O_50,N_2965,N_2953);
nand UO_51 (O_51,N_2972,N_2994);
xor UO_52 (O_52,N_2969,N_2975);
nor UO_53 (O_53,N_2997,N_2975);
nand UO_54 (O_54,N_2999,N_2968);
nor UO_55 (O_55,N_2967,N_2993);
nor UO_56 (O_56,N_2966,N_2960);
xor UO_57 (O_57,N_2974,N_2992);
and UO_58 (O_58,N_2934,N_2942);
and UO_59 (O_59,N_2947,N_2969);
nand UO_60 (O_60,N_2939,N_2978);
nand UO_61 (O_61,N_2959,N_2987);
or UO_62 (O_62,N_2985,N_2962);
or UO_63 (O_63,N_2929,N_2984);
nor UO_64 (O_64,N_2994,N_2955);
or UO_65 (O_65,N_2984,N_2925);
or UO_66 (O_66,N_2966,N_2994);
and UO_67 (O_67,N_2973,N_2936);
nand UO_68 (O_68,N_2956,N_2968);
xnor UO_69 (O_69,N_2925,N_2959);
nand UO_70 (O_70,N_2988,N_2976);
nor UO_71 (O_71,N_2927,N_2974);
or UO_72 (O_72,N_2925,N_2981);
nand UO_73 (O_73,N_2927,N_2930);
or UO_74 (O_74,N_2982,N_2987);
xor UO_75 (O_75,N_2960,N_2975);
nor UO_76 (O_76,N_2927,N_2968);
or UO_77 (O_77,N_2931,N_2989);
nor UO_78 (O_78,N_2936,N_2992);
nand UO_79 (O_79,N_2939,N_2963);
xnor UO_80 (O_80,N_2987,N_2995);
nor UO_81 (O_81,N_2962,N_2927);
xnor UO_82 (O_82,N_2972,N_2978);
or UO_83 (O_83,N_2989,N_2965);
xnor UO_84 (O_84,N_2956,N_2993);
xor UO_85 (O_85,N_2943,N_2977);
xnor UO_86 (O_86,N_2984,N_2998);
nor UO_87 (O_87,N_2952,N_2984);
nand UO_88 (O_88,N_2947,N_2937);
nand UO_89 (O_89,N_2941,N_2946);
xor UO_90 (O_90,N_2964,N_2966);
nand UO_91 (O_91,N_2945,N_2999);
and UO_92 (O_92,N_2986,N_2978);
or UO_93 (O_93,N_2991,N_2935);
and UO_94 (O_94,N_2945,N_2954);
or UO_95 (O_95,N_2941,N_2969);
nand UO_96 (O_96,N_2972,N_2965);
and UO_97 (O_97,N_2993,N_2952);
nor UO_98 (O_98,N_2985,N_2968);
nor UO_99 (O_99,N_2943,N_2954);
nor UO_100 (O_100,N_2977,N_2959);
and UO_101 (O_101,N_2952,N_2956);
and UO_102 (O_102,N_2957,N_2982);
xnor UO_103 (O_103,N_2986,N_2963);
or UO_104 (O_104,N_2952,N_2940);
and UO_105 (O_105,N_2941,N_2989);
or UO_106 (O_106,N_2991,N_2980);
and UO_107 (O_107,N_2987,N_2948);
xor UO_108 (O_108,N_2958,N_2937);
or UO_109 (O_109,N_2942,N_2927);
nor UO_110 (O_110,N_2935,N_2976);
or UO_111 (O_111,N_2996,N_2958);
nor UO_112 (O_112,N_2980,N_2938);
and UO_113 (O_113,N_2963,N_2992);
nand UO_114 (O_114,N_2938,N_2969);
xnor UO_115 (O_115,N_2926,N_2971);
xor UO_116 (O_116,N_2964,N_2967);
and UO_117 (O_117,N_2992,N_2998);
xor UO_118 (O_118,N_2949,N_2966);
nor UO_119 (O_119,N_2987,N_2980);
nor UO_120 (O_120,N_2972,N_2935);
or UO_121 (O_121,N_2997,N_2933);
nor UO_122 (O_122,N_2976,N_2947);
nor UO_123 (O_123,N_2930,N_2953);
nor UO_124 (O_124,N_2953,N_2942);
xnor UO_125 (O_125,N_2979,N_2990);
xnor UO_126 (O_126,N_2943,N_2959);
nor UO_127 (O_127,N_2944,N_2984);
and UO_128 (O_128,N_2960,N_2992);
xor UO_129 (O_129,N_2943,N_2974);
xnor UO_130 (O_130,N_2927,N_2987);
nor UO_131 (O_131,N_2934,N_2952);
or UO_132 (O_132,N_2943,N_2970);
and UO_133 (O_133,N_2971,N_2950);
xor UO_134 (O_134,N_2940,N_2966);
xnor UO_135 (O_135,N_2992,N_2929);
or UO_136 (O_136,N_2971,N_2937);
or UO_137 (O_137,N_2959,N_2973);
nor UO_138 (O_138,N_2926,N_2949);
and UO_139 (O_139,N_2998,N_2951);
xor UO_140 (O_140,N_2961,N_2995);
xnor UO_141 (O_141,N_2975,N_2988);
or UO_142 (O_142,N_2960,N_2933);
and UO_143 (O_143,N_2953,N_2985);
xor UO_144 (O_144,N_2979,N_2931);
nor UO_145 (O_145,N_2993,N_2982);
and UO_146 (O_146,N_2974,N_2949);
xnor UO_147 (O_147,N_2926,N_2953);
nor UO_148 (O_148,N_2973,N_2944);
nor UO_149 (O_149,N_2947,N_2990);
and UO_150 (O_150,N_2931,N_2978);
nor UO_151 (O_151,N_2999,N_2998);
xnor UO_152 (O_152,N_2960,N_2946);
xnor UO_153 (O_153,N_2934,N_2979);
nand UO_154 (O_154,N_2935,N_2954);
or UO_155 (O_155,N_2945,N_2965);
and UO_156 (O_156,N_2979,N_2939);
nand UO_157 (O_157,N_2938,N_2949);
nand UO_158 (O_158,N_2946,N_2956);
or UO_159 (O_159,N_2991,N_2939);
and UO_160 (O_160,N_2990,N_2952);
and UO_161 (O_161,N_2948,N_2951);
and UO_162 (O_162,N_2978,N_2983);
nor UO_163 (O_163,N_2928,N_2983);
and UO_164 (O_164,N_2928,N_2986);
nor UO_165 (O_165,N_2999,N_2952);
xor UO_166 (O_166,N_2986,N_2970);
nand UO_167 (O_167,N_2934,N_2949);
xnor UO_168 (O_168,N_2980,N_2926);
or UO_169 (O_169,N_2957,N_2994);
nand UO_170 (O_170,N_2993,N_2931);
nor UO_171 (O_171,N_2963,N_2969);
xor UO_172 (O_172,N_2995,N_2996);
or UO_173 (O_173,N_2949,N_2987);
nand UO_174 (O_174,N_2965,N_2970);
or UO_175 (O_175,N_2983,N_2946);
nor UO_176 (O_176,N_2978,N_2943);
and UO_177 (O_177,N_2944,N_2982);
nand UO_178 (O_178,N_2941,N_2931);
nor UO_179 (O_179,N_2977,N_2941);
nand UO_180 (O_180,N_2985,N_2929);
nor UO_181 (O_181,N_2984,N_2992);
xor UO_182 (O_182,N_2964,N_2944);
and UO_183 (O_183,N_2966,N_2972);
nand UO_184 (O_184,N_2971,N_2975);
nor UO_185 (O_185,N_2989,N_2955);
nor UO_186 (O_186,N_2994,N_2960);
or UO_187 (O_187,N_2973,N_2987);
or UO_188 (O_188,N_2992,N_2999);
and UO_189 (O_189,N_2961,N_2946);
nand UO_190 (O_190,N_2947,N_2939);
and UO_191 (O_191,N_2995,N_2964);
nor UO_192 (O_192,N_2991,N_2961);
or UO_193 (O_193,N_2960,N_2970);
and UO_194 (O_194,N_2956,N_2959);
and UO_195 (O_195,N_2998,N_2932);
and UO_196 (O_196,N_2928,N_2979);
and UO_197 (O_197,N_2993,N_2995);
and UO_198 (O_198,N_2980,N_2997);
nor UO_199 (O_199,N_2968,N_2991);
or UO_200 (O_200,N_2994,N_2940);
xnor UO_201 (O_201,N_2997,N_2977);
xnor UO_202 (O_202,N_2953,N_2938);
xor UO_203 (O_203,N_2926,N_2962);
nor UO_204 (O_204,N_2999,N_2966);
xnor UO_205 (O_205,N_2980,N_2941);
xnor UO_206 (O_206,N_2932,N_2955);
or UO_207 (O_207,N_2995,N_2981);
nand UO_208 (O_208,N_2998,N_2933);
nor UO_209 (O_209,N_2989,N_2937);
xor UO_210 (O_210,N_2950,N_2934);
nand UO_211 (O_211,N_2926,N_2977);
nand UO_212 (O_212,N_2993,N_2987);
nand UO_213 (O_213,N_2934,N_2963);
or UO_214 (O_214,N_2945,N_2982);
nor UO_215 (O_215,N_2997,N_2955);
xnor UO_216 (O_216,N_2971,N_2943);
nor UO_217 (O_217,N_2949,N_2935);
and UO_218 (O_218,N_2953,N_2950);
nand UO_219 (O_219,N_2937,N_2942);
nand UO_220 (O_220,N_2994,N_2984);
nor UO_221 (O_221,N_2937,N_2984);
nor UO_222 (O_222,N_2966,N_2986);
nor UO_223 (O_223,N_2954,N_2979);
nor UO_224 (O_224,N_2967,N_2974);
and UO_225 (O_225,N_2995,N_2992);
xor UO_226 (O_226,N_2979,N_2933);
nand UO_227 (O_227,N_2947,N_2933);
or UO_228 (O_228,N_2937,N_2959);
xor UO_229 (O_229,N_2950,N_2970);
or UO_230 (O_230,N_2959,N_2935);
xnor UO_231 (O_231,N_2942,N_2997);
xor UO_232 (O_232,N_2992,N_2970);
xnor UO_233 (O_233,N_2929,N_2977);
or UO_234 (O_234,N_2990,N_2944);
and UO_235 (O_235,N_2992,N_2961);
and UO_236 (O_236,N_2934,N_2976);
nand UO_237 (O_237,N_2926,N_2943);
nand UO_238 (O_238,N_2944,N_2952);
and UO_239 (O_239,N_2949,N_2953);
xor UO_240 (O_240,N_2949,N_2948);
nand UO_241 (O_241,N_2986,N_2932);
or UO_242 (O_242,N_2939,N_2935);
nand UO_243 (O_243,N_2937,N_2936);
xnor UO_244 (O_244,N_2941,N_2951);
and UO_245 (O_245,N_2988,N_2964);
and UO_246 (O_246,N_2944,N_2960);
or UO_247 (O_247,N_2958,N_2942);
or UO_248 (O_248,N_2970,N_2985);
nand UO_249 (O_249,N_2963,N_2948);
or UO_250 (O_250,N_2954,N_2967);
or UO_251 (O_251,N_2999,N_2988);
nor UO_252 (O_252,N_2960,N_2928);
nor UO_253 (O_253,N_2930,N_2961);
nor UO_254 (O_254,N_2991,N_2932);
xnor UO_255 (O_255,N_2974,N_2971);
nand UO_256 (O_256,N_2952,N_2973);
and UO_257 (O_257,N_2964,N_2997);
and UO_258 (O_258,N_2925,N_2958);
and UO_259 (O_259,N_2949,N_2970);
and UO_260 (O_260,N_2928,N_2969);
and UO_261 (O_261,N_2935,N_2993);
nor UO_262 (O_262,N_2951,N_2982);
and UO_263 (O_263,N_2949,N_2973);
xor UO_264 (O_264,N_2936,N_2955);
xor UO_265 (O_265,N_2960,N_2990);
nand UO_266 (O_266,N_2975,N_2944);
and UO_267 (O_267,N_2996,N_2992);
nor UO_268 (O_268,N_2963,N_2993);
nand UO_269 (O_269,N_2985,N_2999);
xnor UO_270 (O_270,N_2955,N_2940);
nor UO_271 (O_271,N_2937,N_2930);
xnor UO_272 (O_272,N_2994,N_2933);
nor UO_273 (O_273,N_2934,N_2941);
or UO_274 (O_274,N_2936,N_2940);
nor UO_275 (O_275,N_2943,N_2939);
or UO_276 (O_276,N_2966,N_2963);
nor UO_277 (O_277,N_2943,N_2980);
nor UO_278 (O_278,N_2932,N_2960);
and UO_279 (O_279,N_2958,N_2967);
or UO_280 (O_280,N_2988,N_2926);
nor UO_281 (O_281,N_2977,N_2994);
xnor UO_282 (O_282,N_2974,N_2929);
nand UO_283 (O_283,N_2989,N_2977);
nand UO_284 (O_284,N_2981,N_2933);
or UO_285 (O_285,N_2998,N_2953);
nand UO_286 (O_286,N_2969,N_2974);
xor UO_287 (O_287,N_2963,N_2999);
and UO_288 (O_288,N_2947,N_2936);
and UO_289 (O_289,N_2941,N_2972);
nor UO_290 (O_290,N_2938,N_2958);
nand UO_291 (O_291,N_2972,N_2993);
and UO_292 (O_292,N_2942,N_2983);
nor UO_293 (O_293,N_2964,N_2965);
and UO_294 (O_294,N_2932,N_2966);
or UO_295 (O_295,N_2987,N_2946);
nor UO_296 (O_296,N_2967,N_2930);
nand UO_297 (O_297,N_2944,N_2926);
nor UO_298 (O_298,N_2994,N_2989);
or UO_299 (O_299,N_2926,N_2940);
nand UO_300 (O_300,N_2947,N_2997);
or UO_301 (O_301,N_2972,N_2979);
or UO_302 (O_302,N_2989,N_2996);
xor UO_303 (O_303,N_2986,N_2939);
or UO_304 (O_304,N_2964,N_2940);
nor UO_305 (O_305,N_2981,N_2994);
nand UO_306 (O_306,N_2967,N_2957);
xnor UO_307 (O_307,N_2945,N_2967);
nand UO_308 (O_308,N_2993,N_2965);
xnor UO_309 (O_309,N_2985,N_2945);
nand UO_310 (O_310,N_2976,N_2953);
nand UO_311 (O_311,N_2966,N_2977);
nand UO_312 (O_312,N_2994,N_2982);
nor UO_313 (O_313,N_2965,N_2980);
or UO_314 (O_314,N_2948,N_2992);
and UO_315 (O_315,N_2935,N_2929);
xnor UO_316 (O_316,N_2975,N_2951);
or UO_317 (O_317,N_2986,N_2954);
nand UO_318 (O_318,N_2937,N_2998);
or UO_319 (O_319,N_2947,N_2961);
nand UO_320 (O_320,N_2936,N_2977);
nand UO_321 (O_321,N_2965,N_2955);
or UO_322 (O_322,N_2928,N_2965);
xor UO_323 (O_323,N_2977,N_2988);
xor UO_324 (O_324,N_2948,N_2927);
and UO_325 (O_325,N_2974,N_2937);
and UO_326 (O_326,N_2959,N_2995);
nor UO_327 (O_327,N_2974,N_2935);
and UO_328 (O_328,N_2973,N_2958);
xor UO_329 (O_329,N_2985,N_2983);
xor UO_330 (O_330,N_2947,N_2973);
or UO_331 (O_331,N_2933,N_2925);
and UO_332 (O_332,N_2944,N_2933);
or UO_333 (O_333,N_2947,N_2996);
nand UO_334 (O_334,N_2990,N_2926);
or UO_335 (O_335,N_2958,N_2932);
xnor UO_336 (O_336,N_2978,N_2962);
nand UO_337 (O_337,N_2928,N_2990);
or UO_338 (O_338,N_2957,N_2948);
xnor UO_339 (O_339,N_2981,N_2992);
or UO_340 (O_340,N_2955,N_2976);
and UO_341 (O_341,N_2987,N_2932);
xnor UO_342 (O_342,N_2947,N_2995);
nor UO_343 (O_343,N_2947,N_2987);
nor UO_344 (O_344,N_2943,N_2984);
xor UO_345 (O_345,N_2989,N_2968);
nand UO_346 (O_346,N_2960,N_2949);
or UO_347 (O_347,N_2929,N_2934);
nor UO_348 (O_348,N_2999,N_2986);
nor UO_349 (O_349,N_2953,N_2928);
nand UO_350 (O_350,N_2932,N_2965);
and UO_351 (O_351,N_2997,N_2931);
xor UO_352 (O_352,N_2964,N_2978);
or UO_353 (O_353,N_2943,N_2952);
or UO_354 (O_354,N_2989,N_2945);
or UO_355 (O_355,N_2961,N_2981);
nor UO_356 (O_356,N_2947,N_2970);
and UO_357 (O_357,N_2949,N_2993);
or UO_358 (O_358,N_2967,N_2935);
nor UO_359 (O_359,N_2974,N_2996);
or UO_360 (O_360,N_2930,N_2976);
nand UO_361 (O_361,N_2953,N_2983);
nor UO_362 (O_362,N_2942,N_2988);
and UO_363 (O_363,N_2974,N_2987);
and UO_364 (O_364,N_2982,N_2939);
nand UO_365 (O_365,N_2953,N_2931);
nor UO_366 (O_366,N_2937,N_2925);
xor UO_367 (O_367,N_2931,N_2992);
nor UO_368 (O_368,N_2990,N_2980);
nand UO_369 (O_369,N_2964,N_2938);
or UO_370 (O_370,N_2992,N_2967);
nor UO_371 (O_371,N_2986,N_2938);
or UO_372 (O_372,N_2979,N_2994);
nor UO_373 (O_373,N_2952,N_2988);
nand UO_374 (O_374,N_2982,N_2935);
xor UO_375 (O_375,N_2925,N_2977);
xor UO_376 (O_376,N_2947,N_2979);
nand UO_377 (O_377,N_2956,N_2992);
nand UO_378 (O_378,N_2953,N_2959);
nor UO_379 (O_379,N_2956,N_2943);
nor UO_380 (O_380,N_2957,N_2985);
or UO_381 (O_381,N_2945,N_2959);
and UO_382 (O_382,N_2988,N_2943);
nor UO_383 (O_383,N_2962,N_2931);
or UO_384 (O_384,N_2936,N_2953);
xor UO_385 (O_385,N_2970,N_2951);
and UO_386 (O_386,N_2969,N_2971);
or UO_387 (O_387,N_2959,N_2942);
or UO_388 (O_388,N_2944,N_2985);
nor UO_389 (O_389,N_2969,N_2987);
and UO_390 (O_390,N_2987,N_2933);
or UO_391 (O_391,N_2927,N_2957);
nor UO_392 (O_392,N_2945,N_2962);
nand UO_393 (O_393,N_2925,N_2975);
nand UO_394 (O_394,N_2951,N_2997);
nor UO_395 (O_395,N_2955,N_2966);
nand UO_396 (O_396,N_2970,N_2927);
and UO_397 (O_397,N_2983,N_2980);
and UO_398 (O_398,N_2954,N_2958);
nor UO_399 (O_399,N_2990,N_2932);
xor UO_400 (O_400,N_2955,N_2999);
nor UO_401 (O_401,N_2961,N_2975);
nand UO_402 (O_402,N_2932,N_2961);
nand UO_403 (O_403,N_2941,N_2982);
and UO_404 (O_404,N_2964,N_2955);
or UO_405 (O_405,N_2948,N_2973);
or UO_406 (O_406,N_2925,N_2965);
or UO_407 (O_407,N_2982,N_2969);
and UO_408 (O_408,N_2938,N_2934);
nand UO_409 (O_409,N_2986,N_2983);
nand UO_410 (O_410,N_2960,N_2930);
and UO_411 (O_411,N_2980,N_2949);
or UO_412 (O_412,N_2982,N_2928);
nand UO_413 (O_413,N_2937,N_2932);
nand UO_414 (O_414,N_2970,N_2993);
nand UO_415 (O_415,N_2940,N_2968);
nand UO_416 (O_416,N_2974,N_2991);
nand UO_417 (O_417,N_2926,N_2956);
or UO_418 (O_418,N_2995,N_2985);
nor UO_419 (O_419,N_2951,N_2925);
and UO_420 (O_420,N_2975,N_2979);
and UO_421 (O_421,N_2988,N_2968);
nor UO_422 (O_422,N_2978,N_2968);
xor UO_423 (O_423,N_2964,N_2960);
or UO_424 (O_424,N_2970,N_2989);
xor UO_425 (O_425,N_2975,N_2943);
xnor UO_426 (O_426,N_2949,N_2946);
or UO_427 (O_427,N_2953,N_2939);
and UO_428 (O_428,N_2951,N_2944);
nor UO_429 (O_429,N_2976,N_2994);
xnor UO_430 (O_430,N_2997,N_2998);
nor UO_431 (O_431,N_2939,N_2925);
nor UO_432 (O_432,N_2956,N_2961);
and UO_433 (O_433,N_2984,N_2993);
nor UO_434 (O_434,N_2933,N_2995);
and UO_435 (O_435,N_2947,N_2992);
nor UO_436 (O_436,N_2963,N_2989);
and UO_437 (O_437,N_2975,N_2987);
nand UO_438 (O_438,N_2972,N_2954);
or UO_439 (O_439,N_2930,N_2966);
nand UO_440 (O_440,N_2993,N_2966);
or UO_441 (O_441,N_2951,N_2969);
or UO_442 (O_442,N_2991,N_2949);
nor UO_443 (O_443,N_2951,N_2979);
nor UO_444 (O_444,N_2959,N_2951);
nand UO_445 (O_445,N_2960,N_2937);
xor UO_446 (O_446,N_2968,N_2941);
or UO_447 (O_447,N_2941,N_2950);
xnor UO_448 (O_448,N_2990,N_2955);
nand UO_449 (O_449,N_2930,N_2951);
and UO_450 (O_450,N_2997,N_2971);
and UO_451 (O_451,N_2927,N_2963);
or UO_452 (O_452,N_2951,N_2965);
xnor UO_453 (O_453,N_2969,N_2986);
or UO_454 (O_454,N_2964,N_2949);
nor UO_455 (O_455,N_2945,N_2963);
nor UO_456 (O_456,N_2962,N_2993);
nor UO_457 (O_457,N_2942,N_2932);
nand UO_458 (O_458,N_2973,N_2953);
nand UO_459 (O_459,N_2944,N_2945);
xnor UO_460 (O_460,N_2999,N_2975);
xor UO_461 (O_461,N_2990,N_2993);
and UO_462 (O_462,N_2961,N_2969);
xor UO_463 (O_463,N_2964,N_2961);
or UO_464 (O_464,N_2983,N_2934);
nor UO_465 (O_465,N_2942,N_2949);
xor UO_466 (O_466,N_2959,N_2991);
and UO_467 (O_467,N_2957,N_2944);
and UO_468 (O_468,N_2946,N_2968);
xnor UO_469 (O_469,N_2991,N_2942);
or UO_470 (O_470,N_2937,N_2934);
nor UO_471 (O_471,N_2937,N_2943);
or UO_472 (O_472,N_2928,N_2945);
or UO_473 (O_473,N_2941,N_2945);
xor UO_474 (O_474,N_2964,N_2958);
xor UO_475 (O_475,N_2951,N_2994);
or UO_476 (O_476,N_2991,N_2944);
nor UO_477 (O_477,N_2998,N_2964);
nor UO_478 (O_478,N_2970,N_2994);
and UO_479 (O_479,N_2950,N_2956);
and UO_480 (O_480,N_2973,N_2979);
xnor UO_481 (O_481,N_2960,N_2947);
nor UO_482 (O_482,N_2987,N_2964);
nand UO_483 (O_483,N_2992,N_2939);
xor UO_484 (O_484,N_2959,N_2992);
nor UO_485 (O_485,N_2958,N_2999);
nor UO_486 (O_486,N_2984,N_2973);
nor UO_487 (O_487,N_2994,N_2991);
nand UO_488 (O_488,N_2990,N_2968);
or UO_489 (O_489,N_2984,N_2956);
nand UO_490 (O_490,N_2969,N_2945);
or UO_491 (O_491,N_2967,N_2931);
xor UO_492 (O_492,N_2968,N_2938);
xor UO_493 (O_493,N_2945,N_2949);
and UO_494 (O_494,N_2960,N_2953);
and UO_495 (O_495,N_2948,N_2930);
and UO_496 (O_496,N_2982,N_2991);
or UO_497 (O_497,N_2940,N_2981);
and UO_498 (O_498,N_2971,N_2925);
nor UO_499 (O_499,N_2931,N_2944);
endmodule