module basic_1000_10000_1500_2_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5004,N_5005,N_5008,N_5009,N_5010,N_5011,N_5013,N_5015,N_5016,N_5018,N_5021,N_5022,N_5023,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5039,N_5041,N_5044,N_5045,N_5047,N_5049,N_5050,N_5051,N_5052,N_5056,N_5057,N_5058,N_5059,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5068,N_5071,N_5073,N_5074,N_5076,N_5079,N_5080,N_5081,N_5082,N_5084,N_5087,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5098,N_5099,N_5101,N_5103,N_5106,N_5111,N_5112,N_5114,N_5116,N_5118,N_5119,N_5122,N_5123,N_5127,N_5128,N_5129,N_5130,N_5131,N_5135,N_5136,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5151,N_5152,N_5153,N_5155,N_5156,N_5157,N_5159,N_5160,N_5162,N_5163,N_5164,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5177,N_5178,N_5179,N_5180,N_5182,N_5183,N_5186,N_5187,N_5190,N_5195,N_5196,N_5197,N_5199,N_5202,N_5203,N_5205,N_5206,N_5207,N_5208,N_5209,N_5211,N_5213,N_5214,N_5216,N_5218,N_5219,N_5221,N_5224,N_5225,N_5226,N_5227,N_5228,N_5230,N_5231,N_5232,N_5234,N_5236,N_5240,N_5243,N_5247,N_5248,N_5249,N_5252,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5271,N_5272,N_5273,N_5274,N_5278,N_5280,N_5281,N_5282,N_5285,N_5286,N_5288,N_5290,N_5292,N_5293,N_5294,N_5295,N_5296,N_5300,N_5302,N_5307,N_5308,N_5311,N_5313,N_5317,N_5319,N_5323,N_5326,N_5328,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5338,N_5339,N_5341,N_5342,N_5343,N_5345,N_5346,N_5347,N_5349,N_5352,N_5353,N_5354,N_5356,N_5357,N_5360,N_5361,N_5362,N_5363,N_5364,N_5367,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5376,N_5377,N_5378,N_5379,N_5382,N_5385,N_5386,N_5387,N_5388,N_5392,N_5393,N_5394,N_5395,N_5399,N_5400,N_5402,N_5404,N_5405,N_5406,N_5407,N_5408,N_5410,N_5411,N_5412,N_5414,N_5416,N_5417,N_5419,N_5420,N_5421,N_5422,N_5424,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5435,N_5437,N_5439,N_5440,N_5441,N_5442,N_5444,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5453,N_5454,N_5455,N_5458,N_5460,N_5462,N_5464,N_5466,N_5468,N_5469,N_5472,N_5473,N_5474,N_5475,N_5479,N_5480,N_5483,N_5484,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5500,N_5501,N_5503,N_5504,N_5505,N_5507,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5518,N_5521,N_5522,N_5524,N_5525,N_5526,N_5528,N_5529,N_5531,N_5532,N_5533,N_5534,N_5535,N_5538,N_5539,N_5541,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5553,N_5554,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5569,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5582,N_5583,N_5586,N_5588,N_5589,N_5590,N_5591,N_5592,N_5595,N_5596,N_5598,N_5600,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5610,N_5612,N_5615,N_5618,N_5620,N_5621,N_5622,N_5628,N_5630,N_5631,N_5636,N_5637,N_5639,N_5642,N_5644,N_5645,N_5648,N_5651,N_5652,N_5657,N_5658,N_5660,N_5662,N_5663,N_5664,N_5665,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5676,N_5679,N_5680,N_5682,N_5686,N_5687,N_5689,N_5690,N_5694,N_5697,N_5698,N_5699,N_5701,N_5702,N_5703,N_5705,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5735,N_5736,N_5738,N_5740,N_5741,N_5742,N_5743,N_5746,N_5747,N_5749,N_5751,N_5752,N_5753,N_5754,N_5756,N_5757,N_5759,N_5761,N_5762,N_5763,N_5764,N_5766,N_5767,N_5769,N_5770,N_5771,N_5774,N_5775,N_5776,N_5777,N_5779,N_5780,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5791,N_5793,N_5795,N_5796,N_5798,N_5802,N_5803,N_5807,N_5811,N_5812,N_5815,N_5818,N_5820,N_5823,N_5824,N_5825,N_5827,N_5828,N_5829,N_5831,N_5833,N_5835,N_5836,N_5837,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5848,N_5849,N_5851,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5863,N_5866,N_5867,N_5868,N_5869,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5882,N_5883,N_5884,N_5886,N_5887,N_5888,N_5890,N_5893,N_5896,N_5899,N_5900,N_5902,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5911,N_5914,N_5915,N_5917,N_5918,N_5921,N_5922,N_5923,N_5925,N_5927,N_5928,N_5930,N_5932,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5942,N_5945,N_5946,N_5947,N_5949,N_5951,N_5952,N_5954,N_5955,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5971,N_5973,N_5974,N_5976,N_5977,N_5980,N_5983,N_5984,N_5986,N_5989,N_5992,N_5994,N_5995,N_5996,N_5999,N_6000,N_6002,N_6003,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6012,N_6013,N_6014,N_6015,N_6018,N_6019,N_6021,N_6022,N_6023,N_6030,N_6031,N_6032,N_6034,N_6035,N_6036,N_6037,N_6042,N_6043,N_6045,N_6046,N_6048,N_6049,N_6050,N_6051,N_6053,N_6054,N_6056,N_6057,N_6058,N_6059,N_6061,N_6062,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6072,N_6073,N_6074,N_6075,N_6076,N_6080,N_6081,N_6082,N_6083,N_6087,N_6091,N_6094,N_6095,N_6096,N_6098,N_6100,N_6102,N_6104,N_6106,N_6107,N_6108,N_6110,N_6112,N_6114,N_6115,N_6117,N_6118,N_6119,N_6122,N_6123,N_6124,N_6125,N_6128,N_6129,N_6131,N_6132,N_6134,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6148,N_6150,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6162,N_6163,N_6164,N_6165,N_6170,N_6171,N_6172,N_6173,N_6174,N_6177,N_6178,N_6179,N_6180,N_6183,N_6184,N_6185,N_6186,N_6188,N_6189,N_6193,N_6195,N_6197,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6208,N_6209,N_6210,N_6211,N_6212,N_6214,N_6218,N_6219,N_6222,N_6223,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6238,N_6241,N_6242,N_6244,N_6245,N_6247,N_6253,N_6254,N_6255,N_6257,N_6258,N_6260,N_6261,N_6262,N_6264,N_6266,N_6267,N_6268,N_6270,N_6271,N_6272,N_6273,N_6274,N_6278,N_6282,N_6283,N_6284,N_6285,N_6286,N_6288,N_6289,N_6291,N_6292,N_6293,N_6294,N_6295,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6308,N_6310,N_6313,N_6315,N_6316,N_6318,N_6320,N_6321,N_6322,N_6323,N_6324,N_6326,N_6327,N_6330,N_6331,N_6333,N_6334,N_6336,N_6337,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6354,N_6357,N_6360,N_6361,N_6363,N_6366,N_6367,N_6368,N_6370,N_6371,N_6372,N_6373,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6382,N_6383,N_6385,N_6387,N_6389,N_6390,N_6393,N_6396,N_6400,N_6403,N_6405,N_6409,N_6410,N_6415,N_6416,N_6417,N_6421,N_6422,N_6423,N_6424,N_6428,N_6430,N_6431,N_6432,N_6433,N_6436,N_6437,N_6438,N_6440,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6449,N_6450,N_6452,N_6455,N_6457,N_6459,N_6460,N_6461,N_6464,N_6465,N_6466,N_6468,N_6472,N_6473,N_6477,N_6478,N_6480,N_6482,N_6483,N_6486,N_6487,N_6488,N_6489,N_6491,N_6492,N_6493,N_6494,N_6495,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6504,N_6505,N_6506,N_6509,N_6512,N_6514,N_6516,N_6518,N_6519,N_6520,N_6521,N_6522,N_6524,N_6525,N_6526,N_6528,N_6529,N_6530,N_6535,N_6537,N_6542,N_6543,N_6544,N_6545,N_6547,N_6549,N_6551,N_6552,N_6553,N_6554,N_6557,N_6558,N_6566,N_6567,N_6568,N_6569,N_6575,N_6576,N_6578,N_6579,N_6583,N_6584,N_6586,N_6587,N_6588,N_6591,N_6592,N_6593,N_6595,N_6596,N_6598,N_6599,N_6601,N_6602,N_6605,N_6606,N_6608,N_6609,N_6610,N_6611,N_6613,N_6615,N_6616,N_6619,N_6620,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6633,N_6635,N_6637,N_6639,N_6640,N_6641,N_6647,N_6648,N_6649,N_6651,N_6652,N_6653,N_6655,N_6656,N_6660,N_6662,N_6663,N_6665,N_6668,N_6670,N_6672,N_6674,N_6676,N_6678,N_6679,N_6681,N_6684,N_6685,N_6686,N_6688,N_6691,N_6692,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6703,N_6704,N_6709,N_6711,N_6713,N_6714,N_6715,N_6717,N_6718,N_6719,N_6720,N_6721,N_6724,N_6725,N_6727,N_6729,N_6730,N_6733,N_6734,N_6737,N_6740,N_6741,N_6745,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6755,N_6757,N_6758,N_6759,N_6762,N_6763,N_6764,N_6767,N_6770,N_6771,N_6772,N_6774,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6788,N_6791,N_6794,N_6796,N_6800,N_6803,N_6804,N_6805,N_6806,N_6808,N_6809,N_6810,N_6811,N_6812,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6821,N_6822,N_6823,N_6825,N_6827,N_6828,N_6829,N_6830,N_6833,N_6835,N_6837,N_6838,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6849,N_6850,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6866,N_6867,N_6868,N_6869,N_6870,N_6873,N_6876,N_6877,N_6879,N_6880,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6897,N_6898,N_6900,N_6901,N_6902,N_6903,N_6904,N_6907,N_6908,N_6910,N_6914,N_6915,N_6917,N_6918,N_6921,N_6923,N_6924,N_6925,N_6927,N_6928,N_6929,N_6930,N_6932,N_6934,N_6935,N_6939,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6950,N_6952,N_6954,N_6956,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6966,N_6967,N_6968,N_6969,N_6970,N_6973,N_6974,N_6975,N_6976,N_6978,N_6981,N_6982,N_6985,N_6989,N_6990,N_6991,N_6993,N_6994,N_6999,N_7000,N_7002,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7012,N_7015,N_7019,N_7021,N_7024,N_7025,N_7027,N_7030,N_7031,N_7033,N_7034,N_7035,N_7036,N_7037,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7049,N_7050,N_7051,N_7052,N_7054,N_7055,N_7057,N_7059,N_7061,N_7062,N_7064,N_7068,N_7069,N_7070,N_7072,N_7074,N_7075,N_7076,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7088,N_7091,N_7094,N_7097,N_7099,N_7100,N_7101,N_7103,N_7104,N_7110,N_7111,N_7112,N_7114,N_7115,N_7116,N_7117,N_7118,N_7120,N_7121,N_7122,N_7123,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7133,N_7134,N_7135,N_7136,N_7138,N_7139,N_7140,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7152,N_7153,N_7156,N_7157,N_7158,N_7160,N_7161,N_7163,N_7165,N_7166,N_7167,N_7168,N_7169,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7181,N_7182,N_7184,N_7190,N_7193,N_7196,N_7197,N_7198,N_7200,N_7202,N_7205,N_7206,N_7207,N_7211,N_7212,N_7214,N_7215,N_7218,N_7220,N_7221,N_7224,N_7225,N_7227,N_7230,N_7231,N_7233,N_7234,N_7236,N_7241,N_7243,N_7244,N_7246,N_7248,N_7249,N_7250,N_7251,N_7253,N_7254,N_7256,N_7257,N_7258,N_7262,N_7263,N_7267,N_7268,N_7269,N_7270,N_7271,N_7273,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7287,N_7288,N_7290,N_7291,N_7293,N_7294,N_7295,N_7296,N_7302,N_7303,N_7304,N_7305,N_7306,N_7309,N_7314,N_7315,N_7318,N_7320,N_7321,N_7326,N_7327,N_7328,N_7331,N_7333,N_7334,N_7336,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7348,N_7349,N_7350,N_7351,N_7352,N_7355,N_7358,N_7360,N_7361,N_7363,N_7365,N_7366,N_7367,N_7369,N_7373,N_7376,N_7377,N_7378,N_7382,N_7383,N_7385,N_7386,N_7387,N_7389,N_7390,N_7391,N_7394,N_7395,N_7396,N_7397,N_7399,N_7401,N_7402,N_7404,N_7405,N_7406,N_7409,N_7410,N_7413,N_7415,N_7419,N_7421,N_7423,N_7425,N_7426,N_7428,N_7430,N_7431,N_7432,N_7433,N_7435,N_7436,N_7438,N_7439,N_7440,N_7445,N_7446,N_7447,N_7448,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7464,N_7467,N_7470,N_7472,N_7473,N_7476,N_7478,N_7480,N_7481,N_7482,N_7483,N_7484,N_7486,N_7488,N_7490,N_7494,N_7498,N_7499,N_7500,N_7501,N_7503,N_7504,N_7505,N_7506,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7518,N_7519,N_7522,N_7523,N_7524,N_7525,N_7527,N_7528,N_7529,N_7530,N_7532,N_7534,N_7536,N_7541,N_7542,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7553,N_7554,N_7555,N_7556,N_7557,N_7559,N_7560,N_7562,N_7563,N_7565,N_7566,N_7567,N_7572,N_7573,N_7575,N_7576,N_7579,N_7581,N_7582,N_7584,N_7586,N_7588,N_7594,N_7596,N_7597,N_7598,N_7601,N_7603,N_7606,N_7608,N_7609,N_7611,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7627,N_7630,N_7633,N_7634,N_7637,N_7638,N_7639,N_7640,N_7643,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7654,N_7656,N_7658,N_7660,N_7663,N_7665,N_7666,N_7667,N_7668,N_7670,N_7671,N_7672,N_7675,N_7677,N_7680,N_7683,N_7684,N_7685,N_7688,N_7690,N_7694,N_7695,N_7696,N_7699,N_7702,N_7703,N_7704,N_7706,N_7707,N_7708,N_7709,N_7710,N_7712,N_7713,N_7714,N_7715,N_7716,N_7720,N_7721,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7733,N_7738,N_7740,N_7741,N_7744,N_7746,N_7747,N_7748,N_7750,N_7751,N_7752,N_7756,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7765,N_7768,N_7769,N_7770,N_7772,N_7775,N_7776,N_7779,N_7782,N_7785,N_7786,N_7788,N_7789,N_7790,N_7793,N_7794,N_7795,N_7798,N_7799,N_7800,N_7801,N_7803,N_7805,N_7807,N_7808,N_7809,N_7810,N_7811,N_7813,N_7814,N_7815,N_7816,N_7817,N_7819,N_7820,N_7821,N_7824,N_7825,N_7826,N_7827,N_7829,N_7830,N_7831,N_7832,N_7834,N_7835,N_7836,N_7838,N_7839,N_7840,N_7842,N_7845,N_7846,N_7847,N_7850,N_7852,N_7853,N_7854,N_7855,N_7857,N_7858,N_7859,N_7860,N_7861,N_7865,N_7866,N_7869,N_7870,N_7871,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7890,N_7891,N_7892,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7909,N_7910,N_7911,N_7912,N_7914,N_7915,N_7918,N_7919,N_7923,N_7927,N_7932,N_7935,N_7936,N_7938,N_7940,N_7942,N_7944,N_7945,N_7946,N_7948,N_7951,N_7952,N_7953,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7965,N_7966,N_7967,N_7971,N_7972,N_7973,N_7974,N_7975,N_7977,N_7978,N_7980,N_7982,N_7984,N_7985,N_7987,N_7988,N_7990,N_7992,N_7994,N_7995,N_8003,N_8006,N_8007,N_8009,N_8010,N_8012,N_8013,N_8016,N_8018,N_8022,N_8023,N_8024,N_8027,N_8028,N_8029,N_8030,N_8031,N_8033,N_8034,N_8035,N_8038,N_8039,N_8040,N_8043,N_8045,N_8046,N_8047,N_8048,N_8049,N_8051,N_8052,N_8055,N_8056,N_8057,N_8060,N_8062,N_8063,N_8066,N_8067,N_8072,N_8074,N_8076,N_8079,N_8086,N_8087,N_8088,N_8089,N_8091,N_8095,N_8096,N_8097,N_8098,N_8099,N_8102,N_8103,N_8104,N_8106,N_8107,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8120,N_8122,N_8123,N_8124,N_8126,N_8128,N_8130,N_8131,N_8133,N_8135,N_8136,N_8137,N_8138,N_8140,N_8142,N_8143,N_8144,N_8145,N_8146,N_8150,N_8152,N_8155,N_8156,N_8157,N_8159,N_8161,N_8162,N_8164,N_8165,N_8169,N_8172,N_8174,N_8175,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8189,N_8190,N_8192,N_8194,N_8195,N_8197,N_8200,N_8202,N_8203,N_8205,N_8210,N_8211,N_8212,N_8213,N_8214,N_8217,N_8220,N_8221,N_8222,N_8227,N_8228,N_8229,N_8232,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8242,N_8243,N_8244,N_8247,N_8248,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8261,N_8262,N_8263,N_8264,N_8266,N_8269,N_8274,N_8275,N_8276,N_8279,N_8280,N_8283,N_8286,N_8287,N_8288,N_8289,N_8291,N_8294,N_8295,N_8296,N_8297,N_8299,N_8300,N_8301,N_8303,N_8305,N_8306,N_8308,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8319,N_8320,N_8321,N_8323,N_8326,N_8328,N_8329,N_8330,N_8332,N_8333,N_8335,N_8338,N_8342,N_8343,N_8344,N_8345,N_8348,N_8349,N_8350,N_8356,N_8357,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8368,N_8369,N_8371,N_8373,N_8374,N_8376,N_8377,N_8380,N_8381,N_8384,N_8385,N_8386,N_8387,N_8389,N_8391,N_8393,N_8396,N_8398,N_8399,N_8400,N_8403,N_8405,N_8407,N_8408,N_8409,N_8410,N_8411,N_8416,N_8417,N_8418,N_8419,N_8421,N_8422,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8436,N_8439,N_8441,N_8442,N_8447,N_8449,N_8450,N_8451,N_8452,N_8455,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8466,N_8468,N_8469,N_8470,N_8471,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8490,N_8492,N_8493,N_8494,N_8495,N_8497,N_8498,N_8499,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8508,N_8509,N_8510,N_8512,N_8514,N_8516,N_8517,N_8518,N_8519,N_8520,N_8522,N_8523,N_8524,N_8525,N_8527,N_8529,N_8530,N_8531,N_8533,N_8535,N_8536,N_8537,N_8540,N_8543,N_8545,N_8547,N_8548,N_8553,N_8555,N_8557,N_8559,N_8560,N_8566,N_8568,N_8569,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8578,N_8580,N_8582,N_8583,N_8586,N_8587,N_8588,N_8589,N_8590,N_8592,N_8594,N_8595,N_8597,N_8600,N_8601,N_8602,N_8604,N_8606,N_8607,N_8609,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8619,N_8620,N_8625,N_8626,N_8627,N_8628,N_8629,N_8631,N_8632,N_8633,N_8636,N_8638,N_8639,N_8640,N_8641,N_8646,N_8647,N_8649,N_8651,N_8652,N_8653,N_8655,N_8656,N_8658,N_8659,N_8662,N_8663,N_8666,N_8667,N_8669,N_8671,N_8673,N_8675,N_8676,N_8677,N_8680,N_8681,N_8682,N_8684,N_8685,N_8686,N_8688,N_8690,N_8691,N_8692,N_8693,N_8698,N_8699,N_8700,N_8701,N_8703,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8714,N_8718,N_8719,N_8721,N_8722,N_8725,N_8726,N_8727,N_8728,N_8730,N_8731,N_8734,N_8735,N_8736,N_8737,N_8738,N_8741,N_8745,N_8747,N_8749,N_8752,N_8753,N_8755,N_8756,N_8758,N_8759,N_8761,N_8762,N_8764,N_8767,N_8768,N_8769,N_8772,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8789,N_8791,N_8793,N_8794,N_8795,N_8796,N_8798,N_8799,N_8802,N_8803,N_8806,N_8807,N_8808,N_8809,N_8810,N_8813,N_8814,N_8818,N_8821,N_8822,N_8824,N_8825,N_8826,N_8828,N_8829,N_8831,N_8832,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8854,N_8855,N_8857,N_8859,N_8861,N_8862,N_8864,N_8867,N_8869,N_8870,N_8871,N_8872,N_8874,N_8875,N_8876,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8886,N_8891,N_8892,N_8893,N_8895,N_8896,N_8897,N_8898,N_8900,N_8901,N_8902,N_8904,N_8906,N_8908,N_8909,N_8911,N_8912,N_8913,N_8915,N_8916,N_8917,N_8919,N_8921,N_8922,N_8925,N_8928,N_8929,N_8933,N_8934,N_8935,N_8937,N_8939,N_8943,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8953,N_8954,N_8955,N_8956,N_8958,N_8959,N_8960,N_8961,N_8962,N_8965,N_8967,N_8968,N_8969,N_8970,N_8971,N_8973,N_8974,N_8976,N_8977,N_8979,N_8980,N_8981,N_8982,N_8986,N_8987,N_8990,N_8992,N_8993,N_8996,N_8998,N_8999,N_9002,N_9004,N_9006,N_9009,N_9012,N_9014,N_9015,N_9017,N_9019,N_9020,N_9021,N_9022,N_9024,N_9025,N_9028,N_9032,N_9034,N_9037,N_9039,N_9043,N_9044,N_9045,N_9049,N_9050,N_9051,N_9056,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9069,N_9071,N_9072,N_9073,N_9074,N_9076,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9086,N_9087,N_9088,N_9089,N_9090,N_9094,N_9097,N_9098,N_9099,N_9103,N_9105,N_9106,N_9107,N_9108,N_9110,N_9111,N_9113,N_9114,N_9116,N_9125,N_9128,N_9129,N_9130,N_9134,N_9135,N_9136,N_9139,N_9141,N_9146,N_9147,N_9148,N_9149,N_9152,N_9153,N_9154,N_9155,N_9156,N_9159,N_9160,N_9163,N_9164,N_9165,N_9166,N_9168,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9185,N_9186,N_9192,N_9193,N_9194,N_9196,N_9197,N_9198,N_9200,N_9202,N_9203,N_9204,N_9206,N_9209,N_9212,N_9214,N_9215,N_9217,N_9218,N_9220,N_9221,N_9223,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9235,N_9237,N_9238,N_9241,N_9245,N_9246,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9259,N_9262,N_9264,N_9267,N_9270,N_9272,N_9273,N_9275,N_9276,N_9278,N_9279,N_9280,N_9282,N_9283,N_9286,N_9288,N_9290,N_9292,N_9294,N_9296,N_9301,N_9305,N_9306,N_9309,N_9311,N_9313,N_9314,N_9315,N_9316,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9328,N_9329,N_9330,N_9332,N_9333,N_9334,N_9335,N_9337,N_9338,N_9343,N_9344,N_9345,N_9352,N_9354,N_9356,N_9358,N_9359,N_9361,N_9362,N_9363,N_9365,N_9366,N_9367,N_9372,N_9373,N_9374,N_9376,N_9377,N_9378,N_9380,N_9381,N_9383,N_9385,N_9387,N_9389,N_9390,N_9391,N_9393,N_9397,N_9400,N_9401,N_9402,N_9403,N_9405,N_9406,N_9407,N_9408,N_9410,N_9411,N_9412,N_9413,N_9415,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9425,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9435,N_9437,N_9438,N_9441,N_9442,N_9444,N_9445,N_9446,N_9448,N_9449,N_9450,N_9454,N_9455,N_9457,N_9458,N_9461,N_9464,N_9466,N_9469,N_9471,N_9472,N_9473,N_9475,N_9478,N_9479,N_9481,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9493,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9507,N_9508,N_9510,N_9512,N_9513,N_9514,N_9516,N_9517,N_9518,N_9519,N_9521,N_9522,N_9523,N_9525,N_9527,N_9529,N_9530,N_9532,N_9533,N_9537,N_9538,N_9539,N_9540,N_9541,N_9544,N_9547,N_9548,N_9549,N_9551,N_9552,N_9557,N_9558,N_9560,N_9561,N_9566,N_9567,N_9568,N_9569,N_9570,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9581,N_9584,N_9585,N_9586,N_9587,N_9588,N_9590,N_9591,N_9592,N_9593,N_9594,N_9596,N_9597,N_9599,N_9600,N_9602,N_9603,N_9605,N_9612,N_9613,N_9616,N_9617,N_9618,N_9619,N_9620,N_9632,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9647,N_9648,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9661,N_9662,N_9664,N_9665,N_9667,N_9668,N_9672,N_9673,N_9675,N_9680,N_9682,N_9684,N_9685,N_9686,N_9687,N_9688,N_9690,N_9691,N_9692,N_9695,N_9696,N_9697,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9710,N_9712,N_9713,N_9714,N_9715,N_9716,N_9719,N_9720,N_9721,N_9722,N_9724,N_9727,N_9728,N_9729,N_9730,N_9731,N_9734,N_9737,N_9738,N_9739,N_9741,N_9743,N_9744,N_9745,N_9749,N_9750,N_9755,N_9756,N_9758,N_9760,N_9761,N_9762,N_9765,N_9766,N_9768,N_9769,N_9771,N_9772,N_9776,N_9777,N_9778,N_9780,N_9782,N_9784,N_9785,N_9786,N_9788,N_9789,N_9792,N_9797,N_9801,N_9802,N_9807,N_9808,N_9809,N_9810,N_9812,N_9813,N_9815,N_9816,N_9817,N_9819,N_9821,N_9825,N_9828,N_9830,N_9831,N_9832,N_9834,N_9836,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9845,N_9847,N_9848,N_9849,N_9850,N_9852,N_9854,N_9858,N_9859,N_9861,N_9863,N_9864,N_9865,N_9866,N_9867,N_9869,N_9871,N_9872,N_9874,N_9875,N_9876,N_9877,N_9880,N_9882,N_9886,N_9887,N_9888,N_9889,N_9894,N_9897,N_9898,N_9902,N_9903,N_9906,N_9907,N_9908,N_9909,N_9910,N_9912,N_9914,N_9915,N_9917,N_9921,N_9922,N_9923,N_9924,N_9925,N_9928,N_9933,N_9934,N_9935,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9944,N_9946,N_9948,N_9949,N_9951,N_9952,N_9954,N_9955,N_9956,N_9957,N_9959,N_9960,N_9961,N_9962,N_9963,N_9966,N_9967,N_9968,N_9970,N_9973,N_9976,N_9977,N_9978,N_9979,N_9983,N_9984,N_9986,N_9987,N_9990,N_9993,N_9996,N_9997,N_9999;
or U0 (N_0,In_43,In_664);
and U1 (N_1,In_22,In_706);
xnor U2 (N_2,In_169,In_646);
or U3 (N_3,In_80,In_615);
nor U4 (N_4,In_831,In_593);
nor U5 (N_5,In_60,In_724);
and U6 (N_6,In_946,In_901);
or U7 (N_7,In_549,In_960);
or U8 (N_8,In_819,In_32);
nor U9 (N_9,In_363,In_384);
xnor U10 (N_10,In_457,In_443);
nor U11 (N_11,In_364,In_353);
xnor U12 (N_12,In_699,In_514);
and U13 (N_13,In_663,In_25);
and U14 (N_14,In_841,In_975);
nor U15 (N_15,In_280,In_647);
nand U16 (N_16,In_405,In_648);
and U17 (N_17,In_4,In_544);
nor U18 (N_18,In_705,In_127);
or U19 (N_19,In_698,In_866);
or U20 (N_20,In_753,In_279);
nor U21 (N_21,In_190,In_522);
nor U22 (N_22,In_387,In_134);
nand U23 (N_23,In_145,In_553);
or U24 (N_24,In_128,In_587);
nand U25 (N_25,In_490,In_407);
nor U26 (N_26,In_47,In_650);
xor U27 (N_27,In_761,In_661);
xnor U28 (N_28,In_287,In_267);
and U29 (N_29,In_162,In_478);
nor U30 (N_30,In_362,In_390);
and U31 (N_31,In_981,In_868);
or U32 (N_32,In_36,In_210);
or U33 (N_33,In_18,In_933);
and U34 (N_34,In_50,In_247);
or U35 (N_35,In_30,In_800);
xor U36 (N_36,In_114,In_432);
nand U37 (N_37,In_158,In_397);
nor U38 (N_38,In_777,In_431);
nor U39 (N_39,In_968,In_602);
nand U40 (N_40,In_228,In_61);
xnor U41 (N_41,In_335,In_899);
and U42 (N_42,In_305,In_847);
xnor U43 (N_43,In_389,In_613);
or U44 (N_44,In_111,In_969);
or U45 (N_45,In_248,In_829);
and U46 (N_46,In_535,In_133);
and U47 (N_47,In_886,In_910);
nor U48 (N_48,In_294,In_143);
nor U49 (N_49,In_324,In_555);
nor U50 (N_50,In_726,In_898);
or U51 (N_51,In_500,In_160);
and U52 (N_52,In_897,In_23);
xnor U53 (N_53,In_953,In_419);
nand U54 (N_54,In_772,In_409);
or U55 (N_55,In_307,In_207);
or U56 (N_56,In_934,In_244);
xor U57 (N_57,In_468,In_386);
nand U58 (N_58,In_193,In_654);
and U59 (N_59,In_343,In_971);
xnor U60 (N_60,In_963,In_548);
and U61 (N_61,In_674,In_852);
xor U62 (N_62,In_673,In_356);
and U63 (N_63,In_635,In_872);
and U64 (N_64,In_941,In_271);
xnor U65 (N_65,In_843,In_687);
and U66 (N_66,In_856,In_179);
nand U67 (N_67,In_129,In_752);
nor U68 (N_68,In_321,In_561);
or U69 (N_69,In_985,In_166);
xor U70 (N_70,In_930,In_282);
nand U71 (N_71,In_967,In_449);
xnor U72 (N_72,In_49,In_911);
nor U73 (N_73,In_541,In_113);
and U74 (N_74,In_542,In_949);
or U75 (N_75,In_670,In_936);
and U76 (N_76,In_218,In_896);
and U77 (N_77,In_685,In_315);
or U78 (N_78,In_88,In_77);
nand U79 (N_79,In_436,In_251);
nand U80 (N_80,In_148,In_433);
and U81 (N_81,In_680,In_16);
nand U82 (N_82,In_543,In_918);
or U83 (N_83,In_684,In_204);
nand U84 (N_84,In_888,In_454);
and U85 (N_85,In_823,In_82);
and U86 (N_86,In_329,In_222);
or U87 (N_87,In_89,In_839);
and U88 (N_88,In_453,In_281);
xnor U89 (N_89,In_95,In_558);
nand U90 (N_90,In_511,In_887);
xnor U91 (N_91,In_580,In_26);
or U92 (N_92,In_869,In_229);
nor U93 (N_93,In_764,In_885);
or U94 (N_94,In_825,In_672);
xor U95 (N_95,In_678,In_711);
nor U96 (N_96,In_702,In_827);
and U97 (N_97,In_573,In_117);
or U98 (N_98,In_442,In_665);
nor U99 (N_99,In_970,In_340);
or U100 (N_100,In_197,In_607);
and U101 (N_101,In_520,In_72);
or U102 (N_102,In_401,In_631);
or U103 (N_103,In_574,In_632);
and U104 (N_104,In_810,In_504);
and U105 (N_105,In_8,In_494);
and U106 (N_106,In_171,In_37);
xnor U107 (N_107,In_177,In_225);
nor U108 (N_108,In_458,In_644);
nor U109 (N_109,In_299,In_150);
xor U110 (N_110,In_983,In_174);
xor U111 (N_111,In_217,In_475);
nand U112 (N_112,In_880,In_200);
and U113 (N_113,In_594,In_691);
xor U114 (N_114,In_917,In_756);
nand U115 (N_115,In_242,In_944);
xnor U116 (N_116,In_545,In_404);
xor U117 (N_117,In_750,In_400);
nand U118 (N_118,In_695,In_601);
xor U119 (N_119,In_516,In_130);
nand U120 (N_120,In_205,In_559);
nand U121 (N_121,In_184,In_283);
xnor U122 (N_122,In_894,In_451);
nor U123 (N_123,In_815,In_491);
and U124 (N_124,In_444,In_336);
xor U125 (N_125,In_368,In_378);
nand U126 (N_126,In_802,In_290);
nand U127 (N_127,In_54,In_477);
and U128 (N_128,In_260,In_849);
or U129 (N_129,In_583,In_199);
nand U130 (N_130,In_487,In_604);
or U131 (N_131,In_943,In_828);
nor U132 (N_132,In_308,In_392);
and U133 (N_133,In_306,In_838);
nand U134 (N_134,In_338,In_783);
nand U135 (N_135,In_572,In_793);
and U136 (N_136,In_135,In_620);
nand U137 (N_137,In_560,In_935);
or U138 (N_138,In_125,In_662);
nand U139 (N_139,In_703,In_618);
xor U140 (N_140,In_277,In_103);
xnor U141 (N_141,In_124,In_568);
and U142 (N_142,In_332,In_515);
xor U143 (N_143,In_743,In_424);
and U144 (N_144,In_211,In_126);
nand U145 (N_145,In_70,In_79);
xnor U146 (N_146,In_653,In_639);
and U147 (N_147,In_239,In_27);
and U148 (N_148,In_311,In_940);
xnor U149 (N_149,In_579,In_569);
or U150 (N_150,In_131,In_465);
and U151 (N_151,In_682,In_638);
nand U152 (N_152,In_221,In_909);
xnor U153 (N_153,In_339,In_472);
and U154 (N_154,In_67,In_649);
and U155 (N_155,In_224,In_581);
and U156 (N_156,In_12,In_105);
xor U157 (N_157,In_984,In_996);
nor U158 (N_158,In_817,In_964);
nor U159 (N_159,In_584,In_645);
nand U160 (N_160,In_448,In_293);
and U161 (N_161,In_13,In_881);
xor U162 (N_162,In_196,In_275);
nor U163 (N_163,In_634,In_320);
or U164 (N_164,In_0,In_657);
nor U165 (N_165,In_990,In_626);
and U166 (N_166,In_878,In_689);
nand U167 (N_167,In_519,In_907);
nand U168 (N_168,In_300,In_995);
xnor U169 (N_169,In_789,In_754);
and U170 (N_170,In_992,In_201);
or U171 (N_171,In_883,In_922);
nand U172 (N_172,In_534,In_877);
nor U173 (N_173,In_942,In_73);
or U174 (N_174,In_745,In_671);
and U175 (N_175,In_809,In_302);
nor U176 (N_176,In_844,In_816);
or U177 (N_177,In_213,In_342);
nand U178 (N_178,In_774,In_327);
nand U179 (N_179,In_156,In_110);
nand U180 (N_180,In_216,In_509);
nor U181 (N_181,In_873,In_485);
xor U182 (N_182,In_906,In_628);
nand U183 (N_183,In_15,In_86);
nand U184 (N_184,In_667,In_346);
nor U185 (N_185,In_379,In_413);
xnor U186 (N_186,In_483,In_735);
nand U187 (N_187,In_10,In_437);
nand U188 (N_188,In_845,In_312);
and U189 (N_189,In_425,In_314);
nand U190 (N_190,In_227,In_796);
or U191 (N_191,In_467,In_265);
or U192 (N_192,In_525,In_704);
and U193 (N_193,In_982,In_867);
nand U194 (N_194,In_694,In_729);
and U195 (N_195,In_417,In_440);
xor U196 (N_196,In_163,In_24);
or U197 (N_197,In_571,In_323);
or U198 (N_198,In_147,In_318);
xor U199 (N_199,In_220,In_484);
nand U200 (N_200,In_513,In_142);
nand U201 (N_201,In_68,In_997);
nand U202 (N_202,In_980,In_57);
xnor U203 (N_203,In_84,In_551);
nor U204 (N_204,In_479,In_482);
xor U205 (N_205,In_406,In_118);
nand U206 (N_206,In_837,In_2);
nor U207 (N_207,In_599,In_232);
or U208 (N_208,In_596,In_394);
and U209 (N_209,In_766,In_721);
xnor U210 (N_210,In_506,In_666);
and U211 (N_211,In_590,In_352);
xor U212 (N_212,In_798,In_209);
nor U213 (N_213,In_429,In_564);
nand U214 (N_214,In_427,In_759);
and U215 (N_215,In_144,In_245);
nand U216 (N_216,In_688,In_931);
nor U217 (N_217,In_42,In_556);
nand U218 (N_218,In_787,In_176);
nor U219 (N_219,In_832,In_263);
nand U220 (N_220,In_459,In_576);
nor U221 (N_221,In_316,In_999);
nand U222 (N_222,In_616,In_773);
nor U223 (N_223,In_187,In_624);
nor U224 (N_224,In_230,In_366);
or U225 (N_225,In_399,In_619);
xor U226 (N_226,In_755,In_799);
nand U227 (N_227,In_322,In_871);
and U228 (N_228,In_589,In_464);
nor U229 (N_229,In_234,In_769);
nor U230 (N_230,In_98,In_853);
nand U231 (N_231,In_334,In_902);
nor U232 (N_232,In_760,In_603);
xnor U233 (N_233,In_474,In_188);
or U234 (N_234,In_617,In_929);
and U235 (N_235,In_659,In_375);
nor U236 (N_236,In_337,In_198);
xor U237 (N_237,In_585,In_857);
nor U238 (N_238,In_780,In_391);
xnor U239 (N_239,In_497,In_412);
nor U240 (N_240,In_720,In_807);
nand U241 (N_241,In_591,In_182);
nand U242 (N_242,In_480,In_434);
nand U243 (N_243,In_505,In_836);
nor U244 (N_244,In_716,In_529);
and U245 (N_245,In_466,In_779);
nor U246 (N_246,In_998,In_805);
nand U247 (N_247,In_132,In_567);
or U248 (N_248,In_108,In_499);
and U249 (N_249,In_7,In_627);
nand U250 (N_250,In_701,In_508);
and U251 (N_251,In_882,In_722);
and U252 (N_252,In_994,In_859);
xnor U253 (N_253,In_233,In_446);
or U254 (N_254,In_369,In_903);
and U255 (N_255,In_778,In_347);
nor U256 (N_256,In_732,In_547);
xor U257 (N_257,In_101,In_889);
and U258 (N_258,In_139,In_582);
nor U259 (N_259,In_87,In_633);
nor U260 (N_260,In_532,In_530);
nand U261 (N_261,In_851,In_250);
and U262 (N_262,In_149,In_566);
and U263 (N_263,In_246,In_395);
nand U264 (N_264,In_81,In_396);
nor U265 (N_265,In_660,In_421);
nand U266 (N_266,In_115,In_501);
and U267 (N_267,In_261,In_492);
or U268 (N_268,In_104,In_846);
or U269 (N_269,In_374,In_119);
nor U270 (N_270,In_797,In_834);
or U271 (N_271,In_575,In_655);
or U272 (N_272,In_939,In_526);
xor U273 (N_273,In_266,In_58);
xor U274 (N_274,In_577,In_862);
or U275 (N_275,In_292,In_262);
nor U276 (N_276,In_916,In_758);
nor U277 (N_277,In_328,In_53);
xnor U278 (N_278,In_785,In_355);
or U279 (N_279,In_527,In_173);
xnor U280 (N_280,In_537,In_977);
and U281 (N_281,In_192,In_690);
nand U282 (N_282,In_636,In_238);
xnor U283 (N_283,In_813,In_164);
nor U284 (N_284,In_159,In_373);
nand U285 (N_285,In_710,In_937);
or U286 (N_286,In_154,In_622);
xnor U287 (N_287,In_393,In_681);
xnor U288 (N_288,In_383,In_202);
xnor U289 (N_289,In_713,In_989);
xnor U290 (N_290,In_712,In_489);
xor U291 (N_291,In_725,In_297);
nand U292 (N_292,In_170,In_826);
or U293 (N_293,In_563,In_254);
xor U294 (N_294,In_470,In_333);
nor U295 (N_295,In_462,In_959);
and U296 (N_296,In_71,In_600);
xor U297 (N_297,In_709,In_503);
nand U298 (N_298,In_614,In_641);
nand U299 (N_299,In_122,In_736);
and U300 (N_300,In_870,In_625);
xnor U301 (N_301,In_782,In_249);
or U302 (N_302,In_33,In_208);
xor U303 (N_303,In_276,In_748);
or U304 (N_304,In_658,In_137);
or U305 (N_305,In_675,In_765);
and U306 (N_306,In_606,In_153);
nor U307 (N_307,In_884,In_676);
nor U308 (N_308,In_498,In_730);
xor U309 (N_309,In_908,In_83);
nand U310 (N_310,In_295,In_966);
and U311 (N_311,In_97,In_264);
or U312 (N_312,In_788,In_415);
and U313 (N_313,In_31,In_441);
or U314 (N_314,In_140,In_330);
nand U315 (N_315,In_255,In_848);
or U316 (N_316,In_3,In_598);
or U317 (N_317,In_811,In_528);
nor U318 (N_318,In_69,In_28);
and U319 (N_319,In_411,In_874);
nand U320 (N_320,In_377,In_350);
nor U321 (N_321,In_957,In_426);
nor U322 (N_322,In_303,In_643);
nor U323 (N_323,In_398,In_90);
and U324 (N_324,In_152,In_29);
nand U325 (N_325,In_359,In_728);
and U326 (N_326,In_165,In_102);
xnor U327 (N_327,In_1,In_319);
xnor U328 (N_328,In_151,In_956);
or U329 (N_329,In_422,In_919);
xor U330 (N_330,In_733,In_741);
nand U331 (N_331,In_310,In_818);
nor U332 (N_332,In_240,In_178);
nor U333 (N_333,In_767,In_538);
and U334 (N_334,In_540,In_850);
xor U335 (N_335,In_21,In_189);
or U336 (N_336,In_469,In_679);
nand U337 (N_337,In_948,In_235);
nand U338 (N_338,In_637,In_418);
nand U339 (N_339,In_840,In_588);
xor U340 (N_340,In_253,In_175);
nor U341 (N_341,In_821,In_301);
and U342 (N_342,In_879,In_56);
xor U343 (N_343,In_35,In_146);
xor U344 (N_344,In_812,In_291);
xnor U345 (N_345,In_354,In_270);
nor U346 (N_346,In_219,In_241);
nand U347 (N_347,In_737,In_430);
xnor U348 (N_348,In_52,In_123);
and U349 (N_349,In_770,In_268);
xor U350 (N_350,In_740,In_928);
nor U351 (N_351,In_380,In_206);
nor U352 (N_352,In_172,In_447);
nor U353 (N_353,In_461,In_360);
or U354 (N_354,In_776,In_34);
xor U355 (N_355,In_286,In_993);
nor U356 (N_356,In_388,In_988);
nand U357 (N_357,In_900,In_860);
nor U358 (N_358,In_63,In_517);
or U359 (N_359,In_237,In_361);
xor U360 (N_360,In_259,In_801);
nor U361 (N_361,In_45,In_611);
nand U362 (N_362,In_257,In_858);
nor U363 (N_363,In_865,In_9);
or U364 (N_364,In_912,In_518);
and U365 (N_365,In_806,In_203);
xor U366 (N_366,In_592,In_371);
xor U367 (N_367,In_138,In_855);
or U368 (N_368,In_351,In_791);
or U369 (N_369,In_693,In_804);
nand U370 (N_370,In_236,In_44);
or U371 (N_371,In_357,In_195);
xnor U372 (N_372,In_313,In_326);
and U373 (N_373,In_920,In_742);
xnor U374 (N_374,In_803,In_775);
nor U375 (N_375,In_345,In_605);
nand U376 (N_376,In_652,In_925);
and U377 (N_377,In_183,In_367);
xor U378 (N_378,In_420,In_381);
nor U379 (N_379,In_94,In_621);
nand U380 (N_380,In_623,In_488);
nor U381 (N_381,In_309,In_784);
and U382 (N_382,In_141,In_521);
or U383 (N_383,In_550,In_414);
and U384 (N_384,In_794,In_93);
nand U385 (N_385,In_155,In_974);
xor U386 (N_386,In_385,In_372);
or U387 (N_387,In_820,In_973);
xor U388 (N_388,In_6,In_987);
and U389 (N_389,In_40,In_100);
nand U390 (N_390,In_830,In_452);
and U391 (N_391,In_692,In_757);
nand U392 (N_392,In_11,In_686);
nand U393 (N_393,In_486,In_445);
nor U394 (N_394,In_76,In_792);
and U395 (N_395,In_38,In_476);
xnor U396 (N_396,In_835,In_814);
xor U397 (N_397,In_473,In_284);
and U398 (N_398,In_921,In_121);
or U399 (N_399,In_289,In_924);
nor U400 (N_400,In_382,In_370);
or U401 (N_401,In_258,In_586);
or U402 (N_402,In_612,In_904);
or U403 (N_403,In_91,In_256);
nand U404 (N_404,In_744,In_822);
xnor U405 (N_405,In_546,In_428);
and U406 (N_406,In_578,In_194);
or U407 (N_407,In_214,In_640);
nor U408 (N_408,In_344,In_298);
xnor U409 (N_409,In_231,In_651);
or U410 (N_410,In_331,In_288);
xor U411 (N_411,In_629,In_471);
nand U412 (N_412,In_423,In_186);
and U413 (N_413,In_48,In_296);
xor U414 (N_414,In_875,In_668);
nand U415 (N_415,In_895,In_463);
or U416 (N_416,In_972,In_683);
and U417 (N_417,In_278,In_348);
and U418 (N_418,In_496,In_945);
xor U419 (N_419,In_439,In_642);
xor U420 (N_420,In_986,In_608);
and U421 (N_421,In_768,In_403);
and U422 (N_422,In_609,In_677);
or U423 (N_423,In_718,In_595);
xor U424 (N_424,In_630,In_926);
xor U425 (N_425,In_842,In_17);
xor U426 (N_426,In_99,In_274);
nor U427 (N_427,In_107,In_533);
xor U428 (N_428,In_191,In_978);
and U429 (N_429,In_876,In_531);
nand U430 (N_430,In_927,In_738);
and U431 (N_431,In_749,In_507);
nand U432 (N_432,In_106,In_954);
nand U433 (N_433,In_707,In_854);
xor U434 (N_434,In_700,In_961);
and U435 (N_435,In_243,In_955);
xor U436 (N_436,In_965,In_349);
nand U437 (N_437,In_304,In_763);
nor U438 (N_438,In_727,In_109);
nor U439 (N_439,In_435,In_915);
and U440 (N_440,In_958,In_65);
or U441 (N_441,In_923,In_656);
xor U442 (N_442,In_19,In_951);
nand U443 (N_443,In_493,In_116);
and U444 (N_444,In_512,In_891);
nand U445 (N_445,In_950,In_455);
nor U446 (N_446,In_747,In_358);
nor U447 (N_447,In_795,In_136);
xor U448 (N_448,In_46,In_952);
nor U449 (N_449,In_410,In_947);
nand U450 (N_450,In_762,In_481);
nand U451 (N_451,In_864,In_402);
or U452 (N_452,In_833,In_565);
nand U453 (N_453,In_78,In_719);
xor U454 (N_454,In_438,In_962);
xnor U455 (N_455,In_714,In_523);
or U456 (N_456,In_215,In_708);
nor U457 (N_457,In_450,In_610);
xnor U458 (N_458,In_552,In_252);
nand U459 (N_459,In_408,In_75);
or U460 (N_460,In_717,In_739);
xor U461 (N_461,In_786,In_991);
nor U462 (N_462,In_905,In_5);
nand U463 (N_463,In_696,In_64);
or U464 (N_464,In_539,In_562);
xnor U465 (N_465,In_59,In_85);
xor U466 (N_466,In_226,In_502);
nor U467 (N_467,In_39,In_14);
nand U468 (N_468,In_376,In_554);
or U469 (N_469,In_20,In_341);
or U470 (N_470,In_890,In_861);
xor U471 (N_471,In_272,In_892);
xor U472 (N_472,In_790,In_167);
nor U473 (N_473,In_913,In_92);
or U474 (N_474,In_524,In_161);
nand U475 (N_475,In_597,In_863);
nand U476 (N_476,In_74,In_66);
and U477 (N_477,In_697,In_62);
nand U478 (N_478,In_51,In_893);
or U479 (N_479,In_223,In_460);
and U480 (N_480,In_669,In_495);
nand U481 (N_481,In_570,In_55);
nor U482 (N_482,In_41,In_180);
xor U483 (N_483,In_96,In_771);
nor U484 (N_484,In_536,In_365);
or U485 (N_485,In_181,In_112);
or U486 (N_486,In_824,In_185);
nor U487 (N_487,In_976,In_120);
xor U488 (N_488,In_734,In_273);
nand U489 (N_489,In_751,In_269);
and U490 (N_490,In_979,In_746);
and U491 (N_491,In_317,In_781);
and U492 (N_492,In_212,In_168);
nand U493 (N_493,In_731,In_808);
or U494 (N_494,In_416,In_723);
or U495 (N_495,In_510,In_932);
and U496 (N_496,In_456,In_557);
and U497 (N_497,In_157,In_325);
nor U498 (N_498,In_715,In_938);
and U499 (N_499,In_914,In_285);
or U500 (N_500,In_120,In_89);
nand U501 (N_501,In_783,In_593);
xor U502 (N_502,In_97,In_652);
or U503 (N_503,In_339,In_457);
and U504 (N_504,In_879,In_967);
xor U505 (N_505,In_411,In_689);
nand U506 (N_506,In_543,In_803);
nor U507 (N_507,In_419,In_854);
or U508 (N_508,In_699,In_459);
xnor U509 (N_509,In_17,In_611);
xnor U510 (N_510,In_648,In_733);
nor U511 (N_511,In_16,In_167);
and U512 (N_512,In_922,In_340);
or U513 (N_513,In_839,In_251);
nand U514 (N_514,In_376,In_791);
and U515 (N_515,In_704,In_807);
or U516 (N_516,In_756,In_480);
and U517 (N_517,In_243,In_113);
nand U518 (N_518,In_468,In_876);
nand U519 (N_519,In_922,In_515);
nand U520 (N_520,In_562,In_851);
or U521 (N_521,In_208,In_753);
xor U522 (N_522,In_610,In_247);
or U523 (N_523,In_288,In_136);
nor U524 (N_524,In_358,In_886);
nor U525 (N_525,In_782,In_422);
nor U526 (N_526,In_712,In_454);
nor U527 (N_527,In_22,In_835);
xnor U528 (N_528,In_100,In_369);
xnor U529 (N_529,In_624,In_668);
and U530 (N_530,In_471,In_658);
nand U531 (N_531,In_526,In_42);
nor U532 (N_532,In_182,In_36);
or U533 (N_533,In_781,In_660);
nor U534 (N_534,In_567,In_18);
xnor U535 (N_535,In_974,In_116);
nand U536 (N_536,In_516,In_378);
and U537 (N_537,In_119,In_792);
or U538 (N_538,In_686,In_746);
and U539 (N_539,In_501,In_947);
or U540 (N_540,In_81,In_579);
xor U541 (N_541,In_476,In_264);
nor U542 (N_542,In_398,In_568);
xor U543 (N_543,In_614,In_777);
and U544 (N_544,In_771,In_750);
or U545 (N_545,In_184,In_507);
or U546 (N_546,In_532,In_322);
xor U547 (N_547,In_637,In_715);
and U548 (N_548,In_596,In_298);
nor U549 (N_549,In_197,In_349);
or U550 (N_550,In_49,In_177);
nand U551 (N_551,In_474,In_759);
nand U552 (N_552,In_447,In_620);
nand U553 (N_553,In_666,In_645);
nor U554 (N_554,In_179,In_869);
or U555 (N_555,In_888,In_733);
and U556 (N_556,In_224,In_670);
and U557 (N_557,In_933,In_546);
nand U558 (N_558,In_277,In_134);
or U559 (N_559,In_202,In_497);
nor U560 (N_560,In_786,In_313);
xnor U561 (N_561,In_851,In_646);
xnor U562 (N_562,In_554,In_361);
nand U563 (N_563,In_146,In_335);
or U564 (N_564,In_758,In_700);
xnor U565 (N_565,In_997,In_890);
xor U566 (N_566,In_166,In_241);
and U567 (N_567,In_359,In_339);
nand U568 (N_568,In_675,In_741);
xnor U569 (N_569,In_266,In_674);
or U570 (N_570,In_796,In_773);
nand U571 (N_571,In_827,In_538);
and U572 (N_572,In_880,In_762);
or U573 (N_573,In_530,In_837);
nand U574 (N_574,In_222,In_394);
and U575 (N_575,In_639,In_577);
nand U576 (N_576,In_800,In_585);
xor U577 (N_577,In_13,In_836);
xnor U578 (N_578,In_371,In_416);
nand U579 (N_579,In_853,In_908);
and U580 (N_580,In_339,In_686);
or U581 (N_581,In_503,In_419);
xor U582 (N_582,In_710,In_815);
xor U583 (N_583,In_854,In_254);
xnor U584 (N_584,In_307,In_511);
or U585 (N_585,In_161,In_589);
xor U586 (N_586,In_389,In_108);
and U587 (N_587,In_856,In_1);
and U588 (N_588,In_298,In_288);
xnor U589 (N_589,In_696,In_259);
and U590 (N_590,In_304,In_372);
and U591 (N_591,In_376,In_711);
or U592 (N_592,In_593,In_172);
nand U593 (N_593,In_701,In_17);
or U594 (N_594,In_504,In_176);
or U595 (N_595,In_554,In_241);
xnor U596 (N_596,In_893,In_888);
and U597 (N_597,In_884,In_286);
or U598 (N_598,In_91,In_908);
nor U599 (N_599,In_461,In_267);
and U600 (N_600,In_628,In_815);
or U601 (N_601,In_706,In_531);
nand U602 (N_602,In_104,In_557);
nand U603 (N_603,In_560,In_634);
nor U604 (N_604,In_565,In_416);
nand U605 (N_605,In_145,In_764);
or U606 (N_606,In_498,In_3);
and U607 (N_607,In_874,In_399);
nor U608 (N_608,In_451,In_159);
or U609 (N_609,In_268,In_982);
nor U610 (N_610,In_508,In_862);
nor U611 (N_611,In_629,In_689);
nor U612 (N_612,In_352,In_678);
nand U613 (N_613,In_667,In_748);
xor U614 (N_614,In_8,In_577);
nor U615 (N_615,In_264,In_123);
xor U616 (N_616,In_682,In_704);
nand U617 (N_617,In_806,In_896);
and U618 (N_618,In_803,In_293);
or U619 (N_619,In_38,In_128);
and U620 (N_620,In_796,In_951);
and U621 (N_621,In_665,In_554);
nand U622 (N_622,In_782,In_598);
or U623 (N_623,In_555,In_736);
nand U624 (N_624,In_891,In_196);
or U625 (N_625,In_696,In_300);
and U626 (N_626,In_982,In_256);
xnor U627 (N_627,In_557,In_713);
nor U628 (N_628,In_188,In_908);
nand U629 (N_629,In_736,In_83);
nand U630 (N_630,In_823,In_781);
or U631 (N_631,In_815,In_317);
and U632 (N_632,In_891,In_546);
or U633 (N_633,In_433,In_12);
or U634 (N_634,In_602,In_931);
and U635 (N_635,In_162,In_958);
nor U636 (N_636,In_444,In_142);
or U637 (N_637,In_138,In_62);
or U638 (N_638,In_573,In_197);
nor U639 (N_639,In_811,In_844);
and U640 (N_640,In_762,In_192);
and U641 (N_641,In_244,In_626);
nor U642 (N_642,In_537,In_231);
nor U643 (N_643,In_705,In_469);
nor U644 (N_644,In_21,In_560);
nand U645 (N_645,In_196,In_822);
nand U646 (N_646,In_785,In_380);
or U647 (N_647,In_167,In_915);
and U648 (N_648,In_739,In_894);
nor U649 (N_649,In_617,In_214);
or U650 (N_650,In_65,In_733);
nor U651 (N_651,In_380,In_123);
or U652 (N_652,In_564,In_784);
nor U653 (N_653,In_594,In_601);
and U654 (N_654,In_563,In_615);
xnor U655 (N_655,In_372,In_235);
xnor U656 (N_656,In_892,In_233);
or U657 (N_657,In_958,In_925);
xor U658 (N_658,In_442,In_277);
and U659 (N_659,In_868,In_164);
nand U660 (N_660,In_892,In_366);
nor U661 (N_661,In_92,In_38);
or U662 (N_662,In_619,In_731);
and U663 (N_663,In_836,In_88);
and U664 (N_664,In_201,In_29);
xor U665 (N_665,In_488,In_480);
and U666 (N_666,In_352,In_411);
nand U667 (N_667,In_871,In_237);
xor U668 (N_668,In_791,In_101);
nor U669 (N_669,In_252,In_675);
xnor U670 (N_670,In_156,In_206);
and U671 (N_671,In_345,In_470);
nor U672 (N_672,In_395,In_960);
xnor U673 (N_673,In_583,In_874);
and U674 (N_674,In_460,In_600);
xor U675 (N_675,In_59,In_459);
nor U676 (N_676,In_659,In_891);
nor U677 (N_677,In_265,In_375);
and U678 (N_678,In_738,In_261);
nand U679 (N_679,In_302,In_490);
nand U680 (N_680,In_273,In_358);
and U681 (N_681,In_857,In_628);
or U682 (N_682,In_509,In_287);
nand U683 (N_683,In_548,In_666);
or U684 (N_684,In_485,In_94);
and U685 (N_685,In_201,In_528);
xor U686 (N_686,In_879,In_951);
and U687 (N_687,In_373,In_926);
nand U688 (N_688,In_131,In_566);
xor U689 (N_689,In_185,In_506);
and U690 (N_690,In_498,In_890);
nand U691 (N_691,In_53,In_892);
xnor U692 (N_692,In_988,In_395);
xnor U693 (N_693,In_792,In_120);
or U694 (N_694,In_257,In_739);
xnor U695 (N_695,In_221,In_90);
and U696 (N_696,In_912,In_833);
or U697 (N_697,In_979,In_463);
and U698 (N_698,In_597,In_375);
or U699 (N_699,In_312,In_486);
nand U700 (N_700,In_716,In_513);
xnor U701 (N_701,In_139,In_387);
and U702 (N_702,In_497,In_186);
nor U703 (N_703,In_236,In_738);
and U704 (N_704,In_725,In_581);
or U705 (N_705,In_969,In_354);
nand U706 (N_706,In_106,In_263);
xor U707 (N_707,In_565,In_438);
nor U708 (N_708,In_499,In_495);
xnor U709 (N_709,In_0,In_937);
xnor U710 (N_710,In_50,In_990);
or U711 (N_711,In_485,In_30);
nand U712 (N_712,In_948,In_75);
nand U713 (N_713,In_455,In_379);
or U714 (N_714,In_36,In_26);
or U715 (N_715,In_564,In_333);
and U716 (N_716,In_278,In_3);
nand U717 (N_717,In_17,In_229);
nand U718 (N_718,In_216,In_406);
or U719 (N_719,In_290,In_604);
nand U720 (N_720,In_260,In_418);
and U721 (N_721,In_368,In_911);
xor U722 (N_722,In_331,In_971);
xor U723 (N_723,In_62,In_257);
xor U724 (N_724,In_17,In_440);
xnor U725 (N_725,In_125,In_613);
nor U726 (N_726,In_583,In_31);
and U727 (N_727,In_393,In_458);
xnor U728 (N_728,In_577,In_953);
xor U729 (N_729,In_531,In_84);
nand U730 (N_730,In_816,In_599);
or U731 (N_731,In_606,In_16);
or U732 (N_732,In_233,In_508);
or U733 (N_733,In_400,In_354);
xnor U734 (N_734,In_951,In_889);
xnor U735 (N_735,In_748,In_931);
or U736 (N_736,In_141,In_798);
nor U737 (N_737,In_353,In_108);
or U738 (N_738,In_240,In_312);
xnor U739 (N_739,In_592,In_506);
xor U740 (N_740,In_671,In_843);
and U741 (N_741,In_136,In_260);
nand U742 (N_742,In_966,In_370);
nand U743 (N_743,In_534,In_462);
nand U744 (N_744,In_118,In_211);
nand U745 (N_745,In_439,In_123);
or U746 (N_746,In_132,In_334);
nand U747 (N_747,In_636,In_865);
or U748 (N_748,In_383,In_755);
and U749 (N_749,In_245,In_899);
and U750 (N_750,In_565,In_525);
and U751 (N_751,In_242,In_614);
and U752 (N_752,In_588,In_12);
nand U753 (N_753,In_33,In_29);
xnor U754 (N_754,In_80,In_821);
or U755 (N_755,In_355,In_787);
nand U756 (N_756,In_468,In_968);
nand U757 (N_757,In_333,In_733);
and U758 (N_758,In_762,In_295);
nor U759 (N_759,In_841,In_567);
nand U760 (N_760,In_316,In_898);
and U761 (N_761,In_256,In_115);
nor U762 (N_762,In_100,In_606);
nor U763 (N_763,In_616,In_270);
nor U764 (N_764,In_215,In_345);
nor U765 (N_765,In_820,In_940);
or U766 (N_766,In_732,In_976);
nand U767 (N_767,In_956,In_407);
or U768 (N_768,In_14,In_271);
xor U769 (N_769,In_458,In_875);
or U770 (N_770,In_99,In_969);
and U771 (N_771,In_842,In_660);
or U772 (N_772,In_190,In_845);
or U773 (N_773,In_301,In_939);
xnor U774 (N_774,In_885,In_732);
and U775 (N_775,In_860,In_729);
nor U776 (N_776,In_801,In_254);
nor U777 (N_777,In_533,In_783);
xor U778 (N_778,In_512,In_457);
nor U779 (N_779,In_814,In_581);
nand U780 (N_780,In_298,In_442);
or U781 (N_781,In_319,In_743);
and U782 (N_782,In_102,In_339);
nand U783 (N_783,In_821,In_46);
xnor U784 (N_784,In_619,In_571);
and U785 (N_785,In_411,In_908);
and U786 (N_786,In_534,In_160);
or U787 (N_787,In_369,In_681);
or U788 (N_788,In_267,In_860);
xor U789 (N_789,In_712,In_797);
and U790 (N_790,In_240,In_21);
nand U791 (N_791,In_205,In_399);
and U792 (N_792,In_262,In_338);
xor U793 (N_793,In_872,In_9);
or U794 (N_794,In_282,In_425);
xnor U795 (N_795,In_140,In_985);
or U796 (N_796,In_269,In_957);
and U797 (N_797,In_844,In_732);
nor U798 (N_798,In_595,In_554);
nor U799 (N_799,In_312,In_483);
nand U800 (N_800,In_235,In_571);
or U801 (N_801,In_359,In_450);
nor U802 (N_802,In_582,In_769);
nand U803 (N_803,In_803,In_276);
nor U804 (N_804,In_508,In_829);
xnor U805 (N_805,In_1,In_816);
nand U806 (N_806,In_428,In_647);
and U807 (N_807,In_383,In_668);
or U808 (N_808,In_745,In_699);
and U809 (N_809,In_941,In_909);
nand U810 (N_810,In_949,In_34);
xor U811 (N_811,In_932,In_474);
and U812 (N_812,In_444,In_293);
nand U813 (N_813,In_222,In_304);
nand U814 (N_814,In_377,In_286);
or U815 (N_815,In_469,In_737);
or U816 (N_816,In_390,In_886);
nor U817 (N_817,In_152,In_934);
nand U818 (N_818,In_88,In_332);
nand U819 (N_819,In_588,In_905);
and U820 (N_820,In_509,In_779);
xnor U821 (N_821,In_38,In_489);
nand U822 (N_822,In_457,In_709);
nor U823 (N_823,In_538,In_410);
nand U824 (N_824,In_828,In_385);
or U825 (N_825,In_276,In_499);
or U826 (N_826,In_452,In_138);
nor U827 (N_827,In_215,In_206);
nor U828 (N_828,In_850,In_573);
xor U829 (N_829,In_348,In_936);
or U830 (N_830,In_532,In_152);
nor U831 (N_831,In_577,In_97);
and U832 (N_832,In_130,In_687);
and U833 (N_833,In_27,In_515);
and U834 (N_834,In_893,In_942);
or U835 (N_835,In_855,In_922);
or U836 (N_836,In_460,In_687);
or U837 (N_837,In_733,In_372);
nand U838 (N_838,In_795,In_277);
and U839 (N_839,In_523,In_991);
and U840 (N_840,In_616,In_126);
nor U841 (N_841,In_193,In_630);
or U842 (N_842,In_322,In_175);
nor U843 (N_843,In_908,In_864);
nand U844 (N_844,In_407,In_309);
or U845 (N_845,In_757,In_279);
xor U846 (N_846,In_686,In_621);
or U847 (N_847,In_204,In_683);
nand U848 (N_848,In_912,In_954);
nor U849 (N_849,In_284,In_750);
nand U850 (N_850,In_959,In_816);
nor U851 (N_851,In_277,In_460);
or U852 (N_852,In_305,In_736);
nor U853 (N_853,In_48,In_163);
nor U854 (N_854,In_646,In_570);
or U855 (N_855,In_723,In_498);
or U856 (N_856,In_313,In_693);
xnor U857 (N_857,In_872,In_788);
and U858 (N_858,In_228,In_969);
and U859 (N_859,In_484,In_335);
or U860 (N_860,In_834,In_92);
xor U861 (N_861,In_901,In_226);
nor U862 (N_862,In_37,In_428);
nand U863 (N_863,In_63,In_215);
xor U864 (N_864,In_604,In_389);
nand U865 (N_865,In_4,In_790);
nand U866 (N_866,In_951,In_512);
nand U867 (N_867,In_416,In_531);
and U868 (N_868,In_968,In_695);
and U869 (N_869,In_450,In_405);
xnor U870 (N_870,In_232,In_930);
nor U871 (N_871,In_383,In_429);
and U872 (N_872,In_593,In_237);
nand U873 (N_873,In_281,In_726);
nand U874 (N_874,In_412,In_598);
nand U875 (N_875,In_298,In_790);
nor U876 (N_876,In_438,In_288);
xnor U877 (N_877,In_428,In_470);
and U878 (N_878,In_989,In_64);
xnor U879 (N_879,In_271,In_109);
nor U880 (N_880,In_483,In_205);
or U881 (N_881,In_184,In_726);
xor U882 (N_882,In_303,In_18);
nand U883 (N_883,In_752,In_812);
or U884 (N_884,In_483,In_199);
nand U885 (N_885,In_892,In_852);
and U886 (N_886,In_988,In_208);
nor U887 (N_887,In_233,In_472);
nor U888 (N_888,In_972,In_728);
and U889 (N_889,In_106,In_252);
nand U890 (N_890,In_391,In_158);
and U891 (N_891,In_387,In_413);
nand U892 (N_892,In_288,In_320);
nor U893 (N_893,In_236,In_179);
or U894 (N_894,In_354,In_771);
nor U895 (N_895,In_186,In_716);
nand U896 (N_896,In_206,In_192);
nor U897 (N_897,In_513,In_970);
nor U898 (N_898,In_21,In_462);
or U899 (N_899,In_117,In_968);
xor U900 (N_900,In_463,In_834);
nor U901 (N_901,In_142,In_651);
xnor U902 (N_902,In_627,In_162);
nor U903 (N_903,In_461,In_749);
nor U904 (N_904,In_731,In_644);
nor U905 (N_905,In_235,In_812);
or U906 (N_906,In_472,In_974);
and U907 (N_907,In_178,In_13);
or U908 (N_908,In_246,In_363);
and U909 (N_909,In_988,In_811);
and U910 (N_910,In_742,In_873);
or U911 (N_911,In_640,In_961);
and U912 (N_912,In_897,In_711);
nor U913 (N_913,In_805,In_772);
nor U914 (N_914,In_312,In_930);
xnor U915 (N_915,In_804,In_624);
xor U916 (N_916,In_886,In_937);
xor U917 (N_917,In_772,In_95);
and U918 (N_918,In_884,In_745);
nand U919 (N_919,In_367,In_723);
nor U920 (N_920,In_285,In_37);
or U921 (N_921,In_543,In_940);
or U922 (N_922,In_777,In_874);
and U923 (N_923,In_472,In_220);
or U924 (N_924,In_517,In_104);
nand U925 (N_925,In_737,In_370);
xnor U926 (N_926,In_90,In_744);
nor U927 (N_927,In_880,In_772);
or U928 (N_928,In_340,In_520);
and U929 (N_929,In_444,In_800);
or U930 (N_930,In_142,In_232);
nor U931 (N_931,In_471,In_789);
nand U932 (N_932,In_344,In_160);
nor U933 (N_933,In_157,In_433);
and U934 (N_934,In_820,In_332);
nand U935 (N_935,In_607,In_822);
nor U936 (N_936,In_378,In_90);
or U937 (N_937,In_774,In_540);
or U938 (N_938,In_896,In_781);
nand U939 (N_939,In_86,In_474);
and U940 (N_940,In_731,In_435);
nor U941 (N_941,In_3,In_367);
xnor U942 (N_942,In_928,In_290);
or U943 (N_943,In_638,In_944);
or U944 (N_944,In_169,In_823);
nor U945 (N_945,In_951,In_443);
nor U946 (N_946,In_14,In_85);
xnor U947 (N_947,In_386,In_937);
xnor U948 (N_948,In_417,In_369);
nand U949 (N_949,In_69,In_17);
or U950 (N_950,In_756,In_783);
nand U951 (N_951,In_34,In_446);
nand U952 (N_952,In_6,In_844);
and U953 (N_953,In_365,In_799);
xnor U954 (N_954,In_705,In_997);
nor U955 (N_955,In_158,In_683);
nor U956 (N_956,In_707,In_628);
nand U957 (N_957,In_148,In_547);
xnor U958 (N_958,In_463,In_909);
or U959 (N_959,In_652,In_661);
and U960 (N_960,In_178,In_200);
and U961 (N_961,In_528,In_321);
nand U962 (N_962,In_130,In_907);
nor U963 (N_963,In_746,In_131);
xor U964 (N_964,In_513,In_219);
and U965 (N_965,In_595,In_808);
or U966 (N_966,In_239,In_887);
nand U967 (N_967,In_710,In_457);
nor U968 (N_968,In_378,In_831);
or U969 (N_969,In_842,In_436);
xor U970 (N_970,In_238,In_401);
xnor U971 (N_971,In_822,In_245);
or U972 (N_972,In_485,In_966);
or U973 (N_973,In_840,In_557);
and U974 (N_974,In_119,In_510);
nor U975 (N_975,In_576,In_503);
or U976 (N_976,In_161,In_444);
nand U977 (N_977,In_931,In_65);
nor U978 (N_978,In_236,In_933);
nor U979 (N_979,In_90,In_432);
nor U980 (N_980,In_482,In_127);
nand U981 (N_981,In_128,In_412);
nor U982 (N_982,In_627,In_532);
and U983 (N_983,In_237,In_76);
nand U984 (N_984,In_322,In_948);
xor U985 (N_985,In_871,In_506);
xor U986 (N_986,In_294,In_304);
xor U987 (N_987,In_305,In_721);
nand U988 (N_988,In_53,In_271);
nor U989 (N_989,In_182,In_295);
and U990 (N_990,In_177,In_136);
and U991 (N_991,In_511,In_841);
or U992 (N_992,In_710,In_128);
nor U993 (N_993,In_32,In_436);
nand U994 (N_994,In_490,In_358);
xor U995 (N_995,In_902,In_425);
xor U996 (N_996,In_906,In_119);
and U997 (N_997,In_946,In_383);
or U998 (N_998,In_779,In_432);
nand U999 (N_999,In_918,In_45);
nor U1000 (N_1000,In_995,In_902);
nand U1001 (N_1001,In_420,In_838);
or U1002 (N_1002,In_554,In_862);
nand U1003 (N_1003,In_472,In_31);
and U1004 (N_1004,In_31,In_58);
and U1005 (N_1005,In_417,In_210);
and U1006 (N_1006,In_141,In_538);
nand U1007 (N_1007,In_876,In_442);
or U1008 (N_1008,In_621,In_415);
nand U1009 (N_1009,In_903,In_147);
xnor U1010 (N_1010,In_814,In_239);
and U1011 (N_1011,In_522,In_254);
xnor U1012 (N_1012,In_264,In_278);
xor U1013 (N_1013,In_620,In_356);
or U1014 (N_1014,In_591,In_613);
nor U1015 (N_1015,In_175,In_138);
or U1016 (N_1016,In_764,In_655);
or U1017 (N_1017,In_283,In_215);
and U1018 (N_1018,In_73,In_654);
or U1019 (N_1019,In_986,In_446);
xor U1020 (N_1020,In_911,In_296);
nand U1021 (N_1021,In_160,In_362);
nor U1022 (N_1022,In_872,In_17);
and U1023 (N_1023,In_725,In_829);
nand U1024 (N_1024,In_317,In_719);
nor U1025 (N_1025,In_735,In_952);
nor U1026 (N_1026,In_993,In_295);
xnor U1027 (N_1027,In_271,In_309);
xnor U1028 (N_1028,In_571,In_26);
and U1029 (N_1029,In_249,In_976);
nor U1030 (N_1030,In_962,In_278);
nand U1031 (N_1031,In_859,In_781);
nand U1032 (N_1032,In_109,In_373);
nand U1033 (N_1033,In_765,In_225);
nor U1034 (N_1034,In_689,In_905);
nand U1035 (N_1035,In_275,In_764);
nand U1036 (N_1036,In_390,In_980);
nand U1037 (N_1037,In_0,In_811);
xnor U1038 (N_1038,In_379,In_605);
or U1039 (N_1039,In_920,In_957);
and U1040 (N_1040,In_530,In_865);
nor U1041 (N_1041,In_46,In_587);
nor U1042 (N_1042,In_198,In_813);
xor U1043 (N_1043,In_767,In_812);
xor U1044 (N_1044,In_61,In_753);
or U1045 (N_1045,In_601,In_470);
and U1046 (N_1046,In_511,In_891);
or U1047 (N_1047,In_626,In_482);
nor U1048 (N_1048,In_96,In_586);
nor U1049 (N_1049,In_777,In_787);
xnor U1050 (N_1050,In_307,In_767);
xor U1051 (N_1051,In_201,In_171);
nor U1052 (N_1052,In_948,In_442);
and U1053 (N_1053,In_541,In_672);
and U1054 (N_1054,In_862,In_799);
or U1055 (N_1055,In_126,In_454);
nor U1056 (N_1056,In_178,In_118);
nor U1057 (N_1057,In_520,In_395);
xor U1058 (N_1058,In_457,In_90);
nor U1059 (N_1059,In_926,In_440);
and U1060 (N_1060,In_602,In_711);
nand U1061 (N_1061,In_796,In_635);
nand U1062 (N_1062,In_16,In_880);
nand U1063 (N_1063,In_326,In_986);
or U1064 (N_1064,In_448,In_372);
nand U1065 (N_1065,In_126,In_357);
and U1066 (N_1066,In_452,In_117);
xor U1067 (N_1067,In_959,In_775);
or U1068 (N_1068,In_616,In_172);
nor U1069 (N_1069,In_518,In_939);
or U1070 (N_1070,In_796,In_856);
nor U1071 (N_1071,In_659,In_487);
and U1072 (N_1072,In_199,In_502);
or U1073 (N_1073,In_406,In_666);
xor U1074 (N_1074,In_230,In_933);
nand U1075 (N_1075,In_361,In_148);
xor U1076 (N_1076,In_999,In_591);
xor U1077 (N_1077,In_855,In_879);
nand U1078 (N_1078,In_313,In_529);
nor U1079 (N_1079,In_846,In_336);
and U1080 (N_1080,In_883,In_252);
and U1081 (N_1081,In_468,In_608);
and U1082 (N_1082,In_423,In_542);
xor U1083 (N_1083,In_590,In_158);
and U1084 (N_1084,In_216,In_920);
nor U1085 (N_1085,In_992,In_191);
nand U1086 (N_1086,In_33,In_96);
xor U1087 (N_1087,In_728,In_974);
nand U1088 (N_1088,In_739,In_335);
or U1089 (N_1089,In_744,In_557);
and U1090 (N_1090,In_89,In_680);
nor U1091 (N_1091,In_134,In_142);
xor U1092 (N_1092,In_956,In_589);
or U1093 (N_1093,In_584,In_761);
nor U1094 (N_1094,In_201,In_273);
nand U1095 (N_1095,In_582,In_735);
or U1096 (N_1096,In_388,In_914);
and U1097 (N_1097,In_961,In_888);
nor U1098 (N_1098,In_416,In_395);
nor U1099 (N_1099,In_851,In_813);
xnor U1100 (N_1100,In_944,In_558);
nand U1101 (N_1101,In_568,In_811);
nand U1102 (N_1102,In_904,In_605);
nand U1103 (N_1103,In_815,In_296);
nor U1104 (N_1104,In_525,In_646);
nor U1105 (N_1105,In_764,In_846);
and U1106 (N_1106,In_268,In_52);
nand U1107 (N_1107,In_541,In_936);
and U1108 (N_1108,In_559,In_500);
and U1109 (N_1109,In_639,In_138);
nor U1110 (N_1110,In_10,In_742);
or U1111 (N_1111,In_795,In_310);
nor U1112 (N_1112,In_214,In_972);
or U1113 (N_1113,In_849,In_881);
nor U1114 (N_1114,In_156,In_714);
nor U1115 (N_1115,In_569,In_800);
xnor U1116 (N_1116,In_286,In_706);
nand U1117 (N_1117,In_349,In_884);
xor U1118 (N_1118,In_124,In_797);
xnor U1119 (N_1119,In_551,In_80);
or U1120 (N_1120,In_145,In_430);
xnor U1121 (N_1121,In_309,In_153);
or U1122 (N_1122,In_166,In_28);
nand U1123 (N_1123,In_700,In_467);
nand U1124 (N_1124,In_229,In_187);
or U1125 (N_1125,In_14,In_410);
nor U1126 (N_1126,In_555,In_363);
nand U1127 (N_1127,In_374,In_244);
and U1128 (N_1128,In_182,In_366);
nor U1129 (N_1129,In_93,In_317);
xnor U1130 (N_1130,In_900,In_525);
and U1131 (N_1131,In_495,In_60);
and U1132 (N_1132,In_136,In_80);
and U1133 (N_1133,In_744,In_901);
xor U1134 (N_1134,In_166,In_873);
and U1135 (N_1135,In_261,In_153);
or U1136 (N_1136,In_633,In_524);
nand U1137 (N_1137,In_380,In_884);
or U1138 (N_1138,In_196,In_112);
and U1139 (N_1139,In_630,In_262);
nor U1140 (N_1140,In_168,In_31);
or U1141 (N_1141,In_489,In_171);
and U1142 (N_1142,In_582,In_334);
nor U1143 (N_1143,In_602,In_670);
nor U1144 (N_1144,In_194,In_50);
and U1145 (N_1145,In_988,In_43);
nand U1146 (N_1146,In_604,In_913);
and U1147 (N_1147,In_92,In_0);
nand U1148 (N_1148,In_772,In_333);
or U1149 (N_1149,In_783,In_39);
nand U1150 (N_1150,In_501,In_712);
nand U1151 (N_1151,In_571,In_726);
nand U1152 (N_1152,In_352,In_203);
xnor U1153 (N_1153,In_663,In_195);
and U1154 (N_1154,In_174,In_867);
nand U1155 (N_1155,In_123,In_581);
nand U1156 (N_1156,In_753,In_378);
nand U1157 (N_1157,In_325,In_482);
and U1158 (N_1158,In_114,In_382);
nand U1159 (N_1159,In_87,In_809);
nand U1160 (N_1160,In_704,In_868);
and U1161 (N_1161,In_499,In_120);
xnor U1162 (N_1162,In_22,In_578);
xnor U1163 (N_1163,In_761,In_305);
xor U1164 (N_1164,In_263,In_105);
nor U1165 (N_1165,In_663,In_509);
nor U1166 (N_1166,In_11,In_319);
and U1167 (N_1167,In_507,In_295);
nor U1168 (N_1168,In_710,In_405);
and U1169 (N_1169,In_350,In_833);
nand U1170 (N_1170,In_242,In_949);
xnor U1171 (N_1171,In_442,In_953);
nand U1172 (N_1172,In_378,In_871);
nand U1173 (N_1173,In_28,In_93);
or U1174 (N_1174,In_429,In_268);
xnor U1175 (N_1175,In_120,In_21);
nor U1176 (N_1176,In_561,In_77);
nand U1177 (N_1177,In_499,In_861);
xnor U1178 (N_1178,In_149,In_153);
nand U1179 (N_1179,In_256,In_751);
or U1180 (N_1180,In_838,In_621);
or U1181 (N_1181,In_818,In_157);
nand U1182 (N_1182,In_618,In_795);
or U1183 (N_1183,In_299,In_274);
nand U1184 (N_1184,In_571,In_956);
or U1185 (N_1185,In_142,In_328);
nor U1186 (N_1186,In_759,In_718);
xnor U1187 (N_1187,In_928,In_988);
xor U1188 (N_1188,In_414,In_537);
xnor U1189 (N_1189,In_740,In_862);
and U1190 (N_1190,In_971,In_370);
nand U1191 (N_1191,In_722,In_229);
nor U1192 (N_1192,In_208,In_4);
or U1193 (N_1193,In_649,In_102);
xor U1194 (N_1194,In_567,In_65);
and U1195 (N_1195,In_520,In_69);
nor U1196 (N_1196,In_551,In_274);
nand U1197 (N_1197,In_729,In_345);
and U1198 (N_1198,In_6,In_90);
and U1199 (N_1199,In_131,In_385);
and U1200 (N_1200,In_66,In_661);
or U1201 (N_1201,In_721,In_450);
and U1202 (N_1202,In_659,In_220);
or U1203 (N_1203,In_691,In_251);
xnor U1204 (N_1204,In_600,In_345);
nand U1205 (N_1205,In_160,In_291);
nand U1206 (N_1206,In_867,In_951);
nand U1207 (N_1207,In_281,In_231);
nor U1208 (N_1208,In_808,In_136);
or U1209 (N_1209,In_493,In_590);
nor U1210 (N_1210,In_114,In_845);
nand U1211 (N_1211,In_176,In_229);
nand U1212 (N_1212,In_862,In_769);
and U1213 (N_1213,In_128,In_435);
xnor U1214 (N_1214,In_683,In_141);
nand U1215 (N_1215,In_84,In_741);
xor U1216 (N_1216,In_434,In_6);
nor U1217 (N_1217,In_293,In_738);
xnor U1218 (N_1218,In_750,In_753);
nand U1219 (N_1219,In_30,In_610);
nor U1220 (N_1220,In_64,In_89);
and U1221 (N_1221,In_883,In_632);
nand U1222 (N_1222,In_348,In_532);
xor U1223 (N_1223,In_38,In_632);
xnor U1224 (N_1224,In_946,In_900);
nand U1225 (N_1225,In_655,In_110);
nand U1226 (N_1226,In_247,In_757);
and U1227 (N_1227,In_698,In_281);
or U1228 (N_1228,In_517,In_667);
and U1229 (N_1229,In_293,In_274);
or U1230 (N_1230,In_568,In_809);
or U1231 (N_1231,In_17,In_850);
or U1232 (N_1232,In_475,In_430);
nand U1233 (N_1233,In_676,In_947);
and U1234 (N_1234,In_873,In_43);
nor U1235 (N_1235,In_633,In_400);
nor U1236 (N_1236,In_904,In_912);
and U1237 (N_1237,In_91,In_161);
and U1238 (N_1238,In_895,In_478);
or U1239 (N_1239,In_553,In_671);
and U1240 (N_1240,In_675,In_72);
and U1241 (N_1241,In_416,In_849);
and U1242 (N_1242,In_884,In_849);
nor U1243 (N_1243,In_522,In_966);
nand U1244 (N_1244,In_614,In_933);
xor U1245 (N_1245,In_408,In_314);
nand U1246 (N_1246,In_796,In_611);
nand U1247 (N_1247,In_690,In_654);
nand U1248 (N_1248,In_17,In_655);
nor U1249 (N_1249,In_249,In_832);
or U1250 (N_1250,In_339,In_891);
or U1251 (N_1251,In_766,In_331);
nor U1252 (N_1252,In_908,In_963);
nand U1253 (N_1253,In_839,In_97);
nand U1254 (N_1254,In_604,In_418);
nor U1255 (N_1255,In_550,In_675);
and U1256 (N_1256,In_254,In_829);
and U1257 (N_1257,In_586,In_414);
or U1258 (N_1258,In_196,In_739);
nand U1259 (N_1259,In_867,In_264);
nand U1260 (N_1260,In_891,In_848);
xnor U1261 (N_1261,In_427,In_223);
xor U1262 (N_1262,In_266,In_421);
nor U1263 (N_1263,In_345,In_929);
nand U1264 (N_1264,In_562,In_358);
xor U1265 (N_1265,In_435,In_885);
xor U1266 (N_1266,In_623,In_274);
xor U1267 (N_1267,In_309,In_852);
or U1268 (N_1268,In_17,In_686);
xor U1269 (N_1269,In_880,In_279);
nor U1270 (N_1270,In_696,In_433);
xor U1271 (N_1271,In_832,In_957);
nand U1272 (N_1272,In_232,In_519);
and U1273 (N_1273,In_640,In_684);
and U1274 (N_1274,In_69,In_490);
nand U1275 (N_1275,In_2,In_591);
and U1276 (N_1276,In_526,In_935);
or U1277 (N_1277,In_407,In_387);
and U1278 (N_1278,In_980,In_159);
nand U1279 (N_1279,In_196,In_497);
nand U1280 (N_1280,In_76,In_171);
nor U1281 (N_1281,In_540,In_969);
and U1282 (N_1282,In_208,In_413);
and U1283 (N_1283,In_389,In_901);
and U1284 (N_1284,In_389,In_793);
or U1285 (N_1285,In_279,In_829);
or U1286 (N_1286,In_637,In_57);
nor U1287 (N_1287,In_622,In_823);
or U1288 (N_1288,In_129,In_52);
and U1289 (N_1289,In_432,In_577);
nand U1290 (N_1290,In_501,In_281);
or U1291 (N_1291,In_669,In_654);
nor U1292 (N_1292,In_510,In_946);
xor U1293 (N_1293,In_210,In_565);
nand U1294 (N_1294,In_914,In_425);
nor U1295 (N_1295,In_719,In_918);
and U1296 (N_1296,In_894,In_353);
xnor U1297 (N_1297,In_228,In_957);
or U1298 (N_1298,In_235,In_925);
nand U1299 (N_1299,In_54,In_483);
nor U1300 (N_1300,In_436,In_27);
nand U1301 (N_1301,In_239,In_300);
and U1302 (N_1302,In_797,In_866);
nor U1303 (N_1303,In_74,In_851);
nand U1304 (N_1304,In_897,In_421);
nor U1305 (N_1305,In_570,In_874);
and U1306 (N_1306,In_984,In_51);
nor U1307 (N_1307,In_37,In_148);
nor U1308 (N_1308,In_926,In_6);
and U1309 (N_1309,In_667,In_806);
xor U1310 (N_1310,In_808,In_502);
nand U1311 (N_1311,In_256,In_504);
nand U1312 (N_1312,In_340,In_791);
nand U1313 (N_1313,In_129,In_837);
nand U1314 (N_1314,In_788,In_647);
or U1315 (N_1315,In_730,In_909);
or U1316 (N_1316,In_312,In_439);
or U1317 (N_1317,In_14,In_928);
or U1318 (N_1318,In_302,In_714);
and U1319 (N_1319,In_815,In_571);
nor U1320 (N_1320,In_28,In_171);
nor U1321 (N_1321,In_621,In_134);
nor U1322 (N_1322,In_799,In_547);
nand U1323 (N_1323,In_456,In_553);
and U1324 (N_1324,In_367,In_680);
or U1325 (N_1325,In_290,In_801);
and U1326 (N_1326,In_968,In_394);
nor U1327 (N_1327,In_143,In_724);
or U1328 (N_1328,In_275,In_45);
xnor U1329 (N_1329,In_726,In_930);
xor U1330 (N_1330,In_929,In_975);
and U1331 (N_1331,In_684,In_713);
xor U1332 (N_1332,In_312,In_803);
xnor U1333 (N_1333,In_149,In_352);
nand U1334 (N_1334,In_279,In_260);
nand U1335 (N_1335,In_740,In_397);
xnor U1336 (N_1336,In_560,In_166);
or U1337 (N_1337,In_384,In_377);
xor U1338 (N_1338,In_962,In_672);
and U1339 (N_1339,In_738,In_721);
or U1340 (N_1340,In_436,In_681);
xor U1341 (N_1341,In_540,In_757);
xor U1342 (N_1342,In_843,In_921);
nor U1343 (N_1343,In_637,In_744);
nand U1344 (N_1344,In_208,In_556);
nor U1345 (N_1345,In_464,In_512);
xor U1346 (N_1346,In_517,In_596);
nand U1347 (N_1347,In_841,In_620);
nand U1348 (N_1348,In_10,In_162);
nand U1349 (N_1349,In_693,In_756);
nand U1350 (N_1350,In_763,In_802);
and U1351 (N_1351,In_628,In_23);
nand U1352 (N_1352,In_800,In_636);
or U1353 (N_1353,In_726,In_918);
xor U1354 (N_1354,In_995,In_987);
xnor U1355 (N_1355,In_651,In_979);
or U1356 (N_1356,In_328,In_319);
and U1357 (N_1357,In_708,In_579);
and U1358 (N_1358,In_272,In_420);
and U1359 (N_1359,In_491,In_882);
or U1360 (N_1360,In_127,In_42);
and U1361 (N_1361,In_588,In_211);
nand U1362 (N_1362,In_619,In_11);
or U1363 (N_1363,In_791,In_677);
or U1364 (N_1364,In_963,In_486);
and U1365 (N_1365,In_776,In_618);
xor U1366 (N_1366,In_937,In_289);
or U1367 (N_1367,In_826,In_842);
nand U1368 (N_1368,In_463,In_102);
and U1369 (N_1369,In_309,In_866);
nand U1370 (N_1370,In_737,In_473);
xor U1371 (N_1371,In_319,In_162);
nor U1372 (N_1372,In_192,In_818);
nor U1373 (N_1373,In_346,In_651);
and U1374 (N_1374,In_832,In_841);
nor U1375 (N_1375,In_485,In_313);
xor U1376 (N_1376,In_68,In_178);
nand U1377 (N_1377,In_339,In_512);
xnor U1378 (N_1378,In_791,In_689);
xor U1379 (N_1379,In_150,In_716);
nand U1380 (N_1380,In_701,In_912);
or U1381 (N_1381,In_297,In_673);
and U1382 (N_1382,In_651,In_934);
nand U1383 (N_1383,In_586,In_757);
nand U1384 (N_1384,In_341,In_626);
nand U1385 (N_1385,In_202,In_846);
nand U1386 (N_1386,In_634,In_531);
and U1387 (N_1387,In_907,In_262);
or U1388 (N_1388,In_372,In_578);
and U1389 (N_1389,In_482,In_688);
xnor U1390 (N_1390,In_774,In_220);
xor U1391 (N_1391,In_706,In_723);
or U1392 (N_1392,In_449,In_89);
or U1393 (N_1393,In_786,In_414);
or U1394 (N_1394,In_394,In_350);
or U1395 (N_1395,In_539,In_254);
or U1396 (N_1396,In_616,In_189);
and U1397 (N_1397,In_868,In_667);
nor U1398 (N_1398,In_314,In_295);
xnor U1399 (N_1399,In_5,In_950);
nand U1400 (N_1400,In_251,In_940);
and U1401 (N_1401,In_799,In_101);
xor U1402 (N_1402,In_51,In_983);
or U1403 (N_1403,In_257,In_158);
or U1404 (N_1404,In_570,In_203);
xnor U1405 (N_1405,In_363,In_800);
or U1406 (N_1406,In_850,In_574);
and U1407 (N_1407,In_532,In_237);
or U1408 (N_1408,In_219,In_30);
and U1409 (N_1409,In_30,In_746);
nand U1410 (N_1410,In_494,In_127);
nand U1411 (N_1411,In_819,In_579);
xor U1412 (N_1412,In_338,In_999);
and U1413 (N_1413,In_857,In_174);
nand U1414 (N_1414,In_837,In_903);
nor U1415 (N_1415,In_576,In_907);
and U1416 (N_1416,In_161,In_755);
and U1417 (N_1417,In_66,In_570);
xnor U1418 (N_1418,In_395,In_240);
nand U1419 (N_1419,In_295,In_550);
nand U1420 (N_1420,In_697,In_768);
xor U1421 (N_1421,In_235,In_476);
nand U1422 (N_1422,In_8,In_825);
and U1423 (N_1423,In_703,In_833);
xnor U1424 (N_1424,In_432,In_629);
nor U1425 (N_1425,In_161,In_954);
or U1426 (N_1426,In_495,In_863);
and U1427 (N_1427,In_935,In_669);
xnor U1428 (N_1428,In_81,In_574);
nor U1429 (N_1429,In_631,In_15);
and U1430 (N_1430,In_152,In_135);
nand U1431 (N_1431,In_275,In_260);
nand U1432 (N_1432,In_583,In_771);
nor U1433 (N_1433,In_183,In_720);
or U1434 (N_1434,In_711,In_10);
or U1435 (N_1435,In_219,In_484);
nand U1436 (N_1436,In_357,In_328);
nand U1437 (N_1437,In_87,In_746);
or U1438 (N_1438,In_430,In_970);
nand U1439 (N_1439,In_967,In_927);
nand U1440 (N_1440,In_70,In_839);
xnor U1441 (N_1441,In_928,In_722);
or U1442 (N_1442,In_729,In_192);
xnor U1443 (N_1443,In_48,In_237);
nor U1444 (N_1444,In_403,In_47);
nand U1445 (N_1445,In_711,In_534);
or U1446 (N_1446,In_950,In_439);
xnor U1447 (N_1447,In_231,In_441);
and U1448 (N_1448,In_494,In_806);
or U1449 (N_1449,In_474,In_902);
xor U1450 (N_1450,In_997,In_355);
xnor U1451 (N_1451,In_707,In_386);
or U1452 (N_1452,In_482,In_202);
and U1453 (N_1453,In_647,In_290);
and U1454 (N_1454,In_183,In_445);
nor U1455 (N_1455,In_370,In_527);
nor U1456 (N_1456,In_872,In_691);
xnor U1457 (N_1457,In_640,In_945);
nor U1458 (N_1458,In_846,In_315);
or U1459 (N_1459,In_137,In_849);
xor U1460 (N_1460,In_751,In_475);
nor U1461 (N_1461,In_229,In_646);
nand U1462 (N_1462,In_967,In_17);
or U1463 (N_1463,In_948,In_969);
and U1464 (N_1464,In_994,In_980);
xnor U1465 (N_1465,In_537,In_448);
and U1466 (N_1466,In_922,In_852);
xor U1467 (N_1467,In_116,In_603);
nand U1468 (N_1468,In_885,In_115);
nor U1469 (N_1469,In_685,In_7);
xor U1470 (N_1470,In_285,In_925);
and U1471 (N_1471,In_25,In_770);
xor U1472 (N_1472,In_441,In_492);
xor U1473 (N_1473,In_170,In_365);
and U1474 (N_1474,In_444,In_73);
nor U1475 (N_1475,In_1,In_821);
nor U1476 (N_1476,In_966,In_553);
nand U1477 (N_1477,In_675,In_442);
nand U1478 (N_1478,In_149,In_95);
and U1479 (N_1479,In_626,In_385);
nor U1480 (N_1480,In_694,In_313);
nor U1481 (N_1481,In_959,In_281);
and U1482 (N_1482,In_597,In_676);
nand U1483 (N_1483,In_709,In_349);
nor U1484 (N_1484,In_578,In_470);
xnor U1485 (N_1485,In_672,In_845);
xnor U1486 (N_1486,In_178,In_316);
nor U1487 (N_1487,In_55,In_324);
xor U1488 (N_1488,In_267,In_61);
nor U1489 (N_1489,In_94,In_524);
and U1490 (N_1490,In_8,In_230);
xor U1491 (N_1491,In_326,In_392);
or U1492 (N_1492,In_334,In_882);
or U1493 (N_1493,In_912,In_582);
nand U1494 (N_1494,In_225,In_535);
nand U1495 (N_1495,In_736,In_821);
and U1496 (N_1496,In_399,In_827);
and U1497 (N_1497,In_77,In_206);
or U1498 (N_1498,In_641,In_363);
xnor U1499 (N_1499,In_439,In_723);
nor U1500 (N_1500,In_526,In_959);
nor U1501 (N_1501,In_535,In_635);
nor U1502 (N_1502,In_724,In_969);
or U1503 (N_1503,In_593,In_896);
and U1504 (N_1504,In_270,In_426);
and U1505 (N_1505,In_16,In_413);
or U1506 (N_1506,In_557,In_247);
and U1507 (N_1507,In_588,In_615);
or U1508 (N_1508,In_895,In_550);
xor U1509 (N_1509,In_679,In_468);
nand U1510 (N_1510,In_934,In_855);
or U1511 (N_1511,In_629,In_982);
and U1512 (N_1512,In_470,In_869);
xor U1513 (N_1513,In_428,In_455);
nor U1514 (N_1514,In_47,In_792);
nor U1515 (N_1515,In_173,In_36);
nand U1516 (N_1516,In_18,In_671);
xor U1517 (N_1517,In_329,In_785);
nor U1518 (N_1518,In_366,In_384);
and U1519 (N_1519,In_93,In_535);
and U1520 (N_1520,In_307,In_495);
and U1521 (N_1521,In_77,In_430);
nand U1522 (N_1522,In_846,In_292);
xnor U1523 (N_1523,In_986,In_688);
nor U1524 (N_1524,In_212,In_955);
and U1525 (N_1525,In_822,In_710);
nand U1526 (N_1526,In_769,In_883);
or U1527 (N_1527,In_556,In_385);
nand U1528 (N_1528,In_923,In_569);
and U1529 (N_1529,In_720,In_669);
and U1530 (N_1530,In_285,In_424);
or U1531 (N_1531,In_807,In_460);
and U1532 (N_1532,In_276,In_412);
xnor U1533 (N_1533,In_382,In_45);
and U1534 (N_1534,In_293,In_658);
nor U1535 (N_1535,In_452,In_920);
nor U1536 (N_1536,In_608,In_194);
nor U1537 (N_1537,In_765,In_846);
nand U1538 (N_1538,In_553,In_439);
xnor U1539 (N_1539,In_787,In_420);
or U1540 (N_1540,In_45,In_780);
or U1541 (N_1541,In_224,In_233);
nor U1542 (N_1542,In_572,In_484);
nor U1543 (N_1543,In_619,In_107);
or U1544 (N_1544,In_495,In_382);
nand U1545 (N_1545,In_927,In_42);
nor U1546 (N_1546,In_422,In_619);
xor U1547 (N_1547,In_718,In_657);
and U1548 (N_1548,In_812,In_768);
nand U1549 (N_1549,In_91,In_253);
nand U1550 (N_1550,In_383,In_999);
nor U1551 (N_1551,In_617,In_665);
and U1552 (N_1552,In_799,In_449);
xor U1553 (N_1553,In_167,In_906);
nand U1554 (N_1554,In_696,In_158);
or U1555 (N_1555,In_997,In_965);
xnor U1556 (N_1556,In_941,In_201);
or U1557 (N_1557,In_160,In_829);
and U1558 (N_1558,In_113,In_787);
xor U1559 (N_1559,In_147,In_181);
or U1560 (N_1560,In_262,In_202);
nand U1561 (N_1561,In_74,In_351);
nor U1562 (N_1562,In_314,In_522);
xor U1563 (N_1563,In_0,In_327);
xnor U1564 (N_1564,In_243,In_881);
xor U1565 (N_1565,In_788,In_657);
xor U1566 (N_1566,In_246,In_914);
and U1567 (N_1567,In_159,In_774);
nor U1568 (N_1568,In_445,In_3);
or U1569 (N_1569,In_958,In_221);
xor U1570 (N_1570,In_312,In_970);
xnor U1571 (N_1571,In_633,In_179);
nor U1572 (N_1572,In_396,In_579);
nand U1573 (N_1573,In_856,In_962);
xor U1574 (N_1574,In_920,In_811);
or U1575 (N_1575,In_503,In_153);
xor U1576 (N_1576,In_248,In_448);
or U1577 (N_1577,In_640,In_272);
and U1578 (N_1578,In_77,In_179);
xnor U1579 (N_1579,In_237,In_801);
nor U1580 (N_1580,In_190,In_208);
nor U1581 (N_1581,In_20,In_877);
and U1582 (N_1582,In_732,In_951);
xnor U1583 (N_1583,In_154,In_45);
nand U1584 (N_1584,In_621,In_339);
nor U1585 (N_1585,In_207,In_661);
nor U1586 (N_1586,In_595,In_662);
or U1587 (N_1587,In_350,In_893);
xnor U1588 (N_1588,In_754,In_626);
and U1589 (N_1589,In_378,In_122);
or U1590 (N_1590,In_778,In_253);
and U1591 (N_1591,In_988,In_402);
nor U1592 (N_1592,In_145,In_679);
nand U1593 (N_1593,In_518,In_788);
nor U1594 (N_1594,In_990,In_833);
xor U1595 (N_1595,In_869,In_242);
or U1596 (N_1596,In_98,In_407);
and U1597 (N_1597,In_201,In_696);
and U1598 (N_1598,In_716,In_963);
nand U1599 (N_1599,In_950,In_325);
nor U1600 (N_1600,In_368,In_628);
and U1601 (N_1601,In_963,In_56);
or U1602 (N_1602,In_978,In_479);
xnor U1603 (N_1603,In_464,In_412);
or U1604 (N_1604,In_979,In_780);
xor U1605 (N_1605,In_306,In_303);
or U1606 (N_1606,In_497,In_759);
or U1607 (N_1607,In_442,In_846);
nand U1608 (N_1608,In_188,In_290);
and U1609 (N_1609,In_569,In_354);
and U1610 (N_1610,In_537,In_70);
nor U1611 (N_1611,In_816,In_964);
xnor U1612 (N_1612,In_445,In_376);
xor U1613 (N_1613,In_851,In_914);
and U1614 (N_1614,In_320,In_313);
or U1615 (N_1615,In_51,In_58);
or U1616 (N_1616,In_844,In_481);
xor U1617 (N_1617,In_898,In_524);
and U1618 (N_1618,In_240,In_241);
nand U1619 (N_1619,In_95,In_359);
nor U1620 (N_1620,In_541,In_129);
xnor U1621 (N_1621,In_219,In_827);
nor U1622 (N_1622,In_90,In_871);
and U1623 (N_1623,In_411,In_604);
and U1624 (N_1624,In_334,In_697);
nor U1625 (N_1625,In_895,In_689);
or U1626 (N_1626,In_807,In_558);
or U1627 (N_1627,In_620,In_984);
xnor U1628 (N_1628,In_991,In_308);
nand U1629 (N_1629,In_683,In_308);
or U1630 (N_1630,In_432,In_159);
nand U1631 (N_1631,In_493,In_43);
xor U1632 (N_1632,In_897,In_670);
and U1633 (N_1633,In_49,In_623);
nand U1634 (N_1634,In_728,In_830);
xnor U1635 (N_1635,In_480,In_626);
nor U1636 (N_1636,In_860,In_152);
or U1637 (N_1637,In_919,In_368);
nand U1638 (N_1638,In_557,In_742);
nand U1639 (N_1639,In_4,In_695);
xor U1640 (N_1640,In_178,In_942);
and U1641 (N_1641,In_87,In_23);
nand U1642 (N_1642,In_688,In_73);
xor U1643 (N_1643,In_808,In_749);
nand U1644 (N_1644,In_480,In_481);
nor U1645 (N_1645,In_749,In_298);
and U1646 (N_1646,In_862,In_388);
nand U1647 (N_1647,In_777,In_188);
or U1648 (N_1648,In_25,In_367);
or U1649 (N_1649,In_593,In_874);
or U1650 (N_1650,In_430,In_901);
and U1651 (N_1651,In_456,In_344);
xnor U1652 (N_1652,In_637,In_948);
nor U1653 (N_1653,In_334,In_653);
nor U1654 (N_1654,In_787,In_845);
nor U1655 (N_1655,In_395,In_457);
nor U1656 (N_1656,In_16,In_434);
nand U1657 (N_1657,In_445,In_343);
and U1658 (N_1658,In_701,In_748);
or U1659 (N_1659,In_412,In_784);
or U1660 (N_1660,In_33,In_914);
or U1661 (N_1661,In_394,In_899);
nand U1662 (N_1662,In_448,In_19);
xor U1663 (N_1663,In_560,In_137);
and U1664 (N_1664,In_387,In_573);
xor U1665 (N_1665,In_144,In_272);
and U1666 (N_1666,In_126,In_238);
or U1667 (N_1667,In_566,In_127);
xnor U1668 (N_1668,In_755,In_309);
xor U1669 (N_1669,In_91,In_520);
or U1670 (N_1670,In_764,In_915);
and U1671 (N_1671,In_8,In_608);
or U1672 (N_1672,In_768,In_949);
nand U1673 (N_1673,In_185,In_288);
and U1674 (N_1674,In_846,In_100);
nand U1675 (N_1675,In_858,In_168);
nor U1676 (N_1676,In_665,In_322);
nand U1677 (N_1677,In_921,In_695);
nor U1678 (N_1678,In_879,In_217);
or U1679 (N_1679,In_155,In_282);
xnor U1680 (N_1680,In_988,In_281);
nor U1681 (N_1681,In_407,In_972);
nor U1682 (N_1682,In_757,In_745);
nand U1683 (N_1683,In_944,In_80);
nor U1684 (N_1684,In_157,In_930);
or U1685 (N_1685,In_165,In_703);
nor U1686 (N_1686,In_46,In_404);
and U1687 (N_1687,In_293,In_878);
or U1688 (N_1688,In_448,In_190);
nand U1689 (N_1689,In_203,In_12);
or U1690 (N_1690,In_637,In_159);
xnor U1691 (N_1691,In_964,In_910);
nand U1692 (N_1692,In_235,In_230);
nand U1693 (N_1693,In_731,In_818);
xor U1694 (N_1694,In_776,In_664);
nand U1695 (N_1695,In_616,In_312);
xnor U1696 (N_1696,In_402,In_140);
xor U1697 (N_1697,In_566,In_79);
or U1698 (N_1698,In_995,In_489);
xor U1699 (N_1699,In_606,In_973);
nand U1700 (N_1700,In_198,In_613);
nand U1701 (N_1701,In_39,In_885);
or U1702 (N_1702,In_641,In_32);
and U1703 (N_1703,In_699,In_430);
nand U1704 (N_1704,In_862,In_211);
nor U1705 (N_1705,In_258,In_414);
or U1706 (N_1706,In_605,In_144);
nor U1707 (N_1707,In_344,In_347);
xor U1708 (N_1708,In_151,In_854);
nand U1709 (N_1709,In_997,In_140);
nand U1710 (N_1710,In_626,In_864);
nand U1711 (N_1711,In_967,In_924);
or U1712 (N_1712,In_292,In_578);
nand U1713 (N_1713,In_170,In_585);
or U1714 (N_1714,In_296,In_427);
xor U1715 (N_1715,In_941,In_403);
and U1716 (N_1716,In_169,In_994);
and U1717 (N_1717,In_523,In_219);
or U1718 (N_1718,In_793,In_291);
or U1719 (N_1719,In_923,In_363);
or U1720 (N_1720,In_317,In_243);
nand U1721 (N_1721,In_337,In_523);
and U1722 (N_1722,In_188,In_393);
or U1723 (N_1723,In_785,In_179);
nor U1724 (N_1724,In_599,In_536);
nor U1725 (N_1725,In_295,In_131);
or U1726 (N_1726,In_629,In_771);
nand U1727 (N_1727,In_898,In_589);
nand U1728 (N_1728,In_30,In_78);
and U1729 (N_1729,In_799,In_250);
xnor U1730 (N_1730,In_314,In_983);
and U1731 (N_1731,In_423,In_274);
or U1732 (N_1732,In_550,In_619);
and U1733 (N_1733,In_954,In_218);
xor U1734 (N_1734,In_186,In_630);
or U1735 (N_1735,In_894,In_760);
or U1736 (N_1736,In_640,In_34);
nand U1737 (N_1737,In_163,In_23);
or U1738 (N_1738,In_105,In_94);
nor U1739 (N_1739,In_777,In_506);
nand U1740 (N_1740,In_529,In_499);
xnor U1741 (N_1741,In_106,In_909);
nand U1742 (N_1742,In_240,In_243);
and U1743 (N_1743,In_582,In_835);
xnor U1744 (N_1744,In_351,In_986);
nor U1745 (N_1745,In_248,In_383);
nor U1746 (N_1746,In_842,In_30);
and U1747 (N_1747,In_332,In_102);
or U1748 (N_1748,In_169,In_835);
and U1749 (N_1749,In_714,In_291);
and U1750 (N_1750,In_142,In_320);
nand U1751 (N_1751,In_251,In_765);
xnor U1752 (N_1752,In_996,In_433);
nand U1753 (N_1753,In_441,In_211);
and U1754 (N_1754,In_641,In_989);
and U1755 (N_1755,In_249,In_887);
and U1756 (N_1756,In_689,In_179);
nor U1757 (N_1757,In_300,In_817);
or U1758 (N_1758,In_194,In_777);
nand U1759 (N_1759,In_0,In_377);
nand U1760 (N_1760,In_526,In_50);
nor U1761 (N_1761,In_659,In_104);
xnor U1762 (N_1762,In_831,In_985);
or U1763 (N_1763,In_227,In_464);
nor U1764 (N_1764,In_896,In_219);
or U1765 (N_1765,In_673,In_255);
nand U1766 (N_1766,In_722,In_844);
nor U1767 (N_1767,In_232,In_177);
or U1768 (N_1768,In_559,In_689);
and U1769 (N_1769,In_375,In_981);
and U1770 (N_1770,In_349,In_501);
and U1771 (N_1771,In_488,In_455);
or U1772 (N_1772,In_102,In_36);
or U1773 (N_1773,In_985,In_573);
and U1774 (N_1774,In_806,In_759);
nor U1775 (N_1775,In_741,In_341);
nor U1776 (N_1776,In_956,In_724);
or U1777 (N_1777,In_526,In_352);
or U1778 (N_1778,In_587,In_752);
or U1779 (N_1779,In_3,In_440);
and U1780 (N_1780,In_278,In_140);
or U1781 (N_1781,In_895,In_806);
or U1782 (N_1782,In_971,In_910);
xnor U1783 (N_1783,In_978,In_496);
and U1784 (N_1784,In_754,In_426);
nand U1785 (N_1785,In_546,In_236);
xnor U1786 (N_1786,In_54,In_792);
and U1787 (N_1787,In_698,In_156);
or U1788 (N_1788,In_42,In_769);
and U1789 (N_1789,In_67,In_731);
nor U1790 (N_1790,In_909,In_940);
or U1791 (N_1791,In_112,In_986);
xor U1792 (N_1792,In_317,In_178);
nand U1793 (N_1793,In_515,In_826);
or U1794 (N_1794,In_396,In_445);
nand U1795 (N_1795,In_21,In_403);
nand U1796 (N_1796,In_46,In_652);
or U1797 (N_1797,In_709,In_473);
xor U1798 (N_1798,In_602,In_778);
nor U1799 (N_1799,In_76,In_230);
or U1800 (N_1800,In_237,In_511);
nand U1801 (N_1801,In_667,In_46);
nor U1802 (N_1802,In_945,In_385);
nand U1803 (N_1803,In_533,In_943);
nand U1804 (N_1804,In_507,In_73);
nand U1805 (N_1805,In_441,In_426);
and U1806 (N_1806,In_899,In_604);
nand U1807 (N_1807,In_673,In_696);
nor U1808 (N_1808,In_30,In_898);
xor U1809 (N_1809,In_570,In_812);
nor U1810 (N_1810,In_533,In_768);
xor U1811 (N_1811,In_730,In_571);
and U1812 (N_1812,In_266,In_301);
nor U1813 (N_1813,In_137,In_306);
nand U1814 (N_1814,In_539,In_811);
nand U1815 (N_1815,In_209,In_333);
or U1816 (N_1816,In_328,In_205);
or U1817 (N_1817,In_639,In_915);
xnor U1818 (N_1818,In_976,In_304);
and U1819 (N_1819,In_835,In_305);
xor U1820 (N_1820,In_421,In_95);
and U1821 (N_1821,In_973,In_969);
nor U1822 (N_1822,In_355,In_226);
nor U1823 (N_1823,In_964,In_585);
and U1824 (N_1824,In_60,In_566);
and U1825 (N_1825,In_593,In_843);
nand U1826 (N_1826,In_207,In_356);
and U1827 (N_1827,In_985,In_320);
xnor U1828 (N_1828,In_750,In_990);
nor U1829 (N_1829,In_872,In_253);
nand U1830 (N_1830,In_366,In_94);
xnor U1831 (N_1831,In_705,In_710);
nor U1832 (N_1832,In_992,In_321);
xnor U1833 (N_1833,In_408,In_610);
xnor U1834 (N_1834,In_597,In_757);
or U1835 (N_1835,In_787,In_552);
or U1836 (N_1836,In_54,In_574);
and U1837 (N_1837,In_238,In_653);
or U1838 (N_1838,In_836,In_437);
and U1839 (N_1839,In_429,In_727);
and U1840 (N_1840,In_525,In_729);
nor U1841 (N_1841,In_157,In_661);
or U1842 (N_1842,In_116,In_859);
xor U1843 (N_1843,In_449,In_860);
or U1844 (N_1844,In_327,In_917);
nand U1845 (N_1845,In_386,In_511);
nand U1846 (N_1846,In_340,In_442);
nand U1847 (N_1847,In_672,In_857);
nor U1848 (N_1848,In_931,In_604);
and U1849 (N_1849,In_236,In_1);
xnor U1850 (N_1850,In_280,In_231);
or U1851 (N_1851,In_269,In_823);
and U1852 (N_1852,In_730,In_967);
xor U1853 (N_1853,In_536,In_541);
xnor U1854 (N_1854,In_570,In_126);
and U1855 (N_1855,In_475,In_536);
or U1856 (N_1856,In_672,In_445);
nand U1857 (N_1857,In_670,In_823);
nand U1858 (N_1858,In_988,In_584);
nor U1859 (N_1859,In_614,In_97);
or U1860 (N_1860,In_468,In_771);
or U1861 (N_1861,In_290,In_993);
xnor U1862 (N_1862,In_53,In_2);
or U1863 (N_1863,In_98,In_43);
nor U1864 (N_1864,In_774,In_906);
and U1865 (N_1865,In_262,In_597);
xor U1866 (N_1866,In_769,In_736);
nand U1867 (N_1867,In_349,In_415);
nand U1868 (N_1868,In_938,In_127);
nor U1869 (N_1869,In_764,In_144);
xor U1870 (N_1870,In_683,In_841);
xor U1871 (N_1871,In_513,In_605);
or U1872 (N_1872,In_771,In_115);
xor U1873 (N_1873,In_639,In_878);
xor U1874 (N_1874,In_385,In_991);
nor U1875 (N_1875,In_67,In_860);
nor U1876 (N_1876,In_16,In_917);
and U1877 (N_1877,In_425,In_308);
nand U1878 (N_1878,In_302,In_604);
nand U1879 (N_1879,In_944,In_762);
and U1880 (N_1880,In_618,In_792);
nand U1881 (N_1881,In_342,In_717);
or U1882 (N_1882,In_617,In_122);
xor U1883 (N_1883,In_407,In_444);
xor U1884 (N_1884,In_969,In_883);
nor U1885 (N_1885,In_169,In_284);
nor U1886 (N_1886,In_249,In_176);
xnor U1887 (N_1887,In_799,In_229);
nand U1888 (N_1888,In_702,In_433);
nor U1889 (N_1889,In_752,In_88);
and U1890 (N_1890,In_431,In_873);
xnor U1891 (N_1891,In_616,In_954);
nor U1892 (N_1892,In_446,In_292);
nand U1893 (N_1893,In_333,In_387);
nand U1894 (N_1894,In_469,In_669);
nand U1895 (N_1895,In_446,In_467);
and U1896 (N_1896,In_462,In_837);
or U1897 (N_1897,In_981,In_46);
xnor U1898 (N_1898,In_522,In_738);
and U1899 (N_1899,In_247,In_731);
and U1900 (N_1900,In_108,In_669);
xor U1901 (N_1901,In_199,In_14);
nand U1902 (N_1902,In_478,In_777);
or U1903 (N_1903,In_794,In_188);
nand U1904 (N_1904,In_491,In_66);
nor U1905 (N_1905,In_164,In_235);
or U1906 (N_1906,In_193,In_350);
nor U1907 (N_1907,In_695,In_10);
nand U1908 (N_1908,In_145,In_549);
nand U1909 (N_1909,In_796,In_630);
or U1910 (N_1910,In_120,In_956);
or U1911 (N_1911,In_82,In_644);
xor U1912 (N_1912,In_17,In_996);
nor U1913 (N_1913,In_715,In_324);
or U1914 (N_1914,In_152,In_169);
nor U1915 (N_1915,In_762,In_787);
nor U1916 (N_1916,In_479,In_470);
and U1917 (N_1917,In_944,In_237);
nor U1918 (N_1918,In_528,In_208);
nand U1919 (N_1919,In_347,In_241);
nand U1920 (N_1920,In_915,In_127);
nor U1921 (N_1921,In_444,In_475);
xnor U1922 (N_1922,In_264,In_68);
xnor U1923 (N_1923,In_425,In_138);
and U1924 (N_1924,In_521,In_308);
nand U1925 (N_1925,In_975,In_231);
and U1926 (N_1926,In_574,In_357);
or U1927 (N_1927,In_693,In_831);
nand U1928 (N_1928,In_133,In_514);
or U1929 (N_1929,In_980,In_58);
nor U1930 (N_1930,In_428,In_618);
nand U1931 (N_1931,In_18,In_377);
and U1932 (N_1932,In_738,In_737);
or U1933 (N_1933,In_655,In_879);
nor U1934 (N_1934,In_408,In_828);
nand U1935 (N_1935,In_293,In_891);
nor U1936 (N_1936,In_718,In_668);
nor U1937 (N_1937,In_476,In_627);
or U1938 (N_1938,In_51,In_446);
xnor U1939 (N_1939,In_545,In_460);
nand U1940 (N_1940,In_901,In_958);
or U1941 (N_1941,In_841,In_333);
and U1942 (N_1942,In_28,In_761);
and U1943 (N_1943,In_49,In_650);
or U1944 (N_1944,In_928,In_305);
and U1945 (N_1945,In_703,In_84);
xnor U1946 (N_1946,In_254,In_93);
nor U1947 (N_1947,In_727,In_925);
xnor U1948 (N_1948,In_40,In_104);
xor U1949 (N_1949,In_252,In_582);
nand U1950 (N_1950,In_624,In_280);
nor U1951 (N_1951,In_797,In_690);
nand U1952 (N_1952,In_866,In_694);
xor U1953 (N_1953,In_47,In_458);
xnor U1954 (N_1954,In_290,In_656);
nor U1955 (N_1955,In_599,In_438);
xnor U1956 (N_1956,In_222,In_876);
or U1957 (N_1957,In_714,In_403);
nand U1958 (N_1958,In_809,In_730);
xor U1959 (N_1959,In_801,In_765);
nand U1960 (N_1960,In_123,In_606);
xor U1961 (N_1961,In_539,In_133);
xor U1962 (N_1962,In_17,In_34);
xor U1963 (N_1963,In_837,In_685);
nand U1964 (N_1964,In_848,In_168);
or U1965 (N_1965,In_678,In_38);
or U1966 (N_1966,In_177,In_664);
or U1967 (N_1967,In_435,In_179);
nor U1968 (N_1968,In_748,In_286);
or U1969 (N_1969,In_531,In_97);
nor U1970 (N_1970,In_315,In_361);
and U1971 (N_1971,In_542,In_746);
nor U1972 (N_1972,In_978,In_964);
nor U1973 (N_1973,In_662,In_775);
xor U1974 (N_1974,In_996,In_69);
nand U1975 (N_1975,In_437,In_431);
xnor U1976 (N_1976,In_266,In_332);
xnor U1977 (N_1977,In_66,In_690);
and U1978 (N_1978,In_849,In_103);
or U1979 (N_1979,In_148,In_120);
and U1980 (N_1980,In_784,In_640);
and U1981 (N_1981,In_456,In_157);
nand U1982 (N_1982,In_214,In_946);
and U1983 (N_1983,In_523,In_437);
or U1984 (N_1984,In_586,In_492);
or U1985 (N_1985,In_235,In_367);
or U1986 (N_1986,In_390,In_665);
nand U1987 (N_1987,In_616,In_959);
xnor U1988 (N_1988,In_522,In_807);
nand U1989 (N_1989,In_254,In_792);
nor U1990 (N_1990,In_202,In_959);
nand U1991 (N_1991,In_729,In_273);
nor U1992 (N_1992,In_385,In_540);
nand U1993 (N_1993,In_878,In_50);
xor U1994 (N_1994,In_478,In_674);
xor U1995 (N_1995,In_82,In_791);
xor U1996 (N_1996,In_205,In_272);
or U1997 (N_1997,In_265,In_996);
and U1998 (N_1998,In_898,In_949);
and U1999 (N_1999,In_874,In_641);
nor U2000 (N_2000,In_733,In_500);
nand U2001 (N_2001,In_928,In_103);
xor U2002 (N_2002,In_174,In_634);
xor U2003 (N_2003,In_789,In_788);
and U2004 (N_2004,In_749,In_566);
nor U2005 (N_2005,In_169,In_112);
nor U2006 (N_2006,In_749,In_91);
and U2007 (N_2007,In_58,In_886);
nand U2008 (N_2008,In_128,In_408);
xor U2009 (N_2009,In_946,In_210);
nor U2010 (N_2010,In_835,In_336);
nand U2011 (N_2011,In_68,In_344);
nor U2012 (N_2012,In_991,In_883);
xor U2013 (N_2013,In_950,In_123);
nor U2014 (N_2014,In_826,In_565);
xnor U2015 (N_2015,In_186,In_713);
nor U2016 (N_2016,In_314,In_219);
and U2017 (N_2017,In_682,In_108);
xnor U2018 (N_2018,In_56,In_117);
or U2019 (N_2019,In_650,In_627);
xnor U2020 (N_2020,In_561,In_804);
or U2021 (N_2021,In_243,In_673);
nor U2022 (N_2022,In_895,In_245);
nor U2023 (N_2023,In_845,In_170);
and U2024 (N_2024,In_735,In_982);
xor U2025 (N_2025,In_583,In_662);
or U2026 (N_2026,In_232,In_804);
or U2027 (N_2027,In_945,In_837);
and U2028 (N_2028,In_719,In_611);
xor U2029 (N_2029,In_365,In_910);
nor U2030 (N_2030,In_15,In_11);
or U2031 (N_2031,In_880,In_563);
and U2032 (N_2032,In_440,In_769);
and U2033 (N_2033,In_721,In_800);
or U2034 (N_2034,In_642,In_427);
or U2035 (N_2035,In_665,In_263);
and U2036 (N_2036,In_493,In_121);
or U2037 (N_2037,In_440,In_547);
and U2038 (N_2038,In_287,In_844);
and U2039 (N_2039,In_525,In_202);
and U2040 (N_2040,In_556,In_15);
and U2041 (N_2041,In_658,In_104);
or U2042 (N_2042,In_916,In_396);
xor U2043 (N_2043,In_231,In_208);
or U2044 (N_2044,In_868,In_976);
xor U2045 (N_2045,In_178,In_620);
and U2046 (N_2046,In_120,In_297);
and U2047 (N_2047,In_868,In_289);
nand U2048 (N_2048,In_811,In_236);
nand U2049 (N_2049,In_215,In_891);
xnor U2050 (N_2050,In_872,In_645);
nand U2051 (N_2051,In_699,In_887);
and U2052 (N_2052,In_410,In_946);
xnor U2053 (N_2053,In_978,In_72);
and U2054 (N_2054,In_270,In_229);
xor U2055 (N_2055,In_443,In_8);
or U2056 (N_2056,In_958,In_865);
or U2057 (N_2057,In_227,In_378);
nor U2058 (N_2058,In_131,In_21);
or U2059 (N_2059,In_92,In_166);
or U2060 (N_2060,In_639,In_49);
and U2061 (N_2061,In_823,In_292);
and U2062 (N_2062,In_810,In_388);
and U2063 (N_2063,In_197,In_656);
or U2064 (N_2064,In_421,In_519);
xor U2065 (N_2065,In_239,In_699);
or U2066 (N_2066,In_780,In_753);
and U2067 (N_2067,In_815,In_408);
nand U2068 (N_2068,In_257,In_306);
nand U2069 (N_2069,In_44,In_288);
xnor U2070 (N_2070,In_68,In_889);
and U2071 (N_2071,In_800,In_951);
xor U2072 (N_2072,In_530,In_541);
nor U2073 (N_2073,In_408,In_5);
or U2074 (N_2074,In_845,In_182);
nand U2075 (N_2075,In_593,In_406);
or U2076 (N_2076,In_290,In_568);
nand U2077 (N_2077,In_794,In_52);
nand U2078 (N_2078,In_609,In_778);
xor U2079 (N_2079,In_339,In_700);
nand U2080 (N_2080,In_329,In_919);
or U2081 (N_2081,In_324,In_398);
nor U2082 (N_2082,In_543,In_283);
nand U2083 (N_2083,In_164,In_587);
nor U2084 (N_2084,In_285,In_768);
or U2085 (N_2085,In_55,In_158);
and U2086 (N_2086,In_543,In_887);
nand U2087 (N_2087,In_916,In_221);
xnor U2088 (N_2088,In_399,In_828);
or U2089 (N_2089,In_612,In_245);
and U2090 (N_2090,In_555,In_881);
nor U2091 (N_2091,In_166,In_22);
nand U2092 (N_2092,In_113,In_361);
nor U2093 (N_2093,In_111,In_640);
and U2094 (N_2094,In_339,In_206);
nor U2095 (N_2095,In_14,In_90);
nor U2096 (N_2096,In_189,In_947);
nor U2097 (N_2097,In_479,In_910);
xor U2098 (N_2098,In_316,In_591);
or U2099 (N_2099,In_700,In_587);
and U2100 (N_2100,In_177,In_417);
xnor U2101 (N_2101,In_788,In_939);
xor U2102 (N_2102,In_100,In_213);
nor U2103 (N_2103,In_236,In_428);
nand U2104 (N_2104,In_847,In_477);
and U2105 (N_2105,In_370,In_887);
xnor U2106 (N_2106,In_35,In_989);
nor U2107 (N_2107,In_145,In_238);
nand U2108 (N_2108,In_655,In_374);
nand U2109 (N_2109,In_428,In_484);
nor U2110 (N_2110,In_842,In_865);
nand U2111 (N_2111,In_24,In_666);
nor U2112 (N_2112,In_625,In_235);
xor U2113 (N_2113,In_48,In_394);
and U2114 (N_2114,In_394,In_572);
xor U2115 (N_2115,In_769,In_342);
or U2116 (N_2116,In_37,In_24);
and U2117 (N_2117,In_989,In_545);
or U2118 (N_2118,In_84,In_185);
or U2119 (N_2119,In_395,In_345);
and U2120 (N_2120,In_716,In_264);
xnor U2121 (N_2121,In_385,In_162);
nand U2122 (N_2122,In_204,In_729);
xnor U2123 (N_2123,In_218,In_342);
nor U2124 (N_2124,In_487,In_218);
and U2125 (N_2125,In_273,In_97);
xor U2126 (N_2126,In_688,In_990);
or U2127 (N_2127,In_321,In_58);
nor U2128 (N_2128,In_425,In_61);
and U2129 (N_2129,In_371,In_151);
nand U2130 (N_2130,In_760,In_806);
nor U2131 (N_2131,In_544,In_624);
xor U2132 (N_2132,In_716,In_533);
nand U2133 (N_2133,In_988,In_189);
or U2134 (N_2134,In_677,In_431);
xnor U2135 (N_2135,In_131,In_524);
and U2136 (N_2136,In_105,In_541);
nand U2137 (N_2137,In_442,In_34);
xor U2138 (N_2138,In_228,In_690);
nand U2139 (N_2139,In_983,In_2);
nand U2140 (N_2140,In_697,In_207);
or U2141 (N_2141,In_992,In_545);
and U2142 (N_2142,In_610,In_699);
and U2143 (N_2143,In_405,In_730);
nor U2144 (N_2144,In_896,In_766);
nor U2145 (N_2145,In_240,In_456);
nand U2146 (N_2146,In_283,In_645);
and U2147 (N_2147,In_230,In_680);
xnor U2148 (N_2148,In_916,In_358);
and U2149 (N_2149,In_502,In_292);
xnor U2150 (N_2150,In_5,In_81);
and U2151 (N_2151,In_365,In_142);
nor U2152 (N_2152,In_640,In_49);
xor U2153 (N_2153,In_396,In_54);
xor U2154 (N_2154,In_17,In_748);
xor U2155 (N_2155,In_468,In_178);
or U2156 (N_2156,In_133,In_606);
and U2157 (N_2157,In_135,In_635);
and U2158 (N_2158,In_69,In_281);
nand U2159 (N_2159,In_423,In_995);
nor U2160 (N_2160,In_41,In_281);
and U2161 (N_2161,In_829,In_353);
nor U2162 (N_2162,In_699,In_553);
nand U2163 (N_2163,In_263,In_508);
nor U2164 (N_2164,In_131,In_183);
nand U2165 (N_2165,In_292,In_902);
xor U2166 (N_2166,In_103,In_26);
nand U2167 (N_2167,In_438,In_956);
or U2168 (N_2168,In_835,In_328);
nor U2169 (N_2169,In_321,In_775);
nor U2170 (N_2170,In_19,In_466);
xor U2171 (N_2171,In_932,In_781);
and U2172 (N_2172,In_926,In_928);
or U2173 (N_2173,In_21,In_561);
nand U2174 (N_2174,In_491,In_960);
and U2175 (N_2175,In_688,In_971);
and U2176 (N_2176,In_617,In_261);
nand U2177 (N_2177,In_601,In_330);
xnor U2178 (N_2178,In_361,In_777);
xor U2179 (N_2179,In_222,In_71);
or U2180 (N_2180,In_226,In_698);
or U2181 (N_2181,In_674,In_742);
nand U2182 (N_2182,In_374,In_280);
or U2183 (N_2183,In_929,In_22);
and U2184 (N_2184,In_715,In_149);
or U2185 (N_2185,In_151,In_139);
or U2186 (N_2186,In_862,In_998);
xnor U2187 (N_2187,In_437,In_355);
nand U2188 (N_2188,In_804,In_530);
nand U2189 (N_2189,In_53,In_580);
or U2190 (N_2190,In_140,In_385);
nand U2191 (N_2191,In_613,In_820);
or U2192 (N_2192,In_640,In_595);
xnor U2193 (N_2193,In_140,In_792);
and U2194 (N_2194,In_726,In_139);
nand U2195 (N_2195,In_775,In_245);
and U2196 (N_2196,In_734,In_342);
and U2197 (N_2197,In_487,In_618);
or U2198 (N_2198,In_351,In_862);
xnor U2199 (N_2199,In_496,In_454);
nand U2200 (N_2200,In_684,In_560);
nor U2201 (N_2201,In_906,In_509);
or U2202 (N_2202,In_667,In_273);
or U2203 (N_2203,In_86,In_646);
nand U2204 (N_2204,In_182,In_723);
or U2205 (N_2205,In_115,In_37);
and U2206 (N_2206,In_156,In_456);
or U2207 (N_2207,In_190,In_697);
nand U2208 (N_2208,In_494,In_902);
xor U2209 (N_2209,In_869,In_299);
nor U2210 (N_2210,In_133,In_941);
and U2211 (N_2211,In_983,In_277);
nand U2212 (N_2212,In_128,In_349);
nor U2213 (N_2213,In_490,In_455);
xnor U2214 (N_2214,In_779,In_116);
and U2215 (N_2215,In_574,In_381);
xnor U2216 (N_2216,In_491,In_181);
xor U2217 (N_2217,In_337,In_956);
nand U2218 (N_2218,In_146,In_135);
nor U2219 (N_2219,In_710,In_554);
and U2220 (N_2220,In_108,In_329);
nor U2221 (N_2221,In_267,In_885);
nor U2222 (N_2222,In_844,In_772);
xnor U2223 (N_2223,In_841,In_952);
xnor U2224 (N_2224,In_739,In_60);
nand U2225 (N_2225,In_12,In_166);
and U2226 (N_2226,In_588,In_209);
or U2227 (N_2227,In_189,In_770);
or U2228 (N_2228,In_468,In_499);
and U2229 (N_2229,In_89,In_210);
and U2230 (N_2230,In_77,In_394);
nand U2231 (N_2231,In_365,In_359);
and U2232 (N_2232,In_693,In_875);
or U2233 (N_2233,In_68,In_265);
nor U2234 (N_2234,In_531,In_795);
nand U2235 (N_2235,In_402,In_365);
xor U2236 (N_2236,In_511,In_199);
nor U2237 (N_2237,In_729,In_863);
or U2238 (N_2238,In_643,In_641);
nor U2239 (N_2239,In_95,In_405);
xnor U2240 (N_2240,In_76,In_118);
and U2241 (N_2241,In_558,In_491);
nand U2242 (N_2242,In_274,In_844);
nor U2243 (N_2243,In_660,In_184);
xor U2244 (N_2244,In_416,In_130);
or U2245 (N_2245,In_593,In_305);
and U2246 (N_2246,In_407,In_200);
nand U2247 (N_2247,In_597,In_95);
nor U2248 (N_2248,In_842,In_944);
xor U2249 (N_2249,In_481,In_215);
and U2250 (N_2250,In_548,In_3);
or U2251 (N_2251,In_129,In_920);
nand U2252 (N_2252,In_948,In_297);
nor U2253 (N_2253,In_511,In_759);
nand U2254 (N_2254,In_204,In_905);
and U2255 (N_2255,In_638,In_827);
and U2256 (N_2256,In_171,In_106);
and U2257 (N_2257,In_491,In_649);
and U2258 (N_2258,In_810,In_832);
nand U2259 (N_2259,In_354,In_365);
nand U2260 (N_2260,In_194,In_169);
or U2261 (N_2261,In_62,In_607);
xnor U2262 (N_2262,In_37,In_734);
and U2263 (N_2263,In_339,In_831);
and U2264 (N_2264,In_711,In_743);
and U2265 (N_2265,In_71,In_49);
or U2266 (N_2266,In_834,In_19);
and U2267 (N_2267,In_488,In_106);
xor U2268 (N_2268,In_309,In_981);
or U2269 (N_2269,In_166,In_911);
nand U2270 (N_2270,In_777,In_325);
nor U2271 (N_2271,In_897,In_965);
nand U2272 (N_2272,In_737,In_64);
and U2273 (N_2273,In_667,In_293);
xor U2274 (N_2274,In_648,In_175);
xnor U2275 (N_2275,In_949,In_508);
xor U2276 (N_2276,In_873,In_855);
and U2277 (N_2277,In_43,In_490);
nor U2278 (N_2278,In_49,In_508);
xnor U2279 (N_2279,In_517,In_190);
or U2280 (N_2280,In_946,In_686);
or U2281 (N_2281,In_208,In_428);
and U2282 (N_2282,In_619,In_248);
nand U2283 (N_2283,In_637,In_95);
nand U2284 (N_2284,In_551,In_986);
xnor U2285 (N_2285,In_331,In_245);
nand U2286 (N_2286,In_243,In_43);
or U2287 (N_2287,In_74,In_849);
and U2288 (N_2288,In_392,In_445);
xor U2289 (N_2289,In_240,In_79);
xnor U2290 (N_2290,In_500,In_405);
or U2291 (N_2291,In_678,In_994);
nor U2292 (N_2292,In_784,In_761);
nand U2293 (N_2293,In_420,In_900);
nor U2294 (N_2294,In_759,In_794);
or U2295 (N_2295,In_408,In_457);
and U2296 (N_2296,In_786,In_517);
and U2297 (N_2297,In_490,In_72);
or U2298 (N_2298,In_928,In_168);
or U2299 (N_2299,In_398,In_608);
and U2300 (N_2300,In_432,In_191);
xor U2301 (N_2301,In_183,In_148);
nor U2302 (N_2302,In_441,In_163);
or U2303 (N_2303,In_765,In_916);
xnor U2304 (N_2304,In_651,In_177);
and U2305 (N_2305,In_504,In_167);
nand U2306 (N_2306,In_914,In_2);
or U2307 (N_2307,In_376,In_448);
nand U2308 (N_2308,In_571,In_586);
and U2309 (N_2309,In_131,In_822);
xnor U2310 (N_2310,In_382,In_184);
nand U2311 (N_2311,In_55,In_444);
nor U2312 (N_2312,In_631,In_946);
and U2313 (N_2313,In_340,In_266);
nand U2314 (N_2314,In_602,In_187);
nor U2315 (N_2315,In_89,In_239);
or U2316 (N_2316,In_439,In_258);
or U2317 (N_2317,In_780,In_240);
nor U2318 (N_2318,In_337,In_361);
and U2319 (N_2319,In_535,In_189);
or U2320 (N_2320,In_638,In_411);
or U2321 (N_2321,In_276,In_459);
xnor U2322 (N_2322,In_389,In_607);
nand U2323 (N_2323,In_428,In_0);
xor U2324 (N_2324,In_289,In_684);
nor U2325 (N_2325,In_7,In_89);
and U2326 (N_2326,In_270,In_728);
or U2327 (N_2327,In_48,In_483);
nor U2328 (N_2328,In_883,In_861);
or U2329 (N_2329,In_761,In_562);
and U2330 (N_2330,In_409,In_156);
or U2331 (N_2331,In_229,In_161);
nand U2332 (N_2332,In_763,In_436);
nor U2333 (N_2333,In_142,In_537);
and U2334 (N_2334,In_537,In_336);
nor U2335 (N_2335,In_809,In_162);
nand U2336 (N_2336,In_806,In_434);
and U2337 (N_2337,In_163,In_940);
nand U2338 (N_2338,In_495,In_53);
xor U2339 (N_2339,In_507,In_72);
nor U2340 (N_2340,In_302,In_408);
or U2341 (N_2341,In_263,In_62);
nand U2342 (N_2342,In_136,In_624);
and U2343 (N_2343,In_292,In_665);
and U2344 (N_2344,In_952,In_487);
nor U2345 (N_2345,In_281,In_933);
nand U2346 (N_2346,In_438,In_993);
nand U2347 (N_2347,In_867,In_193);
nor U2348 (N_2348,In_404,In_568);
nor U2349 (N_2349,In_674,In_924);
or U2350 (N_2350,In_707,In_469);
and U2351 (N_2351,In_390,In_154);
or U2352 (N_2352,In_181,In_881);
and U2353 (N_2353,In_379,In_588);
or U2354 (N_2354,In_505,In_890);
nor U2355 (N_2355,In_381,In_864);
nor U2356 (N_2356,In_284,In_39);
and U2357 (N_2357,In_847,In_580);
and U2358 (N_2358,In_224,In_755);
and U2359 (N_2359,In_822,In_259);
xor U2360 (N_2360,In_221,In_26);
and U2361 (N_2361,In_494,In_195);
and U2362 (N_2362,In_68,In_397);
nand U2363 (N_2363,In_667,In_60);
and U2364 (N_2364,In_806,In_18);
or U2365 (N_2365,In_875,In_226);
or U2366 (N_2366,In_657,In_480);
nor U2367 (N_2367,In_490,In_884);
or U2368 (N_2368,In_884,In_386);
nor U2369 (N_2369,In_245,In_74);
or U2370 (N_2370,In_256,In_300);
nand U2371 (N_2371,In_635,In_250);
and U2372 (N_2372,In_924,In_775);
or U2373 (N_2373,In_230,In_49);
and U2374 (N_2374,In_634,In_785);
or U2375 (N_2375,In_397,In_392);
and U2376 (N_2376,In_755,In_128);
nor U2377 (N_2377,In_146,In_929);
xor U2378 (N_2378,In_867,In_917);
or U2379 (N_2379,In_12,In_924);
and U2380 (N_2380,In_176,In_768);
and U2381 (N_2381,In_225,In_34);
and U2382 (N_2382,In_275,In_245);
nor U2383 (N_2383,In_51,In_280);
xnor U2384 (N_2384,In_285,In_366);
nand U2385 (N_2385,In_814,In_427);
xor U2386 (N_2386,In_558,In_81);
and U2387 (N_2387,In_560,In_565);
and U2388 (N_2388,In_233,In_984);
xnor U2389 (N_2389,In_699,In_397);
or U2390 (N_2390,In_969,In_693);
nand U2391 (N_2391,In_312,In_515);
xor U2392 (N_2392,In_712,In_371);
xor U2393 (N_2393,In_45,In_153);
nand U2394 (N_2394,In_789,In_144);
xor U2395 (N_2395,In_752,In_274);
nand U2396 (N_2396,In_925,In_22);
or U2397 (N_2397,In_338,In_595);
or U2398 (N_2398,In_506,In_332);
or U2399 (N_2399,In_167,In_4);
and U2400 (N_2400,In_912,In_63);
nand U2401 (N_2401,In_18,In_261);
or U2402 (N_2402,In_310,In_724);
xor U2403 (N_2403,In_430,In_278);
or U2404 (N_2404,In_194,In_150);
xnor U2405 (N_2405,In_6,In_394);
or U2406 (N_2406,In_765,In_864);
nor U2407 (N_2407,In_150,In_65);
or U2408 (N_2408,In_802,In_975);
or U2409 (N_2409,In_445,In_227);
nor U2410 (N_2410,In_819,In_808);
and U2411 (N_2411,In_400,In_873);
xnor U2412 (N_2412,In_889,In_351);
xnor U2413 (N_2413,In_891,In_388);
and U2414 (N_2414,In_606,In_403);
xor U2415 (N_2415,In_994,In_503);
and U2416 (N_2416,In_332,In_106);
or U2417 (N_2417,In_944,In_721);
and U2418 (N_2418,In_197,In_837);
nand U2419 (N_2419,In_691,In_886);
nand U2420 (N_2420,In_670,In_388);
and U2421 (N_2421,In_473,In_677);
or U2422 (N_2422,In_404,In_965);
or U2423 (N_2423,In_281,In_210);
nor U2424 (N_2424,In_939,In_553);
or U2425 (N_2425,In_620,In_838);
xnor U2426 (N_2426,In_593,In_448);
or U2427 (N_2427,In_294,In_253);
nor U2428 (N_2428,In_217,In_731);
or U2429 (N_2429,In_444,In_196);
nand U2430 (N_2430,In_34,In_305);
nor U2431 (N_2431,In_683,In_431);
nand U2432 (N_2432,In_836,In_15);
nor U2433 (N_2433,In_775,In_208);
nand U2434 (N_2434,In_994,In_52);
or U2435 (N_2435,In_313,In_695);
nand U2436 (N_2436,In_479,In_310);
xnor U2437 (N_2437,In_348,In_71);
xor U2438 (N_2438,In_5,In_185);
xnor U2439 (N_2439,In_904,In_852);
or U2440 (N_2440,In_942,In_635);
nand U2441 (N_2441,In_950,In_9);
and U2442 (N_2442,In_838,In_484);
nor U2443 (N_2443,In_230,In_246);
nor U2444 (N_2444,In_56,In_846);
xor U2445 (N_2445,In_292,In_395);
nor U2446 (N_2446,In_193,In_400);
nand U2447 (N_2447,In_668,In_376);
nor U2448 (N_2448,In_8,In_788);
or U2449 (N_2449,In_918,In_957);
and U2450 (N_2450,In_79,In_277);
and U2451 (N_2451,In_636,In_794);
or U2452 (N_2452,In_15,In_194);
xnor U2453 (N_2453,In_56,In_19);
or U2454 (N_2454,In_649,In_635);
nor U2455 (N_2455,In_55,In_655);
and U2456 (N_2456,In_230,In_877);
or U2457 (N_2457,In_53,In_247);
nor U2458 (N_2458,In_954,In_792);
or U2459 (N_2459,In_598,In_198);
or U2460 (N_2460,In_149,In_32);
or U2461 (N_2461,In_190,In_211);
xor U2462 (N_2462,In_133,In_619);
or U2463 (N_2463,In_741,In_253);
or U2464 (N_2464,In_908,In_360);
nand U2465 (N_2465,In_628,In_673);
and U2466 (N_2466,In_989,In_505);
nand U2467 (N_2467,In_418,In_545);
nand U2468 (N_2468,In_809,In_350);
xnor U2469 (N_2469,In_86,In_946);
nor U2470 (N_2470,In_577,In_444);
nand U2471 (N_2471,In_975,In_640);
nand U2472 (N_2472,In_484,In_559);
xnor U2473 (N_2473,In_950,In_899);
or U2474 (N_2474,In_877,In_241);
nand U2475 (N_2475,In_416,In_784);
xor U2476 (N_2476,In_615,In_708);
and U2477 (N_2477,In_523,In_146);
and U2478 (N_2478,In_952,In_259);
xor U2479 (N_2479,In_960,In_412);
or U2480 (N_2480,In_33,In_730);
or U2481 (N_2481,In_809,In_862);
and U2482 (N_2482,In_783,In_683);
nor U2483 (N_2483,In_899,In_689);
or U2484 (N_2484,In_198,In_832);
xor U2485 (N_2485,In_961,In_150);
xnor U2486 (N_2486,In_133,In_604);
and U2487 (N_2487,In_838,In_320);
nand U2488 (N_2488,In_620,In_250);
xor U2489 (N_2489,In_228,In_478);
or U2490 (N_2490,In_897,In_74);
nand U2491 (N_2491,In_764,In_98);
nand U2492 (N_2492,In_950,In_984);
and U2493 (N_2493,In_331,In_736);
or U2494 (N_2494,In_310,In_980);
and U2495 (N_2495,In_680,In_378);
xnor U2496 (N_2496,In_695,In_923);
or U2497 (N_2497,In_549,In_799);
nand U2498 (N_2498,In_864,In_658);
xor U2499 (N_2499,In_181,In_538);
or U2500 (N_2500,In_32,In_364);
and U2501 (N_2501,In_886,In_758);
or U2502 (N_2502,In_460,In_881);
nor U2503 (N_2503,In_803,In_648);
nand U2504 (N_2504,In_899,In_559);
xnor U2505 (N_2505,In_623,In_923);
nand U2506 (N_2506,In_937,In_362);
nand U2507 (N_2507,In_173,In_548);
nor U2508 (N_2508,In_320,In_405);
nand U2509 (N_2509,In_648,In_772);
xnor U2510 (N_2510,In_108,In_830);
nand U2511 (N_2511,In_779,In_712);
nor U2512 (N_2512,In_903,In_68);
nand U2513 (N_2513,In_764,In_967);
nand U2514 (N_2514,In_98,In_183);
xor U2515 (N_2515,In_161,In_606);
or U2516 (N_2516,In_427,In_121);
nand U2517 (N_2517,In_355,In_7);
xor U2518 (N_2518,In_387,In_361);
nand U2519 (N_2519,In_315,In_141);
nand U2520 (N_2520,In_28,In_119);
or U2521 (N_2521,In_602,In_371);
or U2522 (N_2522,In_298,In_184);
nand U2523 (N_2523,In_566,In_189);
or U2524 (N_2524,In_386,In_232);
or U2525 (N_2525,In_239,In_536);
or U2526 (N_2526,In_655,In_13);
nand U2527 (N_2527,In_951,In_299);
nand U2528 (N_2528,In_562,In_80);
nor U2529 (N_2529,In_5,In_90);
xor U2530 (N_2530,In_674,In_739);
or U2531 (N_2531,In_673,In_516);
or U2532 (N_2532,In_916,In_41);
nor U2533 (N_2533,In_664,In_989);
xnor U2534 (N_2534,In_752,In_56);
xor U2535 (N_2535,In_428,In_202);
nor U2536 (N_2536,In_671,In_52);
and U2537 (N_2537,In_410,In_669);
or U2538 (N_2538,In_545,In_995);
nand U2539 (N_2539,In_308,In_382);
or U2540 (N_2540,In_399,In_914);
xnor U2541 (N_2541,In_466,In_368);
nand U2542 (N_2542,In_581,In_938);
and U2543 (N_2543,In_77,In_622);
xnor U2544 (N_2544,In_983,In_750);
nor U2545 (N_2545,In_327,In_133);
nor U2546 (N_2546,In_484,In_491);
nor U2547 (N_2547,In_165,In_306);
and U2548 (N_2548,In_619,In_830);
nor U2549 (N_2549,In_254,In_570);
nand U2550 (N_2550,In_399,In_278);
nor U2551 (N_2551,In_583,In_68);
nand U2552 (N_2552,In_523,In_912);
nand U2553 (N_2553,In_748,In_209);
nand U2554 (N_2554,In_309,In_512);
or U2555 (N_2555,In_308,In_896);
and U2556 (N_2556,In_14,In_755);
or U2557 (N_2557,In_959,In_707);
xor U2558 (N_2558,In_750,In_708);
nand U2559 (N_2559,In_646,In_302);
nand U2560 (N_2560,In_724,In_266);
xor U2561 (N_2561,In_350,In_664);
nor U2562 (N_2562,In_792,In_485);
and U2563 (N_2563,In_704,In_575);
and U2564 (N_2564,In_581,In_588);
nor U2565 (N_2565,In_58,In_234);
or U2566 (N_2566,In_69,In_950);
nor U2567 (N_2567,In_210,In_139);
nor U2568 (N_2568,In_7,In_715);
nor U2569 (N_2569,In_463,In_344);
nand U2570 (N_2570,In_939,In_635);
nand U2571 (N_2571,In_821,In_401);
or U2572 (N_2572,In_987,In_559);
and U2573 (N_2573,In_13,In_892);
or U2574 (N_2574,In_318,In_669);
xor U2575 (N_2575,In_942,In_640);
xnor U2576 (N_2576,In_200,In_970);
nor U2577 (N_2577,In_108,In_577);
and U2578 (N_2578,In_572,In_728);
xnor U2579 (N_2579,In_601,In_606);
and U2580 (N_2580,In_117,In_993);
xnor U2581 (N_2581,In_676,In_474);
or U2582 (N_2582,In_595,In_325);
nor U2583 (N_2583,In_871,In_877);
nor U2584 (N_2584,In_102,In_688);
nand U2585 (N_2585,In_575,In_251);
or U2586 (N_2586,In_728,In_752);
nand U2587 (N_2587,In_751,In_186);
or U2588 (N_2588,In_498,In_162);
xnor U2589 (N_2589,In_270,In_948);
xor U2590 (N_2590,In_949,In_30);
nor U2591 (N_2591,In_566,In_38);
nand U2592 (N_2592,In_724,In_834);
nor U2593 (N_2593,In_671,In_346);
and U2594 (N_2594,In_530,In_307);
xor U2595 (N_2595,In_895,In_398);
nand U2596 (N_2596,In_224,In_635);
nand U2597 (N_2597,In_577,In_687);
xnor U2598 (N_2598,In_138,In_358);
and U2599 (N_2599,In_42,In_645);
and U2600 (N_2600,In_987,In_464);
nor U2601 (N_2601,In_360,In_481);
nor U2602 (N_2602,In_461,In_143);
nor U2603 (N_2603,In_120,In_429);
nor U2604 (N_2604,In_814,In_77);
and U2605 (N_2605,In_27,In_718);
xnor U2606 (N_2606,In_232,In_255);
xnor U2607 (N_2607,In_15,In_388);
nor U2608 (N_2608,In_559,In_178);
xor U2609 (N_2609,In_696,In_686);
nor U2610 (N_2610,In_122,In_203);
nand U2611 (N_2611,In_767,In_51);
and U2612 (N_2612,In_655,In_49);
or U2613 (N_2613,In_344,In_900);
or U2614 (N_2614,In_121,In_60);
nor U2615 (N_2615,In_617,In_872);
nor U2616 (N_2616,In_132,In_492);
nand U2617 (N_2617,In_678,In_981);
or U2618 (N_2618,In_884,In_567);
xnor U2619 (N_2619,In_324,In_21);
nand U2620 (N_2620,In_301,In_851);
nand U2621 (N_2621,In_887,In_852);
and U2622 (N_2622,In_818,In_805);
xor U2623 (N_2623,In_652,In_11);
nor U2624 (N_2624,In_841,In_694);
xor U2625 (N_2625,In_926,In_691);
xnor U2626 (N_2626,In_750,In_953);
and U2627 (N_2627,In_584,In_434);
and U2628 (N_2628,In_716,In_719);
nand U2629 (N_2629,In_622,In_535);
nand U2630 (N_2630,In_169,In_524);
or U2631 (N_2631,In_998,In_62);
or U2632 (N_2632,In_797,In_11);
and U2633 (N_2633,In_71,In_29);
or U2634 (N_2634,In_987,In_749);
and U2635 (N_2635,In_971,In_15);
nor U2636 (N_2636,In_212,In_271);
nor U2637 (N_2637,In_414,In_199);
or U2638 (N_2638,In_976,In_371);
nand U2639 (N_2639,In_75,In_61);
nor U2640 (N_2640,In_586,In_726);
and U2641 (N_2641,In_582,In_531);
and U2642 (N_2642,In_810,In_360);
or U2643 (N_2643,In_350,In_574);
and U2644 (N_2644,In_2,In_715);
nor U2645 (N_2645,In_296,In_546);
nand U2646 (N_2646,In_13,In_501);
and U2647 (N_2647,In_927,In_605);
nor U2648 (N_2648,In_654,In_599);
or U2649 (N_2649,In_402,In_610);
and U2650 (N_2650,In_19,In_59);
xnor U2651 (N_2651,In_532,In_754);
nor U2652 (N_2652,In_370,In_614);
nor U2653 (N_2653,In_658,In_895);
nand U2654 (N_2654,In_32,In_299);
or U2655 (N_2655,In_669,In_522);
xor U2656 (N_2656,In_244,In_149);
and U2657 (N_2657,In_244,In_756);
or U2658 (N_2658,In_864,In_373);
and U2659 (N_2659,In_130,In_115);
and U2660 (N_2660,In_533,In_395);
xor U2661 (N_2661,In_305,In_810);
nor U2662 (N_2662,In_160,In_663);
xor U2663 (N_2663,In_909,In_69);
and U2664 (N_2664,In_8,In_128);
nand U2665 (N_2665,In_141,In_27);
nor U2666 (N_2666,In_2,In_649);
or U2667 (N_2667,In_314,In_915);
or U2668 (N_2668,In_374,In_591);
nor U2669 (N_2669,In_777,In_64);
nor U2670 (N_2670,In_419,In_44);
and U2671 (N_2671,In_344,In_695);
nand U2672 (N_2672,In_438,In_679);
xnor U2673 (N_2673,In_488,In_402);
and U2674 (N_2674,In_398,In_240);
nor U2675 (N_2675,In_17,In_649);
nor U2676 (N_2676,In_741,In_893);
nor U2677 (N_2677,In_868,In_70);
nand U2678 (N_2678,In_131,In_740);
nand U2679 (N_2679,In_832,In_992);
xnor U2680 (N_2680,In_60,In_33);
or U2681 (N_2681,In_917,In_943);
nor U2682 (N_2682,In_411,In_751);
nand U2683 (N_2683,In_586,In_107);
nor U2684 (N_2684,In_335,In_237);
or U2685 (N_2685,In_482,In_876);
xor U2686 (N_2686,In_766,In_24);
or U2687 (N_2687,In_594,In_200);
nand U2688 (N_2688,In_54,In_879);
or U2689 (N_2689,In_493,In_141);
nand U2690 (N_2690,In_384,In_403);
or U2691 (N_2691,In_362,In_964);
xor U2692 (N_2692,In_193,In_454);
or U2693 (N_2693,In_413,In_668);
or U2694 (N_2694,In_622,In_862);
and U2695 (N_2695,In_127,In_903);
nand U2696 (N_2696,In_923,In_726);
nand U2697 (N_2697,In_834,In_585);
nor U2698 (N_2698,In_600,In_142);
or U2699 (N_2699,In_405,In_289);
xor U2700 (N_2700,In_453,In_8);
xor U2701 (N_2701,In_377,In_672);
nand U2702 (N_2702,In_638,In_452);
or U2703 (N_2703,In_975,In_795);
nand U2704 (N_2704,In_392,In_431);
nor U2705 (N_2705,In_91,In_517);
nor U2706 (N_2706,In_192,In_641);
or U2707 (N_2707,In_12,In_94);
nand U2708 (N_2708,In_677,In_467);
nand U2709 (N_2709,In_895,In_792);
xor U2710 (N_2710,In_727,In_69);
or U2711 (N_2711,In_768,In_452);
nand U2712 (N_2712,In_885,In_275);
and U2713 (N_2713,In_16,In_191);
nor U2714 (N_2714,In_780,In_470);
nand U2715 (N_2715,In_857,In_431);
and U2716 (N_2716,In_341,In_931);
and U2717 (N_2717,In_42,In_183);
or U2718 (N_2718,In_873,In_241);
nand U2719 (N_2719,In_644,In_553);
or U2720 (N_2720,In_86,In_27);
and U2721 (N_2721,In_669,In_774);
nand U2722 (N_2722,In_814,In_256);
nand U2723 (N_2723,In_522,In_922);
nor U2724 (N_2724,In_850,In_157);
or U2725 (N_2725,In_687,In_694);
nor U2726 (N_2726,In_862,In_503);
and U2727 (N_2727,In_989,In_763);
nor U2728 (N_2728,In_963,In_744);
nand U2729 (N_2729,In_542,In_600);
and U2730 (N_2730,In_220,In_59);
nor U2731 (N_2731,In_756,In_790);
nor U2732 (N_2732,In_586,In_484);
or U2733 (N_2733,In_671,In_920);
xor U2734 (N_2734,In_595,In_30);
nor U2735 (N_2735,In_382,In_201);
or U2736 (N_2736,In_671,In_808);
and U2737 (N_2737,In_558,In_930);
nand U2738 (N_2738,In_755,In_254);
and U2739 (N_2739,In_358,In_558);
and U2740 (N_2740,In_722,In_658);
nand U2741 (N_2741,In_424,In_65);
and U2742 (N_2742,In_25,In_524);
xnor U2743 (N_2743,In_88,In_299);
nand U2744 (N_2744,In_571,In_948);
xor U2745 (N_2745,In_846,In_302);
xor U2746 (N_2746,In_472,In_982);
nand U2747 (N_2747,In_63,In_240);
nor U2748 (N_2748,In_922,In_949);
xnor U2749 (N_2749,In_376,In_93);
xor U2750 (N_2750,In_26,In_447);
and U2751 (N_2751,In_266,In_984);
and U2752 (N_2752,In_514,In_129);
nor U2753 (N_2753,In_911,In_684);
and U2754 (N_2754,In_114,In_115);
xnor U2755 (N_2755,In_134,In_720);
nand U2756 (N_2756,In_552,In_961);
nand U2757 (N_2757,In_766,In_250);
nor U2758 (N_2758,In_123,In_0);
and U2759 (N_2759,In_991,In_665);
xor U2760 (N_2760,In_408,In_138);
or U2761 (N_2761,In_66,In_2);
xor U2762 (N_2762,In_561,In_45);
and U2763 (N_2763,In_322,In_147);
and U2764 (N_2764,In_299,In_328);
nor U2765 (N_2765,In_897,In_294);
nand U2766 (N_2766,In_717,In_352);
nand U2767 (N_2767,In_926,In_818);
xor U2768 (N_2768,In_259,In_437);
and U2769 (N_2769,In_461,In_423);
nand U2770 (N_2770,In_718,In_842);
and U2771 (N_2771,In_329,In_906);
nand U2772 (N_2772,In_290,In_865);
xnor U2773 (N_2773,In_365,In_391);
xor U2774 (N_2774,In_896,In_242);
and U2775 (N_2775,In_905,In_314);
or U2776 (N_2776,In_437,In_807);
nor U2777 (N_2777,In_463,In_780);
xor U2778 (N_2778,In_868,In_686);
and U2779 (N_2779,In_966,In_72);
and U2780 (N_2780,In_697,In_254);
nor U2781 (N_2781,In_53,In_140);
nor U2782 (N_2782,In_734,In_182);
nand U2783 (N_2783,In_186,In_233);
and U2784 (N_2784,In_0,In_986);
nor U2785 (N_2785,In_110,In_896);
xnor U2786 (N_2786,In_652,In_836);
and U2787 (N_2787,In_27,In_638);
xnor U2788 (N_2788,In_673,In_518);
or U2789 (N_2789,In_917,In_168);
and U2790 (N_2790,In_438,In_610);
nor U2791 (N_2791,In_508,In_851);
and U2792 (N_2792,In_66,In_306);
and U2793 (N_2793,In_760,In_698);
nand U2794 (N_2794,In_702,In_957);
nand U2795 (N_2795,In_657,In_942);
and U2796 (N_2796,In_731,In_965);
xor U2797 (N_2797,In_8,In_36);
xnor U2798 (N_2798,In_465,In_296);
and U2799 (N_2799,In_695,In_437);
nand U2800 (N_2800,In_555,In_838);
nor U2801 (N_2801,In_817,In_109);
or U2802 (N_2802,In_816,In_77);
and U2803 (N_2803,In_697,In_351);
or U2804 (N_2804,In_731,In_745);
or U2805 (N_2805,In_719,In_325);
nor U2806 (N_2806,In_491,In_192);
xnor U2807 (N_2807,In_834,In_177);
and U2808 (N_2808,In_323,In_572);
nand U2809 (N_2809,In_682,In_74);
nor U2810 (N_2810,In_892,In_331);
xnor U2811 (N_2811,In_397,In_625);
or U2812 (N_2812,In_805,In_932);
nand U2813 (N_2813,In_290,In_252);
xor U2814 (N_2814,In_160,In_255);
nor U2815 (N_2815,In_544,In_293);
nor U2816 (N_2816,In_125,In_650);
nand U2817 (N_2817,In_844,In_380);
nor U2818 (N_2818,In_111,In_269);
xor U2819 (N_2819,In_271,In_837);
nand U2820 (N_2820,In_291,In_132);
nor U2821 (N_2821,In_860,In_747);
nand U2822 (N_2822,In_843,In_94);
or U2823 (N_2823,In_824,In_684);
nand U2824 (N_2824,In_427,In_649);
and U2825 (N_2825,In_803,In_842);
xor U2826 (N_2826,In_930,In_331);
and U2827 (N_2827,In_540,In_527);
nand U2828 (N_2828,In_197,In_890);
or U2829 (N_2829,In_597,In_864);
and U2830 (N_2830,In_923,In_783);
nand U2831 (N_2831,In_94,In_396);
or U2832 (N_2832,In_61,In_150);
xor U2833 (N_2833,In_227,In_149);
nor U2834 (N_2834,In_267,In_332);
xnor U2835 (N_2835,In_451,In_184);
or U2836 (N_2836,In_241,In_450);
nand U2837 (N_2837,In_810,In_661);
and U2838 (N_2838,In_588,In_47);
and U2839 (N_2839,In_953,In_859);
xor U2840 (N_2840,In_127,In_536);
and U2841 (N_2841,In_235,In_245);
nand U2842 (N_2842,In_848,In_995);
xnor U2843 (N_2843,In_691,In_503);
nor U2844 (N_2844,In_939,In_504);
nand U2845 (N_2845,In_594,In_71);
nand U2846 (N_2846,In_504,In_513);
xnor U2847 (N_2847,In_869,In_744);
xnor U2848 (N_2848,In_278,In_398);
nand U2849 (N_2849,In_379,In_327);
nor U2850 (N_2850,In_327,In_323);
or U2851 (N_2851,In_45,In_517);
xnor U2852 (N_2852,In_9,In_984);
nand U2853 (N_2853,In_763,In_829);
xor U2854 (N_2854,In_353,In_60);
xnor U2855 (N_2855,In_181,In_741);
or U2856 (N_2856,In_823,In_456);
or U2857 (N_2857,In_778,In_522);
or U2858 (N_2858,In_926,In_536);
nor U2859 (N_2859,In_527,In_308);
or U2860 (N_2860,In_243,In_901);
or U2861 (N_2861,In_532,In_179);
or U2862 (N_2862,In_709,In_492);
and U2863 (N_2863,In_239,In_213);
nand U2864 (N_2864,In_866,In_68);
and U2865 (N_2865,In_418,In_54);
xor U2866 (N_2866,In_188,In_459);
nand U2867 (N_2867,In_29,In_566);
nor U2868 (N_2868,In_545,In_739);
or U2869 (N_2869,In_118,In_426);
xnor U2870 (N_2870,In_791,In_733);
and U2871 (N_2871,In_358,In_681);
nand U2872 (N_2872,In_707,In_543);
nand U2873 (N_2873,In_237,In_244);
xor U2874 (N_2874,In_567,In_997);
or U2875 (N_2875,In_938,In_181);
or U2876 (N_2876,In_820,In_794);
nor U2877 (N_2877,In_39,In_724);
nor U2878 (N_2878,In_935,In_879);
or U2879 (N_2879,In_655,In_520);
nor U2880 (N_2880,In_109,In_694);
or U2881 (N_2881,In_467,In_385);
and U2882 (N_2882,In_69,In_665);
xnor U2883 (N_2883,In_509,In_938);
nor U2884 (N_2884,In_953,In_924);
nor U2885 (N_2885,In_9,In_138);
xor U2886 (N_2886,In_774,In_539);
or U2887 (N_2887,In_611,In_194);
nor U2888 (N_2888,In_495,In_286);
and U2889 (N_2889,In_227,In_28);
nor U2890 (N_2890,In_852,In_252);
nor U2891 (N_2891,In_846,In_851);
or U2892 (N_2892,In_937,In_762);
and U2893 (N_2893,In_785,In_827);
and U2894 (N_2894,In_764,In_324);
nor U2895 (N_2895,In_556,In_127);
nand U2896 (N_2896,In_76,In_392);
or U2897 (N_2897,In_13,In_813);
nor U2898 (N_2898,In_157,In_917);
nor U2899 (N_2899,In_273,In_891);
and U2900 (N_2900,In_914,In_69);
nor U2901 (N_2901,In_4,In_614);
xor U2902 (N_2902,In_396,In_354);
xnor U2903 (N_2903,In_742,In_572);
nand U2904 (N_2904,In_224,In_171);
nand U2905 (N_2905,In_998,In_359);
and U2906 (N_2906,In_39,In_114);
xnor U2907 (N_2907,In_269,In_824);
xor U2908 (N_2908,In_959,In_481);
and U2909 (N_2909,In_512,In_555);
nor U2910 (N_2910,In_912,In_476);
xor U2911 (N_2911,In_308,In_656);
nand U2912 (N_2912,In_310,In_802);
xor U2913 (N_2913,In_257,In_259);
or U2914 (N_2914,In_107,In_844);
and U2915 (N_2915,In_49,In_47);
or U2916 (N_2916,In_574,In_679);
nand U2917 (N_2917,In_571,In_986);
nand U2918 (N_2918,In_6,In_20);
xor U2919 (N_2919,In_185,In_936);
nor U2920 (N_2920,In_721,In_750);
or U2921 (N_2921,In_792,In_505);
or U2922 (N_2922,In_926,In_509);
nor U2923 (N_2923,In_928,In_137);
nand U2924 (N_2924,In_656,In_469);
nand U2925 (N_2925,In_68,In_868);
or U2926 (N_2926,In_465,In_265);
xor U2927 (N_2927,In_437,In_769);
nor U2928 (N_2928,In_630,In_106);
nand U2929 (N_2929,In_508,In_686);
nor U2930 (N_2930,In_86,In_898);
nor U2931 (N_2931,In_861,In_636);
nand U2932 (N_2932,In_58,In_743);
and U2933 (N_2933,In_71,In_640);
or U2934 (N_2934,In_933,In_588);
and U2935 (N_2935,In_500,In_314);
or U2936 (N_2936,In_518,In_903);
xnor U2937 (N_2937,In_361,In_814);
or U2938 (N_2938,In_689,In_682);
or U2939 (N_2939,In_212,In_708);
nand U2940 (N_2940,In_881,In_914);
nor U2941 (N_2941,In_305,In_225);
or U2942 (N_2942,In_874,In_877);
nand U2943 (N_2943,In_906,In_317);
nand U2944 (N_2944,In_624,In_729);
nand U2945 (N_2945,In_556,In_584);
xnor U2946 (N_2946,In_380,In_71);
nor U2947 (N_2947,In_808,In_381);
or U2948 (N_2948,In_11,In_699);
and U2949 (N_2949,In_364,In_660);
nor U2950 (N_2950,In_637,In_261);
and U2951 (N_2951,In_632,In_114);
xnor U2952 (N_2952,In_553,In_446);
and U2953 (N_2953,In_760,In_362);
and U2954 (N_2954,In_985,In_27);
nand U2955 (N_2955,In_145,In_758);
nand U2956 (N_2956,In_714,In_954);
or U2957 (N_2957,In_837,In_698);
and U2958 (N_2958,In_226,In_813);
or U2959 (N_2959,In_787,In_494);
or U2960 (N_2960,In_322,In_626);
and U2961 (N_2961,In_160,In_68);
nor U2962 (N_2962,In_288,In_222);
nand U2963 (N_2963,In_369,In_519);
or U2964 (N_2964,In_254,In_889);
nor U2965 (N_2965,In_39,In_879);
xnor U2966 (N_2966,In_862,In_642);
nor U2967 (N_2967,In_437,In_444);
nand U2968 (N_2968,In_366,In_500);
or U2969 (N_2969,In_237,In_268);
xor U2970 (N_2970,In_329,In_337);
nor U2971 (N_2971,In_520,In_298);
or U2972 (N_2972,In_52,In_351);
nand U2973 (N_2973,In_771,In_781);
and U2974 (N_2974,In_666,In_438);
xor U2975 (N_2975,In_124,In_549);
and U2976 (N_2976,In_169,In_862);
or U2977 (N_2977,In_484,In_797);
and U2978 (N_2978,In_183,In_259);
xor U2979 (N_2979,In_717,In_490);
nand U2980 (N_2980,In_157,In_617);
and U2981 (N_2981,In_380,In_913);
or U2982 (N_2982,In_807,In_678);
and U2983 (N_2983,In_787,In_536);
xor U2984 (N_2984,In_507,In_754);
xnor U2985 (N_2985,In_206,In_401);
or U2986 (N_2986,In_852,In_911);
nand U2987 (N_2987,In_44,In_78);
and U2988 (N_2988,In_724,In_570);
nor U2989 (N_2989,In_492,In_700);
nor U2990 (N_2990,In_697,In_12);
xor U2991 (N_2991,In_819,In_575);
and U2992 (N_2992,In_584,In_121);
xor U2993 (N_2993,In_173,In_973);
and U2994 (N_2994,In_442,In_872);
nor U2995 (N_2995,In_617,In_323);
nand U2996 (N_2996,In_603,In_916);
and U2997 (N_2997,In_678,In_626);
xnor U2998 (N_2998,In_320,In_593);
nor U2999 (N_2999,In_117,In_58);
nor U3000 (N_3000,In_410,In_77);
xor U3001 (N_3001,In_487,In_24);
or U3002 (N_3002,In_550,In_806);
and U3003 (N_3003,In_343,In_708);
nand U3004 (N_3004,In_908,In_833);
nor U3005 (N_3005,In_108,In_944);
nand U3006 (N_3006,In_489,In_120);
nor U3007 (N_3007,In_992,In_634);
xnor U3008 (N_3008,In_631,In_822);
xnor U3009 (N_3009,In_559,In_459);
and U3010 (N_3010,In_133,In_69);
or U3011 (N_3011,In_384,In_369);
or U3012 (N_3012,In_302,In_97);
nor U3013 (N_3013,In_405,In_377);
and U3014 (N_3014,In_574,In_915);
xor U3015 (N_3015,In_513,In_149);
or U3016 (N_3016,In_512,In_43);
or U3017 (N_3017,In_853,In_794);
and U3018 (N_3018,In_592,In_576);
and U3019 (N_3019,In_990,In_26);
and U3020 (N_3020,In_65,In_663);
and U3021 (N_3021,In_465,In_561);
xor U3022 (N_3022,In_47,In_636);
xor U3023 (N_3023,In_587,In_412);
and U3024 (N_3024,In_624,In_350);
and U3025 (N_3025,In_266,In_478);
nor U3026 (N_3026,In_270,In_495);
or U3027 (N_3027,In_500,In_778);
xnor U3028 (N_3028,In_954,In_930);
nand U3029 (N_3029,In_608,In_273);
or U3030 (N_3030,In_211,In_898);
nor U3031 (N_3031,In_369,In_766);
or U3032 (N_3032,In_247,In_282);
xnor U3033 (N_3033,In_168,In_210);
nand U3034 (N_3034,In_614,In_896);
nor U3035 (N_3035,In_682,In_212);
and U3036 (N_3036,In_735,In_276);
nand U3037 (N_3037,In_571,In_855);
nand U3038 (N_3038,In_565,In_709);
or U3039 (N_3039,In_850,In_568);
or U3040 (N_3040,In_87,In_285);
xnor U3041 (N_3041,In_815,In_643);
and U3042 (N_3042,In_509,In_448);
nand U3043 (N_3043,In_879,In_95);
nor U3044 (N_3044,In_734,In_61);
nand U3045 (N_3045,In_472,In_665);
nand U3046 (N_3046,In_694,In_331);
nor U3047 (N_3047,In_784,In_469);
xnor U3048 (N_3048,In_59,In_415);
xor U3049 (N_3049,In_976,In_63);
or U3050 (N_3050,In_15,In_357);
and U3051 (N_3051,In_535,In_44);
nand U3052 (N_3052,In_221,In_489);
nor U3053 (N_3053,In_639,In_355);
nand U3054 (N_3054,In_943,In_86);
nand U3055 (N_3055,In_945,In_208);
nand U3056 (N_3056,In_405,In_535);
xor U3057 (N_3057,In_876,In_216);
xnor U3058 (N_3058,In_489,In_360);
xor U3059 (N_3059,In_674,In_469);
xor U3060 (N_3060,In_565,In_823);
nand U3061 (N_3061,In_86,In_851);
and U3062 (N_3062,In_141,In_994);
or U3063 (N_3063,In_900,In_526);
or U3064 (N_3064,In_464,In_134);
and U3065 (N_3065,In_250,In_364);
nor U3066 (N_3066,In_972,In_145);
nor U3067 (N_3067,In_843,In_267);
or U3068 (N_3068,In_354,In_546);
or U3069 (N_3069,In_149,In_665);
nor U3070 (N_3070,In_964,In_342);
nand U3071 (N_3071,In_929,In_531);
or U3072 (N_3072,In_611,In_208);
xor U3073 (N_3073,In_427,In_650);
or U3074 (N_3074,In_382,In_598);
or U3075 (N_3075,In_444,In_999);
and U3076 (N_3076,In_89,In_504);
and U3077 (N_3077,In_310,In_483);
nand U3078 (N_3078,In_672,In_212);
nor U3079 (N_3079,In_482,In_270);
nor U3080 (N_3080,In_576,In_271);
and U3081 (N_3081,In_870,In_857);
xnor U3082 (N_3082,In_118,In_782);
or U3083 (N_3083,In_683,In_762);
nand U3084 (N_3084,In_739,In_450);
or U3085 (N_3085,In_3,In_56);
and U3086 (N_3086,In_209,In_515);
xnor U3087 (N_3087,In_259,In_517);
nand U3088 (N_3088,In_335,In_616);
nor U3089 (N_3089,In_827,In_349);
xnor U3090 (N_3090,In_865,In_25);
nand U3091 (N_3091,In_142,In_300);
and U3092 (N_3092,In_568,In_742);
nor U3093 (N_3093,In_32,In_182);
nand U3094 (N_3094,In_504,In_747);
or U3095 (N_3095,In_492,In_66);
nand U3096 (N_3096,In_405,In_502);
or U3097 (N_3097,In_736,In_640);
or U3098 (N_3098,In_361,In_233);
and U3099 (N_3099,In_74,In_659);
or U3100 (N_3100,In_472,In_301);
and U3101 (N_3101,In_472,In_928);
xnor U3102 (N_3102,In_147,In_202);
nor U3103 (N_3103,In_899,In_4);
or U3104 (N_3104,In_986,In_58);
nand U3105 (N_3105,In_967,In_719);
xnor U3106 (N_3106,In_227,In_386);
nand U3107 (N_3107,In_429,In_520);
nand U3108 (N_3108,In_237,In_998);
nand U3109 (N_3109,In_351,In_455);
or U3110 (N_3110,In_800,In_740);
xnor U3111 (N_3111,In_327,In_270);
xnor U3112 (N_3112,In_478,In_137);
nor U3113 (N_3113,In_745,In_76);
nor U3114 (N_3114,In_87,In_486);
xor U3115 (N_3115,In_673,In_911);
or U3116 (N_3116,In_798,In_729);
nor U3117 (N_3117,In_413,In_466);
nor U3118 (N_3118,In_633,In_116);
nand U3119 (N_3119,In_453,In_279);
and U3120 (N_3120,In_623,In_309);
nor U3121 (N_3121,In_150,In_136);
and U3122 (N_3122,In_368,In_445);
and U3123 (N_3123,In_387,In_924);
nand U3124 (N_3124,In_314,In_321);
xor U3125 (N_3125,In_432,In_901);
nand U3126 (N_3126,In_348,In_939);
and U3127 (N_3127,In_436,In_312);
or U3128 (N_3128,In_206,In_987);
nor U3129 (N_3129,In_649,In_626);
nor U3130 (N_3130,In_949,In_656);
xor U3131 (N_3131,In_23,In_8);
nor U3132 (N_3132,In_269,In_492);
nand U3133 (N_3133,In_631,In_995);
nor U3134 (N_3134,In_920,In_849);
nor U3135 (N_3135,In_536,In_232);
or U3136 (N_3136,In_404,In_159);
nand U3137 (N_3137,In_862,In_699);
nor U3138 (N_3138,In_569,In_384);
nor U3139 (N_3139,In_479,In_709);
xor U3140 (N_3140,In_191,In_615);
nand U3141 (N_3141,In_397,In_847);
nor U3142 (N_3142,In_113,In_161);
and U3143 (N_3143,In_231,In_387);
and U3144 (N_3144,In_478,In_558);
and U3145 (N_3145,In_679,In_392);
nand U3146 (N_3146,In_303,In_983);
nand U3147 (N_3147,In_774,In_61);
nor U3148 (N_3148,In_339,In_567);
and U3149 (N_3149,In_620,In_611);
nand U3150 (N_3150,In_796,In_221);
nor U3151 (N_3151,In_488,In_900);
xor U3152 (N_3152,In_335,In_808);
and U3153 (N_3153,In_301,In_348);
xnor U3154 (N_3154,In_677,In_555);
nand U3155 (N_3155,In_325,In_846);
nand U3156 (N_3156,In_148,In_24);
xor U3157 (N_3157,In_457,In_423);
xnor U3158 (N_3158,In_920,In_624);
nor U3159 (N_3159,In_730,In_195);
nand U3160 (N_3160,In_474,In_830);
nor U3161 (N_3161,In_43,In_433);
nor U3162 (N_3162,In_441,In_376);
and U3163 (N_3163,In_525,In_809);
xor U3164 (N_3164,In_297,In_867);
xnor U3165 (N_3165,In_369,In_242);
xor U3166 (N_3166,In_243,In_7);
and U3167 (N_3167,In_269,In_932);
xor U3168 (N_3168,In_751,In_938);
nor U3169 (N_3169,In_379,In_751);
xor U3170 (N_3170,In_478,In_79);
and U3171 (N_3171,In_732,In_83);
nor U3172 (N_3172,In_403,In_781);
or U3173 (N_3173,In_526,In_312);
nand U3174 (N_3174,In_795,In_193);
nor U3175 (N_3175,In_240,In_514);
nand U3176 (N_3176,In_677,In_705);
nor U3177 (N_3177,In_347,In_985);
nand U3178 (N_3178,In_106,In_76);
nand U3179 (N_3179,In_402,In_158);
nand U3180 (N_3180,In_527,In_94);
nand U3181 (N_3181,In_828,In_504);
nand U3182 (N_3182,In_965,In_390);
or U3183 (N_3183,In_217,In_513);
and U3184 (N_3184,In_469,In_84);
and U3185 (N_3185,In_227,In_762);
and U3186 (N_3186,In_163,In_269);
or U3187 (N_3187,In_835,In_268);
and U3188 (N_3188,In_867,In_108);
or U3189 (N_3189,In_989,In_94);
or U3190 (N_3190,In_757,In_652);
nor U3191 (N_3191,In_986,In_522);
and U3192 (N_3192,In_158,In_234);
nand U3193 (N_3193,In_637,In_408);
nor U3194 (N_3194,In_510,In_325);
nand U3195 (N_3195,In_79,In_11);
or U3196 (N_3196,In_261,In_566);
nand U3197 (N_3197,In_856,In_994);
nor U3198 (N_3198,In_334,In_912);
nor U3199 (N_3199,In_947,In_45);
xnor U3200 (N_3200,In_660,In_335);
nand U3201 (N_3201,In_907,In_291);
xor U3202 (N_3202,In_489,In_325);
nand U3203 (N_3203,In_790,In_62);
and U3204 (N_3204,In_210,In_542);
nand U3205 (N_3205,In_556,In_17);
nand U3206 (N_3206,In_400,In_774);
nand U3207 (N_3207,In_742,In_398);
xor U3208 (N_3208,In_115,In_290);
or U3209 (N_3209,In_151,In_853);
nor U3210 (N_3210,In_62,In_45);
and U3211 (N_3211,In_467,In_303);
and U3212 (N_3212,In_968,In_579);
nand U3213 (N_3213,In_289,In_613);
and U3214 (N_3214,In_210,In_518);
nand U3215 (N_3215,In_912,In_587);
and U3216 (N_3216,In_936,In_140);
nor U3217 (N_3217,In_353,In_711);
nand U3218 (N_3218,In_199,In_256);
xor U3219 (N_3219,In_947,In_778);
nor U3220 (N_3220,In_632,In_336);
nor U3221 (N_3221,In_417,In_72);
nand U3222 (N_3222,In_429,In_996);
or U3223 (N_3223,In_742,In_353);
nor U3224 (N_3224,In_451,In_200);
xor U3225 (N_3225,In_832,In_188);
nor U3226 (N_3226,In_98,In_426);
xor U3227 (N_3227,In_643,In_755);
nor U3228 (N_3228,In_842,In_465);
nor U3229 (N_3229,In_614,In_635);
or U3230 (N_3230,In_195,In_230);
xor U3231 (N_3231,In_702,In_798);
xnor U3232 (N_3232,In_330,In_691);
xnor U3233 (N_3233,In_50,In_960);
nand U3234 (N_3234,In_349,In_483);
xnor U3235 (N_3235,In_846,In_203);
and U3236 (N_3236,In_812,In_264);
nor U3237 (N_3237,In_649,In_231);
nor U3238 (N_3238,In_418,In_909);
nand U3239 (N_3239,In_234,In_517);
nand U3240 (N_3240,In_411,In_850);
nor U3241 (N_3241,In_895,In_209);
and U3242 (N_3242,In_258,In_47);
and U3243 (N_3243,In_728,In_401);
or U3244 (N_3244,In_303,In_999);
xnor U3245 (N_3245,In_181,In_400);
and U3246 (N_3246,In_499,In_855);
and U3247 (N_3247,In_343,In_622);
nor U3248 (N_3248,In_976,In_365);
xor U3249 (N_3249,In_799,In_4);
xor U3250 (N_3250,In_931,In_994);
xnor U3251 (N_3251,In_525,In_271);
and U3252 (N_3252,In_246,In_235);
and U3253 (N_3253,In_333,In_428);
nor U3254 (N_3254,In_989,In_210);
nor U3255 (N_3255,In_519,In_924);
xor U3256 (N_3256,In_381,In_341);
or U3257 (N_3257,In_436,In_759);
xnor U3258 (N_3258,In_198,In_306);
and U3259 (N_3259,In_115,In_621);
xor U3260 (N_3260,In_21,In_74);
or U3261 (N_3261,In_439,In_178);
nand U3262 (N_3262,In_212,In_889);
or U3263 (N_3263,In_703,In_303);
or U3264 (N_3264,In_25,In_552);
nor U3265 (N_3265,In_12,In_47);
xnor U3266 (N_3266,In_777,In_822);
nand U3267 (N_3267,In_889,In_337);
or U3268 (N_3268,In_882,In_8);
or U3269 (N_3269,In_807,In_277);
and U3270 (N_3270,In_532,In_871);
nor U3271 (N_3271,In_170,In_731);
xor U3272 (N_3272,In_962,In_807);
xnor U3273 (N_3273,In_50,In_155);
or U3274 (N_3274,In_721,In_547);
or U3275 (N_3275,In_915,In_175);
or U3276 (N_3276,In_723,In_734);
nand U3277 (N_3277,In_465,In_638);
nor U3278 (N_3278,In_62,In_684);
and U3279 (N_3279,In_443,In_902);
nor U3280 (N_3280,In_737,In_783);
or U3281 (N_3281,In_771,In_955);
nor U3282 (N_3282,In_907,In_495);
and U3283 (N_3283,In_830,In_917);
or U3284 (N_3284,In_373,In_195);
xnor U3285 (N_3285,In_837,In_517);
nand U3286 (N_3286,In_951,In_882);
nand U3287 (N_3287,In_75,In_682);
or U3288 (N_3288,In_554,In_327);
nor U3289 (N_3289,In_475,In_8);
and U3290 (N_3290,In_707,In_391);
nand U3291 (N_3291,In_344,In_430);
or U3292 (N_3292,In_581,In_372);
nand U3293 (N_3293,In_467,In_344);
nand U3294 (N_3294,In_250,In_753);
nor U3295 (N_3295,In_852,In_436);
and U3296 (N_3296,In_860,In_731);
xnor U3297 (N_3297,In_225,In_371);
or U3298 (N_3298,In_339,In_28);
nand U3299 (N_3299,In_550,In_454);
or U3300 (N_3300,In_859,In_5);
nand U3301 (N_3301,In_158,In_963);
xnor U3302 (N_3302,In_670,In_503);
nand U3303 (N_3303,In_965,In_907);
or U3304 (N_3304,In_658,In_697);
xor U3305 (N_3305,In_61,In_645);
nand U3306 (N_3306,In_11,In_90);
xor U3307 (N_3307,In_723,In_550);
nor U3308 (N_3308,In_873,In_233);
or U3309 (N_3309,In_551,In_541);
or U3310 (N_3310,In_930,In_207);
xnor U3311 (N_3311,In_514,In_517);
nand U3312 (N_3312,In_790,In_723);
or U3313 (N_3313,In_699,In_465);
nand U3314 (N_3314,In_674,In_106);
nor U3315 (N_3315,In_381,In_544);
xor U3316 (N_3316,In_990,In_302);
nor U3317 (N_3317,In_896,In_208);
xor U3318 (N_3318,In_834,In_831);
nand U3319 (N_3319,In_697,In_727);
xnor U3320 (N_3320,In_553,In_777);
xor U3321 (N_3321,In_846,In_789);
or U3322 (N_3322,In_838,In_330);
or U3323 (N_3323,In_193,In_420);
nor U3324 (N_3324,In_953,In_21);
or U3325 (N_3325,In_327,In_965);
and U3326 (N_3326,In_745,In_106);
or U3327 (N_3327,In_675,In_865);
and U3328 (N_3328,In_984,In_886);
and U3329 (N_3329,In_1,In_947);
and U3330 (N_3330,In_740,In_334);
and U3331 (N_3331,In_70,In_989);
xor U3332 (N_3332,In_392,In_208);
nor U3333 (N_3333,In_767,In_498);
and U3334 (N_3334,In_19,In_155);
nand U3335 (N_3335,In_128,In_955);
nor U3336 (N_3336,In_420,In_104);
or U3337 (N_3337,In_84,In_907);
and U3338 (N_3338,In_133,In_142);
and U3339 (N_3339,In_832,In_408);
and U3340 (N_3340,In_835,In_766);
nand U3341 (N_3341,In_981,In_995);
nor U3342 (N_3342,In_633,In_701);
xor U3343 (N_3343,In_119,In_11);
or U3344 (N_3344,In_858,In_302);
and U3345 (N_3345,In_85,In_803);
or U3346 (N_3346,In_372,In_723);
or U3347 (N_3347,In_784,In_795);
or U3348 (N_3348,In_87,In_879);
and U3349 (N_3349,In_768,In_634);
nor U3350 (N_3350,In_142,In_824);
nand U3351 (N_3351,In_16,In_48);
xnor U3352 (N_3352,In_424,In_834);
and U3353 (N_3353,In_474,In_623);
or U3354 (N_3354,In_693,In_106);
or U3355 (N_3355,In_425,In_893);
and U3356 (N_3356,In_156,In_903);
nor U3357 (N_3357,In_467,In_124);
or U3358 (N_3358,In_403,In_116);
nand U3359 (N_3359,In_567,In_553);
nor U3360 (N_3360,In_544,In_150);
xnor U3361 (N_3361,In_269,In_462);
and U3362 (N_3362,In_68,In_766);
or U3363 (N_3363,In_388,In_488);
xor U3364 (N_3364,In_777,In_701);
nor U3365 (N_3365,In_171,In_122);
nand U3366 (N_3366,In_139,In_217);
nand U3367 (N_3367,In_236,In_421);
nand U3368 (N_3368,In_619,In_678);
nand U3369 (N_3369,In_693,In_846);
or U3370 (N_3370,In_354,In_826);
nor U3371 (N_3371,In_991,In_497);
nor U3372 (N_3372,In_121,In_662);
xnor U3373 (N_3373,In_326,In_712);
or U3374 (N_3374,In_912,In_520);
xnor U3375 (N_3375,In_413,In_504);
or U3376 (N_3376,In_809,In_903);
xor U3377 (N_3377,In_245,In_669);
or U3378 (N_3378,In_73,In_247);
xor U3379 (N_3379,In_973,In_676);
and U3380 (N_3380,In_733,In_706);
and U3381 (N_3381,In_890,In_420);
xnor U3382 (N_3382,In_258,In_186);
nor U3383 (N_3383,In_404,In_952);
xor U3384 (N_3384,In_751,In_52);
nor U3385 (N_3385,In_489,In_179);
and U3386 (N_3386,In_517,In_96);
and U3387 (N_3387,In_339,In_369);
xor U3388 (N_3388,In_377,In_783);
nand U3389 (N_3389,In_623,In_711);
nor U3390 (N_3390,In_5,In_695);
or U3391 (N_3391,In_271,In_418);
and U3392 (N_3392,In_178,In_95);
xnor U3393 (N_3393,In_698,In_542);
nor U3394 (N_3394,In_279,In_481);
xnor U3395 (N_3395,In_556,In_196);
nand U3396 (N_3396,In_147,In_268);
nor U3397 (N_3397,In_149,In_23);
nor U3398 (N_3398,In_980,In_363);
nand U3399 (N_3399,In_869,In_678);
and U3400 (N_3400,In_588,In_752);
nand U3401 (N_3401,In_107,In_862);
and U3402 (N_3402,In_620,In_834);
nand U3403 (N_3403,In_125,In_644);
and U3404 (N_3404,In_51,In_25);
nand U3405 (N_3405,In_367,In_956);
xor U3406 (N_3406,In_877,In_920);
and U3407 (N_3407,In_961,In_871);
nor U3408 (N_3408,In_152,In_994);
and U3409 (N_3409,In_273,In_93);
nor U3410 (N_3410,In_642,In_86);
or U3411 (N_3411,In_92,In_144);
and U3412 (N_3412,In_851,In_631);
and U3413 (N_3413,In_235,In_255);
nor U3414 (N_3414,In_283,In_529);
nor U3415 (N_3415,In_190,In_638);
xor U3416 (N_3416,In_448,In_585);
nor U3417 (N_3417,In_130,In_213);
nand U3418 (N_3418,In_91,In_55);
nor U3419 (N_3419,In_100,In_332);
xnor U3420 (N_3420,In_416,In_417);
nor U3421 (N_3421,In_841,In_117);
or U3422 (N_3422,In_850,In_563);
or U3423 (N_3423,In_477,In_407);
or U3424 (N_3424,In_318,In_748);
nand U3425 (N_3425,In_387,In_340);
nand U3426 (N_3426,In_689,In_107);
nand U3427 (N_3427,In_124,In_226);
and U3428 (N_3428,In_659,In_277);
nor U3429 (N_3429,In_103,In_384);
nand U3430 (N_3430,In_223,In_414);
nor U3431 (N_3431,In_839,In_117);
or U3432 (N_3432,In_551,In_660);
and U3433 (N_3433,In_14,In_226);
nor U3434 (N_3434,In_144,In_858);
nand U3435 (N_3435,In_787,In_316);
and U3436 (N_3436,In_79,In_238);
and U3437 (N_3437,In_866,In_302);
xnor U3438 (N_3438,In_163,In_489);
xnor U3439 (N_3439,In_876,In_19);
nor U3440 (N_3440,In_215,In_395);
nor U3441 (N_3441,In_647,In_573);
or U3442 (N_3442,In_510,In_575);
nor U3443 (N_3443,In_933,In_370);
and U3444 (N_3444,In_311,In_216);
or U3445 (N_3445,In_924,In_280);
or U3446 (N_3446,In_845,In_12);
nor U3447 (N_3447,In_601,In_497);
nor U3448 (N_3448,In_33,In_439);
xor U3449 (N_3449,In_284,In_640);
nor U3450 (N_3450,In_641,In_293);
nand U3451 (N_3451,In_735,In_694);
or U3452 (N_3452,In_297,In_170);
nand U3453 (N_3453,In_623,In_275);
xnor U3454 (N_3454,In_572,In_42);
or U3455 (N_3455,In_302,In_710);
xnor U3456 (N_3456,In_48,In_61);
or U3457 (N_3457,In_288,In_342);
nand U3458 (N_3458,In_655,In_870);
nand U3459 (N_3459,In_247,In_418);
and U3460 (N_3460,In_453,In_290);
nor U3461 (N_3461,In_599,In_139);
or U3462 (N_3462,In_629,In_363);
xor U3463 (N_3463,In_596,In_334);
or U3464 (N_3464,In_726,In_248);
xnor U3465 (N_3465,In_473,In_712);
nand U3466 (N_3466,In_42,In_802);
nor U3467 (N_3467,In_384,In_326);
nor U3468 (N_3468,In_956,In_735);
nor U3469 (N_3469,In_886,In_567);
and U3470 (N_3470,In_896,In_366);
or U3471 (N_3471,In_430,In_911);
and U3472 (N_3472,In_884,In_714);
nand U3473 (N_3473,In_554,In_372);
nand U3474 (N_3474,In_516,In_745);
and U3475 (N_3475,In_878,In_775);
nor U3476 (N_3476,In_829,In_801);
or U3477 (N_3477,In_79,In_245);
or U3478 (N_3478,In_63,In_761);
or U3479 (N_3479,In_681,In_296);
nor U3480 (N_3480,In_342,In_831);
and U3481 (N_3481,In_966,In_254);
and U3482 (N_3482,In_743,In_699);
xnor U3483 (N_3483,In_536,In_235);
or U3484 (N_3484,In_608,In_640);
xnor U3485 (N_3485,In_436,In_143);
xor U3486 (N_3486,In_933,In_454);
nor U3487 (N_3487,In_414,In_562);
nand U3488 (N_3488,In_53,In_28);
or U3489 (N_3489,In_628,In_454);
nand U3490 (N_3490,In_739,In_981);
or U3491 (N_3491,In_995,In_844);
or U3492 (N_3492,In_153,In_266);
or U3493 (N_3493,In_130,In_224);
xnor U3494 (N_3494,In_918,In_439);
xnor U3495 (N_3495,In_729,In_342);
and U3496 (N_3496,In_748,In_801);
nor U3497 (N_3497,In_842,In_827);
nand U3498 (N_3498,In_687,In_440);
xor U3499 (N_3499,In_315,In_72);
xor U3500 (N_3500,In_5,In_349);
nand U3501 (N_3501,In_931,In_933);
nor U3502 (N_3502,In_306,In_797);
xnor U3503 (N_3503,In_167,In_434);
nor U3504 (N_3504,In_368,In_126);
nand U3505 (N_3505,In_906,In_587);
or U3506 (N_3506,In_52,In_277);
and U3507 (N_3507,In_143,In_134);
or U3508 (N_3508,In_254,In_711);
nor U3509 (N_3509,In_705,In_272);
and U3510 (N_3510,In_912,In_778);
or U3511 (N_3511,In_316,In_940);
nor U3512 (N_3512,In_141,In_318);
xnor U3513 (N_3513,In_535,In_668);
and U3514 (N_3514,In_375,In_355);
or U3515 (N_3515,In_269,In_899);
nand U3516 (N_3516,In_680,In_575);
or U3517 (N_3517,In_990,In_185);
xnor U3518 (N_3518,In_407,In_525);
or U3519 (N_3519,In_493,In_178);
nand U3520 (N_3520,In_270,In_740);
xor U3521 (N_3521,In_996,In_307);
xor U3522 (N_3522,In_619,In_553);
xor U3523 (N_3523,In_117,In_145);
nor U3524 (N_3524,In_48,In_856);
nand U3525 (N_3525,In_508,In_874);
and U3526 (N_3526,In_215,In_712);
nand U3527 (N_3527,In_970,In_739);
nor U3528 (N_3528,In_853,In_781);
xnor U3529 (N_3529,In_72,In_166);
xnor U3530 (N_3530,In_905,In_515);
and U3531 (N_3531,In_533,In_161);
nand U3532 (N_3532,In_984,In_114);
xor U3533 (N_3533,In_609,In_107);
or U3534 (N_3534,In_264,In_353);
or U3535 (N_3535,In_132,In_714);
nand U3536 (N_3536,In_409,In_933);
xnor U3537 (N_3537,In_30,In_589);
nand U3538 (N_3538,In_868,In_717);
nand U3539 (N_3539,In_386,In_721);
or U3540 (N_3540,In_937,In_174);
nor U3541 (N_3541,In_324,In_773);
nor U3542 (N_3542,In_850,In_970);
nor U3543 (N_3543,In_24,In_802);
nor U3544 (N_3544,In_567,In_672);
nand U3545 (N_3545,In_554,In_212);
nand U3546 (N_3546,In_143,In_481);
and U3547 (N_3547,In_714,In_293);
nor U3548 (N_3548,In_349,In_735);
or U3549 (N_3549,In_61,In_80);
or U3550 (N_3550,In_680,In_160);
and U3551 (N_3551,In_877,In_984);
and U3552 (N_3552,In_187,In_788);
and U3553 (N_3553,In_648,In_452);
nand U3554 (N_3554,In_641,In_258);
xnor U3555 (N_3555,In_842,In_698);
nand U3556 (N_3556,In_380,In_388);
and U3557 (N_3557,In_73,In_981);
nand U3558 (N_3558,In_820,In_489);
xor U3559 (N_3559,In_730,In_845);
nor U3560 (N_3560,In_90,In_625);
and U3561 (N_3561,In_398,In_336);
and U3562 (N_3562,In_913,In_631);
nand U3563 (N_3563,In_109,In_538);
or U3564 (N_3564,In_882,In_579);
nand U3565 (N_3565,In_846,In_858);
nor U3566 (N_3566,In_212,In_410);
nand U3567 (N_3567,In_392,In_187);
or U3568 (N_3568,In_43,In_565);
nand U3569 (N_3569,In_898,In_427);
or U3570 (N_3570,In_283,In_970);
nor U3571 (N_3571,In_301,In_471);
and U3572 (N_3572,In_382,In_523);
or U3573 (N_3573,In_37,In_533);
or U3574 (N_3574,In_45,In_351);
and U3575 (N_3575,In_421,In_127);
xor U3576 (N_3576,In_643,In_285);
xnor U3577 (N_3577,In_914,In_129);
nand U3578 (N_3578,In_601,In_847);
nor U3579 (N_3579,In_724,In_689);
nand U3580 (N_3580,In_413,In_330);
nand U3581 (N_3581,In_142,In_50);
or U3582 (N_3582,In_29,In_735);
nor U3583 (N_3583,In_468,In_230);
xnor U3584 (N_3584,In_443,In_714);
nor U3585 (N_3585,In_967,In_547);
nand U3586 (N_3586,In_270,In_252);
nand U3587 (N_3587,In_249,In_418);
nand U3588 (N_3588,In_84,In_935);
or U3589 (N_3589,In_429,In_492);
or U3590 (N_3590,In_107,In_454);
nor U3591 (N_3591,In_717,In_492);
or U3592 (N_3592,In_919,In_949);
and U3593 (N_3593,In_81,In_472);
nand U3594 (N_3594,In_482,In_412);
or U3595 (N_3595,In_812,In_37);
or U3596 (N_3596,In_41,In_70);
or U3597 (N_3597,In_365,In_522);
and U3598 (N_3598,In_630,In_154);
nand U3599 (N_3599,In_203,In_216);
and U3600 (N_3600,In_35,In_542);
nor U3601 (N_3601,In_896,In_288);
or U3602 (N_3602,In_253,In_289);
or U3603 (N_3603,In_145,In_69);
nand U3604 (N_3604,In_753,In_431);
and U3605 (N_3605,In_193,In_470);
and U3606 (N_3606,In_987,In_340);
and U3607 (N_3607,In_889,In_164);
nand U3608 (N_3608,In_991,In_363);
and U3609 (N_3609,In_102,In_61);
xnor U3610 (N_3610,In_289,In_562);
nand U3611 (N_3611,In_266,In_325);
nor U3612 (N_3612,In_121,In_638);
and U3613 (N_3613,In_461,In_984);
and U3614 (N_3614,In_956,In_603);
nor U3615 (N_3615,In_713,In_554);
or U3616 (N_3616,In_629,In_369);
or U3617 (N_3617,In_79,In_534);
nor U3618 (N_3618,In_655,In_12);
nor U3619 (N_3619,In_358,In_326);
or U3620 (N_3620,In_955,In_916);
nand U3621 (N_3621,In_691,In_811);
and U3622 (N_3622,In_275,In_706);
nand U3623 (N_3623,In_371,In_744);
and U3624 (N_3624,In_113,In_998);
xnor U3625 (N_3625,In_825,In_114);
nand U3626 (N_3626,In_880,In_87);
nor U3627 (N_3627,In_203,In_897);
nor U3628 (N_3628,In_132,In_447);
nand U3629 (N_3629,In_738,In_556);
and U3630 (N_3630,In_70,In_563);
xor U3631 (N_3631,In_876,In_126);
nand U3632 (N_3632,In_989,In_756);
or U3633 (N_3633,In_152,In_163);
nor U3634 (N_3634,In_178,In_435);
nand U3635 (N_3635,In_774,In_391);
and U3636 (N_3636,In_824,In_994);
or U3637 (N_3637,In_376,In_617);
or U3638 (N_3638,In_415,In_446);
nor U3639 (N_3639,In_210,In_465);
or U3640 (N_3640,In_510,In_778);
nand U3641 (N_3641,In_682,In_939);
or U3642 (N_3642,In_598,In_517);
nor U3643 (N_3643,In_973,In_171);
nor U3644 (N_3644,In_896,In_383);
nand U3645 (N_3645,In_733,In_206);
nand U3646 (N_3646,In_250,In_909);
or U3647 (N_3647,In_456,In_383);
xor U3648 (N_3648,In_639,In_778);
nor U3649 (N_3649,In_722,In_798);
nand U3650 (N_3650,In_611,In_279);
nand U3651 (N_3651,In_608,In_220);
and U3652 (N_3652,In_176,In_833);
and U3653 (N_3653,In_614,In_556);
xor U3654 (N_3654,In_708,In_43);
or U3655 (N_3655,In_700,In_45);
and U3656 (N_3656,In_280,In_434);
or U3657 (N_3657,In_612,In_191);
nand U3658 (N_3658,In_216,In_235);
and U3659 (N_3659,In_968,In_674);
and U3660 (N_3660,In_802,In_723);
xor U3661 (N_3661,In_303,In_214);
xnor U3662 (N_3662,In_522,In_19);
or U3663 (N_3663,In_911,In_751);
and U3664 (N_3664,In_130,In_339);
xor U3665 (N_3665,In_104,In_375);
and U3666 (N_3666,In_585,In_369);
and U3667 (N_3667,In_550,In_134);
nand U3668 (N_3668,In_786,In_732);
nand U3669 (N_3669,In_404,In_649);
or U3670 (N_3670,In_16,In_382);
or U3671 (N_3671,In_195,In_827);
or U3672 (N_3672,In_229,In_11);
or U3673 (N_3673,In_711,In_835);
or U3674 (N_3674,In_743,In_939);
nand U3675 (N_3675,In_115,In_479);
nand U3676 (N_3676,In_777,In_595);
and U3677 (N_3677,In_904,In_132);
xor U3678 (N_3678,In_957,In_648);
and U3679 (N_3679,In_620,In_49);
xor U3680 (N_3680,In_625,In_353);
nor U3681 (N_3681,In_436,In_415);
and U3682 (N_3682,In_691,In_218);
and U3683 (N_3683,In_319,In_644);
nor U3684 (N_3684,In_629,In_473);
nand U3685 (N_3685,In_120,In_185);
xnor U3686 (N_3686,In_252,In_239);
and U3687 (N_3687,In_166,In_730);
xnor U3688 (N_3688,In_523,In_886);
or U3689 (N_3689,In_246,In_884);
nor U3690 (N_3690,In_747,In_603);
nor U3691 (N_3691,In_731,In_864);
and U3692 (N_3692,In_165,In_519);
xor U3693 (N_3693,In_215,In_602);
or U3694 (N_3694,In_933,In_399);
and U3695 (N_3695,In_26,In_726);
xnor U3696 (N_3696,In_61,In_174);
xnor U3697 (N_3697,In_748,In_847);
nor U3698 (N_3698,In_935,In_292);
nor U3699 (N_3699,In_582,In_375);
xor U3700 (N_3700,In_559,In_954);
nand U3701 (N_3701,In_407,In_48);
nor U3702 (N_3702,In_565,In_179);
and U3703 (N_3703,In_766,In_271);
nand U3704 (N_3704,In_685,In_783);
xnor U3705 (N_3705,In_464,In_423);
nor U3706 (N_3706,In_65,In_641);
xnor U3707 (N_3707,In_919,In_206);
and U3708 (N_3708,In_956,In_65);
and U3709 (N_3709,In_245,In_862);
xnor U3710 (N_3710,In_114,In_566);
or U3711 (N_3711,In_925,In_794);
and U3712 (N_3712,In_122,In_380);
and U3713 (N_3713,In_532,In_83);
or U3714 (N_3714,In_18,In_817);
or U3715 (N_3715,In_434,In_549);
nor U3716 (N_3716,In_690,In_994);
nor U3717 (N_3717,In_666,In_227);
or U3718 (N_3718,In_475,In_282);
nand U3719 (N_3719,In_907,In_662);
nor U3720 (N_3720,In_926,In_408);
nor U3721 (N_3721,In_210,In_998);
xnor U3722 (N_3722,In_444,In_889);
xor U3723 (N_3723,In_376,In_578);
or U3724 (N_3724,In_793,In_943);
and U3725 (N_3725,In_894,In_448);
and U3726 (N_3726,In_272,In_241);
or U3727 (N_3727,In_488,In_78);
or U3728 (N_3728,In_81,In_718);
nor U3729 (N_3729,In_727,In_594);
nor U3730 (N_3730,In_593,In_317);
nand U3731 (N_3731,In_211,In_220);
and U3732 (N_3732,In_512,In_334);
or U3733 (N_3733,In_5,In_538);
or U3734 (N_3734,In_367,In_635);
nor U3735 (N_3735,In_850,In_105);
xor U3736 (N_3736,In_709,In_403);
xor U3737 (N_3737,In_972,In_791);
xor U3738 (N_3738,In_663,In_973);
nor U3739 (N_3739,In_920,In_205);
and U3740 (N_3740,In_722,In_183);
or U3741 (N_3741,In_977,In_184);
xor U3742 (N_3742,In_674,In_484);
nand U3743 (N_3743,In_146,In_568);
nor U3744 (N_3744,In_215,In_989);
nor U3745 (N_3745,In_651,In_369);
nand U3746 (N_3746,In_953,In_837);
nand U3747 (N_3747,In_51,In_294);
and U3748 (N_3748,In_437,In_777);
nand U3749 (N_3749,In_539,In_596);
or U3750 (N_3750,In_327,In_997);
nand U3751 (N_3751,In_99,In_859);
and U3752 (N_3752,In_98,In_62);
or U3753 (N_3753,In_262,In_959);
nor U3754 (N_3754,In_667,In_690);
xnor U3755 (N_3755,In_277,In_912);
or U3756 (N_3756,In_920,In_729);
nand U3757 (N_3757,In_596,In_736);
or U3758 (N_3758,In_844,In_667);
and U3759 (N_3759,In_972,In_366);
or U3760 (N_3760,In_753,In_379);
and U3761 (N_3761,In_806,In_440);
nor U3762 (N_3762,In_379,In_691);
nand U3763 (N_3763,In_941,In_397);
xnor U3764 (N_3764,In_95,In_731);
and U3765 (N_3765,In_474,In_15);
nand U3766 (N_3766,In_883,In_68);
nor U3767 (N_3767,In_792,In_297);
nand U3768 (N_3768,In_773,In_206);
nand U3769 (N_3769,In_550,In_380);
nor U3770 (N_3770,In_791,In_754);
nand U3771 (N_3771,In_127,In_965);
nand U3772 (N_3772,In_644,In_234);
xnor U3773 (N_3773,In_734,In_290);
nor U3774 (N_3774,In_695,In_58);
nand U3775 (N_3775,In_745,In_101);
nand U3776 (N_3776,In_966,In_556);
and U3777 (N_3777,In_316,In_774);
nand U3778 (N_3778,In_341,In_84);
xnor U3779 (N_3779,In_196,In_648);
or U3780 (N_3780,In_829,In_24);
nor U3781 (N_3781,In_947,In_177);
nor U3782 (N_3782,In_731,In_650);
and U3783 (N_3783,In_498,In_16);
or U3784 (N_3784,In_177,In_535);
nand U3785 (N_3785,In_845,In_84);
or U3786 (N_3786,In_96,In_746);
nand U3787 (N_3787,In_110,In_763);
and U3788 (N_3788,In_949,In_275);
nor U3789 (N_3789,In_488,In_976);
and U3790 (N_3790,In_142,In_234);
or U3791 (N_3791,In_340,In_744);
and U3792 (N_3792,In_770,In_356);
nor U3793 (N_3793,In_963,In_429);
or U3794 (N_3794,In_246,In_91);
xnor U3795 (N_3795,In_583,In_750);
and U3796 (N_3796,In_119,In_913);
nor U3797 (N_3797,In_128,In_479);
and U3798 (N_3798,In_587,In_33);
xnor U3799 (N_3799,In_312,In_592);
or U3800 (N_3800,In_44,In_451);
nand U3801 (N_3801,In_80,In_772);
nand U3802 (N_3802,In_677,In_152);
nand U3803 (N_3803,In_468,In_113);
nor U3804 (N_3804,In_329,In_984);
and U3805 (N_3805,In_937,In_293);
nand U3806 (N_3806,In_101,In_250);
or U3807 (N_3807,In_989,In_765);
and U3808 (N_3808,In_682,In_226);
xnor U3809 (N_3809,In_810,In_198);
and U3810 (N_3810,In_51,In_272);
nand U3811 (N_3811,In_977,In_213);
xnor U3812 (N_3812,In_710,In_216);
or U3813 (N_3813,In_476,In_199);
nor U3814 (N_3814,In_939,In_731);
and U3815 (N_3815,In_45,In_177);
xnor U3816 (N_3816,In_688,In_562);
nand U3817 (N_3817,In_756,In_380);
or U3818 (N_3818,In_676,In_966);
xor U3819 (N_3819,In_222,In_240);
or U3820 (N_3820,In_226,In_826);
or U3821 (N_3821,In_653,In_826);
and U3822 (N_3822,In_147,In_410);
nor U3823 (N_3823,In_735,In_272);
nor U3824 (N_3824,In_425,In_82);
or U3825 (N_3825,In_822,In_406);
xnor U3826 (N_3826,In_41,In_929);
or U3827 (N_3827,In_526,In_74);
and U3828 (N_3828,In_200,In_924);
and U3829 (N_3829,In_275,In_803);
or U3830 (N_3830,In_871,In_353);
xnor U3831 (N_3831,In_674,In_147);
nand U3832 (N_3832,In_569,In_904);
or U3833 (N_3833,In_797,In_850);
nand U3834 (N_3834,In_353,In_381);
xor U3835 (N_3835,In_821,In_545);
or U3836 (N_3836,In_630,In_657);
xor U3837 (N_3837,In_503,In_390);
nand U3838 (N_3838,In_125,In_964);
and U3839 (N_3839,In_837,In_606);
nor U3840 (N_3840,In_133,In_686);
and U3841 (N_3841,In_988,In_115);
and U3842 (N_3842,In_26,In_865);
xor U3843 (N_3843,In_498,In_436);
or U3844 (N_3844,In_809,In_104);
xor U3845 (N_3845,In_616,In_946);
and U3846 (N_3846,In_501,In_573);
nand U3847 (N_3847,In_629,In_92);
xnor U3848 (N_3848,In_654,In_911);
and U3849 (N_3849,In_338,In_100);
and U3850 (N_3850,In_5,In_916);
nor U3851 (N_3851,In_581,In_416);
or U3852 (N_3852,In_443,In_158);
or U3853 (N_3853,In_373,In_39);
nand U3854 (N_3854,In_462,In_373);
or U3855 (N_3855,In_751,In_381);
xor U3856 (N_3856,In_842,In_216);
and U3857 (N_3857,In_11,In_555);
xnor U3858 (N_3858,In_667,In_191);
nor U3859 (N_3859,In_96,In_956);
and U3860 (N_3860,In_551,In_915);
nor U3861 (N_3861,In_813,In_817);
xnor U3862 (N_3862,In_958,In_495);
and U3863 (N_3863,In_705,In_163);
or U3864 (N_3864,In_41,In_643);
xnor U3865 (N_3865,In_515,In_125);
nand U3866 (N_3866,In_504,In_67);
nor U3867 (N_3867,In_891,In_790);
nor U3868 (N_3868,In_735,In_184);
or U3869 (N_3869,In_816,In_905);
xnor U3870 (N_3870,In_455,In_556);
xnor U3871 (N_3871,In_124,In_396);
xnor U3872 (N_3872,In_106,In_161);
nand U3873 (N_3873,In_677,In_914);
nand U3874 (N_3874,In_965,In_524);
nor U3875 (N_3875,In_775,In_501);
or U3876 (N_3876,In_750,In_729);
and U3877 (N_3877,In_509,In_609);
nand U3878 (N_3878,In_186,In_958);
or U3879 (N_3879,In_155,In_772);
nand U3880 (N_3880,In_196,In_106);
nor U3881 (N_3881,In_479,In_814);
or U3882 (N_3882,In_132,In_484);
and U3883 (N_3883,In_367,In_202);
nor U3884 (N_3884,In_748,In_77);
xnor U3885 (N_3885,In_517,In_224);
and U3886 (N_3886,In_264,In_41);
and U3887 (N_3887,In_620,In_41);
xnor U3888 (N_3888,In_367,In_757);
and U3889 (N_3889,In_113,In_596);
xnor U3890 (N_3890,In_266,In_967);
nand U3891 (N_3891,In_109,In_594);
and U3892 (N_3892,In_336,In_455);
and U3893 (N_3893,In_399,In_513);
or U3894 (N_3894,In_169,In_726);
nor U3895 (N_3895,In_62,In_649);
nand U3896 (N_3896,In_868,In_197);
nand U3897 (N_3897,In_932,In_475);
and U3898 (N_3898,In_677,In_510);
nor U3899 (N_3899,In_614,In_863);
xnor U3900 (N_3900,In_64,In_507);
or U3901 (N_3901,In_154,In_459);
xnor U3902 (N_3902,In_821,In_987);
xnor U3903 (N_3903,In_732,In_92);
xnor U3904 (N_3904,In_235,In_711);
and U3905 (N_3905,In_663,In_979);
nand U3906 (N_3906,In_480,In_426);
xnor U3907 (N_3907,In_875,In_807);
nor U3908 (N_3908,In_321,In_379);
and U3909 (N_3909,In_831,In_142);
or U3910 (N_3910,In_512,In_225);
and U3911 (N_3911,In_480,In_311);
nor U3912 (N_3912,In_641,In_569);
and U3913 (N_3913,In_924,In_329);
nand U3914 (N_3914,In_419,In_2);
or U3915 (N_3915,In_321,In_44);
or U3916 (N_3916,In_92,In_942);
nand U3917 (N_3917,In_982,In_906);
nand U3918 (N_3918,In_823,In_727);
xor U3919 (N_3919,In_318,In_118);
and U3920 (N_3920,In_804,In_429);
nand U3921 (N_3921,In_144,In_419);
or U3922 (N_3922,In_12,In_546);
nand U3923 (N_3923,In_910,In_582);
and U3924 (N_3924,In_621,In_340);
and U3925 (N_3925,In_995,In_485);
nor U3926 (N_3926,In_716,In_900);
and U3927 (N_3927,In_761,In_964);
xnor U3928 (N_3928,In_446,In_241);
xnor U3929 (N_3929,In_300,In_818);
nand U3930 (N_3930,In_366,In_963);
and U3931 (N_3931,In_920,In_143);
nand U3932 (N_3932,In_935,In_920);
and U3933 (N_3933,In_345,In_320);
xor U3934 (N_3934,In_402,In_343);
nand U3935 (N_3935,In_109,In_722);
and U3936 (N_3936,In_689,In_834);
nand U3937 (N_3937,In_956,In_488);
nand U3938 (N_3938,In_611,In_526);
or U3939 (N_3939,In_883,In_425);
and U3940 (N_3940,In_954,In_963);
and U3941 (N_3941,In_319,In_790);
nand U3942 (N_3942,In_574,In_448);
nand U3943 (N_3943,In_581,In_538);
or U3944 (N_3944,In_610,In_277);
or U3945 (N_3945,In_861,In_372);
and U3946 (N_3946,In_322,In_520);
or U3947 (N_3947,In_936,In_710);
xnor U3948 (N_3948,In_926,In_159);
and U3949 (N_3949,In_832,In_278);
nand U3950 (N_3950,In_279,In_561);
or U3951 (N_3951,In_914,In_311);
or U3952 (N_3952,In_479,In_37);
xnor U3953 (N_3953,In_663,In_601);
nor U3954 (N_3954,In_463,In_106);
nand U3955 (N_3955,In_356,In_355);
and U3956 (N_3956,In_51,In_939);
nor U3957 (N_3957,In_855,In_483);
xor U3958 (N_3958,In_184,In_53);
nand U3959 (N_3959,In_302,In_290);
and U3960 (N_3960,In_393,In_657);
xor U3961 (N_3961,In_372,In_872);
or U3962 (N_3962,In_760,In_720);
nor U3963 (N_3963,In_498,In_905);
nand U3964 (N_3964,In_886,In_889);
and U3965 (N_3965,In_54,In_542);
or U3966 (N_3966,In_574,In_342);
xnor U3967 (N_3967,In_272,In_292);
and U3968 (N_3968,In_754,In_928);
nand U3969 (N_3969,In_354,In_879);
xnor U3970 (N_3970,In_327,In_584);
nor U3971 (N_3971,In_2,In_927);
and U3972 (N_3972,In_655,In_497);
and U3973 (N_3973,In_771,In_677);
or U3974 (N_3974,In_212,In_609);
or U3975 (N_3975,In_68,In_890);
nor U3976 (N_3976,In_919,In_268);
or U3977 (N_3977,In_844,In_409);
and U3978 (N_3978,In_542,In_55);
nor U3979 (N_3979,In_36,In_543);
and U3980 (N_3980,In_86,In_931);
nand U3981 (N_3981,In_954,In_672);
nor U3982 (N_3982,In_548,In_10);
xor U3983 (N_3983,In_760,In_819);
nand U3984 (N_3984,In_376,In_963);
nor U3985 (N_3985,In_217,In_307);
nand U3986 (N_3986,In_488,In_706);
xnor U3987 (N_3987,In_693,In_805);
xnor U3988 (N_3988,In_543,In_742);
xnor U3989 (N_3989,In_893,In_354);
or U3990 (N_3990,In_618,In_910);
xnor U3991 (N_3991,In_27,In_234);
or U3992 (N_3992,In_623,In_945);
and U3993 (N_3993,In_201,In_893);
or U3994 (N_3994,In_282,In_732);
and U3995 (N_3995,In_223,In_926);
xnor U3996 (N_3996,In_596,In_24);
nand U3997 (N_3997,In_405,In_416);
nand U3998 (N_3998,In_804,In_851);
nor U3999 (N_3999,In_710,In_973);
and U4000 (N_4000,In_137,In_970);
xor U4001 (N_4001,In_812,In_893);
or U4002 (N_4002,In_744,In_361);
nor U4003 (N_4003,In_48,In_719);
nand U4004 (N_4004,In_918,In_705);
nand U4005 (N_4005,In_926,In_68);
nand U4006 (N_4006,In_289,In_590);
and U4007 (N_4007,In_963,In_451);
nor U4008 (N_4008,In_86,In_668);
and U4009 (N_4009,In_629,In_313);
xnor U4010 (N_4010,In_562,In_893);
or U4011 (N_4011,In_318,In_436);
xnor U4012 (N_4012,In_300,In_382);
nand U4013 (N_4013,In_439,In_571);
nor U4014 (N_4014,In_732,In_58);
or U4015 (N_4015,In_959,In_323);
or U4016 (N_4016,In_885,In_770);
or U4017 (N_4017,In_863,In_885);
xor U4018 (N_4018,In_166,In_820);
xnor U4019 (N_4019,In_89,In_430);
and U4020 (N_4020,In_173,In_589);
or U4021 (N_4021,In_692,In_822);
and U4022 (N_4022,In_470,In_190);
nor U4023 (N_4023,In_681,In_848);
nor U4024 (N_4024,In_557,In_521);
or U4025 (N_4025,In_790,In_608);
nand U4026 (N_4026,In_674,In_101);
nor U4027 (N_4027,In_323,In_154);
xnor U4028 (N_4028,In_772,In_602);
nor U4029 (N_4029,In_852,In_902);
or U4030 (N_4030,In_893,In_468);
and U4031 (N_4031,In_520,In_381);
xor U4032 (N_4032,In_166,In_444);
nor U4033 (N_4033,In_343,In_504);
or U4034 (N_4034,In_876,In_612);
nor U4035 (N_4035,In_310,In_927);
xnor U4036 (N_4036,In_165,In_616);
nand U4037 (N_4037,In_538,In_801);
xnor U4038 (N_4038,In_18,In_425);
or U4039 (N_4039,In_833,In_810);
or U4040 (N_4040,In_105,In_483);
and U4041 (N_4041,In_550,In_290);
and U4042 (N_4042,In_303,In_425);
or U4043 (N_4043,In_509,In_930);
and U4044 (N_4044,In_10,In_894);
nor U4045 (N_4045,In_873,In_67);
and U4046 (N_4046,In_452,In_453);
nor U4047 (N_4047,In_501,In_802);
and U4048 (N_4048,In_55,In_555);
and U4049 (N_4049,In_992,In_468);
and U4050 (N_4050,In_251,In_497);
nand U4051 (N_4051,In_153,In_973);
xnor U4052 (N_4052,In_938,In_306);
nor U4053 (N_4053,In_106,In_650);
and U4054 (N_4054,In_729,In_745);
xor U4055 (N_4055,In_778,In_405);
nand U4056 (N_4056,In_679,In_733);
nand U4057 (N_4057,In_926,In_603);
and U4058 (N_4058,In_567,In_171);
nor U4059 (N_4059,In_306,In_176);
or U4060 (N_4060,In_63,In_606);
nor U4061 (N_4061,In_3,In_660);
or U4062 (N_4062,In_420,In_218);
xnor U4063 (N_4063,In_179,In_984);
xnor U4064 (N_4064,In_386,In_483);
xnor U4065 (N_4065,In_444,In_118);
xnor U4066 (N_4066,In_425,In_316);
nand U4067 (N_4067,In_104,In_886);
nor U4068 (N_4068,In_512,In_556);
nand U4069 (N_4069,In_634,In_567);
nand U4070 (N_4070,In_29,In_165);
xor U4071 (N_4071,In_436,In_961);
nand U4072 (N_4072,In_7,In_937);
nor U4073 (N_4073,In_580,In_548);
nand U4074 (N_4074,In_297,In_484);
and U4075 (N_4075,In_922,In_10);
and U4076 (N_4076,In_97,In_223);
nor U4077 (N_4077,In_407,In_650);
and U4078 (N_4078,In_755,In_228);
and U4079 (N_4079,In_306,In_817);
or U4080 (N_4080,In_464,In_778);
xnor U4081 (N_4081,In_80,In_213);
xor U4082 (N_4082,In_717,In_141);
nor U4083 (N_4083,In_985,In_805);
nor U4084 (N_4084,In_86,In_427);
and U4085 (N_4085,In_201,In_300);
xnor U4086 (N_4086,In_257,In_640);
nor U4087 (N_4087,In_21,In_222);
or U4088 (N_4088,In_254,In_743);
xor U4089 (N_4089,In_254,In_81);
nand U4090 (N_4090,In_172,In_21);
xor U4091 (N_4091,In_571,In_690);
nand U4092 (N_4092,In_221,In_568);
nor U4093 (N_4093,In_770,In_914);
nor U4094 (N_4094,In_265,In_362);
xnor U4095 (N_4095,In_238,In_43);
xor U4096 (N_4096,In_369,In_433);
or U4097 (N_4097,In_906,In_490);
and U4098 (N_4098,In_177,In_42);
xor U4099 (N_4099,In_228,In_501);
xor U4100 (N_4100,In_757,In_434);
and U4101 (N_4101,In_174,In_995);
nor U4102 (N_4102,In_668,In_866);
or U4103 (N_4103,In_393,In_724);
xor U4104 (N_4104,In_346,In_811);
nor U4105 (N_4105,In_251,In_399);
xor U4106 (N_4106,In_739,In_407);
nand U4107 (N_4107,In_844,In_42);
nand U4108 (N_4108,In_361,In_217);
or U4109 (N_4109,In_795,In_536);
xor U4110 (N_4110,In_18,In_414);
nand U4111 (N_4111,In_419,In_151);
nor U4112 (N_4112,In_660,In_775);
nand U4113 (N_4113,In_272,In_485);
nor U4114 (N_4114,In_493,In_690);
nand U4115 (N_4115,In_953,In_852);
xor U4116 (N_4116,In_741,In_367);
nand U4117 (N_4117,In_586,In_969);
xnor U4118 (N_4118,In_409,In_900);
xor U4119 (N_4119,In_653,In_64);
and U4120 (N_4120,In_26,In_37);
nand U4121 (N_4121,In_209,In_604);
nand U4122 (N_4122,In_274,In_273);
and U4123 (N_4123,In_92,In_137);
xor U4124 (N_4124,In_559,In_921);
or U4125 (N_4125,In_836,In_651);
xnor U4126 (N_4126,In_312,In_818);
or U4127 (N_4127,In_132,In_121);
nand U4128 (N_4128,In_661,In_98);
and U4129 (N_4129,In_465,In_620);
nand U4130 (N_4130,In_163,In_871);
nor U4131 (N_4131,In_465,In_903);
xor U4132 (N_4132,In_178,In_418);
and U4133 (N_4133,In_437,In_476);
or U4134 (N_4134,In_5,In_436);
xor U4135 (N_4135,In_375,In_817);
xor U4136 (N_4136,In_900,In_147);
and U4137 (N_4137,In_807,In_263);
xor U4138 (N_4138,In_27,In_198);
nor U4139 (N_4139,In_968,In_638);
xnor U4140 (N_4140,In_187,In_186);
and U4141 (N_4141,In_782,In_436);
and U4142 (N_4142,In_141,In_309);
or U4143 (N_4143,In_15,In_797);
nor U4144 (N_4144,In_483,In_136);
and U4145 (N_4145,In_152,In_900);
xnor U4146 (N_4146,In_942,In_67);
and U4147 (N_4147,In_81,In_827);
or U4148 (N_4148,In_951,In_499);
nand U4149 (N_4149,In_53,In_219);
or U4150 (N_4150,In_110,In_595);
xor U4151 (N_4151,In_409,In_916);
or U4152 (N_4152,In_369,In_124);
and U4153 (N_4153,In_212,In_500);
and U4154 (N_4154,In_96,In_59);
xor U4155 (N_4155,In_133,In_182);
and U4156 (N_4156,In_252,In_289);
and U4157 (N_4157,In_853,In_610);
or U4158 (N_4158,In_288,In_150);
nor U4159 (N_4159,In_58,In_545);
and U4160 (N_4160,In_258,In_236);
or U4161 (N_4161,In_741,In_96);
or U4162 (N_4162,In_996,In_502);
nor U4163 (N_4163,In_787,In_854);
nand U4164 (N_4164,In_785,In_298);
xnor U4165 (N_4165,In_672,In_28);
and U4166 (N_4166,In_935,In_638);
nand U4167 (N_4167,In_578,In_994);
or U4168 (N_4168,In_664,In_367);
or U4169 (N_4169,In_117,In_158);
nor U4170 (N_4170,In_909,In_51);
nor U4171 (N_4171,In_637,In_208);
nand U4172 (N_4172,In_620,In_18);
and U4173 (N_4173,In_647,In_399);
or U4174 (N_4174,In_300,In_180);
or U4175 (N_4175,In_141,In_783);
xnor U4176 (N_4176,In_30,In_381);
or U4177 (N_4177,In_423,In_540);
or U4178 (N_4178,In_786,In_580);
xnor U4179 (N_4179,In_129,In_434);
xnor U4180 (N_4180,In_950,In_363);
and U4181 (N_4181,In_823,In_449);
nor U4182 (N_4182,In_209,In_88);
nand U4183 (N_4183,In_341,In_255);
and U4184 (N_4184,In_487,In_453);
and U4185 (N_4185,In_732,In_857);
and U4186 (N_4186,In_6,In_993);
and U4187 (N_4187,In_171,In_491);
or U4188 (N_4188,In_687,In_809);
or U4189 (N_4189,In_399,In_37);
or U4190 (N_4190,In_743,In_580);
nand U4191 (N_4191,In_396,In_27);
nand U4192 (N_4192,In_76,In_34);
or U4193 (N_4193,In_673,In_616);
or U4194 (N_4194,In_775,In_804);
xor U4195 (N_4195,In_920,In_608);
and U4196 (N_4196,In_150,In_864);
and U4197 (N_4197,In_185,In_891);
nand U4198 (N_4198,In_273,In_861);
or U4199 (N_4199,In_550,In_917);
and U4200 (N_4200,In_674,In_848);
and U4201 (N_4201,In_968,In_535);
xor U4202 (N_4202,In_319,In_150);
and U4203 (N_4203,In_172,In_9);
or U4204 (N_4204,In_802,In_133);
and U4205 (N_4205,In_259,In_875);
nor U4206 (N_4206,In_905,In_595);
nand U4207 (N_4207,In_679,In_644);
and U4208 (N_4208,In_892,In_307);
nor U4209 (N_4209,In_894,In_740);
or U4210 (N_4210,In_438,In_238);
or U4211 (N_4211,In_372,In_930);
xnor U4212 (N_4212,In_586,In_216);
nand U4213 (N_4213,In_169,In_985);
xor U4214 (N_4214,In_350,In_563);
and U4215 (N_4215,In_167,In_226);
xnor U4216 (N_4216,In_726,In_803);
nand U4217 (N_4217,In_786,In_490);
or U4218 (N_4218,In_810,In_981);
xor U4219 (N_4219,In_216,In_231);
nand U4220 (N_4220,In_717,In_104);
nor U4221 (N_4221,In_43,In_112);
nand U4222 (N_4222,In_329,In_851);
and U4223 (N_4223,In_549,In_129);
and U4224 (N_4224,In_65,In_431);
nor U4225 (N_4225,In_411,In_772);
or U4226 (N_4226,In_269,In_676);
and U4227 (N_4227,In_806,In_308);
xnor U4228 (N_4228,In_365,In_535);
and U4229 (N_4229,In_9,In_210);
xnor U4230 (N_4230,In_238,In_332);
and U4231 (N_4231,In_639,In_607);
or U4232 (N_4232,In_910,In_911);
nand U4233 (N_4233,In_929,In_106);
xnor U4234 (N_4234,In_452,In_265);
xnor U4235 (N_4235,In_292,In_764);
or U4236 (N_4236,In_635,In_253);
or U4237 (N_4237,In_611,In_509);
nand U4238 (N_4238,In_291,In_426);
nand U4239 (N_4239,In_52,In_162);
or U4240 (N_4240,In_300,In_894);
or U4241 (N_4241,In_876,In_150);
nor U4242 (N_4242,In_679,In_473);
nor U4243 (N_4243,In_231,In_215);
xnor U4244 (N_4244,In_317,In_589);
and U4245 (N_4245,In_734,In_757);
nand U4246 (N_4246,In_654,In_810);
or U4247 (N_4247,In_105,In_83);
xnor U4248 (N_4248,In_413,In_323);
nand U4249 (N_4249,In_438,In_989);
nand U4250 (N_4250,In_349,In_299);
and U4251 (N_4251,In_969,In_679);
and U4252 (N_4252,In_497,In_12);
xnor U4253 (N_4253,In_409,In_10);
nand U4254 (N_4254,In_203,In_821);
nor U4255 (N_4255,In_181,In_206);
xor U4256 (N_4256,In_391,In_173);
and U4257 (N_4257,In_245,In_924);
or U4258 (N_4258,In_901,In_851);
xnor U4259 (N_4259,In_137,In_521);
and U4260 (N_4260,In_253,In_60);
or U4261 (N_4261,In_485,In_920);
nand U4262 (N_4262,In_343,In_344);
and U4263 (N_4263,In_642,In_315);
nor U4264 (N_4264,In_717,In_152);
nor U4265 (N_4265,In_372,In_599);
or U4266 (N_4266,In_208,In_489);
nor U4267 (N_4267,In_475,In_903);
xor U4268 (N_4268,In_693,In_567);
and U4269 (N_4269,In_922,In_770);
or U4270 (N_4270,In_697,In_364);
nor U4271 (N_4271,In_119,In_603);
nor U4272 (N_4272,In_821,In_129);
nor U4273 (N_4273,In_952,In_334);
or U4274 (N_4274,In_688,In_123);
and U4275 (N_4275,In_8,In_940);
nor U4276 (N_4276,In_467,In_585);
and U4277 (N_4277,In_121,In_527);
nand U4278 (N_4278,In_627,In_860);
nor U4279 (N_4279,In_689,In_449);
and U4280 (N_4280,In_904,In_600);
xnor U4281 (N_4281,In_522,In_489);
and U4282 (N_4282,In_144,In_905);
nand U4283 (N_4283,In_717,In_26);
or U4284 (N_4284,In_940,In_920);
xor U4285 (N_4285,In_582,In_588);
nor U4286 (N_4286,In_418,In_711);
nand U4287 (N_4287,In_380,In_479);
xor U4288 (N_4288,In_234,In_165);
nor U4289 (N_4289,In_902,In_155);
or U4290 (N_4290,In_560,In_354);
xor U4291 (N_4291,In_501,In_929);
or U4292 (N_4292,In_961,In_208);
nand U4293 (N_4293,In_64,In_423);
xor U4294 (N_4294,In_164,In_165);
nand U4295 (N_4295,In_62,In_711);
and U4296 (N_4296,In_632,In_80);
nor U4297 (N_4297,In_957,In_187);
and U4298 (N_4298,In_932,In_338);
xnor U4299 (N_4299,In_239,In_529);
nor U4300 (N_4300,In_832,In_41);
nand U4301 (N_4301,In_127,In_351);
and U4302 (N_4302,In_651,In_460);
and U4303 (N_4303,In_814,In_489);
and U4304 (N_4304,In_139,In_89);
or U4305 (N_4305,In_427,In_419);
or U4306 (N_4306,In_261,In_635);
nor U4307 (N_4307,In_662,In_151);
nor U4308 (N_4308,In_632,In_316);
and U4309 (N_4309,In_362,In_23);
nor U4310 (N_4310,In_550,In_453);
nand U4311 (N_4311,In_760,In_785);
and U4312 (N_4312,In_29,In_504);
xnor U4313 (N_4313,In_60,In_880);
xor U4314 (N_4314,In_248,In_87);
nand U4315 (N_4315,In_702,In_791);
xor U4316 (N_4316,In_272,In_631);
or U4317 (N_4317,In_220,In_942);
nor U4318 (N_4318,In_806,In_30);
or U4319 (N_4319,In_359,In_25);
nor U4320 (N_4320,In_40,In_198);
nand U4321 (N_4321,In_849,In_979);
and U4322 (N_4322,In_816,In_821);
nand U4323 (N_4323,In_992,In_505);
nor U4324 (N_4324,In_869,In_488);
nand U4325 (N_4325,In_688,In_637);
xor U4326 (N_4326,In_348,In_638);
xor U4327 (N_4327,In_388,In_67);
nand U4328 (N_4328,In_420,In_377);
xnor U4329 (N_4329,In_304,In_117);
or U4330 (N_4330,In_185,In_298);
and U4331 (N_4331,In_279,In_486);
nand U4332 (N_4332,In_642,In_859);
xor U4333 (N_4333,In_919,In_689);
or U4334 (N_4334,In_720,In_633);
or U4335 (N_4335,In_155,In_939);
nor U4336 (N_4336,In_826,In_228);
xor U4337 (N_4337,In_828,In_203);
and U4338 (N_4338,In_74,In_362);
xnor U4339 (N_4339,In_430,In_398);
xor U4340 (N_4340,In_314,In_684);
xnor U4341 (N_4341,In_982,In_951);
xnor U4342 (N_4342,In_462,In_496);
xor U4343 (N_4343,In_906,In_799);
xor U4344 (N_4344,In_365,In_11);
xor U4345 (N_4345,In_472,In_935);
or U4346 (N_4346,In_156,In_159);
xor U4347 (N_4347,In_273,In_102);
and U4348 (N_4348,In_962,In_267);
and U4349 (N_4349,In_437,In_752);
nand U4350 (N_4350,In_80,In_71);
nand U4351 (N_4351,In_36,In_41);
and U4352 (N_4352,In_929,In_494);
nor U4353 (N_4353,In_64,In_102);
nor U4354 (N_4354,In_407,In_368);
and U4355 (N_4355,In_793,In_987);
or U4356 (N_4356,In_685,In_884);
nand U4357 (N_4357,In_665,In_243);
nor U4358 (N_4358,In_472,In_473);
or U4359 (N_4359,In_96,In_149);
xnor U4360 (N_4360,In_979,In_67);
nand U4361 (N_4361,In_636,In_854);
and U4362 (N_4362,In_61,In_824);
nor U4363 (N_4363,In_523,In_687);
xor U4364 (N_4364,In_949,In_89);
or U4365 (N_4365,In_133,In_938);
nand U4366 (N_4366,In_429,In_712);
xnor U4367 (N_4367,In_107,In_763);
nor U4368 (N_4368,In_664,In_349);
xor U4369 (N_4369,In_30,In_607);
or U4370 (N_4370,In_640,In_511);
and U4371 (N_4371,In_841,In_75);
nor U4372 (N_4372,In_275,In_686);
nor U4373 (N_4373,In_121,In_691);
nor U4374 (N_4374,In_77,In_569);
and U4375 (N_4375,In_166,In_442);
nand U4376 (N_4376,In_405,In_918);
nor U4377 (N_4377,In_325,In_757);
or U4378 (N_4378,In_622,In_662);
nor U4379 (N_4379,In_18,In_86);
or U4380 (N_4380,In_198,In_909);
xor U4381 (N_4381,In_719,In_8);
xor U4382 (N_4382,In_730,In_428);
nor U4383 (N_4383,In_191,In_319);
nor U4384 (N_4384,In_791,In_823);
and U4385 (N_4385,In_632,In_259);
nand U4386 (N_4386,In_695,In_627);
or U4387 (N_4387,In_221,In_645);
nand U4388 (N_4388,In_659,In_148);
xor U4389 (N_4389,In_621,In_736);
nor U4390 (N_4390,In_211,In_188);
nand U4391 (N_4391,In_256,In_703);
or U4392 (N_4392,In_66,In_664);
and U4393 (N_4393,In_706,In_102);
or U4394 (N_4394,In_806,In_845);
and U4395 (N_4395,In_506,In_920);
xnor U4396 (N_4396,In_170,In_699);
xnor U4397 (N_4397,In_363,In_969);
nor U4398 (N_4398,In_502,In_598);
nor U4399 (N_4399,In_692,In_632);
or U4400 (N_4400,In_468,In_525);
nor U4401 (N_4401,In_338,In_680);
or U4402 (N_4402,In_837,In_179);
nand U4403 (N_4403,In_465,In_855);
xnor U4404 (N_4404,In_951,In_676);
or U4405 (N_4405,In_933,In_499);
or U4406 (N_4406,In_712,In_117);
nor U4407 (N_4407,In_868,In_898);
nand U4408 (N_4408,In_953,In_898);
nand U4409 (N_4409,In_195,In_390);
or U4410 (N_4410,In_943,In_915);
nor U4411 (N_4411,In_711,In_460);
or U4412 (N_4412,In_724,In_660);
nor U4413 (N_4413,In_59,In_9);
nand U4414 (N_4414,In_649,In_730);
or U4415 (N_4415,In_515,In_422);
xor U4416 (N_4416,In_833,In_61);
nor U4417 (N_4417,In_192,In_226);
nand U4418 (N_4418,In_605,In_493);
xor U4419 (N_4419,In_610,In_453);
or U4420 (N_4420,In_128,In_752);
or U4421 (N_4421,In_69,In_500);
and U4422 (N_4422,In_897,In_464);
xnor U4423 (N_4423,In_127,In_995);
nor U4424 (N_4424,In_793,In_72);
and U4425 (N_4425,In_614,In_309);
and U4426 (N_4426,In_140,In_777);
xnor U4427 (N_4427,In_740,In_241);
nor U4428 (N_4428,In_499,In_404);
xnor U4429 (N_4429,In_791,In_460);
and U4430 (N_4430,In_471,In_593);
xnor U4431 (N_4431,In_453,In_214);
or U4432 (N_4432,In_93,In_980);
xor U4433 (N_4433,In_594,In_846);
and U4434 (N_4434,In_2,In_692);
and U4435 (N_4435,In_569,In_315);
nand U4436 (N_4436,In_449,In_235);
nor U4437 (N_4437,In_300,In_859);
and U4438 (N_4438,In_307,In_825);
and U4439 (N_4439,In_339,In_593);
or U4440 (N_4440,In_304,In_909);
nand U4441 (N_4441,In_950,In_257);
and U4442 (N_4442,In_361,In_908);
nor U4443 (N_4443,In_401,In_427);
or U4444 (N_4444,In_53,In_60);
nand U4445 (N_4445,In_904,In_943);
and U4446 (N_4446,In_962,In_68);
nor U4447 (N_4447,In_360,In_931);
nor U4448 (N_4448,In_759,In_628);
or U4449 (N_4449,In_120,In_687);
xor U4450 (N_4450,In_98,In_516);
nor U4451 (N_4451,In_101,In_606);
nand U4452 (N_4452,In_704,In_627);
or U4453 (N_4453,In_207,In_225);
xor U4454 (N_4454,In_292,In_702);
and U4455 (N_4455,In_546,In_466);
nor U4456 (N_4456,In_506,In_6);
or U4457 (N_4457,In_956,In_943);
and U4458 (N_4458,In_823,In_662);
nor U4459 (N_4459,In_874,In_210);
and U4460 (N_4460,In_68,In_869);
or U4461 (N_4461,In_550,In_780);
xor U4462 (N_4462,In_509,In_790);
or U4463 (N_4463,In_998,In_169);
xor U4464 (N_4464,In_386,In_784);
xor U4465 (N_4465,In_207,In_710);
or U4466 (N_4466,In_485,In_592);
or U4467 (N_4467,In_736,In_808);
or U4468 (N_4468,In_682,In_207);
and U4469 (N_4469,In_767,In_815);
nand U4470 (N_4470,In_567,In_757);
nor U4471 (N_4471,In_710,In_10);
nand U4472 (N_4472,In_523,In_639);
or U4473 (N_4473,In_993,In_742);
or U4474 (N_4474,In_739,In_748);
xor U4475 (N_4475,In_140,In_170);
xnor U4476 (N_4476,In_47,In_993);
and U4477 (N_4477,In_738,In_160);
xor U4478 (N_4478,In_781,In_663);
nand U4479 (N_4479,In_8,In_488);
or U4480 (N_4480,In_961,In_89);
xor U4481 (N_4481,In_225,In_760);
xor U4482 (N_4482,In_684,In_671);
nand U4483 (N_4483,In_184,In_638);
nor U4484 (N_4484,In_788,In_478);
nand U4485 (N_4485,In_378,In_854);
and U4486 (N_4486,In_486,In_137);
or U4487 (N_4487,In_921,In_123);
nand U4488 (N_4488,In_606,In_836);
or U4489 (N_4489,In_18,In_963);
and U4490 (N_4490,In_736,In_987);
and U4491 (N_4491,In_527,In_332);
or U4492 (N_4492,In_481,In_739);
nand U4493 (N_4493,In_10,In_786);
xor U4494 (N_4494,In_753,In_626);
nor U4495 (N_4495,In_705,In_578);
nor U4496 (N_4496,In_1,In_652);
xnor U4497 (N_4497,In_717,In_800);
and U4498 (N_4498,In_506,In_352);
and U4499 (N_4499,In_848,In_550);
or U4500 (N_4500,In_183,In_67);
nand U4501 (N_4501,In_921,In_698);
and U4502 (N_4502,In_692,In_84);
and U4503 (N_4503,In_85,In_964);
nand U4504 (N_4504,In_895,In_154);
nor U4505 (N_4505,In_67,In_523);
xnor U4506 (N_4506,In_613,In_950);
and U4507 (N_4507,In_332,In_167);
nor U4508 (N_4508,In_801,In_909);
xor U4509 (N_4509,In_665,In_889);
nand U4510 (N_4510,In_775,In_913);
xor U4511 (N_4511,In_813,In_404);
xor U4512 (N_4512,In_25,In_80);
nor U4513 (N_4513,In_795,In_255);
and U4514 (N_4514,In_340,In_818);
nor U4515 (N_4515,In_598,In_582);
or U4516 (N_4516,In_270,In_880);
nand U4517 (N_4517,In_969,In_233);
nand U4518 (N_4518,In_907,In_404);
or U4519 (N_4519,In_907,In_332);
nand U4520 (N_4520,In_976,In_642);
nand U4521 (N_4521,In_845,In_766);
nor U4522 (N_4522,In_54,In_572);
and U4523 (N_4523,In_783,In_181);
nor U4524 (N_4524,In_230,In_280);
nor U4525 (N_4525,In_228,In_434);
and U4526 (N_4526,In_47,In_550);
xnor U4527 (N_4527,In_852,In_173);
xor U4528 (N_4528,In_407,In_346);
xor U4529 (N_4529,In_3,In_480);
nand U4530 (N_4530,In_195,In_68);
nand U4531 (N_4531,In_427,In_940);
nor U4532 (N_4532,In_692,In_282);
nor U4533 (N_4533,In_0,In_816);
and U4534 (N_4534,In_992,In_260);
nor U4535 (N_4535,In_791,In_880);
nor U4536 (N_4536,In_969,In_971);
xor U4537 (N_4537,In_558,In_640);
and U4538 (N_4538,In_791,In_639);
or U4539 (N_4539,In_700,In_970);
or U4540 (N_4540,In_472,In_406);
nand U4541 (N_4541,In_763,In_787);
nand U4542 (N_4542,In_584,In_377);
xnor U4543 (N_4543,In_153,In_785);
nand U4544 (N_4544,In_839,In_10);
xor U4545 (N_4545,In_32,In_336);
and U4546 (N_4546,In_754,In_837);
nor U4547 (N_4547,In_348,In_761);
nor U4548 (N_4548,In_817,In_683);
or U4549 (N_4549,In_54,In_522);
nand U4550 (N_4550,In_194,In_756);
nor U4551 (N_4551,In_278,In_998);
and U4552 (N_4552,In_759,In_918);
nor U4553 (N_4553,In_876,In_607);
or U4554 (N_4554,In_447,In_665);
and U4555 (N_4555,In_247,In_705);
nor U4556 (N_4556,In_857,In_111);
and U4557 (N_4557,In_409,In_31);
nand U4558 (N_4558,In_367,In_883);
or U4559 (N_4559,In_438,In_366);
nor U4560 (N_4560,In_38,In_309);
and U4561 (N_4561,In_773,In_300);
xor U4562 (N_4562,In_799,In_324);
nand U4563 (N_4563,In_407,In_758);
nor U4564 (N_4564,In_164,In_954);
or U4565 (N_4565,In_16,In_82);
and U4566 (N_4566,In_243,In_667);
and U4567 (N_4567,In_590,In_526);
and U4568 (N_4568,In_635,In_139);
xor U4569 (N_4569,In_979,In_68);
xnor U4570 (N_4570,In_586,In_217);
nand U4571 (N_4571,In_735,In_106);
and U4572 (N_4572,In_926,In_108);
nor U4573 (N_4573,In_711,In_946);
xnor U4574 (N_4574,In_113,In_975);
and U4575 (N_4575,In_617,In_650);
or U4576 (N_4576,In_45,In_764);
nor U4577 (N_4577,In_712,In_141);
nand U4578 (N_4578,In_258,In_120);
and U4579 (N_4579,In_94,In_767);
nand U4580 (N_4580,In_581,In_238);
and U4581 (N_4581,In_688,In_196);
or U4582 (N_4582,In_830,In_835);
nor U4583 (N_4583,In_942,In_613);
xnor U4584 (N_4584,In_203,In_399);
and U4585 (N_4585,In_424,In_392);
or U4586 (N_4586,In_479,In_410);
nand U4587 (N_4587,In_898,In_84);
nor U4588 (N_4588,In_233,In_671);
nand U4589 (N_4589,In_677,In_801);
nor U4590 (N_4590,In_321,In_259);
and U4591 (N_4591,In_146,In_617);
xor U4592 (N_4592,In_133,In_178);
and U4593 (N_4593,In_946,In_74);
and U4594 (N_4594,In_232,In_746);
nand U4595 (N_4595,In_903,In_96);
nand U4596 (N_4596,In_46,In_259);
xor U4597 (N_4597,In_860,In_717);
nand U4598 (N_4598,In_940,In_144);
nor U4599 (N_4599,In_484,In_377);
xor U4600 (N_4600,In_771,In_639);
or U4601 (N_4601,In_523,In_410);
or U4602 (N_4602,In_950,In_570);
or U4603 (N_4603,In_621,In_74);
nor U4604 (N_4604,In_245,In_457);
or U4605 (N_4605,In_738,In_286);
xor U4606 (N_4606,In_811,In_824);
xnor U4607 (N_4607,In_644,In_622);
and U4608 (N_4608,In_437,In_69);
or U4609 (N_4609,In_602,In_66);
xnor U4610 (N_4610,In_711,In_30);
xnor U4611 (N_4611,In_745,In_306);
nand U4612 (N_4612,In_652,In_170);
nand U4613 (N_4613,In_894,In_419);
or U4614 (N_4614,In_539,In_36);
or U4615 (N_4615,In_58,In_224);
nand U4616 (N_4616,In_863,In_275);
or U4617 (N_4617,In_384,In_11);
nand U4618 (N_4618,In_867,In_648);
and U4619 (N_4619,In_247,In_596);
nand U4620 (N_4620,In_205,In_825);
and U4621 (N_4621,In_806,In_637);
and U4622 (N_4622,In_3,In_310);
nor U4623 (N_4623,In_784,In_204);
and U4624 (N_4624,In_419,In_567);
nor U4625 (N_4625,In_409,In_404);
nor U4626 (N_4626,In_89,In_836);
nand U4627 (N_4627,In_125,In_573);
nand U4628 (N_4628,In_854,In_347);
nor U4629 (N_4629,In_918,In_851);
and U4630 (N_4630,In_958,In_454);
nand U4631 (N_4631,In_935,In_929);
xnor U4632 (N_4632,In_375,In_748);
or U4633 (N_4633,In_983,In_762);
nor U4634 (N_4634,In_365,In_622);
and U4635 (N_4635,In_429,In_815);
or U4636 (N_4636,In_945,In_871);
xor U4637 (N_4637,In_166,In_523);
or U4638 (N_4638,In_904,In_178);
and U4639 (N_4639,In_225,In_436);
xor U4640 (N_4640,In_437,In_657);
nand U4641 (N_4641,In_492,In_386);
nor U4642 (N_4642,In_77,In_165);
and U4643 (N_4643,In_730,In_486);
nand U4644 (N_4644,In_311,In_617);
nand U4645 (N_4645,In_305,In_27);
and U4646 (N_4646,In_665,In_530);
xnor U4647 (N_4647,In_418,In_163);
nor U4648 (N_4648,In_31,In_380);
nand U4649 (N_4649,In_72,In_773);
nor U4650 (N_4650,In_915,In_415);
or U4651 (N_4651,In_322,In_616);
xnor U4652 (N_4652,In_155,In_534);
and U4653 (N_4653,In_261,In_973);
nand U4654 (N_4654,In_410,In_721);
nand U4655 (N_4655,In_517,In_967);
and U4656 (N_4656,In_673,In_980);
nor U4657 (N_4657,In_490,In_228);
nand U4658 (N_4658,In_165,In_688);
xor U4659 (N_4659,In_819,In_86);
nand U4660 (N_4660,In_816,In_258);
nand U4661 (N_4661,In_855,In_519);
xnor U4662 (N_4662,In_993,In_270);
and U4663 (N_4663,In_688,In_333);
xnor U4664 (N_4664,In_526,In_548);
xnor U4665 (N_4665,In_176,In_753);
or U4666 (N_4666,In_787,In_191);
nor U4667 (N_4667,In_214,In_628);
nand U4668 (N_4668,In_568,In_123);
xor U4669 (N_4669,In_413,In_687);
nand U4670 (N_4670,In_124,In_895);
xnor U4671 (N_4671,In_701,In_85);
nor U4672 (N_4672,In_637,In_780);
nor U4673 (N_4673,In_228,In_607);
nand U4674 (N_4674,In_803,In_353);
nor U4675 (N_4675,In_830,In_170);
xor U4676 (N_4676,In_567,In_587);
nor U4677 (N_4677,In_952,In_422);
and U4678 (N_4678,In_918,In_725);
and U4679 (N_4679,In_234,In_721);
and U4680 (N_4680,In_571,In_712);
or U4681 (N_4681,In_696,In_242);
nor U4682 (N_4682,In_295,In_435);
nand U4683 (N_4683,In_45,In_261);
xnor U4684 (N_4684,In_802,In_732);
and U4685 (N_4685,In_350,In_995);
xor U4686 (N_4686,In_690,In_569);
nor U4687 (N_4687,In_491,In_551);
or U4688 (N_4688,In_6,In_817);
xnor U4689 (N_4689,In_757,In_888);
nor U4690 (N_4690,In_593,In_390);
xnor U4691 (N_4691,In_46,In_61);
nand U4692 (N_4692,In_843,In_278);
and U4693 (N_4693,In_758,In_510);
or U4694 (N_4694,In_416,In_967);
or U4695 (N_4695,In_484,In_33);
xnor U4696 (N_4696,In_518,In_418);
or U4697 (N_4697,In_89,In_999);
nor U4698 (N_4698,In_23,In_797);
nand U4699 (N_4699,In_80,In_282);
or U4700 (N_4700,In_713,In_7);
nor U4701 (N_4701,In_225,In_146);
or U4702 (N_4702,In_271,In_191);
nand U4703 (N_4703,In_598,In_879);
and U4704 (N_4704,In_595,In_90);
nor U4705 (N_4705,In_143,In_662);
and U4706 (N_4706,In_300,In_612);
xnor U4707 (N_4707,In_520,In_639);
xnor U4708 (N_4708,In_675,In_454);
nand U4709 (N_4709,In_278,In_673);
or U4710 (N_4710,In_242,In_759);
xor U4711 (N_4711,In_832,In_51);
nand U4712 (N_4712,In_801,In_396);
or U4713 (N_4713,In_341,In_6);
nor U4714 (N_4714,In_443,In_270);
or U4715 (N_4715,In_952,In_816);
or U4716 (N_4716,In_795,In_334);
or U4717 (N_4717,In_182,In_417);
nand U4718 (N_4718,In_567,In_869);
nor U4719 (N_4719,In_610,In_805);
or U4720 (N_4720,In_910,In_153);
nand U4721 (N_4721,In_250,In_17);
nand U4722 (N_4722,In_828,In_56);
xnor U4723 (N_4723,In_137,In_695);
xnor U4724 (N_4724,In_853,In_684);
xnor U4725 (N_4725,In_921,In_162);
or U4726 (N_4726,In_191,In_454);
nand U4727 (N_4727,In_715,In_378);
or U4728 (N_4728,In_670,In_263);
and U4729 (N_4729,In_709,In_609);
nor U4730 (N_4730,In_389,In_672);
and U4731 (N_4731,In_266,In_510);
xnor U4732 (N_4732,In_131,In_601);
xnor U4733 (N_4733,In_774,In_162);
or U4734 (N_4734,In_994,In_669);
xnor U4735 (N_4735,In_649,In_525);
xnor U4736 (N_4736,In_377,In_799);
xnor U4737 (N_4737,In_671,In_141);
or U4738 (N_4738,In_903,In_781);
nand U4739 (N_4739,In_290,In_408);
nor U4740 (N_4740,In_852,In_399);
xnor U4741 (N_4741,In_407,In_373);
or U4742 (N_4742,In_98,In_910);
nand U4743 (N_4743,In_948,In_308);
or U4744 (N_4744,In_730,In_7);
nor U4745 (N_4745,In_201,In_191);
nand U4746 (N_4746,In_535,In_492);
nand U4747 (N_4747,In_112,In_879);
xnor U4748 (N_4748,In_873,In_174);
xnor U4749 (N_4749,In_180,In_883);
xnor U4750 (N_4750,In_249,In_327);
and U4751 (N_4751,In_503,In_711);
or U4752 (N_4752,In_741,In_52);
and U4753 (N_4753,In_849,In_916);
nor U4754 (N_4754,In_848,In_863);
xor U4755 (N_4755,In_775,In_121);
nor U4756 (N_4756,In_604,In_417);
or U4757 (N_4757,In_451,In_990);
or U4758 (N_4758,In_490,In_436);
or U4759 (N_4759,In_363,In_639);
xor U4760 (N_4760,In_365,In_595);
nand U4761 (N_4761,In_653,In_898);
xor U4762 (N_4762,In_634,In_314);
nor U4763 (N_4763,In_690,In_699);
xnor U4764 (N_4764,In_224,In_174);
or U4765 (N_4765,In_883,In_108);
and U4766 (N_4766,In_492,In_666);
or U4767 (N_4767,In_667,In_801);
nor U4768 (N_4768,In_167,In_497);
and U4769 (N_4769,In_684,In_811);
or U4770 (N_4770,In_82,In_29);
xor U4771 (N_4771,In_506,In_321);
or U4772 (N_4772,In_186,In_715);
or U4773 (N_4773,In_76,In_686);
nor U4774 (N_4774,In_735,In_334);
and U4775 (N_4775,In_548,In_207);
nand U4776 (N_4776,In_736,In_951);
nor U4777 (N_4777,In_969,In_190);
nand U4778 (N_4778,In_66,In_555);
xnor U4779 (N_4779,In_831,In_939);
or U4780 (N_4780,In_167,In_677);
xnor U4781 (N_4781,In_153,In_574);
and U4782 (N_4782,In_820,In_470);
nand U4783 (N_4783,In_237,In_313);
and U4784 (N_4784,In_332,In_138);
xnor U4785 (N_4785,In_2,In_429);
or U4786 (N_4786,In_204,In_442);
nor U4787 (N_4787,In_698,In_875);
xnor U4788 (N_4788,In_212,In_382);
xor U4789 (N_4789,In_688,In_313);
nand U4790 (N_4790,In_586,In_554);
nor U4791 (N_4791,In_765,In_487);
nand U4792 (N_4792,In_961,In_821);
xnor U4793 (N_4793,In_208,In_809);
xnor U4794 (N_4794,In_84,In_600);
xnor U4795 (N_4795,In_132,In_122);
or U4796 (N_4796,In_688,In_764);
nand U4797 (N_4797,In_423,In_311);
or U4798 (N_4798,In_137,In_751);
or U4799 (N_4799,In_364,In_685);
nor U4800 (N_4800,In_989,In_794);
or U4801 (N_4801,In_339,In_880);
or U4802 (N_4802,In_936,In_48);
or U4803 (N_4803,In_956,In_694);
xor U4804 (N_4804,In_85,In_20);
xnor U4805 (N_4805,In_213,In_544);
and U4806 (N_4806,In_813,In_127);
and U4807 (N_4807,In_979,In_181);
nor U4808 (N_4808,In_14,In_711);
xor U4809 (N_4809,In_37,In_245);
nor U4810 (N_4810,In_471,In_346);
or U4811 (N_4811,In_85,In_577);
or U4812 (N_4812,In_458,In_109);
nor U4813 (N_4813,In_423,In_990);
and U4814 (N_4814,In_561,In_843);
nor U4815 (N_4815,In_679,In_715);
nand U4816 (N_4816,In_857,In_802);
xor U4817 (N_4817,In_681,In_885);
nor U4818 (N_4818,In_485,In_562);
and U4819 (N_4819,In_589,In_840);
or U4820 (N_4820,In_693,In_643);
xnor U4821 (N_4821,In_134,In_967);
xor U4822 (N_4822,In_736,In_30);
nand U4823 (N_4823,In_59,In_377);
nand U4824 (N_4824,In_734,In_511);
or U4825 (N_4825,In_180,In_55);
and U4826 (N_4826,In_992,In_564);
nor U4827 (N_4827,In_774,In_123);
and U4828 (N_4828,In_752,In_220);
nor U4829 (N_4829,In_33,In_941);
nand U4830 (N_4830,In_579,In_681);
and U4831 (N_4831,In_367,In_415);
or U4832 (N_4832,In_199,In_756);
nor U4833 (N_4833,In_558,In_697);
and U4834 (N_4834,In_827,In_609);
nand U4835 (N_4835,In_534,In_249);
nor U4836 (N_4836,In_782,In_220);
and U4837 (N_4837,In_999,In_19);
nor U4838 (N_4838,In_762,In_390);
nand U4839 (N_4839,In_387,In_146);
nor U4840 (N_4840,In_490,In_657);
nand U4841 (N_4841,In_181,In_735);
nor U4842 (N_4842,In_661,In_32);
nand U4843 (N_4843,In_906,In_652);
nor U4844 (N_4844,In_1,In_854);
or U4845 (N_4845,In_709,In_688);
xor U4846 (N_4846,In_82,In_642);
nand U4847 (N_4847,In_569,In_458);
or U4848 (N_4848,In_581,In_893);
and U4849 (N_4849,In_249,In_44);
nor U4850 (N_4850,In_641,In_729);
or U4851 (N_4851,In_950,In_755);
or U4852 (N_4852,In_902,In_97);
nand U4853 (N_4853,In_219,In_691);
nand U4854 (N_4854,In_530,In_40);
nor U4855 (N_4855,In_408,In_868);
nand U4856 (N_4856,In_80,In_958);
or U4857 (N_4857,In_871,In_774);
or U4858 (N_4858,In_573,In_21);
nand U4859 (N_4859,In_453,In_617);
nand U4860 (N_4860,In_315,In_954);
and U4861 (N_4861,In_113,In_722);
and U4862 (N_4862,In_326,In_738);
or U4863 (N_4863,In_520,In_820);
nand U4864 (N_4864,In_49,In_256);
or U4865 (N_4865,In_287,In_276);
nand U4866 (N_4866,In_978,In_165);
or U4867 (N_4867,In_649,In_513);
or U4868 (N_4868,In_282,In_507);
nor U4869 (N_4869,In_307,In_221);
nor U4870 (N_4870,In_208,In_155);
nand U4871 (N_4871,In_516,In_143);
nor U4872 (N_4872,In_369,In_179);
nand U4873 (N_4873,In_369,In_311);
nor U4874 (N_4874,In_156,In_900);
xnor U4875 (N_4875,In_633,In_919);
or U4876 (N_4876,In_25,In_73);
nor U4877 (N_4877,In_584,In_22);
nand U4878 (N_4878,In_432,In_486);
or U4879 (N_4879,In_684,In_311);
nor U4880 (N_4880,In_148,In_185);
or U4881 (N_4881,In_218,In_231);
nor U4882 (N_4882,In_360,In_55);
nor U4883 (N_4883,In_127,In_828);
xnor U4884 (N_4884,In_444,In_681);
nor U4885 (N_4885,In_213,In_622);
nand U4886 (N_4886,In_15,In_402);
and U4887 (N_4887,In_602,In_776);
nor U4888 (N_4888,In_992,In_978);
and U4889 (N_4889,In_742,In_560);
xnor U4890 (N_4890,In_722,In_646);
xor U4891 (N_4891,In_940,In_733);
and U4892 (N_4892,In_969,In_186);
and U4893 (N_4893,In_681,In_412);
and U4894 (N_4894,In_621,In_218);
nand U4895 (N_4895,In_820,In_236);
nor U4896 (N_4896,In_412,In_306);
nand U4897 (N_4897,In_84,In_981);
xnor U4898 (N_4898,In_443,In_566);
and U4899 (N_4899,In_581,In_605);
xor U4900 (N_4900,In_531,In_825);
and U4901 (N_4901,In_339,In_226);
nor U4902 (N_4902,In_631,In_26);
nand U4903 (N_4903,In_650,In_442);
nor U4904 (N_4904,In_184,In_694);
xor U4905 (N_4905,In_922,In_453);
nand U4906 (N_4906,In_543,In_661);
nand U4907 (N_4907,In_637,In_271);
and U4908 (N_4908,In_89,In_184);
and U4909 (N_4909,In_320,In_441);
nor U4910 (N_4910,In_123,In_677);
and U4911 (N_4911,In_877,In_636);
and U4912 (N_4912,In_332,In_912);
or U4913 (N_4913,In_364,In_141);
xnor U4914 (N_4914,In_410,In_996);
nor U4915 (N_4915,In_948,In_521);
xor U4916 (N_4916,In_660,In_135);
nand U4917 (N_4917,In_217,In_958);
or U4918 (N_4918,In_159,In_828);
and U4919 (N_4919,In_701,In_31);
xor U4920 (N_4920,In_8,In_861);
nand U4921 (N_4921,In_621,In_187);
or U4922 (N_4922,In_385,In_762);
and U4923 (N_4923,In_886,In_645);
nand U4924 (N_4924,In_294,In_148);
nor U4925 (N_4925,In_13,In_97);
xnor U4926 (N_4926,In_596,In_38);
nand U4927 (N_4927,In_808,In_920);
nand U4928 (N_4928,In_941,In_402);
nand U4929 (N_4929,In_26,In_163);
xor U4930 (N_4930,In_541,In_901);
or U4931 (N_4931,In_639,In_905);
nand U4932 (N_4932,In_138,In_422);
and U4933 (N_4933,In_994,In_283);
nand U4934 (N_4934,In_288,In_473);
nand U4935 (N_4935,In_467,In_520);
or U4936 (N_4936,In_604,In_511);
nor U4937 (N_4937,In_878,In_443);
and U4938 (N_4938,In_262,In_397);
nand U4939 (N_4939,In_489,In_987);
nand U4940 (N_4940,In_804,In_853);
nor U4941 (N_4941,In_28,In_831);
nor U4942 (N_4942,In_50,In_658);
nand U4943 (N_4943,In_501,In_198);
or U4944 (N_4944,In_959,In_955);
xnor U4945 (N_4945,In_94,In_46);
nand U4946 (N_4946,In_349,In_579);
xnor U4947 (N_4947,In_231,In_853);
nand U4948 (N_4948,In_481,In_760);
nor U4949 (N_4949,In_511,In_179);
or U4950 (N_4950,In_632,In_85);
xor U4951 (N_4951,In_313,In_283);
or U4952 (N_4952,In_991,In_562);
nor U4953 (N_4953,In_177,In_534);
nor U4954 (N_4954,In_890,In_285);
nand U4955 (N_4955,In_756,In_207);
and U4956 (N_4956,In_750,In_383);
xnor U4957 (N_4957,In_892,In_239);
nand U4958 (N_4958,In_201,In_298);
and U4959 (N_4959,In_76,In_545);
nor U4960 (N_4960,In_972,In_957);
nor U4961 (N_4961,In_783,In_637);
xor U4962 (N_4962,In_412,In_745);
nor U4963 (N_4963,In_409,In_533);
or U4964 (N_4964,In_958,In_825);
and U4965 (N_4965,In_393,In_869);
nand U4966 (N_4966,In_44,In_999);
and U4967 (N_4967,In_883,In_276);
xnor U4968 (N_4968,In_543,In_937);
nor U4969 (N_4969,In_332,In_361);
or U4970 (N_4970,In_145,In_176);
nor U4971 (N_4971,In_618,In_760);
and U4972 (N_4972,In_966,In_104);
xor U4973 (N_4973,In_837,In_675);
xor U4974 (N_4974,In_367,In_947);
or U4975 (N_4975,In_746,In_132);
xor U4976 (N_4976,In_425,In_201);
or U4977 (N_4977,In_258,In_720);
or U4978 (N_4978,In_308,In_399);
nor U4979 (N_4979,In_18,In_107);
or U4980 (N_4980,In_264,In_740);
xor U4981 (N_4981,In_14,In_987);
nor U4982 (N_4982,In_62,In_958);
or U4983 (N_4983,In_918,In_351);
or U4984 (N_4984,In_2,In_508);
and U4985 (N_4985,In_718,In_301);
nand U4986 (N_4986,In_33,In_750);
or U4987 (N_4987,In_322,In_63);
and U4988 (N_4988,In_984,In_212);
or U4989 (N_4989,In_362,In_530);
nor U4990 (N_4990,In_28,In_670);
nand U4991 (N_4991,In_656,In_137);
and U4992 (N_4992,In_45,In_818);
or U4993 (N_4993,In_218,In_908);
and U4994 (N_4994,In_947,In_350);
nand U4995 (N_4995,In_143,In_167);
nor U4996 (N_4996,In_638,In_766);
nand U4997 (N_4997,In_813,In_302);
xor U4998 (N_4998,In_860,In_79);
xnor U4999 (N_4999,In_902,In_905);
or U5000 (N_5000,N_1291,N_3273);
or U5001 (N_5001,N_4818,N_3980);
nor U5002 (N_5002,N_3237,N_1192);
xor U5003 (N_5003,N_1882,N_2880);
nand U5004 (N_5004,N_4025,N_2178);
nand U5005 (N_5005,N_1897,N_4766);
and U5006 (N_5006,N_165,N_3061);
nand U5007 (N_5007,N_1797,N_431);
xnor U5008 (N_5008,N_4049,N_99);
xor U5009 (N_5009,N_3462,N_1979);
nor U5010 (N_5010,N_3320,N_3391);
nand U5011 (N_5011,N_2643,N_241);
or U5012 (N_5012,N_2105,N_2249);
nor U5013 (N_5013,N_2440,N_1472);
and U5014 (N_5014,N_3553,N_1095);
and U5015 (N_5015,N_2333,N_2430);
nor U5016 (N_5016,N_2388,N_1776);
or U5017 (N_5017,N_2138,N_203);
nor U5018 (N_5018,N_600,N_2399);
or U5019 (N_5019,N_2513,N_3737);
and U5020 (N_5020,N_1043,N_3685);
xnor U5021 (N_5021,N_1287,N_4703);
or U5022 (N_5022,N_3545,N_3808);
and U5023 (N_5023,N_4753,N_4739);
xor U5024 (N_5024,N_4999,N_3247);
nand U5025 (N_5025,N_3427,N_4849);
or U5026 (N_5026,N_1099,N_153);
nor U5027 (N_5027,N_2370,N_4988);
and U5028 (N_5028,N_4265,N_4691);
and U5029 (N_5029,N_1314,N_3281);
and U5030 (N_5030,N_3001,N_4706);
and U5031 (N_5031,N_4641,N_2039);
or U5032 (N_5032,N_229,N_69);
nor U5033 (N_5033,N_4722,N_1117);
xnor U5034 (N_5034,N_1673,N_3824);
nand U5035 (N_5035,N_874,N_4890);
and U5036 (N_5036,N_1345,N_983);
nor U5037 (N_5037,N_3752,N_3084);
nor U5038 (N_5038,N_2466,N_3866);
or U5039 (N_5039,N_2784,N_4008);
nor U5040 (N_5040,N_4041,N_2207);
nor U5041 (N_5041,N_1297,N_455);
and U5042 (N_5042,N_1143,N_2571);
nand U5043 (N_5043,N_4925,N_1865);
nand U5044 (N_5044,N_307,N_638);
or U5045 (N_5045,N_3726,N_48);
xnor U5046 (N_5046,N_275,N_2248);
and U5047 (N_5047,N_1970,N_1953);
or U5048 (N_5048,N_4102,N_4669);
nor U5049 (N_5049,N_1129,N_2698);
xnor U5050 (N_5050,N_3079,N_1877);
or U5051 (N_5051,N_4770,N_3658);
nand U5052 (N_5052,N_4362,N_4021);
xnor U5053 (N_5053,N_2777,N_38);
and U5054 (N_5054,N_102,N_1694);
and U5055 (N_5055,N_2195,N_1597);
or U5056 (N_5056,N_2739,N_1434);
and U5057 (N_5057,N_2040,N_2840);
and U5058 (N_5058,N_3935,N_1590);
nand U5059 (N_5059,N_3598,N_18);
xnor U5060 (N_5060,N_2812,N_4484);
or U5061 (N_5061,N_1335,N_3385);
nand U5062 (N_5062,N_2584,N_1674);
nor U5063 (N_5063,N_2581,N_1620);
xor U5064 (N_5064,N_1150,N_793);
and U5065 (N_5065,N_296,N_3314);
nand U5066 (N_5066,N_2186,N_3625);
nor U5067 (N_5067,N_2223,N_1672);
xor U5068 (N_5068,N_2029,N_3008);
nand U5069 (N_5069,N_3104,N_847);
xor U5070 (N_5070,N_1457,N_4120);
or U5071 (N_5071,N_986,N_1549);
and U5072 (N_5072,N_42,N_1097);
nand U5073 (N_5073,N_1758,N_3312);
xor U5074 (N_5074,N_4633,N_4570);
nand U5075 (N_5075,N_4915,N_2727);
xnor U5076 (N_5076,N_1699,N_3515);
or U5077 (N_5077,N_4168,N_2920);
nor U5078 (N_5078,N_1679,N_4461);
and U5079 (N_5079,N_3188,N_1578);
or U5080 (N_5080,N_536,N_1639);
nand U5081 (N_5081,N_4400,N_2163);
or U5082 (N_5082,N_2256,N_2637);
or U5083 (N_5083,N_2569,N_4687);
or U5084 (N_5084,N_3843,N_1772);
or U5085 (N_5085,N_4199,N_59);
nor U5086 (N_5086,N_3292,N_4488);
or U5087 (N_5087,N_2200,N_2603);
nand U5088 (N_5088,N_1357,N_292);
nand U5089 (N_5089,N_85,N_794);
and U5090 (N_5090,N_1016,N_255);
xnor U5091 (N_5091,N_4037,N_50);
xor U5092 (N_5092,N_2108,N_3776);
nor U5093 (N_5093,N_4868,N_3175);
and U5094 (N_5094,N_4552,N_2913);
xnor U5095 (N_5095,N_2734,N_3213);
nand U5096 (N_5096,N_304,N_2789);
nor U5097 (N_5097,N_988,N_1141);
or U5098 (N_5098,N_653,N_3123);
and U5099 (N_5099,N_212,N_3224);
and U5100 (N_5100,N_1126,N_1375);
nand U5101 (N_5101,N_3828,N_4177);
xnor U5102 (N_5102,N_795,N_4981);
and U5103 (N_5103,N_439,N_4819);
nand U5104 (N_5104,N_232,N_116);
or U5105 (N_5105,N_4123,N_3634);
nand U5106 (N_5106,N_1596,N_4656);
xnor U5107 (N_5107,N_963,N_4432);
nor U5108 (N_5108,N_3823,N_4824);
nor U5109 (N_5109,N_502,N_4986);
nor U5110 (N_5110,N_4347,N_4939);
nand U5111 (N_5111,N_956,N_1523);
and U5112 (N_5112,N_4697,N_666);
nand U5113 (N_5113,N_1380,N_1256);
nor U5114 (N_5114,N_492,N_1977);
nand U5115 (N_5115,N_4124,N_2180);
xor U5116 (N_5116,N_277,N_2422);
xor U5117 (N_5117,N_194,N_4348);
nand U5118 (N_5118,N_4479,N_444);
nand U5119 (N_5119,N_2053,N_3921);
or U5120 (N_5120,N_4627,N_1064);
or U5121 (N_5121,N_1366,N_4834);
nor U5122 (N_5122,N_3925,N_3420);
nand U5123 (N_5123,N_2374,N_3989);
and U5124 (N_5124,N_806,N_1988);
or U5125 (N_5125,N_1429,N_1969);
xor U5126 (N_5126,N_4052,N_625);
nand U5127 (N_5127,N_3034,N_1248);
or U5128 (N_5128,N_3234,N_122);
nor U5129 (N_5129,N_4243,N_1209);
xnor U5130 (N_5130,N_4022,N_3452);
and U5131 (N_5131,N_3097,N_3495);
and U5132 (N_5132,N_3262,N_2626);
xor U5133 (N_5133,N_2693,N_2470);
nor U5134 (N_5134,N_1516,N_1885);
or U5135 (N_5135,N_3183,N_993);
xnor U5136 (N_5136,N_2315,N_4401);
and U5137 (N_5137,N_3855,N_1640);
nand U5138 (N_5138,N_2420,N_3663);
or U5139 (N_5139,N_1773,N_1086);
xor U5140 (N_5140,N_2051,N_4260);
or U5141 (N_5141,N_2744,N_4816);
or U5142 (N_5142,N_4114,N_1455);
xor U5143 (N_5143,N_2780,N_937);
nand U5144 (N_5144,N_1255,N_3293);
or U5145 (N_5145,N_972,N_97);
xor U5146 (N_5146,N_3159,N_4944);
or U5147 (N_5147,N_282,N_2118);
nand U5148 (N_5148,N_1581,N_1683);
nor U5149 (N_5149,N_907,N_769);
and U5150 (N_5150,N_4178,N_4334);
xnor U5151 (N_5151,N_2402,N_612);
xnor U5152 (N_5152,N_2953,N_4154);
xor U5153 (N_5153,N_4101,N_1187);
or U5154 (N_5154,N_4763,N_737);
and U5155 (N_5155,N_704,N_2891);
nor U5156 (N_5156,N_728,N_204);
and U5157 (N_5157,N_2445,N_4174);
nor U5158 (N_5158,N_1338,N_1042);
xor U5159 (N_5159,N_4920,N_3903);
or U5160 (N_5160,N_1253,N_1689);
nand U5161 (N_5161,N_4899,N_3116);
nand U5162 (N_5162,N_350,N_1480);
and U5163 (N_5163,N_199,N_4665);
xnor U5164 (N_5164,N_4599,N_2621);
xnor U5165 (N_5165,N_1051,N_3103);
nand U5166 (N_5166,N_3645,N_2412);
nand U5167 (N_5167,N_3268,N_2671);
and U5168 (N_5168,N_1591,N_3538);
xnor U5169 (N_5169,N_4952,N_1200);
nor U5170 (N_5170,N_4426,N_683);
nand U5171 (N_5171,N_4853,N_2725);
nor U5172 (N_5172,N_338,N_1738);
nor U5173 (N_5173,N_2524,N_1054);
nor U5174 (N_5174,N_19,N_3200);
and U5175 (N_5175,N_4166,N_2935);
or U5176 (N_5176,N_2602,N_3860);
and U5177 (N_5177,N_4056,N_339);
xnor U5178 (N_5178,N_713,N_1971);
nand U5179 (N_5179,N_897,N_4652);
or U5180 (N_5180,N_2850,N_2799);
nand U5181 (N_5181,N_1462,N_3263);
nand U5182 (N_5182,N_2548,N_3334);
or U5183 (N_5183,N_2993,N_3599);
xnor U5184 (N_5184,N_4924,N_2157);
xor U5185 (N_5185,N_55,N_497);
and U5186 (N_5186,N_4647,N_4233);
nor U5187 (N_5187,N_1404,N_3690);
nor U5188 (N_5188,N_2352,N_1482);
nand U5189 (N_5189,N_2095,N_4678);
or U5190 (N_5190,N_1374,N_2427);
nor U5191 (N_5191,N_1489,N_3751);
xnor U5192 (N_5192,N_4090,N_685);
nand U5193 (N_5193,N_133,N_4989);
and U5194 (N_5194,N_3413,N_3210);
and U5195 (N_5195,N_3446,N_2939);
nor U5196 (N_5196,N_2101,N_2944);
nor U5197 (N_5197,N_1484,N_4745);
nand U5198 (N_5198,N_3643,N_4087);
and U5199 (N_5199,N_2235,N_2484);
xnor U5200 (N_5200,N_2908,N_443);
and U5201 (N_5201,N_1280,N_2984);
nor U5202 (N_5202,N_2194,N_1589);
or U5203 (N_5203,N_4878,N_2305);
nor U5204 (N_5204,N_1166,N_1759);
nor U5205 (N_5205,N_1196,N_826);
nor U5206 (N_5206,N_821,N_835);
xor U5207 (N_5207,N_3622,N_4567);
or U5208 (N_5208,N_920,N_815);
and U5209 (N_5209,N_1492,N_1277);
nor U5210 (N_5210,N_4062,N_4274);
and U5211 (N_5211,N_4940,N_2736);
nor U5212 (N_5212,N_871,N_3729);
xor U5213 (N_5213,N_1083,N_1440);
or U5214 (N_5214,N_3876,N_4425);
and U5215 (N_5215,N_2755,N_3612);
xnor U5216 (N_5216,N_2819,N_488);
nor U5217 (N_5217,N_4074,N_73);
and U5218 (N_5218,N_4538,N_4030);
or U5219 (N_5219,N_3441,N_33);
xor U5220 (N_5220,N_4828,N_4874);
nor U5221 (N_5221,N_184,N_3099);
xor U5222 (N_5222,N_2868,N_3152);
nor U5223 (N_5223,N_1747,N_4203);
or U5224 (N_5224,N_4649,N_127);
or U5225 (N_5225,N_3057,N_481);
or U5226 (N_5226,N_1339,N_1313);
nor U5227 (N_5227,N_1245,N_4359);
xor U5228 (N_5228,N_3535,N_4880);
and U5229 (N_5229,N_7,N_4344);
nor U5230 (N_5230,N_4463,N_4772);
or U5231 (N_5231,N_1461,N_4841);
nor U5232 (N_5232,N_4371,N_4787);
nor U5233 (N_5233,N_346,N_503);
and U5234 (N_5234,N_4974,N_2561);
and U5235 (N_5235,N_4526,N_3684);
or U5236 (N_5236,N_2366,N_1323);
nand U5237 (N_5237,N_4280,N_3907);
nand U5238 (N_5238,N_4388,N_1714);
and U5239 (N_5239,N_1664,N_3922);
xnor U5240 (N_5240,N_4158,N_2469);
xnor U5241 (N_5241,N_80,N_2816);
xor U5242 (N_5242,N_1055,N_1132);
or U5243 (N_5243,N_2444,N_1331);
xor U5244 (N_5244,N_3351,N_53);
or U5245 (N_5245,N_1789,N_2729);
or U5246 (N_5246,N_2049,N_3037);
xnor U5247 (N_5247,N_4176,N_1647);
xor U5248 (N_5248,N_2684,N_3489);
xor U5249 (N_5249,N_3023,N_4593);
or U5250 (N_5250,N_2462,N_4609);
xor U5251 (N_5251,N_1023,N_4934);
nor U5252 (N_5252,N_875,N_1002);
nor U5253 (N_5253,N_1562,N_598);
or U5254 (N_5254,N_3504,N_2222);
or U5255 (N_5255,N_1539,N_2027);
nor U5256 (N_5256,N_804,N_2226);
nand U5257 (N_5257,N_858,N_1751);
or U5258 (N_5258,N_268,N_2865);
and U5259 (N_5259,N_79,N_1537);
or U5260 (N_5260,N_1564,N_2954);
or U5261 (N_5261,N_1641,N_3376);
nor U5262 (N_5262,N_2190,N_423);
or U5263 (N_5263,N_1654,N_4616);
xor U5264 (N_5264,N_1935,N_1949);
or U5265 (N_5265,N_714,N_1299);
nand U5266 (N_5266,N_569,N_2710);
and U5267 (N_5267,N_3290,N_3635);
nor U5268 (N_5268,N_4169,N_2086);
nand U5269 (N_5269,N_2785,N_4962);
nor U5270 (N_5270,N_4222,N_388);
or U5271 (N_5271,N_4556,N_1556);
and U5272 (N_5272,N_2589,N_1534);
and U5273 (N_5273,N_4096,N_3388);
nor U5274 (N_5274,N_4713,N_4332);
nor U5275 (N_5275,N_3770,N_3328);
or U5276 (N_5276,N_992,N_4417);
nand U5277 (N_5277,N_1026,N_2460);
nand U5278 (N_5278,N_3537,N_3680);
nand U5279 (N_5279,N_494,N_2438);
nand U5280 (N_5280,N_294,N_825);
or U5281 (N_5281,N_3275,N_2822);
and U5282 (N_5282,N_4578,N_3570);
nor U5283 (N_5283,N_2692,N_400);
nand U5284 (N_5284,N_3773,N_2308);
xnor U5285 (N_5285,N_2529,N_3558);
nor U5286 (N_5286,N_1835,N_4508);
nand U5287 (N_5287,N_1749,N_1422);
nand U5288 (N_5288,N_3178,N_4572);
xnor U5289 (N_5289,N_911,N_1318);
nand U5290 (N_5290,N_2871,N_3416);
and U5291 (N_5291,N_961,N_558);
or U5292 (N_5292,N_1879,N_3236);
xnor U5293 (N_5293,N_1713,N_915);
nor U5294 (N_5294,N_1621,N_2473);
and U5295 (N_5295,N_2923,N_3755);
nand U5296 (N_5296,N_3594,N_2115);
nor U5297 (N_5297,N_57,N_846);
or U5298 (N_5298,N_745,N_4231);
nor U5299 (N_5299,N_4310,N_4893);
and U5300 (N_5300,N_899,N_865);
xor U5301 (N_5301,N_2081,N_3294);
nor U5302 (N_5302,N_2338,N_3586);
nor U5303 (N_5303,N_4365,N_3045);
xor U5304 (N_5304,N_2225,N_2030);
and U5305 (N_5305,N_2890,N_1329);
or U5306 (N_5306,N_1770,N_3070);
or U5307 (N_5307,N_2910,N_2220);
and U5308 (N_5308,N_3319,N_4554);
and U5309 (N_5309,N_4339,N_1330);
or U5310 (N_5310,N_110,N_58);
nor U5311 (N_5311,N_473,N_4009);
xor U5312 (N_5312,N_1718,N_2770);
xor U5313 (N_5313,N_4564,N_2251);
xnor U5314 (N_5314,N_3662,N_3813);
nor U5315 (N_5315,N_251,N_3472);
xnor U5316 (N_5316,N_2126,N_4643);
nor U5317 (N_5317,N_4854,N_3678);
nand U5318 (N_5318,N_1737,N_4098);
and U5319 (N_5319,N_4821,N_2089);
nor U5320 (N_5320,N_2528,N_4370);
xor U5321 (N_5321,N_3560,N_2535);
and U5322 (N_5322,N_607,N_3355);
xor U5323 (N_5323,N_1409,N_4848);
nor U5324 (N_5324,N_1459,N_1408);
xor U5325 (N_5325,N_4317,N_3246);
xnor U5326 (N_5326,N_4648,N_4683);
xor U5327 (N_5327,N_86,N_3482);
or U5328 (N_5328,N_3068,N_673);
and U5329 (N_5329,N_1981,N_3986);
nor U5330 (N_5330,N_2082,N_4631);
nand U5331 (N_5331,N_1189,N_4437);
or U5332 (N_5332,N_1250,N_1632);
nand U5333 (N_5333,N_4715,N_4885);
and U5334 (N_5334,N_216,N_935);
and U5335 (N_5335,N_3431,N_3932);
or U5336 (N_5336,N_3812,N_873);
xor U5337 (N_5337,N_4596,N_890);
nor U5338 (N_5338,N_4535,N_2236);
nor U5339 (N_5339,N_3888,N_3326);
or U5340 (N_5340,N_2695,N_4246);
nor U5341 (N_5341,N_4137,N_337);
or U5342 (N_5342,N_4950,N_4718);
and U5343 (N_5343,N_4354,N_1225);
or U5344 (N_5344,N_94,N_1553);
xor U5345 (N_5345,N_3258,N_872);
nor U5346 (N_5346,N_4216,N_1940);
xor U5347 (N_5347,N_2351,N_1037);
or U5348 (N_5348,N_2658,N_2015);
nand U5349 (N_5349,N_164,N_3126);
nand U5350 (N_5350,N_2516,N_3050);
nor U5351 (N_5351,N_2281,N_3597);
nor U5352 (N_5352,N_1670,N_4395);
or U5353 (N_5353,N_530,N_1442);
or U5354 (N_5354,N_323,N_2737);
xor U5355 (N_5355,N_4235,N_4394);
xor U5356 (N_5356,N_1242,N_1163);
nand U5357 (N_5357,N_3508,N_3724);
nor U5358 (N_5358,N_1421,N_3802);
and U5359 (N_5359,N_4304,N_3367);
nand U5360 (N_5360,N_2988,N_3566);
or U5361 (N_5361,N_578,N_4086);
nor U5362 (N_5362,N_4660,N_515);
or U5363 (N_5363,N_1697,N_1928);
or U5364 (N_5364,N_4765,N_4855);
or U5365 (N_5365,N_1413,N_3838);
xnor U5366 (N_5366,N_1720,N_2303);
nor U5367 (N_5367,N_1107,N_2512);
or U5368 (N_5368,N_1691,N_3575);
or U5369 (N_5369,N_2002,N_1662);
xor U5370 (N_5370,N_1859,N_1082);
and U5371 (N_5371,N_1198,N_3655);
or U5372 (N_5372,N_1476,N_1659);
nor U5373 (N_5373,N_4071,N_2514);
nand U5374 (N_5374,N_2369,N_1411);
xor U5375 (N_5375,N_3150,N_4415);
xnor U5376 (N_5376,N_1999,N_1114);
or U5377 (N_5377,N_2054,N_818);
and U5378 (N_5378,N_386,N_3248);
xor U5379 (N_5379,N_1398,N_3026);
and U5380 (N_5380,N_3734,N_348);
nand U5381 (N_5381,N_1045,N_4559);
nand U5382 (N_5382,N_2390,N_313);
nor U5383 (N_5383,N_1734,N_930);
xor U5384 (N_5384,N_3691,N_4283);
or U5385 (N_5385,N_4887,N_4613);
nand U5386 (N_5386,N_2999,N_3249);
xor U5387 (N_5387,N_3133,N_1816);
nor U5388 (N_5388,N_3820,N_406);
nor U5389 (N_5389,N_1001,N_1812);
and U5390 (N_5390,N_4423,N_1258);
xor U5391 (N_5391,N_4585,N_1041);
and U5392 (N_5392,N_1385,N_4477);
or U5393 (N_5393,N_3278,N_1505);
nand U5394 (N_5394,N_3603,N_4793);
nor U5395 (N_5395,N_1623,N_4094);
or U5396 (N_5396,N_1552,N_2878);
or U5397 (N_5397,N_3227,N_131);
nor U5398 (N_5398,N_3931,N_512);
xor U5399 (N_5399,N_4852,N_2895);
and U5400 (N_5400,N_1066,N_2102);
nand U5401 (N_5401,N_1487,N_144);
or U5402 (N_5402,N_3804,N_487);
or U5403 (N_5403,N_4290,N_324);
or U5404 (N_5404,N_1658,N_2097);
nor U5405 (N_5405,N_175,N_4193);
and U5406 (N_5406,N_1243,N_3785);
nand U5407 (N_5407,N_924,N_1467);
nand U5408 (N_5408,N_4994,N_3193);
xor U5409 (N_5409,N_2047,N_3827);
xor U5410 (N_5410,N_2916,N_799);
nand U5411 (N_5411,N_3623,N_2213);
and U5412 (N_5412,N_4931,N_2722);
nand U5413 (N_5413,N_1049,N_4412);
xnor U5414 (N_5414,N_3402,N_800);
nand U5415 (N_5415,N_1538,N_4253);
nand U5416 (N_5416,N_531,N_2555);
nand U5417 (N_5417,N_3883,N_4972);
and U5418 (N_5418,N_2656,N_2084);
nor U5419 (N_5419,N_1343,N_3630);
xnor U5420 (N_5420,N_115,N_4615);
xor U5421 (N_5421,N_828,N_3983);
nor U5422 (N_5422,N_4746,N_422);
or U5423 (N_5423,N_1894,N_2879);
or U5424 (N_5424,N_4099,N_1656);
or U5425 (N_5425,N_3170,N_3803);
or U5426 (N_5426,N_1916,N_4330);
xnor U5427 (N_5427,N_2863,N_3805);
or U5428 (N_5428,N_1602,N_1072);
nor U5429 (N_5429,N_1436,N_4001);
and U5430 (N_5430,N_4277,N_2442);
or U5431 (N_5431,N_4392,N_4340);
and U5432 (N_5432,N_1282,N_687);
or U5433 (N_5433,N_308,N_3775);
and U5434 (N_5434,N_3845,N_2218);
nor U5435 (N_5435,N_2751,N_2010);
xnor U5436 (N_5436,N_4055,N_3701);
nand U5437 (N_5437,N_3915,N_1262);
or U5438 (N_5438,N_2848,N_2279);
and U5439 (N_5439,N_256,N_3144);
nand U5440 (N_5440,N_2059,N_2826);
xnor U5441 (N_5441,N_4659,N_2741);
nand U5442 (N_5442,N_3090,N_1349);
or U5443 (N_5443,N_2009,N_844);
and U5444 (N_5444,N_2608,N_228);
xnor U5445 (N_5445,N_4985,N_995);
and U5446 (N_5446,N_3944,N_3530);
nand U5447 (N_5447,N_1238,N_4449);
nor U5448 (N_5448,N_4390,N_676);
nand U5449 (N_5449,N_4503,N_3763);
nor U5450 (N_5450,N_1428,N_4429);
xor U5451 (N_5451,N_3963,N_1908);
xor U5452 (N_5452,N_542,N_3797);
or U5453 (N_5453,N_398,N_2532);
or U5454 (N_5454,N_2099,N_189);
and U5455 (N_5455,N_3578,N_29);
or U5456 (N_5456,N_3880,N_2978);
xor U5457 (N_5457,N_4953,N_4784);
or U5458 (N_5458,N_1279,N_66);
and U5459 (N_5459,N_1730,N_2792);
or U5460 (N_5460,N_1934,N_271);
xnor U5461 (N_5461,N_2992,N_1774);
xor U5462 (N_5462,N_2302,N_3588);
nor U5463 (N_5463,N_4043,N_668);
and U5464 (N_5464,N_1047,N_3517);
nor U5465 (N_5465,N_546,N_3958);
xor U5466 (N_5466,N_4398,N_4551);
nand U5467 (N_5467,N_2318,N_4811);
and U5468 (N_5468,N_582,N_20);
and U5469 (N_5469,N_1191,N_4278);
or U5470 (N_5470,N_1805,N_2133);
nor U5471 (N_5471,N_3716,N_4018);
and U5472 (N_5472,N_2064,N_2856);
and U5473 (N_5473,N_770,N_529);
nand U5474 (N_5474,N_32,N_362);
nand U5475 (N_5475,N_405,N_124);
nor U5476 (N_5476,N_1322,N_3536);
nor U5477 (N_5477,N_4847,N_4605);
nand U5478 (N_5478,N_4312,N_2011);
xor U5479 (N_5479,N_2846,N_3540);
or U5480 (N_5480,N_343,N_1557);
nor U5481 (N_5481,N_4845,N_1864);
xor U5482 (N_5482,N_722,N_250);
nand U5483 (N_5483,N_2129,N_3723);
or U5484 (N_5484,N_197,N_4007);
nor U5485 (N_5485,N_2735,N_2014);
nand U5486 (N_5486,N_2437,N_111);
xor U5487 (N_5487,N_3574,N_2313);
nand U5488 (N_5488,N_1862,N_764);
and U5489 (N_5489,N_1680,N_3185);
xnor U5490 (N_5490,N_3005,N_4827);
nand U5491 (N_5491,N_568,N_1050);
nand U5492 (N_5492,N_1980,N_1405);
and U5493 (N_5493,N_1007,N_877);
or U5494 (N_5494,N_4993,N_4133);
or U5495 (N_5495,N_2344,N_2173);
or U5496 (N_5496,N_1321,N_654);
xor U5497 (N_5497,N_3587,N_3719);
or U5498 (N_5498,N_4205,N_715);
and U5499 (N_5499,N_4015,N_1365);
nand U5500 (N_5500,N_2545,N_4031);
nor U5501 (N_5501,N_2509,N_146);
and U5502 (N_5502,N_1160,N_12);
or U5503 (N_5503,N_3329,N_1604);
nor U5504 (N_5504,N_4217,N_2864);
or U5505 (N_5505,N_2031,N_4714);
xnor U5506 (N_5506,N_120,N_2901);
xor U5507 (N_5507,N_1412,N_60);
and U5508 (N_5508,N_1296,N_154);
or U5509 (N_5509,N_1808,N_1815);
or U5510 (N_5510,N_1838,N_2345);
and U5511 (N_5511,N_2636,N_1918);
or U5512 (N_5512,N_3352,N_3861);
nand U5513 (N_5513,N_1,N_269);
or U5514 (N_5514,N_2424,N_3418);
xnor U5515 (N_5515,N_1902,N_1269);
nor U5516 (N_5516,N_3182,N_134);
or U5517 (N_5517,N_2867,N_4409);
or U5518 (N_5518,N_4575,N_1520);
or U5519 (N_5519,N_2359,N_4012);
or U5520 (N_5520,N_4060,N_247);
or U5521 (N_5521,N_4482,N_4269);
or U5522 (N_5522,N_1402,N_3672);
xnor U5523 (N_5523,N_869,N_1893);
xnor U5524 (N_5524,N_4271,N_2843);
nor U5525 (N_5525,N_2682,N_1362);
and U5526 (N_5526,N_2808,N_4710);
xnor U5527 (N_5527,N_4014,N_200);
or U5528 (N_5528,N_4859,N_615);
and U5529 (N_5529,N_3571,N_3897);
nand U5530 (N_5530,N_4161,N_2021);
xnor U5531 (N_5531,N_3604,N_922);
xor U5532 (N_5532,N_1850,N_3009);
nor U5533 (N_5533,N_1821,N_2058);
nor U5534 (N_5534,N_2111,N_1989);
and U5535 (N_5535,N_2726,N_3736);
nand U5536 (N_5536,N_2151,N_2585);
nand U5537 (N_5537,N_4469,N_1401);
xor U5538 (N_5538,N_4767,N_4964);
nand U5539 (N_5539,N_4755,N_1216);
xnor U5540 (N_5540,N_3284,N_91);
nand U5541 (N_5541,N_4291,N_466);
xnor U5542 (N_5542,N_789,N_1876);
nand U5543 (N_5543,N_4236,N_2093);
or U5544 (N_5544,N_2092,N_694);
nor U5545 (N_5545,N_3215,N_2250);
nand U5546 (N_5546,N_89,N_1400);
nand U5547 (N_5547,N_923,N_4528);
or U5548 (N_5548,N_2900,N_3965);
and U5549 (N_5549,N_773,N_246);
or U5550 (N_5550,N_2884,N_2873);
and U5551 (N_5551,N_1495,N_2216);
and U5552 (N_5552,N_3656,N_4351);
nor U5553 (N_5553,N_1240,N_297);
or U5554 (N_5554,N_1883,N_4282);
xor U5555 (N_5555,N_3131,N_2685);
nand U5556 (N_5556,N_2057,N_1675);
and U5557 (N_5557,N_1426,N_2266);
xor U5558 (N_5558,N_3607,N_3399);
or U5559 (N_5559,N_82,N_565);
xnor U5560 (N_5560,N_845,N_2905);
nor U5561 (N_5561,N_2796,N_1543);
nand U5562 (N_5562,N_757,N_306);
and U5563 (N_5563,N_4932,N_1194);
nand U5564 (N_5564,N_3031,N_4998);
nor U5565 (N_5565,N_948,N_30);
nand U5566 (N_5566,N_2934,N_1769);
and U5567 (N_5567,N_4237,N_4629);
or U5568 (N_5568,N_3145,N_2542);
xor U5569 (N_5569,N_2921,N_4825);
xor U5570 (N_5570,N_2673,N_4764);
nand U5571 (N_5571,N_4884,N_3591);
or U5572 (N_5572,N_1660,N_1491);
and U5573 (N_5573,N_4688,N_2500);
nand U5574 (N_5574,N_3065,N_1878);
and U5575 (N_5575,N_2805,N_1572);
or U5576 (N_5576,N_2273,N_4413);
nor U5577 (N_5577,N_474,N_4289);
nor U5578 (N_5578,N_2615,N_3710);
or U5579 (N_5579,N_1498,N_905);
nor U5580 (N_5580,N_4979,N_1566);
or U5581 (N_5581,N_475,N_4111);
and U5582 (N_5582,N_3373,N_419);
or U5583 (N_5583,N_3956,N_514);
and U5584 (N_5584,N_2598,N_461);
nand U5585 (N_5585,N_262,N_287);
nor U5586 (N_5586,N_888,N_3557);
and U5587 (N_5587,N_2405,N_2264);
nand U5588 (N_5588,N_2620,N_4287);
or U5589 (N_5589,N_3702,N_1568);
nand U5590 (N_5590,N_4574,N_3287);
or U5591 (N_5591,N_1391,N_4214);
nand U5592 (N_5592,N_4628,N_4948);
or U5593 (N_5593,N_4518,N_1706);
nor U5594 (N_5594,N_2122,N_662);
or U5595 (N_5595,N_4107,N_3317);
nand U5596 (N_5596,N_768,N_507);
nand U5597 (N_5597,N_1127,N_2986);
nor U5598 (N_5598,N_3696,N_4314);
and U5599 (N_5599,N_3345,N_2558);
and U5600 (N_5600,N_4150,N_1587);
nor U5601 (N_5601,N_1728,N_604);
nor U5602 (N_5602,N_649,N_4113);
nor U5603 (N_5603,N_2310,N_1358);
nand U5604 (N_5604,N_3467,N_1507);
nor U5605 (N_5605,N_1056,N_4238);
xnor U5606 (N_5606,N_796,N_1425);
or U5607 (N_5607,N_3554,N_4076);
nor U5608 (N_5608,N_1096,N_2373);
nand U5609 (N_5609,N_736,N_2183);
xor U5610 (N_5610,N_541,N_1519);
nand U5611 (N_5611,N_4259,N_3670);
and U5612 (N_5612,N_787,N_1527);
or U5613 (N_5613,N_3444,N_4553);
or U5614 (N_5614,N_1506,N_3782);
nand U5615 (N_5615,N_4396,N_1028);
or U5616 (N_5616,N_3142,N_205);
nand U5617 (N_5617,N_1197,N_2605);
and U5618 (N_5618,N_2679,N_1532);
or U5619 (N_5619,N_3456,N_3493);
xnor U5620 (N_5620,N_622,N_3942);
and U5621 (N_5621,N_726,N_1195);
nor U5622 (N_5622,N_3490,N_1283);
xnor U5623 (N_5623,N_2940,N_1618);
xnor U5624 (N_5624,N_218,N_1524);
nand U5625 (N_5625,N_3245,N_3957);
and U5626 (N_5626,N_4293,N_1497);
xnor U5627 (N_5627,N_564,N_4519);
nand U5628 (N_5628,N_4016,N_4065);
and U5629 (N_5629,N_1724,N_1965);
xnor U5630 (N_5630,N_4721,N_2973);
or U5631 (N_5631,N_3583,N_3135);
or U5632 (N_5632,N_1525,N_2724);
nor U5633 (N_5633,N_594,N_1185);
xnor U5634 (N_5634,N_857,N_3020);
and U5635 (N_5635,N_2543,N_2076);
or U5636 (N_5636,N_3510,N_3503);
xor U5637 (N_5637,N_224,N_2203);
nor U5638 (N_5638,N_1541,N_783);
and U5639 (N_5639,N_2866,N_1130);
and U5640 (N_5640,N_2232,N_1254);
nor U5641 (N_5641,N_4345,N_2958);
nor U5642 (N_5642,N_3119,N_1560);
or U5643 (N_5643,N_2455,N_3197);
xor U5644 (N_5644,N_1188,N_2227);
or U5645 (N_5645,N_562,N_3572);
or U5646 (N_5646,N_2008,N_761);
or U5647 (N_5647,N_4638,N_2001);
nor U5648 (N_5648,N_772,N_1567);
xnor U5649 (N_5649,N_2696,N_4769);
nor U5650 (N_5650,N_1237,N_4104);
or U5651 (N_5651,N_3381,N_445);
and U5652 (N_5652,N_361,N_4229);
nand U5653 (N_5653,N_3532,N_1684);
or U5654 (N_5654,N_1705,N_2837);
nand U5655 (N_5655,N_2155,N_3115);
nor U5656 (N_5656,N_3408,N_4850);
and U5657 (N_5657,N_1184,N_2492);
nand U5658 (N_5658,N_2407,N_1698);
xnor U5659 (N_5659,N_3250,N_2297);
xor U5660 (N_5660,N_4781,N_2560);
xor U5661 (N_5661,N_1057,N_4000);
and U5662 (N_5662,N_4813,N_552);
nand U5663 (N_5663,N_4245,N_2291);
nor U5664 (N_5664,N_2075,N_3445);
or U5665 (N_5665,N_2271,N_1460);
nor U5666 (N_5666,N_776,N_3429);
xnor U5667 (N_5667,N_340,N_206);
and U5668 (N_5668,N_1397,N_1158);
nand U5669 (N_5669,N_1605,N_4897);
or U5670 (N_5670,N_1701,N_3271);
and U5671 (N_5671,N_2229,N_1018);
nand U5672 (N_5672,N_1843,N_1307);
nor U5673 (N_5673,N_107,N_1919);
xnor U5674 (N_5674,N_4201,N_2596);
or U5675 (N_5675,N_4682,N_2104);
and U5676 (N_5676,N_3128,N_3220);
or U5677 (N_5677,N_4809,N_2448);
nand U5678 (N_5678,N_2411,N_3730);
or U5679 (N_5679,N_2556,N_1739);
xnor U5680 (N_5680,N_1104,N_3936);
nand U5681 (N_5681,N_2055,N_1351);
nor U5682 (N_5682,N_4379,N_705);
xor U5683 (N_5683,N_4525,N_1822);
nor U5684 (N_5684,N_1201,N_402);
and U5685 (N_5685,N_1655,N_438);
xor U5686 (N_5686,N_4642,N_172);
nor U5687 (N_5687,N_4978,N_1841);
xnor U5688 (N_5688,N_1565,N_3573);
and U5689 (N_5689,N_3675,N_1081);
nor U5690 (N_5690,N_2748,N_4077);
nor U5691 (N_5691,N_1978,N_266);
nand U5692 (N_5692,N_1149,N_3047);
and U5693 (N_5693,N_2818,N_751);
or U5694 (N_5694,N_1077,N_1278);
or U5695 (N_5695,N_2669,N_3509);
or U5696 (N_5696,N_2286,N_2314);
nand U5697 (N_5697,N_3933,N_4044);
xor U5698 (N_5698,N_257,N_4777);
or U5699 (N_5699,N_2224,N_544);
or U5700 (N_5700,N_4509,N_3694);
nand U5701 (N_5701,N_3787,N_24);
or U5702 (N_5702,N_2959,N_363);
nand U5703 (N_5703,N_3689,N_3229);
nand U5704 (N_5704,N_2408,N_2136);
and U5705 (N_5705,N_3872,N_4759);
or U5706 (N_5706,N_4653,N_4296);
nor U5707 (N_5707,N_1575,N_2161);
or U5708 (N_5708,N_4900,N_1456);
or U5709 (N_5709,N_629,N_631);
and U5710 (N_5710,N_1153,N_4576);
or U5711 (N_5711,N_192,N_3158);
xnor U5712 (N_5712,N_2838,N_1790);
xnor U5713 (N_5713,N_295,N_3960);
or U5714 (N_5714,N_1478,N_3608);
nor U5715 (N_5715,N_4862,N_3681);
nand U5716 (N_5716,N_979,N_1806);
nor U5717 (N_5717,N_1926,N_849);
nor U5718 (N_5718,N_1432,N_4219);
nor U5719 (N_5719,N_2974,N_1115);
or U5720 (N_5720,N_4447,N_2246);
nand U5721 (N_5721,N_1295,N_3796);
or U5722 (N_5722,N_749,N_1985);
and U5723 (N_5723,N_2932,N_3046);
and U5724 (N_5724,N_4324,N_1224);
and U5725 (N_5725,N_1383,N_1260);
or U5726 (N_5726,N_326,N_970);
xnor U5727 (N_5727,N_2520,N_3778);
nor U5728 (N_5728,N_78,N_602);
nor U5729 (N_5729,N_3686,N_290);
or U5730 (N_5730,N_2140,N_4725);
nor U5731 (N_5731,N_1831,N_1952);
or U5732 (N_5732,N_3448,N_3688);
xnor U5733 (N_5733,N_3107,N_3995);
nand U5734 (N_5734,N_4611,N_4108);
nand U5735 (N_5735,N_353,N_4548);
xnor U5736 (N_5736,N_1292,N_2576);
or U5737 (N_5737,N_4035,N_1139);
nand U5738 (N_5738,N_334,N_273);
and U5739 (N_5739,N_534,N_3959);
and U5740 (N_5740,N_4473,N_4655);
or U5741 (N_5741,N_2720,N_3928);
or U5742 (N_5742,N_4145,N_3988);
or U5743 (N_5743,N_2125,N_3289);
nor U5744 (N_5744,N_321,N_3266);
nand U5745 (N_5745,N_3323,N_424);
nand U5746 (N_5746,N_4996,N_1069);
nor U5747 (N_5747,N_1494,N_1819);
xnor U5748 (N_5748,N_453,N_173);
nor U5749 (N_5749,N_252,N_1302);
nand U5750 (N_5750,N_4507,N_1199);
nand U5751 (N_5751,N_2915,N_368);
or U5752 (N_5752,N_2026,N_3952);
xor U5753 (N_5753,N_2574,N_3148);
xnor U5754 (N_5754,N_2311,N_1118);
xor U5755 (N_5755,N_2478,N_2718);
and U5756 (N_5756,N_2874,N_3048);
or U5757 (N_5757,N_143,N_1613);
or U5758 (N_5758,N_2247,N_170);
xor U5759 (N_5759,N_4991,N_605);
or U5760 (N_5760,N_4089,N_950);
or U5761 (N_5761,N_3593,N_3971);
xor U5762 (N_5762,N_4795,N_4569);
nor U5763 (N_5763,N_215,N_2197);
or U5764 (N_5764,N_305,N_40);
nor U5765 (N_5765,N_4408,N_358);
xor U5766 (N_5766,N_731,N_3356);
xnor U5767 (N_5767,N_3641,N_426);
and U5768 (N_5768,N_1229,N_2482);
or U5769 (N_5769,N_4303,N_4496);
xnor U5770 (N_5770,N_2502,N_895);
nor U5771 (N_5771,N_2947,N_940);
or U5772 (N_5772,N_1340,N_2061);
and U5773 (N_5773,N_281,N_4520);
or U5774 (N_5774,N_4587,N_606);
xor U5775 (N_5775,N_3998,N_213);
xnor U5776 (N_5776,N_1686,N_2642);
xnor U5777 (N_5777,N_4497,N_1504);
xnor U5778 (N_5778,N_581,N_456);
xnor U5779 (N_5779,N_489,N_978);
or U5780 (N_5780,N_831,N_207);
xor U5781 (N_5781,N_1550,N_3819);
xor U5782 (N_5782,N_2821,N_2208);
nor U5783 (N_5783,N_420,N_76);
and U5784 (N_5784,N_781,N_2395);
xor U5785 (N_5785,N_1887,N_3790);
xnor U5786 (N_5786,N_2019,N_2544);
nor U5787 (N_5787,N_1062,N_535);
or U5788 (N_5788,N_2565,N_2282);
or U5789 (N_5789,N_820,N_1546);
or U5790 (N_5790,N_3837,N_2036);
and U5791 (N_5791,N_1513,N_3793);
or U5792 (N_5792,N_3064,N_2453);
nand U5793 (N_5793,N_2035,N_2889);
or U5794 (N_5794,N_2593,N_123);
xor U5795 (N_5795,N_2259,N_449);
and U5796 (N_5796,N_3253,N_533);
and U5797 (N_5797,N_4170,N_3822);
nor U5798 (N_5798,N_464,N_962);
nor U5799 (N_5799,N_779,N_312);
or U5800 (N_5800,N_3699,N_4485);
xnor U5801 (N_5801,N_2152,N_4679);
nand U5802 (N_5802,N_1270,N_1943);
xnor U5803 (N_5803,N_974,N_3440);
and U5804 (N_5804,N_4748,N_16);
nor U5805 (N_5805,N_771,N_4881);
nand U5806 (N_5806,N_114,N_4374);
nand U5807 (N_5807,N_2701,N_1888);
nor U5808 (N_5808,N_2335,N_2732);
nor U5809 (N_5809,N_2435,N_4095);
or U5810 (N_5810,N_2631,N_3449);
nor U5811 (N_5811,N_4424,N_371);
xnor U5812 (N_5812,N_904,N_230);
nor U5813 (N_5813,N_4754,N_147);
and U5814 (N_5814,N_1619,N_3466);
and U5815 (N_5815,N_4690,N_1616);
or U5816 (N_5816,N_448,N_1290);
and U5817 (N_5817,N_4421,N_601);
xnor U5818 (N_5818,N_2265,N_2188);
or U5819 (N_5819,N_4911,N_1359);
xnor U5820 (N_5820,N_3592,N_603);
and U5821 (N_5821,N_1175,N_4664);
nor U5822 (N_5822,N_2948,N_4523);
or U5823 (N_5823,N_2769,N_2616);
or U5824 (N_5824,N_1555,N_2982);
nor U5825 (N_5825,N_1628,N_3189);
xor U5826 (N_5826,N_523,N_2361);
nand U5827 (N_5827,N_2705,N_3728);
nor U5828 (N_5828,N_730,N_13);
xor U5829 (N_5829,N_3140,N_3704);
or U5830 (N_5830,N_3494,N_945);
nor U5831 (N_5831,N_4476,N_2094);
xnor U5832 (N_5832,N_2624,N_2330);
nor U5833 (N_5833,N_1501,N_633);
xor U5834 (N_5834,N_2504,N_2461);
and U5835 (N_5835,N_1101,N_498);
or U5836 (N_5836,N_903,N_4967);
and U5837 (N_5837,N_2632,N_263);
xor U5838 (N_5838,N_436,N_2416);
xnor U5839 (N_5839,N_957,N_4961);
and U5840 (N_5840,N_1800,N_2159);
xor U5841 (N_5841,N_1914,N_3307);
nor U5842 (N_5842,N_4844,N_4620);
nand U5843 (N_5843,N_289,N_442);
nor U5844 (N_5844,N_2362,N_1388);
xnor U5845 (N_5845,N_3806,N_537);
xnor U5846 (N_5846,N_4011,N_493);
and U5847 (N_5847,N_4912,N_3774);
xnor U5848 (N_5848,N_4050,N_4320);
xnor U5849 (N_5849,N_650,N_1181);
nand U5850 (N_5850,N_646,N_3967);
xor U5851 (N_5851,N_1276,N_1110);
nand U5852 (N_5852,N_1657,N_4316);
nor U5853 (N_5853,N_3760,N_1371);
nand U5854 (N_5854,N_344,N_2674);
nor U5855 (N_5855,N_4093,N_1464);
nor U5856 (N_5856,N_311,N_4357);
or U5857 (N_5857,N_248,N_3007);
nor U5858 (N_5858,N_623,N_2404);
and U5859 (N_5859,N_1353,N_4673);
and U5860 (N_5860,N_2240,N_553);
and U5861 (N_5861,N_1900,N_4393);
and U5862 (N_5862,N_4202,N_3999);
or U5863 (N_5863,N_2583,N_4148);
nor U5864 (N_5864,N_3749,N_1708);
or U5865 (N_5865,N_4760,N_3633);
nor U5866 (N_5866,N_2677,N_2798);
or U5867 (N_5867,N_4990,N_10);
xnor U5868 (N_5868,N_2580,N_1152);
nor U5869 (N_5869,N_2324,N_1813);
and U5870 (N_5870,N_482,N_1445);
nor U5871 (N_5871,N_3567,N_3618);
or U5872 (N_5872,N_4810,N_2436);
and U5873 (N_5873,N_1503,N_3171);
or U5874 (N_5874,N_2606,N_4833);
or U5875 (N_5875,N_2663,N_3143);
and U5876 (N_5876,N_3404,N_3465);
nor U5877 (N_5877,N_1275,N_477);
xnor U5878 (N_5878,N_1775,N_814);
nor U5879 (N_5879,N_868,N_302);
or U5880 (N_5880,N_1108,N_2886);
and U5881 (N_5881,N_725,N_3638);
xnor U5882 (N_5882,N_381,N_1327);
or U5883 (N_5883,N_4594,N_4160);
xnor U5884 (N_5884,N_4464,N_3789);
and U5885 (N_5885,N_3786,N_446);
and U5886 (N_5886,N_1433,N_345);
and U5887 (N_5887,N_688,N_22);
or U5888 (N_5888,N_1274,N_2763);
and U5889 (N_5889,N_4112,N_70);
nor U5890 (N_5890,N_1223,N_3780);
nand U5891 (N_5891,N_4970,N_2137);
or U5892 (N_5892,N_4433,N_2649);
xnor U5893 (N_5893,N_1271,N_4034);
nand U5894 (N_5894,N_2510,N_579);
or U5895 (N_5895,N_3108,N_1008);
xor U5896 (N_5896,N_4904,N_810);
nor U5897 (N_5897,N_2191,N_1558);
nand U5898 (N_5898,N_3372,N_2123);
or U5899 (N_5899,N_1650,N_680);
and U5900 (N_5900,N_801,N_3311);
nand U5901 (N_5901,N_3891,N_2158);
nand U5902 (N_5902,N_690,N_4942);
xnor U5903 (N_5903,N_4042,N_225);
and U5904 (N_5904,N_4038,N_3412);
or U5905 (N_5905,N_2573,N_2522);
and U5906 (N_5906,N_1744,N_2911);
or U5907 (N_5907,N_432,N_3496);
and U5908 (N_5908,N_1761,N_4971);
and U5909 (N_5909,N_201,N_3849);
nor U5910 (N_5910,N_4505,N_767);
nor U5911 (N_5911,N_3993,N_4651);
and U5912 (N_5912,N_2896,N_3169);
xnor U5913 (N_5913,N_352,N_1036);
nor U5914 (N_5914,N_3695,N_4422);
or U5915 (N_5915,N_1124,N_2307);
nor U5916 (N_5916,N_67,N_394);
or U5917 (N_5917,N_480,N_571);
nand U5918 (N_5918,N_1693,N_2131);
xnor U5919 (N_5919,N_4906,N_1502);
xor U5920 (N_5920,N_1646,N_2141);
nor U5921 (N_5921,N_3792,N_1849);
xnor U5922 (N_5922,N_1094,N_1010);
nand U5923 (N_5923,N_2811,N_4036);
xor U5924 (N_5924,N_580,N_4645);
or U5925 (N_5925,N_4441,N_954);
and U5926 (N_5926,N_3502,N_1178);
nand U5927 (N_5927,N_3163,N_2943);
nand U5928 (N_5928,N_136,N_669);
and U5929 (N_5929,N_479,N_3255);
and U5930 (N_5930,N_4051,N_499);
xor U5931 (N_5931,N_3340,N_1576);
nand U5932 (N_5932,N_1113,N_3235);
or U5933 (N_5933,N_1760,N_3556);
xnor U5934 (N_5934,N_867,N_105);
nand U5935 (N_5935,N_716,N_4969);
nand U5936 (N_5936,N_886,N_921);
xor U5937 (N_5937,N_2498,N_1976);
and U5938 (N_5938,N_710,N_4817);
or U5939 (N_5939,N_3577,N_1328);
xor U5940 (N_5940,N_3129,N_331);
nand U5941 (N_5941,N_614,N_3400);
or U5942 (N_5942,N_4460,N_2768);
and U5943 (N_5943,N_575,N_3242);
xor U5944 (N_5944,N_3889,N_2827);
xnor U5945 (N_5945,N_3718,N_4167);
nor U5946 (N_5946,N_3366,N_3118);
or U5947 (N_5947,N_3380,N_2887);
and U5948 (N_5948,N_1917,N_4720);
nand U5949 (N_5949,N_2629,N_2005);
and U5950 (N_5950,N_3331,N_4127);
or U5951 (N_5951,N_4580,N_1957);
nand U5952 (N_5952,N_2298,N_3000);
xnor U5953 (N_5953,N_3924,N_1592);
and U5954 (N_5954,N_223,N_3260);
nor U5955 (N_5955,N_4516,N_1073);
xor U5956 (N_5956,N_3582,N_11);
nand U5957 (N_5957,N_2274,N_1814);
or U5958 (N_5958,N_2487,N_3887);
nand U5959 (N_5959,N_784,N_1218);
or U5960 (N_5960,N_188,N_2749);
nand U5961 (N_5961,N_3777,N_2659);
nand U5962 (N_5962,N_3914,N_1168);
and U5963 (N_5963,N_2217,N_1837);
nor U5964 (N_5964,N_1930,N_4106);
and U5965 (N_5965,N_2257,N_1745);
nor U5966 (N_5966,N_1347,N_1801);
or U5967 (N_5967,N_1164,N_3369);
or U5968 (N_5968,N_1512,N_1156);
or U5969 (N_5969,N_734,N_4386);
and U5970 (N_5970,N_1753,N_1145);
or U5971 (N_5971,N_260,N_1169);
nor U5972 (N_5972,N_4204,N_4019);
or U5973 (N_5973,N_370,N_2566);
xor U5974 (N_5974,N_1889,N_2347);
and U5975 (N_5975,N_3788,N_2215);
nor U5976 (N_5976,N_1858,N_3451);
and U5977 (N_5977,N_4966,N_1824);
xnor U5978 (N_5978,N_2120,N_4466);
and U5979 (N_5979,N_2902,N_221);
xor U5980 (N_5980,N_525,N_4846);
xnor U5981 (N_5981,N_2662,N_4955);
nand U5982 (N_5982,N_158,N_4363);
nand U5983 (N_5983,N_1676,N_3392);
or U5984 (N_5984,N_2409,N_1875);
nor U5985 (N_5985,N_4864,N_1721);
and U5986 (N_5986,N_1526,N_1499);
nand U5987 (N_5987,N_3707,N_4382);
nor U5988 (N_5988,N_4958,N_274);
xnor U5989 (N_5989,N_4546,N_884);
or U5990 (N_5990,N_822,N_2185);
and U5991 (N_5991,N_545,N_1542);
nand U5992 (N_5992,N_1376,N_4064);
xor U5993 (N_5993,N_2515,N_4487);
or U5994 (N_5994,N_4242,N_3322);
or U5995 (N_5995,N_3093,N_179);
nand U5996 (N_5996,N_743,N_1308);
xor U5997 (N_5997,N_2750,N_2899);
or U5998 (N_5998,N_3996,N_2746);
or U5999 (N_5999,N_679,N_1756);
and U6000 (N_6000,N_3885,N_3961);
or U6001 (N_6001,N_1120,N_1631);
nand U6002 (N_6002,N_1423,N_4159);
or U6003 (N_6003,N_4224,N_2817);
and U6004 (N_6004,N_1963,N_4945);
or U6005 (N_6005,N_2903,N_3121);
nand U6006 (N_6006,N_4109,N_927);
nand U6007 (N_6007,N_4929,N_1622);
and U6008 (N_6008,N_4457,N_616);
xor U6009 (N_6009,N_2517,N_2471);
nand U6010 (N_6010,N_4197,N_695);
nor U6011 (N_6011,N_2456,N_220);
or U6012 (N_6012,N_3395,N_1088);
xnor U6013 (N_6013,N_3966,N_2806);
nor U6014 (N_6014,N_2991,N_2572);
and U6015 (N_6015,N_1352,N_378);
or U6016 (N_6016,N_4696,N_766);
xnor U6017 (N_6017,N_3984,N_2759);
nor U6018 (N_6018,N_3038,N_955);
or U6019 (N_6019,N_732,N_3069);
and U6020 (N_6020,N_4427,N_2854);
nor U6021 (N_6021,N_3470,N_2144);
and U6022 (N_6022,N_4771,N_3029);
and U6023 (N_6023,N_3106,N_4366);
nor U6024 (N_6024,N_1510,N_4226);
and U6025 (N_6025,N_359,N_2165);
and U6026 (N_6026,N_469,N_1786);
or U6027 (N_6027,N_2304,N_1743);
xnor U6028 (N_6028,N_1024,N_1091);
xor U6029 (N_6029,N_333,N_1593);
nand U6030 (N_6030,N_1414,N_3902);
nand U6031 (N_6031,N_26,N_2597);
or U6032 (N_6032,N_1688,N_3060);
or U6033 (N_6033,N_3014,N_2079);
nand U6034 (N_6034,N_1669,N_3130);
nor U6035 (N_6035,N_3342,N_2056);
and U6036 (N_6036,N_3006,N_2065);
xor U6037 (N_6037,N_3228,N_3881);
nor U6038 (N_6038,N_1112,N_4689);
or U6039 (N_6039,N_1205,N_2147);
or U6040 (N_6040,N_1341,N_4891);
nand U6041 (N_6041,N_3081,N_4230);
xnor U6042 (N_6042,N_3717,N_3844);
xnor U6043 (N_6043,N_592,N_4059);
xnor U6044 (N_6044,N_4367,N_430);
and U6045 (N_6045,N_376,N_77);
xor U6046 (N_6046,N_2998,N_3051);
nand U6047 (N_6047,N_982,N_3459);
xnor U6048 (N_6048,N_3315,N_3054);
nor U6049 (N_6049,N_3208,N_3461);
and U6050 (N_6050,N_3977,N_4882);
xor U6051 (N_6051,N_2292,N_3022);
and U6052 (N_6052,N_2860,N_1796);
xor U6053 (N_6053,N_3850,N_4338);
nand U6054 (N_6054,N_1298,N_2000);
and U6055 (N_6055,N_4838,N_2824);
or U6056 (N_6056,N_1171,N_3288);
nand U6057 (N_6057,N_3403,N_1420);
and U6058 (N_6058,N_51,N_885);
nand U6059 (N_6059,N_4561,N_2680);
nand U6060 (N_6060,N_3651,N_4416);
xor U6061 (N_6061,N_1032,N_4336);
or U6062 (N_6062,N_2651,N_159);
and U6063 (N_6063,N_2859,N_4297);
xnor U6064 (N_6064,N_462,N_4152);
nor U6065 (N_6065,N_908,N_3371);
or U6066 (N_6066,N_2738,N_2917);
nor U6067 (N_6067,N_550,N_2117);
nor U6068 (N_6068,N_4155,N_4498);
and U6069 (N_6069,N_1466,N_2683);
nor U6070 (N_6070,N_2421,N_3264);
nand U6071 (N_6071,N_2778,N_1624);
nand U6072 (N_6072,N_2277,N_2278);
nand U6073 (N_6073,N_1966,N_2156);
or U6074 (N_6074,N_1667,N_4797);
and U6075 (N_6075,N_2797,N_384);
nand U6076 (N_6076,N_3363,N_2942);
nand U6077 (N_6077,N_1653,N_3252);
or U6078 (N_6078,N_3713,N_3261);
or U6079 (N_6079,N_949,N_2023);
nand U6080 (N_6080,N_4391,N_942);
nand U6081 (N_6081,N_4830,N_4558);
and U6082 (N_6082,N_1372,N_2689);
and U6083 (N_6083,N_1890,N_367);
nand U6084 (N_6084,N_2145,N_706);
nor U6085 (N_6085,N_1608,N_3017);
or U6086 (N_6086,N_1860,N_994);
nand U6087 (N_6087,N_3839,N_964);
or U6088 (N_6088,N_4405,N_3522);
and U6089 (N_6089,N_4602,N_3609);
nand U6090 (N_6090,N_1920,N_785);
or U6091 (N_6091,N_709,N_2378);
nand U6092 (N_6092,N_3309,N_3549);
xnor U6093 (N_6093,N_98,N_4658);
and U6094 (N_6094,N_392,N_1586);
xor U6095 (N_6095,N_2786,N_4780);
and U6096 (N_6096,N_2505,N_658);
xnor U6097 (N_6097,N_4047,N_3230);
and U6098 (N_6098,N_2400,N_2328);
nor U6099 (N_6099,N_2742,N_1842);
and U6100 (N_6100,N_790,N_1863);
or U6101 (N_6101,N_4032,N_4451);
xnor U6102 (N_6102,N_4375,N_2499);
and U6103 (N_6103,N_4610,N_2530);
or U6104 (N_6104,N_4028,N_478);
or U6105 (N_6105,N_4003,N_4822);
or U6106 (N_6106,N_635,N_2170);
nor U6107 (N_6107,N_2048,N_3937);
and U6108 (N_6108,N_190,N_261);
nand U6109 (N_6109,N_303,N_540);
or U6110 (N_6110,N_3096,N_823);
nand U6111 (N_6111,N_1334,N_4072);
xor U6112 (N_6112,N_513,N_3910);
nor U6113 (N_6113,N_389,N_1968);
or U6114 (N_6114,N_2672,N_2172);
xor U6115 (N_6115,N_1972,N_3550);
or U6116 (N_6116,N_3196,N_1563);
nor U6117 (N_6117,N_3040,N_106);
and U6118 (N_6118,N_391,N_4717);
nand U6119 (N_6119,N_3879,N_3901);
or U6120 (N_6120,N_411,N_156);
and U6121 (N_6121,N_163,N_1696);
xnor U6122 (N_6122,N_149,N_4851);
nand U6123 (N_6123,N_3146,N_4294);
nand U6124 (N_6124,N_4404,N_4951);
and U6125 (N_6125,N_4309,N_1942);
nand U6126 (N_6126,N_1019,N_335);
nor U6127 (N_6127,N_178,N_1766);
nand U6128 (N_6128,N_522,N_1642);
nor U6129 (N_6129,N_1677,N_2526);
nor U6130 (N_6130,N_4544,N_4420);
and U6131 (N_6131,N_1536,N_1973);
xnor U6132 (N_6132,N_1649,N_3484);
or U6133 (N_6133,N_3815,N_258);
nor U6134 (N_6134,N_4858,N_898);
xnor U6135 (N_6135,N_1009,N_2154);
nor U6136 (N_6136,N_4530,N_1488);
nand U6137 (N_6137,N_408,N_3727);
nor U6138 (N_6138,N_1389,N_3280);
nor U6139 (N_6139,N_4165,N_1722);
and U6140 (N_6140,N_2495,N_3475);
or U6141 (N_6141,N_1913,N_3125);
xnor U6142 (N_6142,N_2971,N_980);
and U6143 (N_6143,N_3862,N_2664);
or U6144 (N_6144,N_2113,N_700);
nor U6145 (N_6145,N_4670,N_1202);
xor U6146 (N_6146,N_506,N_2661);
nor U6147 (N_6147,N_3102,N_2198);
or U6148 (N_6148,N_243,N_3979);
nor U6149 (N_6149,N_3127,N_4343);
and U6150 (N_6150,N_2166,N_991);
nor U6151 (N_6151,N_1529,N_4869);
and U6152 (N_6152,N_4215,N_702);
and U6153 (N_6153,N_1886,N_2013);
or U6154 (N_6154,N_2965,N_4194);
or U6155 (N_6155,N_817,N_3272);
nand U6156 (N_6156,N_1554,N_3430);
nand U6157 (N_6157,N_56,N_4483);
nor U6158 (N_6158,N_1193,N_1444);
xor U6159 (N_6159,N_3564,N_4510);
nor U6160 (N_6160,N_735,N_2486);
and U6161 (N_6161,N_1777,N_1921);
and U6162 (N_6162,N_4808,N_627);
or U6163 (N_6163,N_1176,N_2546);
nor U6164 (N_6164,N_1418,N_3580);
and U6165 (N_6165,N_2519,N_2078);
or U6166 (N_6166,N_651,N_4908);
xor U6167 (N_6167,N_280,N_1317);
nand U6168 (N_6168,N_4490,N_3909);
nor U6169 (N_6169,N_412,N_351);
nand U6170 (N_6170,N_1643,N_931);
xnor U6171 (N_6171,N_3821,N_4812);
and U6172 (N_6172,N_2666,N_946);
nand U6173 (N_6173,N_765,N_3968);
nand U6174 (N_6174,N_2381,N_1134);
xnor U6175 (N_6175,N_809,N_1687);
or U6176 (N_6176,N_2350,N_3826);
nor U6177 (N_6177,N_407,N_4480);
xor U6178 (N_6178,N_664,N_3485);
or U6179 (N_6179,N_3180,N_1544);
nor U6180 (N_6180,N_1782,N_396);
or U6181 (N_6181,N_4698,N_4092);
and U6182 (N_6182,N_1736,N_2443);
and U6183 (N_6183,N_532,N_1938);
xor U6184 (N_6184,N_2538,N_62);
nor U6185 (N_6185,N_2536,N_2112);
nor U6186 (N_6186,N_1326,N_8);
xnor U6187 (N_6187,N_2326,N_989);
nor U6188 (N_6188,N_1752,N_4711);
and U6189 (N_6189,N_3934,N_739);
or U6190 (N_6190,N_4740,N_182);
nand U6191 (N_6191,N_2211,N_267);
or U6192 (N_6192,N_3162,N_4129);
xor U6193 (N_6193,N_4943,N_910);
xor U6194 (N_6194,N_4100,N_347);
nor U6195 (N_6195,N_1210,N_4435);
nand U6196 (N_6196,N_619,N_2196);
nor U6197 (N_6197,N_2924,N_567);
xor U6198 (N_6198,N_4121,N_3769);
nor U6199 (N_6199,N_2007,N_1030);
or U6200 (N_6200,N_3436,N_3606);
and U6201 (N_6201,N_1443,N_4029);
and U6202 (N_6202,N_3164,N_320);
and U6203 (N_6203,N_2851,N_3867);
nor U6204 (N_6204,N_587,N_880);
nor U6205 (N_6205,N_936,N_841);
and U6206 (N_6206,N_2667,N_681);
or U6207 (N_6207,N_244,N_2465);
xor U6208 (N_6208,N_3518,N_2447);
or U6209 (N_6209,N_711,N_1700);
and U6210 (N_6210,N_135,N_3665);
and U6211 (N_6211,N_2845,N_1441);
or U6212 (N_6212,N_1381,N_2591);
xnor U6213 (N_6213,N_2160,N_2767);
nor U6214 (N_6214,N_2757,N_2238);
nor U6215 (N_6215,N_750,N_2537);
or U6216 (N_6216,N_1731,N_3647);
or U6217 (N_6217,N_6,N_365);
or U6218 (N_6218,N_4325,N_2132);
nor U6219 (N_6219,N_3507,N_756);
nand U6220 (N_6220,N_4738,N_1493);
or U6221 (N_6221,N_1417,N_2368);
nand U6222 (N_6222,N_4191,N_3087);
and U6223 (N_6223,N_1868,N_3759);
or U6224 (N_6224,N_4820,N_1063);
and U6225 (N_6225,N_3375,N_43);
xnor U6226 (N_6226,N_65,N_617);
nand U6227 (N_6227,N_3712,N_2072);
xnor U6228 (N_6228,N_4517,N_372);
and U6229 (N_6229,N_3276,N_3304);
or U6230 (N_6230,N_1387,N_4636);
or U6231 (N_6231,N_3835,N_3486);
or U6232 (N_6232,N_4381,N_2964);
nor U6233 (N_6233,N_876,N_1651);
nor U6234 (N_6234,N_3579,N_3525);
nor U6235 (N_6235,N_2950,N_2410);
xnor U6236 (N_6236,N_4010,N_4068);
and U6237 (N_6237,N_4210,N_2146);
or U6238 (N_6238,N_856,N_836);
nor U6239 (N_6239,N_990,N_889);
nand U6240 (N_6240,N_758,N_1975);
nor U6241 (N_6241,N_840,N_4666);
xor U6242 (N_6242,N_2446,N_1390);
xnor U6243 (N_6243,N_3306,N_3364);
nand U6244 (N_6244,N_4091,N_2270);
or U6245 (N_6245,N_4735,N_2387);
and U6246 (N_6246,N_4742,N_3499);
xnor U6247 (N_6247,N_4046,N_4407);
or U6248 (N_6248,N_2925,N_4419);
nor U6249 (N_6249,N_3222,N_1588);
xor U6250 (N_6250,N_373,N_2149);
and U6251 (N_6251,N_2164,N_316);
nor U6252 (N_6252,N_2711,N_2810);
nor U6253 (N_6253,N_211,N_4608);
nand U6254 (N_6254,N_3629,N_1909);
nor U6255 (N_6255,N_239,N_3055);
nand U6256 (N_6256,N_1923,N_4511);
nor U6257 (N_6257,N_2756,N_2171);
or U6258 (N_6258,N_1579,N_2293);
and U6259 (N_6259,N_2723,N_1960);
nor U6260 (N_6260,N_2721,N_1427);
and U6261 (N_6261,N_938,N_4406);
or U6262 (N_6262,N_4119,N_4189);
and U6263 (N_6263,N_3927,N_2956);
or U6264 (N_6264,N_4832,N_3565);
nor U6265 (N_6265,N_3865,N_1011);
nand U6266 (N_6266,N_4500,N_3687);
and U6267 (N_6267,N_4829,N_4883);
and U6268 (N_6268,N_4411,N_3923);
xnor U6269 (N_6269,N_35,N_95);
nor U6270 (N_6270,N_4017,N_4192);
nor U6271 (N_6271,N_3147,N_4895);
nor U6272 (N_6272,N_4983,N_4568);
and U6273 (N_6273,N_4750,N_3858);
xnor U6274 (N_6274,N_3086,N_1548);
or U6275 (N_6275,N_2372,N_2507);
and U6276 (N_6276,N_1727,N_4506);
xor U6277 (N_6277,N_3384,N_1465);
nor U6278 (N_6278,N_1431,N_3962);
or U6279 (N_6279,N_2987,N_1901);
nor U6280 (N_6280,N_167,N_3871);
nand U6281 (N_6281,N_1682,N_4583);
and U6282 (N_6282,N_3938,N_1954);
xnor U6283 (N_6283,N_3811,N_1469);
xor U6284 (N_6284,N_2980,N_1912);
xor U6285 (N_6285,N_3559,N_93);
and U6286 (N_6286,N_4305,N_2481);
nor U6287 (N_6287,N_3595,N_2376);
or U6288 (N_6288,N_3552,N_2807);
xnor U6289 (N_6289,N_2630,N_309);
or U6290 (N_6290,N_1454,N_3863);
and U6291 (N_6291,N_4270,N_632);
xor U6292 (N_6292,N_4327,N_1945);
nand U6293 (N_6293,N_2540,N_2414);
xnor U6294 (N_6294,N_440,N_2485);
or U6295 (N_6295,N_3666,N_300);
and U6296 (N_6296,N_3033,N_3244);
or U6297 (N_6297,N_2731,N_1528);
nand U6298 (N_6298,N_2383,N_1630);
xnor U6299 (N_6299,N_3201,N_1870);
nand U6300 (N_6300,N_1485,N_595);
nand U6301 (N_6301,N_763,N_3649);
xnor U6302 (N_6302,N_4521,N_4907);
or U6303 (N_6303,N_4730,N_3204);
xor U6304 (N_6304,N_1415,N_4331);
nor U6305 (N_6305,N_1964,N_2367);
xnor U6306 (N_6306,N_74,N_2193);
or U6307 (N_6307,N_3768,N_418);
or U6308 (N_6308,N_3653,N_4188);
or U6309 (N_6309,N_965,N_3480);
nand U6310 (N_6310,N_2670,N_3964);
nand U6311 (N_6311,N_2647,N_718);
nor U6312 (N_6312,N_2881,N_4073);
nand U6313 (N_6313,N_792,N_2262);
and U6314 (N_6314,N_1468,N_4549);
nand U6315 (N_6315,N_913,N_1950);
xnor U6316 (N_6316,N_465,N_584);
nor U6317 (N_6317,N_458,N_4239);
xnor U6318 (N_6318,N_1603,N_198);
xor U6319 (N_6319,N_3869,N_4871);
nand U6320 (N_6320,N_2783,N_2483);
nand U6321 (N_6321,N_2644,N_1840);
xor U6322 (N_6322,N_1344,N_3098);
or U6323 (N_6323,N_1071,N_4856);
xor U6324 (N_6324,N_1856,N_283);
nand U6325 (N_6325,N_2610,N_4937);
nor U6326 (N_6326,N_2787,N_3624);
xor U6327 (N_6327,N_3092,N_4831);
and U6328 (N_6328,N_4805,N_4196);
xor U6329 (N_6329,N_2952,N_1473);
and U6330 (N_6330,N_4719,N_2083);
nand U6331 (N_6331,N_3336,N_3325);
nand U6332 (N_6332,N_169,N_2085);
nor U6333 (N_6333,N_2587,N_4387);
or U6334 (N_6334,N_3758,N_4916);
xor U6335 (N_6335,N_2668,N_3851);
xnor U6336 (N_6336,N_3546,N_4634);
nor U6337 (N_6337,N_3095,N_4677);
nand U6338 (N_6338,N_830,N_2325);
nor U6339 (N_6339,N_852,N_4180);
nor U6340 (N_6340,N_1140,N_4492);
nor U6341 (N_6341,N_4956,N_21);
nor U6342 (N_6342,N_4865,N_4281);
nand U6343 (N_6343,N_4443,N_3706);
nand U6344 (N_6344,N_3610,N_3083);
and U6345 (N_6345,N_4872,N_960);
and U6346 (N_6346,N_2494,N_3842);
xnor U6347 (N_6347,N_1360,N_4662);
and U6348 (N_6348,N_834,N_5);
nor U6349 (N_6349,N_108,N_1060);
and U6350 (N_6350,N_4006,N_3683);
and U6351 (N_6351,N_4839,N_231);
xnor U6352 (N_6352,N_452,N_4625);
xnor U6353 (N_6353,N_4947,N_3636);
or U6354 (N_6354,N_2488,N_3948);
and U6355 (N_6355,N_2284,N_81);
or U6356 (N_6356,N_1337,N_3002);
and U6357 (N_6357,N_3321,N_2004);
or U6358 (N_6358,N_1922,N_1895);
nor U6359 (N_6359,N_4252,N_2639);
xnor U6360 (N_6360,N_3895,N_951);
nand U6361 (N_6361,N_2976,N_3192);
and U6362 (N_6362,N_981,N_293);
or U6363 (N_6363,N_3181,N_4965);
xor U6364 (N_6364,N_791,N_2418);
or U6365 (N_6365,N_3269,N_2557);
and U6366 (N_6366,N_233,N_380);
and U6367 (N_6367,N_914,N_628);
and U6368 (N_6368,N_3853,N_1079);
nor U6369 (N_6369,N_777,N_4699);
nor U6370 (N_6370,N_952,N_1395);
nor U6371 (N_6371,N_2559,N_4815);
and U6372 (N_6372,N_1719,N_4328);
and U6373 (N_6373,N_1994,N_4591);
and U6374 (N_6374,N_4372,N_2332);
nand U6375 (N_6375,N_3044,N_2477);
and U6376 (N_6376,N_3157,N_2243);
nand U6377 (N_6377,N_620,N_4261);
nand U6378 (N_6378,N_859,N_824);
xor U6379 (N_6379,N_467,N_4806);
nand U6380 (N_6380,N_2791,N_2823);
or U6381 (N_6381,N_101,N_2398);
nor U6382 (N_6382,N_3203,N_4581);
nand U6383 (N_6383,N_2063,N_2339);
nand U6384 (N_6384,N_647,N_4724);
xnor U6385 (N_6385,N_1438,N_375);
nor U6386 (N_6386,N_2295,N_1221);
nor U6387 (N_6387,N_1937,N_1645);
xnor U6388 (N_6388,N_1142,N_3042);
xor U6389 (N_6389,N_1031,N_2678);
and U6390 (N_6390,N_697,N_1173);
and U6391 (N_6391,N_3434,N_1131);
or U6392 (N_6392,N_3,N_109);
nor U6393 (N_6393,N_4315,N_4110);
or U6394 (N_6394,N_4917,N_754);
nand U6395 (N_6395,N_2393,N_1074);
or U6396 (N_6396,N_4600,N_145);
nand U6397 (N_6397,N_3620,N_1251);
or U6398 (N_6398,N_142,N_4209);
xnor U6399 (N_6399,N_2028,N_3661);
or U6400 (N_6400,N_4491,N_3753);
nor U6401 (N_6401,N_3313,N_953);
or U6402 (N_6402,N_1470,N_3221);
nor U6403 (N_6403,N_4751,N_4876);
xnor U6404 (N_6404,N_1311,N_4619);
or U6405 (N_6405,N_1363,N_2233);
and U6406 (N_6406,N_1873,N_626);
and U6407 (N_6407,N_2712,N_854);
or U6408 (N_6408,N_2782,N_2967);
xor U6409 (N_6409,N_4444,N_2290);
and U6410 (N_6410,N_2139,N_2898);
or U6411 (N_6411,N_4118,N_4494);
and U6412 (N_6412,N_1211,N_1846);
xor U6413 (N_6413,N_1927,N_3542);
nand U6414 (N_6414,N_1236,N_829);
nand U6415 (N_6415,N_2919,N_1336);
xnor U6416 (N_6416,N_1125,N_1136);
nor U6417 (N_6417,N_723,N_61);
nand U6418 (N_6418,N_839,N_46);
and U6419 (N_6419,N_3551,N_3561);
or U6420 (N_6420,N_947,N_217);
xor U6421 (N_6421,N_3019,N_1182);
and U6422 (N_6422,N_1634,N_3854);
nor U6423 (N_6423,N_1867,N_4577);
nand U6424 (N_6424,N_4,N_3211);
or U6425 (N_6425,N_2268,N_3279);
nand U6426 (N_6426,N_2066,N_3529);
or U6427 (N_6427,N_2745,N_4470);
nand U6428 (N_6428,N_1871,N_349);
nand U6429 (N_6429,N_2753,N_2972);
nand U6430 (N_6430,N_4368,N_3212);
nor U6431 (N_6431,N_3646,N_4183);
xnor U6432 (N_6432,N_3816,N_2454);
nor U6433 (N_6433,N_3132,N_2936);
xnor U6434 (N_6434,N_929,N_4308);
xnor U6435 (N_6435,N_4026,N_3410);
xor U6436 (N_6436,N_3027,N_4105);
and U6437 (N_6437,N_3239,N_14);
and U6438 (N_6438,N_1161,N_285);
xnor U6439 (N_6439,N_3987,N_4002);
and U6440 (N_6440,N_2554,N_2348);
nor U6441 (N_6441,N_4448,N_4930);
nor U6442 (N_6442,N_2665,N_4207);
and U6443 (N_6443,N_3460,N_1135);
xor U6444 (N_6444,N_3076,N_4747);
nand U6445 (N_6445,N_3569,N_572);
or U6446 (N_6446,N_4187,N_4302);
or U6447 (N_6447,N_2922,N_3291);
or U6448 (N_6448,N_1301,N_463);
and U6449 (N_6449,N_3899,N_3947);
or U6450 (N_6450,N_1690,N_1368);
nand U6451 (N_6451,N_1762,N_2945);
nand U6452 (N_6452,N_645,N_193);
and U6453 (N_6453,N_4084,N_3074);
or U6454 (N_6454,N_2549,N_166);
xor U6455 (N_6455,N_703,N_1046);
and U6456 (N_6456,N_1100,N_3217);
and U6457 (N_6457,N_3761,N_3946);
and U6458 (N_6458,N_1281,N_984);
xnor U6459 (N_6459,N_96,N_2458);
xnor U6460 (N_6460,N_2417,N_237);
nor U6461 (N_6461,N_2752,N_4078);
nand U6462 (N_6462,N_1615,N_641);
or U6463 (N_6463,N_4130,N_2985);
or U6464 (N_6464,N_1644,N_68);
xnor U6465 (N_6465,N_3673,N_2358);
nor U6466 (N_6466,N_1122,N_245);
nand U6467 (N_6467,N_2938,N_1090);
nand U6468 (N_6468,N_2142,N_1967);
and U6469 (N_6469,N_2842,N_3972);
nor U6470 (N_6470,N_1611,N_1839);
xnor U6471 (N_6471,N_3955,N_1167);
or U6472 (N_6472,N_3940,N_2433);
nand U6473 (N_6473,N_264,N_1102);
and U6474 (N_6474,N_4650,N_270);
nand U6475 (N_6475,N_3830,N_1742);
nand U6476 (N_6476,N_3950,N_665);
or U6477 (N_6477,N_3750,N_1599);
and U6478 (N_6478,N_1768,N_3379);
nor U6479 (N_6479,N_2853,N_3383);
and U6480 (N_6480,N_3520,N_2255);
nor U6481 (N_6481,N_2135,N_1247);
xnor U6482 (N_6482,N_447,N_652);
and U6483 (N_6483,N_1369,N_1946);
nor U6484 (N_6484,N_2687,N_1306);
xor U6485 (N_6485,N_4200,N_4980);
xor U6486 (N_6486,N_180,N_2607);
xor U6487 (N_6487,N_137,N_2790);
and U6488 (N_6488,N_1717,N_1061);
nand U6489 (N_6489,N_4258,N_4153);
xor U6490 (N_6490,N_1732,N_3506);
nand U6491 (N_6491,N_2979,N_3360);
nand U6492 (N_6492,N_2121,N_2611);
nand U6493 (N_6493,N_573,N_2794);
or U6494 (N_6494,N_2441,N_208);
or U6495 (N_6495,N_1711,N_1832);
and U6496 (N_6496,N_1092,N_2391);
or U6497 (N_6497,N_36,N_4534);
nor U6498 (N_6498,N_4923,N_4318);
and U6499 (N_6499,N_755,N_286);
or U6500 (N_6500,N_590,N_92);
nand U6501 (N_6501,N_1803,N_1475);
xnor U6502 (N_6502,N_3282,N_4802);
nand U6503 (N_6503,N_2704,N_2957);
xnor U6504 (N_6504,N_2272,N_3206);
and U6505 (N_6505,N_3767,N_3473);
and U6506 (N_6506,N_3748,N_4067);
nor U6507 (N_6507,N_88,N_2088);
nor U6508 (N_6508,N_3601,N_4639);
or U6509 (N_6509,N_1795,N_2206);
or U6510 (N_6510,N_727,N_3362);
xnor U6511 (N_6511,N_2018,N_1810);
xnor U6512 (N_6512,N_4465,N_3300);
or U6513 (N_6513,N_2489,N_3085);
and U6514 (N_6514,N_1471,N_1021);
and U6515 (N_6515,N_196,N_3544);
and U6516 (N_6516,N_2575,N_299);
nor U6517 (N_6517,N_3878,N_891);
xor U6518 (N_6518,N_4149,N_427);
nand U6519 (N_6519,N_943,N_414);
or U6520 (N_6520,N_2577,N_2022);
nand U6521 (N_6521,N_3975,N_2815);
nor U6522 (N_6522,N_2933,N_2493);
nand U6523 (N_6523,N_3016,N_4782);
or U6524 (N_6524,N_4672,N_4935);
and U6525 (N_6525,N_4045,N_1213);
and U6526 (N_6526,N_4814,N_4537);
nor U6527 (N_6527,N_1144,N_4295);
xor U6528 (N_6528,N_2429,N_1617);
nor U6529 (N_6529,N_2981,N_2275);
and U6530 (N_6530,N_2340,N_1386);
xor U6531 (N_6531,N_1809,N_4142);
or U6532 (N_6532,N_3120,N_3600);
and U6533 (N_6533,N_3101,N_1931);
nand U6534 (N_6534,N_4800,N_3186);
or U6535 (N_6535,N_2904,N_4749);
xor U6536 (N_6536,N_4175,N_1017);
nand U6537 (N_6537,N_3742,N_4307);
or U6538 (N_6538,N_1379,N_2386);
nor U6539 (N_6539,N_1259,N_509);
and U6540 (N_6540,N_4708,N_1265);
xnor U6541 (N_6541,N_906,N_1446);
nand U6542 (N_6542,N_4901,N_1986);
and U6543 (N_6543,N_636,N_1625);
nand U6544 (N_6544,N_3809,N_3285);
or U6545 (N_6545,N_129,N_4300);
nor U6546 (N_6546,N_2708,N_2174);
and U6547 (N_6547,N_4450,N_1450);
xnor U6548 (N_6548,N_4588,N_3394);
xor U6549 (N_6549,N_4866,N_2855);
or U6550 (N_6550,N_3310,N_3764);
nand U6551 (N_6551,N_589,N_3117);
nand U6552 (N_6552,N_3257,N_1354);
nand U6553 (N_6553,N_117,N_2464);
and U6554 (N_6554,N_4266,N_2380);
xnor U6555 (N_6555,N_557,N_3511);
xor U6556 (N_6556,N_3240,N_3857);
nor U6557 (N_6557,N_1709,N_610);
or U6558 (N_6558,N_4632,N_3063);
nand U6559 (N_6559,N_774,N_4571);
or U6560 (N_6560,N_655,N_689);
and U6561 (N_6561,N_4657,N_3791);
xnor U6562 (N_6562,N_4533,N_1452);
nor U6563 (N_6563,N_3425,N_2087);
and U6564 (N_6564,N_4081,N_4741);
nand U6565 (N_6565,N_3072,N_4515);
xnor U6566 (N_6566,N_4644,N_1740);
nand U6567 (N_6567,N_2107,N_387);
or U6568 (N_6568,N_3637,N_1241);
and U6569 (N_6569,N_939,N_2877);
and U6570 (N_6570,N_912,N_382);
and U6571 (N_6571,N_3900,N_4788);
and U6572 (N_6572,N_3852,N_3267);
nor U6573 (N_6573,N_2564,N_2309);
or U6574 (N_6574,N_2527,N_3720);
or U6575 (N_6575,N_1570,N_807);
nor U6576 (N_6576,N_1183,N_3209);
or U6577 (N_6577,N_717,N_4249);
or U6578 (N_6578,N_139,N_3859);
nand U6579 (N_6579,N_4791,N_1533);
and U6580 (N_6580,N_4256,N_1703);
nand U6581 (N_6581,N_1128,N_2450);
or U6582 (N_6582,N_3875,N_4597);
and U6583 (N_6583,N_2839,N_3154);
nor U6584 (N_6584,N_3270,N_3632);
xor U6585 (N_6585,N_3848,N_1078);
and U6586 (N_6586,N_618,N_3659);
nand U6587 (N_6587,N_1983,N_3299);
or U6588 (N_6588,N_4607,N_1392);
xor U6589 (N_6589,N_2415,N_3043);
xnor U6590 (N_6590,N_759,N_327);
xor U6591 (N_6591,N_1093,N_1148);
or U6592 (N_6592,N_3709,N_3338);
xnor U6593 (N_6593,N_103,N_762);
and U6594 (N_6594,N_1067,N_4478);
nor U6595 (N_6595,N_3794,N_742);
and U6596 (N_6596,N_644,N_3036);
and U6597 (N_6597,N_2975,N_1530);
and U6598 (N_6598,N_2894,N_3817);
or U6599 (N_6599,N_4385,N_4140);
and U6600 (N_6600,N_3335,N_4240);
xnor U6601 (N_6601,N_966,N_2634);
or U6602 (N_6602,N_2060,N_3166);
nor U6603 (N_6603,N_4873,N_2800);
xor U6604 (N_6604,N_1818,N_3066);
xor U6605 (N_6605,N_3500,N_4079);
and U6606 (N_6606,N_2260,N_4048);
and U6607 (N_6607,N_1106,N_2681);
and U6608 (N_6608,N_4712,N_4729);
nor U6609 (N_6609,N_672,N_113);
xor U6610 (N_6610,N_2103,N_2849);
nor U6611 (N_6611,N_161,N_4195);
nor U6612 (N_6612,N_4132,N_998);
nand U6613 (N_6613,N_656,N_1561);
nor U6614 (N_6614,N_2385,N_630);
or U6615 (N_6615,N_3795,N_959);
and U6616 (N_6616,N_848,N_833);
or U6617 (N_6617,N_3698,N_3739);
or U6618 (N_6618,N_1763,N_1147);
nand U6619 (N_6619,N_2714,N_4823);
or U6620 (N_6620,N_574,N_1830);
and U6621 (N_6621,N_4514,N_3997);
or U6622 (N_6622,N_4399,N_1208);
or U6623 (N_6623,N_3390,N_3476);
xnor U6624 (N_6624,N_3296,N_2563);
xnor U6625 (N_6625,N_4555,N_4566);
or U6626 (N_6626,N_4211,N_2622);
and U6627 (N_6627,N_741,N_2396);
or U6628 (N_6628,N_1828,N_364);
xnor U6629 (N_6629,N_2106,N_3011);
or U6630 (N_6630,N_2650,N_1852);
nand U6631 (N_6631,N_177,N_1044);
and U6632 (N_6632,N_3614,N_3137);
and U6633 (N_6633,N_3358,N_3974);
nor U6634 (N_6634,N_3139,N_2518);
and U6635 (N_6635,N_1305,N_3693);
nor U6636 (N_6636,N_2716,N_3053);
and U6637 (N_6637,N_2906,N_4346);
and U6638 (N_6638,N_1855,N_4959);
nor U6639 (N_6639,N_3464,N_1941);
or U6640 (N_6640,N_4702,N_3519);
and U6641 (N_6641,N_1424,N_4311);
or U6642 (N_6642,N_4117,N_850);
and U6643 (N_6643,N_3233,N_3318);
nor U6644 (N_6644,N_1547,N_1678);
nand U6645 (N_6645,N_2551,N_2428);
xor U6646 (N_6646,N_2694,N_385);
nor U6647 (N_6647,N_4377,N_3477);
nor U6648 (N_6648,N_4263,N_4542);
nand U6649 (N_6649,N_4349,N_1377);
nor U6650 (N_6650,N_1406,N_4220);
nor U6651 (N_6651,N_3333,N_1799);
or U6652 (N_6652,N_3176,N_3697);
or U6653 (N_6653,N_1496,N_2254);
nand U6654 (N_6654,N_4323,N_917);
or U6655 (N_6655,N_4803,N_2660);
nor U6656 (N_6656,N_90,N_401);
nor U6657 (N_6657,N_4992,N_2204);
nor U6658 (N_6658,N_3492,N_3904);
nand U6659 (N_6659,N_3585,N_3640);
xor U6660 (N_6660,N_2888,N_4489);
nand U6661 (N_6661,N_1755,N_265);
xnor U6662 (N_6662,N_4313,N_2212);
nand U6663 (N_6663,N_1070,N_1956);
or U6664 (N_6664,N_2321,N_1715);
xor U6665 (N_6665,N_2317,N_1109);
xnor U6666 (N_6666,N_3153,N_3030);
and U6667 (N_6667,N_3912,N_1612);
nor U6668 (N_6668,N_433,N_2280);
or U6669 (N_6669,N_3501,N_2703);
or U6670 (N_6670,N_4982,N_437);
xor U6671 (N_6671,N_2037,N_2043);
xor U6672 (N_6672,N_2201,N_701);
or U6673 (N_6673,N_3534,N_1924);
xor U6674 (N_6674,N_586,N_3437);
or U6675 (N_6675,N_3705,N_2675);
or U6676 (N_6676,N_1300,N_2876);
nor U6677 (N_6677,N_3664,N_2990);
and U6678 (N_6678,N_4543,N_2977);
and U6679 (N_6679,N_4737,N_1364);
nand U6680 (N_6680,N_2457,N_2167);
or U6681 (N_6681,N_577,N_425);
and U6682 (N_6682,N_4326,N_2252);
nand U6683 (N_6683,N_3168,N_1997);
nand U6684 (N_6684,N_4635,N_3207);
nor U6685 (N_6685,N_1155,N_520);
nand U6686 (N_6686,N_599,N_4082);
xnor U6687 (N_6687,N_3513,N_1246);
or U6688 (N_6688,N_1511,N_3949);
and U6689 (N_6689,N_3173,N_2406);
xnor U6690 (N_6690,N_1707,N_1312);
xor U6691 (N_6691,N_2646,N_235);
xnor U6692 (N_6692,N_1325,N_4428);
nand U6693 (N_6693,N_49,N_3781);
nand U6694 (N_6694,N_2285,N_2983);
xor U6695 (N_6695,N_3722,N_693);
and U6696 (N_6696,N_4061,N_4039);
xor U6697 (N_6697,N_4531,N_2012);
xor U6698 (N_6698,N_812,N_2006);
and U6699 (N_6699,N_4936,N_1844);
xor U6700 (N_6700,N_2609,N_2363);
nor U6701 (N_6701,N_3589,N_1685);
xnor U6702 (N_6702,N_928,N_1996);
and U6703 (N_6703,N_2521,N_3348);
xor U6704 (N_6704,N_1607,N_3874);
nand U6705 (N_6705,N_4626,N_678);
or U6706 (N_6706,N_902,N_1378);
nand U6707 (N_6707,N_1948,N_2331);
nor U6708 (N_6708,N_4116,N_933);
nor U6709 (N_6709,N_1933,N_1435);
nand U6710 (N_6710,N_4601,N_1854);
and U6711 (N_6711,N_2124,N_2143);
and U6712 (N_6712,N_548,N_3075);
or U6713 (N_6713,N_4977,N_518);
or U6714 (N_6714,N_2841,N_1746);
nand U6715 (N_6715,N_1286,N_4728);
nor U6716 (N_6716,N_1447,N_3732);
nand U6717 (N_6717,N_4301,N_4867);
nor U6718 (N_6718,N_1729,N_3406);
xor U6719 (N_6719,N_1080,N_3943);
nand U6720 (N_6720,N_1103,N_1000);
nor U6721 (N_6721,N_3798,N_3973);
nor U6722 (N_6722,N_2761,N_4501);
nor U6723 (N_6723,N_2962,N_4963);
nand U6724 (N_6724,N_4254,N_4182);
xor U6725 (N_6725,N_4146,N_4063);
nor U6726 (N_6726,N_2825,N_837);
xnor U6727 (N_6727,N_862,N_1939);
nor U6728 (N_6728,N_3421,N_4695);
nand U6729 (N_6729,N_3771,N_944);
nor U6730 (N_6730,N_3012,N_1783);
nand U6731 (N_6731,N_2926,N_526);
and U6732 (N_6732,N_1027,N_121);
xor U6733 (N_6733,N_4875,N_3231);
nor U6734 (N_6734,N_3028,N_2715);
nor U6735 (N_6735,N_125,N_4536);
nand U6736 (N_6736,N_2912,N_1356);
or U6737 (N_6737,N_3951,N_4122);
and U6738 (N_6738,N_1905,N_1319);
or U6739 (N_6739,N_2804,N_238);
nor U6740 (N_6740,N_3405,N_3216);
xnor U6741 (N_6741,N_2127,N_3286);
nand U6742 (N_6742,N_3393,N_2192);
nand U6743 (N_6743,N_2401,N_2834);
or U6744 (N_6744,N_1998,N_288);
nor U6745 (N_6745,N_3524,N_4358);
or U6746 (N_6746,N_4612,N_585);
nand U6747 (N_6747,N_1936,N_4941);
xor U6748 (N_6748,N_2862,N_3277);
nand U6749 (N_6749,N_560,N_2276);
nand U6750 (N_6750,N_696,N_1569);
or U6751 (N_6751,N_1778,N_317);
nand U6752 (N_6752,N_4898,N_1712);
nor U6753 (N_6753,N_87,N_3682);
nor U6754 (N_6754,N_692,N_4726);
or U6755 (N_6755,N_3428,N_3991);
or U6756 (N_6756,N_999,N_2645);
nor U6757 (N_6757,N_4843,N_3457);
nand U6758 (N_6758,N_3414,N_643);
and U6759 (N_6759,N_3308,N_892);
xnor U6760 (N_6760,N_4654,N_1065);
and U6761 (N_6761,N_2771,N_2431);
nand U6762 (N_6762,N_1794,N_3512);
or U6763 (N_6763,N_2918,N_1303);
or U6764 (N_6764,N_1157,N_2857);
nor U6765 (N_6765,N_457,N_1235);
or U6766 (N_6766,N_3067,N_2199);
nor U6767 (N_6767,N_1784,N_851);
xor U6768 (N_6768,N_3397,N_1266);
nor U6769 (N_6769,N_4598,N_222);
nor U6770 (N_6770,N_648,N_4499);
or U6771 (N_6771,N_1540,N_3297);
nor U6772 (N_6772,N_314,N_1098);
nand U6773 (N_6773,N_2781,N_3339);
nand U6774 (N_6774,N_4251,N_2434);
or U6775 (N_6775,N_3562,N_4198);
xnor U6776 (N_6776,N_4762,N_4403);
nand U6777 (N_6777,N_3138,N_1648);
and U6778 (N_6778,N_2451,N_2210);
or U6779 (N_6779,N_3886,N_4736);
or U6780 (N_6780,N_2346,N_4212);
nor U6781 (N_6781,N_28,N_4134);
nand U6782 (N_6782,N_1449,N_3745);
and U6783 (N_6783,N_4621,N_2994);
and U6784 (N_6784,N_3639,N_284);
xor U6785 (N_6785,N_2169,N_3669);
nand U6786 (N_6786,N_1228,N_733);
nor U6787 (N_6787,N_3836,N_3032);
or U6788 (N_6788,N_4896,N_1396);
nand U6789 (N_6789,N_2641,N_2389);
nor U6790 (N_6790,N_3194,N_1121);
nand U6791 (N_6791,N_3469,N_729);
nand U6792 (N_6792,N_2747,N_2809);
nand U6793 (N_6793,N_4442,N_4275);
nor U6794 (N_6794,N_3994,N_3468);
xnor U6795 (N_6795,N_2628,N_4565);
nor U6796 (N_6796,N_977,N_490);
or U6797 (N_6797,N_254,N_3241);
and U6798 (N_6798,N_744,N_1165);
xor U6799 (N_6799,N_969,N_3010);
and U6800 (N_6800,N_4285,N_3378);
xnor U6801 (N_6801,N_4773,N_2623);
nand U6802 (N_6802,N_1958,N_660);
nand U6803 (N_6803,N_1003,N_591);
or U6804 (N_6804,N_3738,N_3911);
nand U6805 (N_6805,N_2312,N_3018);
nor U6806 (N_6806,N_4675,N_2261);
nor U6807 (N_6807,N_3353,N_342);
and U6808 (N_6808,N_3330,N_1089);
nor U6809 (N_6809,N_160,N_1944);
and U6810 (N_6810,N_4589,N_3514);
or U6811 (N_6811,N_4894,N_3743);
and U6812 (N_6812,N_210,N_355);
or U6813 (N_6813,N_4139,N_27);
xor U6814 (N_6814,N_1573,N_2377);
or U6815 (N_6815,N_4414,N_4083);
nor U6816 (N_6816,N_4445,N_226);
xnor U6817 (N_6817,N_4995,N_3626);
xnor U6818 (N_6818,N_126,N_1571);
nand U6819 (N_6819,N_4768,N_1932);
xnor U6820 (N_6820,N_3035,N_3725);
xnor U6821 (N_6821,N_3893,N_3783);
or U6822 (N_6822,N_1226,N_2128);
and U6823 (N_6823,N_2550,N_3218);
and U6824 (N_6824,N_460,N_3344);
xnor U6825 (N_6825,N_1907,N_788);
nand U6826 (N_6826,N_2237,N_279);
and U6827 (N_6827,N_3071,N_472);
nor U6828 (N_6828,N_4946,N_1961);
or U6829 (N_6829,N_4527,N_4918);
or U6830 (N_6830,N_3611,N_15);
or U6831 (N_6831,N_1681,N_2946);
nor U6832 (N_6832,N_2927,N_1990);
xor U6833 (N_6833,N_2764,N_4547);
nand U6834 (N_6834,N_2719,N_4069);
nor U6835 (N_6835,N_659,N_2449);
nand U6836 (N_6836,N_3894,N_4973);
xor U6837 (N_6837,N_4284,N_3953);
and U6838 (N_6838,N_4586,N_4752);
nor U6839 (N_6839,N_4502,N_1320);
and U6840 (N_6840,N_1268,N_4783);
and U6841 (N_6841,N_4700,N_4232);
nand U6842 (N_6842,N_4151,N_4744);
or U6843 (N_6843,N_2802,N_4493);
or U6844 (N_6844,N_712,N_4306);
xor U6845 (N_6845,N_132,N_4734);
or U6846 (N_6846,N_2969,N_2052);
xnor U6847 (N_6847,N_1637,N_253);
xnor U6848 (N_6848,N_3856,N_2829);
and U6849 (N_6849,N_3303,N_4582);
xor U6850 (N_6850,N_2365,N_1059);
nor U6851 (N_6851,N_2728,N_4905);
nand U6852 (N_6852,N_1899,N_195);
nand U6853 (N_6853,N_4671,N_23);
and U6854 (N_6854,N_3439,N_3160);
xor U6855 (N_6855,N_4223,N_84);
xnor U6856 (N_6856,N_1013,N_2319);
and U6857 (N_6857,N_1430,N_738);
nand U6858 (N_6858,N_3841,N_3361);
and U6859 (N_6859,N_2525,N_2966);
nor U6860 (N_6860,N_4033,N_1627);
nor U6861 (N_6861,N_3198,N_1439);
nand U6862 (N_6862,N_369,N_318);
xnor U6863 (N_6863,N_468,N_1874);
xnor U6864 (N_6864,N_112,N_435);
nand U6865 (N_6865,N_4870,N_9);
xnor U6866 (N_6866,N_2426,N_3398);
or U6867 (N_6867,N_3327,N_4685);
and U6868 (N_6868,N_3155,N_104);
xor U6869 (N_6869,N_155,N_1034);
nor U6870 (N_6870,N_2590,N_3747);
and U6871 (N_6871,N_3926,N_3094);
nand U6872 (N_6872,N_1382,N_47);
nand U6873 (N_6873,N_925,N_17);
nor U6874 (N_6874,N_675,N_1203);
nor U6875 (N_6875,N_2968,N_2);
or U6876 (N_6876,N_4776,N_811);
xnor U6877 (N_6877,N_3265,N_2024);
nor U6878 (N_6878,N_1264,N_1798);
and U6879 (N_6879,N_4761,N_1025);
xnor U6880 (N_6880,N_3089,N_1006);
xor U6881 (N_6881,N_4341,N_1177);
and U6882 (N_6882,N_3621,N_3568);
xnor U6883 (N_6883,N_2474,N_2187);
nand U6884 (N_6884,N_329,N_1233);
xor U6885 (N_6885,N_608,N_909);
nor U6886 (N_6886,N_3617,N_4004);
nor U6887 (N_6887,N_2883,N_593);
or U6888 (N_6888,N_3721,N_3463);
xor U6889 (N_6889,N_2793,N_4126);
xnor U6890 (N_6890,N_2779,N_3301);
or U6891 (N_6891,N_4860,N_1244);
or U6892 (N_6892,N_3714,N_2852);
nand U6893 (N_6893,N_2119,N_547);
or U6894 (N_6894,N_861,N_3374);
nor U6895 (N_6895,N_1222,N_1853);
or U6896 (N_6896,N_1817,N_34);
nand U6897 (N_6897,N_1807,N_918);
or U6898 (N_6898,N_4040,N_1159);
nor U6899 (N_6899,N_2334,N_1151);
nand U6900 (N_6900,N_3167,N_1373);
nor U6901 (N_6901,N_583,N_25);
xor U6902 (N_6902,N_2941,N_3191);
and U6903 (N_6903,N_2337,N_1053);
or U6904 (N_6904,N_399,N_2930);
or U6905 (N_6905,N_2300,N_551);
xnor U6906 (N_6906,N_3174,N_4522);
and U6907 (N_6907,N_2241,N_2073);
nand U6908 (N_6908,N_819,N_3238);
xor U6909 (N_6909,N_2067,N_2439);
xor U6910 (N_6910,N_4023,N_2153);
or U6911 (N_6911,N_209,N_3411);
nand U6912 (N_6912,N_3368,N_4910);
nor U6913 (N_6913,N_3013,N_2595);
or U6914 (N_6914,N_3602,N_797);
nor U6915 (N_6915,N_3251,N_2425);
or U6916 (N_6916,N_4173,N_2588);
or U6917 (N_6917,N_1257,N_1190);
and U6918 (N_6918,N_4949,N_63);
xnor U6919 (N_6919,N_516,N_2730);
nor U6920 (N_6920,N_3846,N_3810);
and U6921 (N_6921,N_2601,N_171);
and U6922 (N_6922,N_3917,N_2955);
nor U6923 (N_6923,N_2604,N_778);
or U6924 (N_6924,N_4369,N_1361);
xnor U6925 (N_6925,N_808,N_3350);
xnor U6926 (N_6926,N_2861,N_484);
xnor U6927 (N_6927,N_3644,N_44);
and U6928 (N_6928,N_1898,N_1075);
or U6929 (N_6929,N_3015,N_2496);
nor U6930 (N_6930,N_1884,N_4524);
or U6931 (N_6931,N_3214,N_357);
or U6932 (N_6932,N_576,N_752);
xnor U6933 (N_6933,N_838,N_2929);
and U6934 (N_6934,N_1342,N_2774);
or U6935 (N_6935,N_2468,N_4156);
and U6936 (N_6936,N_395,N_4836);
nor U6937 (N_6937,N_4147,N_4842);
and U6938 (N_6938,N_4640,N_4434);
or U6939 (N_6939,N_2403,N_2080);
xor U6940 (N_6940,N_2754,N_2600);
nor U6941 (N_6941,N_2306,N_183);
nor U6942 (N_6942,N_2253,N_561);
nor U6943 (N_6943,N_3807,N_2830);
nor U6944 (N_6944,N_2995,N_1836);
or U6945 (N_6945,N_2294,N_4329);
and U6946 (N_6946,N_450,N_4115);
nor U6947 (N_6947,N_1035,N_2594);
nor U6948 (N_6948,N_4440,N_2836);
nor U6949 (N_6949,N_3676,N_2949);
nand U6950 (N_6950,N_4590,N_2042);
nor U6951 (N_6951,N_4020,N_4785);
and U6952 (N_6952,N_152,N_4786);
nor U6953 (N_6953,N_3754,N_2016);
or U6954 (N_6954,N_1911,N_393);
and U6955 (N_6955,N_4430,N_4563);
nor U6956 (N_6956,N_3898,N_4131);
xnor U6957 (N_6957,N_3523,N_3505);
nand U6958 (N_6958,N_2032,N_3913);
xor U6959 (N_6959,N_4272,N_3305);
or U6960 (N_6960,N_1955,N_2472);
nand U6961 (N_6961,N_4459,N_3814);
nand U6962 (N_6962,N_202,N_870);
nand U6963 (N_6963,N_4775,N_2706);
nor U6964 (N_6964,N_4826,N_301);
or U6965 (N_6965,N_2847,N_41);
nand U6966 (N_6966,N_336,N_1757);
xnor U6967 (N_6967,N_3382,N_3905);
or U6968 (N_6968,N_554,N_4352);
and U6969 (N_6969,N_4144,N_1038);
nor U6970 (N_6970,N_185,N_2267);
and U6971 (N_6971,N_4054,N_661);
and U6972 (N_6972,N_2459,N_2766);
nand U6973 (N_6973,N_4097,N_2928);
or U6974 (N_6974,N_987,N_3772);
or U6975 (N_6975,N_2740,N_682);
or U6976 (N_6976,N_2184,N_3389);
nand U6977 (N_6977,N_686,N_3124);
nand U6978 (N_6978,N_2179,N_1780);
and U6979 (N_6979,N_1661,N_1767);
or U6980 (N_6980,N_1896,N_1174);
xor U6981 (N_6981,N_54,N_958);
nand U6982 (N_6982,N_2419,N_259);
or U6983 (N_6983,N_2354,N_2833);
nor U6984 (N_6984,N_879,N_4646);
nand U6985 (N_6985,N_3829,N_3056);
nand U6986 (N_6986,N_3134,N_2713);
or U6987 (N_6987,N_1483,N_1215);
xnor U6988 (N_6988,N_2828,N_2989);
and U6989 (N_6989,N_2100,N_4179);
nor U6990 (N_6990,N_2316,N_3890);
xnor U6991 (N_6991,N_2176,N_3149);
xor U6992 (N_6992,N_3818,N_4024);
and U6993 (N_6993,N_4668,N_1453);
nand U6994 (N_6994,N_3497,N_527);
and U6995 (N_6995,N_2221,N_2511);
xnor U6996 (N_6996,N_4057,N_4902);
xor U6997 (N_6997,N_1052,N_1582);
nor U6998 (N_6998,N_2803,N_4088);
or U6999 (N_6999,N_2760,N_1370);
xnor U7000 (N_7000,N_4877,N_2168);
or U7001 (N_7001,N_328,N_4255);
or U7002 (N_7002,N_1848,N_4418);
and U7003 (N_7003,N_3341,N_900);
or U7004 (N_7004,N_3744,N_4058);
and U7005 (N_7005,N_4879,N_45);
nor U7006 (N_7006,N_1906,N_434);
nand U7007 (N_7007,N_3343,N_3833);
xnor U7008 (N_7008,N_1288,N_1087);
nand U7009 (N_7009,N_2074,N_4213);
or U7010 (N_7010,N_2765,N_3407);
or U7011 (N_7011,N_3896,N_555);
and U7012 (N_7012,N_971,N_1033);
and U7013 (N_7013,N_3243,N_4273);
and U7014 (N_7014,N_1845,N_168);
and U7015 (N_7015,N_119,N_3982);
or U7016 (N_7016,N_276,N_2686);
xor U7017 (N_7017,N_3834,N_1518);
or U7018 (N_7018,N_4540,N_64);
or U7019 (N_7019,N_2091,N_724);
or U7020 (N_7020,N_3930,N_3077);
xnor U7021 (N_7021,N_1458,N_3111);
xnor U7022 (N_7022,N_4439,N_4337);
or U7023 (N_7023,N_4954,N_3731);
xor U7024 (N_7024,N_2432,N_3920);
xnor U7025 (N_7025,N_4692,N_3831);
nand U7026 (N_7026,N_782,N_4857);
or U7027 (N_7027,N_3939,N_2700);
nor U7028 (N_7028,N_1219,N_1750);
and U7029 (N_7029,N_2625,N_2539);
nor U7030 (N_7030,N_4550,N_3453);
nand U7031 (N_7031,N_1551,N_2961);
nor U7032 (N_7032,N_1881,N_2617);
xnor U7033 (N_7033,N_832,N_3223);
nor U7034 (N_7034,N_2182,N_1123);
nor U7035 (N_7035,N_157,N_1626);
xor U7036 (N_7036,N_2497,N_1515);
nor U7037 (N_7037,N_798,N_4462);
xor U7038 (N_7038,N_2202,N_1261);
xor U7039 (N_7039,N_3800,N_130);
or U7040 (N_7040,N_4262,N_1574);
nand U7041 (N_7041,N_1514,N_1741);
and U7042 (N_7042,N_671,N_3179);
xor U7043 (N_7043,N_2892,N_2287);
and U7044 (N_7044,N_4976,N_748);
nor U7045 (N_7045,N_3642,N_1020);
and U7046 (N_7046,N_1585,N_803);
nor U7047 (N_7047,N_3359,N_4267);
nand U7048 (N_7048,N_2619,N_753);
and U7049 (N_7049,N_3498,N_3110);
or U7050 (N_7050,N_403,N_1249);
and U7051 (N_7051,N_72,N_1272);
nand U7052 (N_7052,N_2033,N_4676);
nor U7053 (N_7053,N_563,N_1600);
nand U7054 (N_7054,N_611,N_2960);
and U7055 (N_7055,N_1609,N_4975);
and U7056 (N_7056,N_2062,N_4380);
nand U7057 (N_7057,N_3454,N_2541);
xnor U7058 (N_7058,N_3840,N_4143);
and U7059 (N_7059,N_1823,N_2547);
or U7060 (N_7060,N_2613,N_2044);
nand U7061 (N_7061,N_1474,N_332);
nand U7062 (N_7062,N_416,N_1162);
and U7063 (N_7063,N_390,N_3226);
xnor U7064 (N_7064,N_1610,N_2423);
or U7065 (N_7065,N_1710,N_3555);
nand U7066 (N_7066,N_2392,N_4241);
xor U7067 (N_7067,N_2758,N_4163);
or U7068 (N_7068,N_3386,N_2743);
nor U7069 (N_7069,N_2479,N_4321);
nand U7070 (N_7070,N_1633,N_4733);
and U7071 (N_7071,N_118,N_663);
and U7072 (N_7072,N_3202,N_2697);
or U7073 (N_7073,N_2690,N_1310);
xnor U7074 (N_7074,N_524,N_613);
or U7075 (N_7075,N_3423,N_322);
or U7076 (N_7076,N_1725,N_2177);
and U7077 (N_7077,N_556,N_3113);
xnor U7078 (N_7078,N_4921,N_151);
xor U7079 (N_7079,N_1490,N_3615);
or U7080 (N_7080,N_2323,N_1509);
and U7081 (N_7081,N_2688,N_1138);
or U7082 (N_7082,N_1394,N_3576);
or U7083 (N_7083,N_1407,N_3039);
and U7084 (N_7084,N_4486,N_4886);
or U7085 (N_7085,N_1869,N_1508);
xor U7086 (N_7086,N_2552,N_4704);
and U7087 (N_7087,N_52,N_4268);
nand U7088 (N_7088,N_1726,N_1820);
or U7089 (N_7089,N_83,N_1076);
and U7090 (N_7090,N_4579,N_4545);
nand U7091 (N_7091,N_4560,N_1521);
xor U7092 (N_7092,N_1754,N_3415);
nor U7093 (N_7093,N_1531,N_2181);
or U7094 (N_7094,N_3548,N_3981);
nand U7095 (N_7095,N_2523,N_1595);
nand U7096 (N_7096,N_1598,N_2717);
nand U7097 (N_7097,N_1695,N_893);
or U7098 (N_7098,N_2508,N_597);
nor U7099 (N_7099,N_967,N_3784);
and U7100 (N_7100,N_1982,N_827);
and U7101 (N_7101,N_505,N_1535);
and U7102 (N_7102,N_3349,N_1785);
and U7103 (N_7103,N_1214,N_3799);
nand U7104 (N_7104,N_538,N_4436);
and U7105 (N_7105,N_1663,N_500);
xnor U7106 (N_7106,N_816,N_242);
xor U7107 (N_7107,N_3442,N_1671);
nand U7108 (N_7108,N_4701,N_4513);
xor U7109 (N_7109,N_1827,N_4532);
nand U7110 (N_7110,N_3884,N_4926);
xor U7111 (N_7111,N_1704,N_3491);
or U7112 (N_7112,N_4125,N_1180);
nand U7113 (N_7113,N_4288,N_2003);
nor U7114 (N_7114,N_1702,N_3195);
nand U7115 (N_7115,N_4103,N_354);
xor U7116 (N_7116,N_863,N_1594);
or U7117 (N_7117,N_4472,N_4727);
nand U7118 (N_7118,N_2382,N_4438);
nand U7119 (N_7119,N_1992,N_2219);
nor U7120 (N_7120,N_3156,N_4085);
or U7121 (N_7121,N_1500,N_3563);
or U7122 (N_7122,N_4227,N_1668);
and U7123 (N_7123,N_2322,N_298);
or U7124 (N_7124,N_1316,N_4027);
xnor U7125 (N_7125,N_1891,N_559);
nand U7126 (N_7126,N_2907,N_3409);
and U7127 (N_7127,N_1040,N_3870);
nor U7128 (N_7128,N_2788,N_1227);
and U7129 (N_7129,N_4584,N_1974);
xor U7130 (N_7130,N_471,N_2283);
xnor U7131 (N_7131,N_2869,N_4622);
xnor U7132 (N_7132,N_4592,N_2343);
xnor U7133 (N_7133,N_2997,N_760);
and U7134 (N_7134,N_1393,N_508);
nor U7135 (N_7135,N_1105,N_3058);
xor U7136 (N_7136,N_3447,N_4225);
nor U7137 (N_7137,N_3708,N_2676);
or U7138 (N_7138,N_639,N_214);
nand U7139 (N_7139,N_0,N_1355);
nor U7140 (N_7140,N_3357,N_3976);
or U7141 (N_7141,N_887,N_4623);
xor U7142 (N_7142,N_543,N_2364);
nor U7143 (N_7143,N_3225,N_2801);
nor U7144 (N_7144,N_3078,N_1995);
nand U7145 (N_7145,N_2150,N_2909);
or U7146 (N_7146,N_2586,N_2239);
nor U7147 (N_7147,N_3478,N_4790);
nor U7148 (N_7148,N_3387,N_234);
nor U7149 (N_7149,N_4758,N_3941);
or U7150 (N_7150,N_3733,N_3432);
and U7151 (N_7151,N_1220,N_3471);
nand U7152 (N_7152,N_3847,N_1333);
nor U7153 (N_7153,N_4184,N_4360);
xnor U7154 (N_7154,N_896,N_2501);
nor U7155 (N_7155,N_2068,N_4162);
xnor U7156 (N_7156,N_2329,N_3919);
nand U7157 (N_7157,N_4474,N_719);
and U7158 (N_7158,N_4512,N_3141);
xor U7159 (N_7159,N_3970,N_4732);
xor U7160 (N_7160,N_483,N_4562);
or U7161 (N_7161,N_2475,N_2570);
xnor U7162 (N_7162,N_4292,N_3929);
and U7163 (N_7163,N_4756,N_2707);
nand U7164 (N_7164,N_4674,N_4389);
nor U7165 (N_7165,N_3674,N_330);
nor U7166 (N_7166,N_4141,N_2353);
xor U7167 (N_7167,N_634,N_4228);
nor U7168 (N_7168,N_511,N_2110);
and U7169 (N_7169,N_4135,N_2568);
nand U7170 (N_7170,N_4684,N_4539);
nand U7171 (N_7171,N_4164,N_3422);
nor U7172 (N_7172,N_2384,N_588);
and U7173 (N_7173,N_2635,N_2034);
and U7174 (N_7174,N_3172,N_4264);
nor U7175 (N_7175,N_4997,N_4190);
xor U7176 (N_7176,N_2776,N_2937);
xor U7177 (N_7177,N_1170,N_3024);
xor U7178 (N_7178,N_1765,N_1252);
nor U7179 (N_7179,N_1309,N_383);
nand U7180 (N_7180,N_1764,N_802);
or U7181 (N_7181,N_539,N_3190);
or U7182 (N_7182,N_100,N_1991);
or U7183 (N_7183,N_4244,N_187);
nor U7184 (N_7184,N_624,N_707);
nand U7185 (N_7185,N_319,N_1267);
nand U7186 (N_7186,N_4468,N_4467);
and U7187 (N_7187,N_4356,N_4172);
nor U7188 (N_7188,N_4397,N_1085);
or U7189 (N_7189,N_2775,N_2533);
nand U7190 (N_7190,N_4630,N_4128);
nor U7191 (N_7191,N_377,N_1022);
xnor U7192 (N_7192,N_941,N_1802);
nand U7193 (N_7193,N_2038,N_379);
and U7194 (N_7194,N_4624,N_1833);
or U7195 (N_7195,N_4319,N_2534);
nor U7196 (N_7196,N_2773,N_3114);
and U7197 (N_7197,N_1285,N_1346);
nor U7198 (N_7198,N_4299,N_1666);
xnor U7199 (N_7199,N_459,N_3302);
and U7200 (N_7200,N_4922,N_2506);
xnor U7201 (N_7201,N_3324,N_315);
or U7202 (N_7202,N_1119,N_3832);
and U7203 (N_7203,N_2413,N_3762);
and U7204 (N_7204,N_3654,N_1068);
and U7205 (N_7205,N_3882,N_4618);
or U7206 (N_7206,N_4384,N_2134);
xnor U7207 (N_7207,N_1665,N_4928);
xor U7208 (N_7208,N_476,N_1947);
xnor U7209 (N_7209,N_1179,N_4804);
xor U7210 (N_7210,N_2263,N_4257);
or U7211 (N_7211,N_2327,N_3528);
xor U7212 (N_7212,N_3088,N_3100);
and U7213 (N_7213,N_501,N_864);
or U7214 (N_7214,N_2503,N_4383);
nor U7215 (N_7215,N_3433,N_510);
nor U7216 (N_7216,N_901,N_1012);
and U7217 (N_7217,N_1217,N_2627);
nand U7218 (N_7218,N_4218,N_3105);
or U7219 (N_7219,N_609,N_2772);
and U7220 (N_7220,N_637,N_1811);
or U7221 (N_7221,N_786,N_2096);
nor U7222 (N_7222,N_1004,N_417);
or U7223 (N_7223,N_2050,N_4452);
nor U7224 (N_7224,N_3527,N_1350);
or U7225 (N_7225,N_2230,N_4789);
xnor U7226 (N_7226,N_325,N_1084);
and U7227 (N_7227,N_2360,N_71);
or U7228 (N_7228,N_3596,N_4957);
and U7229 (N_7229,N_4938,N_4376);
xor U7230 (N_7230,N_128,N_4661);
or U7231 (N_7231,N_4663,N_1294);
xnor U7232 (N_7232,N_3401,N_3679);
and U7233 (N_7233,N_3992,N_698);
nand U7234 (N_7234,N_4458,N_3041);
xnor U7235 (N_7235,N_813,N_1029);
and U7236 (N_7236,N_1186,N_882);
and U7237 (N_7237,N_1993,N_3438);
xnor U7238 (N_7238,N_3892,N_4234);
xnor U7239 (N_7239,N_2090,N_521);
nor U7240 (N_7240,N_519,N_1481);
and U7241 (N_7241,N_3531,N_894);
xor U7242 (N_7242,N_4350,N_227);
and U7243 (N_7243,N_4743,N_4933);
nand U7244 (N_7244,N_805,N_4709);
and U7245 (N_7245,N_4693,N_4322);
nor U7246 (N_7246,N_4604,N_2041);
nor U7247 (N_7247,N_2357,N_3354);
or U7248 (N_7248,N_2963,N_3091);
nor U7249 (N_7249,N_1133,N_2109);
or U7250 (N_7250,N_3908,N_2296);
xor U7251 (N_7251,N_2657,N_454);
nand U7252 (N_7252,N_3283,N_3259);
or U7253 (N_7253,N_1451,N_2567);
and U7254 (N_7254,N_428,N_4617);
xnor U7255 (N_7255,N_4181,N_2299);
and U7256 (N_7256,N_4801,N_4446);
and U7257 (N_7257,N_2077,N_360);
or U7258 (N_7258,N_4863,N_1206);
or U7259 (N_7259,N_4557,N_429);
nor U7260 (N_7260,N_4402,N_2885);
and U7261 (N_7261,N_3479,N_842);
and U7262 (N_7262,N_141,N_677);
nand U7263 (N_7263,N_3516,N_1154);
and U7264 (N_7264,N_4250,N_3062);
xor U7265 (N_7265,N_670,N_4138);
or U7266 (N_7266,N_3052,N_3616);
nor U7267 (N_7267,N_4136,N_1234);
or U7268 (N_7268,N_866,N_1116);
nand U7269 (N_7269,N_415,N_1716);
and U7270 (N_7270,N_140,N_2872);
nand U7271 (N_7271,N_3628,N_4373);
and U7272 (N_7272,N_1367,N_1692);
nor U7273 (N_7273,N_4364,N_3740);
and U7274 (N_7274,N_4707,N_596);
xnor U7275 (N_7275,N_1207,N_4861);
or U7276 (N_7276,N_3346,N_747);
or U7277 (N_7277,N_1733,N_2831);
nor U7278 (N_7278,N_916,N_2592);
xnor U7279 (N_7279,N_2452,N_3627);
and U7280 (N_7280,N_2071,N_3256);
nor U7281 (N_7281,N_3969,N_1614);
xnor U7282 (N_7282,N_3337,N_4778);
nor U7283 (N_7283,N_3677,N_2951);
and U7284 (N_7284,N_1399,N_973);
nor U7285 (N_7285,N_3605,N_2795);
xnor U7286 (N_7286,N_1723,N_1652);
or U7287 (N_7287,N_1172,N_75);
xnor U7288 (N_7288,N_3700,N_2931);
and U7289 (N_7289,N_2231,N_1910);
or U7290 (N_7290,N_2655,N_2288);
or U7291 (N_7291,N_2242,N_878);
or U7292 (N_7292,N_374,N_2480);
or U7293 (N_7293,N_4185,N_3735);
and U7294 (N_7294,N_3487,N_2258);
nor U7295 (N_7295,N_3648,N_1403);
nor U7296 (N_7296,N_549,N_3703);
or U7297 (N_7297,N_4595,N_3004);
nor U7298 (N_7298,N_3756,N_4914);
and U7299 (N_7299,N_4799,N_1866);
nand U7300 (N_7300,N_3825,N_2582);
xor U7301 (N_7301,N_2046,N_4171);
and U7302 (N_7302,N_1826,N_517);
or U7303 (N_7303,N_780,N_4731);
nand U7304 (N_7304,N_3539,N_3003);
nor U7305 (N_7305,N_1880,N_3347);
or U7306 (N_7306,N_3526,N_3059);
and U7307 (N_7307,N_4286,N_3424);
xor U7308 (N_7308,N_2844,N_3488);
and U7309 (N_7309,N_3426,N_2371);
or U7310 (N_7310,N_3316,N_2638);
nand U7311 (N_7311,N_240,N_4066);
or U7312 (N_7312,N_2553,N_1204);
or U7313 (N_7313,N_775,N_491);
and U7314 (N_7314,N_3954,N_2320);
xor U7315 (N_7315,N_3112,N_720);
or U7316 (N_7316,N_3435,N_2970);
or U7317 (N_7317,N_2341,N_1315);
or U7318 (N_7318,N_1477,N_1230);
and U7319 (N_7319,N_2375,N_843);
xor U7320 (N_7320,N_3584,N_2342);
and U7321 (N_7321,N_3918,N_176);
or U7322 (N_7322,N_1847,N_3295);
nor U7323 (N_7323,N_3177,N_4013);
or U7324 (N_7324,N_39,N_1273);
or U7325 (N_7325,N_2875,N_31);
or U7326 (N_7326,N_3541,N_2069);
nor U7327 (N_7327,N_2490,N_3474);
and U7328 (N_7328,N_2562,N_1959);
xor U7329 (N_7329,N_291,N_1293);
or U7330 (N_7330,N_2813,N_1416);
or U7331 (N_7331,N_4606,N_3906);
nand U7332 (N_7332,N_3711,N_1606);
nand U7333 (N_7333,N_3945,N_1332);
xor U7334 (N_7334,N_570,N_1987);
nor U7335 (N_7335,N_2640,N_3199);
xor U7336 (N_7336,N_1212,N_2205);
or U7337 (N_7337,N_1111,N_4504);
and U7338 (N_7338,N_640,N_1629);
nand U7339 (N_7339,N_2858,N_2234);
nand U7340 (N_7340,N_1584,N_1857);
nor U7341 (N_7341,N_1463,N_1014);
and U7342 (N_7342,N_148,N_2762);
and U7343 (N_7343,N_2269,N_2476);
and U7344 (N_7344,N_4248,N_2070);
and U7345 (N_7345,N_1635,N_4837);
and U7346 (N_7346,N_2467,N_4221);
nand U7347 (N_7347,N_1137,N_1861);
or U7348 (N_7348,N_404,N_4903);
nand U7349 (N_7349,N_1583,N_1925);
nand U7350 (N_7350,N_4208,N_3873);
xor U7351 (N_7351,N_3521,N_881);
and U7352 (N_7352,N_37,N_2914);
and U7353 (N_7353,N_3692,N_968);
nor U7354 (N_7354,N_4892,N_2835);
nor U7355 (N_7355,N_853,N_667);
or U7356 (N_7356,N_1577,N_2733);
nor U7357 (N_7357,N_3715,N_496);
xnor U7358 (N_7358,N_674,N_855);
and U7359 (N_7359,N_2020,N_3619);
nand U7360 (N_7360,N_642,N_1231);
and U7361 (N_7361,N_3766,N_1748);
and U7362 (N_7362,N_2652,N_3165);
xor U7363 (N_7363,N_2618,N_3122);
xor U7364 (N_7364,N_2897,N_4927);
and U7365 (N_7365,N_451,N_3652);
nand U7366 (N_7366,N_4541,N_976);
xor U7367 (N_7367,N_3877,N_2612);
nand U7368 (N_7368,N_3481,N_2162);
and U7369 (N_7369,N_4680,N_4723);
nor U7370 (N_7370,N_3109,N_3483);
nand U7371 (N_7371,N_3377,N_441);
xor U7372 (N_7372,N_3581,N_1324);
nand U7373 (N_7373,N_3533,N_4774);
xnor U7374 (N_7374,N_2653,N_4342);
xnor U7375 (N_7375,N_4667,N_4361);
nand U7376 (N_7376,N_684,N_1448);
xnor U7377 (N_7377,N_708,N_1559);
nand U7378 (N_7378,N_1384,N_1793);
xor U7379 (N_7379,N_3274,N_1348);
nand U7380 (N_7380,N_272,N_4840);
nor U7381 (N_7381,N_996,N_883);
xnor U7382 (N_7382,N_3455,N_470);
nand U7383 (N_7383,N_1545,N_2114);
and U7384 (N_7384,N_162,N_3631);
or U7385 (N_7385,N_4206,N_4984);
nand U7386 (N_7386,N_4157,N_3458);
and U7387 (N_7387,N_1437,N_2379);
nor U7388 (N_7388,N_3187,N_413);
or U7389 (N_7389,N_860,N_4410);
xnor U7390 (N_7390,N_4186,N_740);
and U7391 (N_7391,N_3332,N_3161);
nor U7392 (N_7392,N_4075,N_4779);
and U7393 (N_7393,N_2599,N_310);
nand U7394 (N_7394,N_1787,N_1781);
and U7395 (N_7395,N_174,N_2702);
nand U7396 (N_7396,N_3543,N_249);
nor U7397 (N_7397,N_4807,N_4298);
nand U7398 (N_7398,N_1239,N_4355);
and U7399 (N_7399,N_3916,N_1479);
or U7400 (N_7400,N_4353,N_1486);
nand U7401 (N_7401,N_2633,N_2045);
and U7402 (N_7402,N_3254,N_4968);
nand U7403 (N_7403,N_919,N_2228);
nor U7404 (N_7404,N_1304,N_4686);
nand U7405 (N_7405,N_2397,N_1419);
nand U7406 (N_7406,N_1892,N_2116);
xor U7407 (N_7407,N_1005,N_2017);
xor U7408 (N_7408,N_566,N_2301);
xor U7409 (N_7409,N_409,N_2244);
nor U7410 (N_7410,N_3298,N_4279);
xor U7411 (N_7411,N_4694,N_2691);
and U7412 (N_7412,N_2870,N_932);
nor U7413 (N_7413,N_3082,N_4796);
nor U7414 (N_7414,N_3049,N_2098);
or U7415 (N_7415,N_1791,N_3757);
or U7416 (N_7416,N_2394,N_1636);
xor U7417 (N_7417,N_1771,N_3205);
nand U7418 (N_7418,N_2349,N_4471);
nand U7419 (N_7419,N_2356,N_4909);
xnor U7420 (N_7420,N_1638,N_746);
and U7421 (N_7421,N_2175,N_3864);
nand U7422 (N_7422,N_1284,N_1580);
or U7423 (N_7423,N_2882,N_699);
or U7424 (N_7424,N_2214,N_1825);
or U7425 (N_7425,N_4475,N_421);
xnor U7426 (N_7426,N_138,N_1903);
and U7427 (N_7427,N_4431,N_1735);
nand U7428 (N_7428,N_3025,N_997);
nor U7429 (N_7429,N_3232,N_1951);
nand U7430 (N_7430,N_341,N_2654);
xnor U7431 (N_7431,N_4757,N_1039);
nor U7432 (N_7432,N_2578,N_219);
and U7433 (N_7433,N_1522,N_3365);
nor U7434 (N_7434,N_4792,N_3547);
and U7435 (N_7435,N_3868,N_3613);
or U7436 (N_7436,N_1904,N_366);
or U7437 (N_7437,N_4070,N_3021);
nand U7438 (N_7438,N_150,N_3219);
and U7439 (N_7439,N_1984,N_2148);
nor U7440 (N_7440,N_1048,N_3650);
or U7441 (N_7441,N_4455,N_2648);
or U7442 (N_7442,N_621,N_1915);
or U7443 (N_7443,N_3136,N_181);
xnor U7444 (N_7444,N_4835,N_3779);
or U7445 (N_7445,N_3671,N_2893);
xor U7446 (N_7446,N_1601,N_4335);
nand U7447 (N_7447,N_3417,N_1792);
nor U7448 (N_7448,N_4247,N_2699);
nor U7449 (N_7449,N_2491,N_3978);
nor U7450 (N_7450,N_3370,N_4276);
and U7451 (N_7451,N_4481,N_1289);
or U7452 (N_7452,N_2289,N_4919);
and U7453 (N_7453,N_3184,N_3746);
nor U7454 (N_7454,N_1517,N_1015);
and U7455 (N_7455,N_1872,N_3590);
or U7456 (N_7456,N_1788,N_1851);
or U7457 (N_7457,N_4495,N_2336);
and U7458 (N_7458,N_926,N_3450);
nor U7459 (N_7459,N_3667,N_4681);
xnor U7460 (N_7460,N_2245,N_3151);
or U7461 (N_7461,N_934,N_4529);
nor U7462 (N_7462,N_2614,N_2709);
and U7463 (N_7463,N_397,N_2814);
nand U7464 (N_7464,N_4637,N_356);
nor U7465 (N_7465,N_186,N_3073);
nor U7466 (N_7466,N_3080,N_3741);
and U7467 (N_7467,N_691,N_485);
nand U7468 (N_7468,N_3657,N_2579);
and U7469 (N_7469,N_4794,N_4603);
nor U7470 (N_7470,N_4080,N_1232);
nand U7471 (N_7471,N_2209,N_657);
and U7472 (N_7472,N_975,N_2832);
nor U7473 (N_7473,N_2820,N_4798);
or U7474 (N_7474,N_3396,N_4614);
xnor U7475 (N_7475,N_1929,N_2189);
nand U7476 (N_7476,N_4454,N_3660);
and U7477 (N_7477,N_4333,N_495);
nor U7478 (N_7478,N_2355,N_4960);
nand U7479 (N_7479,N_3985,N_2996);
or U7480 (N_7480,N_528,N_278);
nor U7481 (N_7481,N_3419,N_3668);
nor U7482 (N_7482,N_1834,N_4005);
xnor U7483 (N_7483,N_1410,N_3990);
nor U7484 (N_7484,N_4913,N_2130);
xor U7485 (N_7485,N_4053,N_236);
or U7486 (N_7486,N_2025,N_4889);
or U7487 (N_7487,N_721,N_1263);
or U7488 (N_7488,N_4716,N_1962);
or U7489 (N_7489,N_985,N_3443);
xor U7490 (N_7490,N_2463,N_1146);
nand U7491 (N_7491,N_2531,N_4888);
and U7492 (N_7492,N_4456,N_1829);
and U7493 (N_7493,N_4987,N_4453);
nor U7494 (N_7494,N_191,N_4378);
nor U7495 (N_7495,N_410,N_1058);
nor U7496 (N_7496,N_1804,N_3765);
nand U7497 (N_7497,N_486,N_1779);
nand U7498 (N_7498,N_4573,N_3801);
nand U7499 (N_7499,N_504,N_4705);
nor U7500 (N_7500,N_1249,N_3054);
and U7501 (N_7501,N_1454,N_2889);
nor U7502 (N_7502,N_3317,N_2179);
xor U7503 (N_7503,N_2487,N_2858);
or U7504 (N_7504,N_1042,N_3376);
xor U7505 (N_7505,N_1593,N_4428);
nand U7506 (N_7506,N_2535,N_104);
nor U7507 (N_7507,N_2364,N_1900);
or U7508 (N_7508,N_4238,N_4771);
and U7509 (N_7509,N_4155,N_3226);
and U7510 (N_7510,N_686,N_64);
or U7511 (N_7511,N_1916,N_1523);
or U7512 (N_7512,N_1991,N_526);
or U7513 (N_7513,N_4719,N_44);
or U7514 (N_7514,N_1869,N_3118);
xnor U7515 (N_7515,N_352,N_2336);
xnor U7516 (N_7516,N_3993,N_4114);
and U7517 (N_7517,N_3014,N_3554);
nand U7518 (N_7518,N_2417,N_838);
or U7519 (N_7519,N_1058,N_2684);
xor U7520 (N_7520,N_739,N_2937);
or U7521 (N_7521,N_2083,N_1428);
and U7522 (N_7522,N_4522,N_2981);
nand U7523 (N_7523,N_1033,N_2887);
and U7524 (N_7524,N_1558,N_911);
and U7525 (N_7525,N_1199,N_15);
and U7526 (N_7526,N_2783,N_1727);
nand U7527 (N_7527,N_3751,N_1099);
and U7528 (N_7528,N_1395,N_1274);
nor U7529 (N_7529,N_1499,N_3623);
xnor U7530 (N_7530,N_3583,N_4433);
nand U7531 (N_7531,N_3803,N_1996);
nor U7532 (N_7532,N_1496,N_1305);
nand U7533 (N_7533,N_214,N_926);
nor U7534 (N_7534,N_3721,N_1743);
or U7535 (N_7535,N_4841,N_2887);
or U7536 (N_7536,N_4906,N_1922);
xor U7537 (N_7537,N_412,N_3536);
nor U7538 (N_7538,N_3931,N_2282);
nand U7539 (N_7539,N_2393,N_3425);
nand U7540 (N_7540,N_3265,N_4758);
nand U7541 (N_7541,N_1960,N_4351);
nor U7542 (N_7542,N_378,N_2855);
nor U7543 (N_7543,N_2870,N_3833);
nor U7544 (N_7544,N_280,N_312);
nand U7545 (N_7545,N_2547,N_3394);
or U7546 (N_7546,N_4823,N_1999);
nand U7547 (N_7547,N_2577,N_4790);
nor U7548 (N_7548,N_1358,N_2141);
xor U7549 (N_7549,N_2253,N_4917);
or U7550 (N_7550,N_2404,N_534);
xor U7551 (N_7551,N_30,N_3740);
nand U7552 (N_7552,N_2839,N_4683);
and U7553 (N_7553,N_463,N_3270);
nor U7554 (N_7554,N_366,N_807);
xnor U7555 (N_7555,N_4541,N_539);
and U7556 (N_7556,N_289,N_67);
and U7557 (N_7557,N_463,N_1414);
and U7558 (N_7558,N_18,N_1297);
nand U7559 (N_7559,N_174,N_2154);
and U7560 (N_7560,N_1061,N_21);
nor U7561 (N_7561,N_2985,N_4432);
and U7562 (N_7562,N_2984,N_4528);
and U7563 (N_7563,N_4703,N_875);
and U7564 (N_7564,N_4591,N_4666);
or U7565 (N_7565,N_2517,N_3356);
or U7566 (N_7566,N_2119,N_369);
nor U7567 (N_7567,N_4469,N_1552);
xor U7568 (N_7568,N_4615,N_2245);
xnor U7569 (N_7569,N_484,N_2640);
xor U7570 (N_7570,N_2996,N_773);
nand U7571 (N_7571,N_236,N_4314);
nand U7572 (N_7572,N_3959,N_2949);
and U7573 (N_7573,N_494,N_622);
nor U7574 (N_7574,N_1011,N_4092);
or U7575 (N_7575,N_1227,N_3139);
nor U7576 (N_7576,N_452,N_4237);
and U7577 (N_7577,N_663,N_2388);
nor U7578 (N_7578,N_892,N_4946);
or U7579 (N_7579,N_3488,N_959);
xnor U7580 (N_7580,N_430,N_3722);
nand U7581 (N_7581,N_2575,N_4433);
xor U7582 (N_7582,N_1593,N_4291);
and U7583 (N_7583,N_150,N_891);
and U7584 (N_7584,N_64,N_2196);
and U7585 (N_7585,N_4885,N_4474);
and U7586 (N_7586,N_527,N_3924);
or U7587 (N_7587,N_1727,N_2833);
nor U7588 (N_7588,N_2954,N_4346);
nor U7589 (N_7589,N_2994,N_1540);
or U7590 (N_7590,N_464,N_758);
or U7591 (N_7591,N_1206,N_724);
nor U7592 (N_7592,N_3243,N_4973);
or U7593 (N_7593,N_4581,N_115);
xnor U7594 (N_7594,N_2601,N_1083);
nor U7595 (N_7595,N_4415,N_1374);
xnor U7596 (N_7596,N_894,N_3195);
xor U7597 (N_7597,N_1244,N_546);
nor U7598 (N_7598,N_3435,N_885);
xor U7599 (N_7599,N_2230,N_4862);
nor U7600 (N_7600,N_2901,N_427);
or U7601 (N_7601,N_566,N_3058);
and U7602 (N_7602,N_3449,N_4104);
and U7603 (N_7603,N_3975,N_4935);
nand U7604 (N_7604,N_1075,N_595);
and U7605 (N_7605,N_1733,N_2072);
xor U7606 (N_7606,N_4038,N_359);
and U7607 (N_7607,N_1997,N_4835);
nand U7608 (N_7608,N_838,N_3950);
or U7609 (N_7609,N_2092,N_3398);
or U7610 (N_7610,N_4868,N_2325);
nand U7611 (N_7611,N_25,N_4786);
nand U7612 (N_7612,N_360,N_4335);
nor U7613 (N_7613,N_263,N_3073);
xor U7614 (N_7614,N_873,N_2685);
and U7615 (N_7615,N_2096,N_1719);
and U7616 (N_7616,N_841,N_2169);
nor U7617 (N_7617,N_2690,N_253);
xnor U7618 (N_7618,N_2520,N_3781);
or U7619 (N_7619,N_2641,N_4433);
and U7620 (N_7620,N_2255,N_4853);
and U7621 (N_7621,N_1994,N_348);
or U7622 (N_7622,N_4297,N_2225);
xnor U7623 (N_7623,N_4587,N_4268);
or U7624 (N_7624,N_2227,N_3571);
nor U7625 (N_7625,N_501,N_1490);
and U7626 (N_7626,N_443,N_521);
or U7627 (N_7627,N_3752,N_2209);
nand U7628 (N_7628,N_3930,N_769);
or U7629 (N_7629,N_24,N_2604);
nor U7630 (N_7630,N_1141,N_1639);
xnor U7631 (N_7631,N_3215,N_3065);
nor U7632 (N_7632,N_2831,N_846);
or U7633 (N_7633,N_1823,N_3340);
nand U7634 (N_7634,N_510,N_2676);
and U7635 (N_7635,N_4825,N_2060);
xor U7636 (N_7636,N_820,N_3406);
or U7637 (N_7637,N_2041,N_73);
and U7638 (N_7638,N_468,N_972);
and U7639 (N_7639,N_796,N_3731);
xnor U7640 (N_7640,N_2588,N_3900);
xnor U7641 (N_7641,N_229,N_955);
nand U7642 (N_7642,N_3405,N_2277);
nor U7643 (N_7643,N_1145,N_2675);
or U7644 (N_7644,N_4215,N_2990);
nor U7645 (N_7645,N_1934,N_3298);
xor U7646 (N_7646,N_4644,N_1112);
nand U7647 (N_7647,N_1869,N_730);
nor U7648 (N_7648,N_4203,N_2625);
nor U7649 (N_7649,N_1606,N_1684);
nand U7650 (N_7650,N_3465,N_2486);
and U7651 (N_7651,N_4623,N_3780);
and U7652 (N_7652,N_4938,N_869);
nand U7653 (N_7653,N_1301,N_1152);
nor U7654 (N_7654,N_276,N_1289);
and U7655 (N_7655,N_980,N_4010);
or U7656 (N_7656,N_1065,N_2391);
and U7657 (N_7657,N_4757,N_3287);
xnor U7658 (N_7658,N_2912,N_4519);
and U7659 (N_7659,N_311,N_1552);
or U7660 (N_7660,N_2876,N_1042);
or U7661 (N_7661,N_1168,N_3941);
nand U7662 (N_7662,N_1179,N_3526);
and U7663 (N_7663,N_4347,N_2297);
nor U7664 (N_7664,N_2823,N_857);
or U7665 (N_7665,N_2318,N_919);
or U7666 (N_7666,N_4573,N_1303);
nor U7667 (N_7667,N_2929,N_3025);
or U7668 (N_7668,N_1517,N_4511);
xor U7669 (N_7669,N_4574,N_3925);
and U7670 (N_7670,N_3291,N_431);
nor U7671 (N_7671,N_3656,N_1787);
or U7672 (N_7672,N_3293,N_918);
xor U7673 (N_7673,N_1672,N_4566);
or U7674 (N_7674,N_2469,N_4959);
nand U7675 (N_7675,N_4306,N_2280);
or U7676 (N_7676,N_1959,N_2446);
or U7677 (N_7677,N_3126,N_1505);
or U7678 (N_7678,N_4771,N_1384);
and U7679 (N_7679,N_4471,N_2985);
and U7680 (N_7680,N_2666,N_3111);
and U7681 (N_7681,N_861,N_4226);
nand U7682 (N_7682,N_4463,N_1589);
or U7683 (N_7683,N_1780,N_1443);
and U7684 (N_7684,N_42,N_3557);
and U7685 (N_7685,N_4116,N_4205);
nor U7686 (N_7686,N_1818,N_494);
and U7687 (N_7687,N_1648,N_3018);
nor U7688 (N_7688,N_1604,N_2331);
nor U7689 (N_7689,N_4467,N_3194);
and U7690 (N_7690,N_2198,N_1417);
xnor U7691 (N_7691,N_4163,N_620);
nand U7692 (N_7692,N_3890,N_404);
nor U7693 (N_7693,N_3807,N_2590);
xnor U7694 (N_7694,N_819,N_4981);
xor U7695 (N_7695,N_288,N_1209);
xnor U7696 (N_7696,N_918,N_3254);
nand U7697 (N_7697,N_719,N_3787);
or U7698 (N_7698,N_1454,N_1285);
and U7699 (N_7699,N_674,N_3499);
or U7700 (N_7700,N_3590,N_696);
and U7701 (N_7701,N_1041,N_1621);
and U7702 (N_7702,N_1479,N_2232);
xor U7703 (N_7703,N_1838,N_1159);
xor U7704 (N_7704,N_1260,N_374);
and U7705 (N_7705,N_4155,N_4898);
or U7706 (N_7706,N_3795,N_4898);
nor U7707 (N_7707,N_2103,N_1147);
nor U7708 (N_7708,N_2574,N_1044);
and U7709 (N_7709,N_2459,N_379);
or U7710 (N_7710,N_4167,N_1819);
nand U7711 (N_7711,N_1117,N_2710);
and U7712 (N_7712,N_3988,N_3469);
or U7713 (N_7713,N_3321,N_3044);
xor U7714 (N_7714,N_3583,N_1742);
xor U7715 (N_7715,N_4420,N_576);
nand U7716 (N_7716,N_3006,N_231);
or U7717 (N_7717,N_4001,N_2898);
nand U7718 (N_7718,N_4329,N_3735);
nand U7719 (N_7719,N_1437,N_890);
or U7720 (N_7720,N_2525,N_4697);
nand U7721 (N_7721,N_3344,N_4081);
nand U7722 (N_7722,N_3307,N_782);
and U7723 (N_7723,N_4085,N_3893);
and U7724 (N_7724,N_2213,N_3478);
xnor U7725 (N_7725,N_1564,N_2151);
or U7726 (N_7726,N_1237,N_2148);
nor U7727 (N_7727,N_4703,N_4504);
nor U7728 (N_7728,N_4611,N_2813);
nand U7729 (N_7729,N_2565,N_213);
nor U7730 (N_7730,N_2315,N_470);
or U7731 (N_7731,N_1616,N_3280);
and U7732 (N_7732,N_1341,N_4687);
and U7733 (N_7733,N_136,N_4567);
nor U7734 (N_7734,N_984,N_2080);
xnor U7735 (N_7735,N_3370,N_2829);
and U7736 (N_7736,N_808,N_171);
nor U7737 (N_7737,N_771,N_4677);
nand U7738 (N_7738,N_284,N_2011);
xnor U7739 (N_7739,N_3992,N_1778);
xor U7740 (N_7740,N_4538,N_2057);
and U7741 (N_7741,N_3175,N_4896);
nand U7742 (N_7742,N_1358,N_2902);
and U7743 (N_7743,N_3181,N_4105);
nor U7744 (N_7744,N_126,N_3472);
and U7745 (N_7745,N_308,N_3512);
xor U7746 (N_7746,N_1165,N_1869);
and U7747 (N_7747,N_2172,N_2564);
and U7748 (N_7748,N_722,N_440);
nand U7749 (N_7749,N_4453,N_4684);
or U7750 (N_7750,N_3348,N_1807);
xor U7751 (N_7751,N_4410,N_3754);
or U7752 (N_7752,N_2566,N_171);
nand U7753 (N_7753,N_4924,N_3222);
or U7754 (N_7754,N_3883,N_3895);
nor U7755 (N_7755,N_4741,N_1006);
and U7756 (N_7756,N_516,N_3193);
xnor U7757 (N_7757,N_3410,N_3047);
nand U7758 (N_7758,N_1699,N_1674);
or U7759 (N_7759,N_4420,N_3811);
or U7760 (N_7760,N_3701,N_3412);
nand U7761 (N_7761,N_2496,N_1028);
xor U7762 (N_7762,N_3606,N_3019);
nor U7763 (N_7763,N_224,N_893);
or U7764 (N_7764,N_832,N_4699);
nor U7765 (N_7765,N_3942,N_340);
nor U7766 (N_7766,N_1698,N_3491);
nor U7767 (N_7767,N_3557,N_713);
xnor U7768 (N_7768,N_1090,N_540);
xor U7769 (N_7769,N_3847,N_1550);
nor U7770 (N_7770,N_4618,N_632);
and U7771 (N_7771,N_4124,N_358);
or U7772 (N_7772,N_1486,N_2285);
or U7773 (N_7773,N_2294,N_1555);
and U7774 (N_7774,N_2846,N_968);
or U7775 (N_7775,N_1067,N_1936);
or U7776 (N_7776,N_4573,N_4265);
nor U7777 (N_7777,N_828,N_1740);
or U7778 (N_7778,N_3791,N_155);
or U7779 (N_7779,N_1483,N_3889);
nor U7780 (N_7780,N_3409,N_3892);
nor U7781 (N_7781,N_173,N_1503);
or U7782 (N_7782,N_2246,N_4253);
nand U7783 (N_7783,N_4689,N_2635);
or U7784 (N_7784,N_2466,N_2211);
and U7785 (N_7785,N_3649,N_3574);
nor U7786 (N_7786,N_2832,N_4248);
xnor U7787 (N_7787,N_2726,N_2748);
xnor U7788 (N_7788,N_3504,N_3814);
nand U7789 (N_7789,N_2298,N_1521);
or U7790 (N_7790,N_2214,N_1156);
or U7791 (N_7791,N_3824,N_224);
nand U7792 (N_7792,N_4612,N_953);
nand U7793 (N_7793,N_4480,N_3194);
nor U7794 (N_7794,N_1389,N_574);
or U7795 (N_7795,N_4846,N_4927);
xor U7796 (N_7796,N_1026,N_2974);
nor U7797 (N_7797,N_2572,N_356);
and U7798 (N_7798,N_3068,N_866);
and U7799 (N_7799,N_833,N_360);
nor U7800 (N_7800,N_3082,N_1936);
nor U7801 (N_7801,N_1682,N_3618);
nor U7802 (N_7802,N_1371,N_2302);
or U7803 (N_7803,N_1451,N_1999);
nand U7804 (N_7804,N_1417,N_3517);
nor U7805 (N_7805,N_3612,N_357);
and U7806 (N_7806,N_3325,N_1341);
nor U7807 (N_7807,N_4029,N_4579);
or U7808 (N_7808,N_713,N_4354);
and U7809 (N_7809,N_1475,N_2884);
nor U7810 (N_7810,N_4825,N_809);
nor U7811 (N_7811,N_4524,N_2120);
or U7812 (N_7812,N_1519,N_4346);
or U7813 (N_7813,N_2177,N_3700);
xnor U7814 (N_7814,N_2823,N_541);
and U7815 (N_7815,N_1538,N_3825);
nand U7816 (N_7816,N_3072,N_3731);
and U7817 (N_7817,N_519,N_4235);
nor U7818 (N_7818,N_933,N_2918);
or U7819 (N_7819,N_741,N_2041);
or U7820 (N_7820,N_2354,N_4986);
xor U7821 (N_7821,N_4724,N_405);
nor U7822 (N_7822,N_2931,N_3971);
xor U7823 (N_7823,N_376,N_73);
nand U7824 (N_7824,N_2865,N_3617);
xnor U7825 (N_7825,N_3527,N_1459);
or U7826 (N_7826,N_4009,N_1826);
and U7827 (N_7827,N_2981,N_3453);
and U7828 (N_7828,N_3938,N_829);
and U7829 (N_7829,N_3850,N_2389);
xor U7830 (N_7830,N_1223,N_2660);
or U7831 (N_7831,N_4882,N_2157);
nor U7832 (N_7832,N_3694,N_4779);
nor U7833 (N_7833,N_2796,N_813);
nand U7834 (N_7834,N_2564,N_4613);
xnor U7835 (N_7835,N_2890,N_1555);
or U7836 (N_7836,N_4881,N_300);
nand U7837 (N_7837,N_4745,N_3023);
nor U7838 (N_7838,N_575,N_2301);
and U7839 (N_7839,N_4229,N_999);
nor U7840 (N_7840,N_2638,N_103);
nor U7841 (N_7841,N_3365,N_561);
xor U7842 (N_7842,N_3215,N_2599);
nand U7843 (N_7843,N_4900,N_2131);
nor U7844 (N_7844,N_1559,N_2385);
xor U7845 (N_7845,N_2563,N_2241);
xor U7846 (N_7846,N_3877,N_961);
and U7847 (N_7847,N_1665,N_2770);
nand U7848 (N_7848,N_190,N_82);
or U7849 (N_7849,N_1528,N_1952);
and U7850 (N_7850,N_70,N_3539);
and U7851 (N_7851,N_662,N_2882);
nand U7852 (N_7852,N_2691,N_3578);
nand U7853 (N_7853,N_4599,N_501);
xnor U7854 (N_7854,N_1336,N_1462);
nand U7855 (N_7855,N_3791,N_1047);
and U7856 (N_7856,N_712,N_3107);
or U7857 (N_7857,N_4606,N_3502);
xor U7858 (N_7858,N_1473,N_1690);
nand U7859 (N_7859,N_4208,N_4897);
and U7860 (N_7860,N_4203,N_4291);
nor U7861 (N_7861,N_2536,N_1803);
or U7862 (N_7862,N_50,N_2531);
and U7863 (N_7863,N_1093,N_2317);
nor U7864 (N_7864,N_2384,N_1113);
nor U7865 (N_7865,N_3538,N_3725);
nor U7866 (N_7866,N_4149,N_153);
nor U7867 (N_7867,N_3485,N_3107);
xnor U7868 (N_7868,N_238,N_619);
or U7869 (N_7869,N_4923,N_4201);
and U7870 (N_7870,N_976,N_4741);
nand U7871 (N_7871,N_3881,N_4408);
and U7872 (N_7872,N_2558,N_4434);
or U7873 (N_7873,N_1863,N_522);
nor U7874 (N_7874,N_1243,N_3070);
and U7875 (N_7875,N_749,N_4714);
or U7876 (N_7876,N_3110,N_2754);
nand U7877 (N_7877,N_3734,N_1662);
nand U7878 (N_7878,N_213,N_3453);
or U7879 (N_7879,N_1540,N_4242);
nor U7880 (N_7880,N_4754,N_2781);
and U7881 (N_7881,N_1847,N_3219);
nor U7882 (N_7882,N_1603,N_568);
xnor U7883 (N_7883,N_18,N_1696);
and U7884 (N_7884,N_3085,N_4032);
or U7885 (N_7885,N_1621,N_4167);
and U7886 (N_7886,N_3188,N_954);
and U7887 (N_7887,N_1939,N_4706);
or U7888 (N_7888,N_2444,N_3518);
or U7889 (N_7889,N_4416,N_2061);
nand U7890 (N_7890,N_3320,N_2738);
and U7891 (N_7891,N_2687,N_129);
and U7892 (N_7892,N_2648,N_2984);
or U7893 (N_7893,N_2080,N_3260);
nand U7894 (N_7894,N_2218,N_1614);
nor U7895 (N_7895,N_2037,N_2297);
xor U7896 (N_7896,N_4294,N_1320);
or U7897 (N_7897,N_2206,N_2820);
nand U7898 (N_7898,N_1297,N_1810);
nand U7899 (N_7899,N_3805,N_3051);
and U7900 (N_7900,N_711,N_784);
xor U7901 (N_7901,N_3112,N_4592);
or U7902 (N_7902,N_2487,N_2646);
nand U7903 (N_7903,N_4316,N_3209);
nor U7904 (N_7904,N_2815,N_2941);
nand U7905 (N_7905,N_3904,N_2041);
nand U7906 (N_7906,N_431,N_1829);
xnor U7907 (N_7907,N_3688,N_2710);
nor U7908 (N_7908,N_577,N_3233);
xnor U7909 (N_7909,N_4737,N_971);
nand U7910 (N_7910,N_3406,N_1692);
nand U7911 (N_7911,N_1740,N_3201);
xor U7912 (N_7912,N_4798,N_1856);
nand U7913 (N_7913,N_1372,N_2522);
or U7914 (N_7914,N_2236,N_2290);
nor U7915 (N_7915,N_4712,N_4278);
xnor U7916 (N_7916,N_4921,N_1575);
xor U7917 (N_7917,N_324,N_1330);
and U7918 (N_7918,N_3597,N_4749);
xnor U7919 (N_7919,N_4102,N_2393);
and U7920 (N_7920,N_3492,N_469);
or U7921 (N_7921,N_1296,N_1185);
nand U7922 (N_7922,N_1056,N_4976);
nand U7923 (N_7923,N_669,N_309);
xnor U7924 (N_7924,N_2569,N_4024);
and U7925 (N_7925,N_26,N_870);
and U7926 (N_7926,N_523,N_1950);
xor U7927 (N_7927,N_4154,N_2471);
nand U7928 (N_7928,N_2125,N_2593);
nor U7929 (N_7929,N_2331,N_1633);
nor U7930 (N_7930,N_480,N_1393);
nand U7931 (N_7931,N_1512,N_4746);
xor U7932 (N_7932,N_3442,N_790);
xor U7933 (N_7933,N_1330,N_2626);
nand U7934 (N_7934,N_4918,N_3570);
nand U7935 (N_7935,N_2535,N_4702);
nor U7936 (N_7936,N_2458,N_1248);
nand U7937 (N_7937,N_1378,N_3300);
or U7938 (N_7938,N_4837,N_220);
nor U7939 (N_7939,N_2510,N_3776);
nor U7940 (N_7940,N_1458,N_3454);
or U7941 (N_7941,N_90,N_816);
nor U7942 (N_7942,N_4359,N_414);
xnor U7943 (N_7943,N_3471,N_855);
nor U7944 (N_7944,N_1949,N_4123);
nand U7945 (N_7945,N_230,N_1949);
xnor U7946 (N_7946,N_4184,N_2221);
nor U7947 (N_7947,N_925,N_3328);
nand U7948 (N_7948,N_3205,N_4141);
and U7949 (N_7949,N_1101,N_4603);
and U7950 (N_7950,N_1353,N_2310);
or U7951 (N_7951,N_4821,N_726);
or U7952 (N_7952,N_3741,N_1134);
xor U7953 (N_7953,N_610,N_586);
nand U7954 (N_7954,N_1535,N_2638);
xnor U7955 (N_7955,N_1177,N_1584);
or U7956 (N_7956,N_3978,N_3396);
nor U7957 (N_7957,N_2547,N_2258);
nor U7958 (N_7958,N_3495,N_335);
xnor U7959 (N_7959,N_2222,N_63);
nand U7960 (N_7960,N_3177,N_380);
xor U7961 (N_7961,N_2572,N_3811);
and U7962 (N_7962,N_830,N_3010);
nand U7963 (N_7963,N_3532,N_760);
or U7964 (N_7964,N_767,N_2462);
or U7965 (N_7965,N_1744,N_3736);
nor U7966 (N_7966,N_4085,N_2303);
xor U7967 (N_7967,N_3414,N_4932);
or U7968 (N_7968,N_2526,N_633);
nand U7969 (N_7969,N_3706,N_503);
nor U7970 (N_7970,N_836,N_4825);
or U7971 (N_7971,N_575,N_4888);
nand U7972 (N_7972,N_3355,N_4552);
and U7973 (N_7973,N_3163,N_2798);
nor U7974 (N_7974,N_232,N_176);
or U7975 (N_7975,N_2600,N_4981);
or U7976 (N_7976,N_3739,N_2266);
xnor U7977 (N_7977,N_4836,N_2651);
or U7978 (N_7978,N_4729,N_2784);
nor U7979 (N_7979,N_1192,N_3776);
or U7980 (N_7980,N_4590,N_3017);
or U7981 (N_7981,N_3532,N_4908);
or U7982 (N_7982,N_3078,N_870);
nor U7983 (N_7983,N_925,N_4172);
nor U7984 (N_7984,N_2148,N_1978);
or U7985 (N_7985,N_1281,N_4528);
nand U7986 (N_7986,N_709,N_3220);
and U7987 (N_7987,N_4822,N_1607);
nand U7988 (N_7988,N_1520,N_2864);
nand U7989 (N_7989,N_2977,N_369);
nor U7990 (N_7990,N_3379,N_3983);
or U7991 (N_7991,N_2274,N_2827);
nor U7992 (N_7992,N_732,N_4226);
nor U7993 (N_7993,N_2416,N_4116);
and U7994 (N_7994,N_4048,N_800);
nor U7995 (N_7995,N_4346,N_3719);
nand U7996 (N_7996,N_3632,N_391);
and U7997 (N_7997,N_3106,N_652);
xnor U7998 (N_7998,N_2256,N_2197);
and U7999 (N_7999,N_1862,N_1987);
nand U8000 (N_8000,N_91,N_3973);
nor U8001 (N_8001,N_3210,N_1017);
nor U8002 (N_8002,N_2118,N_4544);
or U8003 (N_8003,N_2634,N_405);
nand U8004 (N_8004,N_1313,N_1917);
and U8005 (N_8005,N_3495,N_1629);
nand U8006 (N_8006,N_2758,N_2772);
and U8007 (N_8007,N_3927,N_1815);
or U8008 (N_8008,N_4503,N_4091);
or U8009 (N_8009,N_2541,N_4238);
or U8010 (N_8010,N_2576,N_2927);
nor U8011 (N_8011,N_1896,N_1102);
and U8012 (N_8012,N_3077,N_4357);
and U8013 (N_8013,N_3433,N_4155);
nand U8014 (N_8014,N_3934,N_711);
nand U8015 (N_8015,N_1691,N_56);
and U8016 (N_8016,N_128,N_2486);
xnor U8017 (N_8017,N_2633,N_393);
and U8018 (N_8018,N_2438,N_1250);
nor U8019 (N_8019,N_4359,N_3078);
or U8020 (N_8020,N_3805,N_4929);
or U8021 (N_8021,N_2149,N_837);
xor U8022 (N_8022,N_2386,N_4309);
xnor U8023 (N_8023,N_3104,N_1828);
and U8024 (N_8024,N_2074,N_687);
xor U8025 (N_8025,N_1230,N_2707);
nor U8026 (N_8026,N_1121,N_1755);
and U8027 (N_8027,N_4475,N_2421);
xnor U8028 (N_8028,N_4519,N_2989);
and U8029 (N_8029,N_2011,N_689);
and U8030 (N_8030,N_259,N_4149);
and U8031 (N_8031,N_4671,N_2469);
xor U8032 (N_8032,N_3354,N_2090);
and U8033 (N_8033,N_3739,N_310);
or U8034 (N_8034,N_3115,N_4782);
and U8035 (N_8035,N_972,N_4026);
nand U8036 (N_8036,N_725,N_1234);
xor U8037 (N_8037,N_537,N_305);
nand U8038 (N_8038,N_72,N_1498);
nand U8039 (N_8039,N_2349,N_2152);
nor U8040 (N_8040,N_1785,N_3117);
and U8041 (N_8041,N_4358,N_759);
nand U8042 (N_8042,N_2867,N_3182);
and U8043 (N_8043,N_496,N_3370);
nand U8044 (N_8044,N_3206,N_1596);
or U8045 (N_8045,N_4118,N_2061);
nor U8046 (N_8046,N_1136,N_1991);
nand U8047 (N_8047,N_4299,N_1490);
nand U8048 (N_8048,N_3238,N_87);
xnor U8049 (N_8049,N_1398,N_1367);
xor U8050 (N_8050,N_4818,N_3294);
nor U8051 (N_8051,N_1554,N_3848);
nor U8052 (N_8052,N_2583,N_2497);
nand U8053 (N_8053,N_2899,N_2261);
nand U8054 (N_8054,N_2801,N_1107);
xor U8055 (N_8055,N_949,N_570);
nor U8056 (N_8056,N_4075,N_3838);
nor U8057 (N_8057,N_3910,N_2303);
xnor U8058 (N_8058,N_1010,N_4182);
and U8059 (N_8059,N_1596,N_72);
xor U8060 (N_8060,N_2510,N_405);
xor U8061 (N_8061,N_3483,N_416);
xor U8062 (N_8062,N_3262,N_2498);
or U8063 (N_8063,N_2420,N_3095);
xnor U8064 (N_8064,N_148,N_4306);
xor U8065 (N_8065,N_605,N_4684);
xnor U8066 (N_8066,N_2446,N_2260);
nand U8067 (N_8067,N_3285,N_4754);
and U8068 (N_8068,N_3350,N_526);
and U8069 (N_8069,N_4839,N_4366);
xnor U8070 (N_8070,N_2185,N_3186);
and U8071 (N_8071,N_3362,N_4037);
nor U8072 (N_8072,N_4703,N_366);
nor U8073 (N_8073,N_3356,N_1768);
nor U8074 (N_8074,N_504,N_691);
nand U8075 (N_8075,N_3682,N_2441);
or U8076 (N_8076,N_2509,N_3402);
nor U8077 (N_8077,N_4827,N_233);
or U8078 (N_8078,N_668,N_1405);
or U8079 (N_8079,N_797,N_11);
nor U8080 (N_8080,N_155,N_4856);
xor U8081 (N_8081,N_2455,N_2580);
and U8082 (N_8082,N_1092,N_4411);
nand U8083 (N_8083,N_2430,N_3197);
or U8084 (N_8084,N_278,N_2281);
nand U8085 (N_8085,N_4463,N_437);
and U8086 (N_8086,N_2412,N_2191);
and U8087 (N_8087,N_2828,N_4756);
xor U8088 (N_8088,N_4910,N_353);
nand U8089 (N_8089,N_2239,N_1055);
xor U8090 (N_8090,N_955,N_3632);
nor U8091 (N_8091,N_37,N_3858);
nand U8092 (N_8092,N_2280,N_3772);
or U8093 (N_8093,N_1094,N_4158);
and U8094 (N_8094,N_1025,N_2177);
nand U8095 (N_8095,N_2877,N_1601);
xor U8096 (N_8096,N_2364,N_3117);
nor U8097 (N_8097,N_312,N_3104);
nand U8098 (N_8098,N_2735,N_3859);
nor U8099 (N_8099,N_1713,N_2079);
or U8100 (N_8100,N_4145,N_471);
nor U8101 (N_8101,N_3596,N_752);
or U8102 (N_8102,N_607,N_3599);
and U8103 (N_8103,N_2273,N_1498);
or U8104 (N_8104,N_1351,N_4140);
or U8105 (N_8105,N_2358,N_2473);
xnor U8106 (N_8106,N_2315,N_2474);
nand U8107 (N_8107,N_3937,N_3965);
xor U8108 (N_8108,N_499,N_4068);
and U8109 (N_8109,N_1488,N_4610);
or U8110 (N_8110,N_4906,N_4875);
nand U8111 (N_8111,N_4736,N_3767);
and U8112 (N_8112,N_2495,N_3917);
and U8113 (N_8113,N_836,N_1166);
xnor U8114 (N_8114,N_2901,N_156);
xor U8115 (N_8115,N_977,N_2277);
xnor U8116 (N_8116,N_3586,N_1364);
xnor U8117 (N_8117,N_3618,N_2642);
nand U8118 (N_8118,N_3777,N_2162);
and U8119 (N_8119,N_2025,N_2722);
nor U8120 (N_8120,N_2234,N_1446);
and U8121 (N_8121,N_2299,N_768);
xor U8122 (N_8122,N_1719,N_3159);
nor U8123 (N_8123,N_2613,N_654);
and U8124 (N_8124,N_3086,N_4536);
nor U8125 (N_8125,N_2293,N_2864);
and U8126 (N_8126,N_3478,N_4391);
xnor U8127 (N_8127,N_3100,N_1919);
nand U8128 (N_8128,N_1946,N_2910);
xnor U8129 (N_8129,N_810,N_2711);
and U8130 (N_8130,N_3834,N_565);
or U8131 (N_8131,N_4734,N_4649);
nor U8132 (N_8132,N_3801,N_3434);
nor U8133 (N_8133,N_1866,N_3308);
and U8134 (N_8134,N_3255,N_4011);
nand U8135 (N_8135,N_2039,N_2859);
and U8136 (N_8136,N_4074,N_2628);
xnor U8137 (N_8137,N_1658,N_3457);
and U8138 (N_8138,N_3956,N_1045);
nand U8139 (N_8139,N_1804,N_1822);
or U8140 (N_8140,N_719,N_469);
nor U8141 (N_8141,N_1222,N_2459);
xnor U8142 (N_8142,N_567,N_2949);
nor U8143 (N_8143,N_3948,N_2151);
and U8144 (N_8144,N_4992,N_3819);
nor U8145 (N_8145,N_3118,N_4801);
or U8146 (N_8146,N_3275,N_4782);
nor U8147 (N_8147,N_3958,N_2891);
or U8148 (N_8148,N_1295,N_1629);
and U8149 (N_8149,N_1394,N_4920);
and U8150 (N_8150,N_4970,N_3842);
or U8151 (N_8151,N_2171,N_4222);
or U8152 (N_8152,N_4638,N_4402);
xnor U8153 (N_8153,N_2121,N_120);
xnor U8154 (N_8154,N_4818,N_3485);
and U8155 (N_8155,N_2408,N_639);
or U8156 (N_8156,N_546,N_1102);
nor U8157 (N_8157,N_811,N_1434);
and U8158 (N_8158,N_126,N_46);
nand U8159 (N_8159,N_1420,N_4783);
or U8160 (N_8160,N_3367,N_3185);
or U8161 (N_8161,N_2506,N_1078);
or U8162 (N_8162,N_4477,N_4175);
nand U8163 (N_8163,N_1478,N_1694);
nor U8164 (N_8164,N_929,N_4360);
and U8165 (N_8165,N_1274,N_2919);
nor U8166 (N_8166,N_1742,N_3052);
and U8167 (N_8167,N_3919,N_4253);
and U8168 (N_8168,N_1525,N_3398);
xnor U8169 (N_8169,N_3173,N_1978);
and U8170 (N_8170,N_252,N_337);
nor U8171 (N_8171,N_1564,N_1557);
or U8172 (N_8172,N_2246,N_3568);
and U8173 (N_8173,N_21,N_782);
nor U8174 (N_8174,N_290,N_4281);
or U8175 (N_8175,N_673,N_50);
nor U8176 (N_8176,N_1904,N_3413);
nor U8177 (N_8177,N_4426,N_3224);
nand U8178 (N_8178,N_4113,N_1532);
nor U8179 (N_8179,N_3501,N_1041);
and U8180 (N_8180,N_3271,N_1120);
nor U8181 (N_8181,N_1546,N_2007);
and U8182 (N_8182,N_101,N_4999);
and U8183 (N_8183,N_2443,N_2678);
xor U8184 (N_8184,N_3449,N_333);
and U8185 (N_8185,N_3723,N_3070);
nand U8186 (N_8186,N_1656,N_4595);
or U8187 (N_8187,N_4989,N_2646);
and U8188 (N_8188,N_779,N_1760);
xor U8189 (N_8189,N_416,N_4959);
nor U8190 (N_8190,N_281,N_4959);
or U8191 (N_8191,N_1090,N_4054);
or U8192 (N_8192,N_2935,N_1);
xnor U8193 (N_8193,N_4810,N_4155);
xnor U8194 (N_8194,N_4771,N_4884);
nor U8195 (N_8195,N_4311,N_1096);
nor U8196 (N_8196,N_1891,N_4715);
xnor U8197 (N_8197,N_3221,N_1120);
and U8198 (N_8198,N_773,N_4840);
nand U8199 (N_8199,N_4538,N_2956);
and U8200 (N_8200,N_1657,N_1422);
xor U8201 (N_8201,N_1950,N_4251);
nand U8202 (N_8202,N_1273,N_1874);
nand U8203 (N_8203,N_2132,N_2996);
nand U8204 (N_8204,N_818,N_2356);
xnor U8205 (N_8205,N_1906,N_3377);
nand U8206 (N_8206,N_1042,N_3799);
nand U8207 (N_8207,N_3773,N_3956);
xnor U8208 (N_8208,N_2053,N_1332);
or U8209 (N_8209,N_1048,N_2183);
nand U8210 (N_8210,N_1715,N_1331);
nand U8211 (N_8211,N_2921,N_560);
nand U8212 (N_8212,N_3380,N_1307);
xor U8213 (N_8213,N_3118,N_3490);
xnor U8214 (N_8214,N_2647,N_3310);
or U8215 (N_8215,N_4416,N_1372);
nand U8216 (N_8216,N_3886,N_4455);
nand U8217 (N_8217,N_4876,N_3788);
xor U8218 (N_8218,N_4186,N_2018);
nor U8219 (N_8219,N_4580,N_3000);
and U8220 (N_8220,N_2429,N_356);
or U8221 (N_8221,N_1655,N_2284);
xnor U8222 (N_8222,N_93,N_2012);
and U8223 (N_8223,N_4938,N_4992);
nand U8224 (N_8224,N_2488,N_419);
and U8225 (N_8225,N_1716,N_189);
or U8226 (N_8226,N_3206,N_1204);
nand U8227 (N_8227,N_425,N_3617);
and U8228 (N_8228,N_731,N_3092);
nand U8229 (N_8229,N_2612,N_1772);
nor U8230 (N_8230,N_3576,N_1465);
nor U8231 (N_8231,N_4251,N_4895);
nand U8232 (N_8232,N_1309,N_4423);
xor U8233 (N_8233,N_3726,N_498);
xor U8234 (N_8234,N_3944,N_3443);
nor U8235 (N_8235,N_2364,N_3819);
nand U8236 (N_8236,N_2889,N_1901);
nand U8237 (N_8237,N_958,N_239);
and U8238 (N_8238,N_2755,N_4020);
xnor U8239 (N_8239,N_4723,N_69);
nand U8240 (N_8240,N_4280,N_4299);
nor U8241 (N_8241,N_4002,N_4587);
nand U8242 (N_8242,N_4446,N_2332);
or U8243 (N_8243,N_1367,N_3328);
and U8244 (N_8244,N_638,N_1648);
and U8245 (N_8245,N_3962,N_1862);
nor U8246 (N_8246,N_409,N_2314);
and U8247 (N_8247,N_1449,N_1989);
and U8248 (N_8248,N_3056,N_3187);
nor U8249 (N_8249,N_1265,N_957);
xnor U8250 (N_8250,N_230,N_3090);
nor U8251 (N_8251,N_2425,N_4991);
nand U8252 (N_8252,N_224,N_1889);
nand U8253 (N_8253,N_3560,N_977);
nand U8254 (N_8254,N_4363,N_153);
or U8255 (N_8255,N_3990,N_1838);
xnor U8256 (N_8256,N_4802,N_192);
nand U8257 (N_8257,N_4129,N_1549);
and U8258 (N_8258,N_1128,N_4785);
nor U8259 (N_8259,N_1862,N_553);
or U8260 (N_8260,N_4295,N_3292);
nand U8261 (N_8261,N_4998,N_811);
or U8262 (N_8262,N_4401,N_3819);
and U8263 (N_8263,N_877,N_3454);
nor U8264 (N_8264,N_4985,N_2486);
nand U8265 (N_8265,N_3304,N_4100);
and U8266 (N_8266,N_3056,N_1632);
nor U8267 (N_8267,N_1704,N_3733);
and U8268 (N_8268,N_1020,N_1538);
xnor U8269 (N_8269,N_0,N_1751);
nand U8270 (N_8270,N_986,N_3294);
xnor U8271 (N_8271,N_158,N_1881);
and U8272 (N_8272,N_4644,N_1513);
nand U8273 (N_8273,N_395,N_3193);
and U8274 (N_8274,N_1032,N_920);
and U8275 (N_8275,N_1156,N_3037);
and U8276 (N_8276,N_387,N_473);
nor U8277 (N_8277,N_2224,N_3346);
or U8278 (N_8278,N_969,N_3170);
nand U8279 (N_8279,N_554,N_621);
and U8280 (N_8280,N_1856,N_4903);
xnor U8281 (N_8281,N_3062,N_2087);
nand U8282 (N_8282,N_233,N_3100);
or U8283 (N_8283,N_3645,N_4537);
and U8284 (N_8284,N_2211,N_337);
xor U8285 (N_8285,N_3229,N_3452);
or U8286 (N_8286,N_4142,N_567);
and U8287 (N_8287,N_124,N_1085);
xor U8288 (N_8288,N_636,N_726);
and U8289 (N_8289,N_3473,N_212);
and U8290 (N_8290,N_156,N_256);
xnor U8291 (N_8291,N_3306,N_4458);
nand U8292 (N_8292,N_430,N_3631);
nand U8293 (N_8293,N_571,N_4488);
nand U8294 (N_8294,N_1186,N_1711);
xor U8295 (N_8295,N_519,N_195);
nor U8296 (N_8296,N_1615,N_522);
xnor U8297 (N_8297,N_1514,N_1065);
xor U8298 (N_8298,N_3387,N_1982);
xnor U8299 (N_8299,N_1319,N_2565);
and U8300 (N_8300,N_367,N_4721);
nor U8301 (N_8301,N_2873,N_2590);
or U8302 (N_8302,N_410,N_34);
nand U8303 (N_8303,N_4558,N_3932);
nand U8304 (N_8304,N_4603,N_394);
nand U8305 (N_8305,N_4509,N_3138);
nor U8306 (N_8306,N_4277,N_1154);
xnor U8307 (N_8307,N_2194,N_3922);
xor U8308 (N_8308,N_1439,N_729);
nor U8309 (N_8309,N_4906,N_964);
and U8310 (N_8310,N_1973,N_1204);
and U8311 (N_8311,N_4507,N_3362);
and U8312 (N_8312,N_3023,N_3863);
or U8313 (N_8313,N_1573,N_3685);
xnor U8314 (N_8314,N_1531,N_896);
and U8315 (N_8315,N_4921,N_2032);
nor U8316 (N_8316,N_4963,N_4309);
or U8317 (N_8317,N_873,N_3141);
and U8318 (N_8318,N_94,N_4452);
nor U8319 (N_8319,N_2338,N_4398);
nor U8320 (N_8320,N_3319,N_3038);
nor U8321 (N_8321,N_2988,N_2425);
and U8322 (N_8322,N_3007,N_3043);
nand U8323 (N_8323,N_4228,N_3943);
nor U8324 (N_8324,N_2399,N_1367);
xnor U8325 (N_8325,N_1371,N_4432);
and U8326 (N_8326,N_3386,N_273);
nand U8327 (N_8327,N_1167,N_3758);
nand U8328 (N_8328,N_197,N_4677);
xnor U8329 (N_8329,N_4911,N_4299);
nor U8330 (N_8330,N_2927,N_4825);
and U8331 (N_8331,N_2240,N_2463);
nand U8332 (N_8332,N_4627,N_444);
and U8333 (N_8333,N_4272,N_111);
or U8334 (N_8334,N_4260,N_4167);
and U8335 (N_8335,N_746,N_675);
nor U8336 (N_8336,N_496,N_2010);
nor U8337 (N_8337,N_2321,N_1983);
nand U8338 (N_8338,N_990,N_4373);
or U8339 (N_8339,N_2269,N_1832);
nor U8340 (N_8340,N_2668,N_2990);
or U8341 (N_8341,N_448,N_2269);
and U8342 (N_8342,N_2277,N_2082);
nor U8343 (N_8343,N_2795,N_4221);
nand U8344 (N_8344,N_585,N_2508);
xor U8345 (N_8345,N_1868,N_839);
nand U8346 (N_8346,N_2388,N_989);
xnor U8347 (N_8347,N_4854,N_2458);
xnor U8348 (N_8348,N_4893,N_298);
xnor U8349 (N_8349,N_3318,N_587);
nand U8350 (N_8350,N_3380,N_833);
nor U8351 (N_8351,N_3537,N_1818);
xnor U8352 (N_8352,N_607,N_3551);
xnor U8353 (N_8353,N_4772,N_4689);
and U8354 (N_8354,N_3204,N_1038);
nor U8355 (N_8355,N_3055,N_1918);
nand U8356 (N_8356,N_3897,N_30);
and U8357 (N_8357,N_4933,N_1612);
nand U8358 (N_8358,N_3736,N_3817);
xnor U8359 (N_8359,N_766,N_1554);
xor U8360 (N_8360,N_721,N_2050);
or U8361 (N_8361,N_604,N_2173);
nand U8362 (N_8362,N_1635,N_2471);
or U8363 (N_8363,N_2531,N_1479);
nand U8364 (N_8364,N_2892,N_1997);
or U8365 (N_8365,N_2286,N_4506);
nand U8366 (N_8366,N_1971,N_4944);
and U8367 (N_8367,N_4591,N_3350);
or U8368 (N_8368,N_1288,N_3548);
and U8369 (N_8369,N_235,N_1581);
or U8370 (N_8370,N_4904,N_3991);
nor U8371 (N_8371,N_1527,N_889);
and U8372 (N_8372,N_4515,N_1437);
nand U8373 (N_8373,N_3055,N_3753);
and U8374 (N_8374,N_3687,N_3462);
nor U8375 (N_8375,N_116,N_3554);
nand U8376 (N_8376,N_4597,N_3367);
nor U8377 (N_8377,N_2319,N_134);
nand U8378 (N_8378,N_2139,N_305);
nand U8379 (N_8379,N_1107,N_4100);
nor U8380 (N_8380,N_469,N_2111);
xnor U8381 (N_8381,N_3095,N_3613);
nor U8382 (N_8382,N_2995,N_3298);
xnor U8383 (N_8383,N_2921,N_3743);
xor U8384 (N_8384,N_3070,N_4093);
nand U8385 (N_8385,N_3022,N_1482);
nor U8386 (N_8386,N_3486,N_1961);
nor U8387 (N_8387,N_3708,N_1935);
nor U8388 (N_8388,N_2975,N_2490);
or U8389 (N_8389,N_3256,N_4047);
nand U8390 (N_8390,N_80,N_1129);
nor U8391 (N_8391,N_4252,N_897);
nand U8392 (N_8392,N_3282,N_502);
and U8393 (N_8393,N_710,N_186);
xnor U8394 (N_8394,N_678,N_3315);
or U8395 (N_8395,N_4382,N_1580);
nand U8396 (N_8396,N_526,N_3838);
nor U8397 (N_8397,N_2900,N_769);
nand U8398 (N_8398,N_1076,N_2623);
or U8399 (N_8399,N_2175,N_1568);
xor U8400 (N_8400,N_4654,N_433);
and U8401 (N_8401,N_3988,N_2237);
nand U8402 (N_8402,N_736,N_3556);
nor U8403 (N_8403,N_2163,N_4819);
nand U8404 (N_8404,N_1206,N_4237);
nor U8405 (N_8405,N_3385,N_2955);
nand U8406 (N_8406,N_4199,N_2564);
and U8407 (N_8407,N_2838,N_471);
nand U8408 (N_8408,N_2557,N_4543);
nand U8409 (N_8409,N_3028,N_2376);
or U8410 (N_8410,N_2884,N_3547);
or U8411 (N_8411,N_3318,N_1937);
xor U8412 (N_8412,N_3620,N_1790);
nor U8413 (N_8413,N_3254,N_3101);
and U8414 (N_8414,N_3614,N_1414);
nand U8415 (N_8415,N_152,N_2910);
and U8416 (N_8416,N_543,N_4819);
or U8417 (N_8417,N_1228,N_474);
xor U8418 (N_8418,N_3033,N_931);
or U8419 (N_8419,N_1773,N_3726);
nand U8420 (N_8420,N_1267,N_74);
and U8421 (N_8421,N_3746,N_581);
nand U8422 (N_8422,N_343,N_2885);
xnor U8423 (N_8423,N_334,N_4793);
or U8424 (N_8424,N_1760,N_3514);
or U8425 (N_8425,N_470,N_572);
or U8426 (N_8426,N_3177,N_4894);
xor U8427 (N_8427,N_1116,N_1678);
or U8428 (N_8428,N_2424,N_1499);
or U8429 (N_8429,N_3396,N_1194);
or U8430 (N_8430,N_2773,N_3475);
nand U8431 (N_8431,N_3611,N_3964);
nor U8432 (N_8432,N_2170,N_740);
xor U8433 (N_8433,N_4131,N_3472);
and U8434 (N_8434,N_1151,N_4841);
or U8435 (N_8435,N_111,N_1795);
or U8436 (N_8436,N_3262,N_3746);
or U8437 (N_8437,N_2301,N_4777);
xnor U8438 (N_8438,N_3722,N_1221);
and U8439 (N_8439,N_3120,N_4595);
or U8440 (N_8440,N_1873,N_2959);
nor U8441 (N_8441,N_3367,N_2377);
or U8442 (N_8442,N_920,N_4661);
and U8443 (N_8443,N_2465,N_4054);
nor U8444 (N_8444,N_3204,N_19);
and U8445 (N_8445,N_2983,N_4014);
or U8446 (N_8446,N_4969,N_1520);
xor U8447 (N_8447,N_4307,N_3990);
and U8448 (N_8448,N_1277,N_1923);
nor U8449 (N_8449,N_1110,N_1556);
xor U8450 (N_8450,N_3329,N_4060);
nand U8451 (N_8451,N_4352,N_1916);
nand U8452 (N_8452,N_4079,N_1510);
nor U8453 (N_8453,N_2459,N_1991);
xnor U8454 (N_8454,N_3064,N_930);
nor U8455 (N_8455,N_4967,N_4787);
nand U8456 (N_8456,N_3990,N_2510);
nor U8457 (N_8457,N_337,N_3121);
nor U8458 (N_8458,N_4590,N_4691);
or U8459 (N_8459,N_2915,N_4117);
nand U8460 (N_8460,N_660,N_666);
xor U8461 (N_8461,N_535,N_4684);
nor U8462 (N_8462,N_373,N_1865);
or U8463 (N_8463,N_119,N_3420);
and U8464 (N_8464,N_1852,N_4226);
or U8465 (N_8465,N_4366,N_3000);
or U8466 (N_8466,N_3233,N_4994);
nand U8467 (N_8467,N_4751,N_53);
xor U8468 (N_8468,N_1203,N_189);
or U8469 (N_8469,N_2912,N_1554);
nor U8470 (N_8470,N_1395,N_4072);
xnor U8471 (N_8471,N_1177,N_3125);
xor U8472 (N_8472,N_3772,N_789);
nand U8473 (N_8473,N_3921,N_2754);
or U8474 (N_8474,N_4839,N_761);
xor U8475 (N_8475,N_4317,N_3781);
and U8476 (N_8476,N_3604,N_2549);
nor U8477 (N_8477,N_670,N_2950);
and U8478 (N_8478,N_2087,N_3593);
nor U8479 (N_8479,N_353,N_1917);
or U8480 (N_8480,N_1159,N_1336);
xnor U8481 (N_8481,N_2200,N_1007);
and U8482 (N_8482,N_3455,N_4733);
or U8483 (N_8483,N_1638,N_435);
xnor U8484 (N_8484,N_3315,N_1701);
and U8485 (N_8485,N_3959,N_3373);
nand U8486 (N_8486,N_1862,N_4947);
nand U8487 (N_8487,N_792,N_1284);
nand U8488 (N_8488,N_3055,N_2672);
nand U8489 (N_8489,N_1592,N_1135);
xor U8490 (N_8490,N_2144,N_1315);
nor U8491 (N_8491,N_81,N_2904);
nand U8492 (N_8492,N_297,N_4998);
xor U8493 (N_8493,N_2118,N_4006);
or U8494 (N_8494,N_3819,N_330);
xnor U8495 (N_8495,N_1192,N_4537);
and U8496 (N_8496,N_4004,N_3489);
and U8497 (N_8497,N_4152,N_194);
or U8498 (N_8498,N_3080,N_148);
nand U8499 (N_8499,N_2550,N_3038);
xnor U8500 (N_8500,N_4747,N_2046);
nor U8501 (N_8501,N_1830,N_369);
nand U8502 (N_8502,N_2094,N_1889);
and U8503 (N_8503,N_3121,N_871);
nand U8504 (N_8504,N_4331,N_1032);
or U8505 (N_8505,N_575,N_3835);
nor U8506 (N_8506,N_4486,N_3664);
nor U8507 (N_8507,N_1870,N_827);
or U8508 (N_8508,N_721,N_3144);
xor U8509 (N_8509,N_4224,N_4614);
nand U8510 (N_8510,N_3832,N_2977);
nor U8511 (N_8511,N_4555,N_303);
xor U8512 (N_8512,N_2458,N_2411);
or U8513 (N_8513,N_1403,N_3781);
nor U8514 (N_8514,N_3098,N_6);
and U8515 (N_8515,N_1919,N_2297);
nor U8516 (N_8516,N_1577,N_2305);
xor U8517 (N_8517,N_1007,N_4980);
nor U8518 (N_8518,N_151,N_1384);
xor U8519 (N_8519,N_4709,N_3389);
or U8520 (N_8520,N_565,N_25);
nand U8521 (N_8521,N_139,N_2321);
or U8522 (N_8522,N_3502,N_4742);
or U8523 (N_8523,N_3489,N_986);
and U8524 (N_8524,N_265,N_4125);
or U8525 (N_8525,N_4258,N_3733);
xnor U8526 (N_8526,N_2128,N_4787);
or U8527 (N_8527,N_1718,N_840);
xor U8528 (N_8528,N_3290,N_4898);
or U8529 (N_8529,N_4380,N_2600);
nand U8530 (N_8530,N_3133,N_3053);
nor U8531 (N_8531,N_2872,N_942);
xor U8532 (N_8532,N_1602,N_973);
nand U8533 (N_8533,N_3365,N_2586);
and U8534 (N_8534,N_601,N_100);
and U8535 (N_8535,N_691,N_2046);
nand U8536 (N_8536,N_2914,N_3806);
xnor U8537 (N_8537,N_4822,N_541);
xor U8538 (N_8538,N_4679,N_698);
or U8539 (N_8539,N_1245,N_605);
nand U8540 (N_8540,N_4722,N_648);
or U8541 (N_8541,N_4717,N_149);
nand U8542 (N_8542,N_3583,N_2335);
or U8543 (N_8543,N_241,N_3618);
nor U8544 (N_8544,N_1890,N_4535);
or U8545 (N_8545,N_2327,N_4115);
and U8546 (N_8546,N_1433,N_4346);
nor U8547 (N_8547,N_2040,N_1390);
xor U8548 (N_8548,N_2950,N_84);
nand U8549 (N_8549,N_3468,N_4888);
and U8550 (N_8550,N_1421,N_4875);
nor U8551 (N_8551,N_603,N_1972);
nor U8552 (N_8552,N_2185,N_2397);
nand U8553 (N_8553,N_1992,N_4584);
nor U8554 (N_8554,N_1915,N_3581);
nand U8555 (N_8555,N_193,N_1209);
nor U8556 (N_8556,N_870,N_3241);
xnor U8557 (N_8557,N_4357,N_1239);
nand U8558 (N_8558,N_4726,N_3654);
and U8559 (N_8559,N_3152,N_745);
and U8560 (N_8560,N_1893,N_4806);
nor U8561 (N_8561,N_2830,N_1529);
or U8562 (N_8562,N_2112,N_3294);
nand U8563 (N_8563,N_4054,N_4052);
nand U8564 (N_8564,N_4318,N_4355);
and U8565 (N_8565,N_3286,N_1831);
nor U8566 (N_8566,N_420,N_687);
nor U8567 (N_8567,N_1889,N_76);
and U8568 (N_8568,N_2099,N_3484);
xnor U8569 (N_8569,N_3088,N_4757);
xor U8570 (N_8570,N_296,N_4545);
or U8571 (N_8571,N_3468,N_1763);
or U8572 (N_8572,N_1739,N_1581);
nor U8573 (N_8573,N_1770,N_4583);
and U8574 (N_8574,N_2466,N_19);
xor U8575 (N_8575,N_3187,N_3565);
and U8576 (N_8576,N_676,N_4568);
and U8577 (N_8577,N_3981,N_563);
and U8578 (N_8578,N_1896,N_1357);
nand U8579 (N_8579,N_1107,N_3867);
or U8580 (N_8580,N_4869,N_4783);
xor U8581 (N_8581,N_4027,N_2559);
and U8582 (N_8582,N_1398,N_1728);
nor U8583 (N_8583,N_3510,N_1825);
or U8584 (N_8584,N_972,N_4435);
nand U8585 (N_8585,N_2717,N_1334);
and U8586 (N_8586,N_605,N_3879);
or U8587 (N_8587,N_2508,N_1869);
or U8588 (N_8588,N_4743,N_2097);
nand U8589 (N_8589,N_3785,N_3438);
nor U8590 (N_8590,N_4427,N_4733);
nand U8591 (N_8591,N_3603,N_398);
nand U8592 (N_8592,N_1596,N_4821);
xor U8593 (N_8593,N_271,N_3004);
xor U8594 (N_8594,N_817,N_2444);
and U8595 (N_8595,N_3986,N_2666);
and U8596 (N_8596,N_2884,N_4855);
nor U8597 (N_8597,N_594,N_3681);
and U8598 (N_8598,N_56,N_10);
or U8599 (N_8599,N_2018,N_2987);
xnor U8600 (N_8600,N_779,N_38);
or U8601 (N_8601,N_1959,N_2068);
nor U8602 (N_8602,N_2610,N_2944);
and U8603 (N_8603,N_3671,N_4518);
xnor U8604 (N_8604,N_664,N_4327);
nor U8605 (N_8605,N_3395,N_1527);
xnor U8606 (N_8606,N_527,N_533);
xnor U8607 (N_8607,N_95,N_2608);
nand U8608 (N_8608,N_3802,N_3201);
or U8609 (N_8609,N_2595,N_2360);
nor U8610 (N_8610,N_4520,N_2031);
nand U8611 (N_8611,N_1680,N_1466);
nand U8612 (N_8612,N_4503,N_1668);
nand U8613 (N_8613,N_277,N_2313);
xor U8614 (N_8614,N_375,N_4178);
or U8615 (N_8615,N_4202,N_1872);
xor U8616 (N_8616,N_4488,N_483);
and U8617 (N_8617,N_3255,N_196);
xnor U8618 (N_8618,N_2372,N_3141);
and U8619 (N_8619,N_4888,N_3381);
nand U8620 (N_8620,N_803,N_4752);
xnor U8621 (N_8621,N_387,N_2157);
nand U8622 (N_8622,N_4055,N_3946);
nand U8623 (N_8623,N_892,N_2044);
xor U8624 (N_8624,N_1808,N_2670);
or U8625 (N_8625,N_2305,N_4389);
and U8626 (N_8626,N_2971,N_498);
nand U8627 (N_8627,N_842,N_1044);
nand U8628 (N_8628,N_4816,N_218);
xnor U8629 (N_8629,N_2900,N_1334);
and U8630 (N_8630,N_4888,N_711);
nor U8631 (N_8631,N_2680,N_3943);
or U8632 (N_8632,N_4027,N_2115);
nor U8633 (N_8633,N_27,N_4156);
nor U8634 (N_8634,N_1404,N_2123);
xnor U8635 (N_8635,N_316,N_4631);
nand U8636 (N_8636,N_3909,N_1860);
and U8637 (N_8637,N_1462,N_778);
or U8638 (N_8638,N_1446,N_3712);
nand U8639 (N_8639,N_84,N_3383);
and U8640 (N_8640,N_1168,N_1355);
or U8641 (N_8641,N_1133,N_4140);
nor U8642 (N_8642,N_261,N_2011);
or U8643 (N_8643,N_4656,N_4688);
and U8644 (N_8644,N_861,N_3236);
nor U8645 (N_8645,N_4240,N_3237);
or U8646 (N_8646,N_1247,N_1591);
or U8647 (N_8647,N_2880,N_1081);
nor U8648 (N_8648,N_384,N_1017);
nor U8649 (N_8649,N_3834,N_3639);
or U8650 (N_8650,N_1584,N_2670);
nand U8651 (N_8651,N_4315,N_3364);
nor U8652 (N_8652,N_4072,N_1717);
nand U8653 (N_8653,N_807,N_4677);
nand U8654 (N_8654,N_2302,N_1186);
or U8655 (N_8655,N_3959,N_4483);
and U8656 (N_8656,N_4708,N_439);
nand U8657 (N_8657,N_4134,N_3086);
nor U8658 (N_8658,N_4388,N_815);
xor U8659 (N_8659,N_1368,N_2941);
or U8660 (N_8660,N_1949,N_1635);
nand U8661 (N_8661,N_4763,N_1862);
or U8662 (N_8662,N_4000,N_1464);
and U8663 (N_8663,N_775,N_159);
and U8664 (N_8664,N_3003,N_2827);
nand U8665 (N_8665,N_2696,N_4870);
nand U8666 (N_8666,N_599,N_1103);
or U8667 (N_8667,N_4668,N_2528);
or U8668 (N_8668,N_4995,N_4500);
xnor U8669 (N_8669,N_1678,N_2042);
or U8670 (N_8670,N_4646,N_377);
nand U8671 (N_8671,N_235,N_2403);
nor U8672 (N_8672,N_4919,N_3749);
nand U8673 (N_8673,N_148,N_828);
or U8674 (N_8674,N_1888,N_4875);
xor U8675 (N_8675,N_2315,N_3051);
nand U8676 (N_8676,N_216,N_4610);
nand U8677 (N_8677,N_528,N_3604);
nor U8678 (N_8678,N_4889,N_4017);
or U8679 (N_8679,N_1134,N_1360);
xnor U8680 (N_8680,N_4374,N_1908);
xnor U8681 (N_8681,N_7,N_948);
and U8682 (N_8682,N_672,N_3364);
or U8683 (N_8683,N_1527,N_3912);
xnor U8684 (N_8684,N_4180,N_3623);
nand U8685 (N_8685,N_1613,N_4699);
or U8686 (N_8686,N_2520,N_2163);
nor U8687 (N_8687,N_2380,N_524);
nor U8688 (N_8688,N_2773,N_2636);
and U8689 (N_8689,N_4485,N_17);
nor U8690 (N_8690,N_2044,N_1924);
xor U8691 (N_8691,N_4114,N_848);
and U8692 (N_8692,N_2882,N_4144);
xor U8693 (N_8693,N_3904,N_713);
and U8694 (N_8694,N_77,N_3495);
or U8695 (N_8695,N_2899,N_1644);
xnor U8696 (N_8696,N_2138,N_4944);
and U8697 (N_8697,N_4761,N_3304);
or U8698 (N_8698,N_645,N_280);
xor U8699 (N_8699,N_292,N_142);
and U8700 (N_8700,N_4193,N_4371);
nand U8701 (N_8701,N_325,N_3604);
xor U8702 (N_8702,N_4624,N_1789);
xnor U8703 (N_8703,N_4745,N_2472);
xor U8704 (N_8704,N_2722,N_3214);
nand U8705 (N_8705,N_168,N_82);
xor U8706 (N_8706,N_2081,N_69);
or U8707 (N_8707,N_3651,N_3230);
and U8708 (N_8708,N_383,N_2868);
and U8709 (N_8709,N_2322,N_3145);
xor U8710 (N_8710,N_447,N_769);
and U8711 (N_8711,N_455,N_4123);
and U8712 (N_8712,N_2188,N_1209);
and U8713 (N_8713,N_1421,N_1264);
and U8714 (N_8714,N_4972,N_175);
xnor U8715 (N_8715,N_1296,N_4009);
or U8716 (N_8716,N_230,N_537);
and U8717 (N_8717,N_894,N_4483);
and U8718 (N_8718,N_3934,N_4510);
xnor U8719 (N_8719,N_4907,N_2739);
nor U8720 (N_8720,N_4703,N_4146);
xnor U8721 (N_8721,N_348,N_2987);
nand U8722 (N_8722,N_2087,N_67);
and U8723 (N_8723,N_2531,N_1584);
or U8724 (N_8724,N_4021,N_670);
or U8725 (N_8725,N_2295,N_491);
xnor U8726 (N_8726,N_3655,N_2610);
xor U8727 (N_8727,N_1359,N_2226);
and U8728 (N_8728,N_1198,N_4171);
xor U8729 (N_8729,N_3583,N_1098);
or U8730 (N_8730,N_3225,N_3165);
nor U8731 (N_8731,N_563,N_2580);
or U8732 (N_8732,N_855,N_4052);
and U8733 (N_8733,N_1094,N_1853);
xor U8734 (N_8734,N_902,N_501);
nand U8735 (N_8735,N_4217,N_1720);
nor U8736 (N_8736,N_4621,N_3497);
xor U8737 (N_8737,N_3293,N_2790);
or U8738 (N_8738,N_3984,N_1973);
nor U8739 (N_8739,N_2934,N_4330);
nand U8740 (N_8740,N_3825,N_2884);
nand U8741 (N_8741,N_3828,N_2473);
nor U8742 (N_8742,N_2094,N_4535);
nand U8743 (N_8743,N_2413,N_3028);
or U8744 (N_8744,N_4174,N_2597);
nor U8745 (N_8745,N_2844,N_4995);
nand U8746 (N_8746,N_1873,N_3260);
nand U8747 (N_8747,N_577,N_1170);
xor U8748 (N_8748,N_1511,N_4438);
xnor U8749 (N_8749,N_814,N_834);
nand U8750 (N_8750,N_2377,N_1645);
and U8751 (N_8751,N_4141,N_2238);
and U8752 (N_8752,N_2307,N_4390);
nand U8753 (N_8753,N_4649,N_4265);
and U8754 (N_8754,N_4348,N_1951);
or U8755 (N_8755,N_3910,N_2990);
nor U8756 (N_8756,N_283,N_579);
or U8757 (N_8757,N_737,N_3640);
nand U8758 (N_8758,N_58,N_2942);
or U8759 (N_8759,N_1832,N_884);
xnor U8760 (N_8760,N_1107,N_2980);
nor U8761 (N_8761,N_521,N_22);
nor U8762 (N_8762,N_4737,N_4124);
xor U8763 (N_8763,N_4922,N_2071);
nand U8764 (N_8764,N_4381,N_4265);
nand U8765 (N_8765,N_2032,N_160);
nand U8766 (N_8766,N_4063,N_4627);
or U8767 (N_8767,N_374,N_3835);
or U8768 (N_8768,N_1372,N_762);
xnor U8769 (N_8769,N_352,N_2605);
nand U8770 (N_8770,N_1441,N_2493);
nand U8771 (N_8771,N_3928,N_993);
nor U8772 (N_8772,N_2251,N_487);
nand U8773 (N_8773,N_3371,N_207);
nand U8774 (N_8774,N_1724,N_3477);
nand U8775 (N_8775,N_3408,N_3449);
and U8776 (N_8776,N_2938,N_3485);
or U8777 (N_8777,N_2519,N_4383);
nor U8778 (N_8778,N_1071,N_1480);
and U8779 (N_8779,N_4592,N_4035);
or U8780 (N_8780,N_63,N_2216);
or U8781 (N_8781,N_3316,N_3570);
and U8782 (N_8782,N_410,N_1548);
and U8783 (N_8783,N_4336,N_3653);
and U8784 (N_8784,N_597,N_4042);
and U8785 (N_8785,N_295,N_90);
nor U8786 (N_8786,N_1979,N_4494);
and U8787 (N_8787,N_4009,N_4713);
nand U8788 (N_8788,N_3531,N_1300);
and U8789 (N_8789,N_2125,N_111);
xor U8790 (N_8790,N_339,N_113);
and U8791 (N_8791,N_4148,N_4753);
nor U8792 (N_8792,N_2745,N_1051);
and U8793 (N_8793,N_3701,N_4484);
xnor U8794 (N_8794,N_602,N_2376);
nand U8795 (N_8795,N_1999,N_2191);
xor U8796 (N_8796,N_3992,N_442);
and U8797 (N_8797,N_4523,N_4940);
or U8798 (N_8798,N_1663,N_1820);
nand U8799 (N_8799,N_3805,N_435);
nor U8800 (N_8800,N_4915,N_4191);
or U8801 (N_8801,N_4135,N_203);
nor U8802 (N_8802,N_2147,N_183);
xor U8803 (N_8803,N_1467,N_4755);
nor U8804 (N_8804,N_821,N_144);
nor U8805 (N_8805,N_1268,N_2633);
xor U8806 (N_8806,N_3397,N_1740);
xnor U8807 (N_8807,N_1467,N_2274);
and U8808 (N_8808,N_3363,N_1683);
nand U8809 (N_8809,N_4723,N_3465);
or U8810 (N_8810,N_4287,N_3341);
nand U8811 (N_8811,N_274,N_455);
and U8812 (N_8812,N_1630,N_4199);
or U8813 (N_8813,N_2651,N_1522);
xor U8814 (N_8814,N_678,N_2295);
nor U8815 (N_8815,N_1515,N_178);
or U8816 (N_8816,N_4208,N_3255);
nand U8817 (N_8817,N_3640,N_994);
nor U8818 (N_8818,N_4223,N_733);
nand U8819 (N_8819,N_73,N_4455);
and U8820 (N_8820,N_131,N_2861);
and U8821 (N_8821,N_3126,N_591);
xor U8822 (N_8822,N_1415,N_4890);
or U8823 (N_8823,N_2472,N_1680);
or U8824 (N_8824,N_1632,N_1574);
and U8825 (N_8825,N_4585,N_1885);
nand U8826 (N_8826,N_4571,N_3065);
or U8827 (N_8827,N_4409,N_2351);
or U8828 (N_8828,N_922,N_1259);
nor U8829 (N_8829,N_940,N_471);
xnor U8830 (N_8830,N_4061,N_4340);
and U8831 (N_8831,N_1116,N_3991);
nand U8832 (N_8832,N_3743,N_4211);
and U8833 (N_8833,N_278,N_3353);
nand U8834 (N_8834,N_979,N_4990);
nand U8835 (N_8835,N_4171,N_3758);
nor U8836 (N_8836,N_1519,N_3701);
xor U8837 (N_8837,N_1374,N_1826);
or U8838 (N_8838,N_37,N_3945);
or U8839 (N_8839,N_3618,N_1356);
nor U8840 (N_8840,N_2523,N_1050);
nor U8841 (N_8841,N_3706,N_3914);
nor U8842 (N_8842,N_399,N_4081);
xnor U8843 (N_8843,N_2744,N_212);
nand U8844 (N_8844,N_4906,N_4363);
and U8845 (N_8845,N_4841,N_385);
xnor U8846 (N_8846,N_2394,N_1904);
nor U8847 (N_8847,N_3984,N_1637);
xor U8848 (N_8848,N_2991,N_1267);
nand U8849 (N_8849,N_3244,N_1674);
nand U8850 (N_8850,N_2667,N_3382);
and U8851 (N_8851,N_4939,N_3644);
nand U8852 (N_8852,N_3635,N_733);
xor U8853 (N_8853,N_1474,N_174);
nand U8854 (N_8854,N_770,N_1980);
or U8855 (N_8855,N_3649,N_3137);
or U8856 (N_8856,N_3970,N_1624);
nor U8857 (N_8857,N_1054,N_2689);
xnor U8858 (N_8858,N_4811,N_4940);
xnor U8859 (N_8859,N_2013,N_3678);
nand U8860 (N_8860,N_3370,N_4135);
and U8861 (N_8861,N_3975,N_4604);
and U8862 (N_8862,N_2218,N_4480);
nand U8863 (N_8863,N_2363,N_673);
nand U8864 (N_8864,N_2363,N_1098);
and U8865 (N_8865,N_2140,N_2894);
xnor U8866 (N_8866,N_3274,N_4372);
nor U8867 (N_8867,N_94,N_4860);
nor U8868 (N_8868,N_1603,N_1628);
and U8869 (N_8869,N_2295,N_4932);
or U8870 (N_8870,N_706,N_4948);
or U8871 (N_8871,N_610,N_272);
and U8872 (N_8872,N_2180,N_3313);
and U8873 (N_8873,N_3391,N_3795);
nor U8874 (N_8874,N_4812,N_1099);
xnor U8875 (N_8875,N_4630,N_750);
and U8876 (N_8876,N_2462,N_1421);
or U8877 (N_8877,N_2217,N_1832);
xnor U8878 (N_8878,N_2197,N_1714);
nand U8879 (N_8879,N_3941,N_2157);
xor U8880 (N_8880,N_528,N_3952);
xnor U8881 (N_8881,N_2875,N_3734);
xnor U8882 (N_8882,N_3565,N_219);
nor U8883 (N_8883,N_4927,N_3401);
xnor U8884 (N_8884,N_1841,N_4893);
nand U8885 (N_8885,N_1875,N_410);
nand U8886 (N_8886,N_2469,N_1707);
nor U8887 (N_8887,N_775,N_3081);
or U8888 (N_8888,N_2697,N_4479);
nor U8889 (N_8889,N_4324,N_3242);
nor U8890 (N_8890,N_2898,N_2913);
nand U8891 (N_8891,N_3086,N_3927);
nand U8892 (N_8892,N_368,N_3902);
and U8893 (N_8893,N_2811,N_4550);
and U8894 (N_8894,N_1741,N_4231);
xnor U8895 (N_8895,N_4220,N_2563);
nor U8896 (N_8896,N_3347,N_13);
or U8897 (N_8897,N_2159,N_4046);
or U8898 (N_8898,N_229,N_3867);
nor U8899 (N_8899,N_3181,N_748);
or U8900 (N_8900,N_4333,N_2945);
or U8901 (N_8901,N_4538,N_2987);
nand U8902 (N_8902,N_296,N_979);
xor U8903 (N_8903,N_2462,N_964);
or U8904 (N_8904,N_1104,N_112);
or U8905 (N_8905,N_3704,N_1066);
and U8906 (N_8906,N_1540,N_1152);
and U8907 (N_8907,N_1266,N_3492);
and U8908 (N_8908,N_3310,N_176);
xnor U8909 (N_8909,N_95,N_2355);
nor U8910 (N_8910,N_2441,N_4864);
xnor U8911 (N_8911,N_3537,N_1241);
nor U8912 (N_8912,N_4086,N_4244);
xor U8913 (N_8913,N_2229,N_4763);
xnor U8914 (N_8914,N_1966,N_469);
and U8915 (N_8915,N_669,N_3798);
and U8916 (N_8916,N_1419,N_333);
xnor U8917 (N_8917,N_74,N_2284);
nor U8918 (N_8918,N_4968,N_1960);
nor U8919 (N_8919,N_766,N_4452);
xnor U8920 (N_8920,N_3613,N_2914);
nor U8921 (N_8921,N_3917,N_1303);
nand U8922 (N_8922,N_3446,N_1183);
and U8923 (N_8923,N_2440,N_15);
xor U8924 (N_8924,N_2999,N_3790);
nand U8925 (N_8925,N_1454,N_3734);
nor U8926 (N_8926,N_795,N_4521);
and U8927 (N_8927,N_1385,N_1846);
and U8928 (N_8928,N_2966,N_4405);
and U8929 (N_8929,N_4287,N_884);
xor U8930 (N_8930,N_1480,N_1435);
nor U8931 (N_8931,N_1479,N_2640);
and U8932 (N_8932,N_574,N_4523);
nor U8933 (N_8933,N_2973,N_1415);
xor U8934 (N_8934,N_2778,N_941);
nor U8935 (N_8935,N_3764,N_2958);
or U8936 (N_8936,N_4046,N_4273);
nand U8937 (N_8937,N_3815,N_4298);
nand U8938 (N_8938,N_2073,N_2242);
and U8939 (N_8939,N_4851,N_740);
xor U8940 (N_8940,N_228,N_3851);
nor U8941 (N_8941,N_2487,N_769);
nor U8942 (N_8942,N_3360,N_971);
nand U8943 (N_8943,N_1602,N_1480);
nand U8944 (N_8944,N_2414,N_819);
xor U8945 (N_8945,N_868,N_1397);
xnor U8946 (N_8946,N_1368,N_1975);
or U8947 (N_8947,N_1546,N_660);
xnor U8948 (N_8948,N_2292,N_1580);
nand U8949 (N_8949,N_1059,N_1868);
nand U8950 (N_8950,N_173,N_1540);
nor U8951 (N_8951,N_4538,N_1656);
xor U8952 (N_8952,N_30,N_2981);
nor U8953 (N_8953,N_288,N_1606);
nand U8954 (N_8954,N_3717,N_4023);
nor U8955 (N_8955,N_349,N_1755);
and U8956 (N_8956,N_3052,N_731);
or U8957 (N_8957,N_3369,N_3324);
or U8958 (N_8958,N_1633,N_2745);
or U8959 (N_8959,N_3018,N_2525);
nor U8960 (N_8960,N_2489,N_3544);
and U8961 (N_8961,N_1561,N_2362);
nand U8962 (N_8962,N_3618,N_3217);
and U8963 (N_8963,N_2074,N_1427);
and U8964 (N_8964,N_2366,N_23);
nor U8965 (N_8965,N_982,N_3135);
and U8966 (N_8966,N_4859,N_4386);
xor U8967 (N_8967,N_2423,N_4470);
xnor U8968 (N_8968,N_3761,N_511);
nand U8969 (N_8969,N_3939,N_4249);
or U8970 (N_8970,N_2978,N_2961);
or U8971 (N_8971,N_2031,N_3902);
nand U8972 (N_8972,N_3882,N_903);
nor U8973 (N_8973,N_1104,N_82);
nor U8974 (N_8974,N_2471,N_569);
nor U8975 (N_8975,N_3422,N_4760);
xor U8976 (N_8976,N_18,N_4632);
xor U8977 (N_8977,N_151,N_2063);
and U8978 (N_8978,N_1076,N_2448);
nor U8979 (N_8979,N_945,N_2592);
nor U8980 (N_8980,N_3108,N_4664);
or U8981 (N_8981,N_4209,N_908);
nor U8982 (N_8982,N_68,N_2598);
and U8983 (N_8983,N_4780,N_2460);
nor U8984 (N_8984,N_3332,N_2350);
nor U8985 (N_8985,N_3646,N_4256);
nand U8986 (N_8986,N_4086,N_835);
nor U8987 (N_8987,N_2479,N_4293);
xnor U8988 (N_8988,N_3954,N_4466);
xor U8989 (N_8989,N_2997,N_2710);
and U8990 (N_8990,N_2109,N_4887);
or U8991 (N_8991,N_1085,N_1834);
nand U8992 (N_8992,N_2272,N_4382);
nand U8993 (N_8993,N_2441,N_2870);
nor U8994 (N_8994,N_4507,N_4733);
xor U8995 (N_8995,N_3177,N_1018);
nand U8996 (N_8996,N_1742,N_3151);
xor U8997 (N_8997,N_3124,N_1180);
nor U8998 (N_8998,N_2173,N_1740);
nor U8999 (N_8999,N_4335,N_3520);
nand U9000 (N_9000,N_4514,N_3467);
nand U9001 (N_9001,N_513,N_3504);
and U9002 (N_9002,N_671,N_1513);
or U9003 (N_9003,N_4426,N_2014);
nand U9004 (N_9004,N_217,N_3757);
xor U9005 (N_9005,N_3398,N_2129);
or U9006 (N_9006,N_4069,N_1425);
or U9007 (N_9007,N_1671,N_1292);
and U9008 (N_9008,N_587,N_346);
or U9009 (N_9009,N_3066,N_3185);
nor U9010 (N_9010,N_4334,N_4712);
or U9011 (N_9011,N_3482,N_2670);
nor U9012 (N_9012,N_4494,N_4090);
nand U9013 (N_9013,N_1543,N_4865);
or U9014 (N_9014,N_3443,N_1389);
nor U9015 (N_9015,N_4297,N_1889);
xnor U9016 (N_9016,N_3319,N_729);
nand U9017 (N_9017,N_1006,N_3691);
nand U9018 (N_9018,N_4178,N_1845);
or U9019 (N_9019,N_1886,N_3094);
and U9020 (N_9020,N_2788,N_4437);
xor U9021 (N_9021,N_2705,N_3119);
nor U9022 (N_9022,N_3696,N_1790);
nand U9023 (N_9023,N_3439,N_1905);
nor U9024 (N_9024,N_4715,N_4733);
nor U9025 (N_9025,N_4488,N_1756);
and U9026 (N_9026,N_128,N_2440);
nor U9027 (N_9027,N_4168,N_3871);
nand U9028 (N_9028,N_3841,N_4608);
nand U9029 (N_9029,N_4841,N_2962);
nor U9030 (N_9030,N_2846,N_2177);
nor U9031 (N_9031,N_4120,N_2071);
xnor U9032 (N_9032,N_4507,N_4522);
xor U9033 (N_9033,N_4102,N_4062);
or U9034 (N_9034,N_4520,N_4109);
and U9035 (N_9035,N_4865,N_2450);
nand U9036 (N_9036,N_1924,N_3876);
nor U9037 (N_9037,N_1392,N_3885);
or U9038 (N_9038,N_1341,N_1998);
xor U9039 (N_9039,N_2634,N_1674);
or U9040 (N_9040,N_3672,N_2762);
or U9041 (N_9041,N_2603,N_4852);
nor U9042 (N_9042,N_228,N_1944);
or U9043 (N_9043,N_3001,N_1776);
xor U9044 (N_9044,N_2984,N_3009);
nor U9045 (N_9045,N_1247,N_3824);
and U9046 (N_9046,N_2201,N_2884);
nand U9047 (N_9047,N_4030,N_3631);
and U9048 (N_9048,N_2977,N_1411);
nor U9049 (N_9049,N_2839,N_1270);
and U9050 (N_9050,N_3260,N_3592);
and U9051 (N_9051,N_2205,N_382);
nand U9052 (N_9052,N_1574,N_3829);
and U9053 (N_9053,N_4897,N_1590);
or U9054 (N_9054,N_1218,N_1459);
nand U9055 (N_9055,N_3492,N_1966);
nor U9056 (N_9056,N_3538,N_1928);
nand U9057 (N_9057,N_2507,N_1674);
nor U9058 (N_9058,N_1674,N_4605);
nand U9059 (N_9059,N_857,N_1837);
or U9060 (N_9060,N_7,N_2368);
xor U9061 (N_9061,N_2004,N_4106);
xnor U9062 (N_9062,N_2458,N_1253);
nand U9063 (N_9063,N_1413,N_4419);
and U9064 (N_9064,N_2623,N_1528);
xor U9065 (N_9065,N_1754,N_3380);
nor U9066 (N_9066,N_1450,N_1395);
nor U9067 (N_9067,N_3607,N_1332);
xnor U9068 (N_9068,N_3537,N_1036);
and U9069 (N_9069,N_4730,N_3406);
or U9070 (N_9070,N_1739,N_2452);
xor U9071 (N_9071,N_3009,N_4559);
nor U9072 (N_9072,N_3012,N_4608);
and U9073 (N_9073,N_665,N_1891);
nand U9074 (N_9074,N_2709,N_136);
and U9075 (N_9075,N_1232,N_3228);
nor U9076 (N_9076,N_1785,N_4616);
or U9077 (N_9077,N_421,N_1235);
xor U9078 (N_9078,N_1637,N_1773);
nand U9079 (N_9079,N_1814,N_2641);
and U9080 (N_9080,N_1283,N_4448);
nand U9081 (N_9081,N_4489,N_456);
nor U9082 (N_9082,N_1988,N_1056);
nand U9083 (N_9083,N_4567,N_151);
or U9084 (N_9084,N_1028,N_4211);
xnor U9085 (N_9085,N_574,N_3551);
or U9086 (N_9086,N_1223,N_228);
and U9087 (N_9087,N_1838,N_4718);
and U9088 (N_9088,N_2861,N_601);
nand U9089 (N_9089,N_3763,N_1037);
nand U9090 (N_9090,N_4864,N_962);
nor U9091 (N_9091,N_2980,N_3562);
xnor U9092 (N_9092,N_3352,N_922);
and U9093 (N_9093,N_3414,N_3642);
xor U9094 (N_9094,N_2233,N_2130);
nor U9095 (N_9095,N_1134,N_2543);
xnor U9096 (N_9096,N_1314,N_1785);
nor U9097 (N_9097,N_1442,N_2633);
and U9098 (N_9098,N_2191,N_975);
nand U9099 (N_9099,N_3287,N_4719);
nand U9100 (N_9100,N_1536,N_4635);
nor U9101 (N_9101,N_3339,N_2486);
and U9102 (N_9102,N_2938,N_2753);
and U9103 (N_9103,N_2896,N_3663);
nand U9104 (N_9104,N_959,N_387);
and U9105 (N_9105,N_941,N_344);
nand U9106 (N_9106,N_4293,N_3831);
nand U9107 (N_9107,N_4358,N_1751);
or U9108 (N_9108,N_488,N_298);
nand U9109 (N_9109,N_3942,N_3410);
and U9110 (N_9110,N_1429,N_3992);
and U9111 (N_9111,N_2871,N_2564);
and U9112 (N_9112,N_2997,N_3634);
xor U9113 (N_9113,N_4818,N_122);
xor U9114 (N_9114,N_3055,N_2636);
and U9115 (N_9115,N_1612,N_4366);
nor U9116 (N_9116,N_1026,N_823);
and U9117 (N_9117,N_809,N_4186);
or U9118 (N_9118,N_2625,N_3434);
or U9119 (N_9119,N_615,N_2693);
and U9120 (N_9120,N_2201,N_4568);
xor U9121 (N_9121,N_3163,N_1706);
or U9122 (N_9122,N_2031,N_1349);
nand U9123 (N_9123,N_4173,N_3155);
and U9124 (N_9124,N_2590,N_3240);
or U9125 (N_9125,N_4949,N_574);
nand U9126 (N_9126,N_4510,N_3529);
and U9127 (N_9127,N_2825,N_313);
nand U9128 (N_9128,N_4304,N_4481);
xnor U9129 (N_9129,N_2084,N_2312);
xnor U9130 (N_9130,N_3058,N_2744);
and U9131 (N_9131,N_1845,N_4344);
nor U9132 (N_9132,N_3819,N_623);
or U9133 (N_9133,N_4314,N_2637);
and U9134 (N_9134,N_1998,N_2831);
and U9135 (N_9135,N_725,N_819);
and U9136 (N_9136,N_3080,N_4923);
nand U9137 (N_9137,N_3201,N_2639);
nor U9138 (N_9138,N_4621,N_2006);
nand U9139 (N_9139,N_3177,N_3154);
nand U9140 (N_9140,N_442,N_1663);
or U9141 (N_9141,N_1787,N_4964);
nor U9142 (N_9142,N_4722,N_4708);
xor U9143 (N_9143,N_3326,N_3232);
xnor U9144 (N_9144,N_2960,N_206);
xnor U9145 (N_9145,N_4490,N_3838);
or U9146 (N_9146,N_1335,N_3609);
nor U9147 (N_9147,N_1853,N_1913);
xor U9148 (N_9148,N_2157,N_1587);
nand U9149 (N_9149,N_3242,N_2943);
xnor U9150 (N_9150,N_2081,N_4970);
nand U9151 (N_9151,N_3537,N_877);
and U9152 (N_9152,N_1952,N_1661);
xor U9153 (N_9153,N_4064,N_547);
nor U9154 (N_9154,N_2744,N_1320);
or U9155 (N_9155,N_1433,N_1080);
or U9156 (N_9156,N_2344,N_1215);
xor U9157 (N_9157,N_4142,N_2980);
nand U9158 (N_9158,N_1497,N_2246);
nand U9159 (N_9159,N_3093,N_4409);
nor U9160 (N_9160,N_2311,N_4978);
nor U9161 (N_9161,N_2130,N_4893);
and U9162 (N_9162,N_32,N_2429);
xnor U9163 (N_9163,N_4069,N_2383);
or U9164 (N_9164,N_4671,N_1286);
xnor U9165 (N_9165,N_1714,N_2334);
or U9166 (N_9166,N_1472,N_249);
nor U9167 (N_9167,N_3389,N_3147);
nand U9168 (N_9168,N_2479,N_3163);
and U9169 (N_9169,N_1539,N_402);
xor U9170 (N_9170,N_2248,N_3149);
xnor U9171 (N_9171,N_2777,N_3221);
xnor U9172 (N_9172,N_1895,N_2150);
or U9173 (N_9173,N_2143,N_4463);
nor U9174 (N_9174,N_3804,N_366);
xnor U9175 (N_9175,N_3370,N_4064);
nand U9176 (N_9176,N_1841,N_2118);
xnor U9177 (N_9177,N_4390,N_4057);
or U9178 (N_9178,N_1348,N_4106);
xor U9179 (N_9179,N_2088,N_1558);
and U9180 (N_9180,N_3892,N_3517);
and U9181 (N_9181,N_4845,N_590);
or U9182 (N_9182,N_1780,N_1746);
and U9183 (N_9183,N_4449,N_538);
nor U9184 (N_9184,N_3723,N_3505);
nand U9185 (N_9185,N_853,N_257);
or U9186 (N_9186,N_2380,N_4748);
nand U9187 (N_9187,N_4542,N_2841);
nand U9188 (N_9188,N_2553,N_3443);
nand U9189 (N_9189,N_590,N_3513);
xnor U9190 (N_9190,N_4059,N_3258);
xnor U9191 (N_9191,N_2812,N_2604);
nand U9192 (N_9192,N_2183,N_1037);
and U9193 (N_9193,N_3422,N_4920);
or U9194 (N_9194,N_2675,N_3509);
nand U9195 (N_9195,N_1934,N_3944);
nor U9196 (N_9196,N_22,N_3040);
and U9197 (N_9197,N_4709,N_1235);
nand U9198 (N_9198,N_808,N_609);
nand U9199 (N_9199,N_557,N_4941);
and U9200 (N_9200,N_2055,N_1282);
nor U9201 (N_9201,N_3484,N_4695);
and U9202 (N_9202,N_2279,N_65);
or U9203 (N_9203,N_3129,N_3392);
xor U9204 (N_9204,N_3683,N_2154);
nor U9205 (N_9205,N_4322,N_1099);
and U9206 (N_9206,N_1901,N_1597);
nor U9207 (N_9207,N_3784,N_534);
xor U9208 (N_9208,N_2010,N_600);
or U9209 (N_9209,N_192,N_4728);
or U9210 (N_9210,N_4676,N_2445);
and U9211 (N_9211,N_2026,N_2348);
or U9212 (N_9212,N_117,N_1908);
and U9213 (N_9213,N_2709,N_1463);
nand U9214 (N_9214,N_65,N_1531);
xnor U9215 (N_9215,N_721,N_1845);
nor U9216 (N_9216,N_674,N_286);
nand U9217 (N_9217,N_326,N_3620);
or U9218 (N_9218,N_3675,N_3914);
or U9219 (N_9219,N_3766,N_305);
or U9220 (N_9220,N_2892,N_4832);
or U9221 (N_9221,N_3317,N_2248);
nand U9222 (N_9222,N_1584,N_439);
and U9223 (N_9223,N_3549,N_1383);
nor U9224 (N_9224,N_2208,N_347);
and U9225 (N_9225,N_4489,N_4730);
or U9226 (N_9226,N_1708,N_628);
or U9227 (N_9227,N_1754,N_367);
or U9228 (N_9228,N_1450,N_4793);
xnor U9229 (N_9229,N_1967,N_1176);
nand U9230 (N_9230,N_3642,N_4861);
xnor U9231 (N_9231,N_2806,N_2311);
or U9232 (N_9232,N_4923,N_1093);
xnor U9233 (N_9233,N_4708,N_3513);
nor U9234 (N_9234,N_611,N_2290);
and U9235 (N_9235,N_2229,N_3354);
and U9236 (N_9236,N_2718,N_2105);
nand U9237 (N_9237,N_951,N_2105);
nor U9238 (N_9238,N_2023,N_2294);
or U9239 (N_9239,N_4595,N_4819);
or U9240 (N_9240,N_4594,N_182);
nand U9241 (N_9241,N_113,N_3642);
xor U9242 (N_9242,N_96,N_4514);
or U9243 (N_9243,N_4350,N_4106);
nand U9244 (N_9244,N_1612,N_4535);
and U9245 (N_9245,N_942,N_3869);
and U9246 (N_9246,N_2687,N_4300);
and U9247 (N_9247,N_809,N_1994);
or U9248 (N_9248,N_2658,N_3071);
and U9249 (N_9249,N_3915,N_3769);
nand U9250 (N_9250,N_412,N_1271);
xnor U9251 (N_9251,N_1566,N_1774);
and U9252 (N_9252,N_4691,N_3751);
nand U9253 (N_9253,N_1463,N_1891);
or U9254 (N_9254,N_214,N_537);
and U9255 (N_9255,N_1608,N_4518);
or U9256 (N_9256,N_3349,N_2349);
nor U9257 (N_9257,N_2693,N_1858);
and U9258 (N_9258,N_164,N_4140);
nand U9259 (N_9259,N_3759,N_1367);
nand U9260 (N_9260,N_4794,N_4674);
nor U9261 (N_9261,N_4195,N_553);
nor U9262 (N_9262,N_4318,N_495);
nor U9263 (N_9263,N_969,N_417);
nand U9264 (N_9264,N_2889,N_1935);
nand U9265 (N_9265,N_2449,N_4746);
or U9266 (N_9266,N_2910,N_3761);
or U9267 (N_9267,N_2717,N_615);
or U9268 (N_9268,N_1892,N_907);
and U9269 (N_9269,N_4085,N_3015);
nor U9270 (N_9270,N_4429,N_1150);
nand U9271 (N_9271,N_3755,N_2385);
xnor U9272 (N_9272,N_1487,N_1469);
nor U9273 (N_9273,N_3386,N_965);
xor U9274 (N_9274,N_4869,N_2968);
nor U9275 (N_9275,N_4736,N_1036);
xor U9276 (N_9276,N_789,N_1994);
xor U9277 (N_9277,N_2285,N_2546);
nor U9278 (N_9278,N_400,N_1150);
and U9279 (N_9279,N_965,N_3189);
nor U9280 (N_9280,N_928,N_402);
xnor U9281 (N_9281,N_2079,N_487);
xnor U9282 (N_9282,N_1622,N_2398);
or U9283 (N_9283,N_1308,N_3203);
and U9284 (N_9284,N_2677,N_2034);
nand U9285 (N_9285,N_4341,N_2723);
and U9286 (N_9286,N_1171,N_80);
or U9287 (N_9287,N_4396,N_1340);
and U9288 (N_9288,N_2245,N_3193);
and U9289 (N_9289,N_3274,N_4954);
nand U9290 (N_9290,N_3546,N_3822);
nand U9291 (N_9291,N_1578,N_1520);
nand U9292 (N_9292,N_1135,N_1546);
nand U9293 (N_9293,N_3112,N_4361);
xnor U9294 (N_9294,N_4748,N_3517);
or U9295 (N_9295,N_1463,N_2355);
or U9296 (N_9296,N_883,N_1803);
or U9297 (N_9297,N_4389,N_1468);
nand U9298 (N_9298,N_3713,N_383);
nor U9299 (N_9299,N_2301,N_4913);
nand U9300 (N_9300,N_4446,N_511);
or U9301 (N_9301,N_4853,N_4436);
or U9302 (N_9302,N_2634,N_513);
nand U9303 (N_9303,N_4473,N_2161);
nor U9304 (N_9304,N_3749,N_3975);
and U9305 (N_9305,N_1428,N_388);
nand U9306 (N_9306,N_4378,N_4058);
nor U9307 (N_9307,N_3411,N_544);
xor U9308 (N_9308,N_1564,N_4703);
nand U9309 (N_9309,N_619,N_3579);
xor U9310 (N_9310,N_2384,N_1582);
or U9311 (N_9311,N_3060,N_849);
or U9312 (N_9312,N_2626,N_1078);
xnor U9313 (N_9313,N_379,N_2238);
and U9314 (N_9314,N_3543,N_4469);
nor U9315 (N_9315,N_809,N_3957);
nor U9316 (N_9316,N_124,N_4754);
and U9317 (N_9317,N_1720,N_4106);
nor U9318 (N_9318,N_1929,N_4974);
or U9319 (N_9319,N_1900,N_1720);
nor U9320 (N_9320,N_3904,N_1090);
xor U9321 (N_9321,N_106,N_2999);
nor U9322 (N_9322,N_4319,N_3457);
and U9323 (N_9323,N_2816,N_3833);
or U9324 (N_9324,N_362,N_3986);
nand U9325 (N_9325,N_2851,N_3831);
and U9326 (N_9326,N_1792,N_3455);
nand U9327 (N_9327,N_2903,N_1471);
or U9328 (N_9328,N_4034,N_3941);
nor U9329 (N_9329,N_917,N_819);
nor U9330 (N_9330,N_2361,N_2246);
nor U9331 (N_9331,N_3512,N_3274);
nand U9332 (N_9332,N_3274,N_1564);
and U9333 (N_9333,N_449,N_2961);
nor U9334 (N_9334,N_4634,N_832);
nor U9335 (N_9335,N_4859,N_1036);
or U9336 (N_9336,N_2692,N_3073);
nand U9337 (N_9337,N_339,N_1833);
xnor U9338 (N_9338,N_447,N_1260);
xor U9339 (N_9339,N_4816,N_756);
xnor U9340 (N_9340,N_463,N_678);
or U9341 (N_9341,N_1017,N_646);
and U9342 (N_9342,N_3461,N_3960);
nand U9343 (N_9343,N_4416,N_4651);
nor U9344 (N_9344,N_732,N_56);
nand U9345 (N_9345,N_1698,N_3178);
or U9346 (N_9346,N_1051,N_1074);
xnor U9347 (N_9347,N_3448,N_995);
or U9348 (N_9348,N_1561,N_943);
or U9349 (N_9349,N_734,N_687);
xor U9350 (N_9350,N_2725,N_1073);
and U9351 (N_9351,N_222,N_1420);
xnor U9352 (N_9352,N_1708,N_181);
xor U9353 (N_9353,N_3155,N_323);
and U9354 (N_9354,N_2383,N_645);
and U9355 (N_9355,N_1056,N_458);
nor U9356 (N_9356,N_212,N_998);
and U9357 (N_9357,N_3117,N_4936);
or U9358 (N_9358,N_759,N_2080);
and U9359 (N_9359,N_872,N_1589);
and U9360 (N_9360,N_3406,N_3055);
xor U9361 (N_9361,N_2572,N_2519);
nor U9362 (N_9362,N_3609,N_189);
xnor U9363 (N_9363,N_1831,N_4843);
xnor U9364 (N_9364,N_732,N_1808);
and U9365 (N_9365,N_859,N_3392);
xor U9366 (N_9366,N_4240,N_1154);
nand U9367 (N_9367,N_3151,N_2302);
nand U9368 (N_9368,N_1880,N_2668);
or U9369 (N_9369,N_3645,N_2406);
nor U9370 (N_9370,N_1498,N_1673);
nand U9371 (N_9371,N_1243,N_2395);
nor U9372 (N_9372,N_404,N_1324);
nor U9373 (N_9373,N_4522,N_4150);
and U9374 (N_9374,N_3559,N_4738);
or U9375 (N_9375,N_423,N_4136);
nand U9376 (N_9376,N_1594,N_2013);
nand U9377 (N_9377,N_2547,N_134);
and U9378 (N_9378,N_3923,N_4761);
and U9379 (N_9379,N_1842,N_518);
xor U9380 (N_9380,N_2750,N_4094);
xnor U9381 (N_9381,N_3484,N_1872);
nor U9382 (N_9382,N_4513,N_3407);
or U9383 (N_9383,N_1419,N_657);
nor U9384 (N_9384,N_417,N_465);
and U9385 (N_9385,N_2627,N_1356);
or U9386 (N_9386,N_3084,N_875);
or U9387 (N_9387,N_3783,N_379);
nor U9388 (N_9388,N_3240,N_181);
or U9389 (N_9389,N_1556,N_3709);
and U9390 (N_9390,N_4666,N_1069);
or U9391 (N_9391,N_3046,N_4994);
nor U9392 (N_9392,N_4271,N_3744);
and U9393 (N_9393,N_3012,N_3267);
nor U9394 (N_9394,N_4022,N_1708);
xor U9395 (N_9395,N_3976,N_831);
nor U9396 (N_9396,N_79,N_4585);
xnor U9397 (N_9397,N_2977,N_2237);
or U9398 (N_9398,N_2592,N_3151);
nor U9399 (N_9399,N_4243,N_2113);
or U9400 (N_9400,N_4882,N_2387);
and U9401 (N_9401,N_3585,N_2155);
and U9402 (N_9402,N_1393,N_1826);
or U9403 (N_9403,N_4531,N_1340);
nor U9404 (N_9404,N_3361,N_3286);
or U9405 (N_9405,N_4238,N_4419);
or U9406 (N_9406,N_1611,N_1694);
or U9407 (N_9407,N_547,N_3349);
and U9408 (N_9408,N_302,N_2538);
and U9409 (N_9409,N_1326,N_4708);
and U9410 (N_9410,N_4811,N_122);
and U9411 (N_9411,N_2797,N_2862);
xor U9412 (N_9412,N_3899,N_3636);
or U9413 (N_9413,N_3317,N_238);
nor U9414 (N_9414,N_3117,N_1664);
nor U9415 (N_9415,N_1550,N_2696);
and U9416 (N_9416,N_4248,N_4632);
or U9417 (N_9417,N_1189,N_4557);
nand U9418 (N_9418,N_594,N_433);
xor U9419 (N_9419,N_61,N_4834);
xnor U9420 (N_9420,N_1553,N_1660);
and U9421 (N_9421,N_4099,N_4875);
and U9422 (N_9422,N_2835,N_1570);
nand U9423 (N_9423,N_4925,N_2066);
nand U9424 (N_9424,N_1066,N_775);
and U9425 (N_9425,N_764,N_1440);
and U9426 (N_9426,N_1083,N_4982);
and U9427 (N_9427,N_1543,N_113);
nor U9428 (N_9428,N_4347,N_3622);
and U9429 (N_9429,N_491,N_2521);
or U9430 (N_9430,N_4653,N_3991);
and U9431 (N_9431,N_1255,N_3906);
and U9432 (N_9432,N_4145,N_445);
xor U9433 (N_9433,N_4405,N_249);
and U9434 (N_9434,N_478,N_1783);
or U9435 (N_9435,N_4292,N_2435);
and U9436 (N_9436,N_53,N_2817);
nor U9437 (N_9437,N_1524,N_524);
nand U9438 (N_9438,N_2968,N_895);
nor U9439 (N_9439,N_4420,N_3076);
nand U9440 (N_9440,N_3745,N_3243);
nand U9441 (N_9441,N_2196,N_1644);
or U9442 (N_9442,N_2570,N_2111);
nor U9443 (N_9443,N_213,N_1701);
and U9444 (N_9444,N_54,N_2614);
and U9445 (N_9445,N_4982,N_771);
nand U9446 (N_9446,N_1492,N_638);
xnor U9447 (N_9447,N_1185,N_3738);
nand U9448 (N_9448,N_2396,N_1010);
or U9449 (N_9449,N_634,N_1780);
or U9450 (N_9450,N_3004,N_2743);
nor U9451 (N_9451,N_1019,N_4264);
xnor U9452 (N_9452,N_1734,N_1113);
nor U9453 (N_9453,N_2317,N_2082);
nor U9454 (N_9454,N_519,N_2686);
nor U9455 (N_9455,N_4908,N_675);
xnor U9456 (N_9456,N_2971,N_4134);
xnor U9457 (N_9457,N_4386,N_1706);
nor U9458 (N_9458,N_3251,N_3388);
and U9459 (N_9459,N_3819,N_3576);
xnor U9460 (N_9460,N_747,N_1137);
nand U9461 (N_9461,N_2754,N_1179);
or U9462 (N_9462,N_3259,N_3767);
nor U9463 (N_9463,N_1861,N_2826);
or U9464 (N_9464,N_1650,N_3469);
xor U9465 (N_9465,N_642,N_3505);
or U9466 (N_9466,N_3764,N_1926);
nand U9467 (N_9467,N_286,N_459);
or U9468 (N_9468,N_722,N_3568);
or U9469 (N_9469,N_1884,N_3366);
and U9470 (N_9470,N_4935,N_2586);
nor U9471 (N_9471,N_4903,N_687);
or U9472 (N_9472,N_3421,N_2999);
nor U9473 (N_9473,N_1160,N_2085);
and U9474 (N_9474,N_3859,N_1991);
and U9475 (N_9475,N_537,N_4005);
nand U9476 (N_9476,N_4413,N_2314);
and U9477 (N_9477,N_4989,N_643);
nand U9478 (N_9478,N_3586,N_241);
and U9479 (N_9479,N_1729,N_2894);
xnor U9480 (N_9480,N_1694,N_1722);
nor U9481 (N_9481,N_3334,N_2136);
or U9482 (N_9482,N_964,N_4762);
xor U9483 (N_9483,N_3643,N_4162);
nor U9484 (N_9484,N_1729,N_4720);
or U9485 (N_9485,N_679,N_3956);
and U9486 (N_9486,N_4264,N_355);
xor U9487 (N_9487,N_2581,N_4743);
nand U9488 (N_9488,N_2312,N_413);
or U9489 (N_9489,N_1925,N_3197);
xnor U9490 (N_9490,N_3313,N_1705);
or U9491 (N_9491,N_402,N_4044);
xnor U9492 (N_9492,N_3951,N_4348);
nand U9493 (N_9493,N_4813,N_3777);
nor U9494 (N_9494,N_3787,N_1030);
and U9495 (N_9495,N_650,N_301);
or U9496 (N_9496,N_2697,N_2369);
nor U9497 (N_9497,N_3252,N_2601);
nand U9498 (N_9498,N_3736,N_3586);
nor U9499 (N_9499,N_2159,N_2271);
nor U9500 (N_9500,N_271,N_2120);
and U9501 (N_9501,N_3045,N_3503);
and U9502 (N_9502,N_3058,N_769);
xor U9503 (N_9503,N_2085,N_2311);
nor U9504 (N_9504,N_3306,N_4577);
or U9505 (N_9505,N_1341,N_4560);
nor U9506 (N_9506,N_2828,N_2036);
nor U9507 (N_9507,N_2295,N_3131);
nand U9508 (N_9508,N_4561,N_4023);
or U9509 (N_9509,N_390,N_4146);
and U9510 (N_9510,N_1514,N_3139);
xor U9511 (N_9511,N_2956,N_4245);
or U9512 (N_9512,N_927,N_605);
and U9513 (N_9513,N_3616,N_2538);
and U9514 (N_9514,N_2868,N_1356);
and U9515 (N_9515,N_2533,N_1454);
and U9516 (N_9516,N_3127,N_2749);
nand U9517 (N_9517,N_4622,N_4198);
xnor U9518 (N_9518,N_2072,N_4842);
nand U9519 (N_9519,N_4202,N_3165);
nor U9520 (N_9520,N_2867,N_1007);
and U9521 (N_9521,N_4077,N_2401);
or U9522 (N_9522,N_2275,N_2092);
nor U9523 (N_9523,N_2462,N_2439);
or U9524 (N_9524,N_2476,N_3102);
xnor U9525 (N_9525,N_4868,N_1363);
nor U9526 (N_9526,N_401,N_2863);
or U9527 (N_9527,N_4535,N_2548);
xor U9528 (N_9528,N_788,N_2141);
and U9529 (N_9529,N_871,N_4805);
nand U9530 (N_9530,N_2946,N_3977);
nor U9531 (N_9531,N_2724,N_2729);
nor U9532 (N_9532,N_2479,N_3500);
nand U9533 (N_9533,N_1886,N_19);
xor U9534 (N_9534,N_2338,N_3602);
xnor U9535 (N_9535,N_4287,N_709);
nand U9536 (N_9536,N_1131,N_4603);
xor U9537 (N_9537,N_1735,N_1884);
or U9538 (N_9538,N_1048,N_3729);
nor U9539 (N_9539,N_3141,N_3953);
nand U9540 (N_9540,N_4226,N_107);
nand U9541 (N_9541,N_437,N_4637);
nand U9542 (N_9542,N_4735,N_933);
nand U9543 (N_9543,N_2935,N_3984);
or U9544 (N_9544,N_2762,N_791);
nor U9545 (N_9545,N_4288,N_2256);
and U9546 (N_9546,N_4561,N_4339);
and U9547 (N_9547,N_287,N_4012);
or U9548 (N_9548,N_4454,N_3479);
and U9549 (N_9549,N_2229,N_1389);
nor U9550 (N_9550,N_4312,N_1002);
xor U9551 (N_9551,N_870,N_1249);
nand U9552 (N_9552,N_2145,N_4708);
xnor U9553 (N_9553,N_1992,N_3148);
nand U9554 (N_9554,N_1336,N_3386);
xor U9555 (N_9555,N_311,N_2169);
xor U9556 (N_9556,N_4430,N_4371);
or U9557 (N_9557,N_4494,N_112);
and U9558 (N_9558,N_2616,N_3765);
nor U9559 (N_9559,N_4352,N_1806);
nand U9560 (N_9560,N_3652,N_2120);
nand U9561 (N_9561,N_2710,N_587);
xnor U9562 (N_9562,N_1758,N_2901);
and U9563 (N_9563,N_2625,N_1892);
or U9564 (N_9564,N_698,N_706);
nor U9565 (N_9565,N_540,N_3510);
or U9566 (N_9566,N_1901,N_4945);
and U9567 (N_9567,N_3652,N_3470);
or U9568 (N_9568,N_4966,N_3426);
and U9569 (N_9569,N_2315,N_244);
or U9570 (N_9570,N_3044,N_230);
nor U9571 (N_9571,N_1844,N_4390);
and U9572 (N_9572,N_1259,N_3685);
nand U9573 (N_9573,N_3625,N_4550);
or U9574 (N_9574,N_4257,N_2455);
xor U9575 (N_9575,N_1854,N_3256);
nand U9576 (N_9576,N_4813,N_2291);
xor U9577 (N_9577,N_4326,N_370);
and U9578 (N_9578,N_3724,N_573);
xor U9579 (N_9579,N_268,N_1429);
xnor U9580 (N_9580,N_3259,N_1784);
xnor U9581 (N_9581,N_3865,N_27);
nand U9582 (N_9582,N_4286,N_2036);
xor U9583 (N_9583,N_4041,N_2120);
and U9584 (N_9584,N_4574,N_802);
nor U9585 (N_9585,N_659,N_1430);
and U9586 (N_9586,N_3812,N_4197);
and U9587 (N_9587,N_2032,N_797);
or U9588 (N_9588,N_2815,N_4116);
nor U9589 (N_9589,N_2660,N_97);
and U9590 (N_9590,N_122,N_4232);
nor U9591 (N_9591,N_2697,N_1513);
nand U9592 (N_9592,N_1787,N_3600);
xnor U9593 (N_9593,N_2351,N_3719);
nor U9594 (N_9594,N_1325,N_2386);
nand U9595 (N_9595,N_1459,N_4230);
and U9596 (N_9596,N_3218,N_2474);
or U9597 (N_9597,N_521,N_2922);
and U9598 (N_9598,N_1529,N_841);
and U9599 (N_9599,N_156,N_1467);
and U9600 (N_9600,N_1047,N_2156);
or U9601 (N_9601,N_2552,N_2471);
nand U9602 (N_9602,N_4935,N_2032);
and U9603 (N_9603,N_4838,N_4080);
nor U9604 (N_9604,N_1359,N_2698);
nand U9605 (N_9605,N_258,N_3332);
nor U9606 (N_9606,N_2736,N_1669);
and U9607 (N_9607,N_4750,N_2088);
or U9608 (N_9608,N_4000,N_2068);
xnor U9609 (N_9609,N_2832,N_541);
and U9610 (N_9610,N_1620,N_2398);
or U9611 (N_9611,N_4691,N_3361);
or U9612 (N_9612,N_1882,N_679);
nand U9613 (N_9613,N_2590,N_2490);
or U9614 (N_9614,N_3583,N_151);
nand U9615 (N_9615,N_3653,N_2158);
xor U9616 (N_9616,N_912,N_3630);
xnor U9617 (N_9617,N_38,N_3390);
or U9618 (N_9618,N_169,N_41);
nand U9619 (N_9619,N_2421,N_2570);
or U9620 (N_9620,N_4511,N_1256);
nand U9621 (N_9621,N_1998,N_3770);
or U9622 (N_9622,N_3016,N_45);
and U9623 (N_9623,N_3081,N_2233);
or U9624 (N_9624,N_245,N_660);
nand U9625 (N_9625,N_680,N_4065);
or U9626 (N_9626,N_2555,N_2278);
or U9627 (N_9627,N_2252,N_1745);
xnor U9628 (N_9628,N_3480,N_3519);
nand U9629 (N_9629,N_3174,N_4421);
nor U9630 (N_9630,N_4557,N_755);
nand U9631 (N_9631,N_116,N_73);
nor U9632 (N_9632,N_2556,N_3348);
or U9633 (N_9633,N_2308,N_753);
nor U9634 (N_9634,N_4524,N_4077);
nand U9635 (N_9635,N_2355,N_2598);
or U9636 (N_9636,N_471,N_4640);
and U9637 (N_9637,N_2047,N_721);
or U9638 (N_9638,N_876,N_4778);
nand U9639 (N_9639,N_2822,N_2076);
nand U9640 (N_9640,N_2016,N_3701);
and U9641 (N_9641,N_4315,N_325);
or U9642 (N_9642,N_772,N_2282);
or U9643 (N_9643,N_2444,N_2670);
and U9644 (N_9644,N_3030,N_3041);
nand U9645 (N_9645,N_1048,N_308);
xnor U9646 (N_9646,N_2617,N_2360);
xnor U9647 (N_9647,N_3198,N_2120);
or U9648 (N_9648,N_4705,N_4260);
nand U9649 (N_9649,N_1162,N_3639);
xnor U9650 (N_9650,N_756,N_946);
or U9651 (N_9651,N_628,N_2590);
nand U9652 (N_9652,N_666,N_2660);
xor U9653 (N_9653,N_4217,N_1084);
and U9654 (N_9654,N_747,N_925);
xor U9655 (N_9655,N_1739,N_1706);
or U9656 (N_9656,N_2183,N_1090);
xnor U9657 (N_9657,N_663,N_122);
nand U9658 (N_9658,N_4686,N_4241);
xnor U9659 (N_9659,N_671,N_206);
and U9660 (N_9660,N_4114,N_4418);
nand U9661 (N_9661,N_1912,N_417);
or U9662 (N_9662,N_170,N_4815);
and U9663 (N_9663,N_1495,N_719);
and U9664 (N_9664,N_3583,N_271);
or U9665 (N_9665,N_1272,N_4433);
and U9666 (N_9666,N_4398,N_4587);
nand U9667 (N_9667,N_2631,N_4315);
and U9668 (N_9668,N_3240,N_4576);
or U9669 (N_9669,N_1996,N_4601);
nand U9670 (N_9670,N_2195,N_843);
or U9671 (N_9671,N_299,N_4714);
nor U9672 (N_9672,N_2171,N_4941);
nor U9673 (N_9673,N_1758,N_3866);
nand U9674 (N_9674,N_920,N_4098);
nand U9675 (N_9675,N_3953,N_962);
or U9676 (N_9676,N_143,N_4151);
and U9677 (N_9677,N_4721,N_3610);
and U9678 (N_9678,N_2879,N_107);
nand U9679 (N_9679,N_3785,N_3673);
or U9680 (N_9680,N_984,N_4972);
and U9681 (N_9681,N_4832,N_2641);
or U9682 (N_9682,N_981,N_2534);
nor U9683 (N_9683,N_3742,N_2212);
xnor U9684 (N_9684,N_525,N_208);
nor U9685 (N_9685,N_519,N_588);
and U9686 (N_9686,N_4044,N_3956);
nor U9687 (N_9687,N_2254,N_3329);
and U9688 (N_9688,N_1386,N_1506);
xnor U9689 (N_9689,N_1196,N_3200);
and U9690 (N_9690,N_2863,N_187);
xor U9691 (N_9691,N_3275,N_4241);
or U9692 (N_9692,N_2135,N_1855);
xor U9693 (N_9693,N_204,N_1436);
xor U9694 (N_9694,N_4618,N_4323);
nor U9695 (N_9695,N_4709,N_3853);
nand U9696 (N_9696,N_2434,N_152);
and U9697 (N_9697,N_2733,N_4211);
or U9698 (N_9698,N_441,N_4463);
nand U9699 (N_9699,N_2166,N_3131);
xor U9700 (N_9700,N_4187,N_2418);
or U9701 (N_9701,N_4263,N_3291);
nand U9702 (N_9702,N_4838,N_1980);
nand U9703 (N_9703,N_3417,N_2469);
or U9704 (N_9704,N_388,N_3790);
nor U9705 (N_9705,N_374,N_4098);
xor U9706 (N_9706,N_4928,N_2703);
nor U9707 (N_9707,N_1762,N_2791);
nor U9708 (N_9708,N_3364,N_3326);
nand U9709 (N_9709,N_2559,N_836);
xor U9710 (N_9710,N_4347,N_3703);
and U9711 (N_9711,N_4376,N_1391);
nor U9712 (N_9712,N_3789,N_3749);
xnor U9713 (N_9713,N_2588,N_3221);
nand U9714 (N_9714,N_1376,N_1444);
xor U9715 (N_9715,N_3847,N_2031);
xor U9716 (N_9716,N_3561,N_4008);
nor U9717 (N_9717,N_306,N_3481);
and U9718 (N_9718,N_653,N_716);
xnor U9719 (N_9719,N_3766,N_3189);
nor U9720 (N_9720,N_2301,N_1981);
and U9721 (N_9721,N_352,N_475);
or U9722 (N_9722,N_193,N_4303);
and U9723 (N_9723,N_2379,N_4617);
xor U9724 (N_9724,N_1132,N_714);
nor U9725 (N_9725,N_1906,N_1054);
nand U9726 (N_9726,N_4222,N_3985);
xnor U9727 (N_9727,N_4294,N_257);
and U9728 (N_9728,N_414,N_4631);
nor U9729 (N_9729,N_1138,N_4308);
nor U9730 (N_9730,N_3149,N_4731);
nor U9731 (N_9731,N_4488,N_2018);
xnor U9732 (N_9732,N_3781,N_3873);
nor U9733 (N_9733,N_3297,N_86);
nor U9734 (N_9734,N_1866,N_1503);
xnor U9735 (N_9735,N_3970,N_4451);
and U9736 (N_9736,N_2820,N_967);
or U9737 (N_9737,N_466,N_4789);
or U9738 (N_9738,N_4738,N_2845);
and U9739 (N_9739,N_1397,N_748);
and U9740 (N_9740,N_3273,N_2061);
nor U9741 (N_9741,N_3611,N_350);
xnor U9742 (N_9742,N_2880,N_1859);
nand U9743 (N_9743,N_3230,N_643);
or U9744 (N_9744,N_1249,N_731);
nand U9745 (N_9745,N_1450,N_3319);
nor U9746 (N_9746,N_3668,N_3694);
nand U9747 (N_9747,N_3698,N_947);
nand U9748 (N_9748,N_2622,N_730);
nand U9749 (N_9749,N_2353,N_72);
and U9750 (N_9750,N_2587,N_3016);
nand U9751 (N_9751,N_3451,N_1523);
or U9752 (N_9752,N_661,N_2488);
nand U9753 (N_9753,N_1455,N_328);
xor U9754 (N_9754,N_797,N_401);
or U9755 (N_9755,N_3715,N_4019);
or U9756 (N_9756,N_2931,N_3474);
nand U9757 (N_9757,N_4050,N_4132);
or U9758 (N_9758,N_2391,N_567);
or U9759 (N_9759,N_772,N_2078);
nand U9760 (N_9760,N_1086,N_2764);
or U9761 (N_9761,N_24,N_3598);
nor U9762 (N_9762,N_2349,N_2861);
nand U9763 (N_9763,N_4254,N_885);
xnor U9764 (N_9764,N_4692,N_928);
or U9765 (N_9765,N_4677,N_3884);
nor U9766 (N_9766,N_4347,N_1534);
nand U9767 (N_9767,N_4553,N_2804);
xnor U9768 (N_9768,N_627,N_2567);
nand U9769 (N_9769,N_1622,N_696);
and U9770 (N_9770,N_4234,N_4981);
nand U9771 (N_9771,N_4900,N_387);
and U9772 (N_9772,N_3789,N_2802);
or U9773 (N_9773,N_447,N_1032);
xnor U9774 (N_9774,N_2584,N_1542);
xnor U9775 (N_9775,N_4121,N_3001);
nand U9776 (N_9776,N_1564,N_2245);
nor U9777 (N_9777,N_890,N_3566);
nand U9778 (N_9778,N_1282,N_144);
and U9779 (N_9779,N_183,N_1443);
nor U9780 (N_9780,N_2140,N_4384);
and U9781 (N_9781,N_128,N_549);
nand U9782 (N_9782,N_3780,N_3666);
or U9783 (N_9783,N_4263,N_4350);
xnor U9784 (N_9784,N_4308,N_2766);
nor U9785 (N_9785,N_1317,N_1607);
xor U9786 (N_9786,N_579,N_1361);
or U9787 (N_9787,N_3311,N_1651);
and U9788 (N_9788,N_2172,N_2537);
nor U9789 (N_9789,N_1856,N_1776);
nor U9790 (N_9790,N_2942,N_3889);
nand U9791 (N_9791,N_4392,N_4355);
and U9792 (N_9792,N_3564,N_3806);
or U9793 (N_9793,N_852,N_4472);
nand U9794 (N_9794,N_1664,N_973);
nand U9795 (N_9795,N_4905,N_2327);
and U9796 (N_9796,N_665,N_2041);
or U9797 (N_9797,N_703,N_4614);
xor U9798 (N_9798,N_1602,N_3343);
xor U9799 (N_9799,N_1389,N_63);
xnor U9800 (N_9800,N_1583,N_3594);
or U9801 (N_9801,N_622,N_558);
or U9802 (N_9802,N_3520,N_763);
nor U9803 (N_9803,N_1738,N_4388);
xnor U9804 (N_9804,N_1532,N_4220);
nor U9805 (N_9805,N_3681,N_1488);
nand U9806 (N_9806,N_3310,N_3237);
nand U9807 (N_9807,N_3415,N_1139);
nand U9808 (N_9808,N_3834,N_1980);
or U9809 (N_9809,N_3477,N_3584);
and U9810 (N_9810,N_1418,N_2858);
or U9811 (N_9811,N_704,N_2661);
or U9812 (N_9812,N_124,N_2705);
nor U9813 (N_9813,N_3615,N_4827);
xnor U9814 (N_9814,N_3776,N_2179);
and U9815 (N_9815,N_228,N_3681);
nor U9816 (N_9816,N_4297,N_2857);
nor U9817 (N_9817,N_4550,N_4306);
and U9818 (N_9818,N_2073,N_3992);
nor U9819 (N_9819,N_3312,N_4190);
xor U9820 (N_9820,N_2087,N_983);
xnor U9821 (N_9821,N_1123,N_3553);
or U9822 (N_9822,N_1133,N_3708);
nand U9823 (N_9823,N_1700,N_4221);
xnor U9824 (N_9824,N_3935,N_3557);
and U9825 (N_9825,N_3798,N_1308);
xnor U9826 (N_9826,N_1648,N_2019);
nor U9827 (N_9827,N_1850,N_4731);
xor U9828 (N_9828,N_1990,N_657);
nand U9829 (N_9829,N_965,N_841);
nand U9830 (N_9830,N_182,N_2454);
and U9831 (N_9831,N_605,N_80);
and U9832 (N_9832,N_2091,N_1508);
nor U9833 (N_9833,N_4870,N_2459);
nor U9834 (N_9834,N_3485,N_3403);
and U9835 (N_9835,N_520,N_1249);
or U9836 (N_9836,N_283,N_2359);
and U9837 (N_9837,N_1274,N_1529);
and U9838 (N_9838,N_2929,N_2692);
and U9839 (N_9839,N_3432,N_1950);
nand U9840 (N_9840,N_2772,N_252);
or U9841 (N_9841,N_1936,N_894);
and U9842 (N_9842,N_3179,N_4990);
nor U9843 (N_9843,N_550,N_1389);
nand U9844 (N_9844,N_3814,N_871);
xnor U9845 (N_9845,N_1297,N_2821);
nor U9846 (N_9846,N_1094,N_391);
or U9847 (N_9847,N_2768,N_2277);
and U9848 (N_9848,N_3177,N_668);
nor U9849 (N_9849,N_2116,N_1347);
or U9850 (N_9850,N_3856,N_4606);
or U9851 (N_9851,N_1406,N_4811);
xnor U9852 (N_9852,N_3771,N_71);
nand U9853 (N_9853,N_4092,N_2569);
or U9854 (N_9854,N_2502,N_3669);
or U9855 (N_9855,N_4133,N_92);
or U9856 (N_9856,N_2415,N_3950);
or U9857 (N_9857,N_1814,N_1518);
or U9858 (N_9858,N_366,N_2555);
xnor U9859 (N_9859,N_4808,N_1356);
nor U9860 (N_9860,N_3482,N_2960);
xor U9861 (N_9861,N_4785,N_4212);
xnor U9862 (N_9862,N_2681,N_1778);
or U9863 (N_9863,N_2489,N_674);
xor U9864 (N_9864,N_4590,N_1917);
and U9865 (N_9865,N_2561,N_3400);
or U9866 (N_9866,N_3971,N_2071);
or U9867 (N_9867,N_3946,N_3883);
nand U9868 (N_9868,N_492,N_401);
or U9869 (N_9869,N_2649,N_3715);
xnor U9870 (N_9870,N_1909,N_295);
nand U9871 (N_9871,N_4973,N_3254);
nand U9872 (N_9872,N_3847,N_4857);
nor U9873 (N_9873,N_1765,N_1891);
nor U9874 (N_9874,N_3404,N_195);
xnor U9875 (N_9875,N_471,N_1068);
nand U9876 (N_9876,N_2429,N_1247);
nand U9877 (N_9877,N_4954,N_2938);
and U9878 (N_9878,N_1117,N_3366);
nor U9879 (N_9879,N_3385,N_498);
and U9880 (N_9880,N_3777,N_3941);
nand U9881 (N_9881,N_4049,N_1245);
and U9882 (N_9882,N_4759,N_3932);
and U9883 (N_9883,N_4403,N_2757);
or U9884 (N_9884,N_3014,N_1754);
nor U9885 (N_9885,N_344,N_2651);
and U9886 (N_9886,N_4754,N_2059);
or U9887 (N_9887,N_52,N_4422);
nand U9888 (N_9888,N_2125,N_3201);
nor U9889 (N_9889,N_1703,N_942);
and U9890 (N_9890,N_2020,N_2995);
or U9891 (N_9891,N_87,N_433);
nand U9892 (N_9892,N_3877,N_2395);
nor U9893 (N_9893,N_3909,N_2324);
or U9894 (N_9894,N_3982,N_930);
nor U9895 (N_9895,N_103,N_4543);
nand U9896 (N_9896,N_2718,N_15);
nor U9897 (N_9897,N_702,N_1120);
or U9898 (N_9898,N_479,N_3112);
xnor U9899 (N_9899,N_849,N_3831);
xnor U9900 (N_9900,N_2708,N_16);
xnor U9901 (N_9901,N_2709,N_255);
or U9902 (N_9902,N_4601,N_479);
nand U9903 (N_9903,N_1122,N_3587);
xnor U9904 (N_9904,N_4702,N_2745);
nor U9905 (N_9905,N_2305,N_4206);
nand U9906 (N_9906,N_4258,N_2917);
or U9907 (N_9907,N_1192,N_4375);
and U9908 (N_9908,N_551,N_1863);
and U9909 (N_9909,N_622,N_4590);
xor U9910 (N_9910,N_790,N_4864);
nand U9911 (N_9911,N_1659,N_4980);
nand U9912 (N_9912,N_4161,N_2292);
and U9913 (N_9913,N_3924,N_953);
xor U9914 (N_9914,N_4539,N_2445);
and U9915 (N_9915,N_3750,N_247);
and U9916 (N_9916,N_48,N_2824);
nor U9917 (N_9917,N_2621,N_4542);
nand U9918 (N_9918,N_4909,N_3409);
or U9919 (N_9919,N_1044,N_3543);
xnor U9920 (N_9920,N_2586,N_4107);
xor U9921 (N_9921,N_3341,N_116);
xor U9922 (N_9922,N_2218,N_978);
nand U9923 (N_9923,N_2927,N_1942);
and U9924 (N_9924,N_2684,N_2043);
xor U9925 (N_9925,N_4197,N_2785);
or U9926 (N_9926,N_3006,N_4842);
xnor U9927 (N_9927,N_1258,N_640);
nor U9928 (N_9928,N_303,N_4699);
or U9929 (N_9929,N_2495,N_4064);
or U9930 (N_9930,N_4369,N_2186);
xnor U9931 (N_9931,N_1074,N_4269);
or U9932 (N_9932,N_1607,N_2103);
nand U9933 (N_9933,N_1711,N_2417);
nand U9934 (N_9934,N_327,N_268);
and U9935 (N_9935,N_782,N_1248);
xor U9936 (N_9936,N_1995,N_4595);
nand U9937 (N_9937,N_278,N_744);
xor U9938 (N_9938,N_4425,N_3595);
nand U9939 (N_9939,N_4347,N_3388);
or U9940 (N_9940,N_1226,N_2262);
or U9941 (N_9941,N_1950,N_3697);
or U9942 (N_9942,N_2274,N_4715);
nand U9943 (N_9943,N_1224,N_647);
nand U9944 (N_9944,N_1512,N_4031);
and U9945 (N_9945,N_3046,N_3062);
or U9946 (N_9946,N_2788,N_2214);
nor U9947 (N_9947,N_3055,N_3649);
or U9948 (N_9948,N_2367,N_1464);
xnor U9949 (N_9949,N_3340,N_786);
nor U9950 (N_9950,N_930,N_26);
xnor U9951 (N_9951,N_1746,N_2672);
and U9952 (N_9952,N_2377,N_439);
and U9953 (N_9953,N_109,N_716);
or U9954 (N_9954,N_4152,N_1431);
xnor U9955 (N_9955,N_2206,N_3981);
nor U9956 (N_9956,N_4220,N_4319);
and U9957 (N_9957,N_322,N_4623);
xor U9958 (N_9958,N_1066,N_826);
or U9959 (N_9959,N_202,N_59);
xor U9960 (N_9960,N_3707,N_1481);
nor U9961 (N_9961,N_2200,N_1732);
nand U9962 (N_9962,N_1135,N_1747);
or U9963 (N_9963,N_1359,N_4809);
and U9964 (N_9964,N_664,N_4941);
xnor U9965 (N_9965,N_3603,N_4276);
or U9966 (N_9966,N_3517,N_2002);
or U9967 (N_9967,N_4476,N_884);
xnor U9968 (N_9968,N_3135,N_1126);
or U9969 (N_9969,N_636,N_1210);
or U9970 (N_9970,N_1179,N_88);
and U9971 (N_9971,N_1201,N_1159);
xor U9972 (N_9972,N_3160,N_4318);
and U9973 (N_9973,N_4948,N_3424);
nor U9974 (N_9974,N_3589,N_464);
nor U9975 (N_9975,N_2845,N_3);
xnor U9976 (N_9976,N_1487,N_1447);
xnor U9977 (N_9977,N_3893,N_2925);
xnor U9978 (N_9978,N_3502,N_3148);
and U9979 (N_9979,N_345,N_3900);
and U9980 (N_9980,N_2206,N_4011);
nand U9981 (N_9981,N_1692,N_181);
nor U9982 (N_9982,N_814,N_4840);
nor U9983 (N_9983,N_1396,N_3520);
xnor U9984 (N_9984,N_1532,N_3864);
nor U9985 (N_9985,N_3753,N_1444);
nand U9986 (N_9986,N_2215,N_4268);
nor U9987 (N_9987,N_1016,N_4110);
nand U9988 (N_9988,N_4287,N_423);
and U9989 (N_9989,N_3273,N_285);
nand U9990 (N_9990,N_3666,N_1347);
xor U9991 (N_9991,N_2375,N_4012);
nand U9992 (N_9992,N_2408,N_2137);
xnor U9993 (N_9993,N_2836,N_3791);
xor U9994 (N_9994,N_4281,N_2235);
nand U9995 (N_9995,N_3167,N_4193);
nand U9996 (N_9996,N_2685,N_205);
xnor U9997 (N_9997,N_849,N_3535);
nand U9998 (N_9998,N_4977,N_1102);
xor U9999 (N_9999,N_1756,N_3412);
and UO_0 (O_0,N_8676,N_7690);
and UO_1 (O_1,N_6641,N_9712);
xnor UO_2 (O_2,N_5547,N_5509);
nor UO_3 (O_3,N_5367,N_8063);
xnor UO_4 (O_4,N_5272,N_8861);
xnor UO_5 (O_5,N_9074,N_7383);
nand UO_6 (O_6,N_7153,N_5582);
nor UO_7 (O_7,N_5484,N_7205);
xor UO_8 (O_8,N_9887,N_6371);
nand UO_9 (O_9,N_8529,N_7305);
nand UO_10 (O_10,N_9959,N_9643);
nor UO_11 (O_11,N_6258,N_8275);
xnor UO_12 (O_12,N_9097,N_8776);
nand UO_13 (O_13,N_5472,N_9889);
nor UO_14 (O_14,N_9600,N_9691);
or UO_15 (O_15,N_9957,N_9397);
or UO_16 (O_16,N_9682,N_8762);
nor UO_17 (O_17,N_8986,N_9065);
xnor UO_18 (O_18,N_7729,N_7320);
nor UO_19 (O_19,N_7504,N_8469);
nand UO_20 (O_20,N_6969,N_6007);
nand UO_21 (O_21,N_8221,N_6410);
nand UO_22 (O_22,N_6148,N_6791);
and UO_23 (O_23,N_5563,N_7706);
nand UO_24 (O_24,N_9852,N_7820);
and UO_25 (O_25,N_8422,N_9817);
nand UO_26 (O_26,N_8091,N_7294);
nor UO_27 (O_27,N_6110,N_6160);
nor UO_28 (O_28,N_6737,N_5182);
and UO_29 (O_29,N_9858,N_5877);
and UO_30 (O_30,N_9301,N_6639);
nand UO_31 (O_31,N_7894,N_9325);
nor UO_32 (O_32,N_5525,N_5343);
and UO_33 (O_33,N_9737,N_6593);
nand UO_34 (O_34,N_8764,N_8364);
and UO_35 (O_35,N_9516,N_7458);
or UO_36 (O_36,N_5961,N_9193);
and UO_37 (O_37,N_8839,N_8238);
and UO_38 (O_38,N_9088,N_6460);
nand UO_39 (O_39,N_5541,N_7702);
nand UO_40 (O_40,N_6437,N_9322);
xor UO_41 (O_41,N_8338,N_6030);
xnor UO_42 (O_42,N_8104,N_9081);
or UO_43 (O_43,N_6067,N_9662);
or UO_44 (O_44,N_9206,N_5076);
nor UO_45 (O_45,N_8755,N_6069);
or UO_46 (O_46,N_8316,N_5848);
or UO_47 (O_47,N_8509,N_6779);
nor UO_48 (O_48,N_5178,N_9192);
and UO_49 (O_49,N_5963,N_8747);
nor UO_50 (O_50,N_7935,N_8416);
and UO_51 (O_51,N_5363,N_5399);
and UO_52 (O_52,N_7763,N_9071);
nor UO_53 (O_53,N_6119,N_8955);
nor UO_54 (O_54,N_5844,N_6858);
nor UO_55 (O_55,N_6363,N_7044);
and UO_56 (O_56,N_8409,N_9836);
nor UO_57 (O_57,N_8214,N_7622);
and UO_58 (O_58,N_6633,N_9938);
and UO_59 (O_59,N_6863,N_7859);
and UO_60 (O_60,N_9908,N_6153);
xnor UO_61 (O_61,N_5573,N_7169);
and UO_62 (O_62,N_6389,N_6351);
nand UO_63 (O_63,N_5777,N_7280);
nor UO_64 (O_64,N_5501,N_7877);
or UO_65 (O_65,N_9345,N_8133);
nor UO_66 (O_66,N_7142,N_9160);
or UO_67 (O_67,N_9106,N_9329);
and UO_68 (O_68,N_8627,N_5658);
nand UO_69 (O_69,N_7532,N_6554);
nand UO_70 (O_70,N_9262,N_9586);
or UO_71 (O_71,N_9229,N_9320);
xor UO_72 (O_72,N_7290,N_9393);
nand UO_73 (O_73,N_7470,N_7834);
nor UO_74 (O_74,N_9116,N_7051);
or UO_75 (O_75,N_8772,N_8150);
or UO_76 (O_76,N_9421,N_9238);
xnor UO_77 (O_77,N_9802,N_6142);
and UO_78 (O_78,N_5995,N_7033);
and UO_79 (O_79,N_8306,N_8893);
or UO_80 (O_80,N_7122,N_5720);
nand UO_81 (O_81,N_5202,N_5846);
nor UO_82 (O_82,N_5560,N_5334);
nand UO_83 (O_83,N_7212,N_9696);
or UO_84 (O_84,N_7481,N_6444);
xor UO_85 (O_85,N_8400,N_9859);
and UO_86 (O_86,N_8212,N_6227);
or UO_87 (O_87,N_7448,N_9592);
or UO_88 (O_88,N_7524,N_8048);
nand UO_89 (O_89,N_9294,N_6947);
and UO_90 (O_90,N_5909,N_9865);
and UO_91 (O_91,N_6291,N_9306);
nor UO_92 (O_92,N_7891,N_6729);
and UO_93 (O_93,N_5829,N_9588);
or UO_94 (O_94,N_7115,N_8646);
nor UO_95 (O_95,N_5741,N_8428);
or UO_96 (O_96,N_7103,N_7302);
or UO_97 (O_97,N_5945,N_6994);
xnor UO_98 (O_98,N_9530,N_6465);
and UO_99 (O_99,N_6350,N_6908);
xnor UO_100 (O_100,N_7097,N_6373);
xor UO_101 (O_101,N_9313,N_9637);
xor UO_102 (O_102,N_5561,N_5569);
nor UO_103 (O_103,N_7911,N_7342);
xor UO_104 (O_104,N_8345,N_8468);
and UO_105 (O_105,N_8540,N_8097);
xor UO_106 (O_106,N_7746,N_8791);
or UO_107 (O_107,N_5216,N_5711);
nor UO_108 (O_108,N_8759,N_5129);
nor UO_109 (O_109,N_7041,N_8320);
and UO_110 (O_110,N_8494,N_5374);
xor UO_111 (O_111,N_7365,N_8752);
nor UO_112 (O_112,N_7256,N_9275);
xnor UO_113 (O_113,N_8911,N_6012);
and UO_114 (O_114,N_8821,N_5332);
or UO_115 (O_115,N_6210,N_5783);
and UO_116 (O_116,N_5247,N_5749);
nor UO_117 (O_117,N_6183,N_7572);
xor UO_118 (O_118,N_9727,N_7099);
nor UO_119 (O_119,N_6700,N_9508);
xor UO_120 (O_120,N_8837,N_5699);
nor UO_121 (O_121,N_6383,N_9907);
or UO_122 (O_122,N_5317,N_7052);
or UO_123 (O_123,N_6586,N_5971);
nor UO_124 (O_124,N_9069,N_6171);
and UO_125 (O_125,N_8901,N_5400);
xnor UO_126 (O_126,N_5762,N_7875);
nor UO_127 (O_127,N_5930,N_6960);
or UO_128 (O_128,N_8369,N_9510);
or UO_129 (O_129,N_7402,N_6050);
and UO_130 (O_130,N_5010,N_7126);
xor UO_131 (O_131,N_6271,N_6963);
xor UO_132 (O_132,N_5153,N_8183);
xor UO_133 (O_133,N_9906,N_7582);
xor UO_134 (O_134,N_6656,N_9025);
nand UO_135 (O_135,N_7726,N_7880);
nand UO_136 (O_136,N_7522,N_8426);
nand UO_137 (O_137,N_5973,N_6676);
nand UO_138 (O_138,N_7483,N_5227);
nand UO_139 (O_139,N_8350,N_7573);
and UO_140 (O_140,N_7425,N_5514);
nor UO_141 (O_141,N_8841,N_7919);
and UO_142 (O_142,N_5293,N_9356);
or UO_143 (O_143,N_7519,N_7083);
and UO_144 (O_144,N_7410,N_5127);
and UO_145 (O_145,N_5424,N_7835);
nand UO_146 (O_146,N_8708,N_5353);
or UO_147 (O_147,N_7436,N_5789);
xnor UO_148 (O_148,N_6115,N_8425);
nor UO_149 (O_149,N_5271,N_8295);
nor UO_150 (O_150,N_7494,N_8518);
or UO_151 (O_151,N_5904,N_8010);
and UO_152 (O_152,N_9225,N_7068);
and UO_153 (O_153,N_7846,N_8578);
nand UO_154 (O_154,N_8313,N_8789);
xnor UO_155 (O_155,N_6446,N_9828);
nor UO_156 (O_156,N_5964,N_7269);
and UO_157 (O_157,N_5689,N_5557);
nor UO_158 (O_158,N_6008,N_8291);
nor UO_159 (O_159,N_9248,N_9180);
nor UO_160 (O_160,N_6415,N_5905);
nor UO_161 (O_161,N_8510,N_7744);
xor UO_162 (O_162,N_6195,N_5092);
and UO_163 (O_163,N_8194,N_5387);
nand UO_164 (O_164,N_9656,N_6921);
nand UO_165 (O_165,N_9871,N_9834);
nand UO_166 (O_166,N_8822,N_6883);
or UO_167 (O_167,N_5906,N_6313);
nand UO_168 (O_168,N_8162,N_6747);
and UO_169 (O_169,N_8701,N_9361);
nor UO_170 (O_170,N_9960,N_5421);
or UO_171 (O_171,N_9654,N_9673);
nand UO_172 (O_172,N_7547,N_9235);
nor UO_173 (O_173,N_9680,N_5488);
and UO_174 (O_174,N_5009,N_9552);
nand UO_175 (O_175,N_7057,N_6321);
xnor UO_176 (O_176,N_6156,N_7246);
and UO_177 (O_177,N_7860,N_7511);
nand UO_178 (O_178,N_7249,N_7615);
and UO_179 (O_179,N_6730,N_9478);
or UO_180 (O_180,N_5377,N_5663);
xor UO_181 (O_181,N_7640,N_6901);
nand UO_182 (O_182,N_8365,N_5664);
xnor UO_183 (O_183,N_6771,N_9695);
and UO_184 (O_184,N_5411,N_7938);
or UO_185 (O_185,N_5589,N_6849);
nor UO_186 (O_186,N_8785,N_7457);
and UO_187 (O_187,N_6932,N_8012);
or UO_188 (O_188,N_5295,N_9561);
xnor UO_189 (O_189,N_6861,N_8667);
and UO_190 (O_190,N_5360,N_6900);
nand UO_191 (O_191,N_9410,N_6770);
and UO_192 (O_192,N_6343,N_5490);
nor UO_193 (O_193,N_5323,N_5853);
xnor UO_194 (O_194,N_7055,N_5914);
or UO_195 (O_195,N_9935,N_6320);
or UO_196 (O_196,N_8326,N_8712);
xor UO_197 (O_197,N_5952,N_6719);
nor UO_198 (O_198,N_6610,N_8685);
or UO_199 (O_199,N_8009,N_5785);
and UO_200 (O_200,N_9761,N_5249);
nor UO_201 (O_201,N_7128,N_5240);
nor UO_202 (O_202,N_6718,N_8734);
and UO_203 (O_203,N_6609,N_6037);
nor UO_204 (O_204,N_7227,N_5767);
xnor UO_205 (O_205,N_7287,N_6179);
or UO_206 (O_206,N_6337,N_5857);
or UO_207 (O_207,N_7086,N_6023);
nand UO_208 (O_208,N_9776,N_8451);
and UO_209 (O_209,N_9049,N_8332);
or UO_210 (O_210,N_5673,N_9221);
and UO_211 (O_211,N_8569,N_9343);
nor UO_212 (O_212,N_5453,N_6035);
xnor UO_213 (O_213,N_6750,N_7015);
xnor UO_214 (O_214,N_9642,N_8143);
nand UO_215 (O_215,N_8190,N_8883);
and UO_216 (O_216,N_6724,N_9448);
xor UO_217 (O_217,N_5899,N_6974);
or UO_218 (O_218,N_7873,N_5596);
or UO_219 (O_219,N_7897,N_5566);
or UO_220 (O_220,N_6129,N_5143);
nand UO_221 (O_221,N_7406,N_9481);
nor UO_222 (O_222,N_9766,N_9241);
and UO_223 (O_223,N_9044,N_9159);
xnor UO_224 (O_224,N_7775,N_8045);
and UO_225 (O_225,N_8296,N_9602);
nor UO_226 (O_226,N_9400,N_6396);
nand UO_227 (O_227,N_5214,N_5729);
nand UO_228 (O_228,N_9502,N_9672);
and UO_229 (O_229,N_7882,N_9864);
nor UO_230 (O_230,N_8089,N_6428);
nand UO_231 (O_231,N_6066,N_5902);
xor UO_232 (O_232,N_6602,N_5187);
or UO_233 (O_233,N_5228,N_7043);
or UO_234 (O_234,N_7459,N_7688);
or UO_235 (O_235,N_5845,N_9863);
and UO_236 (O_236,N_9970,N_7545);
and UO_237 (O_237,N_9212,N_8118);
nand UO_238 (O_238,N_9639,N_7832);
or UO_239 (O_239,N_7760,N_6222);
nand UO_240 (O_240,N_6794,N_8006);
and UO_241 (O_241,N_8583,N_7638);
nand UO_242 (O_242,N_7855,N_6189);
or UO_243 (O_243,N_6812,N_6850);
nor UO_244 (O_244,N_8138,N_9540);
xor UO_245 (O_245,N_9914,N_7598);
xor UO_246 (O_246,N_8498,N_7010);
nand UO_247 (O_247,N_9512,N_5248);
or UO_248 (O_248,N_9413,N_9484);
and UO_249 (O_249,N_9541,N_6315);
nand UO_250 (O_250,N_6230,N_7900);
nand UO_251 (O_251,N_8824,N_5513);
and UO_252 (O_252,N_9490,N_9432);
xnor UO_253 (O_253,N_8671,N_9194);
or UO_254 (O_254,N_7801,N_6625);
or UO_255 (O_255,N_5405,N_7386);
nand UO_256 (O_256,N_5410,N_8303);
xnor UO_257 (O_257,N_5066,N_7236);
nor UO_258 (O_258,N_9560,N_6613);
and UO_259 (O_259,N_9164,N_5690);
or UO_260 (O_260,N_7838,N_8749);
xnor UO_261 (O_261,N_6910,N_7836);
nor UO_262 (O_262,N_9292,N_7932);
xor UO_263 (O_263,N_6713,N_8490);
nand UO_264 (O_264,N_9141,N_6464);
xor UO_265 (O_265,N_9758,N_9147);
xor UO_266 (O_266,N_9984,N_8182);
nand UO_267 (O_267,N_7405,N_8027);
nor UO_268 (O_268,N_9173,N_7291);
nor UO_269 (O_269,N_8485,N_9489);
or UO_270 (O_270,N_7988,N_9067);
nor UO_271 (O_271,N_9037,N_8613);
or UO_272 (O_272,N_7197,N_5049);
xor UO_273 (O_273,N_5576,N_9529);
nor UO_274 (O_274,N_9438,N_6616);
nor UO_275 (O_275,N_9408,N_6962);
nand UO_276 (O_276,N_7350,N_5869);
xor UO_277 (O_277,N_6976,N_6918);
xor UO_278 (O_278,N_6745,N_7857);
or UO_279 (O_279,N_7069,N_8031);
xnor UO_280 (O_280,N_8756,N_6543);
and UO_281 (O_281,N_5872,N_5186);
nor UO_282 (O_282,N_9789,N_9574);
and UO_283 (O_283,N_6509,N_5980);
or UO_284 (O_284,N_8227,N_6270);
nand UO_285 (O_285,N_8297,N_6755);
nor UO_286 (O_286,N_5580,N_6999);
nor UO_287 (O_287,N_9128,N_5718);
xor UO_288 (O_288,N_5866,N_6537);
and UO_289 (O_289,N_8928,N_9728);
and UO_290 (O_290,N_6758,N_8410);
nand UO_291 (O_291,N_9877,N_6679);
or UO_292 (O_292,N_9772,N_7035);
nor UO_293 (O_293,N_9149,N_6211);
xor UO_294 (O_294,N_5422,N_9278);
and UO_295 (O_295,N_8916,N_8710);
xnor UO_296 (O_296,N_9978,N_8993);
and UO_297 (O_297,N_7439,N_7140);
xor UO_298 (O_298,N_6043,N_6734);
nand UO_299 (O_299,N_5723,N_5080);
nand UO_300 (O_300,N_9708,N_7432);
nand UO_301 (O_301,N_6430,N_9154);
nor UO_302 (O_302,N_6942,N_5151);
nor UO_303 (O_303,N_7952,N_9028);
and UO_304 (O_304,N_6289,N_8213);
nand UO_305 (O_305,N_8959,N_8777);
nand UO_306 (O_306,N_5023,N_7318);
nand UO_307 (O_307,N_8474,N_5056);
or UO_308 (O_308,N_9082,N_6504);
and UO_309 (O_309,N_7328,N_9267);
xor UO_310 (O_310,N_5033,N_8688);
nor UO_311 (O_311,N_6628,N_7327);
nor UO_312 (O_312,N_8203,N_8692);
nor UO_313 (O_313,N_6423,N_6950);
nor UO_314 (O_314,N_5759,N_5116);
and UO_315 (O_315,N_8572,N_6013);
xnor UO_316 (O_316,N_9171,N_8461);
nor UO_317 (O_317,N_9925,N_7215);
and UO_318 (O_318,N_5258,N_7799);
nand UO_319 (O_319,N_5884,N_8626);
nand UO_320 (O_320,N_8874,N_7121);
and UO_321 (O_321,N_8652,N_7007);
xor UO_322 (O_322,N_6303,N_5775);
nor UO_323 (O_323,N_7168,N_7819);
nor UO_324 (O_324,N_7163,N_7127);
nand UO_325 (O_325,N_5915,N_6547);
and UO_326 (O_326,N_9996,N_8908);
xor UO_327 (O_327,N_8374,N_6882);
nand UO_328 (O_328,N_6163,N_7936);
nand UO_329 (O_329,N_5064,N_7136);
nor UO_330 (O_330,N_8604,N_7961);
and UO_331 (O_331,N_8432,N_7391);
nand UO_332 (O_332,N_8047,N_9365);
nand UO_333 (O_333,N_6898,N_6112);
xnor UO_334 (O_334,N_8996,N_6887);
xnor UO_335 (O_335,N_9165,N_8519);
nand UO_336 (O_336,N_7476,N_5782);
or UO_337 (O_337,N_5578,N_7942);
nand UO_338 (O_338,N_9903,N_6238);
or UO_339 (O_339,N_7431,N_5111);
and UO_340 (O_340,N_7884,N_5179);
nor UO_341 (O_341,N_6197,N_7627);
xor UO_342 (O_342,N_6274,N_8442);
nor UO_343 (O_343,N_9785,N_8686);
nor UO_344 (O_344,N_7747,N_6229);
xor UO_345 (O_345,N_8536,N_7528);
and UO_346 (O_346,N_7321,N_5965);
nand UO_347 (O_347,N_8393,N_5392);
xor UO_348 (O_348,N_9485,N_6273);
xor UO_349 (O_349,N_7861,N_6568);
xor UO_350 (O_350,N_6627,N_6341);
xnor UO_351 (O_351,N_8029,N_9850);
nand UO_352 (O_352,N_8880,N_9372);
nand UO_353 (O_353,N_6422,N_6975);
and UO_354 (O_354,N_6934,N_7740);
nor UO_355 (O_355,N_9665,N_9072);
xnor UO_356 (O_356,N_7143,N_9523);
nor UO_357 (O_357,N_9973,N_8935);
nor UO_358 (O_358,N_7453,N_8917);
nand UO_359 (O_359,N_9715,N_8102);
and UO_360 (O_360,N_9569,N_7360);
or UO_361 (O_361,N_7173,N_6075);
xnor UO_362 (O_362,N_5812,N_9098);
nand UO_363 (O_363,N_8049,N_6003);
nand UO_364 (O_364,N_8655,N_9423);
or UO_365 (O_365,N_7814,N_5140);
nor UO_366 (O_366,N_9445,N_5098);
or UO_367 (O_367,N_5917,N_7870);
nor UO_368 (O_368,N_8921,N_8482);
xnor UO_369 (O_369,N_6301,N_6902);
xnor UO_370 (O_370,N_5887,N_6822);
and UO_371 (O_371,N_7896,N_5259);
nand UO_372 (O_372,N_9493,N_7647);
nand UO_373 (O_373,N_5890,N_7040);
xor UO_374 (O_374,N_9064,N_9909);
or UO_375 (O_375,N_9999,N_9704);
xor UO_376 (O_376,N_9910,N_6829);
xor UO_377 (O_377,N_9500,N_5435);
xor UO_378 (O_378,N_5743,N_9094);
or UO_379 (O_379,N_7385,N_6477);
nand UO_380 (O_380,N_5694,N_6626);
nand UO_381 (O_381,N_8913,N_7196);
xor UO_382 (O_382,N_6840,N_7254);
nand UO_383 (O_383,N_5896,N_6967);
nor UO_384 (O_384,N_6440,N_8195);
and UO_385 (O_385,N_7858,N_8079);
or UO_386 (O_386,N_5642,N_6118);
nor UO_387 (O_387,N_5326,N_6842);
nand UO_388 (O_388,N_6082,N_7072);
nor UO_389 (O_389,N_7309,N_8473);
xnor UO_390 (O_390,N_9146,N_6703);
nand UO_391 (O_391,N_6095,N_8156);
nand UO_392 (O_392,N_7094,N_7667);
and UO_393 (O_393,N_8795,N_7824);
or UO_394 (O_394,N_7306,N_5173);
nand UO_395 (O_395,N_9768,N_7518);
or UO_396 (O_396,N_9979,N_5479);
and UO_397 (O_397,N_9664,N_7576);
nand UO_398 (O_398,N_9418,N_9380);
xnor UO_399 (O_399,N_9056,N_9427);
and UO_400 (O_400,N_6954,N_5395);
and UO_401 (O_401,N_8405,N_6058);
xnor UO_402 (O_402,N_6473,N_5559);
nand UO_403 (O_403,N_7117,N_9721);
or UO_404 (O_404,N_8236,N_8775);
nor UO_405 (O_405,N_5029,N_5044);
nor UO_406 (O_406,N_8460,N_6601);
and UO_407 (O_407,N_5152,N_9652);
and UO_408 (O_408,N_5356,N_6108);
and UO_409 (O_409,N_9223,N_9457);
nor UO_410 (O_410,N_6545,N_9383);
or UO_411 (O_411,N_5651,N_9020);
xor UO_412 (O_412,N_5784,N_9114);
nor UO_413 (O_413,N_8371,N_5606);
xnor UO_414 (O_414,N_6991,N_6973);
nor UO_415 (O_415,N_7050,N_6825);
nand UO_416 (O_416,N_6087,N_7125);
nor UO_417 (O_417,N_6529,N_8875);
or UO_418 (O_418,N_7005,N_5082);
nand UO_419 (O_419,N_9568,N_9566);
or UO_420 (O_420,N_7694,N_5715);
xnor UO_421 (O_421,N_7455,N_5280);
nand UO_422 (O_422,N_7120,N_7076);
and UO_423 (O_423,N_7770,N_5437);
xor UO_424 (O_424,N_8501,N_9335);
nor UO_425 (O_425,N_9022,N_5878);
xnor UO_426 (O_426,N_8620,N_6357);
nor UO_427 (O_427,N_8649,N_8202);
or UO_428 (O_428,N_7728,N_8055);
xnor UO_429 (O_429,N_5454,N_6698);
nor UO_430 (O_430,N_5190,N_6907);
or UO_431 (O_431,N_8937,N_7395);
nor UO_432 (O_432,N_6978,N_5786);
and UO_433 (O_433,N_8252,N_9968);
xor UO_434 (O_434,N_8169,N_7452);
nand UO_435 (O_435,N_8838,N_8131);
nand UO_436 (O_436,N_7886,N_8180);
nand UO_437 (O_437,N_8741,N_6002);
nand UO_438 (O_438,N_5084,N_7892);
xor UO_439 (O_439,N_8826,N_6528);
nor UO_440 (O_440,N_5145,N_8951);
and UO_441 (O_441,N_5208,N_9473);
nand UO_442 (O_442,N_6804,N_5724);
nand UO_443 (O_443,N_8633,N_6193);
nor UO_444 (O_444,N_9831,N_7088);
xnor UO_445 (O_445,N_5030,N_8310);
nand UO_446 (O_446,N_9990,N_5432);
or UO_447 (O_447,N_7314,N_8813);
nand UO_448 (O_448,N_8758,N_7421);
nand UO_449 (O_449,N_7145,N_7135);
nand UO_450 (O_450,N_9921,N_6982);
or UO_451 (O_451,N_5747,N_6295);
or UO_452 (O_452,N_7623,N_9498);
nor UO_453 (O_453,N_9178,N_6096);
or UO_454 (O_454,N_7243,N_7658);
or UO_455 (O_455,N_8043,N_7639);
nand UO_456 (O_456,N_5458,N_5716);
nor UO_457 (O_457,N_8974,N_9603);
and UO_458 (O_458,N_8506,N_8287);
and UO_459 (O_459,N_8262,N_9750);
or UO_460 (O_460,N_7987,N_9076);
nor UO_461 (O_461,N_6122,N_6711);
xor UO_462 (O_462,N_5947,N_7671);
and UO_463 (O_463,N_7975,N_5442);
nand UO_464 (O_464,N_7901,N_6873);
nor UO_465 (O_465,N_5590,N_6228);
xor UO_466 (O_466,N_7019,N_5081);
and UO_467 (O_467,N_8525,N_9174);
nor UO_468 (O_468,N_6500,N_6117);
nand UO_469 (O_469,N_7918,N_5731);
and UO_470 (O_470,N_9288,N_6877);
xor UO_471 (O_471,N_5062,N_7684);
or UO_472 (O_472,N_8730,N_9840);
or UO_473 (O_473,N_5996,N_5412);
nand UO_474 (O_474,N_9204,N_9196);
or UO_475 (O_475,N_8503,N_6809);
and UO_476 (O_476,N_5698,N_7536);
and UO_477 (O_477,N_7293,N_9373);
and UO_478 (O_478,N_6686,N_5079);
nand UO_479 (O_479,N_6218,N_6009);
nand UO_480 (O_480,N_6624,N_6605);
nand UO_481 (O_481,N_5888,N_8956);
nand UO_482 (O_482,N_6150,N_5512);
and UO_483 (O_483,N_6544,N_8484);
xor UO_484 (O_484,N_6125,N_6821);
nor UO_485 (O_485,N_8380,N_8782);
xor UO_486 (O_486,N_5177,N_5807);
or UO_487 (O_487,N_9801,N_7940);
xor UO_488 (O_488,N_9272,N_6385);
nand UO_489 (O_489,N_7027,N_8034);
nand UO_490 (O_490,N_6623,N_6284);
and UO_491 (O_491,N_6891,N_8235);
nor UO_492 (O_492,N_5371,N_9324);
and UO_493 (O_493,N_9730,N_7966);
and UO_494 (O_494,N_6046,N_8205);
nor UO_495 (O_495,N_5882,N_9788);
and UO_496 (O_496,N_9406,N_5440);
xnor UO_497 (O_497,N_6330,N_8641);
and UO_498 (O_498,N_9045,N_7351);
nor UO_499 (O_499,N_9062,N_9533);
or UO_500 (O_500,N_9366,N_9825);
xnor UO_501 (O_501,N_8631,N_6685);
and UO_502 (O_502,N_6501,N_5313);
or UO_503 (O_503,N_7634,N_5357);
nand UO_504 (O_504,N_5288,N_8140);
xnor UO_505 (O_505,N_5071,N_8897);
xnor UO_506 (O_506,N_9993,N_9934);
or UO_507 (O_507,N_7885,N_8934);
nand UO_508 (O_508,N_8919,N_7198);
nand UO_509 (O_509,N_5672,N_5522);
or UO_510 (O_510,N_9882,N_6903);
or UO_511 (O_511,N_5095,N_6045);
and UO_512 (O_512,N_7464,N_5533);
xnor UO_513 (O_513,N_5157,N_5263);
and UO_514 (O_514,N_7376,N_9251);
and UO_515 (O_515,N_6068,N_8735);
or UO_516 (O_516,N_8007,N_9501);
and UO_517 (O_517,N_7369,N_6785);
xnor UO_518 (O_518,N_8636,N_9567);
nor UO_519 (O_519,N_9479,N_5841);
nand UO_520 (O_520,N_9249,N_5264);
nor UO_521 (O_521,N_7472,N_5393);
xor UO_522 (O_522,N_9644,N_7874);
and UO_523 (O_523,N_8612,N_7842);
or UO_524 (O_524,N_6442,N_8896);
nor UO_525 (O_525,N_7971,N_5577);
and UO_526 (O_526,N_7899,N_7250);
and UO_527 (O_527,N_9939,N_9807);
or UO_528 (O_528,N_5662,N_6278);
nand UO_529 (O_529,N_8074,N_6344);
or UO_530 (O_530,N_8793,N_8607);
or UO_531 (O_531,N_9332,N_9111);
or UO_532 (O_532,N_8809,N_7588);
xnor UO_533 (O_533,N_8172,N_9245);
or UO_534 (O_534,N_5871,N_9311);
xor UO_535 (O_535,N_8721,N_9217);
and UO_536 (O_536,N_9464,N_8517);
or UO_537 (O_537,N_5670,N_6774);
nand UO_538 (O_538,N_8136,N_6674);
nand UO_539 (O_539,N_8232,N_9966);
nor UO_540 (O_540,N_9455,N_5203);
xnor UO_541 (O_541,N_5620,N_7501);
or UO_542 (O_542,N_8269,N_6817);
and UO_543 (O_543,N_5230,N_5873);
xor UO_544 (O_544,N_6611,N_9558);
nand UO_545 (O_545,N_7651,N_7630);
and UO_546 (O_546,N_6447,N_8130);
nand UO_547 (O_547,N_9956,N_5068);
nand UO_548 (O_548,N_5282,N_9815);
nand UO_549 (O_549,N_7514,N_9591);
nor UO_550 (O_550,N_9270,N_6579);
and UO_551 (O_551,N_8362,N_6170);
and UO_552 (O_552,N_7789,N_7304);
or UO_553 (O_553,N_7396,N_9549);
and UO_554 (O_554,N_8595,N_6445);
xnor UO_555 (O_555,N_7813,N_6818);
xor UO_556 (O_556,N_7786,N_8038);
and UO_557 (O_557,N_5261,N_6223);
and UO_558 (O_558,N_6062,N_8126);
nor UO_559 (O_559,N_9525,N_6772);
xor UO_560 (O_560,N_7904,N_9576);
xor UO_561 (O_561,N_5605,N_7000);
or UO_562 (O_562,N_6361,N_5754);
or UO_563 (O_563,N_9359,N_6349);
or UO_564 (O_564,N_5949,N_9135);
and UO_565 (O_565,N_5726,N_6557);
nor UO_566 (O_566,N_5701,N_8906);
xor UO_567 (O_567,N_5564,N_5827);
xor UO_568 (O_568,N_5556,N_9688);
xnor UO_569 (O_569,N_8228,N_9961);
or UO_570 (O_570,N_7551,N_6692);
nand UO_571 (O_571,N_9618,N_8958);
and UO_572 (O_572,N_9797,N_5735);
xor UO_573 (O_573,N_9286,N_6497);
nand UO_574 (O_574,N_8559,N_6525);
or UO_575 (O_575,N_6241,N_8707);
or UO_576 (O_576,N_7850,N_6752);
and UO_577 (O_577,N_7363,N_6144);
xor UO_578 (O_578,N_9729,N_6526);
and UO_579 (O_579,N_8728,N_8222);
and UO_580 (O_580,N_6345,N_5296);
nor UO_581 (O_581,N_8576,N_7211);
xnor UO_582 (O_582,N_5148,N_7488);
and UO_583 (O_583,N_8458,N_9648);
and UO_584 (O_584,N_8962,N_6959);
and UO_585 (O_585,N_9087,N_6370);
or UO_586 (O_586,N_7696,N_7621);
xnor UO_587 (O_587,N_9632,N_7149);
or UO_588 (O_588,N_5600,N_6846);
nand UO_589 (O_589,N_5994,N_8165);
or UO_590 (O_590,N_6845,N_5147);
and UO_591 (O_591,N_9946,N_7008);
or UO_592 (O_592,N_5094,N_6749);
nand UO_593 (O_593,N_7974,N_7967);
nand UO_594 (O_594,N_7510,N_6268);
and UO_595 (O_595,N_6049,N_5199);
or UO_596 (O_596,N_9279,N_7982);
nor UO_597 (O_597,N_5746,N_9330);
and UO_598 (O_598,N_8321,N_5273);
xnor UO_599 (O_599,N_6830,N_9875);
nor UO_600 (O_600,N_5534,N_7563);
or UO_601 (O_601,N_5427,N_6468);
xnor UO_602 (O_602,N_7584,N_8859);
nor UO_603 (O_603,N_7123,N_6741);
xor UO_604 (O_604,N_8349,N_8492);
nor UO_605 (O_605,N_9816,N_9200);
and UO_606 (O_606,N_7565,N_5835);
and UO_607 (O_607,N_8949,N_6498);
or UO_608 (O_608,N_9017,N_6542);
xnor UO_609 (O_609,N_6941,N_8968);
nor UO_610 (O_610,N_5836,N_8806);
nand UO_611 (O_611,N_8783,N_6051);
and UO_612 (O_612,N_9152,N_7161);
nor UO_613 (O_613,N_5146,N_6870);
nor UO_614 (O_614,N_7257,N_9220);
nand UO_615 (O_615,N_7482,N_6022);
nor UO_616 (O_616,N_9697,N_8681);
xor UO_617 (O_617,N_8283,N_7133);
or UO_618 (O_618,N_7275,N_7980);
and UO_619 (O_619,N_6260,N_5290);
or UO_620 (O_620,N_9183,N_8886);
xnor UO_621 (O_621,N_7233,N_8719);
or UO_622 (O_622,N_9412,N_9170);
nand UO_623 (O_623,N_5369,N_7959);
xor UO_624 (O_624,N_6715,N_5631);
xor UO_625 (O_625,N_8954,N_7049);
xor UO_626 (O_626,N_5722,N_8960);
or UO_627 (O_627,N_6282,N_9471);
xor UO_628 (O_628,N_5163,N_6788);
xnor UO_629 (O_629,N_6584,N_6433);
xor UO_630 (O_630,N_5535,N_9703);
and UO_631 (O_631,N_7447,N_5406);
xnor UO_632 (O_632,N_6663,N_5621);
nand UO_633 (O_633,N_6486,N_5128);
or UO_634 (O_634,N_6010,N_5430);
nand UO_635 (O_635,N_8259,N_9983);
nand UO_636 (O_636,N_5034,N_6816);
or UO_637 (O_637,N_9954,N_9578);
nand UO_638 (O_638,N_8611,N_7478);
xnor UO_639 (O_639,N_8925,N_7506);
and UO_640 (O_640,N_6219,N_8737);
or UO_641 (O_641,N_7910,N_9444);
and UO_642 (O_642,N_5636,N_6376);
nor UO_643 (O_643,N_9692,N_9316);
nand UO_644 (O_644,N_6177,N_5960);
nor UO_645 (O_645,N_5588,N_7852);
nor UO_646 (O_646,N_8115,N_7751);
and UO_647 (O_647,N_9469,N_5849);
or UO_648 (O_648,N_6864,N_8625);
and UO_649 (O_649,N_6637,N_8738);
and UO_650 (O_650,N_9377,N_5420);
or UO_651 (O_651,N_5039,N_5740);
nor UO_652 (O_652,N_8575,N_7869);
nor UO_653 (O_653,N_7677,N_7633);
nand UO_654 (O_654,N_5652,N_6064);
and UO_655 (O_655,N_8470,N_5061);
and UO_656 (O_656,N_9867,N_9517);
nor UO_657 (O_657,N_9941,N_8308);
xnor UO_658 (O_658,N_8947,N_6596);
xor UO_659 (O_659,N_6981,N_7349);
or UO_660 (O_660,N_5550,N_5548);
xnor UO_661 (O_661,N_9050,N_8185);
xor UO_662 (O_662,N_8900,N_6480);
nand UO_663 (O_663,N_6514,N_5031);
nor UO_664 (O_664,N_8051,N_6591);
or UO_665 (O_665,N_9771,N_9254);
nand UO_666 (O_666,N_5507,N_5883);
nor UO_667 (O_667,N_8555,N_6588);
nor UO_668 (O_668,N_7654,N_5668);
and UO_669 (O_669,N_7147,N_9869);
and UO_670 (O_670,N_7611,N_6929);
or UO_671 (O_671,N_8431,N_8342);
nand UO_672 (O_672,N_9250,N_5946);
nand UO_673 (O_673,N_5851,N_6805);
and UO_674 (O_674,N_8486,N_9792);
xnor UO_675 (O_675,N_6576,N_5579);
nor UO_676 (O_676,N_7829,N_9389);
and UO_677 (O_677,N_7955,N_5531);
nor UO_678 (O_678,N_7618,N_5455);
or UO_679 (O_679,N_5697,N_6930);
and UO_680 (O_680,N_5934,N_9218);
nor UO_681 (O_681,N_9429,N_5922);
nor UO_682 (O_682,N_6323,N_5657);
nand UO_683 (O_683,N_8359,N_8560);
nor UO_684 (O_684,N_5252,N_9519);
nand UO_685 (O_685,N_9700,N_8706);
or UO_686 (O_686,N_5101,N_8003);
nand UO_687 (O_687,N_5532,N_6810);
or UO_688 (O_688,N_9731,N_8520);
xnor UO_689 (O_689,N_5345,N_5175);
nor UO_690 (O_690,N_7175,N_7712);
and UO_691 (O_691,N_8441,N_5615);
nor UO_692 (O_692,N_5639,N_5373);
nor UO_693 (O_693,N_9496,N_9962);
and UO_694 (O_694,N_8463,N_6266);
or UO_695 (O_695,N_8682,N_8950);
nor UO_696 (O_696,N_9738,N_6660);
nor UO_697 (O_697,N_7527,N_6297);
or UO_698 (O_698,N_8373,N_6018);
xnor UO_699 (O_699,N_6174,N_5342);
or UO_700 (O_700,N_5492,N_8725);
xnor UO_701 (O_701,N_6054,N_8895);
and UO_702 (O_702,N_8116,N_8035);
and UO_703 (O_703,N_8466,N_5854);
and UO_704 (O_704,N_6495,N_8112);
nor UO_705 (O_705,N_8573,N_9861);
xor UO_706 (O_706,N_5977,N_9387);
nand UO_707 (O_707,N_6387,N_5962);
xnor UO_708 (O_708,N_5063,N_5942);
nor UO_709 (O_709,N_5761,N_9156);
or UO_710 (O_710,N_6048,N_8266);
xnor UO_711 (O_711,N_9963,N_7756);
and UO_712 (O_712,N_8013,N_9179);
nor UO_713 (O_713,N_8016,N_8124);
and UO_714 (O_714,N_7944,N_7134);
and UO_715 (O_715,N_9587,N_9522);
and UO_716 (O_716,N_9830,N_7104);
nor UO_717 (O_717,N_7382,N_5226);
nor UO_718 (O_718,N_8137,N_5680);
and UO_719 (O_719,N_8512,N_6173);
xnor UO_720 (O_720,N_5285,N_9845);
and UO_721 (O_721,N_7438,N_7708);
nand UO_722 (O_722,N_6493,N_5311);
xnor UO_723 (O_723,N_7581,N_6308);
and UO_724 (O_724,N_8300,N_5546);
xor UO_725 (O_725,N_8459,N_9090);
or UO_726 (O_726,N_6876,N_7262);
xor UO_727 (O_727,N_9612,N_6164);
or UO_728 (O_728,N_7157,N_7782);
xnor UO_729 (O_729,N_5591,N_9066);
or UO_730 (O_730,N_7182,N_5439);
or UO_731 (O_731,N_6599,N_7172);
nand UO_732 (O_732,N_6232,N_9209);
nor UO_733 (O_733,N_7091,N_7399);
and UO_734 (O_734,N_9685,N_7378);
nor UO_735 (O_735,N_8256,N_9215);
or UO_736 (O_736,N_6866,N_9403);
and UO_737 (O_737,N_7672,N_8769);
and UO_738 (O_738,N_5727,N_5232);
or UO_739 (O_739,N_5172,N_6714);
nand UO_740 (O_740,N_8639,N_8480);
and UO_741 (O_741,N_8690,N_6587);
nand UO_742 (O_742,N_6031,N_8122);
and UO_743 (O_743,N_5554,N_5004);
nor UO_744 (O_744,N_5843,N_9548);
or UO_745 (O_745,N_8408,N_9838);
or UO_746 (O_746,N_6209,N_5763);
xor UO_747 (O_747,N_8450,N_8098);
or UO_748 (O_748,N_6757,N_9734);
nand UO_749 (O_749,N_9253,N_7348);
nand UO_750 (O_750,N_6516,N_7114);
xor UO_751 (O_751,N_8606,N_9951);
nor UO_752 (O_752,N_9441,N_6566);
and UO_753 (O_753,N_6032,N_7895);
xnor UO_754 (O_754,N_9782,N_5462);
and UO_755 (O_755,N_8829,N_6253);
or UO_756 (O_756,N_8018,N_7951);
and UO_757 (O_757,N_8714,N_7225);
nand UO_758 (O_758,N_7548,N_5195);
xor UO_759 (O_759,N_6204,N_9113);
nand UO_760 (O_760,N_7597,N_8586);
nor UO_761 (O_761,N_9381,N_6518);
xnor UO_762 (O_762,N_6868,N_8680);
nor UO_763 (O_763,N_8892,N_5414);
xor UO_764 (O_764,N_6489,N_8872);
and UO_765 (O_765,N_9079,N_6699);
and UO_766 (O_766,N_8123,N_6178);
nand UO_767 (O_767,N_8274,N_9778);
xor UO_768 (O_768,N_8363,N_6970);
nand UO_769 (O_769,N_7193,N_9495);
or UO_770 (O_770,N_7346,N_8711);
xnor UO_771 (O_771,N_7788,N_9551);
or UO_772 (O_772,N_9280,N_7887);
nor UO_773 (O_773,N_6502,N_8537);
or UO_774 (O_774,N_7129,N_8096);
or UO_775 (O_775,N_6662,N_6796);
nor UO_776 (O_776,N_7500,N_9107);
or UO_777 (O_777,N_9105,N_6036);
or UO_778 (O_778,N_8691,N_5159);
or UO_779 (O_779,N_7643,N_6952);
nor UO_780 (O_780,N_6214,N_8200);
and UO_781 (O_781,N_8421,N_9084);
and UO_782 (O_782,N_5856,N_8505);
xnor UO_783 (O_783,N_8870,N_5863);
nor UO_784 (O_784,N_6334,N_6324);
xnor UO_785 (O_785,N_6524,N_7484);
or UO_786 (O_786,N_6553,N_9296);
and UO_787 (O_787,N_6721,N_5091);
nand UO_788 (O_788,N_8781,N_9130);
nand UO_789 (O_789,N_8709,N_5013);
or UO_790 (O_790,N_5976,N_9458);
and UO_791 (O_791,N_9362,N_9391);
nand UO_792 (O_792,N_6059,N_7542);
nand UO_793 (O_793,N_8871,N_8197);
and UO_794 (O_794,N_7946,N_6254);
nor UO_795 (O_795,N_7994,N_6299);
nand UO_796 (O_796,N_8286,N_8419);
or UO_797 (O_797,N_8898,N_5207);
and UO_798 (O_798,N_9808,N_9952);
nor UO_799 (O_799,N_8876,N_6647);
nor UO_800 (O_800,N_8497,N_6862);
xor UO_801 (O_801,N_9503,N_7992);
nor UO_802 (O_802,N_5867,N_9309);
nand UO_803 (O_803,N_8703,N_9922);
xnor UO_804 (O_804,N_6808,N_8301);
xnor UO_805 (O_805,N_6482,N_7358);
nand UO_806 (O_806,N_6635,N_7798);
nand UO_807 (O_807,N_6316,N_9720);
and UO_808 (O_808,N_7958,N_7075);
and UO_809 (O_809,N_8028,N_5346);
or UO_810 (O_810,N_7344,N_7840);
and UO_811 (O_811,N_7710,N_5466);
xnor UO_812 (O_812,N_9228,N_5211);
or UO_813 (O_813,N_9176,N_7084);
xnor UO_814 (O_814,N_5234,N_6380);
nand UO_815 (O_815,N_6964,N_9442);
and UO_816 (O_816,N_5710,N_6681);
and UO_817 (O_817,N_7435,N_8263);
xnor UO_818 (O_818,N_7158,N_5574);
nor UO_819 (O_819,N_6104,N_8981);
xnor UO_820 (O_820,N_7758,N_7030);
or UO_821 (O_821,N_5622,N_8391);
or UO_822 (O_822,N_5999,N_5779);
nand UO_823 (O_823,N_7912,N_8247);
nand UO_824 (O_824,N_7445,N_5028);
nor UO_825 (O_825,N_9832,N_6764);
nor UO_826 (O_826,N_7515,N_9086);
xor UO_827 (O_827,N_8146,N_8836);
nor UO_828 (O_828,N_8722,N_8155);
nand UO_829 (O_829,N_6583,N_9282);
xnor UO_830 (O_830,N_8386,N_6894);
nor UO_831 (O_831,N_7156,N_6879);
or UO_832 (O_832,N_8429,N_9762);
nor UO_833 (O_833,N_6298,N_8376);
xnor UO_834 (O_834,N_9338,N_9866);
or UO_835 (O_835,N_5798,N_9475);
xor UO_836 (O_836,N_6782,N_7064);
nor UO_837 (O_837,N_6472,N_8254);
xnor UO_838 (O_838,N_8979,N_6065);
nor UO_839 (O_839,N_7244,N_7575);
nor UO_840 (O_840,N_8179,N_7646);
nand UO_841 (O_841,N_7953,N_5428);
and UO_842 (O_842,N_6759,N_6522);
or UO_843 (O_843,N_6074,N_5774);
or UO_844 (O_844,N_7707,N_5155);
nand UO_845 (O_845,N_8799,N_5005);
and UO_846 (O_846,N_7345,N_6670);
nor UO_847 (O_847,N_6530,N_7815);
nor UO_848 (O_848,N_8329,N_7720);
nand UO_849 (O_849,N_9155,N_8430);
nor UO_850 (O_850,N_5090,N_5341);
xnor UO_851 (O_851,N_9166,N_8475);
nor UO_852 (O_852,N_6748,N_6598);
nor UO_853 (O_853,N_6827,N_8658);
and UO_854 (O_854,N_9819,N_6172);
nor UO_855 (O_855,N_6304,N_5687);
xnor UO_856 (O_856,N_5219,N_8787);
or UO_857 (O_857,N_8319,N_9198);
nand UO_858 (O_858,N_5021,N_8825);
or UO_859 (O_859,N_5932,N_7433);
nor UO_860 (O_860,N_9264,N_6927);
nor UO_861 (O_861,N_9593,N_6696);
xor UO_862 (O_862,N_6459,N_5274);
nand UO_863 (O_863,N_6184,N_8784);
and UO_864 (O_864,N_9110,N_8933);
or UO_865 (O_865,N_7190,N_9744);
xnor UO_866 (O_866,N_7152,N_5483);
nor UO_867 (O_867,N_5702,N_9417);
xnor UO_868 (O_868,N_6837,N_8181);
or UO_869 (O_869,N_7839,N_8718);
nor UO_870 (O_870,N_7499,N_8157);
xor UO_871 (O_871,N_5645,N_5407);
and UO_872 (O_872,N_9449,N_8600);
nor UO_873 (O_873,N_9197,N_9129);
nand UO_874 (O_874,N_8659,N_8675);
and UO_875 (O_875,N_8417,N_7343);
or UO_876 (O_876,N_5139,N_6763);
xnor UO_877 (O_877,N_9786,N_8891);
or UO_878 (O_878,N_7373,N_9942);
xnor UO_879 (O_879,N_6034,N_9912);
and UO_880 (O_880,N_5618,N_8548);
and UO_881 (O_881,N_6457,N_8522);
xnor UO_882 (O_882,N_5665,N_9276);
xnor UO_883 (O_883,N_9012,N_5328);
nand UO_884 (O_884,N_7100,N_7725);
nand UO_885 (O_885,N_7112,N_7554);
or UO_886 (O_886,N_5286,N_6487);
nand UO_887 (O_887,N_5174,N_6552);
nand UO_888 (O_888,N_9821,N_9880);
and UO_889 (O_889,N_6649,N_5354);
and UO_890 (O_890,N_5676,N_9315);
nor UO_891 (O_891,N_8945,N_8663);
and UO_892 (O_892,N_6727,N_8381);
or UO_893 (O_893,N_6786,N_5637);
nor UO_894 (O_894,N_5225,N_7251);
nor UO_895 (O_895,N_7281,N_7042);
nor UO_896 (O_896,N_6141,N_5347);
and UO_897 (O_897,N_6107,N_9902);
nor UO_898 (O_898,N_7490,N_7074);
nor UO_899 (O_899,N_5376,N_7902);
nor UO_900 (O_900,N_5099,N_9599);
nand UO_901 (O_901,N_6622,N_5144);
nor UO_902 (O_902,N_7741,N_9702);
and UO_903 (O_903,N_6367,N_5123);
nand UO_904 (O_904,N_9755,N_7656);
nand UO_905 (O_905,N_7415,N_7505);
and UO_906 (O_906,N_5719,N_5164);
nand UO_907 (O_907,N_6886,N_8848);
or UO_908 (O_908,N_7341,N_7790);
xor UO_909 (O_909,N_6678,N_8343);
nor UO_910 (O_910,N_6904,N_8768);
or UO_911 (O_911,N_8294,N_7241);
and UO_912 (O_912,N_7214,N_8418);
nor UO_913 (O_913,N_8842,N_9420);
and UO_914 (O_914,N_9933,N_8217);
xor UO_915 (O_915,N_5608,N_9641);
and UO_916 (O_916,N_8387,N_7167);
nor UO_917 (O_917,N_9613,N_6186);
nor UO_918 (O_918,N_6506,N_5583);
xor UO_919 (O_919,N_7248,N_7258);
nor UO_920 (O_920,N_7009,N_6185);
or UO_921 (O_921,N_9488,N_5766);
or UO_922 (O_922,N_5855,N_7166);
xnor UO_923 (O_923,N_6847,N_5923);
xor UO_924 (O_924,N_7650,N_5811);
or UO_925 (O_925,N_7785,N_8088);
nor UO_926 (O_926,N_9849,N_7847);
nor UO_927 (O_927,N_8449,N_5595);
or UO_928 (O_928,N_5364,N_5769);
and UO_929 (O_929,N_9461,N_8471);
and UO_930 (O_930,N_6535,N_7498);
and UO_931 (O_931,N_8344,N_9940);
or UO_932 (O_932,N_7649,N_6595);
nor UO_933 (O_933,N_9713,N_8533);
or UO_934 (O_934,N_8999,N_8514);
nor UO_935 (O_935,N_5183,N_8192);
and UO_936 (O_936,N_7230,N_9638);
or UO_937 (O_937,N_5224,N_5828);
nor UO_938 (O_938,N_8864,N_7039);
nand UO_939 (O_939,N_9232,N_9741);
nor UO_940 (O_940,N_6780,N_5831);
xor UO_941 (O_941,N_8189,N_5510);
or UO_942 (O_942,N_9976,N_6205);
nor UO_943 (O_943,N_9894,N_9544);
nor UO_944 (O_944,N_9765,N_6784);
xor UO_945 (O_945,N_8818,N_8502);
xor UO_946 (O_946,N_7606,N_7059);
and UO_947 (O_947,N_5300,N_6811);
nor UO_948 (O_948,N_8447,N_7486);
nand UO_949 (O_949,N_7461,N_6382);
xor UO_950 (O_950,N_7945,N_8328);
nor UO_951 (O_951,N_7404,N_8971);
xnor UO_952 (O_952,N_8943,N_8847);
nor UO_953 (O_953,N_5842,N_5243);
and UO_954 (O_954,N_7101,N_7031);
or UO_955 (O_955,N_5875,N_6201);
or UO_956 (O_956,N_8046,N_7730);
and UO_957 (O_957,N_8483,N_5728);
xnor UO_958 (O_958,N_7276,N_7146);
or UO_959 (O_959,N_6819,N_7361);
nor UO_960 (O_960,N_8977,N_6188);
and UO_961 (O_961,N_6990,N_7503);
xnor UO_962 (O_962,N_6053,N_8398);
nand UO_963 (O_963,N_5433,N_8939);
and UO_964 (O_964,N_5444,N_8589);
nor UO_965 (O_965,N_8389,N_8399);
and UO_966 (O_966,N_5526,N_9647);
and UO_967 (O_967,N_7525,N_5162);
xor UO_968 (O_968,N_5984,N_5669);
or UO_969 (O_969,N_9019,N_6366);
nor UO_970 (O_970,N_6575,N_5256);
xnor UO_971 (O_971,N_9435,N_5955);
or UO_972 (O_972,N_5379,N_6648);
or UO_973 (O_973,N_5058,N_9148);
or UO_974 (O_974,N_9809,N_5416);
xnor UO_975 (O_975,N_8992,N_8462);
xor UO_976 (O_976,N_9273,N_5974);
or UO_977 (O_977,N_8066,N_8407);
xnor UO_978 (O_978,N_7666,N_8164);
and UO_979 (O_979,N_5378,N_6165);
nor UO_980 (O_980,N_5468,N_8684);
or UO_981 (O_981,N_6688,N_8862);
xnor UO_982 (O_982,N_9924,N_5473);
xnor UO_983 (O_983,N_8909,N_8794);
or UO_984 (O_984,N_9937,N_7648);
nand UO_985 (O_985,N_6285,N_5494);
nand UO_986 (O_986,N_6806,N_8023);
or UO_987 (O_987,N_9810,N_5713);
nor UO_988 (O_988,N_7377,N_6924);
xnor UO_989 (O_989,N_8638,N_8736);
or UO_990 (O_990,N_8761,N_8656);
xnor UO_991 (O_991,N_5780,N_7914);
nor UO_992 (O_992,N_8647,N_8727);
and UO_993 (O_993,N_7277,N_6283);
nand UO_994 (O_994,N_6569,N_7762);
and UO_995 (O_995,N_9847,N_8411);
nor UO_996 (O_996,N_7070,N_8840);
xor UO_997 (O_997,N_6342,N_7733);
nand UO_998 (O_998,N_6081,N_7426);
xnor UO_999 (O_999,N_5679,N_7456);
nor UO_1000 (O_1000,N_5907,N_6379);
nor UO_1001 (O_1001,N_8879,N_7845);
and UO_1002 (O_1002,N_5671,N_7769);
and UO_1003 (O_1003,N_7460,N_5603);
nor UO_1004 (O_1004,N_5141,N_5549);
nand UO_1005 (O_1005,N_7668,N_8479);
or UO_1006 (O_1006,N_8384,N_7428);
and UO_1007 (O_1007,N_6294,N_5752);
nand UO_1008 (O_1008,N_6833,N_6923);
nor UO_1009 (O_1009,N_5868,N_6890);
and UO_1010 (O_1010,N_8545,N_5142);
xor UO_1011 (O_1011,N_7024,N_6835);
and UO_1012 (O_1012,N_7118,N_9707);
nor UO_1013 (O_1013,N_6432,N_8566);
nor UO_1014 (O_1014,N_7915,N_7972);
or UO_1015 (O_1015,N_7202,N_8289);
and UO_1016 (O_1016,N_5648,N_5528);
or UO_1017 (O_1017,N_6346,N_7817);
nor UO_1018 (O_1018,N_5751,N_7221);
nand UO_1019 (O_1019,N_9374,N_5180);
and UO_1020 (O_1020,N_6300,N_9419);
nor UO_1021 (O_1021,N_5776,N_7962);
nor UO_1022 (O_1022,N_8033,N_5787);
nor UO_1023 (O_1023,N_9483,N_7807);
xor UO_1024 (O_1024,N_9651,N_8535);
or UO_1025 (O_1025,N_7685,N_6450);
and UO_1026 (O_1026,N_9450,N_7713);
nor UO_1027 (O_1027,N_8424,N_5417);
and UO_1028 (O_1028,N_9428,N_5937);
and UO_1029 (O_1029,N_5770,N_9472);
nor UO_1030 (O_1030,N_7660,N_9575);
nor UO_1031 (O_1031,N_9136,N_6961);
nand UO_1032 (O_1032,N_5795,N_8368);
or UO_1033 (O_1033,N_9099,N_5575);
or UO_1034 (O_1034,N_9842,N_6958);
and UO_1035 (O_1035,N_7727,N_7680);
nor UO_1036 (O_1036,N_5886,N_6620);
and UO_1037 (O_1037,N_7614,N_5221);
and UO_1038 (O_1038,N_7883,N_6867);
nand UO_1039 (O_1039,N_6242,N_6897);
or UO_1040 (O_1040,N_5333,N_7586);
or UO_1041 (O_1041,N_6114,N_6488);
xor UO_1042 (O_1042,N_7116,N_5592);
or UO_1043 (O_1043,N_9231,N_9230);
and UO_1044 (O_1044,N_9186,N_6293);
xnor UO_1045 (O_1045,N_5402,N_6157);
xor UO_1046 (O_1046,N_9290,N_6928);
nand UO_1047 (O_1047,N_5921,N_9955);
xnor UO_1048 (O_1048,N_8998,N_9006);
or UO_1049 (O_1049,N_6519,N_9653);
or UO_1050 (O_1050,N_8590,N_8142);
nand UO_1051 (O_1051,N_5983,N_5660);
nor UO_1052 (O_1052,N_6483,N_5319);
and UO_1053 (O_1053,N_7905,N_9898);
xnor UO_1054 (O_1054,N_6057,N_8312);
or UO_1055 (O_1055,N_7534,N_8786);
xor UO_1056 (O_1056,N_5825,N_9977);
or UO_1057 (O_1057,N_6652,N_9585);
nor UO_1058 (O_1058,N_7923,N_6322);
or UO_1059 (O_1059,N_8753,N_6264);
xor UO_1060 (O_1060,N_9521,N_7513);
or UO_1061 (O_1061,N_7752,N_6668);
nor UO_1062 (O_1062,N_9486,N_8481);
xor UO_1063 (O_1063,N_5992,N_8651);
and UO_1064 (O_1064,N_6378,N_9640);
and UO_1065 (O_1065,N_5119,N_9514);
nor UO_1066 (O_1066,N_9454,N_8615);
or UO_1067 (O_1067,N_5160,N_7881);
and UO_1068 (O_1068,N_9182,N_8987);
or UO_1069 (O_1069,N_9917,N_6098);
and UO_1070 (O_1070,N_9367,N_8237);
or UO_1071 (O_1071,N_6261,N_5051);
nand UO_1072 (O_1072,N_7772,N_8700);
nand UO_1073 (O_1073,N_6815,N_5131);
nor UO_1074 (O_1074,N_8832,N_8052);
or UO_1075 (O_1075,N_7963,N_9466);
xnor UO_1076 (O_1076,N_5122,N_7334);
xnor UO_1077 (O_1077,N_8062,N_8099);
xnor UO_1078 (O_1078,N_9491,N_5022);
xnor UO_1079 (O_1079,N_8030,N_9716);
nand UO_1080 (O_1080,N_6856,N_8814);
xnor UO_1081 (O_1081,N_8348,N_8594);
or UO_1082 (O_1082,N_6520,N_8807);
or UO_1083 (O_1083,N_7220,N_6466);
xor UO_1084 (O_1084,N_9255,N_5598);
nand UO_1085 (O_1085,N_9363,N_9668);
or UO_1086 (O_1086,N_9163,N_7423);
nand UO_1087 (O_1087,N_9425,N_7148);
and UO_1088 (O_1088,N_9015,N_7352);
and UO_1089 (O_1089,N_8970,N_8976);
nand UO_1090 (O_1090,N_6704,N_6019);
nor UO_1091 (O_1091,N_7231,N_5302);
and UO_1092 (O_1092,N_6512,N_7550);
and UO_1093 (O_1093,N_8305,N_5815);
nand UO_1094 (O_1094,N_5135,N_6005);
xnor UO_1095 (O_1095,N_9848,N_6478);
xnor UO_1096 (O_1096,N_7419,N_8922);
xnor UO_1097 (O_1097,N_9344,N_5757);
nand UO_1098 (O_1098,N_9507,N_7803);
or UO_1099 (O_1099,N_7805,N_6106);
and UO_1100 (O_1100,N_9655,N_8677);
nand UO_1101 (O_1101,N_8478,N_6375);
or UO_1102 (O_1102,N_7480,N_6272);
and UO_1103 (O_1103,N_7795,N_5112);
and UO_1104 (O_1104,N_7002,N_6154);
nor UO_1105 (O_1105,N_6778,N_8699);
or UO_1106 (O_1106,N_6651,N_9876);
and UO_1107 (O_1107,N_7207,N_9581);
and UO_1108 (O_1108,N_7336,N_5820);
or UO_1109 (O_1109,N_8946,N_7956);
or UO_1110 (O_1110,N_9415,N_9928);
nand UO_1111 (O_1111,N_6492,N_7139);
nand UO_1112 (O_1112,N_6403,N_9722);
nor UO_1113 (O_1113,N_8597,N_7326);
nand UO_1114 (O_1114,N_7620,N_9487);
nand UO_1115 (O_1115,N_5515,N_8144);
nor UO_1116 (O_1116,N_5802,N_6372);
nor UO_1117 (O_1117,N_6944,N_6869);
and UO_1118 (O_1118,N_6753,N_8884);
nand UO_1119 (O_1119,N_6989,N_8508);
and UO_1120 (O_1120,N_6895,N_7825);
nor UO_1121 (O_1121,N_6844,N_5607);
xor UO_1122 (O_1122,N_8464,N_6491);
and UO_1123 (O_1123,N_6208,N_6438);
xnor UO_1124 (O_1124,N_7776,N_7695);
nor UO_1125 (O_1125,N_8980,N_8588);
nand UO_1126 (O_1126,N_9986,N_7866);
and UO_1127 (O_1127,N_8253,N_8333);
nand UO_1128 (O_1128,N_7809,N_9352);
or UO_1129 (O_1129,N_5446,N_8779);
xnor UO_1130 (O_1130,N_6331,N_5231);
and UO_1131 (O_1131,N_9854,N_7409);
nor UO_1132 (O_1132,N_8882,N_7553);
and UO_1133 (O_1133,N_8731,N_7263);
and UO_1134 (O_1134,N_7224,N_9874);
nor UO_1135 (O_1135,N_8850,N_7984);
xnor UO_1136 (O_1136,N_8152,N_5480);
xor UO_1137 (O_1137,N_6348,N_8628);
nor UO_1138 (O_1138,N_9431,N_9843);
or UO_1139 (O_1139,N_8095,N_5016);
and UO_1140 (O_1140,N_5027,N_5450);
nor UO_1141 (O_1141,N_8427,N_6968);
nor UO_1142 (O_1142,N_6159,N_6935);
xnor UO_1143 (O_1143,N_8849,N_7355);
xor UO_1144 (O_1144,N_9103,N_5572);
and UO_1145 (O_1145,N_6945,N_5824);
nor UO_1146 (O_1146,N_7562,N_7890);
nor UO_1147 (O_1147,N_7541,N_5382);
nor UO_1148 (O_1148,N_7973,N_5518);
and UO_1149 (O_1149,N_6828,N_9002);
and UO_1150 (O_1150,N_9323,N_6015);
or UO_1151 (O_1151,N_9745,N_5408);
and UO_1152 (O_1152,N_8229,N_8969);
nor UO_1153 (O_1153,N_5730,N_5331);
and UO_1154 (O_1154,N_9089,N_6461);
nand UO_1155 (O_1155,N_6006,N_8662);
and UO_1156 (O_1156,N_8929,N_9739);
xnor UO_1157 (O_1157,N_7876,N_7995);
xnor UO_1158 (O_1158,N_8990,N_5106);
or UO_1159 (O_1159,N_5196,N_9949);
and UO_1160 (O_1160,N_8056,N_7977);
nor UO_1161 (O_1161,N_8557,N_8803);
and UO_1162 (O_1162,N_9134,N_6615);
nor UO_1163 (O_1163,N_5732,N_9948);
xor UO_1164 (O_1164,N_7985,N_6145);
nand UO_1165 (O_1165,N_7176,N_6892);
nor UO_1166 (O_1166,N_6893,N_8852);
nor UO_1167 (O_1167,N_6558,N_9777);
nand UO_1168 (O_1168,N_9888,N_8798);
nand UO_1169 (O_1169,N_9407,N_6347);
and UO_1170 (O_1170,N_5918,N_5388);
nand UO_1171 (O_1171,N_7062,N_9328);
nand UO_1172 (O_1172,N_5103,N_5460);
or UO_1173 (O_1173,N_8592,N_6709);
or UO_1174 (O_1174,N_8965,N_6823);
nor UO_1175 (O_1175,N_7957,N_9051);
and UO_1176 (O_1176,N_8067,N_8211);
and UO_1177 (O_1177,N_7670,N_8767);
nand UO_1178 (O_1178,N_9687,N_6234);
nand UO_1179 (O_1179,N_9749,N_8114);
xnor UO_1180 (O_1180,N_9617,N_6860);
and UO_1181 (O_1181,N_5197,N_7034);
nand UO_1182 (O_1182,N_6449,N_5803);
xor UO_1183 (O_1183,N_6124,N_7271);
and UO_1184 (O_1184,N_9923,N_8315);
nand UO_1185 (O_1185,N_9705,N_7529);
nor UO_1186 (O_1186,N_7579,N_8982);
nand UO_1187 (O_1187,N_6452,N_6180);
xnor UO_1188 (O_1188,N_6354,N_8299);
or UO_1189 (O_1189,N_9139,N_5045);
nor UO_1190 (O_1190,N_6021,N_7714);
xor UO_1191 (O_1191,N_8178,N_5294);
and UO_1192 (O_1192,N_6292,N_5764);
nand UO_1193 (O_1193,N_9915,N_5002);
nand UO_1194 (O_1194,N_6855,N_8248);
and UO_1195 (O_1195,N_8361,N_5431);
nor UO_1196 (O_1196,N_8087,N_9513);
nand UO_1197 (O_1197,N_8640,N_7779);
and UO_1198 (O_1198,N_5936,N_6162);
nand UO_1199 (O_1199,N_8530,N_5018);
or UO_1200 (O_1200,N_7715,N_9684);
nor UO_1201 (O_1201,N_8311,N_5925);
or UO_1202 (O_1202,N_9080,N_6333);
nor UO_1203 (O_1203,N_9616,N_8948);
nor UO_1204 (O_1204,N_9813,N_7138);
and UO_1205 (O_1205,N_9504,N_8601);
nand UO_1206 (O_1206,N_7295,N_9620);
nor UO_1207 (O_1207,N_6993,N_6360);
or UO_1208 (O_1208,N_7566,N_8632);
and UO_1209 (O_1209,N_6549,N_9358);
and UO_1210 (O_1210,N_5449,N_9987);
and UO_1211 (O_1211,N_7296,N_9743);
and UO_1212 (O_1212,N_5558,N_9168);
and UO_1213 (O_1213,N_5551,N_9181);
nor UO_1214 (O_1214,N_8261,N_5874);
or UO_1215 (O_1215,N_6094,N_7171);
or UO_1216 (O_1216,N_8854,N_7546);
xor UO_1217 (O_1217,N_9083,N_5951);
xnor UO_1218 (O_1218,N_7037,N_9570);
xor UO_1219 (O_1219,N_7927,N_6915);
or UO_1220 (O_1220,N_6310,N_5788);
nor UO_1221 (O_1221,N_6783,N_7699);
and UO_1222 (O_1222,N_6494,N_9246);
xnor UO_1223 (O_1223,N_8076,N_5260);
nand UO_1224 (O_1224,N_8961,N_6717);
or UO_1225 (O_1225,N_9584,N_7601);
nor UO_1226 (O_1226,N_6939,N_5308);
nand UO_1227 (O_1227,N_6076,N_8614);
xnor UO_1228 (O_1228,N_5793,N_6212);
xor UO_1229 (O_1229,N_6841,N_7430);
nand UO_1230 (O_1230,N_5089,N_8531);
xnor UO_1231 (O_1231,N_5349,N_8619);
nor UO_1232 (O_1232,N_5011,N_5796);
nand UO_1233 (O_1233,N_5205,N_7821);
or UO_1234 (O_1234,N_8973,N_9405);
nand UO_1235 (O_1235,N_8778,N_5136);
or UO_1236 (O_1236,N_8524,N_7397);
nor UO_1237 (O_1237,N_7387,N_7394);
nor UO_1238 (O_1238,N_7567,N_7333);
xnor UO_1239 (O_1239,N_5330,N_9497);
nor UO_1240 (O_1240,N_9009,N_6072);
nand UO_1241 (O_1241,N_6684,N_5876);
nand UO_1242 (O_1242,N_7234,N_5738);
nor UO_1243 (O_1243,N_7206,N_6014);
nor UO_1244 (O_1244,N_9378,N_7594);
or UO_1245 (O_1245,N_9537,N_5939);
or UO_1246 (O_1246,N_8024,N_6326);
or UO_1247 (O_1247,N_8571,N_6262);
and UO_1248 (O_1248,N_9390,N_7331);
xnor UO_1249 (O_1249,N_8967,N_9252);
xor UO_1250 (O_1250,N_6985,N_5705);
nor UO_1251 (O_1251,N_6143,N_5307);
or UO_1252 (O_1252,N_6733,N_5927);
xor UO_1253 (O_1253,N_7160,N_8855);
nand UO_1254 (O_1254,N_7596,N_6640);
nor UO_1255 (O_1255,N_6443,N_6725);
or UO_1256 (O_1256,N_8057,N_8436);
nand UO_1257 (O_1257,N_6336,N_9769);
nand UO_1258 (O_1258,N_8280,N_5553);
and UO_1259 (O_1259,N_7765,N_9784);
nand UO_1260 (O_1260,N_6691,N_8403);
and UO_1261 (O_1261,N_6885,N_6158);
nand UO_1262 (O_1262,N_9667,N_7174);
nor UO_1263 (O_1263,N_6305,N_5714);
nand UO_1264 (O_1264,N_6377,N_7200);
and UO_1265 (O_1265,N_8881,N_6267);
and UO_1266 (O_1266,N_7273,N_8547);
or UO_1267 (O_1267,N_8609,N_6843);
nand UO_1268 (O_1268,N_7165,N_8802);
and UO_1269 (O_1269,N_9021,N_5001);
nor UO_1270 (O_1270,N_5721,N_9177);
and UO_1271 (O_1271,N_8587,N_7560);
nand UO_1272 (O_1272,N_8264,N_7253);
nor UO_1273 (O_1273,N_9499,N_8666);
or UO_1274 (O_1274,N_5156,N_8745);
or UO_1275 (O_1275,N_9314,N_5372);
xor UO_1276 (O_1276,N_6140,N_6102);
or UO_1277 (O_1277,N_8867,N_9063);
xnor UO_1278 (O_1278,N_8357,N_6838);
nand UO_1279 (O_1279,N_8439,N_6655);
nor UO_1280 (O_1280,N_6061,N_5911);
nor UO_1281 (O_1281,N_7446,N_7990);
nor UO_1282 (O_1282,N_5093,N_9596);
or UO_1283 (O_1283,N_5441,N_8244);
or UO_1284 (O_1284,N_5352,N_7675);
nor UO_1285 (O_1285,N_9039,N_8673);
or UO_1286 (O_1286,N_9259,N_6914);
or UO_1287 (O_1287,N_9897,N_7826);
xor UO_1288 (O_1288,N_9686,N_8060);
or UO_1289 (O_1289,N_9333,N_9619);
or UO_1290 (O_1290,N_7467,N_8653);
nand UO_1291 (O_1291,N_5209,N_9760);
xnor UO_1292 (O_1292,N_5041,N_5447);
nor UO_1293 (O_1293,N_8808,N_7616);
xor UO_1294 (O_1294,N_5362,N_7965);
and UO_1295 (O_1295,N_6128,N_9446);
or UO_1296 (O_1296,N_9402,N_5335);
or UO_1297 (O_1297,N_9430,N_5338);
or UO_1298 (O_1298,N_9043,N_8323);
xnor UO_1299 (O_1299,N_8022,N_5130);
nor UO_1300 (O_1300,N_5057,N_8377);
xor UO_1301 (O_1301,N_6131,N_9437);
and UO_1302 (O_1302,N_6400,N_5612);
xor UO_1303 (O_1303,N_7278,N_5900);
and UO_1304 (O_1304,N_5114,N_5630);
or UO_1305 (O_1305,N_9108,N_9675);
nand UO_1306 (O_1306,N_8574,N_7663);
or UO_1307 (O_1307,N_7530,N_6499);
xnor UO_1308 (O_1308,N_6767,N_7609);
nor UO_1309 (O_1309,N_7619,N_6042);
nand UO_1310 (O_1310,N_9706,N_6257);
xnor UO_1311 (O_1311,N_8726,N_8902);
nand UO_1312 (O_1312,N_7960,N_8360);
nor UO_1313 (O_1313,N_6455,N_9886);
and UO_1314 (O_1314,N_8669,N_6697);
and UO_1315 (O_1315,N_7721,N_9172);
or UO_1316 (O_1316,N_6592,N_7144);
and UO_1317 (O_1317,N_9227,N_7288);
nor UO_1318 (O_1318,N_8356,N_6409);
nor UO_1319 (O_1319,N_6619,N_8828);
nor UO_1320 (O_1320,N_5236,N_7800);
or UO_1321 (O_1321,N_5823,N_6567);
xnor UO_1322 (O_1322,N_6288,N_9061);
or UO_1323 (O_1323,N_5171,N_5394);
xor UO_1324 (O_1324,N_7110,N_7556);
nand UO_1325 (O_1325,N_6884,N_6226);
nand UO_1326 (O_1326,N_5015,N_7948);
and UO_1327 (O_1327,N_5292,N_9756);
and UO_1328 (O_1328,N_6200,N_6781);
xnor UO_1329 (O_1329,N_7267,N_6421);
nand UO_1330 (O_1330,N_6417,N_6073);
nand UO_1331 (O_1331,N_7549,N_8582);
or UO_1332 (O_1332,N_5538,N_9034);
or UO_1333 (O_1333,N_5052,N_7978);
or UO_1334 (O_1334,N_7898,N_9337);
and UO_1335 (O_1335,N_8385,N_9839);
nand UO_1336 (O_1336,N_7888,N_6083);
nor UO_1337 (O_1337,N_5935,N_8698);
xor UO_1338 (O_1338,N_7473,N_5958);
nor UO_1339 (O_1339,N_8276,N_5475);
and UO_1340 (O_1340,N_9401,N_7865);
xnor UO_1341 (O_1341,N_7831,N_5966);
xnor UO_1342 (O_1342,N_9690,N_8912);
nor UO_1343 (O_1343,N_9321,N_7909);
nor UO_1344 (O_1344,N_5833,N_5386);
and UO_1345 (O_1345,N_7761,N_6245);
and UO_1346 (O_1346,N_7853,N_8159);
or UO_1347 (O_1347,N_6390,N_7082);
xnor UO_1348 (O_1348,N_8039,N_6857);
and UO_1349 (O_1349,N_9202,N_6629);
and UO_1350 (O_1350,N_8568,N_5682);
or UO_1351 (O_1351,N_5928,N_6286);
or UO_1352 (O_1352,N_5954,N_7704);
nand UO_1353 (O_1353,N_5959,N_6966);
nor UO_1354 (O_1354,N_8279,N_9547);
nand UO_1355 (O_1355,N_6551,N_6800);
nand UO_1356 (O_1356,N_6416,N_7523);
and UO_1357 (O_1357,N_6244,N_5505);
nor UO_1358 (O_1358,N_5059,N_5464);
xor UO_1359 (O_1359,N_6814,N_9073);
or UO_1360 (O_1360,N_8629,N_5213);
or UO_1361 (O_1361,N_9326,N_7557);
or UO_1362 (O_1362,N_9385,N_8616);
nor UO_1363 (O_1363,N_6132,N_7608);
or UO_1364 (O_1364,N_7830,N_5404);
and UO_1365 (O_1365,N_6247,N_8161);
nand UO_1366 (O_1366,N_5008,N_8499);
nor UO_1367 (O_1367,N_6155,N_8953);
xor UO_1368 (O_1368,N_5703,N_5753);
xnor UO_1369 (O_1369,N_8602,N_9532);
xnor UO_1370 (O_1370,N_8113,N_6000);
and UO_1371 (O_1371,N_8106,N_6859);
nand UO_1372 (O_1372,N_9635,N_5073);
nor UO_1373 (O_1373,N_7440,N_8796);
xor UO_1374 (O_1374,N_8580,N_6608);
nor UO_1375 (O_1375,N_5429,N_5489);
xor UO_1376 (O_1376,N_5087,N_8543);
or UO_1377 (O_1377,N_6925,N_8175);
nand UO_1378 (O_1378,N_5529,N_8495);
or UO_1379 (O_1379,N_6203,N_6327);
nor UO_1380 (O_1380,N_7268,N_7703);
nand UO_1381 (O_1381,N_7181,N_8493);
and UO_1382 (O_1382,N_8314,N_5989);
and UO_1383 (O_1383,N_9004,N_7111);
xnor UO_1384 (O_1384,N_7270,N_8904);
nor UO_1385 (O_1385,N_9812,N_9153);
xor UO_1386 (O_1386,N_8317,N_9661);
or UO_1387 (O_1387,N_5712,N_8693);
and UO_1388 (O_1388,N_9411,N_9422);
or UO_1389 (O_1389,N_5524,N_8869);
nand UO_1390 (O_1390,N_7315,N_5521);
nor UO_1391 (O_1391,N_9214,N_9203);
and UO_1392 (O_1392,N_8523,N_9539);
nand UO_1393 (O_1393,N_6653,N_7366);
or UO_1394 (O_1394,N_5504,N_7716);
nand UO_1395 (O_1395,N_9944,N_6318);
xnor UO_1396 (O_1396,N_7080,N_5736);
and UO_1397 (O_1397,N_8851,N_5858);
nor UO_1398 (O_1398,N_5278,N_5170);
xnor UO_1399 (O_1399,N_7184,N_8174);
and UO_1400 (O_1400,N_6505,N_9334);
or UO_1401 (O_1401,N_6405,N_7389);
or UO_1402 (O_1402,N_8452,N_7683);
nand UO_1403 (O_1403,N_6091,N_8857);
nand UO_1404 (O_1404,N_9354,N_6255);
nor UO_1405 (O_1405,N_5065,N_7054);
nor UO_1406 (O_1406,N_9305,N_8135);
or UO_1407 (O_1407,N_8117,N_5511);
nand UO_1408 (O_1408,N_9175,N_7367);
nor UO_1409 (O_1409,N_9719,N_9967);
xor UO_1410 (O_1410,N_7816,N_9634);
or UO_1411 (O_1411,N_9841,N_8831);
xor UO_1412 (O_1412,N_7559,N_5000);
nand UO_1413 (O_1413,N_9283,N_6695);
or UO_1414 (O_1414,N_5370,N_9226);
xor UO_1415 (O_1415,N_9872,N_8810);
nand UO_1416 (O_1416,N_6231,N_7555);
xnor UO_1417 (O_1417,N_9714,N_5419);
nand UO_1418 (O_1418,N_7401,N_7794);
nand UO_1419 (O_1419,N_7021,N_7004);
and UO_1420 (O_1420,N_8243,N_6880);
xnor UO_1421 (O_1421,N_6431,N_5893);
nand UO_1422 (O_1422,N_5361,N_5047);
and UO_1423 (O_1423,N_7012,N_7512);
or UO_1424 (O_1424,N_8477,N_9710);
nor UO_1425 (O_1425,N_9538,N_6521);
xnor UO_1426 (O_1426,N_5791,N_9024);
nor UO_1427 (O_1427,N_8255,N_5771);
nand UO_1428 (O_1428,N_8145,N_7854);
and UO_1429 (O_1429,N_5837,N_8553);
xnor UO_1430 (O_1430,N_6100,N_8210);
nand UO_1431 (O_1431,N_8915,N_5074);
or UO_1432 (O_1432,N_9125,N_9237);
or UO_1433 (O_1433,N_9701,N_6393);
or UO_1434 (O_1434,N_6368,N_8455);
xor UO_1435 (O_1435,N_6740,N_7827);
or UO_1436 (O_1436,N_7025,N_7625);
xor UO_1437 (O_1437,N_6302,N_8220);
xnor UO_1438 (O_1438,N_9605,N_5604);
nand UO_1439 (O_1439,N_5218,N_5118);
nor UO_1440 (O_1440,N_8120,N_6080);
or UO_1441 (O_1441,N_8103,N_5206);
or UO_1442 (O_1442,N_6606,N_5628);
or UO_1443 (O_1443,N_8330,N_7793);
and UO_1444 (O_1444,N_6803,N_8184);
nand UO_1445 (O_1445,N_9594,N_5493);
or UO_1446 (O_1446,N_7603,N_7036);
and UO_1447 (O_1447,N_7768,N_7006);
nor UO_1448 (O_1448,N_7454,N_6917);
xor UO_1449 (O_1449,N_9557,N_7811);
or UO_1450 (O_1450,N_8086,N_8239);
nand UO_1451 (O_1451,N_5539,N_8504);
or UO_1452 (O_1452,N_8476,N_9997);
nand UO_1453 (O_1453,N_5448,N_8040);
nor UO_1454 (O_1454,N_7738,N_9518);
or UO_1455 (O_1455,N_8780,N_5986);
nand UO_1456 (O_1456,N_9577,N_5756);
xor UO_1457 (O_1457,N_6436,N_9376);
and UO_1458 (O_1458,N_8288,N_6056);
xor UO_1459 (O_1459,N_9032,N_8128);
and UO_1460 (O_1460,N_9597,N_8240);
and UO_1461 (O_1461,N_9185,N_5562);
and UO_1462 (O_1462,N_5050,N_7279);
and UO_1463 (O_1463,N_8257,N_6720);
nand UO_1464 (O_1464,N_7130,N_7303);
nor UO_1465 (O_1465,N_8335,N_7748);
and UO_1466 (O_1466,N_5644,N_5469);
nor UO_1467 (O_1467,N_8527,N_6672);
or UO_1468 (O_1468,N_7665,N_5451);
nand UO_1469 (O_1469,N_7413,N_5500);
and UO_1470 (O_1470,N_5818,N_8072);
xor UO_1471 (O_1471,N_6202,N_7624);
nand UO_1472 (O_1472,N_5938,N_5474);
xnor UO_1473 (O_1473,N_9780,N_9014);
or UO_1474 (O_1474,N_8516,N_8396);
nand UO_1475 (O_1475,N_9579,N_7218);
nor UO_1476 (O_1476,N_7810,N_6134);
or UO_1477 (O_1477,N_5908,N_6956);
nor UO_1478 (O_1478,N_7903,N_7081);
or UO_1479 (O_1479,N_6424,N_6751);
xnor UO_1480 (O_1480,N_9724,N_5586);
and UO_1481 (O_1481,N_7617,N_7808);
nand UO_1482 (O_1482,N_7878,N_5686);
nor UO_1483 (O_1483,N_9590,N_6665);
nand UO_1484 (O_1484,N_5742,N_6762);
xor UO_1485 (O_1485,N_5565,N_7085);
and UO_1486 (O_1486,N_7709,N_5610);
xnor UO_1487 (O_1487,N_5265,N_7871);
nand UO_1488 (O_1488,N_6123,N_7390);
nor UO_1489 (O_1489,N_8107,N_7061);
nand UO_1490 (O_1490,N_6233,N_6946);
nand UO_1491 (O_1491,N_5281,N_9527);
nor UO_1492 (O_1492,N_8258,N_7637);
xnor UO_1493 (O_1493,N_5385,N_9636);
nor UO_1494 (O_1494,N_5503,N_5491);
xnor UO_1495 (O_1495,N_5257,N_7759);
and UO_1496 (O_1496,N_6943,N_5426);
xor UO_1497 (O_1497,N_7750,N_8242);
nand UO_1498 (O_1498,N_6578,N_5032);
nor UO_1499 (O_1499,N_5262,N_5339);
endmodule