module basic_500_3000_500_40_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_13,In_142);
and U1 (N_1,In_265,In_445);
and U2 (N_2,In_38,In_143);
nor U3 (N_3,In_192,In_106);
nor U4 (N_4,In_468,In_76);
or U5 (N_5,In_286,In_408);
nand U6 (N_6,In_206,In_128);
or U7 (N_7,In_1,In_341);
xor U8 (N_8,In_260,In_419);
nor U9 (N_9,In_239,In_209);
or U10 (N_10,In_384,In_91);
or U11 (N_11,In_197,In_22);
nor U12 (N_12,In_162,In_233);
nor U13 (N_13,In_362,In_159);
nor U14 (N_14,In_495,In_418);
nand U15 (N_15,In_194,In_37);
nor U16 (N_16,In_393,In_67);
or U17 (N_17,In_114,In_139);
or U18 (N_18,In_325,In_88);
and U19 (N_19,In_157,In_476);
nor U20 (N_20,In_3,In_25);
xor U21 (N_21,In_285,In_43);
and U22 (N_22,In_52,In_41);
or U23 (N_23,In_327,In_296);
or U24 (N_24,In_211,In_44);
nand U25 (N_25,In_299,In_245);
nor U26 (N_26,In_112,In_494);
and U27 (N_27,In_219,In_116);
nand U28 (N_28,In_102,In_144);
and U29 (N_29,In_496,In_361);
xor U30 (N_30,In_94,In_170);
nand U31 (N_31,In_349,In_326);
nor U32 (N_32,In_30,In_431);
nand U33 (N_33,In_90,In_357);
and U34 (N_34,In_228,In_229);
and U35 (N_35,In_140,In_26);
nand U36 (N_36,In_372,In_356);
and U37 (N_37,In_263,In_50);
and U38 (N_38,In_0,In_173);
or U39 (N_39,In_31,In_230);
nand U40 (N_40,In_183,In_342);
nor U41 (N_41,In_380,In_89);
nor U42 (N_42,In_389,In_123);
nand U43 (N_43,In_334,In_352);
and U44 (N_44,In_291,In_332);
nand U45 (N_45,In_413,In_166);
xnor U46 (N_46,In_121,In_359);
nand U47 (N_47,In_451,In_218);
or U48 (N_48,In_127,In_227);
and U49 (N_49,In_403,In_18);
xnor U50 (N_50,In_369,In_45);
or U51 (N_51,In_117,In_175);
xnor U52 (N_52,In_274,In_104);
nor U53 (N_53,In_270,In_367);
and U54 (N_54,In_93,In_257);
and U55 (N_55,In_81,In_204);
nor U56 (N_56,In_379,In_399);
or U57 (N_57,In_436,In_35);
nor U58 (N_58,In_467,In_344);
nand U59 (N_59,In_382,In_168);
or U60 (N_60,In_338,In_92);
nand U61 (N_61,In_289,In_199);
nor U62 (N_62,In_484,In_32);
or U63 (N_63,In_15,In_475);
and U64 (N_64,In_259,In_256);
nand U65 (N_65,In_111,In_234);
nor U66 (N_66,In_46,In_63);
nor U67 (N_67,In_115,In_450);
nor U68 (N_68,In_61,In_130);
or U69 (N_69,In_150,In_388);
nand U70 (N_70,In_411,In_179);
and U71 (N_71,In_201,In_207);
nor U72 (N_72,In_360,In_283);
or U73 (N_73,In_442,In_138);
nand U74 (N_74,In_141,In_315);
or U75 (N_75,In_16,In_188);
nor U76 (N_76,In_276,In_282);
and U77 (N_77,N_24,In_428);
nand U78 (N_78,In_86,N_45);
nand U79 (N_79,N_8,In_290);
nor U80 (N_80,In_136,In_264);
nor U81 (N_81,In_232,In_96);
or U82 (N_82,N_26,In_486);
nor U83 (N_83,In_350,In_103);
nand U84 (N_84,In_180,In_237);
and U85 (N_85,In_202,In_12);
nand U86 (N_86,In_156,In_308);
nor U87 (N_87,In_490,N_38);
nand U88 (N_88,In_298,In_297);
nand U89 (N_89,In_160,N_43);
and U90 (N_90,In_246,In_371);
nand U91 (N_91,In_163,In_288);
nor U92 (N_92,In_322,N_58);
nor U93 (N_93,In_73,In_345);
or U94 (N_94,N_59,In_80);
xor U95 (N_95,In_107,In_307);
nor U96 (N_96,In_383,In_7);
or U97 (N_97,In_225,In_177);
and U98 (N_98,In_217,N_32);
nor U99 (N_99,In_244,In_433);
xnor U100 (N_100,In_205,In_129);
nor U101 (N_101,In_462,N_33);
and U102 (N_102,In_165,In_196);
nand U103 (N_103,In_365,In_184);
or U104 (N_104,In_465,In_493);
nand U105 (N_105,N_53,In_429);
nor U106 (N_106,In_58,N_66);
nor U107 (N_107,N_18,In_385);
nor U108 (N_108,In_97,In_459);
nor U109 (N_109,In_323,In_24);
nand U110 (N_110,In_453,In_421);
or U111 (N_111,N_54,In_85);
nor U112 (N_112,In_152,In_28);
nor U113 (N_113,In_294,In_272);
or U114 (N_114,In_321,In_249);
and U115 (N_115,In_118,In_19);
and U116 (N_116,In_251,N_40);
xnor U117 (N_117,In_377,In_443);
xnor U118 (N_118,In_71,In_409);
nor U119 (N_119,In_198,In_9);
and U120 (N_120,In_463,In_69);
and U121 (N_121,In_448,In_222);
nand U122 (N_122,N_49,In_119);
or U123 (N_123,In_303,In_392);
or U124 (N_124,In_213,In_223);
or U125 (N_125,In_471,In_376);
nor U126 (N_126,In_269,In_72);
and U127 (N_127,In_499,In_330);
nand U128 (N_128,In_478,In_191);
xor U129 (N_129,In_231,In_34);
xnor U130 (N_130,In_423,N_7);
and U131 (N_131,In_224,In_410);
nand U132 (N_132,N_36,N_65);
or U133 (N_133,N_17,In_62);
xor U134 (N_134,In_253,In_149);
or U135 (N_135,In_311,In_238);
and U136 (N_136,In_275,In_295);
nand U137 (N_137,In_64,N_41);
nor U138 (N_138,In_407,In_491);
xor U139 (N_139,In_262,N_74);
nand U140 (N_140,In_59,N_31);
and U141 (N_141,N_15,In_487);
xnor U142 (N_142,In_439,In_266);
xor U143 (N_143,N_73,In_440);
or U144 (N_144,In_355,In_182);
and U145 (N_145,In_398,In_187);
and U146 (N_146,In_454,In_461);
xnor U147 (N_147,In_381,N_19);
nor U148 (N_148,In_447,In_279);
and U149 (N_149,N_13,In_489);
nand U150 (N_150,N_9,In_248);
nor U151 (N_151,In_422,In_36);
nand U152 (N_152,N_105,N_30);
and U153 (N_153,In_5,N_0);
or U154 (N_154,In_126,N_145);
xnor U155 (N_155,In_414,In_66);
or U156 (N_156,In_135,In_108);
nor U157 (N_157,N_111,In_425);
nor U158 (N_158,N_137,N_34);
nor U159 (N_159,In_100,In_220);
nand U160 (N_160,N_142,N_2);
nor U161 (N_161,N_101,N_104);
nand U162 (N_162,N_89,In_420);
or U163 (N_163,In_171,In_292);
nand U164 (N_164,In_20,In_470);
nand U165 (N_165,In_354,In_124);
nand U166 (N_166,In_56,In_75);
or U167 (N_167,In_99,N_4);
and U168 (N_168,N_100,In_455);
xnor U169 (N_169,N_80,In_469);
or U170 (N_170,N_124,In_84);
or U171 (N_171,N_84,N_109);
or U172 (N_172,N_5,N_23);
and U173 (N_173,N_88,N_126);
and U174 (N_174,N_76,N_21);
nand U175 (N_175,In_95,In_319);
nand U176 (N_176,In_415,In_146);
and U177 (N_177,N_6,In_333);
nor U178 (N_178,N_46,In_373);
xor U179 (N_179,In_181,In_302);
nand U180 (N_180,In_60,N_44);
nand U181 (N_181,In_17,In_23);
or U182 (N_182,In_57,N_1);
nor U183 (N_183,N_78,N_42);
nor U184 (N_184,N_92,N_48);
or U185 (N_185,N_120,In_200);
and U186 (N_186,In_4,N_81);
or U187 (N_187,In_479,In_472);
and U188 (N_188,In_261,In_424);
nand U189 (N_189,In_167,N_68);
xnor U190 (N_190,In_27,N_91);
nand U191 (N_191,In_132,N_144);
xnor U192 (N_192,N_148,In_174);
and U193 (N_193,N_116,In_329);
and U194 (N_194,In_314,In_460);
and U195 (N_195,In_358,N_106);
nor U196 (N_196,In_391,In_313);
nand U197 (N_197,In_430,In_161);
nor U198 (N_198,N_136,In_301);
nand U199 (N_199,In_87,In_435);
or U200 (N_200,In_318,In_390);
or U201 (N_201,N_14,In_397);
nand U202 (N_202,N_130,In_169);
xnor U203 (N_203,In_33,In_396);
nor U204 (N_204,N_39,In_304);
nand U205 (N_205,In_401,In_221);
nand U206 (N_206,N_128,In_14);
xnor U207 (N_207,N_110,In_214);
or U208 (N_208,In_458,In_79);
nand U209 (N_209,In_190,In_82);
nor U210 (N_210,In_426,In_189);
xnor U211 (N_211,N_51,N_83);
or U212 (N_212,In_151,In_226);
or U213 (N_213,In_497,In_153);
nand U214 (N_214,In_400,In_364);
or U215 (N_215,N_50,In_306);
nand U216 (N_216,In_434,N_134);
nand U217 (N_217,In_6,In_77);
xor U218 (N_218,In_477,In_216);
or U219 (N_219,In_186,In_368);
xor U220 (N_220,N_67,In_155);
xor U221 (N_221,In_178,In_394);
nand U222 (N_222,In_483,In_29);
and U223 (N_223,N_141,In_176);
nand U224 (N_224,In_281,N_125);
or U225 (N_225,In_247,In_481);
and U226 (N_226,In_148,In_147);
and U227 (N_227,N_61,N_209);
nand U228 (N_228,N_168,In_164);
nand U229 (N_229,In_54,In_331);
nand U230 (N_230,In_98,N_97);
xor U231 (N_231,In_212,N_161);
xor U232 (N_232,In_48,N_96);
nand U233 (N_233,N_196,N_29);
nor U234 (N_234,In_474,In_335);
or U235 (N_235,N_223,In_339);
or U236 (N_236,In_109,N_79);
nand U237 (N_237,In_485,In_437);
nand U238 (N_238,N_25,N_198);
nand U239 (N_239,In_386,In_416);
nand U240 (N_240,In_193,In_277);
nor U241 (N_241,In_449,N_164);
nor U242 (N_242,N_153,N_173);
or U243 (N_243,In_498,N_163);
and U244 (N_244,In_122,N_113);
and U245 (N_245,N_191,In_125);
nor U246 (N_246,N_149,N_155);
or U247 (N_247,In_324,In_83);
nand U248 (N_248,In_195,In_271);
nand U249 (N_249,N_205,In_404);
and U250 (N_250,N_69,In_11);
nand U251 (N_251,N_98,In_74);
or U252 (N_252,N_129,In_406);
nand U253 (N_253,In_51,In_105);
nand U254 (N_254,In_466,In_438);
nand U255 (N_255,In_137,N_221);
nand U256 (N_256,In_480,N_139);
nand U257 (N_257,N_176,In_351);
nand U258 (N_258,In_492,In_236);
nor U259 (N_259,N_140,In_235);
nor U260 (N_260,N_211,N_202);
nand U261 (N_261,N_199,N_143);
or U262 (N_262,N_216,N_28);
nor U263 (N_263,In_417,In_252);
nor U264 (N_264,In_208,N_82);
or U265 (N_265,In_346,In_267);
xnor U266 (N_266,In_39,N_102);
nor U267 (N_267,In_293,In_405);
and U268 (N_268,N_62,N_218);
xnor U269 (N_269,N_107,In_133);
nand U270 (N_270,In_456,N_219);
nor U271 (N_271,N_184,N_171);
nand U272 (N_272,N_115,N_154);
nand U273 (N_273,N_206,N_174);
nor U274 (N_274,In_215,N_224);
and U275 (N_275,N_204,In_70);
and U276 (N_276,In_395,N_132);
nand U277 (N_277,In_457,In_242);
xnor U278 (N_278,N_10,N_11);
nand U279 (N_279,N_103,N_179);
nor U280 (N_280,In_370,In_65);
or U281 (N_281,In_240,N_158);
or U282 (N_282,N_60,In_441);
or U283 (N_283,N_150,N_27);
xnor U284 (N_284,In_482,In_47);
nand U285 (N_285,N_94,N_190);
and U286 (N_286,In_268,In_158);
nor U287 (N_287,N_56,N_222);
nor U288 (N_288,In_273,N_117);
nand U289 (N_289,In_203,N_20);
nor U290 (N_290,N_119,In_375);
and U291 (N_291,N_182,N_63);
and U292 (N_292,N_70,N_159);
xor U293 (N_293,N_162,N_180);
or U294 (N_294,In_255,N_72);
nor U295 (N_295,In_374,N_112);
and U296 (N_296,N_95,N_75);
xor U297 (N_297,In_250,In_340);
nand U298 (N_298,N_93,N_217);
or U299 (N_299,In_473,In_172);
or U300 (N_300,In_258,N_284);
or U301 (N_301,N_157,In_378);
nand U302 (N_302,N_178,In_78);
or U303 (N_303,N_254,N_251);
nand U304 (N_304,N_114,N_127);
nor U305 (N_305,N_22,N_203);
or U306 (N_306,In_402,N_274);
or U307 (N_307,N_279,N_247);
nand U308 (N_308,N_269,N_283);
and U309 (N_309,N_87,N_280);
xnor U310 (N_310,N_186,N_241);
nand U311 (N_311,N_256,N_282);
and U312 (N_312,N_257,In_464);
or U313 (N_313,N_135,N_273);
nand U314 (N_314,N_122,N_121);
nor U315 (N_315,N_200,In_284);
or U316 (N_316,N_194,N_267);
and U317 (N_317,N_172,N_210);
or U318 (N_318,N_264,N_201);
and U319 (N_319,In_312,In_131);
nor U320 (N_320,In_134,N_290);
or U321 (N_321,N_208,In_363);
nand U322 (N_322,N_12,N_220);
or U323 (N_323,In_243,N_170);
nand U324 (N_324,In_444,In_387);
or U325 (N_325,N_275,N_252);
and U326 (N_326,N_146,N_212);
nor U327 (N_327,In_353,N_213);
or U328 (N_328,N_238,N_214);
and U329 (N_329,N_240,N_165);
nand U330 (N_330,N_298,N_152);
nor U331 (N_331,In_427,In_278);
and U332 (N_332,N_183,In_53);
or U333 (N_333,In_366,N_86);
or U334 (N_334,N_193,N_227);
nand U335 (N_335,N_295,N_248);
or U336 (N_336,N_77,N_57);
nor U337 (N_337,N_271,N_243);
and U338 (N_338,N_297,In_305);
and U339 (N_339,N_225,In_317);
or U340 (N_340,N_244,N_286);
nor U341 (N_341,In_113,In_10);
xor U342 (N_342,In_185,N_187);
or U343 (N_343,In_348,In_300);
and U344 (N_344,In_2,N_233);
nor U345 (N_345,N_90,N_293);
or U346 (N_346,N_262,N_250);
and U347 (N_347,N_185,N_16);
nor U348 (N_348,N_277,In_343);
xor U349 (N_349,N_3,In_49);
and U350 (N_350,In_210,N_242);
xnor U351 (N_351,N_245,In_42);
or U352 (N_352,N_167,N_268);
xnor U353 (N_353,N_37,In_309);
and U354 (N_354,N_188,N_292);
and U355 (N_355,N_237,N_263);
nor U356 (N_356,In_310,N_260);
nand U357 (N_357,In_488,In_154);
nand U358 (N_358,N_133,In_241);
and U359 (N_359,N_235,N_47);
nor U360 (N_360,N_299,N_123);
or U361 (N_361,N_195,In_280);
xor U362 (N_362,N_215,N_239);
nor U363 (N_363,In_21,N_265);
nand U364 (N_364,In_120,N_236);
nor U365 (N_365,N_138,N_71);
nand U366 (N_366,In_68,N_166);
or U367 (N_367,N_287,In_336);
nor U368 (N_368,N_85,N_276);
and U369 (N_369,N_229,N_64);
nand U370 (N_370,N_255,In_287);
nand U371 (N_371,In_328,N_234);
and U372 (N_372,N_131,In_316);
nor U373 (N_373,N_160,In_446);
or U374 (N_374,N_288,N_285);
or U375 (N_375,N_325,N_338);
or U376 (N_376,N_309,N_359);
nor U377 (N_377,In_452,N_281);
nor U378 (N_378,N_228,N_355);
nor U379 (N_379,N_348,N_326);
nor U380 (N_380,N_339,N_312);
or U381 (N_381,N_311,In_55);
or U382 (N_382,N_361,N_327);
and U383 (N_383,N_337,In_8);
and U384 (N_384,N_345,N_335);
nand U385 (N_385,In_110,N_302);
or U386 (N_386,N_266,N_347);
xor U387 (N_387,N_181,N_356);
nor U388 (N_388,N_371,N_336);
and U389 (N_389,N_317,N_52);
nor U390 (N_390,N_253,N_272);
nor U391 (N_391,N_99,N_278);
and U392 (N_392,N_362,N_333);
nor U393 (N_393,In_145,N_343);
nor U394 (N_394,N_319,N_249);
nand U395 (N_395,N_324,N_156);
xor U396 (N_396,In_347,N_310);
and U397 (N_397,N_351,N_357);
and U398 (N_398,N_330,N_332);
nand U399 (N_399,N_342,N_364);
xnor U400 (N_400,N_55,N_353);
nand U401 (N_401,N_307,N_341);
nand U402 (N_402,N_316,N_372);
nand U403 (N_403,N_314,N_313);
or U404 (N_404,N_360,N_323);
nor U405 (N_405,N_291,N_308);
nand U406 (N_406,N_261,N_374);
nor U407 (N_407,N_35,N_340);
xnor U408 (N_408,N_352,N_147);
or U409 (N_409,N_350,N_349);
or U410 (N_410,N_151,N_118);
or U411 (N_411,N_346,N_303);
xnor U412 (N_412,N_363,N_258);
nor U413 (N_413,N_369,N_270);
and U414 (N_414,N_197,In_40);
nor U415 (N_415,N_232,In_101);
nand U416 (N_416,N_354,N_300);
or U417 (N_417,N_230,N_315);
nand U418 (N_418,N_334,N_108);
and U419 (N_419,N_305,N_177);
nor U420 (N_420,N_306,N_370);
xnor U421 (N_421,N_296,N_358);
and U422 (N_422,N_373,N_321);
nor U423 (N_423,N_304,N_231);
nand U424 (N_424,N_328,N_289);
and U425 (N_425,N_322,N_365);
nand U426 (N_426,In_432,N_329);
or U427 (N_427,N_207,N_175);
or U428 (N_428,In_337,N_259);
and U429 (N_429,N_320,N_192);
xnor U430 (N_430,In_412,N_367);
and U431 (N_431,N_189,N_331);
nand U432 (N_432,N_169,N_294);
xor U433 (N_433,In_320,N_344);
and U434 (N_434,N_366,N_226);
or U435 (N_435,N_318,In_254);
nand U436 (N_436,N_301,N_368);
xnor U437 (N_437,N_246,N_278);
or U438 (N_438,N_361,N_304);
xor U439 (N_439,N_357,N_347);
nand U440 (N_440,N_192,N_52);
nor U441 (N_441,N_361,N_169);
nand U442 (N_442,N_347,N_345);
nor U443 (N_443,N_175,N_151);
or U444 (N_444,In_40,N_331);
and U445 (N_445,N_307,N_231);
and U446 (N_446,In_55,N_333);
and U447 (N_447,N_313,N_353);
nand U448 (N_448,N_361,N_344);
nand U449 (N_449,N_360,N_52);
nor U450 (N_450,N_421,N_422);
or U451 (N_451,N_436,N_398);
and U452 (N_452,N_443,N_376);
or U453 (N_453,N_449,N_419);
and U454 (N_454,N_390,N_439);
and U455 (N_455,N_432,N_413);
xnor U456 (N_456,N_402,N_375);
nand U457 (N_457,N_442,N_445);
or U458 (N_458,N_438,N_394);
xor U459 (N_459,N_407,N_386);
nor U460 (N_460,N_429,N_417);
nand U461 (N_461,N_396,N_378);
nand U462 (N_462,N_400,N_389);
nor U463 (N_463,N_401,N_412);
xor U464 (N_464,N_399,N_385);
xor U465 (N_465,N_448,N_427);
or U466 (N_466,N_393,N_377);
nand U467 (N_467,N_411,N_392);
nand U468 (N_468,N_388,N_403);
nor U469 (N_469,N_395,N_444);
nand U470 (N_470,N_404,N_384);
nor U471 (N_471,N_416,N_434);
nand U472 (N_472,N_428,N_426);
and U473 (N_473,N_435,N_415);
nand U474 (N_474,N_414,N_446);
nand U475 (N_475,N_440,N_405);
or U476 (N_476,N_409,N_406);
or U477 (N_477,N_397,N_423);
or U478 (N_478,N_437,N_430);
or U479 (N_479,N_447,N_387);
or U480 (N_480,N_379,N_382);
nand U481 (N_481,N_380,N_431);
xnor U482 (N_482,N_441,N_418);
nand U483 (N_483,N_408,N_425);
and U484 (N_484,N_383,N_381);
and U485 (N_485,N_424,N_420);
and U486 (N_486,N_410,N_391);
and U487 (N_487,N_433,N_386);
or U488 (N_488,N_382,N_406);
nor U489 (N_489,N_415,N_408);
nor U490 (N_490,N_403,N_438);
nand U491 (N_491,N_448,N_377);
or U492 (N_492,N_379,N_388);
xor U493 (N_493,N_420,N_413);
xnor U494 (N_494,N_417,N_407);
nand U495 (N_495,N_411,N_402);
nor U496 (N_496,N_412,N_446);
nor U497 (N_497,N_410,N_405);
xnor U498 (N_498,N_439,N_427);
nor U499 (N_499,N_412,N_424);
and U500 (N_500,N_434,N_445);
nand U501 (N_501,N_431,N_395);
nand U502 (N_502,N_449,N_416);
nor U503 (N_503,N_411,N_383);
and U504 (N_504,N_416,N_440);
and U505 (N_505,N_394,N_409);
nand U506 (N_506,N_424,N_392);
xnor U507 (N_507,N_412,N_436);
xor U508 (N_508,N_380,N_430);
nor U509 (N_509,N_377,N_389);
and U510 (N_510,N_407,N_393);
or U511 (N_511,N_382,N_444);
nor U512 (N_512,N_449,N_393);
and U513 (N_513,N_413,N_449);
nand U514 (N_514,N_430,N_391);
or U515 (N_515,N_442,N_449);
nand U516 (N_516,N_425,N_395);
and U517 (N_517,N_382,N_411);
or U518 (N_518,N_400,N_442);
nor U519 (N_519,N_398,N_385);
nand U520 (N_520,N_419,N_418);
or U521 (N_521,N_413,N_376);
and U522 (N_522,N_382,N_408);
nand U523 (N_523,N_434,N_402);
and U524 (N_524,N_379,N_414);
or U525 (N_525,N_463,N_458);
nand U526 (N_526,N_487,N_477);
or U527 (N_527,N_508,N_462);
nand U528 (N_528,N_509,N_488);
nand U529 (N_529,N_489,N_514);
or U530 (N_530,N_473,N_453);
nand U531 (N_531,N_516,N_504);
and U532 (N_532,N_479,N_505);
nor U533 (N_533,N_497,N_524);
nor U534 (N_534,N_486,N_481);
nor U535 (N_535,N_459,N_498);
nor U536 (N_536,N_490,N_511);
nor U537 (N_537,N_468,N_470);
and U538 (N_538,N_456,N_455);
and U539 (N_539,N_467,N_520);
nor U540 (N_540,N_496,N_502);
or U541 (N_541,N_466,N_469);
nor U542 (N_542,N_450,N_491);
nor U543 (N_543,N_465,N_460);
xor U544 (N_544,N_503,N_451);
nand U545 (N_545,N_501,N_452);
nand U546 (N_546,N_454,N_484);
nand U547 (N_547,N_475,N_521);
or U548 (N_548,N_478,N_485);
and U549 (N_549,N_483,N_480);
xor U550 (N_550,N_518,N_515);
nor U551 (N_551,N_495,N_507);
nand U552 (N_552,N_464,N_512);
nor U553 (N_553,N_523,N_474);
nor U554 (N_554,N_513,N_461);
nand U555 (N_555,N_492,N_499);
and U556 (N_556,N_472,N_500);
or U557 (N_557,N_506,N_519);
or U558 (N_558,N_510,N_457);
or U559 (N_559,N_493,N_494);
nor U560 (N_560,N_471,N_482);
nand U561 (N_561,N_476,N_517);
nor U562 (N_562,N_522,N_466);
nor U563 (N_563,N_485,N_502);
xor U564 (N_564,N_477,N_485);
or U565 (N_565,N_524,N_488);
nor U566 (N_566,N_494,N_477);
and U567 (N_567,N_460,N_517);
nor U568 (N_568,N_471,N_477);
xor U569 (N_569,N_521,N_479);
and U570 (N_570,N_490,N_503);
xor U571 (N_571,N_469,N_461);
nor U572 (N_572,N_488,N_466);
or U573 (N_573,N_463,N_512);
nand U574 (N_574,N_481,N_497);
nand U575 (N_575,N_485,N_499);
and U576 (N_576,N_466,N_486);
xor U577 (N_577,N_460,N_468);
xnor U578 (N_578,N_520,N_474);
nand U579 (N_579,N_465,N_510);
nor U580 (N_580,N_489,N_459);
and U581 (N_581,N_474,N_502);
xnor U582 (N_582,N_477,N_458);
nor U583 (N_583,N_513,N_473);
nor U584 (N_584,N_475,N_500);
xor U585 (N_585,N_521,N_522);
or U586 (N_586,N_498,N_491);
or U587 (N_587,N_497,N_455);
nor U588 (N_588,N_459,N_470);
nor U589 (N_589,N_473,N_456);
and U590 (N_590,N_505,N_503);
and U591 (N_591,N_487,N_471);
and U592 (N_592,N_465,N_514);
nor U593 (N_593,N_516,N_468);
and U594 (N_594,N_450,N_523);
nand U595 (N_595,N_514,N_511);
nor U596 (N_596,N_485,N_515);
nor U597 (N_597,N_488,N_516);
nor U598 (N_598,N_466,N_517);
nand U599 (N_599,N_520,N_482);
or U600 (N_600,N_552,N_543);
nand U601 (N_601,N_550,N_547);
nor U602 (N_602,N_585,N_590);
or U603 (N_603,N_598,N_587);
nor U604 (N_604,N_536,N_558);
nand U605 (N_605,N_593,N_599);
or U606 (N_606,N_535,N_531);
nand U607 (N_607,N_584,N_554);
nand U608 (N_608,N_576,N_572);
or U609 (N_609,N_575,N_542);
and U610 (N_610,N_557,N_594);
or U611 (N_611,N_528,N_563);
xnor U612 (N_612,N_568,N_577);
nor U613 (N_613,N_553,N_562);
nor U614 (N_614,N_586,N_541);
nor U615 (N_615,N_573,N_589);
nand U616 (N_616,N_527,N_525);
nand U617 (N_617,N_597,N_592);
or U618 (N_618,N_595,N_546);
or U619 (N_619,N_551,N_533);
nand U620 (N_620,N_544,N_588);
nand U621 (N_621,N_555,N_579);
nor U622 (N_622,N_545,N_560);
nand U623 (N_623,N_549,N_564);
nor U624 (N_624,N_596,N_574);
and U625 (N_625,N_566,N_569);
or U626 (N_626,N_578,N_529);
xor U627 (N_627,N_526,N_591);
and U628 (N_628,N_559,N_565);
nor U629 (N_629,N_530,N_534);
and U630 (N_630,N_539,N_538);
or U631 (N_631,N_561,N_537);
nor U632 (N_632,N_581,N_556);
and U633 (N_633,N_571,N_548);
nor U634 (N_634,N_567,N_583);
xor U635 (N_635,N_570,N_582);
xnor U636 (N_636,N_580,N_532);
nor U637 (N_637,N_540,N_599);
or U638 (N_638,N_574,N_550);
or U639 (N_639,N_530,N_546);
nand U640 (N_640,N_539,N_568);
xor U641 (N_641,N_570,N_529);
and U642 (N_642,N_585,N_565);
or U643 (N_643,N_544,N_590);
nor U644 (N_644,N_533,N_574);
or U645 (N_645,N_559,N_583);
and U646 (N_646,N_583,N_593);
and U647 (N_647,N_540,N_552);
nand U648 (N_648,N_533,N_559);
nor U649 (N_649,N_529,N_598);
nor U650 (N_650,N_546,N_541);
nor U651 (N_651,N_557,N_564);
nand U652 (N_652,N_528,N_590);
nor U653 (N_653,N_530,N_594);
nand U654 (N_654,N_579,N_538);
nor U655 (N_655,N_537,N_527);
nand U656 (N_656,N_538,N_559);
or U657 (N_657,N_593,N_548);
xnor U658 (N_658,N_594,N_553);
or U659 (N_659,N_558,N_540);
nand U660 (N_660,N_559,N_527);
and U661 (N_661,N_543,N_530);
or U662 (N_662,N_533,N_557);
nand U663 (N_663,N_580,N_584);
or U664 (N_664,N_562,N_584);
nand U665 (N_665,N_562,N_585);
or U666 (N_666,N_591,N_535);
or U667 (N_667,N_549,N_538);
and U668 (N_668,N_559,N_591);
nand U669 (N_669,N_551,N_526);
nor U670 (N_670,N_582,N_544);
nand U671 (N_671,N_575,N_565);
xor U672 (N_672,N_526,N_559);
or U673 (N_673,N_574,N_527);
and U674 (N_674,N_564,N_563);
nor U675 (N_675,N_644,N_657);
or U676 (N_676,N_631,N_659);
and U677 (N_677,N_661,N_601);
and U678 (N_678,N_669,N_658);
nand U679 (N_679,N_611,N_637);
or U680 (N_680,N_635,N_647);
nand U681 (N_681,N_652,N_629);
nor U682 (N_682,N_630,N_616);
nand U683 (N_683,N_656,N_633);
or U684 (N_684,N_615,N_639);
or U685 (N_685,N_606,N_660);
nor U686 (N_686,N_672,N_636);
or U687 (N_687,N_626,N_649);
and U688 (N_688,N_655,N_627);
nand U689 (N_689,N_620,N_641);
nand U690 (N_690,N_628,N_618);
nor U691 (N_691,N_623,N_668);
nand U692 (N_692,N_663,N_662);
nand U693 (N_693,N_673,N_624);
nor U694 (N_694,N_670,N_612);
and U695 (N_695,N_665,N_600);
nand U696 (N_696,N_674,N_621);
nor U697 (N_697,N_642,N_625);
nand U698 (N_698,N_632,N_634);
or U699 (N_699,N_653,N_671);
nor U700 (N_700,N_650,N_608);
nor U701 (N_701,N_654,N_643);
xor U702 (N_702,N_648,N_646);
nand U703 (N_703,N_617,N_651);
nor U704 (N_704,N_605,N_607);
and U705 (N_705,N_614,N_610);
nor U706 (N_706,N_638,N_640);
xor U707 (N_707,N_664,N_619);
or U708 (N_708,N_622,N_604);
or U709 (N_709,N_645,N_602);
or U710 (N_710,N_609,N_667);
nor U711 (N_711,N_603,N_613);
or U712 (N_712,N_666,N_669);
nand U713 (N_713,N_612,N_613);
nor U714 (N_714,N_612,N_611);
xnor U715 (N_715,N_643,N_623);
xnor U716 (N_716,N_627,N_602);
or U717 (N_717,N_604,N_673);
nor U718 (N_718,N_634,N_623);
and U719 (N_719,N_612,N_674);
nor U720 (N_720,N_609,N_631);
nor U721 (N_721,N_606,N_647);
and U722 (N_722,N_627,N_606);
nand U723 (N_723,N_647,N_646);
nand U724 (N_724,N_611,N_670);
nor U725 (N_725,N_647,N_674);
and U726 (N_726,N_651,N_622);
or U727 (N_727,N_662,N_646);
or U728 (N_728,N_600,N_605);
nor U729 (N_729,N_645,N_620);
nor U730 (N_730,N_647,N_664);
nand U731 (N_731,N_619,N_623);
or U732 (N_732,N_609,N_674);
nand U733 (N_733,N_614,N_674);
nor U734 (N_734,N_638,N_600);
nand U735 (N_735,N_648,N_605);
or U736 (N_736,N_674,N_606);
or U737 (N_737,N_629,N_673);
nor U738 (N_738,N_642,N_654);
nor U739 (N_739,N_646,N_624);
and U740 (N_740,N_620,N_624);
nor U741 (N_741,N_664,N_623);
or U742 (N_742,N_604,N_652);
nand U743 (N_743,N_629,N_605);
and U744 (N_744,N_660,N_613);
xor U745 (N_745,N_665,N_666);
nor U746 (N_746,N_662,N_600);
and U747 (N_747,N_611,N_640);
xor U748 (N_748,N_653,N_645);
nand U749 (N_749,N_608,N_651);
and U750 (N_750,N_680,N_719);
nor U751 (N_751,N_691,N_714);
xor U752 (N_752,N_699,N_711);
nor U753 (N_753,N_721,N_694);
and U754 (N_754,N_685,N_677);
nor U755 (N_755,N_712,N_749);
nor U756 (N_756,N_684,N_705);
or U757 (N_757,N_713,N_725);
or U758 (N_758,N_703,N_730);
or U759 (N_759,N_746,N_718);
and U760 (N_760,N_698,N_744);
nor U761 (N_761,N_738,N_731);
or U762 (N_762,N_697,N_748);
xnor U763 (N_763,N_720,N_689);
and U764 (N_764,N_681,N_737);
nand U765 (N_765,N_726,N_693);
xor U766 (N_766,N_715,N_722);
and U767 (N_767,N_696,N_727);
nor U768 (N_768,N_692,N_716);
and U769 (N_769,N_717,N_723);
nand U770 (N_770,N_676,N_701);
or U771 (N_771,N_743,N_735);
nand U772 (N_772,N_740,N_739);
nand U773 (N_773,N_736,N_729);
or U774 (N_774,N_742,N_687);
and U775 (N_775,N_690,N_682);
nor U776 (N_776,N_695,N_747);
xnor U777 (N_777,N_708,N_732);
or U778 (N_778,N_728,N_686);
nor U779 (N_779,N_678,N_679);
xnor U780 (N_780,N_724,N_704);
nand U781 (N_781,N_675,N_688);
nor U782 (N_782,N_683,N_734);
and U783 (N_783,N_709,N_741);
and U784 (N_784,N_700,N_745);
or U785 (N_785,N_733,N_702);
nor U786 (N_786,N_706,N_707);
nand U787 (N_787,N_710,N_697);
or U788 (N_788,N_740,N_722);
nand U789 (N_789,N_695,N_743);
or U790 (N_790,N_732,N_693);
and U791 (N_791,N_684,N_715);
nor U792 (N_792,N_728,N_707);
and U793 (N_793,N_728,N_692);
xor U794 (N_794,N_682,N_681);
nand U795 (N_795,N_681,N_707);
or U796 (N_796,N_685,N_696);
and U797 (N_797,N_747,N_739);
nor U798 (N_798,N_684,N_749);
or U799 (N_799,N_698,N_689);
and U800 (N_800,N_726,N_680);
nand U801 (N_801,N_728,N_719);
nor U802 (N_802,N_691,N_725);
or U803 (N_803,N_737,N_698);
or U804 (N_804,N_718,N_698);
xor U805 (N_805,N_688,N_677);
and U806 (N_806,N_698,N_743);
or U807 (N_807,N_706,N_728);
and U808 (N_808,N_714,N_727);
or U809 (N_809,N_747,N_676);
nand U810 (N_810,N_676,N_736);
nand U811 (N_811,N_723,N_696);
and U812 (N_812,N_692,N_715);
xnor U813 (N_813,N_745,N_693);
nor U814 (N_814,N_741,N_689);
nor U815 (N_815,N_677,N_687);
nor U816 (N_816,N_693,N_742);
or U817 (N_817,N_731,N_709);
nor U818 (N_818,N_676,N_702);
nor U819 (N_819,N_737,N_746);
nand U820 (N_820,N_693,N_702);
and U821 (N_821,N_706,N_719);
xnor U822 (N_822,N_687,N_733);
or U823 (N_823,N_723,N_677);
and U824 (N_824,N_697,N_706);
or U825 (N_825,N_819,N_786);
or U826 (N_826,N_777,N_792);
or U827 (N_827,N_762,N_765);
or U828 (N_828,N_764,N_783);
and U829 (N_829,N_784,N_778);
nor U830 (N_830,N_769,N_823);
and U831 (N_831,N_815,N_755);
xor U832 (N_832,N_756,N_788);
nor U833 (N_833,N_809,N_757);
nor U834 (N_834,N_816,N_806);
and U835 (N_835,N_814,N_802);
and U836 (N_836,N_754,N_775);
and U837 (N_837,N_770,N_800);
nand U838 (N_838,N_774,N_807);
and U839 (N_839,N_812,N_752);
nor U840 (N_840,N_798,N_797);
nand U841 (N_841,N_795,N_791);
and U842 (N_842,N_790,N_780);
nor U843 (N_843,N_753,N_804);
xnor U844 (N_844,N_782,N_811);
and U845 (N_845,N_779,N_801);
and U846 (N_846,N_805,N_789);
xnor U847 (N_847,N_771,N_759);
nor U848 (N_848,N_768,N_776);
or U849 (N_849,N_758,N_793);
or U850 (N_850,N_767,N_817);
nor U851 (N_851,N_821,N_824);
and U852 (N_852,N_781,N_772);
and U853 (N_853,N_803,N_763);
or U854 (N_854,N_750,N_822);
nand U855 (N_855,N_766,N_760);
nor U856 (N_856,N_794,N_787);
nand U857 (N_857,N_808,N_818);
xor U858 (N_858,N_773,N_785);
nand U859 (N_859,N_796,N_820);
nand U860 (N_860,N_799,N_813);
or U861 (N_861,N_751,N_761);
and U862 (N_862,N_810,N_773);
and U863 (N_863,N_782,N_787);
nor U864 (N_864,N_812,N_800);
nor U865 (N_865,N_808,N_777);
or U866 (N_866,N_795,N_751);
nand U867 (N_867,N_784,N_819);
nor U868 (N_868,N_815,N_782);
or U869 (N_869,N_766,N_762);
or U870 (N_870,N_756,N_814);
nand U871 (N_871,N_811,N_820);
nand U872 (N_872,N_774,N_795);
or U873 (N_873,N_765,N_784);
nor U874 (N_874,N_777,N_762);
nand U875 (N_875,N_809,N_783);
nor U876 (N_876,N_817,N_775);
or U877 (N_877,N_788,N_762);
or U878 (N_878,N_805,N_824);
and U879 (N_879,N_754,N_793);
and U880 (N_880,N_751,N_812);
nand U881 (N_881,N_799,N_824);
nor U882 (N_882,N_813,N_816);
or U883 (N_883,N_754,N_819);
xor U884 (N_884,N_800,N_753);
nor U885 (N_885,N_750,N_810);
nand U886 (N_886,N_801,N_793);
nor U887 (N_887,N_820,N_764);
and U888 (N_888,N_823,N_772);
nand U889 (N_889,N_771,N_791);
and U890 (N_890,N_822,N_803);
nor U891 (N_891,N_756,N_817);
or U892 (N_892,N_772,N_753);
and U893 (N_893,N_750,N_778);
nand U894 (N_894,N_810,N_790);
or U895 (N_895,N_774,N_789);
or U896 (N_896,N_811,N_823);
nand U897 (N_897,N_790,N_789);
or U898 (N_898,N_810,N_793);
and U899 (N_899,N_779,N_752);
or U900 (N_900,N_859,N_849);
xnor U901 (N_901,N_834,N_829);
nand U902 (N_902,N_847,N_830);
nand U903 (N_903,N_882,N_858);
and U904 (N_904,N_879,N_877);
nand U905 (N_905,N_896,N_840);
xnor U906 (N_906,N_872,N_851);
xor U907 (N_907,N_832,N_899);
or U908 (N_908,N_890,N_897);
and U909 (N_909,N_876,N_871);
xnor U910 (N_910,N_836,N_831);
nand U911 (N_911,N_898,N_850);
nor U912 (N_912,N_865,N_895);
and U913 (N_913,N_846,N_827);
nand U914 (N_914,N_874,N_860);
nand U915 (N_915,N_894,N_825);
and U916 (N_916,N_854,N_828);
nand U917 (N_917,N_843,N_891);
or U918 (N_918,N_856,N_844);
nor U919 (N_919,N_833,N_867);
and U920 (N_920,N_863,N_878);
nand U921 (N_921,N_857,N_861);
xnor U922 (N_922,N_862,N_873);
and U923 (N_923,N_881,N_887);
or U924 (N_924,N_842,N_837);
and U925 (N_925,N_884,N_893);
nor U926 (N_926,N_880,N_826);
and U927 (N_927,N_853,N_875);
and U928 (N_928,N_883,N_864);
or U929 (N_929,N_841,N_845);
xnor U930 (N_930,N_888,N_838);
nor U931 (N_931,N_839,N_848);
nor U932 (N_932,N_835,N_892);
or U933 (N_933,N_868,N_869);
xor U934 (N_934,N_870,N_886);
or U935 (N_935,N_889,N_885);
nand U936 (N_936,N_855,N_852);
and U937 (N_937,N_866,N_842);
nand U938 (N_938,N_867,N_872);
or U939 (N_939,N_831,N_859);
nand U940 (N_940,N_894,N_835);
xor U941 (N_941,N_850,N_881);
or U942 (N_942,N_877,N_833);
nor U943 (N_943,N_843,N_845);
or U944 (N_944,N_836,N_878);
nor U945 (N_945,N_878,N_825);
xor U946 (N_946,N_844,N_837);
nand U947 (N_947,N_856,N_866);
nor U948 (N_948,N_830,N_851);
or U949 (N_949,N_885,N_878);
or U950 (N_950,N_836,N_869);
nor U951 (N_951,N_853,N_876);
nand U952 (N_952,N_864,N_839);
or U953 (N_953,N_872,N_827);
xnor U954 (N_954,N_868,N_886);
and U955 (N_955,N_842,N_881);
xor U956 (N_956,N_839,N_899);
and U957 (N_957,N_832,N_842);
or U958 (N_958,N_860,N_825);
or U959 (N_959,N_863,N_852);
nor U960 (N_960,N_849,N_857);
nand U961 (N_961,N_885,N_834);
or U962 (N_962,N_886,N_853);
and U963 (N_963,N_888,N_882);
or U964 (N_964,N_840,N_876);
and U965 (N_965,N_892,N_877);
nand U966 (N_966,N_890,N_860);
nor U967 (N_967,N_856,N_841);
nor U968 (N_968,N_888,N_853);
and U969 (N_969,N_832,N_841);
and U970 (N_970,N_833,N_857);
xor U971 (N_971,N_841,N_880);
or U972 (N_972,N_838,N_833);
and U973 (N_973,N_883,N_842);
xor U974 (N_974,N_864,N_875);
and U975 (N_975,N_901,N_956);
and U976 (N_976,N_928,N_900);
and U977 (N_977,N_902,N_962);
or U978 (N_978,N_961,N_937);
or U979 (N_979,N_904,N_929);
nor U980 (N_980,N_939,N_959);
and U981 (N_981,N_965,N_963);
or U982 (N_982,N_971,N_923);
or U983 (N_983,N_930,N_953);
or U984 (N_984,N_916,N_908);
and U985 (N_985,N_950,N_915);
nor U986 (N_986,N_967,N_960);
nand U987 (N_987,N_921,N_958);
nand U988 (N_988,N_934,N_947);
or U989 (N_989,N_913,N_942);
nand U990 (N_990,N_938,N_935);
xor U991 (N_991,N_907,N_931);
nor U992 (N_992,N_919,N_924);
xor U993 (N_993,N_945,N_951);
xor U994 (N_994,N_926,N_910);
nor U995 (N_995,N_973,N_969);
and U996 (N_996,N_909,N_972);
or U997 (N_997,N_920,N_917);
or U998 (N_998,N_912,N_911);
nand U999 (N_999,N_954,N_914);
nor U1000 (N_1000,N_966,N_943);
and U1001 (N_1001,N_932,N_940);
nand U1002 (N_1002,N_903,N_970);
or U1003 (N_1003,N_905,N_974);
nor U1004 (N_1004,N_933,N_936);
nor U1005 (N_1005,N_944,N_925);
and U1006 (N_1006,N_964,N_957);
or U1007 (N_1007,N_927,N_955);
xnor U1008 (N_1008,N_946,N_968);
and U1009 (N_1009,N_922,N_941);
or U1010 (N_1010,N_948,N_949);
nor U1011 (N_1011,N_952,N_918);
nand U1012 (N_1012,N_906,N_911);
and U1013 (N_1013,N_912,N_952);
xnor U1014 (N_1014,N_955,N_962);
or U1015 (N_1015,N_938,N_906);
or U1016 (N_1016,N_906,N_952);
nand U1017 (N_1017,N_954,N_949);
and U1018 (N_1018,N_916,N_970);
and U1019 (N_1019,N_950,N_922);
xor U1020 (N_1020,N_967,N_903);
nor U1021 (N_1021,N_961,N_918);
and U1022 (N_1022,N_957,N_939);
and U1023 (N_1023,N_926,N_942);
or U1024 (N_1024,N_956,N_927);
nand U1025 (N_1025,N_901,N_967);
nand U1026 (N_1026,N_940,N_947);
or U1027 (N_1027,N_954,N_972);
nand U1028 (N_1028,N_936,N_929);
nor U1029 (N_1029,N_970,N_907);
xor U1030 (N_1030,N_962,N_972);
nand U1031 (N_1031,N_961,N_928);
and U1032 (N_1032,N_963,N_904);
and U1033 (N_1033,N_952,N_934);
nand U1034 (N_1034,N_969,N_950);
or U1035 (N_1035,N_905,N_960);
nor U1036 (N_1036,N_949,N_931);
and U1037 (N_1037,N_903,N_922);
nand U1038 (N_1038,N_946,N_911);
nand U1039 (N_1039,N_925,N_914);
and U1040 (N_1040,N_943,N_951);
and U1041 (N_1041,N_959,N_935);
and U1042 (N_1042,N_943,N_941);
nand U1043 (N_1043,N_908,N_973);
nand U1044 (N_1044,N_936,N_952);
or U1045 (N_1045,N_911,N_963);
nor U1046 (N_1046,N_964,N_962);
and U1047 (N_1047,N_968,N_943);
nor U1048 (N_1048,N_901,N_922);
or U1049 (N_1049,N_912,N_921);
nor U1050 (N_1050,N_999,N_982);
xor U1051 (N_1051,N_979,N_1032);
and U1052 (N_1052,N_1012,N_1004);
nor U1053 (N_1053,N_1047,N_992);
and U1054 (N_1054,N_1007,N_985);
and U1055 (N_1055,N_1046,N_1011);
xnor U1056 (N_1056,N_980,N_1006);
nor U1057 (N_1057,N_998,N_991);
nand U1058 (N_1058,N_1029,N_975);
nand U1059 (N_1059,N_1038,N_977);
xor U1060 (N_1060,N_984,N_1010);
nor U1061 (N_1061,N_1036,N_1033);
nand U1062 (N_1062,N_1017,N_1044);
nor U1063 (N_1063,N_1031,N_1002);
and U1064 (N_1064,N_990,N_993);
xnor U1065 (N_1065,N_1030,N_1049);
or U1066 (N_1066,N_1015,N_1026);
and U1067 (N_1067,N_1037,N_1014);
nand U1068 (N_1068,N_1025,N_987);
and U1069 (N_1069,N_1021,N_1040);
nand U1070 (N_1070,N_988,N_1041);
nand U1071 (N_1071,N_1016,N_1009);
or U1072 (N_1072,N_996,N_986);
or U1073 (N_1073,N_1023,N_1039);
nand U1074 (N_1074,N_976,N_1000);
nand U1075 (N_1075,N_1018,N_994);
and U1076 (N_1076,N_1008,N_1048);
nand U1077 (N_1077,N_1042,N_1020);
or U1078 (N_1078,N_989,N_1019);
or U1079 (N_1079,N_1045,N_1001);
and U1080 (N_1080,N_1005,N_1013);
nand U1081 (N_1081,N_1043,N_981);
and U1082 (N_1082,N_995,N_1028);
nand U1083 (N_1083,N_978,N_997);
nor U1084 (N_1084,N_1035,N_983);
nand U1085 (N_1085,N_1024,N_1034);
nor U1086 (N_1086,N_1003,N_1022);
nand U1087 (N_1087,N_1027,N_1012);
and U1088 (N_1088,N_1016,N_1012);
nand U1089 (N_1089,N_1027,N_1035);
or U1090 (N_1090,N_977,N_1003);
or U1091 (N_1091,N_1027,N_984);
or U1092 (N_1092,N_1010,N_996);
nor U1093 (N_1093,N_1026,N_1039);
nor U1094 (N_1094,N_1049,N_1022);
nand U1095 (N_1095,N_1003,N_1027);
and U1096 (N_1096,N_1023,N_1014);
nand U1097 (N_1097,N_994,N_1031);
and U1098 (N_1098,N_1002,N_1018);
nand U1099 (N_1099,N_1046,N_1039);
nand U1100 (N_1100,N_1040,N_1002);
and U1101 (N_1101,N_1024,N_1000);
nor U1102 (N_1102,N_1042,N_990);
nand U1103 (N_1103,N_983,N_1023);
nand U1104 (N_1104,N_988,N_1006);
or U1105 (N_1105,N_997,N_1025);
or U1106 (N_1106,N_1003,N_1010);
or U1107 (N_1107,N_1006,N_1046);
nor U1108 (N_1108,N_1041,N_1020);
and U1109 (N_1109,N_1010,N_987);
and U1110 (N_1110,N_994,N_1044);
or U1111 (N_1111,N_1009,N_1027);
or U1112 (N_1112,N_993,N_1011);
or U1113 (N_1113,N_997,N_1038);
nor U1114 (N_1114,N_1011,N_1040);
or U1115 (N_1115,N_1008,N_1012);
nor U1116 (N_1116,N_989,N_1002);
or U1117 (N_1117,N_995,N_1037);
nor U1118 (N_1118,N_1001,N_1039);
or U1119 (N_1119,N_989,N_976);
and U1120 (N_1120,N_982,N_1021);
and U1121 (N_1121,N_982,N_995);
and U1122 (N_1122,N_977,N_986);
nor U1123 (N_1123,N_1011,N_1018);
nor U1124 (N_1124,N_1041,N_1022);
nor U1125 (N_1125,N_1052,N_1091);
and U1126 (N_1126,N_1103,N_1053);
or U1127 (N_1127,N_1065,N_1063);
or U1128 (N_1128,N_1113,N_1092);
nand U1129 (N_1129,N_1111,N_1054);
nand U1130 (N_1130,N_1115,N_1074);
xnor U1131 (N_1131,N_1089,N_1059);
xor U1132 (N_1132,N_1110,N_1116);
nand U1133 (N_1133,N_1075,N_1077);
xor U1134 (N_1134,N_1076,N_1096);
nand U1135 (N_1135,N_1057,N_1108);
or U1136 (N_1136,N_1121,N_1093);
nor U1137 (N_1137,N_1112,N_1073);
and U1138 (N_1138,N_1123,N_1080);
nand U1139 (N_1139,N_1070,N_1101);
and U1140 (N_1140,N_1068,N_1055);
or U1141 (N_1141,N_1124,N_1106);
or U1142 (N_1142,N_1086,N_1083);
nand U1143 (N_1143,N_1072,N_1117);
or U1144 (N_1144,N_1097,N_1079);
or U1145 (N_1145,N_1104,N_1102);
or U1146 (N_1146,N_1060,N_1058);
or U1147 (N_1147,N_1095,N_1098);
and U1148 (N_1148,N_1107,N_1081);
nand U1149 (N_1149,N_1120,N_1114);
or U1150 (N_1150,N_1056,N_1094);
nand U1151 (N_1151,N_1078,N_1071);
or U1152 (N_1152,N_1105,N_1082);
xor U1153 (N_1153,N_1069,N_1087);
nand U1154 (N_1154,N_1119,N_1064);
or U1155 (N_1155,N_1067,N_1122);
nor U1156 (N_1156,N_1109,N_1066);
or U1157 (N_1157,N_1088,N_1099);
nand U1158 (N_1158,N_1084,N_1090);
nor U1159 (N_1159,N_1051,N_1062);
nand U1160 (N_1160,N_1050,N_1118);
and U1161 (N_1161,N_1085,N_1100);
or U1162 (N_1162,N_1061,N_1070);
or U1163 (N_1163,N_1062,N_1089);
or U1164 (N_1164,N_1124,N_1117);
xor U1165 (N_1165,N_1111,N_1123);
or U1166 (N_1166,N_1074,N_1050);
nand U1167 (N_1167,N_1050,N_1096);
or U1168 (N_1168,N_1082,N_1118);
or U1169 (N_1169,N_1106,N_1098);
nand U1170 (N_1170,N_1095,N_1078);
xor U1171 (N_1171,N_1084,N_1101);
or U1172 (N_1172,N_1073,N_1075);
xor U1173 (N_1173,N_1059,N_1083);
nor U1174 (N_1174,N_1090,N_1120);
nand U1175 (N_1175,N_1124,N_1080);
nor U1176 (N_1176,N_1067,N_1104);
nor U1177 (N_1177,N_1093,N_1064);
and U1178 (N_1178,N_1119,N_1118);
and U1179 (N_1179,N_1063,N_1082);
or U1180 (N_1180,N_1061,N_1082);
or U1181 (N_1181,N_1107,N_1124);
and U1182 (N_1182,N_1082,N_1094);
nand U1183 (N_1183,N_1055,N_1099);
xnor U1184 (N_1184,N_1096,N_1118);
nand U1185 (N_1185,N_1105,N_1114);
and U1186 (N_1186,N_1102,N_1071);
nor U1187 (N_1187,N_1068,N_1073);
and U1188 (N_1188,N_1119,N_1075);
or U1189 (N_1189,N_1088,N_1118);
nand U1190 (N_1190,N_1072,N_1053);
nand U1191 (N_1191,N_1081,N_1093);
nor U1192 (N_1192,N_1112,N_1080);
nand U1193 (N_1193,N_1085,N_1104);
xor U1194 (N_1194,N_1074,N_1097);
and U1195 (N_1195,N_1053,N_1058);
nand U1196 (N_1196,N_1063,N_1076);
nor U1197 (N_1197,N_1101,N_1104);
or U1198 (N_1198,N_1051,N_1083);
and U1199 (N_1199,N_1080,N_1059);
nand U1200 (N_1200,N_1141,N_1152);
or U1201 (N_1201,N_1166,N_1161);
and U1202 (N_1202,N_1192,N_1165);
and U1203 (N_1203,N_1169,N_1135);
and U1204 (N_1204,N_1175,N_1183);
nor U1205 (N_1205,N_1140,N_1196);
and U1206 (N_1206,N_1129,N_1139);
or U1207 (N_1207,N_1145,N_1127);
or U1208 (N_1208,N_1193,N_1146);
nor U1209 (N_1209,N_1194,N_1187);
nor U1210 (N_1210,N_1134,N_1197);
nor U1211 (N_1211,N_1163,N_1190);
nor U1212 (N_1212,N_1156,N_1186);
and U1213 (N_1213,N_1151,N_1199);
nor U1214 (N_1214,N_1126,N_1136);
or U1215 (N_1215,N_1144,N_1150);
nor U1216 (N_1216,N_1185,N_1176);
nor U1217 (N_1217,N_1189,N_1180);
nor U1218 (N_1218,N_1154,N_1198);
nor U1219 (N_1219,N_1137,N_1160);
nand U1220 (N_1220,N_1188,N_1174);
nand U1221 (N_1221,N_1131,N_1179);
nor U1222 (N_1222,N_1159,N_1178);
nand U1223 (N_1223,N_1191,N_1167);
and U1224 (N_1224,N_1158,N_1132);
or U1225 (N_1225,N_1125,N_1173);
nand U1226 (N_1226,N_1170,N_1171);
nor U1227 (N_1227,N_1128,N_1142);
or U1228 (N_1228,N_1148,N_1138);
nand U1229 (N_1229,N_1195,N_1162);
xor U1230 (N_1230,N_1164,N_1184);
nor U1231 (N_1231,N_1149,N_1172);
nand U1232 (N_1232,N_1147,N_1168);
nand U1233 (N_1233,N_1182,N_1133);
nand U1234 (N_1234,N_1181,N_1153);
nor U1235 (N_1235,N_1177,N_1155);
or U1236 (N_1236,N_1157,N_1130);
nor U1237 (N_1237,N_1143,N_1167);
xnor U1238 (N_1238,N_1168,N_1146);
nand U1239 (N_1239,N_1129,N_1144);
nor U1240 (N_1240,N_1186,N_1153);
or U1241 (N_1241,N_1126,N_1141);
nor U1242 (N_1242,N_1140,N_1174);
nand U1243 (N_1243,N_1130,N_1199);
or U1244 (N_1244,N_1172,N_1134);
or U1245 (N_1245,N_1129,N_1198);
and U1246 (N_1246,N_1196,N_1192);
or U1247 (N_1247,N_1136,N_1180);
nand U1248 (N_1248,N_1174,N_1195);
nor U1249 (N_1249,N_1142,N_1144);
and U1250 (N_1250,N_1179,N_1162);
and U1251 (N_1251,N_1165,N_1145);
xnor U1252 (N_1252,N_1160,N_1177);
or U1253 (N_1253,N_1138,N_1188);
xor U1254 (N_1254,N_1130,N_1179);
xnor U1255 (N_1255,N_1137,N_1189);
or U1256 (N_1256,N_1146,N_1182);
or U1257 (N_1257,N_1144,N_1166);
or U1258 (N_1258,N_1190,N_1149);
nand U1259 (N_1259,N_1185,N_1179);
nor U1260 (N_1260,N_1198,N_1127);
nand U1261 (N_1261,N_1156,N_1132);
or U1262 (N_1262,N_1154,N_1180);
and U1263 (N_1263,N_1142,N_1195);
nor U1264 (N_1264,N_1172,N_1177);
or U1265 (N_1265,N_1174,N_1171);
nor U1266 (N_1266,N_1134,N_1176);
or U1267 (N_1267,N_1160,N_1130);
xnor U1268 (N_1268,N_1173,N_1136);
and U1269 (N_1269,N_1185,N_1192);
nand U1270 (N_1270,N_1146,N_1133);
and U1271 (N_1271,N_1154,N_1196);
nor U1272 (N_1272,N_1135,N_1151);
nand U1273 (N_1273,N_1197,N_1177);
nor U1274 (N_1274,N_1196,N_1178);
nor U1275 (N_1275,N_1264,N_1200);
nand U1276 (N_1276,N_1258,N_1249);
and U1277 (N_1277,N_1207,N_1231);
and U1278 (N_1278,N_1205,N_1263);
nor U1279 (N_1279,N_1252,N_1206);
nor U1280 (N_1280,N_1255,N_1238);
nand U1281 (N_1281,N_1244,N_1219);
and U1282 (N_1282,N_1271,N_1209);
and U1283 (N_1283,N_1236,N_1226);
nor U1284 (N_1284,N_1246,N_1218);
nand U1285 (N_1285,N_1228,N_1202);
nand U1286 (N_1286,N_1247,N_1245);
and U1287 (N_1287,N_1230,N_1217);
or U1288 (N_1288,N_1274,N_1229);
nor U1289 (N_1289,N_1260,N_1239);
nor U1290 (N_1290,N_1233,N_1232);
and U1291 (N_1291,N_1216,N_1273);
nor U1292 (N_1292,N_1267,N_1211);
nand U1293 (N_1293,N_1254,N_1268);
xor U1294 (N_1294,N_1248,N_1262);
nor U1295 (N_1295,N_1220,N_1235);
nor U1296 (N_1296,N_1215,N_1210);
or U1297 (N_1297,N_1266,N_1223);
and U1298 (N_1298,N_1225,N_1214);
or U1299 (N_1299,N_1250,N_1221);
nand U1300 (N_1300,N_1269,N_1212);
nand U1301 (N_1301,N_1234,N_1204);
nor U1302 (N_1302,N_1208,N_1242);
and U1303 (N_1303,N_1259,N_1251);
and U1304 (N_1304,N_1257,N_1240);
nor U1305 (N_1305,N_1222,N_1270);
and U1306 (N_1306,N_1237,N_1253);
or U1307 (N_1307,N_1203,N_1261);
or U1308 (N_1308,N_1213,N_1201);
and U1309 (N_1309,N_1265,N_1227);
or U1310 (N_1310,N_1243,N_1241);
nand U1311 (N_1311,N_1256,N_1224);
or U1312 (N_1312,N_1272,N_1203);
and U1313 (N_1313,N_1209,N_1217);
and U1314 (N_1314,N_1201,N_1208);
nor U1315 (N_1315,N_1211,N_1204);
or U1316 (N_1316,N_1229,N_1236);
nand U1317 (N_1317,N_1268,N_1219);
and U1318 (N_1318,N_1222,N_1267);
nand U1319 (N_1319,N_1232,N_1217);
nor U1320 (N_1320,N_1223,N_1247);
and U1321 (N_1321,N_1230,N_1246);
and U1322 (N_1322,N_1219,N_1247);
nor U1323 (N_1323,N_1242,N_1262);
and U1324 (N_1324,N_1263,N_1208);
nand U1325 (N_1325,N_1271,N_1265);
nor U1326 (N_1326,N_1212,N_1244);
nand U1327 (N_1327,N_1224,N_1217);
or U1328 (N_1328,N_1230,N_1204);
nand U1329 (N_1329,N_1210,N_1224);
or U1330 (N_1330,N_1201,N_1263);
nor U1331 (N_1331,N_1209,N_1225);
or U1332 (N_1332,N_1226,N_1239);
and U1333 (N_1333,N_1265,N_1232);
and U1334 (N_1334,N_1238,N_1233);
and U1335 (N_1335,N_1210,N_1238);
xor U1336 (N_1336,N_1234,N_1270);
nand U1337 (N_1337,N_1246,N_1213);
xor U1338 (N_1338,N_1226,N_1235);
or U1339 (N_1339,N_1234,N_1265);
xor U1340 (N_1340,N_1224,N_1245);
and U1341 (N_1341,N_1204,N_1208);
nor U1342 (N_1342,N_1251,N_1212);
xor U1343 (N_1343,N_1217,N_1220);
or U1344 (N_1344,N_1229,N_1210);
xor U1345 (N_1345,N_1223,N_1271);
nor U1346 (N_1346,N_1201,N_1251);
nor U1347 (N_1347,N_1237,N_1274);
xor U1348 (N_1348,N_1274,N_1262);
nand U1349 (N_1349,N_1243,N_1256);
and U1350 (N_1350,N_1345,N_1280);
nor U1351 (N_1351,N_1306,N_1342);
and U1352 (N_1352,N_1287,N_1285);
xor U1353 (N_1353,N_1318,N_1294);
and U1354 (N_1354,N_1347,N_1275);
and U1355 (N_1355,N_1321,N_1293);
nand U1356 (N_1356,N_1320,N_1283);
nand U1357 (N_1357,N_1307,N_1301);
nor U1358 (N_1358,N_1302,N_1316);
nor U1359 (N_1359,N_1346,N_1289);
nand U1360 (N_1360,N_1343,N_1281);
or U1361 (N_1361,N_1326,N_1295);
nand U1362 (N_1362,N_1291,N_1311);
xnor U1363 (N_1363,N_1296,N_1310);
and U1364 (N_1364,N_1284,N_1331);
nor U1365 (N_1365,N_1292,N_1344);
xor U1366 (N_1366,N_1334,N_1314);
and U1367 (N_1367,N_1325,N_1317);
nand U1368 (N_1368,N_1323,N_1312);
nand U1369 (N_1369,N_1337,N_1299);
nor U1370 (N_1370,N_1304,N_1297);
or U1371 (N_1371,N_1328,N_1298);
and U1372 (N_1372,N_1290,N_1348);
xnor U1373 (N_1373,N_1340,N_1279);
nor U1374 (N_1374,N_1305,N_1308);
xnor U1375 (N_1375,N_1277,N_1324);
nor U1376 (N_1376,N_1336,N_1332);
and U1377 (N_1377,N_1278,N_1303);
or U1378 (N_1378,N_1276,N_1282);
xnor U1379 (N_1379,N_1322,N_1338);
nor U1380 (N_1380,N_1335,N_1330);
xnor U1381 (N_1381,N_1315,N_1327);
or U1382 (N_1382,N_1349,N_1288);
and U1383 (N_1383,N_1309,N_1319);
nor U1384 (N_1384,N_1339,N_1300);
and U1385 (N_1385,N_1313,N_1286);
nor U1386 (N_1386,N_1333,N_1329);
nand U1387 (N_1387,N_1341,N_1312);
nand U1388 (N_1388,N_1329,N_1294);
nor U1389 (N_1389,N_1334,N_1326);
and U1390 (N_1390,N_1291,N_1313);
or U1391 (N_1391,N_1298,N_1315);
and U1392 (N_1392,N_1317,N_1291);
or U1393 (N_1393,N_1277,N_1310);
nor U1394 (N_1394,N_1322,N_1326);
and U1395 (N_1395,N_1317,N_1321);
or U1396 (N_1396,N_1275,N_1310);
and U1397 (N_1397,N_1302,N_1292);
xor U1398 (N_1398,N_1319,N_1341);
nand U1399 (N_1399,N_1281,N_1292);
nand U1400 (N_1400,N_1324,N_1339);
nor U1401 (N_1401,N_1307,N_1337);
nor U1402 (N_1402,N_1320,N_1338);
nor U1403 (N_1403,N_1307,N_1298);
or U1404 (N_1404,N_1307,N_1323);
nand U1405 (N_1405,N_1296,N_1300);
and U1406 (N_1406,N_1324,N_1293);
or U1407 (N_1407,N_1302,N_1278);
nor U1408 (N_1408,N_1278,N_1344);
xor U1409 (N_1409,N_1329,N_1288);
nand U1410 (N_1410,N_1295,N_1338);
or U1411 (N_1411,N_1306,N_1309);
nor U1412 (N_1412,N_1293,N_1278);
or U1413 (N_1413,N_1317,N_1313);
nor U1414 (N_1414,N_1343,N_1313);
nor U1415 (N_1415,N_1295,N_1299);
nand U1416 (N_1416,N_1343,N_1329);
xnor U1417 (N_1417,N_1332,N_1284);
or U1418 (N_1418,N_1283,N_1335);
or U1419 (N_1419,N_1276,N_1301);
nor U1420 (N_1420,N_1323,N_1294);
nor U1421 (N_1421,N_1336,N_1291);
nand U1422 (N_1422,N_1332,N_1277);
nand U1423 (N_1423,N_1318,N_1344);
or U1424 (N_1424,N_1294,N_1342);
or U1425 (N_1425,N_1381,N_1350);
nand U1426 (N_1426,N_1357,N_1368);
xnor U1427 (N_1427,N_1418,N_1402);
nand U1428 (N_1428,N_1355,N_1392);
nor U1429 (N_1429,N_1395,N_1384);
nor U1430 (N_1430,N_1380,N_1421);
nand U1431 (N_1431,N_1417,N_1351);
nor U1432 (N_1432,N_1416,N_1364);
or U1433 (N_1433,N_1404,N_1397);
nand U1434 (N_1434,N_1391,N_1377);
and U1435 (N_1435,N_1373,N_1385);
nor U1436 (N_1436,N_1401,N_1394);
nor U1437 (N_1437,N_1424,N_1360);
nand U1438 (N_1438,N_1396,N_1409);
xnor U1439 (N_1439,N_1354,N_1359);
or U1440 (N_1440,N_1387,N_1362);
nand U1441 (N_1441,N_1410,N_1412);
nor U1442 (N_1442,N_1419,N_1376);
nand U1443 (N_1443,N_1408,N_1388);
nor U1444 (N_1444,N_1420,N_1400);
or U1445 (N_1445,N_1413,N_1358);
and U1446 (N_1446,N_1423,N_1411);
nand U1447 (N_1447,N_1399,N_1407);
nor U1448 (N_1448,N_1386,N_1414);
nand U1449 (N_1449,N_1422,N_1403);
nor U1450 (N_1450,N_1361,N_1371);
or U1451 (N_1451,N_1366,N_1389);
nand U1452 (N_1452,N_1406,N_1370);
nor U1453 (N_1453,N_1405,N_1379);
and U1454 (N_1454,N_1375,N_1393);
nand U1455 (N_1455,N_1415,N_1352);
nor U1456 (N_1456,N_1367,N_1372);
or U1457 (N_1457,N_1378,N_1363);
nand U1458 (N_1458,N_1369,N_1398);
or U1459 (N_1459,N_1383,N_1353);
nand U1460 (N_1460,N_1356,N_1382);
xnor U1461 (N_1461,N_1390,N_1365);
xor U1462 (N_1462,N_1374,N_1372);
nand U1463 (N_1463,N_1390,N_1361);
nand U1464 (N_1464,N_1362,N_1356);
and U1465 (N_1465,N_1380,N_1409);
nor U1466 (N_1466,N_1360,N_1366);
and U1467 (N_1467,N_1414,N_1373);
nand U1468 (N_1468,N_1409,N_1394);
nand U1469 (N_1469,N_1405,N_1376);
and U1470 (N_1470,N_1373,N_1352);
and U1471 (N_1471,N_1373,N_1424);
nor U1472 (N_1472,N_1416,N_1360);
and U1473 (N_1473,N_1388,N_1366);
nor U1474 (N_1474,N_1405,N_1403);
xor U1475 (N_1475,N_1396,N_1387);
nor U1476 (N_1476,N_1406,N_1399);
or U1477 (N_1477,N_1379,N_1370);
nand U1478 (N_1478,N_1422,N_1389);
or U1479 (N_1479,N_1400,N_1414);
nor U1480 (N_1480,N_1352,N_1396);
and U1481 (N_1481,N_1359,N_1419);
nor U1482 (N_1482,N_1350,N_1411);
nand U1483 (N_1483,N_1373,N_1405);
nand U1484 (N_1484,N_1409,N_1413);
or U1485 (N_1485,N_1396,N_1353);
nand U1486 (N_1486,N_1357,N_1404);
nand U1487 (N_1487,N_1373,N_1366);
nor U1488 (N_1488,N_1352,N_1416);
nor U1489 (N_1489,N_1402,N_1411);
nand U1490 (N_1490,N_1409,N_1414);
nor U1491 (N_1491,N_1367,N_1424);
and U1492 (N_1492,N_1383,N_1412);
xnor U1493 (N_1493,N_1351,N_1385);
or U1494 (N_1494,N_1355,N_1411);
or U1495 (N_1495,N_1409,N_1422);
nand U1496 (N_1496,N_1365,N_1406);
and U1497 (N_1497,N_1356,N_1364);
or U1498 (N_1498,N_1406,N_1416);
and U1499 (N_1499,N_1368,N_1374);
nor U1500 (N_1500,N_1493,N_1471);
and U1501 (N_1501,N_1427,N_1459);
or U1502 (N_1502,N_1482,N_1452);
nand U1503 (N_1503,N_1429,N_1483);
and U1504 (N_1504,N_1438,N_1440);
or U1505 (N_1505,N_1428,N_1433);
nor U1506 (N_1506,N_1487,N_1473);
nand U1507 (N_1507,N_1463,N_1492);
xnor U1508 (N_1508,N_1462,N_1435);
and U1509 (N_1509,N_1481,N_1470);
and U1510 (N_1510,N_1437,N_1461);
or U1511 (N_1511,N_1496,N_1489);
and U1512 (N_1512,N_1449,N_1478);
or U1513 (N_1513,N_1479,N_1450);
xnor U1514 (N_1514,N_1446,N_1484);
nand U1515 (N_1515,N_1474,N_1457);
nand U1516 (N_1516,N_1466,N_1431);
and U1517 (N_1517,N_1455,N_1443);
xnor U1518 (N_1518,N_1434,N_1451);
and U1519 (N_1519,N_1468,N_1488);
nor U1520 (N_1520,N_1445,N_1495);
or U1521 (N_1521,N_1497,N_1486);
and U1522 (N_1522,N_1480,N_1441);
or U1523 (N_1523,N_1475,N_1436);
or U1524 (N_1524,N_1454,N_1485);
and U1525 (N_1525,N_1448,N_1456);
and U1526 (N_1526,N_1472,N_1460);
xnor U1527 (N_1527,N_1430,N_1442);
nand U1528 (N_1528,N_1469,N_1494);
and U1529 (N_1529,N_1476,N_1447);
and U1530 (N_1530,N_1491,N_1477);
xor U1531 (N_1531,N_1453,N_1467);
or U1532 (N_1532,N_1425,N_1432);
and U1533 (N_1533,N_1426,N_1444);
or U1534 (N_1534,N_1465,N_1439);
and U1535 (N_1535,N_1499,N_1464);
and U1536 (N_1536,N_1458,N_1498);
nand U1537 (N_1537,N_1490,N_1463);
nor U1538 (N_1538,N_1436,N_1484);
xor U1539 (N_1539,N_1472,N_1453);
and U1540 (N_1540,N_1459,N_1489);
xor U1541 (N_1541,N_1457,N_1492);
nor U1542 (N_1542,N_1426,N_1465);
or U1543 (N_1543,N_1467,N_1483);
or U1544 (N_1544,N_1490,N_1429);
or U1545 (N_1545,N_1475,N_1467);
or U1546 (N_1546,N_1488,N_1438);
or U1547 (N_1547,N_1434,N_1431);
and U1548 (N_1548,N_1483,N_1472);
nor U1549 (N_1549,N_1484,N_1475);
nor U1550 (N_1550,N_1427,N_1486);
and U1551 (N_1551,N_1470,N_1428);
nor U1552 (N_1552,N_1476,N_1466);
xor U1553 (N_1553,N_1465,N_1471);
nor U1554 (N_1554,N_1464,N_1460);
or U1555 (N_1555,N_1440,N_1499);
nor U1556 (N_1556,N_1478,N_1461);
and U1557 (N_1557,N_1472,N_1496);
nand U1558 (N_1558,N_1498,N_1475);
or U1559 (N_1559,N_1459,N_1482);
and U1560 (N_1560,N_1437,N_1471);
or U1561 (N_1561,N_1492,N_1440);
nand U1562 (N_1562,N_1476,N_1499);
nor U1563 (N_1563,N_1432,N_1479);
or U1564 (N_1564,N_1425,N_1427);
or U1565 (N_1565,N_1498,N_1461);
nor U1566 (N_1566,N_1437,N_1462);
xor U1567 (N_1567,N_1448,N_1446);
and U1568 (N_1568,N_1487,N_1452);
and U1569 (N_1569,N_1447,N_1479);
or U1570 (N_1570,N_1453,N_1496);
nand U1571 (N_1571,N_1453,N_1466);
and U1572 (N_1572,N_1495,N_1428);
nor U1573 (N_1573,N_1457,N_1438);
or U1574 (N_1574,N_1440,N_1489);
nand U1575 (N_1575,N_1501,N_1521);
xor U1576 (N_1576,N_1520,N_1509);
or U1577 (N_1577,N_1549,N_1544);
or U1578 (N_1578,N_1565,N_1557);
nand U1579 (N_1579,N_1507,N_1562);
nand U1580 (N_1580,N_1543,N_1536);
xnor U1581 (N_1581,N_1524,N_1529);
and U1582 (N_1582,N_1566,N_1510);
or U1583 (N_1583,N_1561,N_1518);
nand U1584 (N_1584,N_1563,N_1568);
xor U1585 (N_1585,N_1500,N_1515);
nand U1586 (N_1586,N_1570,N_1574);
nand U1587 (N_1587,N_1571,N_1526);
nor U1588 (N_1588,N_1523,N_1508);
nor U1589 (N_1589,N_1558,N_1531);
and U1590 (N_1590,N_1522,N_1546);
nor U1591 (N_1591,N_1547,N_1556);
xor U1592 (N_1592,N_1569,N_1511);
nand U1593 (N_1593,N_1506,N_1545);
or U1594 (N_1594,N_1539,N_1519);
xnor U1595 (N_1595,N_1527,N_1516);
or U1596 (N_1596,N_1567,N_1554);
or U1597 (N_1597,N_1559,N_1541);
xor U1598 (N_1598,N_1538,N_1530);
xor U1599 (N_1599,N_1514,N_1502);
nor U1600 (N_1600,N_1551,N_1503);
nor U1601 (N_1601,N_1548,N_1572);
nor U1602 (N_1602,N_1552,N_1505);
xor U1603 (N_1603,N_1525,N_1550);
and U1604 (N_1604,N_1535,N_1533);
or U1605 (N_1605,N_1537,N_1553);
nor U1606 (N_1606,N_1504,N_1528);
and U1607 (N_1607,N_1542,N_1517);
and U1608 (N_1608,N_1512,N_1513);
nor U1609 (N_1609,N_1573,N_1560);
nor U1610 (N_1610,N_1564,N_1534);
and U1611 (N_1611,N_1540,N_1555);
xor U1612 (N_1612,N_1532,N_1555);
or U1613 (N_1613,N_1540,N_1502);
nand U1614 (N_1614,N_1536,N_1568);
or U1615 (N_1615,N_1507,N_1560);
and U1616 (N_1616,N_1530,N_1568);
nor U1617 (N_1617,N_1549,N_1518);
nand U1618 (N_1618,N_1517,N_1521);
or U1619 (N_1619,N_1561,N_1513);
and U1620 (N_1620,N_1501,N_1551);
nand U1621 (N_1621,N_1563,N_1532);
xor U1622 (N_1622,N_1513,N_1521);
nand U1623 (N_1623,N_1569,N_1562);
nor U1624 (N_1624,N_1565,N_1539);
nand U1625 (N_1625,N_1517,N_1536);
nor U1626 (N_1626,N_1536,N_1501);
or U1627 (N_1627,N_1502,N_1503);
nand U1628 (N_1628,N_1523,N_1549);
or U1629 (N_1629,N_1548,N_1512);
nor U1630 (N_1630,N_1570,N_1549);
xor U1631 (N_1631,N_1562,N_1508);
nand U1632 (N_1632,N_1549,N_1521);
nor U1633 (N_1633,N_1545,N_1528);
and U1634 (N_1634,N_1516,N_1561);
nor U1635 (N_1635,N_1512,N_1570);
nor U1636 (N_1636,N_1565,N_1511);
and U1637 (N_1637,N_1565,N_1571);
or U1638 (N_1638,N_1537,N_1541);
xor U1639 (N_1639,N_1510,N_1574);
or U1640 (N_1640,N_1550,N_1508);
or U1641 (N_1641,N_1527,N_1526);
nor U1642 (N_1642,N_1573,N_1565);
nand U1643 (N_1643,N_1514,N_1545);
nand U1644 (N_1644,N_1526,N_1510);
or U1645 (N_1645,N_1530,N_1535);
nor U1646 (N_1646,N_1564,N_1510);
nor U1647 (N_1647,N_1512,N_1502);
nand U1648 (N_1648,N_1534,N_1523);
or U1649 (N_1649,N_1525,N_1563);
and U1650 (N_1650,N_1640,N_1637);
nand U1651 (N_1651,N_1626,N_1593);
xnor U1652 (N_1652,N_1596,N_1608);
or U1653 (N_1653,N_1580,N_1620);
nor U1654 (N_1654,N_1594,N_1597);
nor U1655 (N_1655,N_1634,N_1604);
nand U1656 (N_1656,N_1612,N_1601);
and U1657 (N_1657,N_1636,N_1592);
or U1658 (N_1658,N_1611,N_1606);
or U1659 (N_1659,N_1586,N_1635);
nand U1660 (N_1660,N_1613,N_1577);
or U1661 (N_1661,N_1631,N_1642);
and U1662 (N_1662,N_1587,N_1582);
nand U1663 (N_1663,N_1603,N_1645);
or U1664 (N_1664,N_1625,N_1600);
nand U1665 (N_1665,N_1616,N_1581);
or U1666 (N_1666,N_1633,N_1607);
nand U1667 (N_1667,N_1641,N_1609);
nor U1668 (N_1668,N_1638,N_1644);
nor U1669 (N_1669,N_1618,N_1632);
xnor U1670 (N_1670,N_1588,N_1627);
or U1671 (N_1671,N_1615,N_1591);
nor U1672 (N_1672,N_1648,N_1647);
xor U1673 (N_1673,N_1578,N_1576);
and U1674 (N_1674,N_1602,N_1583);
or U1675 (N_1675,N_1621,N_1623);
xor U1676 (N_1676,N_1575,N_1639);
nand U1677 (N_1677,N_1584,N_1649);
nand U1678 (N_1678,N_1622,N_1585);
and U1679 (N_1679,N_1579,N_1630);
nand U1680 (N_1680,N_1614,N_1617);
nor U1681 (N_1681,N_1599,N_1619);
nor U1682 (N_1682,N_1598,N_1646);
and U1683 (N_1683,N_1628,N_1610);
nand U1684 (N_1684,N_1590,N_1589);
and U1685 (N_1685,N_1605,N_1595);
nor U1686 (N_1686,N_1643,N_1624);
nand U1687 (N_1687,N_1629,N_1589);
nor U1688 (N_1688,N_1644,N_1597);
nor U1689 (N_1689,N_1649,N_1629);
nand U1690 (N_1690,N_1616,N_1608);
xor U1691 (N_1691,N_1632,N_1597);
nor U1692 (N_1692,N_1649,N_1643);
nor U1693 (N_1693,N_1625,N_1582);
and U1694 (N_1694,N_1605,N_1646);
nor U1695 (N_1695,N_1588,N_1617);
xor U1696 (N_1696,N_1626,N_1612);
nand U1697 (N_1697,N_1643,N_1642);
or U1698 (N_1698,N_1581,N_1623);
xnor U1699 (N_1699,N_1620,N_1590);
nor U1700 (N_1700,N_1580,N_1612);
and U1701 (N_1701,N_1601,N_1610);
xor U1702 (N_1702,N_1575,N_1605);
and U1703 (N_1703,N_1600,N_1590);
and U1704 (N_1704,N_1579,N_1622);
nand U1705 (N_1705,N_1600,N_1597);
xnor U1706 (N_1706,N_1622,N_1646);
nand U1707 (N_1707,N_1641,N_1634);
or U1708 (N_1708,N_1581,N_1643);
xnor U1709 (N_1709,N_1640,N_1578);
or U1710 (N_1710,N_1639,N_1610);
or U1711 (N_1711,N_1622,N_1613);
xor U1712 (N_1712,N_1622,N_1641);
and U1713 (N_1713,N_1587,N_1633);
or U1714 (N_1714,N_1583,N_1643);
and U1715 (N_1715,N_1623,N_1578);
and U1716 (N_1716,N_1612,N_1632);
nor U1717 (N_1717,N_1597,N_1609);
nor U1718 (N_1718,N_1642,N_1592);
nand U1719 (N_1719,N_1626,N_1603);
and U1720 (N_1720,N_1589,N_1641);
nand U1721 (N_1721,N_1597,N_1584);
and U1722 (N_1722,N_1588,N_1600);
nand U1723 (N_1723,N_1618,N_1604);
nor U1724 (N_1724,N_1642,N_1638);
nand U1725 (N_1725,N_1670,N_1690);
and U1726 (N_1726,N_1662,N_1695);
and U1727 (N_1727,N_1664,N_1671);
or U1728 (N_1728,N_1715,N_1710);
nand U1729 (N_1729,N_1697,N_1707);
and U1730 (N_1730,N_1678,N_1653);
and U1731 (N_1731,N_1655,N_1651);
xor U1732 (N_1732,N_1711,N_1666);
nor U1733 (N_1733,N_1657,N_1689);
nand U1734 (N_1734,N_1658,N_1700);
nor U1735 (N_1735,N_1681,N_1713);
xor U1736 (N_1736,N_1694,N_1701);
and U1737 (N_1737,N_1696,N_1685);
and U1738 (N_1738,N_1676,N_1667);
nand U1739 (N_1739,N_1688,N_1687);
nand U1740 (N_1740,N_1650,N_1677);
nand U1741 (N_1741,N_1714,N_1721);
and U1742 (N_1742,N_1716,N_1712);
nor U1743 (N_1743,N_1675,N_1706);
or U1744 (N_1744,N_1661,N_1724);
or U1745 (N_1745,N_1720,N_1704);
nand U1746 (N_1746,N_1709,N_1663);
nand U1747 (N_1747,N_1684,N_1722);
or U1748 (N_1748,N_1702,N_1673);
and U1749 (N_1749,N_1674,N_1679);
or U1750 (N_1750,N_1669,N_1660);
or U1751 (N_1751,N_1686,N_1665);
nor U1752 (N_1752,N_1693,N_1708);
or U1753 (N_1753,N_1699,N_1659);
nor U1754 (N_1754,N_1672,N_1723);
or U1755 (N_1755,N_1654,N_1692);
nand U1756 (N_1756,N_1683,N_1705);
or U1757 (N_1757,N_1680,N_1691);
and U1758 (N_1758,N_1719,N_1652);
xor U1759 (N_1759,N_1668,N_1703);
or U1760 (N_1760,N_1717,N_1656);
nor U1761 (N_1761,N_1698,N_1682);
nand U1762 (N_1762,N_1718,N_1664);
nand U1763 (N_1763,N_1686,N_1698);
and U1764 (N_1764,N_1702,N_1676);
nand U1765 (N_1765,N_1719,N_1703);
or U1766 (N_1766,N_1703,N_1699);
nor U1767 (N_1767,N_1682,N_1724);
nor U1768 (N_1768,N_1699,N_1711);
or U1769 (N_1769,N_1701,N_1676);
nand U1770 (N_1770,N_1674,N_1663);
nor U1771 (N_1771,N_1697,N_1680);
nor U1772 (N_1772,N_1714,N_1655);
or U1773 (N_1773,N_1687,N_1695);
nor U1774 (N_1774,N_1724,N_1708);
nor U1775 (N_1775,N_1709,N_1687);
nor U1776 (N_1776,N_1663,N_1652);
and U1777 (N_1777,N_1708,N_1663);
xor U1778 (N_1778,N_1678,N_1677);
nor U1779 (N_1779,N_1651,N_1672);
and U1780 (N_1780,N_1714,N_1715);
nor U1781 (N_1781,N_1675,N_1691);
nor U1782 (N_1782,N_1657,N_1679);
or U1783 (N_1783,N_1705,N_1670);
and U1784 (N_1784,N_1717,N_1666);
or U1785 (N_1785,N_1687,N_1683);
nor U1786 (N_1786,N_1661,N_1664);
nor U1787 (N_1787,N_1724,N_1655);
nor U1788 (N_1788,N_1709,N_1676);
nor U1789 (N_1789,N_1715,N_1676);
and U1790 (N_1790,N_1668,N_1716);
nor U1791 (N_1791,N_1707,N_1696);
or U1792 (N_1792,N_1720,N_1724);
xnor U1793 (N_1793,N_1663,N_1661);
or U1794 (N_1794,N_1674,N_1669);
nand U1795 (N_1795,N_1708,N_1692);
and U1796 (N_1796,N_1697,N_1696);
or U1797 (N_1797,N_1659,N_1720);
nand U1798 (N_1798,N_1671,N_1650);
nand U1799 (N_1799,N_1712,N_1696);
or U1800 (N_1800,N_1735,N_1767);
nor U1801 (N_1801,N_1742,N_1756);
or U1802 (N_1802,N_1776,N_1773);
or U1803 (N_1803,N_1746,N_1741);
or U1804 (N_1804,N_1760,N_1762);
nand U1805 (N_1805,N_1770,N_1761);
and U1806 (N_1806,N_1734,N_1736);
or U1807 (N_1807,N_1768,N_1743);
nand U1808 (N_1808,N_1787,N_1780);
or U1809 (N_1809,N_1752,N_1775);
nor U1810 (N_1810,N_1790,N_1759);
and U1811 (N_1811,N_1788,N_1797);
xor U1812 (N_1812,N_1784,N_1748);
or U1813 (N_1813,N_1749,N_1757);
or U1814 (N_1814,N_1731,N_1755);
xnor U1815 (N_1815,N_1739,N_1733);
nor U1816 (N_1816,N_1778,N_1737);
and U1817 (N_1817,N_1763,N_1727);
and U1818 (N_1818,N_1754,N_1728);
or U1819 (N_1819,N_1769,N_1766);
nor U1820 (N_1820,N_1774,N_1747);
and U1821 (N_1821,N_1750,N_1771);
or U1822 (N_1822,N_1782,N_1795);
or U1823 (N_1823,N_1725,N_1793);
xnor U1824 (N_1824,N_1758,N_1729);
nor U1825 (N_1825,N_1772,N_1726);
nand U1826 (N_1826,N_1730,N_1796);
nand U1827 (N_1827,N_1738,N_1779);
and U1828 (N_1828,N_1781,N_1792);
nor U1829 (N_1829,N_1764,N_1732);
and U1830 (N_1830,N_1744,N_1753);
nor U1831 (N_1831,N_1765,N_1789);
nor U1832 (N_1832,N_1791,N_1798);
or U1833 (N_1833,N_1777,N_1785);
and U1834 (N_1834,N_1786,N_1783);
or U1835 (N_1835,N_1794,N_1751);
or U1836 (N_1836,N_1745,N_1799);
or U1837 (N_1837,N_1740,N_1797);
or U1838 (N_1838,N_1759,N_1732);
and U1839 (N_1839,N_1789,N_1775);
xor U1840 (N_1840,N_1769,N_1760);
nor U1841 (N_1841,N_1799,N_1791);
or U1842 (N_1842,N_1778,N_1732);
or U1843 (N_1843,N_1725,N_1731);
or U1844 (N_1844,N_1728,N_1789);
nand U1845 (N_1845,N_1778,N_1750);
and U1846 (N_1846,N_1795,N_1783);
or U1847 (N_1847,N_1769,N_1740);
and U1848 (N_1848,N_1764,N_1734);
xnor U1849 (N_1849,N_1756,N_1764);
and U1850 (N_1850,N_1749,N_1794);
and U1851 (N_1851,N_1746,N_1758);
nor U1852 (N_1852,N_1797,N_1726);
xor U1853 (N_1853,N_1787,N_1766);
nor U1854 (N_1854,N_1739,N_1775);
nand U1855 (N_1855,N_1729,N_1784);
and U1856 (N_1856,N_1737,N_1734);
xnor U1857 (N_1857,N_1774,N_1767);
nand U1858 (N_1858,N_1775,N_1796);
xnor U1859 (N_1859,N_1781,N_1766);
nand U1860 (N_1860,N_1727,N_1758);
xor U1861 (N_1861,N_1764,N_1742);
and U1862 (N_1862,N_1778,N_1781);
and U1863 (N_1863,N_1762,N_1739);
nor U1864 (N_1864,N_1742,N_1788);
and U1865 (N_1865,N_1728,N_1793);
nor U1866 (N_1866,N_1799,N_1760);
and U1867 (N_1867,N_1792,N_1727);
or U1868 (N_1868,N_1765,N_1752);
or U1869 (N_1869,N_1761,N_1799);
nand U1870 (N_1870,N_1752,N_1741);
and U1871 (N_1871,N_1763,N_1789);
or U1872 (N_1872,N_1793,N_1789);
xor U1873 (N_1873,N_1774,N_1789);
nand U1874 (N_1874,N_1754,N_1736);
or U1875 (N_1875,N_1802,N_1839);
xnor U1876 (N_1876,N_1860,N_1824);
or U1877 (N_1877,N_1805,N_1800);
nand U1878 (N_1878,N_1812,N_1807);
nor U1879 (N_1879,N_1810,N_1870);
and U1880 (N_1880,N_1822,N_1834);
nor U1881 (N_1881,N_1825,N_1849);
and U1882 (N_1882,N_1867,N_1850);
or U1883 (N_1883,N_1819,N_1816);
xnor U1884 (N_1884,N_1855,N_1848);
and U1885 (N_1885,N_1846,N_1871);
nand U1886 (N_1886,N_1869,N_1840);
and U1887 (N_1887,N_1803,N_1821);
and U1888 (N_1888,N_1873,N_1808);
nand U1889 (N_1889,N_1854,N_1806);
nor U1890 (N_1890,N_1866,N_1843);
and U1891 (N_1891,N_1827,N_1868);
and U1892 (N_1892,N_1833,N_1823);
xnor U1893 (N_1893,N_1829,N_1864);
nor U1894 (N_1894,N_1857,N_1856);
nor U1895 (N_1895,N_1814,N_1841);
and U1896 (N_1896,N_1861,N_1862);
or U1897 (N_1897,N_1847,N_1842);
nor U1898 (N_1898,N_1835,N_1836);
and U1899 (N_1899,N_1826,N_1811);
or U1900 (N_1900,N_1817,N_1837);
nor U1901 (N_1901,N_1844,N_1865);
nor U1902 (N_1902,N_1831,N_1845);
and U1903 (N_1903,N_1872,N_1874);
nand U1904 (N_1904,N_1853,N_1830);
nor U1905 (N_1905,N_1838,N_1863);
xor U1906 (N_1906,N_1820,N_1809);
nand U1907 (N_1907,N_1852,N_1828);
nand U1908 (N_1908,N_1851,N_1813);
xnor U1909 (N_1909,N_1859,N_1818);
nand U1910 (N_1910,N_1804,N_1801);
nand U1911 (N_1911,N_1815,N_1858);
nor U1912 (N_1912,N_1832,N_1862);
nand U1913 (N_1913,N_1871,N_1823);
nand U1914 (N_1914,N_1871,N_1847);
xor U1915 (N_1915,N_1857,N_1868);
and U1916 (N_1916,N_1817,N_1828);
nand U1917 (N_1917,N_1835,N_1811);
nand U1918 (N_1918,N_1814,N_1874);
xor U1919 (N_1919,N_1865,N_1815);
or U1920 (N_1920,N_1851,N_1836);
nor U1921 (N_1921,N_1808,N_1815);
and U1922 (N_1922,N_1857,N_1853);
xnor U1923 (N_1923,N_1832,N_1831);
or U1924 (N_1924,N_1824,N_1812);
or U1925 (N_1925,N_1855,N_1860);
and U1926 (N_1926,N_1804,N_1813);
nor U1927 (N_1927,N_1843,N_1855);
nor U1928 (N_1928,N_1840,N_1827);
xnor U1929 (N_1929,N_1828,N_1849);
and U1930 (N_1930,N_1817,N_1830);
or U1931 (N_1931,N_1816,N_1811);
xnor U1932 (N_1932,N_1845,N_1862);
nor U1933 (N_1933,N_1860,N_1813);
nor U1934 (N_1934,N_1833,N_1824);
nand U1935 (N_1935,N_1840,N_1846);
nor U1936 (N_1936,N_1818,N_1812);
or U1937 (N_1937,N_1864,N_1823);
xnor U1938 (N_1938,N_1836,N_1853);
nand U1939 (N_1939,N_1852,N_1836);
and U1940 (N_1940,N_1832,N_1852);
and U1941 (N_1941,N_1870,N_1849);
and U1942 (N_1942,N_1801,N_1871);
and U1943 (N_1943,N_1800,N_1818);
nor U1944 (N_1944,N_1803,N_1868);
nand U1945 (N_1945,N_1864,N_1858);
nand U1946 (N_1946,N_1846,N_1850);
and U1947 (N_1947,N_1836,N_1825);
and U1948 (N_1948,N_1850,N_1842);
nand U1949 (N_1949,N_1819,N_1874);
nor U1950 (N_1950,N_1932,N_1901);
nand U1951 (N_1951,N_1937,N_1940);
nand U1952 (N_1952,N_1887,N_1918);
nor U1953 (N_1953,N_1923,N_1922);
and U1954 (N_1954,N_1896,N_1920);
nand U1955 (N_1955,N_1909,N_1915);
nand U1956 (N_1956,N_1942,N_1897);
nor U1957 (N_1957,N_1924,N_1905);
nor U1958 (N_1958,N_1895,N_1889);
or U1959 (N_1959,N_1927,N_1944);
xnor U1960 (N_1960,N_1919,N_1883);
and U1961 (N_1961,N_1912,N_1888);
nand U1962 (N_1962,N_1884,N_1931);
nand U1963 (N_1963,N_1893,N_1904);
nand U1964 (N_1964,N_1921,N_1941);
nand U1965 (N_1965,N_1890,N_1900);
and U1966 (N_1966,N_1934,N_1881);
nand U1967 (N_1967,N_1926,N_1947);
nor U1968 (N_1968,N_1878,N_1929);
nor U1969 (N_1969,N_1891,N_1880);
nor U1970 (N_1970,N_1908,N_1903);
xnor U1971 (N_1971,N_1928,N_1949);
nand U1972 (N_1972,N_1948,N_1875);
nand U1973 (N_1973,N_1898,N_1894);
and U1974 (N_1974,N_1930,N_1945);
nand U1975 (N_1975,N_1911,N_1877);
nor U1976 (N_1976,N_1916,N_1914);
or U1977 (N_1977,N_1892,N_1876);
or U1978 (N_1978,N_1899,N_1936);
nand U1979 (N_1979,N_1943,N_1907);
nor U1980 (N_1980,N_1885,N_1913);
nand U1981 (N_1981,N_1925,N_1935);
nand U1982 (N_1982,N_1946,N_1906);
xor U1983 (N_1983,N_1917,N_1882);
or U1984 (N_1984,N_1939,N_1910);
and U1985 (N_1985,N_1933,N_1879);
or U1986 (N_1986,N_1938,N_1886);
and U1987 (N_1987,N_1902,N_1941);
nand U1988 (N_1988,N_1883,N_1945);
nand U1989 (N_1989,N_1922,N_1926);
nand U1990 (N_1990,N_1898,N_1879);
or U1991 (N_1991,N_1906,N_1912);
and U1992 (N_1992,N_1908,N_1877);
nand U1993 (N_1993,N_1934,N_1875);
and U1994 (N_1994,N_1910,N_1898);
or U1995 (N_1995,N_1930,N_1889);
or U1996 (N_1996,N_1889,N_1942);
nor U1997 (N_1997,N_1919,N_1924);
nand U1998 (N_1998,N_1889,N_1917);
nor U1999 (N_1999,N_1948,N_1907);
or U2000 (N_2000,N_1882,N_1915);
nor U2001 (N_2001,N_1924,N_1881);
nor U2002 (N_2002,N_1902,N_1932);
or U2003 (N_2003,N_1911,N_1943);
nand U2004 (N_2004,N_1884,N_1899);
or U2005 (N_2005,N_1904,N_1898);
nand U2006 (N_2006,N_1949,N_1901);
nand U2007 (N_2007,N_1896,N_1924);
or U2008 (N_2008,N_1914,N_1896);
nand U2009 (N_2009,N_1912,N_1924);
nand U2010 (N_2010,N_1876,N_1887);
nand U2011 (N_2011,N_1911,N_1919);
nand U2012 (N_2012,N_1902,N_1911);
and U2013 (N_2013,N_1890,N_1943);
nor U2014 (N_2014,N_1900,N_1917);
xnor U2015 (N_2015,N_1883,N_1947);
nor U2016 (N_2016,N_1935,N_1890);
and U2017 (N_2017,N_1920,N_1912);
and U2018 (N_2018,N_1949,N_1936);
xor U2019 (N_2019,N_1927,N_1926);
and U2020 (N_2020,N_1875,N_1879);
nor U2021 (N_2021,N_1893,N_1943);
nand U2022 (N_2022,N_1936,N_1890);
nor U2023 (N_2023,N_1892,N_1925);
xnor U2024 (N_2024,N_1928,N_1903);
or U2025 (N_2025,N_2008,N_1992);
or U2026 (N_2026,N_2009,N_1973);
and U2027 (N_2027,N_1966,N_1994);
nand U2028 (N_2028,N_1963,N_1997);
and U2029 (N_2029,N_2020,N_2022);
and U2030 (N_2030,N_1978,N_2004);
and U2031 (N_2031,N_2001,N_1996);
nand U2032 (N_2032,N_1988,N_2024);
xor U2033 (N_2033,N_1958,N_2011);
xnor U2034 (N_2034,N_2010,N_2000);
nand U2035 (N_2035,N_1964,N_1979);
xnor U2036 (N_2036,N_2012,N_1961);
nor U2037 (N_2037,N_1984,N_1977);
and U2038 (N_2038,N_2006,N_1981);
xor U2039 (N_2039,N_1993,N_1980);
nand U2040 (N_2040,N_1967,N_1955);
nor U2041 (N_2041,N_2007,N_1991);
nor U2042 (N_2042,N_1962,N_2003);
nor U2043 (N_2043,N_1972,N_2005);
nor U2044 (N_2044,N_2018,N_2017);
and U2045 (N_2045,N_1975,N_1987);
nand U2046 (N_2046,N_2016,N_1990);
and U2047 (N_2047,N_1956,N_1952);
nand U2048 (N_2048,N_2015,N_1969);
or U2049 (N_2049,N_2013,N_2019);
and U2050 (N_2050,N_2014,N_1971);
nor U2051 (N_2051,N_1995,N_1974);
nor U2052 (N_2052,N_1998,N_1985);
xnor U2053 (N_2053,N_1960,N_1989);
and U2054 (N_2054,N_2002,N_1976);
nand U2055 (N_2055,N_1959,N_1954);
nand U2056 (N_2056,N_2021,N_1986);
and U2057 (N_2057,N_1953,N_1951);
nand U2058 (N_2058,N_1982,N_1950);
nor U2059 (N_2059,N_1968,N_2023);
nor U2060 (N_2060,N_1965,N_1999);
and U2061 (N_2061,N_1983,N_1970);
nand U2062 (N_2062,N_1957,N_1999);
or U2063 (N_2063,N_1950,N_1990);
nand U2064 (N_2064,N_1984,N_2007);
nor U2065 (N_2065,N_2006,N_1991);
or U2066 (N_2066,N_2008,N_1974);
xnor U2067 (N_2067,N_2001,N_1953);
and U2068 (N_2068,N_1982,N_1966);
xor U2069 (N_2069,N_1970,N_1959);
and U2070 (N_2070,N_1977,N_1959);
and U2071 (N_2071,N_2002,N_2015);
nand U2072 (N_2072,N_2000,N_2008);
nor U2073 (N_2073,N_2006,N_1988);
and U2074 (N_2074,N_1999,N_2004);
nand U2075 (N_2075,N_1970,N_1971);
or U2076 (N_2076,N_1989,N_1950);
or U2077 (N_2077,N_1991,N_2008);
or U2078 (N_2078,N_2012,N_2017);
or U2079 (N_2079,N_1988,N_2022);
nand U2080 (N_2080,N_1961,N_1993);
or U2081 (N_2081,N_2017,N_1965);
and U2082 (N_2082,N_1980,N_2019);
nand U2083 (N_2083,N_1986,N_2008);
and U2084 (N_2084,N_2018,N_2014);
xor U2085 (N_2085,N_1962,N_1980);
and U2086 (N_2086,N_1981,N_1976);
and U2087 (N_2087,N_1972,N_2012);
and U2088 (N_2088,N_1991,N_1956);
xnor U2089 (N_2089,N_1967,N_1954);
nor U2090 (N_2090,N_1970,N_1963);
nor U2091 (N_2091,N_2000,N_2004);
nor U2092 (N_2092,N_1978,N_1951);
nor U2093 (N_2093,N_2002,N_1989);
nor U2094 (N_2094,N_1961,N_1952);
xor U2095 (N_2095,N_2005,N_2007);
and U2096 (N_2096,N_1963,N_1990);
nor U2097 (N_2097,N_1968,N_1999);
nand U2098 (N_2098,N_2010,N_2012);
or U2099 (N_2099,N_1964,N_2011);
nand U2100 (N_2100,N_2095,N_2067);
or U2101 (N_2101,N_2071,N_2065);
xor U2102 (N_2102,N_2057,N_2077);
nand U2103 (N_2103,N_2028,N_2027);
xnor U2104 (N_2104,N_2050,N_2073);
or U2105 (N_2105,N_2060,N_2074);
xnor U2106 (N_2106,N_2096,N_2058);
nor U2107 (N_2107,N_2091,N_2035);
or U2108 (N_2108,N_2033,N_2092);
nand U2109 (N_2109,N_2036,N_2061);
and U2110 (N_2110,N_2048,N_2079);
and U2111 (N_2111,N_2039,N_2083);
nand U2112 (N_2112,N_2047,N_2089);
nor U2113 (N_2113,N_2086,N_2051);
nand U2114 (N_2114,N_2099,N_2030);
nand U2115 (N_2115,N_2044,N_2062);
and U2116 (N_2116,N_2059,N_2064);
or U2117 (N_2117,N_2093,N_2055);
nor U2118 (N_2118,N_2040,N_2070);
nand U2119 (N_2119,N_2066,N_2043);
or U2120 (N_2120,N_2097,N_2053);
or U2121 (N_2121,N_2085,N_2041);
and U2122 (N_2122,N_2075,N_2063);
nand U2123 (N_2123,N_2034,N_2090);
or U2124 (N_2124,N_2081,N_2037);
nand U2125 (N_2125,N_2072,N_2082);
or U2126 (N_2126,N_2084,N_2046);
and U2127 (N_2127,N_2087,N_2078);
and U2128 (N_2128,N_2076,N_2025);
and U2129 (N_2129,N_2098,N_2031);
and U2130 (N_2130,N_2032,N_2088);
or U2131 (N_2131,N_2026,N_2049);
xor U2132 (N_2132,N_2069,N_2068);
or U2133 (N_2133,N_2045,N_2029);
and U2134 (N_2134,N_2054,N_2094);
nand U2135 (N_2135,N_2052,N_2080);
or U2136 (N_2136,N_2042,N_2056);
nor U2137 (N_2137,N_2038,N_2095);
xnor U2138 (N_2138,N_2052,N_2090);
nor U2139 (N_2139,N_2041,N_2031);
nand U2140 (N_2140,N_2098,N_2049);
xnor U2141 (N_2141,N_2027,N_2073);
or U2142 (N_2142,N_2072,N_2074);
nand U2143 (N_2143,N_2078,N_2061);
and U2144 (N_2144,N_2059,N_2049);
nand U2145 (N_2145,N_2088,N_2073);
nor U2146 (N_2146,N_2099,N_2041);
nor U2147 (N_2147,N_2058,N_2069);
nor U2148 (N_2148,N_2053,N_2050);
xnor U2149 (N_2149,N_2069,N_2049);
xnor U2150 (N_2150,N_2025,N_2069);
or U2151 (N_2151,N_2075,N_2098);
xnor U2152 (N_2152,N_2088,N_2033);
and U2153 (N_2153,N_2061,N_2046);
and U2154 (N_2154,N_2093,N_2039);
nor U2155 (N_2155,N_2082,N_2052);
nor U2156 (N_2156,N_2038,N_2076);
and U2157 (N_2157,N_2053,N_2081);
nor U2158 (N_2158,N_2051,N_2062);
or U2159 (N_2159,N_2070,N_2099);
nand U2160 (N_2160,N_2041,N_2052);
and U2161 (N_2161,N_2046,N_2085);
and U2162 (N_2162,N_2033,N_2075);
nand U2163 (N_2163,N_2043,N_2070);
or U2164 (N_2164,N_2094,N_2070);
nor U2165 (N_2165,N_2040,N_2031);
or U2166 (N_2166,N_2045,N_2076);
nor U2167 (N_2167,N_2057,N_2062);
and U2168 (N_2168,N_2055,N_2051);
nand U2169 (N_2169,N_2027,N_2090);
or U2170 (N_2170,N_2025,N_2078);
and U2171 (N_2171,N_2063,N_2039);
nand U2172 (N_2172,N_2080,N_2056);
or U2173 (N_2173,N_2046,N_2079);
and U2174 (N_2174,N_2077,N_2098);
or U2175 (N_2175,N_2154,N_2123);
and U2176 (N_2176,N_2130,N_2120);
and U2177 (N_2177,N_2116,N_2144);
and U2178 (N_2178,N_2111,N_2112);
nand U2179 (N_2179,N_2158,N_2102);
and U2180 (N_2180,N_2150,N_2142);
and U2181 (N_2181,N_2159,N_2100);
or U2182 (N_2182,N_2170,N_2151);
xnor U2183 (N_2183,N_2129,N_2107);
or U2184 (N_2184,N_2161,N_2140);
nand U2185 (N_2185,N_2138,N_2171);
or U2186 (N_2186,N_2119,N_2134);
or U2187 (N_2187,N_2131,N_2101);
and U2188 (N_2188,N_2174,N_2121);
and U2189 (N_2189,N_2136,N_2149);
nor U2190 (N_2190,N_2156,N_2108);
or U2191 (N_2191,N_2145,N_2169);
nand U2192 (N_2192,N_2143,N_2133);
xnor U2193 (N_2193,N_2173,N_2152);
or U2194 (N_2194,N_2115,N_2103);
and U2195 (N_2195,N_2126,N_2164);
or U2196 (N_2196,N_2147,N_2157);
xor U2197 (N_2197,N_2118,N_2139);
or U2198 (N_2198,N_2167,N_2114);
nor U2199 (N_2199,N_2146,N_2109);
or U2200 (N_2200,N_2128,N_2160);
and U2201 (N_2201,N_2104,N_2122);
nor U2202 (N_2202,N_2106,N_2168);
nand U2203 (N_2203,N_2148,N_2117);
nor U2204 (N_2204,N_2105,N_2162);
xnor U2205 (N_2205,N_2165,N_2141);
or U2206 (N_2206,N_2127,N_2166);
or U2207 (N_2207,N_2135,N_2132);
or U2208 (N_2208,N_2163,N_2153);
or U2209 (N_2209,N_2110,N_2113);
xor U2210 (N_2210,N_2172,N_2155);
or U2211 (N_2211,N_2137,N_2124);
nand U2212 (N_2212,N_2125,N_2149);
and U2213 (N_2213,N_2107,N_2119);
nor U2214 (N_2214,N_2127,N_2159);
or U2215 (N_2215,N_2108,N_2158);
nor U2216 (N_2216,N_2102,N_2110);
xnor U2217 (N_2217,N_2106,N_2111);
nand U2218 (N_2218,N_2141,N_2136);
and U2219 (N_2219,N_2141,N_2169);
xnor U2220 (N_2220,N_2149,N_2142);
nand U2221 (N_2221,N_2138,N_2109);
and U2222 (N_2222,N_2105,N_2169);
or U2223 (N_2223,N_2169,N_2149);
and U2224 (N_2224,N_2139,N_2130);
and U2225 (N_2225,N_2118,N_2104);
and U2226 (N_2226,N_2107,N_2109);
or U2227 (N_2227,N_2119,N_2169);
nand U2228 (N_2228,N_2167,N_2131);
nand U2229 (N_2229,N_2101,N_2158);
xor U2230 (N_2230,N_2174,N_2146);
nand U2231 (N_2231,N_2126,N_2148);
or U2232 (N_2232,N_2107,N_2169);
nor U2233 (N_2233,N_2106,N_2164);
or U2234 (N_2234,N_2140,N_2101);
and U2235 (N_2235,N_2145,N_2116);
nor U2236 (N_2236,N_2140,N_2174);
nor U2237 (N_2237,N_2153,N_2165);
and U2238 (N_2238,N_2167,N_2152);
nor U2239 (N_2239,N_2111,N_2164);
nor U2240 (N_2240,N_2127,N_2158);
or U2241 (N_2241,N_2127,N_2147);
nand U2242 (N_2242,N_2151,N_2120);
and U2243 (N_2243,N_2109,N_2145);
and U2244 (N_2244,N_2158,N_2149);
nor U2245 (N_2245,N_2125,N_2123);
or U2246 (N_2246,N_2120,N_2138);
xor U2247 (N_2247,N_2123,N_2153);
or U2248 (N_2248,N_2151,N_2147);
and U2249 (N_2249,N_2167,N_2111);
or U2250 (N_2250,N_2193,N_2232);
xor U2251 (N_2251,N_2245,N_2184);
nor U2252 (N_2252,N_2205,N_2237);
nor U2253 (N_2253,N_2224,N_2200);
nor U2254 (N_2254,N_2204,N_2185);
nand U2255 (N_2255,N_2201,N_2214);
nand U2256 (N_2256,N_2246,N_2229);
nor U2257 (N_2257,N_2211,N_2220);
xnor U2258 (N_2258,N_2221,N_2238);
and U2259 (N_2259,N_2217,N_2225);
or U2260 (N_2260,N_2207,N_2191);
and U2261 (N_2261,N_2180,N_2175);
or U2262 (N_2262,N_2186,N_2216);
nand U2263 (N_2263,N_2243,N_2209);
or U2264 (N_2264,N_2240,N_2223);
and U2265 (N_2265,N_2239,N_2195);
xnor U2266 (N_2266,N_2228,N_2192);
nand U2267 (N_2267,N_2234,N_2182);
nor U2268 (N_2268,N_2188,N_2215);
nor U2269 (N_2269,N_2249,N_2181);
or U2270 (N_2270,N_2235,N_2248);
nor U2271 (N_2271,N_2222,N_2183);
or U2272 (N_2272,N_2212,N_2202);
and U2273 (N_2273,N_2208,N_2194);
and U2274 (N_2274,N_2227,N_2210);
nor U2275 (N_2275,N_2179,N_2231);
nand U2276 (N_2276,N_2233,N_2230);
xor U2277 (N_2277,N_2241,N_2197);
nand U2278 (N_2278,N_2236,N_2226);
nand U2279 (N_2279,N_2199,N_2203);
and U2280 (N_2280,N_2219,N_2213);
and U2281 (N_2281,N_2206,N_2189);
or U2282 (N_2282,N_2177,N_2198);
and U2283 (N_2283,N_2218,N_2187);
and U2284 (N_2284,N_2244,N_2242);
and U2285 (N_2285,N_2190,N_2176);
nand U2286 (N_2286,N_2178,N_2196);
xnor U2287 (N_2287,N_2247,N_2205);
nand U2288 (N_2288,N_2190,N_2214);
and U2289 (N_2289,N_2221,N_2180);
nand U2290 (N_2290,N_2212,N_2213);
xnor U2291 (N_2291,N_2188,N_2242);
or U2292 (N_2292,N_2239,N_2198);
and U2293 (N_2293,N_2186,N_2241);
and U2294 (N_2294,N_2178,N_2175);
or U2295 (N_2295,N_2178,N_2192);
nand U2296 (N_2296,N_2183,N_2182);
nor U2297 (N_2297,N_2237,N_2202);
nor U2298 (N_2298,N_2180,N_2208);
nand U2299 (N_2299,N_2195,N_2191);
nor U2300 (N_2300,N_2186,N_2197);
or U2301 (N_2301,N_2179,N_2197);
nor U2302 (N_2302,N_2223,N_2231);
nor U2303 (N_2303,N_2227,N_2224);
xor U2304 (N_2304,N_2240,N_2244);
and U2305 (N_2305,N_2232,N_2226);
nand U2306 (N_2306,N_2227,N_2209);
nor U2307 (N_2307,N_2236,N_2188);
and U2308 (N_2308,N_2206,N_2227);
or U2309 (N_2309,N_2240,N_2229);
and U2310 (N_2310,N_2238,N_2230);
nand U2311 (N_2311,N_2225,N_2195);
or U2312 (N_2312,N_2231,N_2206);
nor U2313 (N_2313,N_2198,N_2203);
nor U2314 (N_2314,N_2233,N_2224);
or U2315 (N_2315,N_2197,N_2238);
nand U2316 (N_2316,N_2177,N_2182);
nand U2317 (N_2317,N_2209,N_2218);
or U2318 (N_2318,N_2215,N_2221);
and U2319 (N_2319,N_2232,N_2203);
xor U2320 (N_2320,N_2241,N_2176);
nor U2321 (N_2321,N_2184,N_2185);
or U2322 (N_2322,N_2200,N_2220);
or U2323 (N_2323,N_2199,N_2212);
or U2324 (N_2324,N_2224,N_2236);
or U2325 (N_2325,N_2253,N_2259);
nor U2326 (N_2326,N_2305,N_2286);
and U2327 (N_2327,N_2300,N_2297);
or U2328 (N_2328,N_2279,N_2304);
or U2329 (N_2329,N_2273,N_2296);
nand U2330 (N_2330,N_2272,N_2282);
nor U2331 (N_2331,N_2261,N_2274);
or U2332 (N_2332,N_2250,N_2291);
or U2333 (N_2333,N_2254,N_2321);
or U2334 (N_2334,N_2320,N_2276);
nand U2335 (N_2335,N_2284,N_2280);
nand U2336 (N_2336,N_2264,N_2319);
nor U2337 (N_2337,N_2313,N_2252);
xnor U2338 (N_2338,N_2256,N_2322);
or U2339 (N_2339,N_2303,N_2307);
nor U2340 (N_2340,N_2324,N_2311);
and U2341 (N_2341,N_2263,N_2294);
and U2342 (N_2342,N_2257,N_2323);
nor U2343 (N_2343,N_2270,N_2308);
nor U2344 (N_2344,N_2306,N_2255);
or U2345 (N_2345,N_2289,N_2283);
and U2346 (N_2346,N_2312,N_2268);
and U2347 (N_2347,N_2260,N_2318);
and U2348 (N_2348,N_2298,N_2251);
or U2349 (N_2349,N_2266,N_2285);
nand U2350 (N_2350,N_2316,N_2262);
or U2351 (N_2351,N_2315,N_2293);
nand U2352 (N_2352,N_2269,N_2309);
nand U2353 (N_2353,N_2275,N_2299);
nor U2354 (N_2354,N_2271,N_2288);
nand U2355 (N_2355,N_2295,N_2258);
xnor U2356 (N_2356,N_2292,N_2277);
xor U2357 (N_2357,N_2317,N_2314);
nand U2358 (N_2358,N_2265,N_2267);
nor U2359 (N_2359,N_2287,N_2290);
xnor U2360 (N_2360,N_2301,N_2281);
nand U2361 (N_2361,N_2310,N_2302);
nor U2362 (N_2362,N_2278,N_2309);
xor U2363 (N_2363,N_2257,N_2288);
or U2364 (N_2364,N_2271,N_2257);
and U2365 (N_2365,N_2295,N_2320);
or U2366 (N_2366,N_2323,N_2315);
and U2367 (N_2367,N_2292,N_2293);
and U2368 (N_2368,N_2265,N_2284);
nand U2369 (N_2369,N_2314,N_2298);
and U2370 (N_2370,N_2319,N_2276);
nor U2371 (N_2371,N_2274,N_2265);
xor U2372 (N_2372,N_2303,N_2290);
nand U2373 (N_2373,N_2258,N_2283);
nand U2374 (N_2374,N_2289,N_2263);
nor U2375 (N_2375,N_2291,N_2257);
and U2376 (N_2376,N_2279,N_2319);
nor U2377 (N_2377,N_2264,N_2252);
and U2378 (N_2378,N_2262,N_2264);
nor U2379 (N_2379,N_2250,N_2307);
nor U2380 (N_2380,N_2298,N_2293);
or U2381 (N_2381,N_2278,N_2269);
nor U2382 (N_2382,N_2258,N_2255);
nand U2383 (N_2383,N_2289,N_2268);
or U2384 (N_2384,N_2305,N_2289);
or U2385 (N_2385,N_2310,N_2299);
nand U2386 (N_2386,N_2290,N_2305);
or U2387 (N_2387,N_2305,N_2295);
or U2388 (N_2388,N_2256,N_2321);
or U2389 (N_2389,N_2280,N_2269);
or U2390 (N_2390,N_2307,N_2297);
or U2391 (N_2391,N_2309,N_2280);
and U2392 (N_2392,N_2292,N_2301);
nand U2393 (N_2393,N_2279,N_2294);
and U2394 (N_2394,N_2298,N_2299);
or U2395 (N_2395,N_2308,N_2293);
nor U2396 (N_2396,N_2282,N_2324);
or U2397 (N_2397,N_2251,N_2264);
and U2398 (N_2398,N_2254,N_2320);
nand U2399 (N_2399,N_2297,N_2310);
nand U2400 (N_2400,N_2395,N_2390);
or U2401 (N_2401,N_2335,N_2329);
nand U2402 (N_2402,N_2381,N_2346);
and U2403 (N_2403,N_2347,N_2398);
nor U2404 (N_2404,N_2341,N_2357);
nand U2405 (N_2405,N_2326,N_2327);
and U2406 (N_2406,N_2325,N_2343);
and U2407 (N_2407,N_2371,N_2367);
or U2408 (N_2408,N_2375,N_2368);
and U2409 (N_2409,N_2364,N_2396);
nor U2410 (N_2410,N_2392,N_2385);
and U2411 (N_2411,N_2344,N_2399);
or U2412 (N_2412,N_2331,N_2382);
nand U2413 (N_2413,N_2360,N_2348);
nand U2414 (N_2414,N_2334,N_2380);
nand U2415 (N_2415,N_2365,N_2351);
or U2416 (N_2416,N_2393,N_2352);
or U2417 (N_2417,N_2362,N_2338);
xor U2418 (N_2418,N_2377,N_2379);
nand U2419 (N_2419,N_2370,N_2342);
nor U2420 (N_2420,N_2328,N_2384);
and U2421 (N_2421,N_2350,N_2391);
nor U2422 (N_2422,N_2374,N_2389);
xnor U2423 (N_2423,N_2356,N_2345);
xor U2424 (N_2424,N_2373,N_2366);
or U2425 (N_2425,N_2397,N_2340);
and U2426 (N_2426,N_2372,N_2330);
and U2427 (N_2427,N_2337,N_2349);
and U2428 (N_2428,N_2353,N_2332);
or U2429 (N_2429,N_2354,N_2376);
and U2430 (N_2430,N_2339,N_2369);
nand U2431 (N_2431,N_2378,N_2361);
nor U2432 (N_2432,N_2358,N_2388);
xor U2433 (N_2433,N_2394,N_2359);
nor U2434 (N_2434,N_2355,N_2387);
nand U2435 (N_2435,N_2333,N_2383);
nand U2436 (N_2436,N_2336,N_2363);
nor U2437 (N_2437,N_2386,N_2369);
nor U2438 (N_2438,N_2398,N_2352);
xnor U2439 (N_2439,N_2396,N_2371);
nand U2440 (N_2440,N_2352,N_2373);
nor U2441 (N_2441,N_2338,N_2391);
nand U2442 (N_2442,N_2335,N_2364);
or U2443 (N_2443,N_2371,N_2385);
and U2444 (N_2444,N_2325,N_2396);
nand U2445 (N_2445,N_2349,N_2393);
nor U2446 (N_2446,N_2359,N_2392);
xor U2447 (N_2447,N_2368,N_2325);
xor U2448 (N_2448,N_2388,N_2368);
nor U2449 (N_2449,N_2373,N_2374);
xor U2450 (N_2450,N_2388,N_2362);
or U2451 (N_2451,N_2330,N_2335);
nor U2452 (N_2452,N_2359,N_2362);
nor U2453 (N_2453,N_2342,N_2390);
nor U2454 (N_2454,N_2365,N_2392);
or U2455 (N_2455,N_2353,N_2345);
nand U2456 (N_2456,N_2360,N_2341);
or U2457 (N_2457,N_2352,N_2350);
nor U2458 (N_2458,N_2349,N_2366);
nor U2459 (N_2459,N_2363,N_2371);
and U2460 (N_2460,N_2393,N_2367);
nand U2461 (N_2461,N_2341,N_2344);
nand U2462 (N_2462,N_2382,N_2378);
and U2463 (N_2463,N_2350,N_2333);
xnor U2464 (N_2464,N_2353,N_2368);
nand U2465 (N_2465,N_2369,N_2382);
and U2466 (N_2466,N_2377,N_2365);
nand U2467 (N_2467,N_2347,N_2373);
nor U2468 (N_2468,N_2383,N_2342);
or U2469 (N_2469,N_2328,N_2337);
nand U2470 (N_2470,N_2351,N_2335);
nand U2471 (N_2471,N_2394,N_2378);
xnor U2472 (N_2472,N_2341,N_2376);
and U2473 (N_2473,N_2366,N_2386);
and U2474 (N_2474,N_2376,N_2334);
and U2475 (N_2475,N_2439,N_2429);
nand U2476 (N_2476,N_2431,N_2420);
or U2477 (N_2477,N_2404,N_2472);
xnor U2478 (N_2478,N_2413,N_2448);
or U2479 (N_2479,N_2453,N_2411);
nor U2480 (N_2480,N_2433,N_2426);
nor U2481 (N_2481,N_2403,N_2418);
nor U2482 (N_2482,N_2467,N_2469);
nor U2483 (N_2483,N_2470,N_2409);
nor U2484 (N_2484,N_2447,N_2461);
or U2485 (N_2485,N_2437,N_2412);
or U2486 (N_2486,N_2444,N_2473);
and U2487 (N_2487,N_2459,N_2424);
and U2488 (N_2488,N_2443,N_2455);
nor U2489 (N_2489,N_2454,N_2425);
or U2490 (N_2490,N_2430,N_2465);
or U2491 (N_2491,N_2457,N_2460);
nor U2492 (N_2492,N_2408,N_2464);
nand U2493 (N_2493,N_2462,N_2442);
nand U2494 (N_2494,N_2449,N_2463);
nand U2495 (N_2495,N_2427,N_2416);
nand U2496 (N_2496,N_2452,N_2428);
nor U2497 (N_2497,N_2474,N_2415);
nor U2498 (N_2498,N_2432,N_2450);
nor U2499 (N_2499,N_2438,N_2446);
or U2500 (N_2500,N_2400,N_2441);
or U2501 (N_2501,N_2419,N_2406);
xnor U2502 (N_2502,N_2422,N_2405);
or U2503 (N_2503,N_2417,N_2456);
or U2504 (N_2504,N_2414,N_2471);
xnor U2505 (N_2505,N_2434,N_2458);
or U2506 (N_2506,N_2410,N_2445);
or U2507 (N_2507,N_2466,N_2402);
or U2508 (N_2508,N_2451,N_2401);
nor U2509 (N_2509,N_2440,N_2435);
and U2510 (N_2510,N_2407,N_2468);
nand U2511 (N_2511,N_2436,N_2421);
and U2512 (N_2512,N_2423,N_2448);
nand U2513 (N_2513,N_2427,N_2466);
xnor U2514 (N_2514,N_2446,N_2440);
and U2515 (N_2515,N_2446,N_2413);
nor U2516 (N_2516,N_2469,N_2468);
or U2517 (N_2517,N_2409,N_2430);
nor U2518 (N_2518,N_2403,N_2432);
nand U2519 (N_2519,N_2415,N_2448);
and U2520 (N_2520,N_2469,N_2407);
and U2521 (N_2521,N_2469,N_2413);
and U2522 (N_2522,N_2402,N_2455);
nand U2523 (N_2523,N_2465,N_2453);
nand U2524 (N_2524,N_2473,N_2468);
or U2525 (N_2525,N_2443,N_2407);
or U2526 (N_2526,N_2452,N_2433);
or U2527 (N_2527,N_2413,N_2471);
nor U2528 (N_2528,N_2441,N_2464);
and U2529 (N_2529,N_2404,N_2471);
nor U2530 (N_2530,N_2443,N_2423);
nor U2531 (N_2531,N_2472,N_2428);
xor U2532 (N_2532,N_2421,N_2400);
or U2533 (N_2533,N_2471,N_2406);
nor U2534 (N_2534,N_2427,N_2445);
nand U2535 (N_2535,N_2441,N_2449);
nor U2536 (N_2536,N_2439,N_2407);
xor U2537 (N_2537,N_2401,N_2404);
xnor U2538 (N_2538,N_2426,N_2460);
or U2539 (N_2539,N_2427,N_2413);
nand U2540 (N_2540,N_2403,N_2469);
nand U2541 (N_2541,N_2411,N_2414);
nand U2542 (N_2542,N_2440,N_2449);
nand U2543 (N_2543,N_2419,N_2403);
and U2544 (N_2544,N_2438,N_2441);
and U2545 (N_2545,N_2439,N_2469);
nand U2546 (N_2546,N_2446,N_2471);
nand U2547 (N_2547,N_2461,N_2450);
nor U2548 (N_2548,N_2447,N_2408);
nor U2549 (N_2549,N_2468,N_2444);
xor U2550 (N_2550,N_2540,N_2514);
or U2551 (N_2551,N_2528,N_2476);
nand U2552 (N_2552,N_2500,N_2527);
nand U2553 (N_2553,N_2522,N_2549);
nor U2554 (N_2554,N_2475,N_2502);
and U2555 (N_2555,N_2525,N_2477);
xor U2556 (N_2556,N_2483,N_2482);
nor U2557 (N_2557,N_2543,N_2490);
xnor U2558 (N_2558,N_2516,N_2536);
or U2559 (N_2559,N_2529,N_2501);
nor U2560 (N_2560,N_2507,N_2491);
and U2561 (N_2561,N_2504,N_2530);
xnor U2562 (N_2562,N_2498,N_2534);
or U2563 (N_2563,N_2524,N_2481);
or U2564 (N_2564,N_2479,N_2486);
and U2565 (N_2565,N_2533,N_2513);
nor U2566 (N_2566,N_2546,N_2485);
nor U2567 (N_2567,N_2545,N_2531);
xnor U2568 (N_2568,N_2532,N_2535);
nand U2569 (N_2569,N_2478,N_2538);
nor U2570 (N_2570,N_2488,N_2519);
nand U2571 (N_2571,N_2518,N_2539);
or U2572 (N_2572,N_2503,N_2541);
and U2573 (N_2573,N_2497,N_2547);
and U2574 (N_2574,N_2484,N_2496);
or U2575 (N_2575,N_2544,N_2520);
and U2576 (N_2576,N_2517,N_2494);
nand U2577 (N_2577,N_2493,N_2510);
nand U2578 (N_2578,N_2489,N_2505);
nor U2579 (N_2579,N_2495,N_2509);
xor U2580 (N_2580,N_2487,N_2508);
or U2581 (N_2581,N_2512,N_2521);
xnor U2582 (N_2582,N_2506,N_2492);
nor U2583 (N_2583,N_2548,N_2480);
nand U2584 (N_2584,N_2523,N_2537);
or U2585 (N_2585,N_2542,N_2511);
nand U2586 (N_2586,N_2526,N_2515);
or U2587 (N_2587,N_2499,N_2546);
or U2588 (N_2588,N_2503,N_2479);
nor U2589 (N_2589,N_2539,N_2504);
and U2590 (N_2590,N_2542,N_2530);
nor U2591 (N_2591,N_2517,N_2525);
nor U2592 (N_2592,N_2547,N_2510);
and U2593 (N_2593,N_2496,N_2537);
and U2594 (N_2594,N_2549,N_2491);
nand U2595 (N_2595,N_2517,N_2501);
nor U2596 (N_2596,N_2506,N_2514);
nand U2597 (N_2597,N_2504,N_2490);
nand U2598 (N_2598,N_2546,N_2535);
nor U2599 (N_2599,N_2539,N_2546);
xor U2600 (N_2600,N_2517,N_2541);
nor U2601 (N_2601,N_2528,N_2534);
nand U2602 (N_2602,N_2521,N_2508);
or U2603 (N_2603,N_2519,N_2477);
and U2604 (N_2604,N_2500,N_2549);
and U2605 (N_2605,N_2487,N_2515);
or U2606 (N_2606,N_2511,N_2496);
and U2607 (N_2607,N_2543,N_2500);
xor U2608 (N_2608,N_2509,N_2534);
nor U2609 (N_2609,N_2487,N_2523);
nand U2610 (N_2610,N_2536,N_2502);
or U2611 (N_2611,N_2486,N_2498);
nand U2612 (N_2612,N_2500,N_2535);
or U2613 (N_2613,N_2529,N_2487);
or U2614 (N_2614,N_2478,N_2521);
xor U2615 (N_2615,N_2485,N_2514);
nor U2616 (N_2616,N_2546,N_2495);
xnor U2617 (N_2617,N_2507,N_2478);
or U2618 (N_2618,N_2530,N_2539);
and U2619 (N_2619,N_2529,N_2512);
nor U2620 (N_2620,N_2513,N_2518);
nor U2621 (N_2621,N_2530,N_2501);
or U2622 (N_2622,N_2531,N_2489);
nor U2623 (N_2623,N_2536,N_2485);
nand U2624 (N_2624,N_2536,N_2549);
nor U2625 (N_2625,N_2618,N_2581);
xor U2626 (N_2626,N_2560,N_2592);
nand U2627 (N_2627,N_2574,N_2616);
and U2628 (N_2628,N_2611,N_2570);
nand U2629 (N_2629,N_2593,N_2569);
xnor U2630 (N_2630,N_2557,N_2621);
nor U2631 (N_2631,N_2580,N_2596);
and U2632 (N_2632,N_2603,N_2575);
xnor U2633 (N_2633,N_2579,N_2588);
nor U2634 (N_2634,N_2553,N_2568);
and U2635 (N_2635,N_2599,N_2615);
nor U2636 (N_2636,N_2619,N_2571);
nor U2637 (N_2637,N_2607,N_2583);
or U2638 (N_2638,N_2598,N_2591);
and U2639 (N_2639,N_2620,N_2595);
or U2640 (N_2640,N_2624,N_2565);
nand U2641 (N_2641,N_2622,N_2556);
or U2642 (N_2642,N_2572,N_2564);
and U2643 (N_2643,N_2601,N_2617);
or U2644 (N_2644,N_2577,N_2563);
and U2645 (N_2645,N_2605,N_2600);
nand U2646 (N_2646,N_2578,N_2555);
or U2647 (N_2647,N_2608,N_2566);
nand U2648 (N_2648,N_2606,N_2561);
xor U2649 (N_2649,N_2602,N_2576);
or U2650 (N_2650,N_2554,N_2551);
nand U2651 (N_2651,N_2573,N_2558);
and U2652 (N_2652,N_2552,N_2597);
and U2653 (N_2653,N_2567,N_2623);
or U2654 (N_2654,N_2587,N_2585);
or U2655 (N_2655,N_2584,N_2562);
nand U2656 (N_2656,N_2613,N_2589);
or U2657 (N_2657,N_2550,N_2609);
xnor U2658 (N_2658,N_2559,N_2612);
or U2659 (N_2659,N_2586,N_2604);
nor U2660 (N_2660,N_2582,N_2614);
or U2661 (N_2661,N_2594,N_2610);
nand U2662 (N_2662,N_2590,N_2584);
or U2663 (N_2663,N_2566,N_2571);
or U2664 (N_2664,N_2562,N_2556);
nor U2665 (N_2665,N_2563,N_2602);
nand U2666 (N_2666,N_2572,N_2553);
nand U2667 (N_2667,N_2596,N_2610);
nor U2668 (N_2668,N_2559,N_2580);
or U2669 (N_2669,N_2594,N_2597);
nor U2670 (N_2670,N_2580,N_2618);
nor U2671 (N_2671,N_2617,N_2598);
nor U2672 (N_2672,N_2601,N_2620);
nand U2673 (N_2673,N_2622,N_2573);
or U2674 (N_2674,N_2577,N_2554);
nor U2675 (N_2675,N_2580,N_2622);
or U2676 (N_2676,N_2572,N_2606);
or U2677 (N_2677,N_2574,N_2557);
nor U2678 (N_2678,N_2569,N_2550);
and U2679 (N_2679,N_2563,N_2600);
or U2680 (N_2680,N_2582,N_2603);
or U2681 (N_2681,N_2568,N_2617);
or U2682 (N_2682,N_2579,N_2603);
or U2683 (N_2683,N_2590,N_2553);
nand U2684 (N_2684,N_2595,N_2622);
or U2685 (N_2685,N_2561,N_2550);
nand U2686 (N_2686,N_2624,N_2591);
nand U2687 (N_2687,N_2550,N_2572);
and U2688 (N_2688,N_2569,N_2565);
and U2689 (N_2689,N_2574,N_2598);
and U2690 (N_2690,N_2611,N_2594);
or U2691 (N_2691,N_2609,N_2603);
nand U2692 (N_2692,N_2563,N_2620);
and U2693 (N_2693,N_2577,N_2616);
nand U2694 (N_2694,N_2585,N_2609);
or U2695 (N_2695,N_2610,N_2614);
nand U2696 (N_2696,N_2581,N_2552);
nand U2697 (N_2697,N_2562,N_2576);
or U2698 (N_2698,N_2605,N_2586);
and U2699 (N_2699,N_2550,N_2595);
and U2700 (N_2700,N_2675,N_2636);
or U2701 (N_2701,N_2649,N_2633);
nor U2702 (N_2702,N_2647,N_2638);
or U2703 (N_2703,N_2678,N_2682);
or U2704 (N_2704,N_2660,N_2658);
xor U2705 (N_2705,N_2690,N_2674);
or U2706 (N_2706,N_2641,N_2696);
nand U2707 (N_2707,N_2694,N_2666);
xor U2708 (N_2708,N_2671,N_2639);
and U2709 (N_2709,N_2688,N_2626);
nand U2710 (N_2710,N_2662,N_2625);
or U2711 (N_2711,N_2655,N_2683);
and U2712 (N_2712,N_2648,N_2691);
and U2713 (N_2713,N_2680,N_2653);
and U2714 (N_2714,N_2686,N_2640);
nand U2715 (N_2715,N_2664,N_2650);
and U2716 (N_2716,N_2663,N_2681);
xor U2717 (N_2717,N_2697,N_2657);
nor U2718 (N_2718,N_2661,N_2668);
or U2719 (N_2719,N_2642,N_2687);
xor U2720 (N_2720,N_2669,N_2654);
and U2721 (N_2721,N_2645,N_2635);
and U2722 (N_2722,N_2679,N_2665);
nand U2723 (N_2723,N_2646,N_2689);
nor U2724 (N_2724,N_2667,N_2634);
and U2725 (N_2725,N_2698,N_2628);
nand U2726 (N_2726,N_2693,N_2637);
xor U2727 (N_2727,N_2629,N_2630);
nand U2728 (N_2728,N_2673,N_2627);
or U2729 (N_2729,N_2692,N_2672);
nand U2730 (N_2730,N_2632,N_2651);
nor U2731 (N_2731,N_2676,N_2685);
and U2732 (N_2732,N_2652,N_2644);
and U2733 (N_2733,N_2677,N_2699);
nand U2734 (N_2734,N_2659,N_2631);
xor U2735 (N_2735,N_2684,N_2656);
nor U2736 (N_2736,N_2643,N_2695);
xor U2737 (N_2737,N_2670,N_2674);
nand U2738 (N_2738,N_2678,N_2655);
nor U2739 (N_2739,N_2630,N_2692);
and U2740 (N_2740,N_2669,N_2638);
and U2741 (N_2741,N_2658,N_2634);
nand U2742 (N_2742,N_2693,N_2669);
nor U2743 (N_2743,N_2654,N_2660);
xnor U2744 (N_2744,N_2636,N_2682);
nor U2745 (N_2745,N_2660,N_2646);
or U2746 (N_2746,N_2635,N_2649);
or U2747 (N_2747,N_2650,N_2682);
xor U2748 (N_2748,N_2627,N_2657);
nand U2749 (N_2749,N_2631,N_2676);
nand U2750 (N_2750,N_2674,N_2630);
and U2751 (N_2751,N_2666,N_2649);
nor U2752 (N_2752,N_2684,N_2626);
nand U2753 (N_2753,N_2637,N_2670);
and U2754 (N_2754,N_2638,N_2639);
or U2755 (N_2755,N_2648,N_2647);
xor U2756 (N_2756,N_2625,N_2633);
or U2757 (N_2757,N_2640,N_2634);
nand U2758 (N_2758,N_2676,N_2694);
nand U2759 (N_2759,N_2648,N_2681);
nand U2760 (N_2760,N_2649,N_2696);
or U2761 (N_2761,N_2636,N_2654);
nor U2762 (N_2762,N_2654,N_2638);
nand U2763 (N_2763,N_2695,N_2650);
or U2764 (N_2764,N_2684,N_2665);
and U2765 (N_2765,N_2697,N_2669);
or U2766 (N_2766,N_2655,N_2671);
and U2767 (N_2767,N_2688,N_2650);
nor U2768 (N_2768,N_2647,N_2688);
nor U2769 (N_2769,N_2635,N_2636);
nand U2770 (N_2770,N_2655,N_2680);
or U2771 (N_2771,N_2658,N_2684);
nor U2772 (N_2772,N_2655,N_2662);
and U2773 (N_2773,N_2676,N_2644);
nand U2774 (N_2774,N_2696,N_2674);
and U2775 (N_2775,N_2714,N_2732);
nor U2776 (N_2776,N_2741,N_2747);
nor U2777 (N_2777,N_2722,N_2752);
xor U2778 (N_2778,N_2721,N_2706);
nor U2779 (N_2779,N_2761,N_2719);
and U2780 (N_2780,N_2708,N_2758);
nand U2781 (N_2781,N_2715,N_2713);
or U2782 (N_2782,N_2772,N_2737);
or U2783 (N_2783,N_2759,N_2764);
xnor U2784 (N_2784,N_2704,N_2762);
nor U2785 (N_2785,N_2733,N_2736);
nor U2786 (N_2786,N_2724,N_2743);
or U2787 (N_2787,N_2744,N_2768);
and U2788 (N_2788,N_2730,N_2757);
or U2789 (N_2789,N_2739,N_2771);
xor U2790 (N_2790,N_2725,N_2734);
xor U2791 (N_2791,N_2750,N_2773);
nor U2792 (N_2792,N_2702,N_2746);
and U2793 (N_2793,N_2738,N_2769);
and U2794 (N_2794,N_2735,N_2770);
or U2795 (N_2795,N_2710,N_2727);
and U2796 (N_2796,N_2700,N_2717);
nand U2797 (N_2797,N_2745,N_2774);
nand U2798 (N_2798,N_2754,N_2716);
xor U2799 (N_2799,N_2740,N_2749);
nor U2800 (N_2800,N_2705,N_2763);
and U2801 (N_2801,N_2711,N_2728);
or U2802 (N_2802,N_2765,N_2767);
nand U2803 (N_2803,N_2729,N_2731);
nand U2804 (N_2804,N_2718,N_2753);
nor U2805 (N_2805,N_2723,N_2755);
or U2806 (N_2806,N_2751,N_2748);
xor U2807 (N_2807,N_2742,N_2707);
nor U2808 (N_2808,N_2726,N_2760);
nor U2809 (N_2809,N_2709,N_2701);
nand U2810 (N_2810,N_2756,N_2712);
or U2811 (N_2811,N_2703,N_2720);
nor U2812 (N_2812,N_2766,N_2735);
or U2813 (N_2813,N_2723,N_2761);
and U2814 (N_2814,N_2713,N_2751);
nand U2815 (N_2815,N_2761,N_2712);
nand U2816 (N_2816,N_2725,N_2750);
nand U2817 (N_2817,N_2772,N_2715);
nor U2818 (N_2818,N_2756,N_2720);
xnor U2819 (N_2819,N_2751,N_2739);
and U2820 (N_2820,N_2758,N_2770);
nand U2821 (N_2821,N_2757,N_2719);
nor U2822 (N_2822,N_2725,N_2721);
nand U2823 (N_2823,N_2717,N_2772);
or U2824 (N_2824,N_2735,N_2743);
nor U2825 (N_2825,N_2750,N_2728);
and U2826 (N_2826,N_2724,N_2721);
nand U2827 (N_2827,N_2705,N_2715);
or U2828 (N_2828,N_2728,N_2703);
nand U2829 (N_2829,N_2739,N_2719);
or U2830 (N_2830,N_2769,N_2720);
nand U2831 (N_2831,N_2729,N_2746);
xor U2832 (N_2832,N_2765,N_2718);
nor U2833 (N_2833,N_2720,N_2773);
nor U2834 (N_2834,N_2744,N_2715);
nor U2835 (N_2835,N_2774,N_2726);
or U2836 (N_2836,N_2763,N_2736);
and U2837 (N_2837,N_2718,N_2701);
or U2838 (N_2838,N_2774,N_2746);
xor U2839 (N_2839,N_2725,N_2745);
and U2840 (N_2840,N_2708,N_2744);
or U2841 (N_2841,N_2741,N_2704);
and U2842 (N_2842,N_2709,N_2761);
nand U2843 (N_2843,N_2754,N_2720);
and U2844 (N_2844,N_2753,N_2743);
nor U2845 (N_2845,N_2761,N_2717);
nor U2846 (N_2846,N_2745,N_2737);
nand U2847 (N_2847,N_2756,N_2761);
nand U2848 (N_2848,N_2748,N_2712);
nor U2849 (N_2849,N_2737,N_2751);
or U2850 (N_2850,N_2838,N_2842);
nand U2851 (N_2851,N_2830,N_2804);
or U2852 (N_2852,N_2841,N_2840);
or U2853 (N_2853,N_2777,N_2833);
and U2854 (N_2854,N_2835,N_2813);
and U2855 (N_2855,N_2825,N_2816);
and U2856 (N_2856,N_2798,N_2844);
xnor U2857 (N_2857,N_2789,N_2809);
and U2858 (N_2858,N_2783,N_2800);
and U2859 (N_2859,N_2826,N_2802);
and U2860 (N_2860,N_2812,N_2803);
nor U2861 (N_2861,N_2815,N_2822);
nor U2862 (N_2862,N_2821,N_2849);
nor U2863 (N_2863,N_2820,N_2787);
nor U2864 (N_2864,N_2778,N_2801);
nor U2865 (N_2865,N_2831,N_2775);
or U2866 (N_2866,N_2827,N_2847);
and U2867 (N_2867,N_2780,N_2814);
and U2868 (N_2868,N_2781,N_2819);
nand U2869 (N_2869,N_2790,N_2799);
and U2870 (N_2870,N_2795,N_2823);
nand U2871 (N_2871,N_2811,N_2794);
and U2872 (N_2872,N_2834,N_2796);
xor U2873 (N_2873,N_2805,N_2791);
and U2874 (N_2874,N_2784,N_2793);
nor U2875 (N_2875,N_2782,N_2845);
nand U2876 (N_2876,N_2848,N_2808);
nor U2877 (N_2877,N_2776,N_2817);
and U2878 (N_2878,N_2786,N_2824);
xor U2879 (N_2879,N_2846,N_2837);
nor U2880 (N_2880,N_2785,N_2807);
or U2881 (N_2881,N_2797,N_2836);
and U2882 (N_2882,N_2843,N_2832);
nor U2883 (N_2883,N_2806,N_2829);
or U2884 (N_2884,N_2792,N_2828);
and U2885 (N_2885,N_2788,N_2810);
nor U2886 (N_2886,N_2779,N_2839);
or U2887 (N_2887,N_2818,N_2795);
nor U2888 (N_2888,N_2827,N_2783);
nor U2889 (N_2889,N_2801,N_2792);
nand U2890 (N_2890,N_2827,N_2795);
nand U2891 (N_2891,N_2831,N_2816);
nand U2892 (N_2892,N_2814,N_2823);
nand U2893 (N_2893,N_2780,N_2832);
nor U2894 (N_2894,N_2776,N_2842);
nor U2895 (N_2895,N_2813,N_2785);
nor U2896 (N_2896,N_2797,N_2845);
or U2897 (N_2897,N_2787,N_2818);
xnor U2898 (N_2898,N_2799,N_2809);
nor U2899 (N_2899,N_2822,N_2798);
nand U2900 (N_2900,N_2776,N_2780);
nand U2901 (N_2901,N_2814,N_2793);
and U2902 (N_2902,N_2822,N_2829);
nand U2903 (N_2903,N_2831,N_2818);
xor U2904 (N_2904,N_2835,N_2802);
or U2905 (N_2905,N_2778,N_2789);
nor U2906 (N_2906,N_2843,N_2803);
nand U2907 (N_2907,N_2808,N_2788);
nand U2908 (N_2908,N_2827,N_2814);
and U2909 (N_2909,N_2820,N_2779);
nand U2910 (N_2910,N_2825,N_2848);
nor U2911 (N_2911,N_2826,N_2791);
xnor U2912 (N_2912,N_2842,N_2790);
xor U2913 (N_2913,N_2818,N_2820);
or U2914 (N_2914,N_2790,N_2845);
nand U2915 (N_2915,N_2816,N_2839);
or U2916 (N_2916,N_2807,N_2814);
nand U2917 (N_2917,N_2776,N_2830);
xnor U2918 (N_2918,N_2842,N_2807);
or U2919 (N_2919,N_2783,N_2834);
xor U2920 (N_2920,N_2842,N_2786);
and U2921 (N_2921,N_2777,N_2849);
and U2922 (N_2922,N_2808,N_2777);
xnor U2923 (N_2923,N_2792,N_2834);
and U2924 (N_2924,N_2789,N_2788);
nor U2925 (N_2925,N_2873,N_2881);
nor U2926 (N_2926,N_2916,N_2851);
or U2927 (N_2927,N_2898,N_2871);
nand U2928 (N_2928,N_2866,N_2854);
xor U2929 (N_2929,N_2909,N_2895);
nand U2930 (N_2930,N_2914,N_2877);
nand U2931 (N_2931,N_2906,N_2903);
and U2932 (N_2932,N_2870,N_2872);
and U2933 (N_2933,N_2856,N_2853);
nor U2934 (N_2934,N_2894,N_2864);
nand U2935 (N_2935,N_2915,N_2850);
and U2936 (N_2936,N_2885,N_2858);
and U2937 (N_2937,N_2922,N_2918);
xor U2938 (N_2938,N_2889,N_2892);
and U2939 (N_2939,N_2876,N_2917);
and U2940 (N_2940,N_2907,N_2857);
nor U2941 (N_2941,N_2861,N_2896);
nor U2942 (N_2942,N_2878,N_2880);
nor U2943 (N_2943,N_2919,N_2882);
and U2944 (N_2944,N_2887,N_2899);
nand U2945 (N_2945,N_2904,N_2921);
or U2946 (N_2946,N_2893,N_2890);
and U2947 (N_2947,N_2900,N_2908);
nand U2948 (N_2948,N_2891,N_2855);
nor U2949 (N_2949,N_2863,N_2883);
and U2950 (N_2950,N_2862,N_2905);
and U2951 (N_2951,N_2913,N_2875);
nand U2952 (N_2952,N_2874,N_2879);
and U2953 (N_2953,N_2869,N_2912);
nor U2954 (N_2954,N_2852,N_2884);
xnor U2955 (N_2955,N_2888,N_2859);
or U2956 (N_2956,N_2860,N_2923);
and U2957 (N_2957,N_2911,N_2920);
and U2958 (N_2958,N_2901,N_2924);
nand U2959 (N_2959,N_2886,N_2868);
and U2960 (N_2960,N_2897,N_2902);
nand U2961 (N_2961,N_2865,N_2867);
and U2962 (N_2962,N_2910,N_2880);
or U2963 (N_2963,N_2859,N_2886);
or U2964 (N_2964,N_2908,N_2890);
nand U2965 (N_2965,N_2916,N_2910);
nand U2966 (N_2966,N_2861,N_2894);
and U2967 (N_2967,N_2920,N_2916);
nor U2968 (N_2968,N_2905,N_2869);
and U2969 (N_2969,N_2898,N_2890);
and U2970 (N_2970,N_2895,N_2886);
and U2971 (N_2971,N_2890,N_2868);
nand U2972 (N_2972,N_2864,N_2909);
nor U2973 (N_2973,N_2882,N_2854);
or U2974 (N_2974,N_2910,N_2850);
nor U2975 (N_2975,N_2872,N_2883);
nand U2976 (N_2976,N_2897,N_2891);
nor U2977 (N_2977,N_2893,N_2871);
nand U2978 (N_2978,N_2855,N_2864);
and U2979 (N_2979,N_2856,N_2885);
nand U2980 (N_2980,N_2886,N_2908);
or U2981 (N_2981,N_2898,N_2869);
nor U2982 (N_2982,N_2908,N_2921);
or U2983 (N_2983,N_2902,N_2875);
and U2984 (N_2984,N_2917,N_2882);
and U2985 (N_2985,N_2855,N_2879);
nor U2986 (N_2986,N_2921,N_2912);
or U2987 (N_2987,N_2875,N_2888);
nand U2988 (N_2988,N_2901,N_2904);
nand U2989 (N_2989,N_2890,N_2879);
nand U2990 (N_2990,N_2890,N_2918);
and U2991 (N_2991,N_2891,N_2895);
nand U2992 (N_2992,N_2906,N_2871);
nand U2993 (N_2993,N_2894,N_2893);
xnor U2994 (N_2994,N_2897,N_2904);
and U2995 (N_2995,N_2893,N_2888);
and U2996 (N_2996,N_2884,N_2916);
and U2997 (N_2997,N_2893,N_2881);
nand U2998 (N_2998,N_2863,N_2921);
nor U2999 (N_2999,N_2898,N_2892);
or UO_0 (O_0,N_2929,N_2982);
and UO_1 (O_1,N_2957,N_2960);
or UO_2 (O_2,N_2954,N_2940);
or UO_3 (O_3,N_2948,N_2934);
nor UO_4 (O_4,N_2980,N_2993);
and UO_5 (O_5,N_2959,N_2943);
and UO_6 (O_6,N_2998,N_2931);
nand UO_7 (O_7,N_2981,N_2997);
xor UO_8 (O_8,N_2994,N_2953);
and UO_9 (O_9,N_2933,N_2937);
and UO_10 (O_10,N_2946,N_2963);
and UO_11 (O_11,N_2927,N_2955);
nor UO_12 (O_12,N_2930,N_2925);
and UO_13 (O_13,N_2991,N_2999);
nor UO_14 (O_14,N_2990,N_2966);
xnor UO_15 (O_15,N_2988,N_2978);
nor UO_16 (O_16,N_2974,N_2992);
or UO_17 (O_17,N_2949,N_2951);
xnor UO_18 (O_18,N_2989,N_2945);
nor UO_19 (O_19,N_2969,N_2944);
nand UO_20 (O_20,N_2975,N_2965);
or UO_21 (O_21,N_2950,N_2926);
or UO_22 (O_22,N_2986,N_2958);
nand UO_23 (O_23,N_2936,N_2983);
nor UO_24 (O_24,N_2996,N_2939);
and UO_25 (O_25,N_2961,N_2942);
or UO_26 (O_26,N_2952,N_2932);
and UO_27 (O_27,N_2970,N_2956);
or UO_28 (O_28,N_2968,N_2977);
or UO_29 (O_29,N_2928,N_2985);
and UO_30 (O_30,N_2947,N_2976);
nand UO_31 (O_31,N_2972,N_2962);
nand UO_32 (O_32,N_2973,N_2964);
or UO_33 (O_33,N_2979,N_2995);
or UO_34 (O_34,N_2941,N_2984);
and UO_35 (O_35,N_2935,N_2971);
nand UO_36 (O_36,N_2967,N_2938);
nor UO_37 (O_37,N_2987,N_2958);
and UO_38 (O_38,N_2941,N_2926);
nor UO_39 (O_39,N_2926,N_2956);
nor UO_40 (O_40,N_2971,N_2967);
xor UO_41 (O_41,N_2956,N_2954);
nor UO_42 (O_42,N_2926,N_2953);
and UO_43 (O_43,N_2927,N_2973);
or UO_44 (O_44,N_2932,N_2933);
and UO_45 (O_45,N_2965,N_2963);
or UO_46 (O_46,N_2957,N_2982);
and UO_47 (O_47,N_2951,N_2945);
nor UO_48 (O_48,N_2995,N_2938);
nor UO_49 (O_49,N_2996,N_2945);
nand UO_50 (O_50,N_2998,N_2938);
nor UO_51 (O_51,N_2957,N_2937);
nand UO_52 (O_52,N_2940,N_2969);
nor UO_53 (O_53,N_2956,N_2987);
nand UO_54 (O_54,N_2939,N_2955);
nor UO_55 (O_55,N_2952,N_2954);
or UO_56 (O_56,N_2940,N_2945);
or UO_57 (O_57,N_2993,N_2985);
nor UO_58 (O_58,N_2974,N_2998);
or UO_59 (O_59,N_2995,N_2966);
and UO_60 (O_60,N_2938,N_2962);
nand UO_61 (O_61,N_2958,N_2992);
xor UO_62 (O_62,N_2991,N_2956);
or UO_63 (O_63,N_2957,N_2963);
nand UO_64 (O_64,N_2951,N_2994);
and UO_65 (O_65,N_2957,N_2948);
nand UO_66 (O_66,N_2971,N_2960);
nand UO_67 (O_67,N_2989,N_2963);
and UO_68 (O_68,N_2934,N_2942);
and UO_69 (O_69,N_2989,N_2955);
and UO_70 (O_70,N_2994,N_2982);
and UO_71 (O_71,N_2945,N_2928);
or UO_72 (O_72,N_2926,N_2981);
or UO_73 (O_73,N_2996,N_2953);
nand UO_74 (O_74,N_2973,N_2929);
or UO_75 (O_75,N_2964,N_2989);
or UO_76 (O_76,N_2939,N_2966);
nor UO_77 (O_77,N_2967,N_2969);
xnor UO_78 (O_78,N_2951,N_2963);
and UO_79 (O_79,N_2950,N_2933);
and UO_80 (O_80,N_2973,N_2965);
or UO_81 (O_81,N_2942,N_2997);
and UO_82 (O_82,N_2935,N_2990);
or UO_83 (O_83,N_2991,N_2980);
xor UO_84 (O_84,N_2961,N_2983);
or UO_85 (O_85,N_2952,N_2979);
and UO_86 (O_86,N_2969,N_2996);
or UO_87 (O_87,N_2938,N_2984);
nor UO_88 (O_88,N_2960,N_2999);
or UO_89 (O_89,N_2963,N_2994);
nand UO_90 (O_90,N_2997,N_2995);
nor UO_91 (O_91,N_2959,N_2990);
or UO_92 (O_92,N_2998,N_2973);
or UO_93 (O_93,N_2943,N_2982);
nor UO_94 (O_94,N_2999,N_2933);
or UO_95 (O_95,N_2952,N_2950);
nand UO_96 (O_96,N_2952,N_2930);
xnor UO_97 (O_97,N_2943,N_2996);
nor UO_98 (O_98,N_2964,N_2938);
and UO_99 (O_99,N_2995,N_2967);
xnor UO_100 (O_100,N_2988,N_2945);
or UO_101 (O_101,N_2964,N_2958);
and UO_102 (O_102,N_2995,N_2980);
and UO_103 (O_103,N_2938,N_2989);
xor UO_104 (O_104,N_2985,N_2995);
nand UO_105 (O_105,N_2992,N_2959);
or UO_106 (O_106,N_2972,N_2946);
nor UO_107 (O_107,N_2952,N_2962);
nor UO_108 (O_108,N_2995,N_2957);
nor UO_109 (O_109,N_2988,N_2942);
and UO_110 (O_110,N_2961,N_2977);
or UO_111 (O_111,N_2935,N_2961);
and UO_112 (O_112,N_2964,N_2929);
or UO_113 (O_113,N_2998,N_2976);
or UO_114 (O_114,N_2958,N_2928);
nor UO_115 (O_115,N_2981,N_2931);
nor UO_116 (O_116,N_2981,N_2965);
or UO_117 (O_117,N_2988,N_2964);
and UO_118 (O_118,N_2992,N_2998);
and UO_119 (O_119,N_2996,N_2978);
or UO_120 (O_120,N_2990,N_2939);
and UO_121 (O_121,N_2996,N_2948);
nor UO_122 (O_122,N_2959,N_2965);
nand UO_123 (O_123,N_2998,N_2949);
nand UO_124 (O_124,N_2964,N_2996);
nand UO_125 (O_125,N_2958,N_2974);
nor UO_126 (O_126,N_2938,N_2969);
or UO_127 (O_127,N_2945,N_2927);
xor UO_128 (O_128,N_2957,N_2964);
and UO_129 (O_129,N_2974,N_2932);
nand UO_130 (O_130,N_2994,N_2991);
nand UO_131 (O_131,N_2984,N_2958);
nand UO_132 (O_132,N_2942,N_2975);
or UO_133 (O_133,N_2925,N_2963);
nand UO_134 (O_134,N_2984,N_2928);
and UO_135 (O_135,N_2989,N_2941);
and UO_136 (O_136,N_2945,N_2964);
and UO_137 (O_137,N_2963,N_2970);
or UO_138 (O_138,N_2960,N_2981);
and UO_139 (O_139,N_2995,N_2971);
or UO_140 (O_140,N_2965,N_2934);
nand UO_141 (O_141,N_2955,N_2938);
or UO_142 (O_142,N_2953,N_2927);
nor UO_143 (O_143,N_2962,N_2993);
nor UO_144 (O_144,N_2933,N_2951);
or UO_145 (O_145,N_2985,N_2979);
nor UO_146 (O_146,N_2959,N_2947);
xor UO_147 (O_147,N_2995,N_2976);
nor UO_148 (O_148,N_2990,N_2982);
nand UO_149 (O_149,N_2953,N_2992);
and UO_150 (O_150,N_2985,N_2981);
or UO_151 (O_151,N_2934,N_2989);
and UO_152 (O_152,N_2949,N_2968);
nand UO_153 (O_153,N_2961,N_2927);
nor UO_154 (O_154,N_2947,N_2952);
nor UO_155 (O_155,N_2973,N_2969);
xnor UO_156 (O_156,N_2993,N_2972);
and UO_157 (O_157,N_2990,N_2942);
nor UO_158 (O_158,N_2975,N_2978);
nand UO_159 (O_159,N_2968,N_2980);
xor UO_160 (O_160,N_2940,N_2936);
nor UO_161 (O_161,N_2973,N_2962);
or UO_162 (O_162,N_2958,N_2982);
nor UO_163 (O_163,N_2937,N_2978);
nor UO_164 (O_164,N_2928,N_2943);
nor UO_165 (O_165,N_2927,N_2942);
nor UO_166 (O_166,N_2976,N_2953);
and UO_167 (O_167,N_2955,N_2935);
nor UO_168 (O_168,N_2976,N_2941);
and UO_169 (O_169,N_2994,N_2926);
xnor UO_170 (O_170,N_2930,N_2947);
and UO_171 (O_171,N_2981,N_2982);
nor UO_172 (O_172,N_2980,N_2947);
nor UO_173 (O_173,N_2966,N_2925);
or UO_174 (O_174,N_2972,N_2982);
and UO_175 (O_175,N_2944,N_2979);
nor UO_176 (O_176,N_2947,N_2942);
nand UO_177 (O_177,N_2959,N_2940);
and UO_178 (O_178,N_2977,N_2943);
nor UO_179 (O_179,N_2952,N_2963);
and UO_180 (O_180,N_2927,N_2964);
nor UO_181 (O_181,N_2977,N_2981);
nand UO_182 (O_182,N_2988,N_2991);
nor UO_183 (O_183,N_2972,N_2942);
nor UO_184 (O_184,N_2956,N_2998);
or UO_185 (O_185,N_2953,N_2999);
or UO_186 (O_186,N_2982,N_2934);
nand UO_187 (O_187,N_2962,N_2932);
xor UO_188 (O_188,N_2963,N_2991);
or UO_189 (O_189,N_2947,N_2982);
and UO_190 (O_190,N_2990,N_2994);
nor UO_191 (O_191,N_2975,N_2992);
nor UO_192 (O_192,N_2995,N_2945);
or UO_193 (O_193,N_2967,N_2986);
xor UO_194 (O_194,N_2940,N_2942);
xor UO_195 (O_195,N_2990,N_2962);
nor UO_196 (O_196,N_2957,N_2928);
nor UO_197 (O_197,N_2962,N_2984);
nand UO_198 (O_198,N_2952,N_2989);
nand UO_199 (O_199,N_2965,N_2993);
nor UO_200 (O_200,N_2979,N_2958);
and UO_201 (O_201,N_2938,N_2977);
or UO_202 (O_202,N_2977,N_2953);
nor UO_203 (O_203,N_2977,N_2988);
nor UO_204 (O_204,N_2935,N_2981);
and UO_205 (O_205,N_2967,N_2972);
nor UO_206 (O_206,N_2960,N_2962);
xnor UO_207 (O_207,N_2981,N_2999);
nor UO_208 (O_208,N_2949,N_2937);
nor UO_209 (O_209,N_2926,N_2951);
or UO_210 (O_210,N_2960,N_2961);
and UO_211 (O_211,N_2988,N_2956);
and UO_212 (O_212,N_2928,N_2983);
and UO_213 (O_213,N_2964,N_2970);
and UO_214 (O_214,N_2967,N_2999);
nor UO_215 (O_215,N_2929,N_2950);
nor UO_216 (O_216,N_2986,N_2977);
nor UO_217 (O_217,N_2965,N_2971);
or UO_218 (O_218,N_2996,N_2942);
and UO_219 (O_219,N_2957,N_2946);
nand UO_220 (O_220,N_2989,N_2987);
nor UO_221 (O_221,N_2930,N_2954);
xnor UO_222 (O_222,N_2980,N_2930);
nor UO_223 (O_223,N_2943,N_2929);
nand UO_224 (O_224,N_2981,N_2937);
and UO_225 (O_225,N_2934,N_2964);
nand UO_226 (O_226,N_2932,N_2958);
nor UO_227 (O_227,N_2997,N_2944);
xnor UO_228 (O_228,N_2943,N_2949);
nand UO_229 (O_229,N_2945,N_2992);
xor UO_230 (O_230,N_2951,N_2952);
nor UO_231 (O_231,N_2990,N_2927);
nor UO_232 (O_232,N_2976,N_2971);
or UO_233 (O_233,N_2991,N_2975);
nor UO_234 (O_234,N_2979,N_2989);
or UO_235 (O_235,N_2982,N_2928);
and UO_236 (O_236,N_2930,N_2944);
nor UO_237 (O_237,N_2958,N_2947);
and UO_238 (O_238,N_2958,N_2991);
xor UO_239 (O_239,N_2940,N_2964);
and UO_240 (O_240,N_2946,N_2981);
nor UO_241 (O_241,N_2959,N_2984);
or UO_242 (O_242,N_2935,N_2977);
nand UO_243 (O_243,N_2969,N_2939);
nand UO_244 (O_244,N_2966,N_2974);
nor UO_245 (O_245,N_2970,N_2952);
nor UO_246 (O_246,N_2997,N_2950);
or UO_247 (O_247,N_2930,N_2938);
and UO_248 (O_248,N_2978,N_2963);
nor UO_249 (O_249,N_2998,N_2975);
xor UO_250 (O_250,N_2938,N_2936);
and UO_251 (O_251,N_2940,N_2985);
or UO_252 (O_252,N_2992,N_2997);
nand UO_253 (O_253,N_2932,N_2950);
or UO_254 (O_254,N_2963,N_2975);
or UO_255 (O_255,N_2930,N_2939);
nor UO_256 (O_256,N_2969,N_2954);
and UO_257 (O_257,N_2926,N_2949);
or UO_258 (O_258,N_2957,N_2972);
or UO_259 (O_259,N_2939,N_2975);
or UO_260 (O_260,N_2942,N_2932);
or UO_261 (O_261,N_2960,N_2956);
nor UO_262 (O_262,N_2944,N_2996);
or UO_263 (O_263,N_2990,N_2969);
nor UO_264 (O_264,N_2967,N_2982);
or UO_265 (O_265,N_2955,N_2995);
nor UO_266 (O_266,N_2932,N_2992);
and UO_267 (O_267,N_2984,N_2936);
or UO_268 (O_268,N_2988,N_2951);
nor UO_269 (O_269,N_2966,N_2926);
or UO_270 (O_270,N_2930,N_2976);
nand UO_271 (O_271,N_2994,N_2998);
nor UO_272 (O_272,N_2984,N_2969);
and UO_273 (O_273,N_2978,N_2964);
and UO_274 (O_274,N_2930,N_2933);
or UO_275 (O_275,N_2986,N_2979);
nand UO_276 (O_276,N_2941,N_2960);
nor UO_277 (O_277,N_2931,N_2966);
xor UO_278 (O_278,N_2963,N_2981);
nor UO_279 (O_279,N_2963,N_2928);
xor UO_280 (O_280,N_2929,N_2984);
and UO_281 (O_281,N_2987,N_2952);
nor UO_282 (O_282,N_2969,N_2953);
or UO_283 (O_283,N_2984,N_2982);
nor UO_284 (O_284,N_2997,N_2965);
or UO_285 (O_285,N_2998,N_2932);
or UO_286 (O_286,N_2934,N_2971);
and UO_287 (O_287,N_2998,N_2962);
and UO_288 (O_288,N_2963,N_2958);
and UO_289 (O_289,N_2926,N_2984);
and UO_290 (O_290,N_2930,N_2955);
nand UO_291 (O_291,N_2985,N_2980);
and UO_292 (O_292,N_2931,N_2944);
and UO_293 (O_293,N_2995,N_2954);
xnor UO_294 (O_294,N_2962,N_2983);
nor UO_295 (O_295,N_2947,N_2979);
or UO_296 (O_296,N_2978,N_2989);
nand UO_297 (O_297,N_2928,N_2995);
nand UO_298 (O_298,N_2974,N_2928);
nand UO_299 (O_299,N_2927,N_2972);
and UO_300 (O_300,N_2957,N_2975);
xor UO_301 (O_301,N_2971,N_2981);
nand UO_302 (O_302,N_2951,N_2992);
nor UO_303 (O_303,N_2977,N_2958);
nand UO_304 (O_304,N_2930,N_2973);
and UO_305 (O_305,N_2942,N_2939);
or UO_306 (O_306,N_2956,N_2985);
and UO_307 (O_307,N_2952,N_2931);
nor UO_308 (O_308,N_2997,N_2959);
nand UO_309 (O_309,N_2961,N_2968);
nor UO_310 (O_310,N_2973,N_2944);
nor UO_311 (O_311,N_2981,N_2945);
and UO_312 (O_312,N_2999,N_2969);
nor UO_313 (O_313,N_2965,N_2938);
nand UO_314 (O_314,N_2993,N_2960);
xor UO_315 (O_315,N_2970,N_2991);
nand UO_316 (O_316,N_2959,N_2958);
or UO_317 (O_317,N_2946,N_2969);
nand UO_318 (O_318,N_2934,N_2959);
or UO_319 (O_319,N_2940,N_2974);
nor UO_320 (O_320,N_2960,N_2996);
xor UO_321 (O_321,N_2975,N_2960);
nor UO_322 (O_322,N_2962,N_2991);
nand UO_323 (O_323,N_2980,N_2926);
nand UO_324 (O_324,N_2954,N_2929);
or UO_325 (O_325,N_2966,N_2970);
nor UO_326 (O_326,N_2928,N_2955);
nand UO_327 (O_327,N_2990,N_2936);
or UO_328 (O_328,N_2976,N_2990);
nand UO_329 (O_329,N_2950,N_2938);
xor UO_330 (O_330,N_2959,N_2957);
xnor UO_331 (O_331,N_2976,N_2931);
or UO_332 (O_332,N_2972,N_2995);
and UO_333 (O_333,N_2950,N_2925);
nor UO_334 (O_334,N_2953,N_2954);
nor UO_335 (O_335,N_2944,N_2955);
nor UO_336 (O_336,N_2971,N_2949);
or UO_337 (O_337,N_2931,N_2964);
or UO_338 (O_338,N_2925,N_2976);
and UO_339 (O_339,N_2982,N_2942);
nor UO_340 (O_340,N_2926,N_2972);
nor UO_341 (O_341,N_2983,N_2969);
and UO_342 (O_342,N_2975,N_2999);
and UO_343 (O_343,N_2992,N_2982);
and UO_344 (O_344,N_2958,N_2995);
nor UO_345 (O_345,N_2983,N_2925);
xnor UO_346 (O_346,N_2966,N_2976);
nor UO_347 (O_347,N_2997,N_2999);
xnor UO_348 (O_348,N_2936,N_2957);
and UO_349 (O_349,N_2925,N_2965);
or UO_350 (O_350,N_2976,N_2992);
xnor UO_351 (O_351,N_2927,N_2936);
nor UO_352 (O_352,N_2980,N_2961);
or UO_353 (O_353,N_2947,N_2946);
xor UO_354 (O_354,N_2988,N_2952);
xnor UO_355 (O_355,N_2938,N_2940);
and UO_356 (O_356,N_2995,N_2977);
and UO_357 (O_357,N_2940,N_2981);
and UO_358 (O_358,N_2957,N_2993);
or UO_359 (O_359,N_2929,N_2994);
or UO_360 (O_360,N_2982,N_2974);
and UO_361 (O_361,N_2946,N_2979);
or UO_362 (O_362,N_2939,N_2998);
xnor UO_363 (O_363,N_2961,N_2978);
nand UO_364 (O_364,N_2981,N_2980);
nand UO_365 (O_365,N_2938,N_2948);
nand UO_366 (O_366,N_2980,N_2962);
or UO_367 (O_367,N_2930,N_2926);
and UO_368 (O_368,N_2994,N_2938);
or UO_369 (O_369,N_2943,N_2979);
and UO_370 (O_370,N_2962,N_2954);
and UO_371 (O_371,N_2962,N_2959);
nand UO_372 (O_372,N_2991,N_2936);
nand UO_373 (O_373,N_2985,N_2929);
nor UO_374 (O_374,N_2931,N_2993);
nand UO_375 (O_375,N_2935,N_2952);
nand UO_376 (O_376,N_2979,N_2977);
nand UO_377 (O_377,N_2953,N_2943);
or UO_378 (O_378,N_2929,N_2951);
nor UO_379 (O_379,N_2925,N_2994);
nor UO_380 (O_380,N_2946,N_2964);
or UO_381 (O_381,N_2996,N_2926);
and UO_382 (O_382,N_2997,N_2949);
and UO_383 (O_383,N_2929,N_2938);
nor UO_384 (O_384,N_2982,N_2931);
nand UO_385 (O_385,N_2932,N_2930);
or UO_386 (O_386,N_2941,N_2945);
nand UO_387 (O_387,N_2997,N_2935);
nand UO_388 (O_388,N_2984,N_2957);
and UO_389 (O_389,N_2973,N_2932);
or UO_390 (O_390,N_2960,N_2925);
or UO_391 (O_391,N_2945,N_2999);
and UO_392 (O_392,N_2935,N_2933);
or UO_393 (O_393,N_2982,N_2977);
nor UO_394 (O_394,N_2993,N_2995);
and UO_395 (O_395,N_2951,N_2980);
xnor UO_396 (O_396,N_2991,N_2929);
nor UO_397 (O_397,N_2933,N_2977);
xor UO_398 (O_398,N_2969,N_2970);
xnor UO_399 (O_399,N_2950,N_2972);
nor UO_400 (O_400,N_2991,N_2992);
and UO_401 (O_401,N_2981,N_2934);
nand UO_402 (O_402,N_2937,N_2997);
nand UO_403 (O_403,N_2950,N_2984);
or UO_404 (O_404,N_2938,N_2973);
nor UO_405 (O_405,N_2961,N_2969);
and UO_406 (O_406,N_2953,N_2964);
nand UO_407 (O_407,N_2983,N_2947);
or UO_408 (O_408,N_2948,N_2988);
and UO_409 (O_409,N_2958,N_2960);
and UO_410 (O_410,N_2977,N_2929);
nand UO_411 (O_411,N_2985,N_2947);
nand UO_412 (O_412,N_2936,N_2951);
and UO_413 (O_413,N_2964,N_2928);
and UO_414 (O_414,N_2998,N_2985);
and UO_415 (O_415,N_2928,N_2971);
xor UO_416 (O_416,N_2961,N_2957);
nor UO_417 (O_417,N_2949,N_2947);
xor UO_418 (O_418,N_2934,N_2939);
or UO_419 (O_419,N_2948,N_2952);
and UO_420 (O_420,N_2976,N_2984);
nand UO_421 (O_421,N_2994,N_2941);
or UO_422 (O_422,N_2958,N_2989);
nor UO_423 (O_423,N_2989,N_2973);
nand UO_424 (O_424,N_2967,N_2984);
and UO_425 (O_425,N_2993,N_2997);
nor UO_426 (O_426,N_2933,N_2996);
nor UO_427 (O_427,N_2985,N_2943);
and UO_428 (O_428,N_2999,N_2950);
and UO_429 (O_429,N_2934,N_2968);
nor UO_430 (O_430,N_2947,N_2991);
or UO_431 (O_431,N_2979,N_2951);
and UO_432 (O_432,N_2966,N_2991);
and UO_433 (O_433,N_2951,N_2986);
nor UO_434 (O_434,N_2952,N_2997);
xor UO_435 (O_435,N_2985,N_2975);
nor UO_436 (O_436,N_2948,N_2986);
nand UO_437 (O_437,N_2963,N_2976);
nor UO_438 (O_438,N_2980,N_2958);
nand UO_439 (O_439,N_2966,N_2999);
or UO_440 (O_440,N_2998,N_2933);
nor UO_441 (O_441,N_2942,N_2998);
nor UO_442 (O_442,N_2949,N_2993);
nand UO_443 (O_443,N_2958,N_2933);
nor UO_444 (O_444,N_2978,N_2979);
xor UO_445 (O_445,N_2952,N_2974);
nor UO_446 (O_446,N_2934,N_2956);
nand UO_447 (O_447,N_2994,N_2946);
or UO_448 (O_448,N_2947,N_2965);
nand UO_449 (O_449,N_2938,N_2987);
nor UO_450 (O_450,N_2997,N_2990);
xor UO_451 (O_451,N_2946,N_2982);
or UO_452 (O_452,N_2977,N_2934);
nand UO_453 (O_453,N_2987,N_2946);
and UO_454 (O_454,N_2935,N_2932);
nand UO_455 (O_455,N_2986,N_2946);
and UO_456 (O_456,N_2981,N_2958);
nand UO_457 (O_457,N_2989,N_2972);
xor UO_458 (O_458,N_2931,N_2954);
nor UO_459 (O_459,N_2929,N_2967);
nand UO_460 (O_460,N_2997,N_2968);
nor UO_461 (O_461,N_2935,N_2986);
and UO_462 (O_462,N_2992,N_2926);
or UO_463 (O_463,N_2965,N_2929);
nor UO_464 (O_464,N_2944,N_2936);
and UO_465 (O_465,N_2971,N_2977);
xnor UO_466 (O_466,N_2994,N_2956);
nor UO_467 (O_467,N_2937,N_2979);
and UO_468 (O_468,N_2968,N_2959);
nand UO_469 (O_469,N_2948,N_2989);
and UO_470 (O_470,N_2970,N_2958);
nand UO_471 (O_471,N_2961,N_2929);
nor UO_472 (O_472,N_2927,N_2951);
nand UO_473 (O_473,N_2932,N_2997);
and UO_474 (O_474,N_2996,N_2936);
or UO_475 (O_475,N_2936,N_2953);
nand UO_476 (O_476,N_2988,N_2946);
nand UO_477 (O_477,N_2944,N_2965);
nor UO_478 (O_478,N_2941,N_2951);
xnor UO_479 (O_479,N_2957,N_2930);
or UO_480 (O_480,N_2987,N_2934);
nor UO_481 (O_481,N_2980,N_2938);
nand UO_482 (O_482,N_2956,N_2955);
nor UO_483 (O_483,N_2938,N_2993);
xnor UO_484 (O_484,N_2942,N_2991);
nand UO_485 (O_485,N_2999,N_2934);
and UO_486 (O_486,N_2972,N_2976);
nor UO_487 (O_487,N_2959,N_2977);
nor UO_488 (O_488,N_2961,N_2946);
and UO_489 (O_489,N_2978,N_2932);
and UO_490 (O_490,N_2929,N_2939);
nor UO_491 (O_491,N_2993,N_2940);
and UO_492 (O_492,N_2955,N_2994);
xor UO_493 (O_493,N_2963,N_2968);
nand UO_494 (O_494,N_2945,N_2925);
or UO_495 (O_495,N_2999,N_2936);
or UO_496 (O_496,N_2977,N_2944);
and UO_497 (O_497,N_2994,N_2954);
or UO_498 (O_498,N_2949,N_2950);
or UO_499 (O_499,N_2982,N_2978);
endmodule