module basic_1000_10000_1500_2_levels_1xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5005,N_5006,N_5007,N_5008,N_5010,N_5012,N_5014,N_5016,N_5017,N_5019,N_5020,N_5022,N_5023,N_5024,N_5026,N_5027,N_5028,N_5033,N_5036,N_5038,N_5040,N_5041,N_5045,N_5046,N_5048,N_5050,N_5051,N_5052,N_5053,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5066,N_5067,N_5068,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5082,N_5086,N_5087,N_5090,N_5091,N_5092,N_5093,N_5096,N_5097,N_5099,N_5100,N_5102,N_5103,N_5105,N_5106,N_5107,N_5109,N_5110,N_5112,N_5114,N_5115,N_5116,N_5117,N_5118,N_5120,N_5121,N_5123,N_5125,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5135,N_5137,N_5138,N_5139,N_5141,N_5142,N_5145,N_5146,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5158,N_5160,N_5161,N_5162,N_5164,N_5165,N_5166,N_5167,N_5169,N_5171,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5181,N_5182,N_5183,N_5184,N_5185,N_5188,N_5189,N_5190,N_5191,N_5196,N_5198,N_5200,N_5202,N_5205,N_5206,N_5209,N_5211,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5221,N_5224,N_5226,N_5228,N_5233,N_5234,N_5237,N_5238,N_5241,N_5242,N_5243,N_5244,N_5246,N_5247,N_5249,N_5251,N_5252,N_5253,N_5254,N_5256,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5278,N_5279,N_5280,N_5283,N_5286,N_5287,N_5288,N_5291,N_5294,N_5295,N_5296,N_5298,N_5299,N_5300,N_5301,N_5302,N_5305,N_5307,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5318,N_5319,N_5323,N_5324,N_5328,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5338,N_5339,N_5340,N_5344,N_5347,N_5348,N_5349,N_5355,N_5357,N_5358,N_5359,N_5360,N_5362,N_5363,N_5366,N_5369,N_5370,N_5371,N_5373,N_5374,N_5375,N_5377,N_5379,N_5380,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5391,N_5394,N_5395,N_5396,N_5397,N_5399,N_5401,N_5402,N_5403,N_5404,N_5407,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5417,N_5420,N_5423,N_5424,N_5425,N_5433,N_5434,N_5436,N_5438,N_5440,N_5441,N_5444,N_5447,N_5449,N_5450,N_5452,N_5453,N_5457,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5466,N_5468,N_5469,N_5470,N_5471,N_5474,N_5475,N_5476,N_5477,N_5478,N_5484,N_5486,N_5487,N_5489,N_5492,N_5494,N_5495,N_5497,N_5499,N_5501,N_5503,N_5505,N_5507,N_5508,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5519,N_5520,N_5521,N_5522,N_5523,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5534,N_5535,N_5536,N_5537,N_5539,N_5540,N_5541,N_5543,N_5549,N_5550,N_5551,N_5553,N_5558,N_5560,N_5562,N_5564,N_5569,N_5570,N_5571,N_5572,N_5574,N_5575,N_5577,N_5578,N_5580,N_5581,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5595,N_5596,N_5597,N_5599,N_5600,N_5601,N_5603,N_5604,N_5605,N_5607,N_5608,N_5609,N_5612,N_5613,N_5616,N_5617,N_5618,N_5619,N_5620,N_5622,N_5623,N_5625,N_5628,N_5629,N_5630,N_5632,N_5633,N_5634,N_5636,N_5637,N_5642,N_5643,N_5646,N_5647,N_5650,N_5653,N_5654,N_5657,N_5658,N_5664,N_5665,N_5669,N_5673,N_5675,N_5676,N_5678,N_5680,N_5685,N_5686,N_5687,N_5688,N_5689,N_5691,N_5693,N_5694,N_5697,N_5698,N_5699,N_5702,N_5704,N_5706,N_5707,N_5709,N_5712,N_5713,N_5715,N_5716,N_5718,N_5721,N_5722,N_5725,N_5726,N_5728,N_5729,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5745,N_5746,N_5748,N_5749,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5759,N_5760,N_5761,N_5762,N_5763,N_5765,N_5766,N_5767,N_5768,N_5770,N_5771,N_5772,N_5773,N_5777,N_5778,N_5779,N_5780,N_5782,N_5784,N_5785,N_5788,N_5789,N_5790,N_5791,N_5792,N_5794,N_5795,N_5796,N_5798,N_5800,N_5802,N_5803,N_5806,N_5807,N_5808,N_5815,N_5820,N_5821,N_5822,N_5823,N_5824,N_5827,N_5828,N_5829,N_5830,N_5831,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5841,N_5843,N_5844,N_5845,N_5849,N_5850,N_5853,N_5856,N_5857,N_5858,N_5859,N_5860,N_5862,N_5863,N_5865,N_5866,N_5867,N_5868,N_5871,N_5872,N_5873,N_5876,N_5877,N_5878,N_5879,N_5880,N_5882,N_5883,N_5884,N_5885,N_5887,N_5888,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5923,N_5925,N_5926,N_5927,N_5928,N_5930,N_5931,N_5933,N_5934,N_5935,N_5938,N_5941,N_5942,N_5945,N_5946,N_5947,N_5949,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5959,N_5961,N_5964,N_5965,N_5967,N_5970,N_5971,N_5972,N_5974,N_5975,N_5977,N_5978,N_5979,N_5980,N_5982,N_5983,N_5985,N_5986,N_5989,N_5990,N_5992,N_5993,N_5994,N_5995,N_5997,N_6000,N_6004,N_6007,N_6009,N_6010,N_6014,N_6016,N_6018,N_6019,N_6020,N_6022,N_6024,N_6025,N_6027,N_6028,N_6029,N_6031,N_6033,N_6035,N_6036,N_6039,N_6040,N_6042,N_6045,N_6046,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6057,N_6058,N_6059,N_6062,N_6065,N_6067,N_6068,N_6069,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6086,N_6088,N_6089,N_6090,N_6091,N_6094,N_6095,N_6096,N_6098,N_6100,N_6101,N_6103,N_6105,N_6106,N_6107,N_6108,N_6113,N_6117,N_6118,N_6119,N_6122,N_6123,N_6124,N_6125,N_6126,N_6128,N_6130,N_6131,N_6133,N_6136,N_6137,N_6138,N_6139,N_6140,N_6142,N_6144,N_6150,N_6151,N_6154,N_6155,N_6156,N_6157,N_6160,N_6161,N_6163,N_6164,N_6165,N_6166,N_6167,N_6169,N_6170,N_6172,N_6173,N_6174,N_6176,N_6177,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6190,N_6192,N_6193,N_6195,N_6197,N_6199,N_6201,N_6202,N_6203,N_6204,N_6205,N_6208,N_6209,N_6210,N_6212,N_6213,N_6215,N_6218,N_6219,N_6222,N_6223,N_6224,N_6227,N_6230,N_6231,N_6232,N_6234,N_6235,N_6237,N_6239,N_6241,N_6242,N_6245,N_6246,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6264,N_6265,N_6268,N_6272,N_6274,N_6275,N_6278,N_6280,N_6282,N_6284,N_6288,N_6289,N_6292,N_6293,N_6295,N_6296,N_6299,N_6300,N_6302,N_6303,N_6306,N_6309,N_6312,N_6313,N_6314,N_6315,N_6317,N_6319,N_6323,N_6324,N_6325,N_6326,N_6329,N_6331,N_6332,N_6333,N_6334,N_6337,N_6338,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6348,N_6350,N_6351,N_6352,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6362,N_6364,N_6365,N_6369,N_6370,N_6371,N_6373,N_6374,N_6375,N_6376,N_6377,N_6379,N_6380,N_6381,N_6382,N_6387,N_6390,N_6391,N_6392,N_6395,N_6396,N_6397,N_6400,N_6402,N_6403,N_6404,N_6410,N_6411,N_6412,N_6413,N_6415,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6425,N_6427,N_6430,N_6431,N_6432,N_6434,N_6435,N_6437,N_6438,N_6439,N_6441,N_6443,N_6444,N_6446,N_6448,N_6450,N_6451,N_6455,N_6456,N_6459,N_6460,N_6462,N_6463,N_6464,N_6467,N_6468,N_6469,N_6471,N_6472,N_6473,N_6474,N_6475,N_6477,N_6478,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6491,N_6492,N_6493,N_6495,N_6497,N_6499,N_6500,N_6501,N_6503,N_6504,N_6506,N_6507,N_6508,N_6512,N_6514,N_6515,N_6516,N_6517,N_6520,N_6523,N_6524,N_6525,N_6526,N_6528,N_6529,N_6530,N_6532,N_6537,N_6539,N_6541,N_6542,N_6543,N_6545,N_6549,N_6550,N_6552,N_6554,N_6555,N_6556,N_6559,N_6560,N_6561,N_6562,N_6565,N_6567,N_6572,N_6576,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6587,N_6588,N_6591,N_6593,N_6598,N_6602,N_6603,N_6604,N_6606,N_6607,N_6608,N_6610,N_6611,N_6612,N_6615,N_6617,N_6619,N_6620,N_6624,N_6625,N_6626,N_6628,N_6629,N_6631,N_6633,N_6634,N_6636,N_6637,N_6638,N_6643,N_6644,N_6645,N_6647,N_6648,N_6650,N_6651,N_6654,N_6655,N_6656,N_6658,N_6660,N_6662,N_6665,N_6667,N_6668,N_6669,N_6672,N_6673,N_6674,N_6675,N_6678,N_6680,N_6683,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6700,N_6702,N_6703,N_6705,N_6706,N_6708,N_6709,N_6712,N_6713,N_6716,N_6718,N_6720,N_6723,N_6724,N_6725,N_6726,N_6727,N_6729,N_6730,N_6731,N_6732,N_6736,N_6738,N_6739,N_6740,N_6742,N_6746,N_6747,N_6748,N_6752,N_6755,N_6757,N_6758,N_6759,N_6761,N_6762,N_6765,N_6766,N_6767,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6787,N_6788,N_6789,N_6793,N_6795,N_6797,N_6799,N_6800,N_6801,N_6802,N_6803,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6814,N_6815,N_6817,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6827,N_6828,N_6831,N_6835,N_6836,N_6837,N_6839,N_6841,N_6842,N_6844,N_6848,N_6849,N_6850,N_6852,N_6854,N_6855,N_6856,N_6857,N_6859,N_6860,N_6861,N_6865,N_6866,N_6868,N_6869,N_6870,N_6872,N_6874,N_6876,N_6877,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6887,N_6888,N_6889,N_6891,N_6892,N_6893,N_6894,N_6895,N_6897,N_6898,N_6901,N_6902,N_6903,N_6905,N_6906,N_6907,N_6909,N_6911,N_6912,N_6913,N_6914,N_6915,N_6917,N_6918,N_6920,N_6923,N_6924,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6933,N_6934,N_6935,N_6936,N_6938,N_6939,N_6940,N_6943,N_6947,N_6948,N_6949,N_6952,N_6955,N_6956,N_6958,N_6959,N_6960,N_6963,N_6964,N_6965,N_6968,N_6969,N_6970,N_6973,N_6978,N_6979,N_6980,N_6982,N_6983,N_6985,N_6987,N_6989,N_6993,N_6996,N_6998,N_6999,N_7000,N_7001,N_7002,N_7004,N_7005,N_7006,N_7010,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7024,N_7025,N_7026,N_7030,N_7032,N_7034,N_7036,N_7038,N_7044,N_7045,N_7047,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7067,N_7070,N_7072,N_7075,N_7076,N_7078,N_7079,N_7080,N_7082,N_7083,N_7086,N_7088,N_7089,N_7090,N_7091,N_7093,N_7094,N_7096,N_7098,N_7103,N_7105,N_7106,N_7108,N_7109,N_7110,N_7111,N_7112,N_7117,N_7121,N_7122,N_7126,N_7127,N_7128,N_7130,N_7137,N_7138,N_7139,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7150,N_7155,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7165,N_7166,N_7169,N_7170,N_7172,N_7174,N_7175,N_7177,N_7179,N_7180,N_7182,N_7183,N_7185,N_7186,N_7187,N_7188,N_7189,N_7193,N_7194,N_7196,N_7197,N_7198,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7207,N_7209,N_7210,N_7212,N_7213,N_7214,N_7216,N_7218,N_7219,N_7220,N_7221,N_7222,N_7224,N_7227,N_7228,N_7229,N_7232,N_7234,N_7236,N_7238,N_7239,N_7240,N_7242,N_7244,N_7245,N_7248,N_7249,N_7250,N_7252,N_7253,N_7254,N_7258,N_7260,N_7263,N_7264,N_7269,N_7271,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7281,N_7282,N_7283,N_7284,N_7286,N_7287,N_7288,N_7290,N_7291,N_7292,N_7294,N_7295,N_7297,N_7298,N_7300,N_7301,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7313,N_7314,N_7315,N_7316,N_7317,N_7319,N_7320,N_7323,N_7325,N_7326,N_7327,N_7328,N_7329,N_7331,N_7332,N_7334,N_7338,N_7341,N_7343,N_7346,N_7347,N_7348,N_7349,N_7351,N_7352,N_7356,N_7357,N_7360,N_7361,N_7363,N_7365,N_7366,N_7369,N_7370,N_7371,N_7373,N_7375,N_7376,N_7377,N_7379,N_7381,N_7382,N_7383,N_7384,N_7385,N_7390,N_7391,N_7392,N_7393,N_7394,N_7397,N_7399,N_7401,N_7402,N_7404,N_7406,N_7407,N_7408,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7417,N_7418,N_7419,N_7420,N_7421,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7431,N_7432,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7445,N_7446,N_7447,N_7450,N_7452,N_7453,N_7455,N_7456,N_7457,N_7459,N_7460,N_7461,N_7462,N_7463,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7472,N_7475,N_7476,N_7480,N_7482,N_7487,N_7488,N_7489,N_7491,N_7493,N_7494,N_7495,N_7496,N_7498,N_7499,N_7500,N_7502,N_7506,N_7507,N_7508,N_7509,N_7511,N_7512,N_7514,N_7515,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7526,N_7527,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7541,N_7544,N_7545,N_7549,N_7550,N_7551,N_7552,N_7555,N_7557,N_7558,N_7559,N_7560,N_7564,N_7567,N_7568,N_7569,N_7571,N_7573,N_7575,N_7578,N_7579,N_7580,N_7581,N_7582,N_7584,N_7585,N_7589,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7598,N_7599,N_7600,N_7602,N_7605,N_7607,N_7610,N_7611,N_7613,N_7614,N_7616,N_7617,N_7618,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7631,N_7633,N_7637,N_7639,N_7640,N_7642,N_7644,N_7645,N_7646,N_7647,N_7649,N_7650,N_7651,N_7652,N_7654,N_7655,N_7656,N_7657,N_7659,N_7661,N_7662,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7671,N_7672,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7687,N_7689,N_7690,N_7692,N_7693,N_7694,N_7695,N_7697,N_7698,N_7699,N_7700,N_7702,N_7706,N_7707,N_7708,N_7709,N_7711,N_7713,N_7716,N_7720,N_7722,N_7723,N_7724,N_7725,N_7730,N_7733,N_7734,N_7737,N_7739,N_7742,N_7743,N_7744,N_7745,N_7748,N_7749,N_7750,N_7751,N_7752,N_7754,N_7755,N_7758,N_7759,N_7762,N_7763,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7777,N_7778,N_7779,N_7780,N_7782,N_7785,N_7791,N_7795,N_7797,N_7800,N_7801,N_7804,N_7805,N_7806,N_7808,N_7809,N_7812,N_7813,N_7814,N_7815,N_7816,N_7818,N_7820,N_7821,N_7825,N_7826,N_7828,N_7829,N_7832,N_7835,N_7836,N_7838,N_7840,N_7842,N_7844,N_7846,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7856,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7868,N_7869,N_7870,N_7873,N_7874,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7897,N_7899,N_7900,N_7903,N_7904,N_7909,N_7910,N_7911,N_7914,N_7919,N_7921,N_7924,N_7927,N_7928,N_7931,N_7932,N_7933,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7946,N_7947,N_7950,N_7951,N_7952,N_7953,N_7954,N_7956,N_7961,N_7963,N_7964,N_7966,N_7969,N_7970,N_7972,N_7974,N_7975,N_7977,N_7978,N_7979,N_7980,N_7982,N_7984,N_7985,N_7988,N_7989,N_7992,N_7993,N_7994,N_7995,N_7996,N_8000,N_8001,N_8005,N_8010,N_8011,N_8012,N_8013,N_8015,N_8017,N_8019,N_8021,N_8023,N_8024,N_8025,N_8027,N_8028,N_8029,N_8031,N_8032,N_8033,N_8034,N_8035,N_8037,N_8038,N_8039,N_8040,N_8041,N_8043,N_8044,N_8045,N_8048,N_8050,N_8054,N_8055,N_8056,N_8057,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8069,N_8070,N_8071,N_8072,N_8074,N_8075,N_8076,N_8077,N_8079,N_8083,N_8084,N_8086,N_8089,N_8091,N_8092,N_8095,N_8099,N_8100,N_8101,N_8102,N_8104,N_8105,N_8106,N_8107,N_8109,N_8110,N_8113,N_8115,N_8118,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8132,N_8136,N_8140,N_8142,N_8144,N_8145,N_8146,N_8147,N_8150,N_8157,N_8158,N_8161,N_8165,N_8167,N_8168,N_8170,N_8171,N_8177,N_8178,N_8180,N_8181,N_8182,N_8184,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8196,N_8197,N_8200,N_8201,N_8205,N_8206,N_8207,N_8208,N_8212,N_8218,N_8219,N_8220,N_8224,N_8226,N_8228,N_8229,N_8230,N_8231,N_8233,N_8234,N_8235,N_8236,N_8238,N_8239,N_8242,N_8244,N_8246,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8258,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8272,N_8273,N_8274,N_8275,N_8278,N_8279,N_8281,N_8283,N_8286,N_8287,N_8289,N_8293,N_8295,N_8297,N_8298,N_8300,N_8302,N_8303,N_8304,N_8305,N_8308,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8318,N_8320,N_8321,N_8324,N_8325,N_8326,N_8327,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8337,N_8340,N_8341,N_8342,N_8345,N_8346,N_8347,N_8349,N_8350,N_8351,N_8355,N_8357,N_8359,N_8360,N_8361,N_8364,N_8366,N_8367,N_8368,N_8370,N_8372,N_8373,N_8374,N_8375,N_8376,N_8378,N_8379,N_8380,N_8382,N_8383,N_8384,N_8385,N_8387,N_8391,N_8392,N_8393,N_8395,N_8400,N_8401,N_8402,N_8404,N_8406,N_8410,N_8415,N_8417,N_8418,N_8419,N_8420,N_8421,N_8424,N_8426,N_8427,N_8428,N_8429,N_8431,N_8433,N_8434,N_8436,N_8439,N_8440,N_8442,N_8443,N_8444,N_8446,N_8447,N_8448,N_8449,N_8450,N_8453,N_8455,N_8456,N_8457,N_8459,N_8460,N_8465,N_8466,N_8468,N_8470,N_8471,N_8472,N_8474,N_8475,N_8478,N_8480,N_8483,N_8486,N_8487,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8497,N_8499,N_8501,N_8503,N_8504,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8513,N_8515,N_8517,N_8518,N_8520,N_8522,N_8523,N_8525,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8535,N_8536,N_8539,N_8540,N_8541,N_8542,N_8543,N_8546,N_8548,N_8550,N_8552,N_8553,N_8557,N_8558,N_8560,N_8562,N_8563,N_8564,N_8565,N_8566,N_8569,N_8570,N_8571,N_8575,N_8577,N_8578,N_8582,N_8584,N_8585,N_8587,N_8588,N_8591,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8602,N_8603,N_8605,N_8606,N_8607,N_8610,N_8613,N_8614,N_8615,N_8616,N_8618,N_8620,N_8621,N_8622,N_8625,N_8626,N_8629,N_8633,N_8634,N_8637,N_8638,N_8639,N_8642,N_8643,N_8644,N_8646,N_8652,N_8657,N_8658,N_8659,N_8661,N_8662,N_8663,N_8665,N_8668,N_8670,N_8676,N_8677,N_8679,N_8680,N_8685,N_8686,N_8690,N_8691,N_8692,N_8694,N_8695,N_8696,N_8699,N_8700,N_8701,N_8702,N_8704,N_8706,N_8707,N_8708,N_8711,N_8713,N_8714,N_8715,N_8716,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8725,N_8726,N_8727,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8739,N_8740,N_8743,N_8744,N_8745,N_8746,N_8748,N_8749,N_8750,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8759,N_8761,N_8766,N_8767,N_8768,N_8771,N_8773,N_8774,N_8775,N_8777,N_8778,N_8780,N_8782,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8792,N_8793,N_8795,N_8796,N_8797,N_8798,N_8799,N_8801,N_8803,N_8805,N_8807,N_8808,N_8809,N_8812,N_8814,N_8815,N_8816,N_8818,N_8819,N_8820,N_8822,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8842,N_8844,N_8845,N_8847,N_8849,N_8852,N_8854,N_8855,N_8857,N_8860,N_8861,N_8862,N_8864,N_8867,N_8869,N_8871,N_8872,N_8873,N_8875,N_8876,N_8878,N_8879,N_8880,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8890,N_8892,N_8893,N_8895,N_8896,N_8898,N_8899,N_8900,N_8903,N_8904,N_8905,N_8907,N_8913,N_8917,N_8919,N_8920,N_8921,N_8923,N_8924,N_8926,N_8927,N_8932,N_8933,N_8934,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8946,N_8948,N_8950,N_8951,N_8952,N_8953,N_8954,N_8956,N_8959,N_8961,N_8962,N_8963,N_8964,N_8965,N_8967,N_8968,N_8970,N_8971,N_8972,N_8974,N_8975,N_8982,N_8983,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8993,N_8996,N_8999,N_9000,N_9003,N_9005,N_9007,N_9008,N_9010,N_9011,N_9012,N_9013,N_9015,N_9016,N_9017,N_9018,N_9019,N_9023,N_9024,N_9027,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9037,N_9038,N_9039,N_9041,N_9042,N_9045,N_9046,N_9048,N_9049,N_9051,N_9053,N_9055,N_9056,N_9057,N_9061,N_9063,N_9064,N_9067,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9078,N_9079,N_9080,N_9082,N_9085,N_9086,N_9087,N_9088,N_9090,N_9091,N_9095,N_9096,N_9097,N_9099,N_9100,N_9101,N_9103,N_9104,N_9106,N_9113,N_9116,N_9118,N_9119,N_9121,N_9123,N_9125,N_9126,N_9131,N_9134,N_9136,N_9137,N_9138,N_9141,N_9145,N_9147,N_9148,N_9150,N_9152,N_9153,N_9154,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9167,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9179,N_9181,N_9182,N_9183,N_9190,N_9191,N_9192,N_9200,N_9201,N_9202,N_9203,N_9204,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9215,N_9216,N_9217,N_9219,N_9220,N_9221,N_9223,N_9226,N_9229,N_9233,N_9237,N_9240,N_9241,N_9242,N_9243,N_9244,N_9246,N_9247,N_9248,N_9251,N_9252,N_9255,N_9256,N_9257,N_9258,N_9259,N_9262,N_9263,N_9264,N_9266,N_9267,N_9270,N_9271,N_9273,N_9274,N_9275,N_9277,N_9278,N_9282,N_9283,N_9284,N_9285,N_9289,N_9291,N_9292,N_9293,N_9294,N_9295,N_9297,N_9299,N_9300,N_9301,N_9304,N_9305,N_9307,N_9311,N_9314,N_9317,N_9318,N_9320,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9332,N_9333,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9343,N_9345,N_9346,N_9347,N_9348,N_9349,N_9351,N_9352,N_9354,N_9356,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9365,N_9370,N_9373,N_9376,N_9377,N_9378,N_9379,N_9382,N_9384,N_9386,N_9389,N_9393,N_9394,N_9396,N_9397,N_9399,N_9400,N_9401,N_9403,N_9407,N_9408,N_9409,N_9411,N_9412,N_9414,N_9416,N_9418,N_9419,N_9420,N_9422,N_9426,N_9427,N_9429,N_9433,N_9434,N_9436,N_9437,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9449,N_9451,N_9453,N_9454,N_9455,N_9457,N_9458,N_9460,N_9464,N_9468,N_9470,N_9471,N_9473,N_9475,N_9476,N_9477,N_9481,N_9482,N_9484,N_9487,N_9488,N_9489,N_9492,N_9494,N_9495,N_9496,N_9498,N_9500,N_9505,N_9507,N_9508,N_9511,N_9513,N_9515,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9529,N_9531,N_9533,N_9534,N_9536,N_9538,N_9540,N_9542,N_9545,N_9546,N_9547,N_9548,N_9551,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9563,N_9564,N_9566,N_9574,N_9575,N_9577,N_9585,N_9587,N_9589,N_9590,N_9591,N_9592,N_9596,N_9597,N_9599,N_9600,N_9601,N_9602,N_9605,N_9606,N_9607,N_9608,N_9610,N_9611,N_9613,N_9614,N_9617,N_9619,N_9620,N_9622,N_9626,N_9630,N_9633,N_9634,N_9636,N_9637,N_9640,N_9641,N_9644,N_9645,N_9646,N_9648,N_9650,N_9651,N_9652,N_9653,N_9654,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9663,N_9665,N_9667,N_9669,N_9670,N_9671,N_9672,N_9674,N_9675,N_9678,N_9679,N_9681,N_9682,N_9684,N_9686,N_9687,N_9688,N_9689,N_9691,N_9693,N_9696,N_9699,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9709,N_9711,N_9714,N_9715,N_9716,N_9717,N_9719,N_9720,N_9721,N_9724,N_9726,N_9727,N_9728,N_9729,N_9731,N_9732,N_9733,N_9737,N_9738,N_9740,N_9741,N_9742,N_9743,N_9744,N_9746,N_9748,N_9749,N_9750,N_9752,N_9754,N_9755,N_9756,N_9757,N_9759,N_9760,N_9763,N_9764,N_9766,N_9767,N_9769,N_9771,N_9772,N_9774,N_9775,N_9780,N_9781,N_9784,N_9786,N_9787,N_9788,N_9790,N_9791,N_9793,N_9795,N_9799,N_9801,N_9802,N_9803,N_9805,N_9806,N_9808,N_9809,N_9811,N_9815,N_9816,N_9820,N_9821,N_9823,N_9824,N_9825,N_9826,N_9828,N_9830,N_9834,N_9835,N_9837,N_9839,N_9840,N_9843,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9853,N_9854,N_9856,N_9857,N_9858,N_9859,N_9861,N_9862,N_9866,N_9871,N_9872,N_9874,N_9875,N_9877,N_9879,N_9881,N_9882,N_9883,N_9884,N_9885,N_9887,N_9888,N_9891,N_9892,N_9894,N_9896,N_9897,N_9900,N_9902,N_9903,N_9904,N_9905,N_9907,N_9908,N_9909,N_9910,N_9912,N_9914,N_9915,N_9919,N_9920,N_9921,N_9923,N_9924,N_9926,N_9934,N_9936,N_9937,N_9938,N_9941,N_9942,N_9943,N_9947,N_9948,N_9949,N_9951,N_9954,N_9955,N_9956,N_9958,N_9960,N_9962,N_9963,N_9965,N_9967,N_9968,N_9969,N_9971,N_9973,N_9974,N_9975,N_9980,N_9981,N_9983,N_9984,N_9986,N_9988,N_9989,N_9993,N_9994,N_9995,N_9997,N_9998,N_9999;
nand U0 (N_0,In_84,In_945);
nand U1 (N_1,In_972,In_97);
nor U2 (N_2,In_474,In_538);
nand U3 (N_3,In_378,In_556);
and U4 (N_4,In_449,In_848);
nand U5 (N_5,In_776,In_9);
nor U6 (N_6,In_570,In_852);
nor U7 (N_7,In_319,In_559);
nor U8 (N_8,In_668,In_112);
nor U9 (N_9,In_147,In_929);
and U10 (N_10,In_573,In_358);
and U11 (N_11,In_694,In_66);
and U12 (N_12,In_989,In_237);
nand U13 (N_13,In_823,In_145);
xor U14 (N_14,In_949,In_311);
or U15 (N_15,In_462,In_824);
nand U16 (N_16,In_234,In_334);
and U17 (N_17,In_325,In_755);
and U18 (N_18,In_995,In_246);
or U19 (N_19,In_298,In_816);
nand U20 (N_20,In_15,In_545);
nor U21 (N_21,In_220,In_692);
nand U22 (N_22,In_11,In_415);
nand U23 (N_23,In_154,In_239);
nor U24 (N_24,In_531,In_447);
and U25 (N_25,In_833,In_926);
nor U26 (N_26,In_895,In_568);
nor U27 (N_27,In_354,In_437);
or U28 (N_28,In_377,In_452);
and U29 (N_29,In_927,In_445);
and U30 (N_30,In_539,In_606);
nor U31 (N_31,In_134,In_240);
and U32 (N_32,In_603,In_365);
nor U33 (N_33,In_841,In_718);
nand U34 (N_34,In_160,In_654);
nand U35 (N_35,In_301,In_83);
and U36 (N_36,In_574,In_255);
and U37 (N_37,In_673,In_578);
or U38 (N_38,In_385,In_674);
nor U39 (N_39,In_269,In_389);
nand U40 (N_40,In_260,In_631);
and U41 (N_41,In_830,In_772);
nand U42 (N_42,In_355,In_178);
or U43 (N_43,In_528,In_324);
nand U44 (N_44,In_189,In_297);
and U45 (N_45,In_300,In_106);
nand U46 (N_46,In_595,In_643);
nor U47 (N_47,In_78,In_119);
or U48 (N_48,In_778,In_894);
nor U49 (N_49,In_33,In_655);
and U50 (N_50,In_96,In_359);
or U51 (N_51,In_457,In_962);
or U52 (N_52,In_318,In_39);
or U53 (N_53,In_336,In_278);
nor U54 (N_54,In_493,In_803);
and U55 (N_55,In_863,In_888);
nand U56 (N_56,In_215,In_524);
nor U57 (N_57,In_845,In_715);
nor U58 (N_58,In_337,In_525);
and U59 (N_59,In_828,In_520);
nand U60 (N_60,In_4,In_717);
and U61 (N_61,In_843,In_596);
nand U62 (N_62,In_304,In_503);
nor U63 (N_63,In_34,In_180);
or U64 (N_64,In_988,In_339);
or U65 (N_65,In_347,In_549);
nand U66 (N_66,In_594,In_345);
or U67 (N_67,In_497,In_948);
nand U68 (N_68,In_349,In_176);
nand U69 (N_69,In_31,In_342);
or U70 (N_70,In_273,In_241);
or U71 (N_71,In_969,In_840);
nand U72 (N_72,In_601,In_79);
nand U73 (N_73,In_95,In_814);
nand U74 (N_74,In_68,In_174);
nand U75 (N_75,In_263,In_314);
and U76 (N_76,In_646,In_495);
nand U77 (N_77,In_741,In_566);
nor U78 (N_78,In_22,In_496);
nand U79 (N_79,In_290,In_481);
and U80 (N_80,In_7,In_429);
nor U81 (N_81,In_282,In_466);
or U82 (N_82,In_941,In_121);
nor U83 (N_83,In_92,In_544);
and U84 (N_84,In_744,In_45);
nand U85 (N_85,In_515,In_100);
or U86 (N_86,In_430,In_720);
or U87 (N_87,In_913,In_5);
nand U88 (N_88,In_422,In_821);
or U89 (N_89,In_861,In_396);
or U90 (N_90,In_149,In_785);
nand U91 (N_91,In_144,In_126);
nand U92 (N_92,In_442,In_25);
and U93 (N_93,In_899,In_439);
nand U94 (N_94,In_40,In_581);
and U95 (N_95,In_571,In_771);
and U96 (N_96,In_48,In_478);
nand U97 (N_97,In_148,In_903);
and U98 (N_98,In_799,In_839);
nand U99 (N_99,In_155,In_883);
and U100 (N_100,In_118,In_219);
or U101 (N_101,In_761,In_217);
and U102 (N_102,In_151,In_680);
nor U103 (N_103,In_187,In_666);
and U104 (N_104,In_804,In_548);
nand U105 (N_105,In_185,In_338);
or U106 (N_106,In_536,In_871);
nor U107 (N_107,In_380,In_383);
xor U108 (N_108,In_274,In_953);
nor U109 (N_109,In_994,In_341);
nor U110 (N_110,In_504,In_990);
nand U111 (N_111,In_87,In_213);
nand U112 (N_112,In_955,In_438);
nand U113 (N_113,In_878,In_560);
nor U114 (N_114,In_296,In_82);
nand U115 (N_115,In_238,In_707);
nand U116 (N_116,In_85,In_133);
and U117 (N_117,In_822,In_272);
and U118 (N_118,In_956,In_867);
and U119 (N_119,In_487,In_513);
and U120 (N_120,In_172,In_932);
or U121 (N_121,In_259,In_173);
or U122 (N_122,In_223,In_880);
and U123 (N_123,In_882,In_944);
nand U124 (N_124,In_617,In_854);
and U125 (N_125,In_41,In_558);
or U126 (N_126,In_609,In_829);
nand U127 (N_127,In_411,In_851);
nor U128 (N_128,In_242,In_786);
nand U129 (N_129,In_689,In_51);
nand U130 (N_130,In_508,In_862);
and U131 (N_131,In_636,In_838);
nor U132 (N_132,In_472,In_564);
or U133 (N_133,In_16,In_930);
nand U134 (N_134,In_293,In_390);
or U135 (N_135,In_317,In_908);
nand U136 (N_136,In_143,In_781);
nand U137 (N_137,In_904,In_977);
nor U138 (N_138,In_991,In_491);
and U139 (N_139,In_868,In_262);
nor U140 (N_140,In_625,In_887);
nor U141 (N_141,In_473,In_667);
or U142 (N_142,In_653,In_323);
nor U143 (N_143,In_167,In_922);
nand U144 (N_144,In_12,In_89);
or U145 (N_145,In_244,In_470);
or U146 (N_146,In_612,In_837);
and U147 (N_147,In_295,In_902);
and U148 (N_148,In_866,In_328);
and U149 (N_149,In_211,In_691);
nand U150 (N_150,In_150,In_376);
nand U151 (N_151,In_494,In_233);
nand U152 (N_152,In_471,In_791);
nor U153 (N_153,In_970,In_627);
and U154 (N_154,In_825,In_693);
or U155 (N_155,In_102,In_251);
nand U156 (N_156,In_918,In_875);
nand U157 (N_157,In_884,In_869);
and U158 (N_158,In_381,In_555);
and U159 (N_159,In_76,In_623);
nand U160 (N_160,In_469,In_247);
and U161 (N_161,In_113,In_737);
nor U162 (N_162,In_114,In_14);
nor U163 (N_163,In_626,In_767);
nor U164 (N_164,In_727,In_811);
nand U165 (N_165,In_346,In_593);
nor U166 (N_166,In_157,In_322);
or U167 (N_167,In_435,In_639);
or U168 (N_168,In_577,In_710);
nor U169 (N_169,In_634,In_218);
nand U170 (N_170,In_881,In_175);
nand U171 (N_171,In_128,In_672);
nor U172 (N_172,In_896,In_584);
xnor U173 (N_173,In_931,In_373);
or U174 (N_174,In_794,In_936);
or U175 (N_175,In_400,In_254);
and U176 (N_176,In_892,In_420);
and U177 (N_177,In_924,In_879);
and U178 (N_178,In_588,In_256);
or U179 (N_179,In_946,In_446);
nand U180 (N_180,In_0,In_543);
nor U181 (N_181,In_214,In_393);
and U182 (N_182,In_731,In_410);
and U183 (N_183,In_414,In_876);
nand U184 (N_184,In_897,In_512);
nand U185 (N_185,In_698,In_532);
or U186 (N_186,In_98,In_912);
and U187 (N_187,In_61,In_925);
or U188 (N_188,In_893,In_850);
or U189 (N_189,In_739,In_464);
nor U190 (N_190,In_764,In_159);
nand U191 (N_191,In_796,In_94);
nand U192 (N_192,In_57,In_960);
and U193 (N_193,In_367,In_281);
nor U194 (N_194,In_788,In_708);
nor U195 (N_195,In_586,In_834);
nor U196 (N_196,In_171,In_770);
or U197 (N_197,In_99,In_505);
nor U198 (N_198,In_424,In_137);
and U199 (N_199,In_406,In_726);
nand U200 (N_200,In_245,In_756);
nand U201 (N_201,In_937,In_745);
nand U202 (N_202,In_227,In_773);
or U203 (N_203,In_206,In_333);
and U204 (N_204,In_506,In_455);
nor U205 (N_205,In_279,In_250);
and U206 (N_206,In_704,In_135);
nand U207 (N_207,In_21,In_20);
nor U208 (N_208,In_987,In_886);
nand U209 (N_209,In_43,In_484);
or U210 (N_210,In_52,In_343);
nand U211 (N_211,In_729,In_364);
nor U212 (N_212,In_50,In_93);
nand U213 (N_213,In_614,In_64);
nand U214 (N_214,In_321,In_961);
or U215 (N_215,In_140,In_73);
nand U216 (N_216,In_266,In_249);
nor U217 (N_217,In_243,In_448);
or U218 (N_218,In_62,In_404);
nand U219 (N_219,In_540,In_855);
nor U220 (N_220,In_71,In_600);
nand U221 (N_221,In_635,In_648);
or U222 (N_222,In_535,In_44);
and U223 (N_223,In_479,In_332);
and U224 (N_224,In_3,In_401);
nand U225 (N_225,In_394,In_194);
or U226 (N_226,In_817,In_374);
or U227 (N_227,In_10,In_65);
nand U228 (N_228,In_488,In_562);
or U229 (N_229,In_230,In_928);
nor U230 (N_230,In_748,In_939);
or U231 (N_231,In_652,In_477);
and U232 (N_232,In_379,In_292);
nand U233 (N_233,In_943,In_919);
and U234 (N_234,In_517,In_516);
nor U235 (N_235,In_69,In_565);
and U236 (N_236,In_117,In_976);
and U237 (N_237,In_552,In_664);
nand U238 (N_238,In_108,In_774);
nand U239 (N_239,In_712,In_819);
nand U240 (N_240,In_60,In_277);
nor U241 (N_241,In_368,In_307);
and U242 (N_242,In_610,In_547);
or U243 (N_243,In_320,In_350);
nand U244 (N_244,In_541,In_709);
nor U245 (N_245,In_125,In_847);
nor U246 (N_246,In_416,In_752);
nand U247 (N_247,In_436,In_724);
nor U248 (N_248,In_658,In_690);
nor U249 (N_249,In_361,In_619);
or U250 (N_250,In_360,In_502);
nor U251 (N_251,In_585,In_344);
or U252 (N_252,In_465,In_6);
nor U253 (N_253,In_809,In_910);
nor U254 (N_254,In_980,In_787);
or U255 (N_255,In_763,In_179);
and U256 (N_256,In_158,In_742);
nand U257 (N_257,In_280,In_370);
nand U258 (N_258,In_975,In_957);
or U259 (N_259,In_901,In_681);
or U260 (N_260,In_63,In_426);
nor U261 (N_261,In_226,In_909);
and U262 (N_262,In_856,In_705);
and U263 (N_263,In_561,In_35);
nor U264 (N_264,In_192,In_808);
and U265 (N_265,In_865,In_202);
and U266 (N_266,In_229,In_801);
nand U267 (N_267,In_372,In_917);
or U268 (N_268,In_188,In_940);
and U269 (N_269,In_993,In_701);
and U270 (N_270,In_141,In_58);
or U271 (N_271,In_56,In_369);
and U272 (N_272,In_23,In_486);
nor U273 (N_273,In_417,In_914);
or U274 (N_274,In_19,In_730);
or U275 (N_275,In_934,In_419);
nand U276 (N_276,In_184,In_340);
nor U277 (N_277,In_751,In_782);
and U278 (N_278,In_951,In_890);
nand U279 (N_279,In_310,In_511);
or U280 (N_280,In_569,In_699);
and U281 (N_281,In_270,In_792);
nor U282 (N_282,In_362,In_706);
or U283 (N_283,In_713,In_978);
nor U284 (N_284,In_399,In_327);
or U285 (N_285,In_659,In_152);
nand U286 (N_286,In_711,In_997);
nor U287 (N_287,In_753,In_971);
and U288 (N_288,In_663,In_754);
and U289 (N_289,In_29,In_351);
and U290 (N_290,In_575,In_526);
or U291 (N_291,In_425,In_567);
nand U292 (N_292,In_597,In_453);
nor U293 (N_293,In_225,In_162);
nand U294 (N_294,In_81,In_74);
nor U295 (N_295,In_507,In_32);
nand U296 (N_296,In_331,In_170);
nor U297 (N_297,In_13,In_521);
or U298 (N_298,In_427,In_732);
or U299 (N_299,In_758,In_454);
and U300 (N_300,In_966,In_352);
and U301 (N_301,In_210,In_458);
or U302 (N_302,In_54,In_687);
nor U303 (N_303,In_762,In_252);
nor U304 (N_304,In_235,In_716);
or U305 (N_305,In_580,In_412);
nor U306 (N_306,In_264,In_67);
nor U307 (N_307,In_17,In_428);
or U308 (N_308,In_200,In_388);
nand U309 (N_309,In_703,In_783);
and U310 (N_310,In_620,In_657);
nor U311 (N_311,In_498,In_222);
nand U312 (N_312,In_421,In_330);
nand U313 (N_313,In_733,In_534);
nand U314 (N_314,In_193,In_678);
or U315 (N_315,In_90,In_797);
nand U316 (N_316,In_27,In_221);
nand U317 (N_317,In_434,In_490);
nand U318 (N_318,In_363,In_191);
xnor U319 (N_319,In_992,In_183);
nor U320 (N_320,In_846,In_463);
and U321 (N_321,In_450,In_387);
nand U322 (N_322,In_366,In_467);
and U323 (N_323,In_554,In_2);
and U324 (N_324,In_408,In_967);
nand U325 (N_325,In_844,In_641);
nand U326 (N_326,In_759,In_287);
and U327 (N_327,In_650,In_138);
nor U328 (N_328,In_697,In_725);
and U329 (N_329,In_813,In_459);
nor U330 (N_330,In_873,In_405);
nand U331 (N_331,In_798,In_38);
nand U332 (N_332,In_624,In_315);
or U333 (N_333,In_679,In_999);
nor U334 (N_334,In_736,In_375);
nand U335 (N_335,In_810,In_289);
nand U336 (N_336,In_199,In_529);
nand U337 (N_337,In_700,In_642);
nand U338 (N_338,In_204,In_224);
and U339 (N_339,In_265,In_291);
nor U340 (N_340,In_858,In_647);
nor U341 (N_341,In_728,In_431);
or U342 (N_342,In_616,In_587);
nand U343 (N_343,In_166,In_686);
nand U344 (N_344,In_661,In_283);
or U345 (N_345,In_77,In_615);
nor U346 (N_346,In_982,In_18);
nor U347 (N_347,In_468,In_36);
and U348 (N_348,In_286,In_831);
nor U349 (N_349,In_815,In_527);
nand U350 (N_350,In_719,In_142);
or U351 (N_351,In_303,In_483);
nand U352 (N_352,In_312,In_127);
nor U353 (N_353,In_308,In_632);
nor U354 (N_354,In_313,In_201);
and U355 (N_355,In_860,In_986);
and U356 (N_356,In_432,In_985);
nand U357 (N_357,In_738,In_386);
nor U358 (N_358,In_104,In_285);
nand U359 (N_359,In_42,In_80);
and U360 (N_360,In_485,In_637);
nor U361 (N_361,In_766,In_443);
or U362 (N_362,In_231,In_123);
nand U363 (N_363,In_784,In_605);
nand U364 (N_364,In_807,In_476);
nor U365 (N_365,In_973,In_870);
nand U366 (N_366,In_115,In_670);
and U367 (N_367,In_981,In_397);
nand U368 (N_368,In_276,In_169);
nor U369 (N_369,In_906,In_460);
or U370 (N_370,In_523,In_550);
nor U371 (N_371,In_177,In_46);
nor U372 (N_372,In_806,In_30);
nand U373 (N_373,In_91,In_853);
nor U374 (N_374,In_129,In_618);
and U375 (N_375,In_409,In_916);
nand U376 (N_376,In_676,In_433);
and U377 (N_377,In_599,In_563);
nor U378 (N_378,In_644,In_907);
nand U379 (N_379,In_489,In_677);
nor U380 (N_380,In_132,In_195);
and U381 (N_381,In_827,In_403);
or U382 (N_382,In_248,In_820);
nor U383 (N_383,In_284,In_418);
and U384 (N_384,In_271,In_398);
or U385 (N_385,In_933,In_258);
and U386 (N_386,In_24,In_921);
nand U387 (N_387,In_722,In_391);
or U388 (N_388,In_335,In_288);
nor U389 (N_389,In_530,In_186);
nor U390 (N_390,In_1,In_604);
nor U391 (N_391,In_103,In_518);
or U392 (N_392,In_836,In_207);
and U393 (N_393,In_522,In_702);
nor U394 (N_394,In_947,In_53);
nand U395 (N_395,In_979,In_26);
and U396 (N_396,In_818,In_105);
nor U397 (N_397,In_675,In_793);
nor U398 (N_398,In_628,In_629);
or U399 (N_399,In_898,In_613);
or U400 (N_400,In_757,In_805);
nand U401 (N_401,In_402,In_557);
or U402 (N_402,In_357,In_735);
nor U403 (N_403,In_590,In_576);
or U404 (N_404,In_130,In_261);
and U405 (N_405,In_622,In_316);
nor U406 (N_406,In_958,In_746);
xnor U407 (N_407,In_382,In_168);
and U408 (N_408,In_826,In_857);
nand U409 (N_409,In_645,In_671);
or U410 (N_410,In_542,In_116);
nand U411 (N_411,In_329,In_920);
and U412 (N_412,In_197,In_768);
nor U413 (N_413,In_591,In_302);
and U414 (N_414,In_911,In_533);
nand U415 (N_415,In_163,In_800);
nor U416 (N_416,In_8,In_682);
or U417 (N_417,In_440,In_146);
nor U418 (N_418,In_514,In_519);
nand U419 (N_419,In_208,In_500);
and U420 (N_420,In_734,In_165);
nand U421 (N_421,In_553,In_294);
and U422 (N_422,In_461,In_630);
nor U423 (N_423,In_499,In_968);
and U424 (N_424,In_684,In_37);
and U425 (N_425,In_608,In_164);
nor U426 (N_426,In_110,In_651);
nand U427 (N_427,In_326,In_216);
or U428 (N_428,In_750,In_72);
and U429 (N_429,In_475,In_501);
or U430 (N_430,In_423,In_779);
and U431 (N_431,In_203,In_583);
nor U432 (N_432,In_905,In_28);
nor U433 (N_433,In_482,In_510);
or U434 (N_434,In_965,In_181);
or U435 (N_435,In_228,In_392);
nor U436 (N_436,In_665,In_638);
nor U437 (N_437,In_891,In_353);
or U438 (N_438,In_662,In_696);
nand U439 (N_439,In_572,In_835);
or U440 (N_440,In_49,In_685);
and U441 (N_441,In_75,In_959);
nand U442 (N_442,In_236,In_582);
nand U443 (N_443,In_107,In_743);
or U444 (N_444,In_942,In_441);
nor U445 (N_445,In_356,In_182);
nand U446 (N_446,In_607,In_889);
and U447 (N_447,In_88,In_780);
nor U448 (N_448,In_589,In_790);
xnor U449 (N_449,In_885,In_395);
nor U450 (N_450,In_101,In_198);
nor U451 (N_451,In_915,In_305);
and U452 (N_452,In_640,In_714);
and U453 (N_453,In_111,In_598);
nand U454 (N_454,In_156,In_740);
and U455 (N_455,In_984,In_384);
nor U456 (N_456,In_695,In_348);
nor U457 (N_457,In_938,In_232);
nor U458 (N_458,In_900,In_688);
or U459 (N_459,In_832,In_775);
nor U460 (N_460,In_974,In_509);
and U461 (N_461,In_546,In_592);
and U462 (N_462,In_795,In_212);
or U463 (N_463,In_723,In_749);
nor U464 (N_464,In_964,In_849);
or U465 (N_465,In_131,In_492);
nand U466 (N_466,In_196,In_275);
or U467 (N_467,In_602,In_55);
nor U468 (N_468,In_59,In_954);
and U469 (N_469,In_309,In_70);
or U470 (N_470,In_413,In_996);
nor U471 (N_471,In_769,In_649);
or U472 (N_472,In_86,In_579);
xnor U473 (N_473,In_923,In_299);
nor U474 (N_474,In_683,In_874);
and U475 (N_475,In_864,In_877);
nand U476 (N_476,In_537,In_407);
nor U477 (N_477,In_253,In_306);
nor U478 (N_478,In_480,In_812);
and U479 (N_479,In_998,In_139);
nand U480 (N_480,In_136,In_444);
and U481 (N_481,In_952,In_721);
nand U482 (N_482,In_656,In_747);
nand U483 (N_483,In_669,In_268);
and U484 (N_484,In_161,In_122);
and U485 (N_485,In_109,In_451);
nor U486 (N_486,In_209,In_190);
and U487 (N_487,In_257,In_765);
nor U488 (N_488,In_267,In_802);
or U489 (N_489,In_47,In_789);
nor U490 (N_490,In_777,In_963);
or U491 (N_491,In_872,In_950);
and U492 (N_492,In_551,In_859);
nor U493 (N_493,In_983,In_456);
nand U494 (N_494,In_660,In_611);
nand U495 (N_495,In_124,In_760);
nor U496 (N_496,In_205,In_120);
and U497 (N_497,In_633,In_935);
nor U498 (N_498,In_621,In_842);
nor U499 (N_499,In_153,In_371);
or U500 (N_500,In_756,In_1);
nor U501 (N_501,In_283,In_592);
nand U502 (N_502,In_407,In_96);
nor U503 (N_503,In_943,In_66);
nor U504 (N_504,In_548,In_574);
xor U505 (N_505,In_850,In_13);
nand U506 (N_506,In_766,In_920);
nor U507 (N_507,In_377,In_715);
nand U508 (N_508,In_329,In_969);
and U509 (N_509,In_653,In_86);
nor U510 (N_510,In_425,In_558);
and U511 (N_511,In_775,In_740);
or U512 (N_512,In_445,In_629);
nand U513 (N_513,In_147,In_136);
nand U514 (N_514,In_2,In_861);
nor U515 (N_515,In_120,In_556);
nor U516 (N_516,In_216,In_474);
and U517 (N_517,In_847,In_130);
or U518 (N_518,In_397,In_519);
and U519 (N_519,In_295,In_165);
or U520 (N_520,In_298,In_185);
nand U521 (N_521,In_368,In_447);
nand U522 (N_522,In_791,In_23);
nand U523 (N_523,In_334,In_563);
nor U524 (N_524,In_196,In_914);
and U525 (N_525,In_154,In_294);
nor U526 (N_526,In_307,In_241);
nand U527 (N_527,In_665,In_780);
nor U528 (N_528,In_196,In_584);
or U529 (N_529,In_516,In_946);
nor U530 (N_530,In_308,In_240);
and U531 (N_531,In_512,In_149);
nand U532 (N_532,In_784,In_818);
nand U533 (N_533,In_821,In_914);
nand U534 (N_534,In_824,In_832);
and U535 (N_535,In_430,In_54);
nand U536 (N_536,In_712,In_728);
and U537 (N_537,In_439,In_944);
nand U538 (N_538,In_190,In_987);
or U539 (N_539,In_572,In_800);
or U540 (N_540,In_113,In_260);
and U541 (N_541,In_462,In_253);
or U542 (N_542,In_932,In_244);
or U543 (N_543,In_124,In_315);
nor U544 (N_544,In_680,In_491);
and U545 (N_545,In_71,In_228);
nor U546 (N_546,In_870,In_988);
or U547 (N_547,In_84,In_561);
nor U548 (N_548,In_141,In_488);
nand U549 (N_549,In_505,In_529);
and U550 (N_550,In_495,In_754);
and U551 (N_551,In_899,In_332);
nor U552 (N_552,In_822,In_511);
nand U553 (N_553,In_220,In_913);
nand U554 (N_554,In_699,In_285);
and U555 (N_555,In_516,In_613);
nand U556 (N_556,In_631,In_983);
nor U557 (N_557,In_720,In_546);
nand U558 (N_558,In_594,In_284);
and U559 (N_559,In_263,In_462);
and U560 (N_560,In_728,In_350);
nor U561 (N_561,In_82,In_158);
or U562 (N_562,In_646,In_274);
nor U563 (N_563,In_750,In_58);
or U564 (N_564,In_702,In_926);
and U565 (N_565,In_460,In_876);
xor U566 (N_566,In_688,In_680);
or U567 (N_567,In_106,In_965);
or U568 (N_568,In_697,In_397);
nand U569 (N_569,In_341,In_780);
nand U570 (N_570,In_492,In_66);
nor U571 (N_571,In_722,In_984);
nand U572 (N_572,In_431,In_386);
and U573 (N_573,In_493,In_188);
or U574 (N_574,In_354,In_266);
or U575 (N_575,In_666,In_609);
or U576 (N_576,In_816,In_546);
and U577 (N_577,In_333,In_515);
and U578 (N_578,In_244,In_634);
nand U579 (N_579,In_212,In_340);
and U580 (N_580,In_62,In_973);
and U581 (N_581,In_163,In_579);
and U582 (N_582,In_780,In_179);
or U583 (N_583,In_195,In_812);
or U584 (N_584,In_23,In_711);
or U585 (N_585,In_648,In_62);
and U586 (N_586,In_570,In_870);
and U587 (N_587,In_788,In_151);
nor U588 (N_588,In_865,In_58);
nand U589 (N_589,In_441,In_546);
nand U590 (N_590,In_956,In_33);
or U591 (N_591,In_498,In_70);
and U592 (N_592,In_600,In_286);
and U593 (N_593,In_946,In_665);
and U594 (N_594,In_760,In_560);
and U595 (N_595,In_939,In_743);
and U596 (N_596,In_183,In_515);
or U597 (N_597,In_478,In_337);
or U598 (N_598,In_785,In_917);
nor U599 (N_599,In_15,In_241);
and U600 (N_600,In_121,In_278);
or U601 (N_601,In_755,In_31);
nand U602 (N_602,In_833,In_910);
or U603 (N_603,In_147,In_829);
or U604 (N_604,In_76,In_314);
nor U605 (N_605,In_204,In_883);
or U606 (N_606,In_270,In_247);
nor U607 (N_607,In_777,In_84);
nand U608 (N_608,In_410,In_791);
nor U609 (N_609,In_32,In_112);
nand U610 (N_610,In_291,In_53);
or U611 (N_611,In_92,In_459);
nand U612 (N_612,In_322,In_703);
and U613 (N_613,In_857,In_61);
and U614 (N_614,In_746,In_650);
and U615 (N_615,In_818,In_502);
nand U616 (N_616,In_631,In_939);
and U617 (N_617,In_211,In_44);
or U618 (N_618,In_62,In_965);
or U619 (N_619,In_539,In_723);
or U620 (N_620,In_101,In_239);
nor U621 (N_621,In_384,In_820);
and U622 (N_622,In_382,In_623);
nor U623 (N_623,In_242,In_656);
nand U624 (N_624,In_184,In_824);
nand U625 (N_625,In_855,In_492);
nand U626 (N_626,In_170,In_51);
and U627 (N_627,In_563,In_919);
and U628 (N_628,In_621,In_393);
nand U629 (N_629,In_887,In_90);
or U630 (N_630,In_976,In_600);
and U631 (N_631,In_990,In_337);
nand U632 (N_632,In_436,In_953);
nor U633 (N_633,In_936,In_621);
or U634 (N_634,In_247,In_5);
nor U635 (N_635,In_884,In_736);
nand U636 (N_636,In_571,In_432);
or U637 (N_637,In_81,In_182);
or U638 (N_638,In_774,In_526);
nor U639 (N_639,In_405,In_889);
and U640 (N_640,In_744,In_484);
nor U641 (N_641,In_622,In_591);
or U642 (N_642,In_989,In_752);
or U643 (N_643,In_614,In_519);
nand U644 (N_644,In_274,In_475);
or U645 (N_645,In_343,In_528);
or U646 (N_646,In_145,In_868);
nand U647 (N_647,In_562,In_370);
nand U648 (N_648,In_233,In_973);
and U649 (N_649,In_403,In_345);
nand U650 (N_650,In_377,In_193);
and U651 (N_651,In_591,In_107);
nand U652 (N_652,In_305,In_377);
or U653 (N_653,In_35,In_87);
nand U654 (N_654,In_15,In_347);
or U655 (N_655,In_788,In_589);
and U656 (N_656,In_59,In_463);
or U657 (N_657,In_614,In_2);
or U658 (N_658,In_10,In_119);
nor U659 (N_659,In_146,In_840);
nand U660 (N_660,In_894,In_889);
nand U661 (N_661,In_485,In_215);
or U662 (N_662,In_213,In_644);
nor U663 (N_663,In_266,In_72);
or U664 (N_664,In_465,In_20);
or U665 (N_665,In_445,In_229);
or U666 (N_666,In_876,In_834);
nand U667 (N_667,In_993,In_194);
and U668 (N_668,In_213,In_980);
nor U669 (N_669,In_730,In_838);
nand U670 (N_670,In_282,In_223);
nand U671 (N_671,In_748,In_427);
nand U672 (N_672,In_659,In_262);
nand U673 (N_673,In_502,In_826);
or U674 (N_674,In_246,In_284);
nor U675 (N_675,In_76,In_237);
or U676 (N_676,In_765,In_609);
nor U677 (N_677,In_991,In_858);
or U678 (N_678,In_977,In_980);
nor U679 (N_679,In_66,In_6);
or U680 (N_680,In_347,In_429);
nor U681 (N_681,In_952,In_955);
nor U682 (N_682,In_818,In_346);
nand U683 (N_683,In_117,In_374);
nor U684 (N_684,In_353,In_716);
nor U685 (N_685,In_636,In_285);
or U686 (N_686,In_204,In_381);
nand U687 (N_687,In_15,In_267);
and U688 (N_688,In_475,In_783);
and U689 (N_689,In_557,In_782);
nor U690 (N_690,In_801,In_421);
nor U691 (N_691,In_102,In_862);
nand U692 (N_692,In_467,In_505);
and U693 (N_693,In_496,In_233);
and U694 (N_694,In_545,In_703);
nand U695 (N_695,In_161,In_459);
and U696 (N_696,In_945,In_748);
nand U697 (N_697,In_703,In_228);
or U698 (N_698,In_218,In_150);
or U699 (N_699,In_964,In_175);
and U700 (N_700,In_699,In_560);
or U701 (N_701,In_366,In_104);
and U702 (N_702,In_165,In_729);
nor U703 (N_703,In_838,In_575);
nor U704 (N_704,In_469,In_841);
and U705 (N_705,In_899,In_123);
nor U706 (N_706,In_525,In_755);
or U707 (N_707,In_866,In_320);
nor U708 (N_708,In_584,In_788);
nor U709 (N_709,In_423,In_158);
and U710 (N_710,In_561,In_667);
and U711 (N_711,In_531,In_669);
and U712 (N_712,In_268,In_897);
and U713 (N_713,In_321,In_514);
or U714 (N_714,In_129,In_236);
nand U715 (N_715,In_351,In_39);
nor U716 (N_716,In_760,In_480);
nor U717 (N_717,In_641,In_534);
nor U718 (N_718,In_451,In_93);
nor U719 (N_719,In_487,In_818);
and U720 (N_720,In_891,In_154);
nor U721 (N_721,In_357,In_202);
and U722 (N_722,In_371,In_885);
or U723 (N_723,In_535,In_482);
nor U724 (N_724,In_788,In_572);
and U725 (N_725,In_27,In_645);
nand U726 (N_726,In_474,In_947);
nand U727 (N_727,In_487,In_173);
nor U728 (N_728,In_175,In_115);
or U729 (N_729,In_606,In_15);
nor U730 (N_730,In_414,In_124);
and U731 (N_731,In_109,In_680);
or U732 (N_732,In_771,In_598);
nand U733 (N_733,In_685,In_108);
nor U734 (N_734,In_184,In_41);
nand U735 (N_735,In_455,In_222);
and U736 (N_736,In_538,In_850);
nor U737 (N_737,In_966,In_920);
nor U738 (N_738,In_485,In_278);
and U739 (N_739,In_739,In_441);
nand U740 (N_740,In_187,In_64);
nand U741 (N_741,In_570,In_760);
and U742 (N_742,In_865,In_971);
nor U743 (N_743,In_747,In_573);
nor U744 (N_744,In_660,In_438);
and U745 (N_745,In_381,In_369);
and U746 (N_746,In_745,In_742);
xnor U747 (N_747,In_251,In_240);
nand U748 (N_748,In_75,In_343);
xnor U749 (N_749,In_640,In_607);
and U750 (N_750,In_417,In_963);
and U751 (N_751,In_580,In_86);
nand U752 (N_752,In_128,In_750);
and U753 (N_753,In_906,In_723);
or U754 (N_754,In_403,In_628);
nor U755 (N_755,In_452,In_311);
nor U756 (N_756,In_838,In_561);
and U757 (N_757,In_769,In_748);
and U758 (N_758,In_624,In_840);
and U759 (N_759,In_867,In_71);
and U760 (N_760,In_443,In_395);
nand U761 (N_761,In_300,In_72);
nand U762 (N_762,In_915,In_663);
and U763 (N_763,In_188,In_956);
nor U764 (N_764,In_644,In_707);
or U765 (N_765,In_271,In_625);
or U766 (N_766,In_745,In_361);
nor U767 (N_767,In_556,In_663);
nor U768 (N_768,In_449,In_608);
and U769 (N_769,In_140,In_182);
and U770 (N_770,In_100,In_492);
nand U771 (N_771,In_491,In_0);
or U772 (N_772,In_2,In_834);
nand U773 (N_773,In_566,In_55);
or U774 (N_774,In_689,In_264);
nor U775 (N_775,In_335,In_313);
nand U776 (N_776,In_803,In_558);
and U777 (N_777,In_606,In_120);
nand U778 (N_778,In_979,In_684);
nand U779 (N_779,In_124,In_296);
nand U780 (N_780,In_939,In_152);
xnor U781 (N_781,In_528,In_471);
and U782 (N_782,In_44,In_116);
nor U783 (N_783,In_56,In_810);
nand U784 (N_784,In_654,In_313);
or U785 (N_785,In_205,In_637);
and U786 (N_786,In_826,In_765);
nand U787 (N_787,In_322,In_657);
nor U788 (N_788,In_627,In_880);
nand U789 (N_789,In_176,In_703);
xnor U790 (N_790,In_595,In_583);
nand U791 (N_791,In_571,In_986);
or U792 (N_792,In_54,In_514);
nand U793 (N_793,In_659,In_328);
or U794 (N_794,In_319,In_476);
and U795 (N_795,In_208,In_212);
nor U796 (N_796,In_293,In_862);
nor U797 (N_797,In_683,In_169);
or U798 (N_798,In_334,In_800);
nand U799 (N_799,In_227,In_234);
nand U800 (N_800,In_422,In_255);
nand U801 (N_801,In_546,In_345);
nand U802 (N_802,In_309,In_529);
and U803 (N_803,In_576,In_936);
and U804 (N_804,In_719,In_597);
nand U805 (N_805,In_546,In_409);
nand U806 (N_806,In_916,In_773);
nor U807 (N_807,In_732,In_526);
or U808 (N_808,In_599,In_922);
nand U809 (N_809,In_859,In_121);
or U810 (N_810,In_670,In_122);
or U811 (N_811,In_64,In_656);
nand U812 (N_812,In_13,In_185);
and U813 (N_813,In_930,In_541);
or U814 (N_814,In_917,In_170);
nand U815 (N_815,In_812,In_112);
nor U816 (N_816,In_92,In_679);
and U817 (N_817,In_981,In_572);
nor U818 (N_818,In_877,In_648);
nor U819 (N_819,In_992,In_563);
or U820 (N_820,In_267,In_989);
nand U821 (N_821,In_992,In_424);
nand U822 (N_822,In_215,In_67);
and U823 (N_823,In_522,In_157);
nand U824 (N_824,In_208,In_423);
xnor U825 (N_825,In_299,In_871);
xnor U826 (N_826,In_442,In_172);
nand U827 (N_827,In_835,In_630);
nor U828 (N_828,In_755,In_926);
and U829 (N_829,In_114,In_827);
or U830 (N_830,In_306,In_143);
nor U831 (N_831,In_131,In_54);
or U832 (N_832,In_124,In_268);
or U833 (N_833,In_826,In_206);
nor U834 (N_834,In_553,In_44);
and U835 (N_835,In_320,In_582);
or U836 (N_836,In_867,In_548);
and U837 (N_837,In_185,In_164);
nand U838 (N_838,In_1,In_103);
or U839 (N_839,In_267,In_558);
and U840 (N_840,In_187,In_356);
and U841 (N_841,In_206,In_871);
xnor U842 (N_842,In_62,In_860);
and U843 (N_843,In_110,In_188);
or U844 (N_844,In_618,In_524);
nor U845 (N_845,In_675,In_754);
or U846 (N_846,In_172,In_877);
nand U847 (N_847,In_868,In_397);
or U848 (N_848,In_178,In_391);
or U849 (N_849,In_576,In_957);
nand U850 (N_850,In_566,In_743);
nand U851 (N_851,In_540,In_107);
nand U852 (N_852,In_897,In_474);
nand U853 (N_853,In_200,In_837);
and U854 (N_854,In_907,In_300);
or U855 (N_855,In_673,In_148);
nand U856 (N_856,In_331,In_564);
nor U857 (N_857,In_927,In_495);
nor U858 (N_858,In_136,In_762);
nor U859 (N_859,In_425,In_662);
or U860 (N_860,In_844,In_193);
nor U861 (N_861,In_854,In_376);
and U862 (N_862,In_208,In_148);
nor U863 (N_863,In_544,In_890);
or U864 (N_864,In_846,In_440);
or U865 (N_865,In_180,In_266);
nor U866 (N_866,In_654,In_405);
or U867 (N_867,In_533,In_96);
nand U868 (N_868,In_675,In_939);
and U869 (N_869,In_684,In_488);
or U870 (N_870,In_511,In_412);
nand U871 (N_871,In_659,In_476);
or U872 (N_872,In_191,In_373);
and U873 (N_873,In_764,In_542);
xnor U874 (N_874,In_843,In_510);
and U875 (N_875,In_166,In_341);
nor U876 (N_876,In_23,In_121);
or U877 (N_877,In_62,In_635);
nand U878 (N_878,In_17,In_997);
and U879 (N_879,In_488,In_882);
and U880 (N_880,In_865,In_950);
or U881 (N_881,In_618,In_432);
nand U882 (N_882,In_481,In_867);
nand U883 (N_883,In_424,In_372);
nor U884 (N_884,In_408,In_537);
nor U885 (N_885,In_500,In_628);
or U886 (N_886,In_241,In_313);
or U887 (N_887,In_164,In_206);
nor U888 (N_888,In_547,In_360);
nand U889 (N_889,In_970,In_896);
nor U890 (N_890,In_367,In_102);
nor U891 (N_891,In_308,In_143);
nor U892 (N_892,In_962,In_937);
nor U893 (N_893,In_569,In_60);
and U894 (N_894,In_315,In_449);
or U895 (N_895,In_544,In_925);
or U896 (N_896,In_631,In_701);
or U897 (N_897,In_628,In_406);
and U898 (N_898,In_360,In_670);
nor U899 (N_899,In_816,In_101);
nand U900 (N_900,In_258,In_528);
or U901 (N_901,In_255,In_149);
and U902 (N_902,In_300,In_797);
nand U903 (N_903,In_612,In_129);
or U904 (N_904,In_279,In_961);
nand U905 (N_905,In_301,In_113);
nand U906 (N_906,In_493,In_524);
nor U907 (N_907,In_574,In_817);
or U908 (N_908,In_407,In_33);
and U909 (N_909,In_39,In_400);
nor U910 (N_910,In_142,In_433);
nand U911 (N_911,In_311,In_373);
and U912 (N_912,In_748,In_717);
or U913 (N_913,In_22,In_357);
nor U914 (N_914,In_720,In_363);
nor U915 (N_915,In_67,In_615);
nand U916 (N_916,In_963,In_518);
nand U917 (N_917,In_528,In_39);
and U918 (N_918,In_672,In_473);
nand U919 (N_919,In_951,In_334);
and U920 (N_920,In_646,In_720);
nand U921 (N_921,In_716,In_422);
or U922 (N_922,In_925,In_155);
or U923 (N_923,In_111,In_910);
nand U924 (N_924,In_462,In_63);
nand U925 (N_925,In_125,In_151);
or U926 (N_926,In_277,In_367);
or U927 (N_927,In_655,In_627);
or U928 (N_928,In_768,In_669);
or U929 (N_929,In_182,In_382);
nand U930 (N_930,In_460,In_148);
nand U931 (N_931,In_526,In_835);
nor U932 (N_932,In_323,In_190);
nor U933 (N_933,In_818,In_275);
and U934 (N_934,In_363,In_240);
or U935 (N_935,In_781,In_503);
nor U936 (N_936,In_126,In_679);
or U937 (N_937,In_126,In_65);
and U938 (N_938,In_58,In_231);
nand U939 (N_939,In_98,In_123);
nand U940 (N_940,In_931,In_992);
or U941 (N_941,In_274,In_137);
and U942 (N_942,In_915,In_755);
nand U943 (N_943,In_968,In_120);
nor U944 (N_944,In_527,In_48);
and U945 (N_945,In_564,In_100);
or U946 (N_946,In_214,In_946);
and U947 (N_947,In_231,In_69);
or U948 (N_948,In_896,In_290);
and U949 (N_949,In_626,In_292);
and U950 (N_950,In_149,In_769);
and U951 (N_951,In_833,In_790);
nor U952 (N_952,In_356,In_138);
nand U953 (N_953,In_604,In_18);
and U954 (N_954,In_712,In_166);
nor U955 (N_955,In_301,In_286);
nor U956 (N_956,In_106,In_866);
and U957 (N_957,In_987,In_236);
nand U958 (N_958,In_539,In_638);
and U959 (N_959,In_495,In_714);
and U960 (N_960,In_773,In_129);
nor U961 (N_961,In_770,In_689);
and U962 (N_962,In_919,In_202);
xnor U963 (N_963,In_928,In_428);
and U964 (N_964,In_284,In_648);
and U965 (N_965,In_887,In_284);
nand U966 (N_966,In_739,In_669);
nor U967 (N_967,In_733,In_292);
and U968 (N_968,In_539,In_768);
and U969 (N_969,In_69,In_429);
nor U970 (N_970,In_651,In_938);
or U971 (N_971,In_516,In_504);
and U972 (N_972,In_183,In_983);
and U973 (N_973,In_181,In_510);
nor U974 (N_974,In_814,In_654);
and U975 (N_975,In_983,In_755);
nand U976 (N_976,In_572,In_331);
nand U977 (N_977,In_199,In_25);
and U978 (N_978,In_134,In_151);
or U979 (N_979,In_335,In_511);
or U980 (N_980,In_352,In_11);
and U981 (N_981,In_576,In_920);
or U982 (N_982,In_742,In_910);
nor U983 (N_983,In_940,In_764);
or U984 (N_984,In_410,In_135);
and U985 (N_985,In_239,In_342);
nor U986 (N_986,In_130,In_763);
nor U987 (N_987,In_347,In_145);
and U988 (N_988,In_295,In_560);
nor U989 (N_989,In_336,In_558);
nand U990 (N_990,In_536,In_385);
or U991 (N_991,In_304,In_799);
nor U992 (N_992,In_430,In_212);
and U993 (N_993,In_628,In_237);
or U994 (N_994,In_264,In_494);
or U995 (N_995,In_728,In_981);
nor U996 (N_996,In_972,In_295);
or U997 (N_997,In_523,In_239);
nor U998 (N_998,In_784,In_162);
nor U999 (N_999,In_913,In_232);
or U1000 (N_1000,In_533,In_209);
or U1001 (N_1001,In_723,In_886);
nand U1002 (N_1002,In_791,In_617);
nand U1003 (N_1003,In_515,In_878);
nand U1004 (N_1004,In_345,In_109);
nor U1005 (N_1005,In_14,In_182);
and U1006 (N_1006,In_106,In_958);
and U1007 (N_1007,In_757,In_788);
nand U1008 (N_1008,In_495,In_847);
nor U1009 (N_1009,In_968,In_467);
and U1010 (N_1010,In_223,In_294);
or U1011 (N_1011,In_744,In_196);
and U1012 (N_1012,In_447,In_201);
and U1013 (N_1013,In_976,In_34);
and U1014 (N_1014,In_668,In_254);
and U1015 (N_1015,In_834,In_150);
or U1016 (N_1016,In_481,In_771);
and U1017 (N_1017,In_707,In_391);
nor U1018 (N_1018,In_290,In_240);
or U1019 (N_1019,In_622,In_888);
nor U1020 (N_1020,In_38,In_361);
nor U1021 (N_1021,In_987,In_647);
nor U1022 (N_1022,In_320,In_969);
and U1023 (N_1023,In_544,In_708);
and U1024 (N_1024,In_735,In_867);
and U1025 (N_1025,In_45,In_928);
nor U1026 (N_1026,In_370,In_439);
nor U1027 (N_1027,In_194,In_524);
nand U1028 (N_1028,In_718,In_258);
nand U1029 (N_1029,In_905,In_822);
nor U1030 (N_1030,In_632,In_478);
nor U1031 (N_1031,In_825,In_819);
and U1032 (N_1032,In_747,In_701);
or U1033 (N_1033,In_930,In_708);
or U1034 (N_1034,In_411,In_589);
nand U1035 (N_1035,In_482,In_391);
and U1036 (N_1036,In_841,In_637);
or U1037 (N_1037,In_624,In_757);
nor U1038 (N_1038,In_653,In_758);
nor U1039 (N_1039,In_742,In_438);
or U1040 (N_1040,In_870,In_701);
or U1041 (N_1041,In_35,In_14);
nor U1042 (N_1042,In_818,In_290);
or U1043 (N_1043,In_155,In_981);
nand U1044 (N_1044,In_124,In_482);
or U1045 (N_1045,In_640,In_596);
and U1046 (N_1046,In_107,In_86);
and U1047 (N_1047,In_711,In_468);
nand U1048 (N_1048,In_88,In_902);
nor U1049 (N_1049,In_68,In_9);
and U1050 (N_1050,In_8,In_637);
nand U1051 (N_1051,In_882,In_724);
nor U1052 (N_1052,In_255,In_370);
and U1053 (N_1053,In_796,In_129);
nand U1054 (N_1054,In_468,In_295);
or U1055 (N_1055,In_970,In_497);
nor U1056 (N_1056,In_900,In_833);
nand U1057 (N_1057,In_12,In_141);
xnor U1058 (N_1058,In_219,In_530);
and U1059 (N_1059,In_942,In_370);
and U1060 (N_1060,In_799,In_750);
or U1061 (N_1061,In_855,In_455);
and U1062 (N_1062,In_23,In_537);
nand U1063 (N_1063,In_461,In_89);
nand U1064 (N_1064,In_302,In_548);
or U1065 (N_1065,In_492,In_697);
nor U1066 (N_1066,In_93,In_517);
nor U1067 (N_1067,In_484,In_509);
and U1068 (N_1068,In_349,In_400);
and U1069 (N_1069,In_73,In_658);
or U1070 (N_1070,In_613,In_6);
and U1071 (N_1071,In_911,In_496);
and U1072 (N_1072,In_621,In_11);
nand U1073 (N_1073,In_268,In_230);
nand U1074 (N_1074,In_316,In_66);
nand U1075 (N_1075,In_177,In_553);
nor U1076 (N_1076,In_626,In_830);
nor U1077 (N_1077,In_988,In_711);
or U1078 (N_1078,In_598,In_604);
or U1079 (N_1079,In_998,In_761);
or U1080 (N_1080,In_415,In_0);
nand U1081 (N_1081,In_173,In_729);
nand U1082 (N_1082,In_647,In_285);
and U1083 (N_1083,In_73,In_989);
nand U1084 (N_1084,In_110,In_634);
and U1085 (N_1085,In_868,In_628);
or U1086 (N_1086,In_790,In_926);
or U1087 (N_1087,In_762,In_499);
nor U1088 (N_1088,In_854,In_695);
nor U1089 (N_1089,In_209,In_643);
and U1090 (N_1090,In_446,In_831);
and U1091 (N_1091,In_697,In_528);
nor U1092 (N_1092,In_608,In_35);
or U1093 (N_1093,In_679,In_764);
nand U1094 (N_1094,In_814,In_135);
nor U1095 (N_1095,In_118,In_19);
nor U1096 (N_1096,In_785,In_165);
nor U1097 (N_1097,In_986,In_184);
or U1098 (N_1098,In_747,In_160);
and U1099 (N_1099,In_584,In_699);
nand U1100 (N_1100,In_621,In_683);
or U1101 (N_1101,In_388,In_109);
nor U1102 (N_1102,In_430,In_92);
nor U1103 (N_1103,In_885,In_117);
nor U1104 (N_1104,In_194,In_67);
nor U1105 (N_1105,In_595,In_549);
and U1106 (N_1106,In_250,In_742);
nand U1107 (N_1107,In_705,In_187);
or U1108 (N_1108,In_572,In_871);
and U1109 (N_1109,In_224,In_233);
nor U1110 (N_1110,In_12,In_469);
and U1111 (N_1111,In_606,In_946);
or U1112 (N_1112,In_671,In_842);
nor U1113 (N_1113,In_803,In_994);
nand U1114 (N_1114,In_247,In_690);
or U1115 (N_1115,In_232,In_598);
nand U1116 (N_1116,In_786,In_809);
and U1117 (N_1117,In_563,In_866);
and U1118 (N_1118,In_750,In_982);
and U1119 (N_1119,In_788,In_263);
or U1120 (N_1120,In_712,In_257);
or U1121 (N_1121,In_359,In_909);
and U1122 (N_1122,In_747,In_962);
nor U1123 (N_1123,In_186,In_328);
nand U1124 (N_1124,In_312,In_573);
nor U1125 (N_1125,In_498,In_447);
nor U1126 (N_1126,In_764,In_29);
and U1127 (N_1127,In_379,In_334);
nand U1128 (N_1128,In_670,In_169);
or U1129 (N_1129,In_784,In_263);
nand U1130 (N_1130,In_896,In_858);
or U1131 (N_1131,In_195,In_411);
and U1132 (N_1132,In_894,In_311);
or U1133 (N_1133,In_952,In_351);
nor U1134 (N_1134,In_228,In_316);
nor U1135 (N_1135,In_560,In_442);
or U1136 (N_1136,In_558,In_9);
and U1137 (N_1137,In_503,In_992);
and U1138 (N_1138,In_179,In_417);
nor U1139 (N_1139,In_575,In_129);
nand U1140 (N_1140,In_237,In_451);
and U1141 (N_1141,In_804,In_87);
and U1142 (N_1142,In_744,In_283);
or U1143 (N_1143,In_111,In_610);
or U1144 (N_1144,In_656,In_632);
nand U1145 (N_1145,In_220,In_139);
or U1146 (N_1146,In_639,In_434);
nor U1147 (N_1147,In_677,In_493);
nand U1148 (N_1148,In_401,In_152);
or U1149 (N_1149,In_981,In_592);
and U1150 (N_1150,In_236,In_113);
nand U1151 (N_1151,In_638,In_711);
or U1152 (N_1152,In_807,In_753);
nand U1153 (N_1153,In_602,In_486);
and U1154 (N_1154,In_799,In_647);
and U1155 (N_1155,In_286,In_435);
nor U1156 (N_1156,In_488,In_287);
nand U1157 (N_1157,In_511,In_285);
nand U1158 (N_1158,In_508,In_36);
nor U1159 (N_1159,In_296,In_761);
nor U1160 (N_1160,In_673,In_772);
nand U1161 (N_1161,In_213,In_244);
and U1162 (N_1162,In_39,In_885);
or U1163 (N_1163,In_71,In_882);
nor U1164 (N_1164,In_206,In_475);
nor U1165 (N_1165,In_651,In_845);
nor U1166 (N_1166,In_995,In_601);
or U1167 (N_1167,In_853,In_957);
nor U1168 (N_1168,In_388,In_152);
nor U1169 (N_1169,In_763,In_459);
and U1170 (N_1170,In_415,In_814);
nand U1171 (N_1171,In_781,In_886);
nand U1172 (N_1172,In_86,In_862);
and U1173 (N_1173,In_546,In_128);
and U1174 (N_1174,In_345,In_229);
nor U1175 (N_1175,In_396,In_939);
nor U1176 (N_1176,In_194,In_239);
nor U1177 (N_1177,In_492,In_541);
nand U1178 (N_1178,In_753,In_605);
or U1179 (N_1179,In_783,In_42);
and U1180 (N_1180,In_246,In_613);
nor U1181 (N_1181,In_864,In_9);
and U1182 (N_1182,In_359,In_811);
and U1183 (N_1183,In_388,In_383);
nor U1184 (N_1184,In_188,In_590);
xor U1185 (N_1185,In_97,In_228);
nor U1186 (N_1186,In_205,In_79);
and U1187 (N_1187,In_444,In_592);
nand U1188 (N_1188,In_965,In_34);
nand U1189 (N_1189,In_181,In_323);
or U1190 (N_1190,In_150,In_664);
nor U1191 (N_1191,In_513,In_603);
nor U1192 (N_1192,In_475,In_198);
nor U1193 (N_1193,In_25,In_903);
nor U1194 (N_1194,In_502,In_935);
nor U1195 (N_1195,In_445,In_723);
nor U1196 (N_1196,In_707,In_93);
or U1197 (N_1197,In_919,In_183);
or U1198 (N_1198,In_440,In_95);
and U1199 (N_1199,In_782,In_877);
nand U1200 (N_1200,In_178,In_699);
and U1201 (N_1201,In_430,In_132);
or U1202 (N_1202,In_702,In_421);
nand U1203 (N_1203,In_696,In_155);
or U1204 (N_1204,In_158,In_31);
nor U1205 (N_1205,In_544,In_790);
nor U1206 (N_1206,In_939,In_823);
and U1207 (N_1207,In_913,In_60);
nor U1208 (N_1208,In_516,In_819);
or U1209 (N_1209,In_416,In_461);
or U1210 (N_1210,In_445,In_486);
xor U1211 (N_1211,In_633,In_415);
nor U1212 (N_1212,In_789,In_29);
nand U1213 (N_1213,In_20,In_763);
nor U1214 (N_1214,In_781,In_632);
nor U1215 (N_1215,In_54,In_205);
or U1216 (N_1216,In_688,In_58);
and U1217 (N_1217,In_894,In_818);
nand U1218 (N_1218,In_345,In_201);
nor U1219 (N_1219,In_851,In_387);
nand U1220 (N_1220,In_563,In_207);
nor U1221 (N_1221,In_778,In_568);
nand U1222 (N_1222,In_340,In_987);
nand U1223 (N_1223,In_675,In_999);
and U1224 (N_1224,In_814,In_584);
and U1225 (N_1225,In_764,In_164);
and U1226 (N_1226,In_176,In_261);
nor U1227 (N_1227,In_722,In_633);
nor U1228 (N_1228,In_44,In_90);
nand U1229 (N_1229,In_456,In_592);
nor U1230 (N_1230,In_956,In_686);
and U1231 (N_1231,In_967,In_109);
nor U1232 (N_1232,In_458,In_71);
nand U1233 (N_1233,In_198,In_197);
and U1234 (N_1234,In_830,In_259);
and U1235 (N_1235,In_233,In_158);
or U1236 (N_1236,In_53,In_574);
nand U1237 (N_1237,In_582,In_564);
and U1238 (N_1238,In_805,In_783);
nand U1239 (N_1239,In_292,In_295);
and U1240 (N_1240,In_332,In_72);
and U1241 (N_1241,In_466,In_285);
nor U1242 (N_1242,In_516,In_818);
or U1243 (N_1243,In_783,In_104);
and U1244 (N_1244,In_109,In_829);
and U1245 (N_1245,In_35,In_125);
and U1246 (N_1246,In_141,In_482);
or U1247 (N_1247,In_272,In_7);
or U1248 (N_1248,In_766,In_628);
nand U1249 (N_1249,In_740,In_278);
and U1250 (N_1250,In_895,In_202);
nor U1251 (N_1251,In_724,In_614);
nand U1252 (N_1252,In_185,In_552);
nor U1253 (N_1253,In_812,In_166);
and U1254 (N_1254,In_558,In_604);
nor U1255 (N_1255,In_988,In_302);
and U1256 (N_1256,In_956,In_950);
nand U1257 (N_1257,In_28,In_128);
or U1258 (N_1258,In_733,In_171);
and U1259 (N_1259,In_52,In_791);
xor U1260 (N_1260,In_940,In_882);
nand U1261 (N_1261,In_844,In_925);
nor U1262 (N_1262,In_290,In_247);
nand U1263 (N_1263,In_280,In_371);
nand U1264 (N_1264,In_66,In_406);
or U1265 (N_1265,In_858,In_859);
nor U1266 (N_1266,In_521,In_897);
nand U1267 (N_1267,In_460,In_790);
or U1268 (N_1268,In_564,In_435);
nand U1269 (N_1269,In_198,In_738);
or U1270 (N_1270,In_106,In_897);
and U1271 (N_1271,In_935,In_271);
nor U1272 (N_1272,In_181,In_215);
or U1273 (N_1273,In_128,In_403);
nor U1274 (N_1274,In_687,In_899);
nor U1275 (N_1275,In_526,In_654);
nor U1276 (N_1276,In_706,In_631);
or U1277 (N_1277,In_765,In_764);
nor U1278 (N_1278,In_194,In_27);
or U1279 (N_1279,In_702,In_436);
xor U1280 (N_1280,In_341,In_461);
or U1281 (N_1281,In_765,In_67);
or U1282 (N_1282,In_14,In_631);
and U1283 (N_1283,In_417,In_855);
or U1284 (N_1284,In_103,In_396);
nor U1285 (N_1285,In_417,In_309);
nor U1286 (N_1286,In_420,In_774);
nor U1287 (N_1287,In_11,In_811);
nor U1288 (N_1288,In_137,In_395);
nand U1289 (N_1289,In_320,In_71);
nor U1290 (N_1290,In_501,In_507);
nor U1291 (N_1291,In_22,In_291);
or U1292 (N_1292,In_997,In_916);
nand U1293 (N_1293,In_910,In_568);
or U1294 (N_1294,In_358,In_389);
nand U1295 (N_1295,In_82,In_521);
or U1296 (N_1296,In_469,In_724);
and U1297 (N_1297,In_990,In_94);
or U1298 (N_1298,In_707,In_898);
nand U1299 (N_1299,In_168,In_909);
nor U1300 (N_1300,In_581,In_9);
nand U1301 (N_1301,In_775,In_100);
and U1302 (N_1302,In_368,In_208);
nor U1303 (N_1303,In_463,In_718);
nor U1304 (N_1304,In_398,In_512);
nand U1305 (N_1305,In_636,In_705);
and U1306 (N_1306,In_56,In_709);
and U1307 (N_1307,In_557,In_623);
and U1308 (N_1308,In_726,In_441);
and U1309 (N_1309,In_182,In_939);
and U1310 (N_1310,In_577,In_248);
and U1311 (N_1311,In_134,In_677);
nand U1312 (N_1312,In_202,In_84);
or U1313 (N_1313,In_406,In_603);
or U1314 (N_1314,In_623,In_72);
nor U1315 (N_1315,In_902,In_998);
nand U1316 (N_1316,In_364,In_842);
and U1317 (N_1317,In_713,In_106);
and U1318 (N_1318,In_770,In_323);
and U1319 (N_1319,In_47,In_233);
and U1320 (N_1320,In_648,In_464);
or U1321 (N_1321,In_801,In_867);
nor U1322 (N_1322,In_656,In_772);
nand U1323 (N_1323,In_104,In_817);
or U1324 (N_1324,In_402,In_197);
and U1325 (N_1325,In_968,In_182);
nor U1326 (N_1326,In_36,In_733);
nand U1327 (N_1327,In_752,In_460);
or U1328 (N_1328,In_814,In_511);
or U1329 (N_1329,In_837,In_949);
nor U1330 (N_1330,In_229,In_278);
nor U1331 (N_1331,In_168,In_436);
nor U1332 (N_1332,In_625,In_805);
or U1333 (N_1333,In_591,In_483);
nor U1334 (N_1334,In_966,In_629);
nor U1335 (N_1335,In_334,In_53);
xor U1336 (N_1336,In_235,In_525);
nand U1337 (N_1337,In_179,In_721);
and U1338 (N_1338,In_207,In_519);
nor U1339 (N_1339,In_30,In_675);
and U1340 (N_1340,In_251,In_906);
nor U1341 (N_1341,In_679,In_457);
nor U1342 (N_1342,In_523,In_584);
or U1343 (N_1343,In_575,In_715);
and U1344 (N_1344,In_718,In_757);
and U1345 (N_1345,In_213,In_272);
and U1346 (N_1346,In_515,In_563);
or U1347 (N_1347,In_950,In_703);
and U1348 (N_1348,In_546,In_306);
or U1349 (N_1349,In_281,In_701);
nor U1350 (N_1350,In_78,In_976);
and U1351 (N_1351,In_938,In_446);
or U1352 (N_1352,In_289,In_385);
nor U1353 (N_1353,In_454,In_34);
or U1354 (N_1354,In_140,In_716);
and U1355 (N_1355,In_815,In_925);
nor U1356 (N_1356,In_402,In_644);
nand U1357 (N_1357,In_935,In_48);
or U1358 (N_1358,In_873,In_813);
nor U1359 (N_1359,In_630,In_285);
and U1360 (N_1360,In_903,In_571);
nor U1361 (N_1361,In_328,In_435);
nor U1362 (N_1362,In_314,In_723);
and U1363 (N_1363,In_803,In_735);
xnor U1364 (N_1364,In_185,In_273);
nand U1365 (N_1365,In_355,In_967);
nor U1366 (N_1366,In_282,In_32);
nor U1367 (N_1367,In_243,In_764);
nand U1368 (N_1368,In_119,In_584);
or U1369 (N_1369,In_834,In_9);
and U1370 (N_1370,In_448,In_407);
nand U1371 (N_1371,In_896,In_976);
nor U1372 (N_1372,In_66,In_922);
nor U1373 (N_1373,In_828,In_580);
or U1374 (N_1374,In_411,In_866);
and U1375 (N_1375,In_812,In_957);
and U1376 (N_1376,In_480,In_913);
nand U1377 (N_1377,In_283,In_10);
nor U1378 (N_1378,In_943,In_916);
or U1379 (N_1379,In_457,In_34);
or U1380 (N_1380,In_533,In_169);
nor U1381 (N_1381,In_142,In_837);
nand U1382 (N_1382,In_420,In_788);
nand U1383 (N_1383,In_875,In_574);
and U1384 (N_1384,In_978,In_504);
or U1385 (N_1385,In_110,In_285);
nor U1386 (N_1386,In_309,In_500);
and U1387 (N_1387,In_196,In_560);
nand U1388 (N_1388,In_701,In_585);
and U1389 (N_1389,In_881,In_216);
nand U1390 (N_1390,In_651,In_658);
and U1391 (N_1391,In_272,In_495);
nor U1392 (N_1392,In_231,In_155);
nand U1393 (N_1393,In_728,In_165);
or U1394 (N_1394,In_122,In_469);
nor U1395 (N_1395,In_718,In_552);
nor U1396 (N_1396,In_672,In_377);
xnor U1397 (N_1397,In_364,In_341);
and U1398 (N_1398,In_507,In_731);
nor U1399 (N_1399,In_241,In_796);
or U1400 (N_1400,In_744,In_645);
nor U1401 (N_1401,In_561,In_488);
and U1402 (N_1402,In_324,In_50);
nand U1403 (N_1403,In_238,In_325);
nand U1404 (N_1404,In_500,In_359);
or U1405 (N_1405,In_992,In_61);
nor U1406 (N_1406,In_435,In_512);
or U1407 (N_1407,In_127,In_769);
nand U1408 (N_1408,In_165,In_199);
nand U1409 (N_1409,In_217,In_840);
or U1410 (N_1410,In_739,In_939);
and U1411 (N_1411,In_611,In_599);
and U1412 (N_1412,In_33,In_186);
or U1413 (N_1413,In_135,In_753);
nor U1414 (N_1414,In_944,In_522);
nor U1415 (N_1415,In_853,In_513);
nor U1416 (N_1416,In_354,In_232);
nor U1417 (N_1417,In_77,In_73);
or U1418 (N_1418,In_56,In_603);
or U1419 (N_1419,In_858,In_522);
nor U1420 (N_1420,In_292,In_973);
nor U1421 (N_1421,In_956,In_83);
and U1422 (N_1422,In_51,In_902);
nor U1423 (N_1423,In_450,In_743);
xnor U1424 (N_1424,In_667,In_538);
and U1425 (N_1425,In_626,In_625);
nor U1426 (N_1426,In_818,In_511);
or U1427 (N_1427,In_619,In_683);
nand U1428 (N_1428,In_218,In_125);
and U1429 (N_1429,In_564,In_905);
and U1430 (N_1430,In_487,In_360);
nand U1431 (N_1431,In_345,In_996);
or U1432 (N_1432,In_142,In_171);
and U1433 (N_1433,In_636,In_861);
or U1434 (N_1434,In_482,In_587);
nand U1435 (N_1435,In_115,In_637);
and U1436 (N_1436,In_387,In_936);
nand U1437 (N_1437,In_818,In_281);
and U1438 (N_1438,In_607,In_193);
and U1439 (N_1439,In_743,In_426);
and U1440 (N_1440,In_919,In_687);
and U1441 (N_1441,In_610,In_791);
nand U1442 (N_1442,In_139,In_980);
and U1443 (N_1443,In_754,In_503);
nand U1444 (N_1444,In_975,In_160);
nand U1445 (N_1445,In_870,In_330);
nand U1446 (N_1446,In_132,In_105);
or U1447 (N_1447,In_359,In_614);
nor U1448 (N_1448,In_344,In_24);
nor U1449 (N_1449,In_847,In_654);
and U1450 (N_1450,In_823,In_507);
and U1451 (N_1451,In_355,In_79);
nand U1452 (N_1452,In_197,In_419);
nor U1453 (N_1453,In_334,In_272);
nor U1454 (N_1454,In_524,In_711);
nand U1455 (N_1455,In_630,In_875);
or U1456 (N_1456,In_699,In_69);
and U1457 (N_1457,In_260,In_442);
and U1458 (N_1458,In_658,In_488);
and U1459 (N_1459,In_379,In_243);
nor U1460 (N_1460,In_85,In_408);
nor U1461 (N_1461,In_96,In_765);
and U1462 (N_1462,In_475,In_543);
nand U1463 (N_1463,In_920,In_350);
nand U1464 (N_1464,In_301,In_575);
and U1465 (N_1465,In_69,In_858);
or U1466 (N_1466,In_700,In_538);
nand U1467 (N_1467,In_209,In_229);
or U1468 (N_1468,In_55,In_624);
or U1469 (N_1469,In_796,In_786);
or U1470 (N_1470,In_262,In_399);
and U1471 (N_1471,In_591,In_184);
and U1472 (N_1472,In_899,In_129);
and U1473 (N_1473,In_791,In_338);
nor U1474 (N_1474,In_142,In_720);
and U1475 (N_1475,In_177,In_377);
and U1476 (N_1476,In_445,In_475);
nand U1477 (N_1477,In_882,In_546);
nor U1478 (N_1478,In_178,In_485);
and U1479 (N_1479,In_246,In_832);
or U1480 (N_1480,In_376,In_413);
nor U1481 (N_1481,In_749,In_590);
or U1482 (N_1482,In_814,In_417);
or U1483 (N_1483,In_40,In_498);
and U1484 (N_1484,In_272,In_779);
and U1485 (N_1485,In_63,In_246);
nor U1486 (N_1486,In_398,In_320);
and U1487 (N_1487,In_788,In_539);
and U1488 (N_1488,In_748,In_810);
or U1489 (N_1489,In_427,In_358);
or U1490 (N_1490,In_344,In_389);
and U1491 (N_1491,In_431,In_23);
nand U1492 (N_1492,In_446,In_972);
nor U1493 (N_1493,In_568,In_879);
nor U1494 (N_1494,In_50,In_278);
or U1495 (N_1495,In_255,In_14);
nand U1496 (N_1496,In_446,In_494);
or U1497 (N_1497,In_306,In_673);
or U1498 (N_1498,In_255,In_361);
or U1499 (N_1499,In_363,In_214);
nor U1500 (N_1500,In_966,In_477);
or U1501 (N_1501,In_964,In_228);
nand U1502 (N_1502,In_153,In_251);
nand U1503 (N_1503,In_90,In_605);
nand U1504 (N_1504,In_448,In_287);
nand U1505 (N_1505,In_659,In_124);
and U1506 (N_1506,In_52,In_877);
nand U1507 (N_1507,In_844,In_680);
and U1508 (N_1508,In_916,In_892);
or U1509 (N_1509,In_471,In_722);
or U1510 (N_1510,In_763,In_584);
and U1511 (N_1511,In_685,In_886);
nor U1512 (N_1512,In_341,In_951);
nor U1513 (N_1513,In_239,In_170);
nor U1514 (N_1514,In_7,In_222);
and U1515 (N_1515,In_688,In_661);
nor U1516 (N_1516,In_188,In_917);
nor U1517 (N_1517,In_373,In_896);
nor U1518 (N_1518,In_665,In_572);
nand U1519 (N_1519,In_63,In_927);
nand U1520 (N_1520,In_227,In_710);
nor U1521 (N_1521,In_955,In_342);
and U1522 (N_1522,In_510,In_304);
or U1523 (N_1523,In_541,In_130);
or U1524 (N_1524,In_732,In_44);
or U1525 (N_1525,In_71,In_192);
nor U1526 (N_1526,In_54,In_487);
nand U1527 (N_1527,In_508,In_187);
and U1528 (N_1528,In_571,In_428);
or U1529 (N_1529,In_641,In_275);
and U1530 (N_1530,In_564,In_289);
nor U1531 (N_1531,In_820,In_379);
and U1532 (N_1532,In_905,In_902);
nor U1533 (N_1533,In_286,In_308);
and U1534 (N_1534,In_398,In_16);
and U1535 (N_1535,In_958,In_664);
nor U1536 (N_1536,In_511,In_376);
nor U1537 (N_1537,In_377,In_951);
nor U1538 (N_1538,In_6,In_552);
nand U1539 (N_1539,In_595,In_639);
or U1540 (N_1540,In_457,In_960);
nor U1541 (N_1541,In_873,In_685);
nor U1542 (N_1542,In_24,In_980);
nor U1543 (N_1543,In_793,In_694);
and U1544 (N_1544,In_712,In_628);
and U1545 (N_1545,In_109,In_843);
or U1546 (N_1546,In_497,In_659);
or U1547 (N_1547,In_127,In_500);
and U1548 (N_1548,In_619,In_492);
or U1549 (N_1549,In_881,In_410);
nand U1550 (N_1550,In_772,In_261);
nand U1551 (N_1551,In_57,In_856);
or U1552 (N_1552,In_496,In_790);
nand U1553 (N_1553,In_547,In_56);
nor U1554 (N_1554,In_232,In_602);
or U1555 (N_1555,In_272,In_508);
or U1556 (N_1556,In_194,In_234);
and U1557 (N_1557,In_741,In_592);
nor U1558 (N_1558,In_991,In_533);
nand U1559 (N_1559,In_18,In_800);
nor U1560 (N_1560,In_732,In_798);
or U1561 (N_1561,In_714,In_812);
nor U1562 (N_1562,In_182,In_645);
and U1563 (N_1563,In_46,In_842);
and U1564 (N_1564,In_675,In_823);
or U1565 (N_1565,In_82,In_698);
and U1566 (N_1566,In_530,In_101);
or U1567 (N_1567,In_473,In_53);
nor U1568 (N_1568,In_986,In_781);
and U1569 (N_1569,In_134,In_799);
and U1570 (N_1570,In_284,In_184);
nand U1571 (N_1571,In_381,In_57);
nand U1572 (N_1572,In_203,In_873);
and U1573 (N_1573,In_772,In_33);
nand U1574 (N_1574,In_325,In_14);
and U1575 (N_1575,In_640,In_796);
and U1576 (N_1576,In_292,In_754);
nor U1577 (N_1577,In_107,In_862);
and U1578 (N_1578,In_722,In_26);
or U1579 (N_1579,In_203,In_564);
nand U1580 (N_1580,In_522,In_86);
and U1581 (N_1581,In_764,In_126);
nand U1582 (N_1582,In_120,In_693);
nand U1583 (N_1583,In_998,In_859);
and U1584 (N_1584,In_628,In_288);
or U1585 (N_1585,In_79,In_964);
or U1586 (N_1586,In_516,In_671);
and U1587 (N_1587,In_359,In_871);
nand U1588 (N_1588,In_35,In_746);
nor U1589 (N_1589,In_406,In_393);
or U1590 (N_1590,In_738,In_766);
or U1591 (N_1591,In_826,In_6);
and U1592 (N_1592,In_539,In_46);
and U1593 (N_1593,In_850,In_740);
xor U1594 (N_1594,In_556,In_980);
or U1595 (N_1595,In_903,In_756);
nor U1596 (N_1596,In_440,In_505);
or U1597 (N_1597,In_131,In_922);
nand U1598 (N_1598,In_949,In_535);
or U1599 (N_1599,In_428,In_315);
nor U1600 (N_1600,In_569,In_868);
nor U1601 (N_1601,In_733,In_503);
or U1602 (N_1602,In_921,In_36);
nand U1603 (N_1603,In_113,In_793);
nor U1604 (N_1604,In_334,In_114);
nor U1605 (N_1605,In_169,In_433);
or U1606 (N_1606,In_360,In_440);
and U1607 (N_1607,In_779,In_590);
or U1608 (N_1608,In_106,In_691);
nand U1609 (N_1609,In_376,In_15);
nor U1610 (N_1610,In_690,In_474);
or U1611 (N_1611,In_620,In_516);
nor U1612 (N_1612,In_620,In_38);
or U1613 (N_1613,In_723,In_838);
nor U1614 (N_1614,In_143,In_824);
and U1615 (N_1615,In_983,In_339);
or U1616 (N_1616,In_336,In_276);
nand U1617 (N_1617,In_355,In_780);
and U1618 (N_1618,In_847,In_323);
nor U1619 (N_1619,In_430,In_600);
nand U1620 (N_1620,In_347,In_329);
nand U1621 (N_1621,In_294,In_392);
nor U1622 (N_1622,In_698,In_972);
nor U1623 (N_1623,In_440,In_572);
or U1624 (N_1624,In_694,In_565);
nor U1625 (N_1625,In_978,In_160);
and U1626 (N_1626,In_333,In_511);
xnor U1627 (N_1627,In_995,In_903);
nor U1628 (N_1628,In_611,In_314);
and U1629 (N_1629,In_505,In_265);
nand U1630 (N_1630,In_709,In_443);
nand U1631 (N_1631,In_541,In_622);
or U1632 (N_1632,In_809,In_920);
and U1633 (N_1633,In_577,In_190);
nand U1634 (N_1634,In_568,In_792);
nor U1635 (N_1635,In_95,In_330);
nor U1636 (N_1636,In_19,In_851);
nor U1637 (N_1637,In_863,In_50);
and U1638 (N_1638,In_647,In_985);
or U1639 (N_1639,In_920,In_1);
and U1640 (N_1640,In_662,In_460);
and U1641 (N_1641,In_687,In_710);
nand U1642 (N_1642,In_528,In_434);
and U1643 (N_1643,In_615,In_507);
and U1644 (N_1644,In_499,In_920);
xor U1645 (N_1645,In_522,In_842);
and U1646 (N_1646,In_928,In_341);
nand U1647 (N_1647,In_160,In_669);
nand U1648 (N_1648,In_675,In_781);
and U1649 (N_1649,In_65,In_184);
and U1650 (N_1650,In_664,In_368);
nor U1651 (N_1651,In_855,In_952);
and U1652 (N_1652,In_708,In_948);
and U1653 (N_1653,In_279,In_57);
nor U1654 (N_1654,In_145,In_975);
nand U1655 (N_1655,In_504,In_823);
and U1656 (N_1656,In_916,In_584);
and U1657 (N_1657,In_43,In_289);
or U1658 (N_1658,In_846,In_493);
or U1659 (N_1659,In_302,In_94);
and U1660 (N_1660,In_881,In_497);
or U1661 (N_1661,In_356,In_129);
nand U1662 (N_1662,In_670,In_990);
nor U1663 (N_1663,In_775,In_463);
nor U1664 (N_1664,In_422,In_76);
or U1665 (N_1665,In_48,In_395);
nor U1666 (N_1666,In_957,In_866);
nor U1667 (N_1667,In_541,In_323);
nor U1668 (N_1668,In_390,In_176);
nand U1669 (N_1669,In_8,In_78);
nor U1670 (N_1670,In_316,In_372);
nor U1671 (N_1671,In_660,In_356);
or U1672 (N_1672,In_768,In_458);
or U1673 (N_1673,In_95,In_947);
nor U1674 (N_1674,In_599,In_469);
or U1675 (N_1675,In_303,In_619);
nand U1676 (N_1676,In_24,In_582);
and U1677 (N_1677,In_908,In_586);
nand U1678 (N_1678,In_510,In_523);
or U1679 (N_1679,In_340,In_84);
nor U1680 (N_1680,In_210,In_226);
nand U1681 (N_1681,In_953,In_631);
or U1682 (N_1682,In_931,In_582);
and U1683 (N_1683,In_871,In_912);
or U1684 (N_1684,In_681,In_408);
nor U1685 (N_1685,In_968,In_747);
and U1686 (N_1686,In_828,In_374);
or U1687 (N_1687,In_82,In_840);
and U1688 (N_1688,In_982,In_752);
or U1689 (N_1689,In_147,In_866);
nor U1690 (N_1690,In_364,In_694);
or U1691 (N_1691,In_5,In_12);
and U1692 (N_1692,In_966,In_46);
nand U1693 (N_1693,In_714,In_88);
nand U1694 (N_1694,In_768,In_644);
nor U1695 (N_1695,In_217,In_399);
nand U1696 (N_1696,In_270,In_57);
and U1697 (N_1697,In_832,In_181);
and U1698 (N_1698,In_249,In_333);
or U1699 (N_1699,In_115,In_852);
nor U1700 (N_1700,In_79,In_813);
and U1701 (N_1701,In_952,In_636);
nand U1702 (N_1702,In_399,In_470);
nand U1703 (N_1703,In_945,In_817);
and U1704 (N_1704,In_571,In_10);
or U1705 (N_1705,In_793,In_704);
nand U1706 (N_1706,In_544,In_435);
xnor U1707 (N_1707,In_415,In_552);
and U1708 (N_1708,In_289,In_359);
or U1709 (N_1709,In_14,In_86);
and U1710 (N_1710,In_51,In_383);
nor U1711 (N_1711,In_667,In_272);
and U1712 (N_1712,In_466,In_802);
and U1713 (N_1713,In_853,In_992);
nor U1714 (N_1714,In_70,In_28);
and U1715 (N_1715,In_748,In_591);
nand U1716 (N_1716,In_643,In_712);
or U1717 (N_1717,In_463,In_732);
nor U1718 (N_1718,In_922,In_785);
nor U1719 (N_1719,In_561,In_804);
and U1720 (N_1720,In_455,In_319);
or U1721 (N_1721,In_977,In_391);
nor U1722 (N_1722,In_767,In_875);
or U1723 (N_1723,In_672,In_560);
and U1724 (N_1724,In_110,In_441);
and U1725 (N_1725,In_413,In_473);
or U1726 (N_1726,In_828,In_168);
nor U1727 (N_1727,In_278,In_478);
or U1728 (N_1728,In_193,In_39);
nor U1729 (N_1729,In_653,In_976);
and U1730 (N_1730,In_371,In_423);
or U1731 (N_1731,In_378,In_571);
and U1732 (N_1732,In_717,In_633);
nor U1733 (N_1733,In_195,In_111);
and U1734 (N_1734,In_9,In_25);
nand U1735 (N_1735,In_198,In_4);
and U1736 (N_1736,In_586,In_273);
nand U1737 (N_1737,In_491,In_18);
nand U1738 (N_1738,In_214,In_428);
nand U1739 (N_1739,In_800,In_937);
nand U1740 (N_1740,In_306,In_879);
nor U1741 (N_1741,In_216,In_597);
or U1742 (N_1742,In_717,In_423);
nand U1743 (N_1743,In_964,In_979);
nor U1744 (N_1744,In_233,In_824);
nand U1745 (N_1745,In_723,In_457);
and U1746 (N_1746,In_256,In_594);
and U1747 (N_1747,In_493,In_510);
and U1748 (N_1748,In_369,In_292);
or U1749 (N_1749,In_540,In_57);
nor U1750 (N_1750,In_84,In_122);
nand U1751 (N_1751,In_730,In_79);
and U1752 (N_1752,In_8,In_2);
or U1753 (N_1753,In_642,In_835);
and U1754 (N_1754,In_592,In_338);
and U1755 (N_1755,In_273,In_94);
nor U1756 (N_1756,In_220,In_583);
or U1757 (N_1757,In_399,In_879);
and U1758 (N_1758,In_563,In_740);
nor U1759 (N_1759,In_244,In_675);
nor U1760 (N_1760,In_168,In_285);
nand U1761 (N_1761,In_615,In_582);
and U1762 (N_1762,In_122,In_800);
nand U1763 (N_1763,In_372,In_717);
nand U1764 (N_1764,In_598,In_480);
and U1765 (N_1765,In_743,In_123);
and U1766 (N_1766,In_370,In_774);
or U1767 (N_1767,In_63,In_157);
and U1768 (N_1768,In_896,In_426);
and U1769 (N_1769,In_626,In_485);
and U1770 (N_1770,In_62,In_526);
nand U1771 (N_1771,In_810,In_353);
and U1772 (N_1772,In_19,In_331);
and U1773 (N_1773,In_65,In_987);
and U1774 (N_1774,In_405,In_11);
nor U1775 (N_1775,In_377,In_587);
nand U1776 (N_1776,In_390,In_905);
or U1777 (N_1777,In_917,In_203);
nand U1778 (N_1778,In_505,In_882);
or U1779 (N_1779,In_762,In_825);
and U1780 (N_1780,In_249,In_260);
and U1781 (N_1781,In_627,In_891);
nand U1782 (N_1782,In_393,In_70);
nand U1783 (N_1783,In_40,In_582);
nand U1784 (N_1784,In_877,In_228);
and U1785 (N_1785,In_474,In_686);
and U1786 (N_1786,In_885,In_436);
nand U1787 (N_1787,In_331,In_897);
or U1788 (N_1788,In_276,In_324);
and U1789 (N_1789,In_712,In_261);
or U1790 (N_1790,In_531,In_270);
or U1791 (N_1791,In_487,In_951);
nor U1792 (N_1792,In_420,In_546);
nor U1793 (N_1793,In_487,In_298);
and U1794 (N_1794,In_243,In_655);
nor U1795 (N_1795,In_980,In_628);
nand U1796 (N_1796,In_717,In_321);
nand U1797 (N_1797,In_356,In_541);
and U1798 (N_1798,In_845,In_690);
or U1799 (N_1799,In_336,In_73);
xor U1800 (N_1800,In_39,In_615);
nor U1801 (N_1801,In_376,In_690);
or U1802 (N_1802,In_497,In_287);
or U1803 (N_1803,In_186,In_689);
or U1804 (N_1804,In_285,In_607);
nor U1805 (N_1805,In_651,In_360);
nor U1806 (N_1806,In_581,In_397);
nor U1807 (N_1807,In_285,In_836);
or U1808 (N_1808,In_357,In_546);
or U1809 (N_1809,In_161,In_638);
or U1810 (N_1810,In_233,In_802);
nand U1811 (N_1811,In_984,In_485);
and U1812 (N_1812,In_848,In_617);
or U1813 (N_1813,In_25,In_694);
nor U1814 (N_1814,In_309,In_607);
nor U1815 (N_1815,In_366,In_265);
or U1816 (N_1816,In_614,In_381);
or U1817 (N_1817,In_59,In_966);
and U1818 (N_1818,In_776,In_839);
nand U1819 (N_1819,In_267,In_226);
nand U1820 (N_1820,In_636,In_160);
nand U1821 (N_1821,In_822,In_387);
or U1822 (N_1822,In_564,In_594);
nand U1823 (N_1823,In_505,In_487);
nand U1824 (N_1824,In_294,In_408);
or U1825 (N_1825,In_995,In_144);
and U1826 (N_1826,In_190,In_203);
nand U1827 (N_1827,In_761,In_601);
nor U1828 (N_1828,In_535,In_534);
or U1829 (N_1829,In_68,In_731);
or U1830 (N_1830,In_609,In_359);
and U1831 (N_1831,In_756,In_577);
nand U1832 (N_1832,In_481,In_77);
nand U1833 (N_1833,In_489,In_559);
and U1834 (N_1834,In_601,In_237);
or U1835 (N_1835,In_650,In_385);
nor U1836 (N_1836,In_691,In_243);
nand U1837 (N_1837,In_715,In_174);
and U1838 (N_1838,In_594,In_17);
nor U1839 (N_1839,In_733,In_604);
and U1840 (N_1840,In_420,In_652);
or U1841 (N_1841,In_386,In_526);
nand U1842 (N_1842,In_546,In_494);
nand U1843 (N_1843,In_822,In_700);
or U1844 (N_1844,In_722,In_922);
nand U1845 (N_1845,In_705,In_38);
and U1846 (N_1846,In_440,In_235);
and U1847 (N_1847,In_928,In_439);
nor U1848 (N_1848,In_229,In_647);
and U1849 (N_1849,In_116,In_580);
or U1850 (N_1850,In_880,In_281);
or U1851 (N_1851,In_14,In_242);
and U1852 (N_1852,In_432,In_856);
or U1853 (N_1853,In_520,In_366);
nand U1854 (N_1854,In_423,In_968);
nand U1855 (N_1855,In_366,In_246);
nand U1856 (N_1856,In_579,In_491);
nand U1857 (N_1857,In_592,In_356);
or U1858 (N_1858,In_337,In_181);
and U1859 (N_1859,In_510,In_943);
or U1860 (N_1860,In_464,In_755);
or U1861 (N_1861,In_713,In_958);
nand U1862 (N_1862,In_830,In_170);
nor U1863 (N_1863,In_412,In_190);
nand U1864 (N_1864,In_938,In_570);
nor U1865 (N_1865,In_415,In_652);
nor U1866 (N_1866,In_568,In_107);
nand U1867 (N_1867,In_272,In_134);
and U1868 (N_1868,In_927,In_42);
and U1869 (N_1869,In_508,In_448);
nor U1870 (N_1870,In_223,In_524);
nand U1871 (N_1871,In_834,In_209);
nor U1872 (N_1872,In_725,In_615);
or U1873 (N_1873,In_638,In_790);
or U1874 (N_1874,In_822,In_453);
or U1875 (N_1875,In_589,In_35);
nand U1876 (N_1876,In_419,In_913);
or U1877 (N_1877,In_90,In_976);
and U1878 (N_1878,In_912,In_964);
and U1879 (N_1879,In_80,In_730);
and U1880 (N_1880,In_462,In_182);
nor U1881 (N_1881,In_901,In_804);
nand U1882 (N_1882,In_986,In_768);
and U1883 (N_1883,In_839,In_954);
nor U1884 (N_1884,In_134,In_444);
nor U1885 (N_1885,In_90,In_829);
and U1886 (N_1886,In_785,In_863);
or U1887 (N_1887,In_246,In_647);
xnor U1888 (N_1888,In_90,In_216);
nand U1889 (N_1889,In_785,In_715);
or U1890 (N_1890,In_304,In_568);
nor U1891 (N_1891,In_852,In_334);
or U1892 (N_1892,In_78,In_271);
nor U1893 (N_1893,In_267,In_62);
and U1894 (N_1894,In_944,In_92);
nor U1895 (N_1895,In_564,In_340);
and U1896 (N_1896,In_606,In_979);
nor U1897 (N_1897,In_266,In_133);
nor U1898 (N_1898,In_163,In_333);
and U1899 (N_1899,In_419,In_614);
nand U1900 (N_1900,In_531,In_977);
or U1901 (N_1901,In_644,In_139);
and U1902 (N_1902,In_719,In_923);
or U1903 (N_1903,In_536,In_6);
nor U1904 (N_1904,In_525,In_547);
nor U1905 (N_1905,In_764,In_381);
and U1906 (N_1906,In_852,In_992);
or U1907 (N_1907,In_661,In_557);
or U1908 (N_1908,In_451,In_794);
and U1909 (N_1909,In_599,In_630);
and U1910 (N_1910,In_373,In_960);
and U1911 (N_1911,In_457,In_863);
and U1912 (N_1912,In_733,In_764);
nor U1913 (N_1913,In_936,In_37);
nand U1914 (N_1914,In_573,In_605);
nor U1915 (N_1915,In_537,In_444);
and U1916 (N_1916,In_313,In_970);
and U1917 (N_1917,In_647,In_648);
nor U1918 (N_1918,In_257,In_6);
nor U1919 (N_1919,In_236,In_559);
nor U1920 (N_1920,In_356,In_823);
and U1921 (N_1921,In_793,In_710);
and U1922 (N_1922,In_518,In_406);
and U1923 (N_1923,In_97,In_151);
or U1924 (N_1924,In_793,In_668);
nor U1925 (N_1925,In_61,In_600);
xor U1926 (N_1926,In_467,In_180);
and U1927 (N_1927,In_193,In_469);
nand U1928 (N_1928,In_990,In_913);
nand U1929 (N_1929,In_937,In_660);
and U1930 (N_1930,In_253,In_218);
or U1931 (N_1931,In_617,In_341);
nor U1932 (N_1932,In_342,In_605);
nor U1933 (N_1933,In_658,In_570);
and U1934 (N_1934,In_424,In_47);
nand U1935 (N_1935,In_811,In_182);
nand U1936 (N_1936,In_63,In_559);
nor U1937 (N_1937,In_288,In_97);
or U1938 (N_1938,In_960,In_876);
nand U1939 (N_1939,In_820,In_467);
and U1940 (N_1940,In_879,In_467);
xor U1941 (N_1941,In_281,In_642);
and U1942 (N_1942,In_766,In_589);
nand U1943 (N_1943,In_568,In_29);
or U1944 (N_1944,In_537,In_536);
nor U1945 (N_1945,In_423,In_359);
nor U1946 (N_1946,In_718,In_76);
or U1947 (N_1947,In_261,In_715);
and U1948 (N_1948,In_763,In_726);
nand U1949 (N_1949,In_257,In_219);
nand U1950 (N_1950,In_258,In_61);
nor U1951 (N_1951,In_328,In_914);
nor U1952 (N_1952,In_386,In_413);
nand U1953 (N_1953,In_571,In_642);
nor U1954 (N_1954,In_954,In_854);
nor U1955 (N_1955,In_459,In_57);
nor U1956 (N_1956,In_479,In_180);
or U1957 (N_1957,In_421,In_499);
or U1958 (N_1958,In_292,In_770);
or U1959 (N_1959,In_131,In_610);
and U1960 (N_1960,In_210,In_685);
nand U1961 (N_1961,In_638,In_929);
nor U1962 (N_1962,In_707,In_403);
and U1963 (N_1963,In_970,In_766);
and U1964 (N_1964,In_397,In_762);
or U1965 (N_1965,In_114,In_272);
and U1966 (N_1966,In_265,In_702);
or U1967 (N_1967,In_125,In_892);
xor U1968 (N_1968,In_207,In_575);
nor U1969 (N_1969,In_91,In_165);
and U1970 (N_1970,In_348,In_705);
nand U1971 (N_1971,In_423,In_313);
or U1972 (N_1972,In_808,In_184);
or U1973 (N_1973,In_652,In_690);
and U1974 (N_1974,In_569,In_650);
or U1975 (N_1975,In_301,In_361);
and U1976 (N_1976,In_456,In_74);
nor U1977 (N_1977,In_582,In_407);
nor U1978 (N_1978,In_796,In_654);
or U1979 (N_1979,In_28,In_617);
and U1980 (N_1980,In_676,In_222);
or U1981 (N_1981,In_660,In_407);
and U1982 (N_1982,In_1,In_909);
nand U1983 (N_1983,In_784,In_227);
or U1984 (N_1984,In_389,In_479);
nand U1985 (N_1985,In_87,In_666);
nand U1986 (N_1986,In_583,In_419);
nand U1987 (N_1987,In_558,In_300);
nor U1988 (N_1988,In_13,In_316);
nand U1989 (N_1989,In_757,In_552);
nand U1990 (N_1990,In_945,In_394);
nor U1991 (N_1991,In_202,In_557);
or U1992 (N_1992,In_527,In_30);
nor U1993 (N_1993,In_181,In_407);
and U1994 (N_1994,In_404,In_682);
nand U1995 (N_1995,In_322,In_110);
nor U1996 (N_1996,In_255,In_108);
nand U1997 (N_1997,In_39,In_113);
nor U1998 (N_1998,In_18,In_356);
and U1999 (N_1999,In_902,In_758);
and U2000 (N_2000,In_340,In_310);
and U2001 (N_2001,In_438,In_706);
and U2002 (N_2002,In_711,In_585);
nor U2003 (N_2003,In_817,In_3);
nand U2004 (N_2004,In_65,In_673);
nand U2005 (N_2005,In_39,In_905);
or U2006 (N_2006,In_694,In_187);
nor U2007 (N_2007,In_143,In_934);
nor U2008 (N_2008,In_534,In_739);
nor U2009 (N_2009,In_742,In_933);
and U2010 (N_2010,In_883,In_996);
nand U2011 (N_2011,In_634,In_837);
nor U2012 (N_2012,In_48,In_709);
and U2013 (N_2013,In_314,In_474);
and U2014 (N_2014,In_89,In_432);
nand U2015 (N_2015,In_222,In_707);
or U2016 (N_2016,In_695,In_84);
and U2017 (N_2017,In_417,In_495);
nand U2018 (N_2018,In_896,In_444);
nand U2019 (N_2019,In_535,In_554);
and U2020 (N_2020,In_841,In_270);
or U2021 (N_2021,In_411,In_541);
or U2022 (N_2022,In_215,In_652);
or U2023 (N_2023,In_600,In_347);
nor U2024 (N_2024,In_527,In_376);
or U2025 (N_2025,In_930,In_297);
and U2026 (N_2026,In_818,In_189);
nand U2027 (N_2027,In_38,In_950);
or U2028 (N_2028,In_122,In_337);
and U2029 (N_2029,In_226,In_559);
or U2030 (N_2030,In_128,In_867);
nand U2031 (N_2031,In_549,In_83);
nand U2032 (N_2032,In_380,In_594);
nor U2033 (N_2033,In_946,In_50);
or U2034 (N_2034,In_932,In_927);
nand U2035 (N_2035,In_15,In_452);
and U2036 (N_2036,In_406,In_754);
and U2037 (N_2037,In_797,In_249);
or U2038 (N_2038,In_822,In_619);
or U2039 (N_2039,In_665,In_915);
nand U2040 (N_2040,In_609,In_55);
or U2041 (N_2041,In_40,In_657);
or U2042 (N_2042,In_51,In_39);
and U2043 (N_2043,In_298,In_506);
nand U2044 (N_2044,In_485,In_240);
xor U2045 (N_2045,In_296,In_133);
or U2046 (N_2046,In_520,In_215);
nor U2047 (N_2047,In_510,In_315);
nand U2048 (N_2048,In_199,In_914);
and U2049 (N_2049,In_822,In_454);
or U2050 (N_2050,In_240,In_520);
nand U2051 (N_2051,In_497,In_920);
nand U2052 (N_2052,In_681,In_567);
nand U2053 (N_2053,In_571,In_235);
or U2054 (N_2054,In_647,In_35);
nand U2055 (N_2055,In_61,In_707);
or U2056 (N_2056,In_96,In_342);
nor U2057 (N_2057,In_6,In_582);
or U2058 (N_2058,In_632,In_238);
nor U2059 (N_2059,In_352,In_904);
and U2060 (N_2060,In_629,In_738);
and U2061 (N_2061,In_53,In_8);
nor U2062 (N_2062,In_717,In_679);
nand U2063 (N_2063,In_656,In_623);
nor U2064 (N_2064,In_12,In_278);
nor U2065 (N_2065,In_830,In_530);
nand U2066 (N_2066,In_614,In_7);
nor U2067 (N_2067,In_273,In_335);
nand U2068 (N_2068,In_754,In_689);
nor U2069 (N_2069,In_812,In_929);
nor U2070 (N_2070,In_277,In_647);
nand U2071 (N_2071,In_146,In_392);
or U2072 (N_2072,In_194,In_187);
and U2073 (N_2073,In_823,In_166);
and U2074 (N_2074,In_181,In_541);
nand U2075 (N_2075,In_673,In_734);
nand U2076 (N_2076,In_422,In_171);
or U2077 (N_2077,In_43,In_956);
or U2078 (N_2078,In_133,In_635);
nor U2079 (N_2079,In_74,In_929);
nand U2080 (N_2080,In_588,In_9);
or U2081 (N_2081,In_188,In_140);
or U2082 (N_2082,In_800,In_125);
or U2083 (N_2083,In_868,In_496);
nand U2084 (N_2084,In_857,In_816);
nand U2085 (N_2085,In_3,In_552);
nand U2086 (N_2086,In_634,In_670);
or U2087 (N_2087,In_23,In_271);
or U2088 (N_2088,In_259,In_582);
or U2089 (N_2089,In_528,In_871);
nand U2090 (N_2090,In_492,In_624);
or U2091 (N_2091,In_175,In_416);
nand U2092 (N_2092,In_727,In_615);
and U2093 (N_2093,In_174,In_32);
nor U2094 (N_2094,In_374,In_124);
nand U2095 (N_2095,In_889,In_672);
and U2096 (N_2096,In_5,In_705);
nand U2097 (N_2097,In_429,In_469);
nand U2098 (N_2098,In_727,In_706);
nor U2099 (N_2099,In_454,In_99);
xnor U2100 (N_2100,In_381,In_543);
or U2101 (N_2101,In_757,In_359);
nor U2102 (N_2102,In_434,In_547);
nor U2103 (N_2103,In_628,In_603);
or U2104 (N_2104,In_422,In_706);
nor U2105 (N_2105,In_700,In_62);
and U2106 (N_2106,In_543,In_778);
or U2107 (N_2107,In_511,In_394);
and U2108 (N_2108,In_631,In_2);
or U2109 (N_2109,In_326,In_61);
nand U2110 (N_2110,In_650,In_564);
nor U2111 (N_2111,In_509,In_720);
or U2112 (N_2112,In_617,In_767);
and U2113 (N_2113,In_874,In_809);
and U2114 (N_2114,In_468,In_183);
nor U2115 (N_2115,In_826,In_550);
nor U2116 (N_2116,In_609,In_824);
or U2117 (N_2117,In_567,In_954);
nor U2118 (N_2118,In_863,In_262);
or U2119 (N_2119,In_800,In_765);
nor U2120 (N_2120,In_346,In_634);
or U2121 (N_2121,In_783,In_991);
nor U2122 (N_2122,In_948,In_900);
nor U2123 (N_2123,In_551,In_511);
and U2124 (N_2124,In_240,In_997);
nand U2125 (N_2125,In_319,In_832);
and U2126 (N_2126,In_666,In_547);
and U2127 (N_2127,In_65,In_675);
nand U2128 (N_2128,In_831,In_366);
or U2129 (N_2129,In_261,In_195);
xnor U2130 (N_2130,In_818,In_179);
and U2131 (N_2131,In_358,In_261);
nor U2132 (N_2132,In_958,In_178);
nand U2133 (N_2133,In_445,In_119);
and U2134 (N_2134,In_302,In_630);
nand U2135 (N_2135,In_537,In_361);
nand U2136 (N_2136,In_799,In_706);
nor U2137 (N_2137,In_950,In_70);
nor U2138 (N_2138,In_190,In_276);
nand U2139 (N_2139,In_513,In_662);
nand U2140 (N_2140,In_366,In_232);
nor U2141 (N_2141,In_857,In_307);
nor U2142 (N_2142,In_955,In_850);
nor U2143 (N_2143,In_357,In_375);
or U2144 (N_2144,In_904,In_261);
nor U2145 (N_2145,In_347,In_652);
nor U2146 (N_2146,In_825,In_98);
nand U2147 (N_2147,In_682,In_259);
nor U2148 (N_2148,In_820,In_401);
or U2149 (N_2149,In_462,In_305);
nor U2150 (N_2150,In_603,In_447);
nor U2151 (N_2151,In_317,In_572);
nor U2152 (N_2152,In_975,In_306);
nand U2153 (N_2153,In_26,In_802);
nor U2154 (N_2154,In_658,In_827);
and U2155 (N_2155,In_901,In_101);
nor U2156 (N_2156,In_913,In_732);
nand U2157 (N_2157,In_829,In_942);
nand U2158 (N_2158,In_396,In_410);
and U2159 (N_2159,In_148,In_771);
nand U2160 (N_2160,In_180,In_957);
nor U2161 (N_2161,In_228,In_194);
nor U2162 (N_2162,In_583,In_38);
or U2163 (N_2163,In_60,In_876);
nand U2164 (N_2164,In_696,In_758);
nand U2165 (N_2165,In_420,In_522);
nor U2166 (N_2166,In_49,In_942);
and U2167 (N_2167,In_921,In_215);
or U2168 (N_2168,In_68,In_918);
nor U2169 (N_2169,In_92,In_911);
or U2170 (N_2170,In_916,In_739);
and U2171 (N_2171,In_238,In_107);
nor U2172 (N_2172,In_91,In_240);
or U2173 (N_2173,In_875,In_512);
and U2174 (N_2174,In_546,In_205);
or U2175 (N_2175,In_698,In_679);
and U2176 (N_2176,In_368,In_915);
nand U2177 (N_2177,In_578,In_525);
nor U2178 (N_2178,In_806,In_456);
or U2179 (N_2179,In_386,In_687);
nor U2180 (N_2180,In_684,In_596);
or U2181 (N_2181,In_480,In_841);
and U2182 (N_2182,In_140,In_334);
nand U2183 (N_2183,In_204,In_808);
and U2184 (N_2184,In_206,In_545);
nand U2185 (N_2185,In_761,In_205);
and U2186 (N_2186,In_168,In_281);
or U2187 (N_2187,In_700,In_74);
and U2188 (N_2188,In_578,In_3);
nand U2189 (N_2189,In_135,In_211);
nand U2190 (N_2190,In_248,In_210);
and U2191 (N_2191,In_715,In_485);
or U2192 (N_2192,In_3,In_279);
nand U2193 (N_2193,In_92,In_332);
nor U2194 (N_2194,In_125,In_470);
or U2195 (N_2195,In_460,In_636);
nor U2196 (N_2196,In_693,In_571);
nand U2197 (N_2197,In_586,In_365);
nor U2198 (N_2198,In_185,In_574);
and U2199 (N_2199,In_361,In_881);
nor U2200 (N_2200,In_110,In_998);
nor U2201 (N_2201,In_437,In_170);
or U2202 (N_2202,In_865,In_238);
or U2203 (N_2203,In_892,In_309);
nor U2204 (N_2204,In_596,In_71);
or U2205 (N_2205,In_316,In_87);
or U2206 (N_2206,In_961,In_801);
or U2207 (N_2207,In_73,In_104);
nand U2208 (N_2208,In_589,In_498);
or U2209 (N_2209,In_566,In_772);
and U2210 (N_2210,In_290,In_19);
nor U2211 (N_2211,In_49,In_374);
nor U2212 (N_2212,In_676,In_77);
and U2213 (N_2213,In_406,In_419);
nand U2214 (N_2214,In_304,In_363);
nor U2215 (N_2215,In_656,In_131);
nand U2216 (N_2216,In_380,In_669);
or U2217 (N_2217,In_376,In_785);
nor U2218 (N_2218,In_751,In_499);
nor U2219 (N_2219,In_511,In_140);
or U2220 (N_2220,In_480,In_535);
nand U2221 (N_2221,In_125,In_479);
or U2222 (N_2222,In_100,In_981);
nand U2223 (N_2223,In_25,In_971);
and U2224 (N_2224,In_365,In_960);
or U2225 (N_2225,In_466,In_242);
nand U2226 (N_2226,In_193,In_853);
and U2227 (N_2227,In_312,In_212);
or U2228 (N_2228,In_710,In_672);
or U2229 (N_2229,In_532,In_791);
nor U2230 (N_2230,In_225,In_629);
nand U2231 (N_2231,In_365,In_796);
nor U2232 (N_2232,In_770,In_416);
and U2233 (N_2233,In_45,In_570);
or U2234 (N_2234,In_128,In_556);
or U2235 (N_2235,In_214,In_152);
nor U2236 (N_2236,In_859,In_55);
nand U2237 (N_2237,In_140,In_796);
and U2238 (N_2238,In_390,In_821);
and U2239 (N_2239,In_253,In_256);
and U2240 (N_2240,In_999,In_732);
or U2241 (N_2241,In_568,In_886);
nand U2242 (N_2242,In_814,In_749);
nor U2243 (N_2243,In_403,In_874);
nand U2244 (N_2244,In_194,In_559);
nand U2245 (N_2245,In_986,In_279);
or U2246 (N_2246,In_25,In_877);
or U2247 (N_2247,In_277,In_784);
nor U2248 (N_2248,In_691,In_178);
nor U2249 (N_2249,In_73,In_468);
nor U2250 (N_2250,In_719,In_348);
nor U2251 (N_2251,In_640,In_438);
nor U2252 (N_2252,In_518,In_632);
nor U2253 (N_2253,In_641,In_605);
nand U2254 (N_2254,In_210,In_584);
or U2255 (N_2255,In_84,In_884);
or U2256 (N_2256,In_790,In_331);
and U2257 (N_2257,In_261,In_122);
nor U2258 (N_2258,In_599,In_392);
nor U2259 (N_2259,In_457,In_117);
and U2260 (N_2260,In_991,In_809);
or U2261 (N_2261,In_465,In_79);
nand U2262 (N_2262,In_26,In_585);
and U2263 (N_2263,In_822,In_261);
nand U2264 (N_2264,In_512,In_710);
and U2265 (N_2265,In_395,In_628);
and U2266 (N_2266,In_837,In_227);
and U2267 (N_2267,In_294,In_995);
nand U2268 (N_2268,In_736,In_764);
nor U2269 (N_2269,In_45,In_209);
or U2270 (N_2270,In_423,In_604);
or U2271 (N_2271,In_40,In_431);
and U2272 (N_2272,In_792,In_392);
nand U2273 (N_2273,In_928,In_421);
and U2274 (N_2274,In_101,In_662);
and U2275 (N_2275,In_770,In_848);
or U2276 (N_2276,In_96,In_576);
nor U2277 (N_2277,In_786,In_602);
and U2278 (N_2278,In_241,In_227);
nor U2279 (N_2279,In_417,In_298);
and U2280 (N_2280,In_984,In_171);
nand U2281 (N_2281,In_674,In_892);
or U2282 (N_2282,In_548,In_993);
nand U2283 (N_2283,In_834,In_51);
nand U2284 (N_2284,In_865,In_842);
nand U2285 (N_2285,In_517,In_104);
nand U2286 (N_2286,In_918,In_845);
nor U2287 (N_2287,In_56,In_713);
or U2288 (N_2288,In_380,In_742);
nor U2289 (N_2289,In_935,In_948);
nand U2290 (N_2290,In_748,In_716);
nor U2291 (N_2291,In_431,In_770);
nor U2292 (N_2292,In_631,In_335);
or U2293 (N_2293,In_141,In_176);
nor U2294 (N_2294,In_840,In_880);
nor U2295 (N_2295,In_908,In_512);
or U2296 (N_2296,In_17,In_668);
and U2297 (N_2297,In_71,In_689);
nor U2298 (N_2298,In_124,In_658);
nor U2299 (N_2299,In_673,In_146);
or U2300 (N_2300,In_112,In_538);
or U2301 (N_2301,In_135,In_816);
nor U2302 (N_2302,In_471,In_133);
nand U2303 (N_2303,In_798,In_348);
nand U2304 (N_2304,In_989,In_404);
nand U2305 (N_2305,In_967,In_470);
nand U2306 (N_2306,In_664,In_671);
nand U2307 (N_2307,In_854,In_774);
or U2308 (N_2308,In_618,In_561);
nand U2309 (N_2309,In_315,In_988);
nor U2310 (N_2310,In_126,In_894);
and U2311 (N_2311,In_358,In_779);
and U2312 (N_2312,In_474,In_69);
and U2313 (N_2313,In_76,In_513);
or U2314 (N_2314,In_344,In_770);
nor U2315 (N_2315,In_8,In_552);
and U2316 (N_2316,In_729,In_663);
or U2317 (N_2317,In_825,In_562);
nor U2318 (N_2318,In_356,In_188);
or U2319 (N_2319,In_32,In_375);
and U2320 (N_2320,In_340,In_59);
nor U2321 (N_2321,In_626,In_614);
or U2322 (N_2322,In_316,In_190);
nand U2323 (N_2323,In_568,In_761);
nand U2324 (N_2324,In_340,In_304);
and U2325 (N_2325,In_834,In_839);
or U2326 (N_2326,In_861,In_834);
nand U2327 (N_2327,In_294,In_758);
or U2328 (N_2328,In_298,In_871);
and U2329 (N_2329,In_741,In_63);
nand U2330 (N_2330,In_168,In_299);
nand U2331 (N_2331,In_86,In_173);
and U2332 (N_2332,In_756,In_84);
nand U2333 (N_2333,In_787,In_978);
and U2334 (N_2334,In_719,In_547);
nor U2335 (N_2335,In_602,In_893);
and U2336 (N_2336,In_318,In_22);
or U2337 (N_2337,In_956,In_542);
and U2338 (N_2338,In_228,In_327);
or U2339 (N_2339,In_673,In_189);
nand U2340 (N_2340,In_366,In_697);
nor U2341 (N_2341,In_732,In_343);
nor U2342 (N_2342,In_923,In_59);
and U2343 (N_2343,In_811,In_378);
and U2344 (N_2344,In_632,In_207);
nand U2345 (N_2345,In_385,In_624);
and U2346 (N_2346,In_36,In_290);
and U2347 (N_2347,In_553,In_465);
nand U2348 (N_2348,In_800,In_640);
or U2349 (N_2349,In_691,In_707);
nor U2350 (N_2350,In_689,In_291);
and U2351 (N_2351,In_37,In_759);
or U2352 (N_2352,In_852,In_730);
or U2353 (N_2353,In_924,In_828);
or U2354 (N_2354,In_860,In_874);
nor U2355 (N_2355,In_41,In_165);
nor U2356 (N_2356,In_204,In_299);
and U2357 (N_2357,In_757,In_947);
or U2358 (N_2358,In_974,In_433);
and U2359 (N_2359,In_996,In_409);
nor U2360 (N_2360,In_621,In_202);
or U2361 (N_2361,In_301,In_457);
and U2362 (N_2362,In_881,In_692);
nand U2363 (N_2363,In_807,In_900);
nor U2364 (N_2364,In_725,In_129);
nor U2365 (N_2365,In_135,In_902);
or U2366 (N_2366,In_505,In_728);
or U2367 (N_2367,In_74,In_739);
or U2368 (N_2368,In_150,In_440);
nand U2369 (N_2369,In_36,In_427);
and U2370 (N_2370,In_386,In_700);
nand U2371 (N_2371,In_757,In_269);
nand U2372 (N_2372,In_716,In_40);
and U2373 (N_2373,In_571,In_469);
nand U2374 (N_2374,In_920,In_895);
nor U2375 (N_2375,In_504,In_847);
nor U2376 (N_2376,In_750,In_663);
and U2377 (N_2377,In_119,In_129);
nor U2378 (N_2378,In_893,In_486);
and U2379 (N_2379,In_609,In_99);
nor U2380 (N_2380,In_840,In_473);
or U2381 (N_2381,In_563,In_561);
or U2382 (N_2382,In_190,In_982);
and U2383 (N_2383,In_859,In_880);
nand U2384 (N_2384,In_978,In_931);
nand U2385 (N_2385,In_289,In_528);
nor U2386 (N_2386,In_5,In_152);
nor U2387 (N_2387,In_67,In_478);
nand U2388 (N_2388,In_219,In_831);
and U2389 (N_2389,In_300,In_783);
and U2390 (N_2390,In_561,In_178);
nor U2391 (N_2391,In_336,In_930);
nor U2392 (N_2392,In_624,In_756);
or U2393 (N_2393,In_416,In_683);
nor U2394 (N_2394,In_560,In_502);
or U2395 (N_2395,In_719,In_345);
and U2396 (N_2396,In_166,In_338);
nand U2397 (N_2397,In_459,In_960);
or U2398 (N_2398,In_187,In_139);
nand U2399 (N_2399,In_686,In_96);
and U2400 (N_2400,In_864,In_486);
nor U2401 (N_2401,In_592,In_46);
nand U2402 (N_2402,In_194,In_437);
nor U2403 (N_2403,In_167,In_881);
and U2404 (N_2404,In_881,In_215);
and U2405 (N_2405,In_70,In_58);
nor U2406 (N_2406,In_227,In_251);
and U2407 (N_2407,In_970,In_653);
or U2408 (N_2408,In_881,In_559);
nor U2409 (N_2409,In_906,In_357);
or U2410 (N_2410,In_655,In_802);
nor U2411 (N_2411,In_505,In_294);
nor U2412 (N_2412,In_369,In_647);
nand U2413 (N_2413,In_874,In_869);
nand U2414 (N_2414,In_0,In_699);
or U2415 (N_2415,In_600,In_590);
and U2416 (N_2416,In_373,In_124);
or U2417 (N_2417,In_868,In_111);
and U2418 (N_2418,In_544,In_949);
or U2419 (N_2419,In_542,In_983);
and U2420 (N_2420,In_303,In_291);
xor U2421 (N_2421,In_126,In_465);
nand U2422 (N_2422,In_118,In_641);
or U2423 (N_2423,In_128,In_711);
nand U2424 (N_2424,In_669,In_317);
or U2425 (N_2425,In_501,In_811);
nor U2426 (N_2426,In_947,In_18);
or U2427 (N_2427,In_6,In_358);
nand U2428 (N_2428,In_344,In_735);
or U2429 (N_2429,In_605,In_120);
or U2430 (N_2430,In_629,In_572);
nor U2431 (N_2431,In_112,In_444);
or U2432 (N_2432,In_78,In_293);
or U2433 (N_2433,In_139,In_245);
or U2434 (N_2434,In_846,In_935);
or U2435 (N_2435,In_753,In_606);
and U2436 (N_2436,In_551,In_69);
and U2437 (N_2437,In_477,In_634);
nor U2438 (N_2438,In_816,In_922);
nor U2439 (N_2439,In_850,In_167);
and U2440 (N_2440,In_165,In_879);
nand U2441 (N_2441,In_755,In_52);
nand U2442 (N_2442,In_812,In_155);
or U2443 (N_2443,In_558,In_910);
or U2444 (N_2444,In_277,In_75);
nand U2445 (N_2445,In_690,In_914);
nor U2446 (N_2446,In_170,In_842);
xor U2447 (N_2447,In_926,In_913);
or U2448 (N_2448,In_564,In_573);
or U2449 (N_2449,In_370,In_80);
nor U2450 (N_2450,In_394,In_209);
nor U2451 (N_2451,In_431,In_641);
or U2452 (N_2452,In_977,In_990);
or U2453 (N_2453,In_700,In_326);
and U2454 (N_2454,In_595,In_733);
or U2455 (N_2455,In_629,In_363);
or U2456 (N_2456,In_955,In_638);
or U2457 (N_2457,In_355,In_231);
and U2458 (N_2458,In_322,In_94);
nand U2459 (N_2459,In_256,In_480);
nor U2460 (N_2460,In_263,In_946);
nor U2461 (N_2461,In_869,In_161);
nor U2462 (N_2462,In_855,In_162);
and U2463 (N_2463,In_683,In_813);
nand U2464 (N_2464,In_377,In_828);
nand U2465 (N_2465,In_141,In_382);
nor U2466 (N_2466,In_41,In_678);
and U2467 (N_2467,In_884,In_282);
nand U2468 (N_2468,In_764,In_938);
nand U2469 (N_2469,In_107,In_200);
or U2470 (N_2470,In_438,In_945);
nand U2471 (N_2471,In_602,In_227);
or U2472 (N_2472,In_383,In_685);
and U2473 (N_2473,In_360,In_524);
nand U2474 (N_2474,In_925,In_417);
and U2475 (N_2475,In_28,In_737);
or U2476 (N_2476,In_633,In_751);
nand U2477 (N_2477,In_759,In_142);
and U2478 (N_2478,In_820,In_905);
and U2479 (N_2479,In_247,In_689);
nor U2480 (N_2480,In_0,In_754);
nor U2481 (N_2481,In_767,In_534);
nor U2482 (N_2482,In_141,In_290);
nand U2483 (N_2483,In_645,In_618);
nor U2484 (N_2484,In_409,In_781);
and U2485 (N_2485,In_684,In_497);
and U2486 (N_2486,In_955,In_460);
or U2487 (N_2487,In_117,In_714);
or U2488 (N_2488,In_970,In_536);
and U2489 (N_2489,In_236,In_150);
nor U2490 (N_2490,In_416,In_314);
nand U2491 (N_2491,In_307,In_725);
and U2492 (N_2492,In_462,In_25);
nand U2493 (N_2493,In_397,In_725);
or U2494 (N_2494,In_973,In_114);
and U2495 (N_2495,In_791,In_234);
and U2496 (N_2496,In_454,In_494);
nor U2497 (N_2497,In_285,In_804);
nor U2498 (N_2498,In_72,In_1);
and U2499 (N_2499,In_348,In_151);
and U2500 (N_2500,In_867,In_179);
nand U2501 (N_2501,In_673,In_780);
nand U2502 (N_2502,In_429,In_298);
nand U2503 (N_2503,In_545,In_656);
nor U2504 (N_2504,In_444,In_217);
or U2505 (N_2505,In_717,In_385);
or U2506 (N_2506,In_6,In_782);
or U2507 (N_2507,In_835,In_679);
nand U2508 (N_2508,In_877,In_651);
or U2509 (N_2509,In_597,In_403);
nand U2510 (N_2510,In_949,In_809);
nand U2511 (N_2511,In_544,In_86);
or U2512 (N_2512,In_251,In_643);
and U2513 (N_2513,In_107,In_794);
or U2514 (N_2514,In_487,In_868);
nand U2515 (N_2515,In_497,In_193);
nand U2516 (N_2516,In_439,In_276);
nand U2517 (N_2517,In_936,In_405);
or U2518 (N_2518,In_853,In_974);
nand U2519 (N_2519,In_22,In_530);
nor U2520 (N_2520,In_450,In_690);
nor U2521 (N_2521,In_222,In_14);
nor U2522 (N_2522,In_782,In_49);
and U2523 (N_2523,In_359,In_256);
nand U2524 (N_2524,In_953,In_774);
or U2525 (N_2525,In_435,In_241);
nor U2526 (N_2526,In_358,In_81);
or U2527 (N_2527,In_597,In_158);
nand U2528 (N_2528,In_735,In_443);
and U2529 (N_2529,In_481,In_442);
or U2530 (N_2530,In_3,In_172);
nand U2531 (N_2531,In_524,In_495);
nor U2532 (N_2532,In_93,In_989);
and U2533 (N_2533,In_310,In_118);
nand U2534 (N_2534,In_880,In_555);
nor U2535 (N_2535,In_144,In_314);
nor U2536 (N_2536,In_326,In_634);
and U2537 (N_2537,In_798,In_378);
and U2538 (N_2538,In_213,In_551);
or U2539 (N_2539,In_877,In_803);
and U2540 (N_2540,In_351,In_462);
or U2541 (N_2541,In_222,In_337);
nor U2542 (N_2542,In_470,In_98);
xor U2543 (N_2543,In_323,In_254);
and U2544 (N_2544,In_569,In_272);
and U2545 (N_2545,In_470,In_196);
and U2546 (N_2546,In_568,In_254);
or U2547 (N_2547,In_227,In_664);
and U2548 (N_2548,In_603,In_98);
or U2549 (N_2549,In_503,In_400);
nand U2550 (N_2550,In_878,In_747);
nand U2551 (N_2551,In_716,In_298);
nor U2552 (N_2552,In_697,In_306);
and U2553 (N_2553,In_768,In_858);
or U2554 (N_2554,In_653,In_385);
or U2555 (N_2555,In_364,In_331);
nand U2556 (N_2556,In_57,In_827);
nand U2557 (N_2557,In_733,In_565);
or U2558 (N_2558,In_874,In_970);
and U2559 (N_2559,In_715,In_624);
and U2560 (N_2560,In_62,In_229);
and U2561 (N_2561,In_235,In_721);
nor U2562 (N_2562,In_686,In_221);
nor U2563 (N_2563,In_901,In_582);
or U2564 (N_2564,In_344,In_720);
nand U2565 (N_2565,In_461,In_935);
nor U2566 (N_2566,In_63,In_674);
or U2567 (N_2567,In_733,In_452);
or U2568 (N_2568,In_885,In_315);
nand U2569 (N_2569,In_834,In_663);
nand U2570 (N_2570,In_70,In_216);
and U2571 (N_2571,In_295,In_768);
or U2572 (N_2572,In_575,In_274);
nor U2573 (N_2573,In_913,In_98);
and U2574 (N_2574,In_621,In_459);
or U2575 (N_2575,In_78,In_745);
nor U2576 (N_2576,In_824,In_380);
and U2577 (N_2577,In_973,In_20);
and U2578 (N_2578,In_25,In_365);
nand U2579 (N_2579,In_510,In_956);
nand U2580 (N_2580,In_183,In_334);
nand U2581 (N_2581,In_228,In_151);
and U2582 (N_2582,In_558,In_687);
nor U2583 (N_2583,In_754,In_313);
nand U2584 (N_2584,In_530,In_579);
or U2585 (N_2585,In_802,In_99);
or U2586 (N_2586,In_975,In_922);
and U2587 (N_2587,In_105,In_519);
or U2588 (N_2588,In_467,In_910);
nor U2589 (N_2589,In_808,In_712);
or U2590 (N_2590,In_9,In_35);
or U2591 (N_2591,In_588,In_465);
nand U2592 (N_2592,In_237,In_703);
or U2593 (N_2593,In_271,In_106);
and U2594 (N_2594,In_50,In_157);
and U2595 (N_2595,In_66,In_364);
or U2596 (N_2596,In_392,In_10);
nand U2597 (N_2597,In_632,In_104);
nor U2598 (N_2598,In_330,In_195);
nand U2599 (N_2599,In_104,In_300);
and U2600 (N_2600,In_331,In_311);
or U2601 (N_2601,In_43,In_475);
or U2602 (N_2602,In_143,In_404);
and U2603 (N_2603,In_260,In_148);
and U2604 (N_2604,In_736,In_517);
nor U2605 (N_2605,In_367,In_103);
xnor U2606 (N_2606,In_495,In_980);
or U2607 (N_2607,In_884,In_378);
nor U2608 (N_2608,In_512,In_533);
nor U2609 (N_2609,In_600,In_64);
and U2610 (N_2610,In_263,In_724);
xnor U2611 (N_2611,In_425,In_826);
or U2612 (N_2612,In_214,In_116);
or U2613 (N_2613,In_621,In_394);
and U2614 (N_2614,In_624,In_950);
nor U2615 (N_2615,In_151,In_610);
nor U2616 (N_2616,In_162,In_461);
nor U2617 (N_2617,In_803,In_421);
and U2618 (N_2618,In_376,In_61);
or U2619 (N_2619,In_439,In_717);
and U2620 (N_2620,In_307,In_826);
nor U2621 (N_2621,In_456,In_473);
xnor U2622 (N_2622,In_141,In_616);
and U2623 (N_2623,In_851,In_158);
nor U2624 (N_2624,In_118,In_892);
nand U2625 (N_2625,In_515,In_917);
nand U2626 (N_2626,In_426,In_945);
and U2627 (N_2627,In_105,In_730);
nor U2628 (N_2628,In_639,In_309);
or U2629 (N_2629,In_720,In_797);
nor U2630 (N_2630,In_76,In_44);
or U2631 (N_2631,In_709,In_824);
nand U2632 (N_2632,In_863,In_876);
and U2633 (N_2633,In_161,In_915);
and U2634 (N_2634,In_402,In_259);
nor U2635 (N_2635,In_833,In_755);
xnor U2636 (N_2636,In_931,In_753);
or U2637 (N_2637,In_323,In_130);
and U2638 (N_2638,In_912,In_805);
nor U2639 (N_2639,In_68,In_725);
or U2640 (N_2640,In_797,In_929);
nand U2641 (N_2641,In_965,In_975);
nand U2642 (N_2642,In_772,In_995);
and U2643 (N_2643,In_149,In_752);
nand U2644 (N_2644,In_338,In_364);
and U2645 (N_2645,In_543,In_71);
or U2646 (N_2646,In_535,In_797);
and U2647 (N_2647,In_690,In_52);
and U2648 (N_2648,In_344,In_838);
nor U2649 (N_2649,In_704,In_271);
and U2650 (N_2650,In_634,In_216);
or U2651 (N_2651,In_250,In_970);
nand U2652 (N_2652,In_721,In_484);
or U2653 (N_2653,In_362,In_316);
nor U2654 (N_2654,In_824,In_70);
xnor U2655 (N_2655,In_209,In_988);
nand U2656 (N_2656,In_626,In_762);
and U2657 (N_2657,In_906,In_766);
nor U2658 (N_2658,In_9,In_526);
and U2659 (N_2659,In_646,In_52);
or U2660 (N_2660,In_377,In_415);
or U2661 (N_2661,In_732,In_871);
nand U2662 (N_2662,In_534,In_975);
nand U2663 (N_2663,In_776,In_323);
and U2664 (N_2664,In_322,In_539);
nor U2665 (N_2665,In_678,In_772);
and U2666 (N_2666,In_842,In_390);
nand U2667 (N_2667,In_427,In_581);
nand U2668 (N_2668,In_89,In_77);
nor U2669 (N_2669,In_701,In_666);
or U2670 (N_2670,In_325,In_244);
and U2671 (N_2671,In_588,In_792);
or U2672 (N_2672,In_964,In_483);
nor U2673 (N_2673,In_10,In_744);
and U2674 (N_2674,In_562,In_242);
nand U2675 (N_2675,In_893,In_984);
nor U2676 (N_2676,In_917,In_13);
and U2677 (N_2677,In_631,In_677);
nor U2678 (N_2678,In_714,In_77);
nor U2679 (N_2679,In_415,In_915);
or U2680 (N_2680,In_793,In_424);
nand U2681 (N_2681,In_223,In_183);
nor U2682 (N_2682,In_944,In_779);
or U2683 (N_2683,In_725,In_111);
nand U2684 (N_2684,In_245,In_929);
or U2685 (N_2685,In_574,In_420);
or U2686 (N_2686,In_895,In_561);
or U2687 (N_2687,In_989,In_629);
nor U2688 (N_2688,In_752,In_933);
nor U2689 (N_2689,In_232,In_541);
or U2690 (N_2690,In_643,In_184);
nor U2691 (N_2691,In_349,In_712);
or U2692 (N_2692,In_795,In_521);
and U2693 (N_2693,In_885,In_336);
nand U2694 (N_2694,In_252,In_793);
nand U2695 (N_2695,In_685,In_420);
and U2696 (N_2696,In_635,In_636);
and U2697 (N_2697,In_213,In_346);
nor U2698 (N_2698,In_576,In_418);
and U2699 (N_2699,In_785,In_685);
and U2700 (N_2700,In_941,In_919);
nor U2701 (N_2701,In_694,In_477);
nand U2702 (N_2702,In_68,In_961);
nor U2703 (N_2703,In_115,In_235);
nor U2704 (N_2704,In_37,In_305);
nor U2705 (N_2705,In_206,In_385);
nand U2706 (N_2706,In_76,In_187);
nor U2707 (N_2707,In_781,In_826);
and U2708 (N_2708,In_601,In_242);
nand U2709 (N_2709,In_921,In_790);
and U2710 (N_2710,In_953,In_580);
and U2711 (N_2711,In_210,In_549);
and U2712 (N_2712,In_365,In_394);
or U2713 (N_2713,In_508,In_314);
or U2714 (N_2714,In_44,In_839);
and U2715 (N_2715,In_462,In_904);
nor U2716 (N_2716,In_237,In_234);
and U2717 (N_2717,In_810,In_874);
and U2718 (N_2718,In_904,In_899);
and U2719 (N_2719,In_914,In_650);
and U2720 (N_2720,In_26,In_816);
nand U2721 (N_2721,In_636,In_10);
or U2722 (N_2722,In_745,In_245);
and U2723 (N_2723,In_566,In_463);
nor U2724 (N_2724,In_577,In_953);
and U2725 (N_2725,In_106,In_991);
nand U2726 (N_2726,In_688,In_770);
or U2727 (N_2727,In_541,In_767);
nor U2728 (N_2728,In_847,In_705);
xor U2729 (N_2729,In_680,In_68);
or U2730 (N_2730,In_740,In_550);
nor U2731 (N_2731,In_272,In_504);
nand U2732 (N_2732,In_221,In_128);
nor U2733 (N_2733,In_833,In_921);
or U2734 (N_2734,In_770,In_720);
nor U2735 (N_2735,In_423,In_264);
and U2736 (N_2736,In_163,In_701);
nand U2737 (N_2737,In_421,In_987);
nand U2738 (N_2738,In_861,In_634);
nor U2739 (N_2739,In_430,In_295);
nand U2740 (N_2740,In_430,In_692);
or U2741 (N_2741,In_456,In_646);
nand U2742 (N_2742,In_796,In_508);
nand U2743 (N_2743,In_585,In_815);
or U2744 (N_2744,In_233,In_621);
and U2745 (N_2745,In_584,In_420);
nand U2746 (N_2746,In_135,In_958);
nand U2747 (N_2747,In_156,In_56);
nor U2748 (N_2748,In_866,In_855);
nor U2749 (N_2749,In_340,In_359);
or U2750 (N_2750,In_292,In_992);
and U2751 (N_2751,In_216,In_631);
and U2752 (N_2752,In_684,In_937);
or U2753 (N_2753,In_994,In_127);
or U2754 (N_2754,In_85,In_51);
and U2755 (N_2755,In_928,In_412);
and U2756 (N_2756,In_270,In_953);
nor U2757 (N_2757,In_668,In_799);
and U2758 (N_2758,In_602,In_488);
nand U2759 (N_2759,In_935,In_423);
and U2760 (N_2760,In_575,In_179);
nand U2761 (N_2761,In_515,In_166);
nor U2762 (N_2762,In_966,In_545);
or U2763 (N_2763,In_737,In_955);
nor U2764 (N_2764,In_635,In_709);
nand U2765 (N_2765,In_803,In_351);
nand U2766 (N_2766,In_714,In_272);
nor U2767 (N_2767,In_685,In_832);
nand U2768 (N_2768,In_882,In_881);
and U2769 (N_2769,In_494,In_545);
or U2770 (N_2770,In_502,In_214);
and U2771 (N_2771,In_332,In_318);
and U2772 (N_2772,In_245,In_99);
nor U2773 (N_2773,In_637,In_84);
nor U2774 (N_2774,In_381,In_212);
and U2775 (N_2775,In_129,In_393);
nor U2776 (N_2776,In_560,In_639);
and U2777 (N_2777,In_839,In_945);
nor U2778 (N_2778,In_512,In_520);
and U2779 (N_2779,In_408,In_435);
and U2780 (N_2780,In_8,In_346);
or U2781 (N_2781,In_387,In_426);
nand U2782 (N_2782,In_155,In_388);
nor U2783 (N_2783,In_869,In_18);
nand U2784 (N_2784,In_760,In_302);
and U2785 (N_2785,In_78,In_60);
or U2786 (N_2786,In_905,In_391);
nand U2787 (N_2787,In_824,In_71);
nor U2788 (N_2788,In_83,In_475);
nand U2789 (N_2789,In_856,In_678);
nand U2790 (N_2790,In_882,In_933);
or U2791 (N_2791,In_705,In_400);
or U2792 (N_2792,In_565,In_968);
nand U2793 (N_2793,In_80,In_369);
or U2794 (N_2794,In_698,In_275);
or U2795 (N_2795,In_199,In_742);
nand U2796 (N_2796,In_726,In_268);
nand U2797 (N_2797,In_182,In_301);
or U2798 (N_2798,In_150,In_872);
nand U2799 (N_2799,In_640,In_975);
nand U2800 (N_2800,In_987,In_427);
and U2801 (N_2801,In_899,In_155);
nand U2802 (N_2802,In_856,In_322);
nand U2803 (N_2803,In_384,In_95);
nor U2804 (N_2804,In_805,In_468);
nor U2805 (N_2805,In_911,In_523);
or U2806 (N_2806,In_944,In_464);
nand U2807 (N_2807,In_741,In_504);
nand U2808 (N_2808,In_426,In_771);
nand U2809 (N_2809,In_313,In_715);
or U2810 (N_2810,In_153,In_11);
nand U2811 (N_2811,In_198,In_241);
and U2812 (N_2812,In_850,In_706);
or U2813 (N_2813,In_551,In_544);
nand U2814 (N_2814,In_744,In_512);
xnor U2815 (N_2815,In_979,In_935);
nor U2816 (N_2816,In_163,In_266);
or U2817 (N_2817,In_388,In_754);
and U2818 (N_2818,In_319,In_811);
or U2819 (N_2819,In_847,In_740);
nand U2820 (N_2820,In_882,In_752);
and U2821 (N_2821,In_882,In_678);
or U2822 (N_2822,In_77,In_897);
nand U2823 (N_2823,In_320,In_602);
nor U2824 (N_2824,In_953,In_573);
or U2825 (N_2825,In_205,In_393);
nand U2826 (N_2826,In_348,In_961);
nor U2827 (N_2827,In_457,In_150);
nand U2828 (N_2828,In_89,In_147);
nor U2829 (N_2829,In_79,In_199);
and U2830 (N_2830,In_266,In_358);
or U2831 (N_2831,In_839,In_971);
nand U2832 (N_2832,In_784,In_214);
nand U2833 (N_2833,In_280,In_537);
nand U2834 (N_2834,In_101,In_77);
or U2835 (N_2835,In_741,In_610);
or U2836 (N_2836,In_522,In_248);
and U2837 (N_2837,In_193,In_224);
or U2838 (N_2838,In_957,In_143);
or U2839 (N_2839,In_21,In_826);
nand U2840 (N_2840,In_361,In_135);
nand U2841 (N_2841,In_974,In_799);
and U2842 (N_2842,In_110,In_603);
and U2843 (N_2843,In_796,In_537);
and U2844 (N_2844,In_27,In_580);
and U2845 (N_2845,In_880,In_444);
or U2846 (N_2846,In_415,In_668);
nor U2847 (N_2847,In_352,In_254);
and U2848 (N_2848,In_496,In_333);
nand U2849 (N_2849,In_150,In_417);
nor U2850 (N_2850,In_53,In_561);
and U2851 (N_2851,In_851,In_685);
or U2852 (N_2852,In_535,In_757);
nor U2853 (N_2853,In_951,In_423);
nor U2854 (N_2854,In_27,In_862);
xnor U2855 (N_2855,In_531,In_172);
nand U2856 (N_2856,In_935,In_73);
nand U2857 (N_2857,In_303,In_882);
nand U2858 (N_2858,In_991,In_66);
nor U2859 (N_2859,In_131,In_901);
nand U2860 (N_2860,In_147,In_77);
and U2861 (N_2861,In_655,In_813);
nand U2862 (N_2862,In_17,In_624);
nor U2863 (N_2863,In_542,In_596);
or U2864 (N_2864,In_29,In_396);
or U2865 (N_2865,In_700,In_423);
and U2866 (N_2866,In_405,In_47);
and U2867 (N_2867,In_990,In_23);
and U2868 (N_2868,In_23,In_36);
and U2869 (N_2869,In_983,In_115);
nor U2870 (N_2870,In_643,In_576);
nand U2871 (N_2871,In_794,In_174);
nor U2872 (N_2872,In_859,In_844);
or U2873 (N_2873,In_244,In_851);
nand U2874 (N_2874,In_278,In_272);
and U2875 (N_2875,In_600,In_319);
nand U2876 (N_2876,In_507,In_244);
or U2877 (N_2877,In_155,In_665);
and U2878 (N_2878,In_97,In_332);
nand U2879 (N_2879,In_814,In_122);
or U2880 (N_2880,In_502,In_219);
or U2881 (N_2881,In_330,In_249);
nor U2882 (N_2882,In_278,In_122);
or U2883 (N_2883,In_658,In_365);
nor U2884 (N_2884,In_917,In_510);
nor U2885 (N_2885,In_803,In_679);
nor U2886 (N_2886,In_936,In_390);
and U2887 (N_2887,In_848,In_499);
nand U2888 (N_2888,In_83,In_869);
and U2889 (N_2889,In_665,In_329);
or U2890 (N_2890,In_313,In_199);
nor U2891 (N_2891,In_488,In_310);
nand U2892 (N_2892,In_679,In_612);
or U2893 (N_2893,In_450,In_230);
nand U2894 (N_2894,In_895,In_676);
nor U2895 (N_2895,In_841,In_863);
nand U2896 (N_2896,In_876,In_868);
or U2897 (N_2897,In_693,In_53);
and U2898 (N_2898,In_742,In_192);
xnor U2899 (N_2899,In_650,In_490);
and U2900 (N_2900,In_686,In_239);
and U2901 (N_2901,In_194,In_494);
or U2902 (N_2902,In_584,In_400);
or U2903 (N_2903,In_63,In_294);
and U2904 (N_2904,In_846,In_243);
nor U2905 (N_2905,In_633,In_754);
nand U2906 (N_2906,In_801,In_858);
and U2907 (N_2907,In_561,In_251);
nand U2908 (N_2908,In_271,In_11);
and U2909 (N_2909,In_717,In_406);
and U2910 (N_2910,In_193,In_886);
nor U2911 (N_2911,In_743,In_540);
or U2912 (N_2912,In_84,In_630);
or U2913 (N_2913,In_170,In_599);
and U2914 (N_2914,In_995,In_356);
nand U2915 (N_2915,In_980,In_664);
nor U2916 (N_2916,In_778,In_994);
or U2917 (N_2917,In_30,In_738);
nand U2918 (N_2918,In_964,In_271);
nand U2919 (N_2919,In_663,In_159);
nand U2920 (N_2920,In_478,In_36);
nor U2921 (N_2921,In_238,In_391);
and U2922 (N_2922,In_817,In_369);
and U2923 (N_2923,In_184,In_959);
nor U2924 (N_2924,In_159,In_491);
and U2925 (N_2925,In_717,In_831);
nor U2926 (N_2926,In_433,In_504);
and U2927 (N_2927,In_330,In_960);
and U2928 (N_2928,In_79,In_372);
nor U2929 (N_2929,In_570,In_116);
nand U2930 (N_2930,In_904,In_369);
or U2931 (N_2931,In_773,In_197);
or U2932 (N_2932,In_423,In_511);
and U2933 (N_2933,In_210,In_614);
nor U2934 (N_2934,In_129,In_212);
nand U2935 (N_2935,In_561,In_702);
and U2936 (N_2936,In_279,In_664);
nand U2937 (N_2937,In_738,In_491);
nor U2938 (N_2938,In_884,In_738);
nor U2939 (N_2939,In_508,In_132);
nor U2940 (N_2940,In_510,In_103);
nand U2941 (N_2941,In_380,In_43);
nor U2942 (N_2942,In_790,In_192);
and U2943 (N_2943,In_147,In_954);
nand U2944 (N_2944,In_597,In_222);
nand U2945 (N_2945,In_285,In_474);
nor U2946 (N_2946,In_745,In_352);
and U2947 (N_2947,In_66,In_597);
nand U2948 (N_2948,In_734,In_742);
nand U2949 (N_2949,In_626,In_731);
nor U2950 (N_2950,In_102,In_662);
and U2951 (N_2951,In_531,In_953);
nor U2952 (N_2952,In_759,In_736);
nand U2953 (N_2953,In_589,In_174);
or U2954 (N_2954,In_861,In_688);
and U2955 (N_2955,In_892,In_657);
or U2956 (N_2956,In_14,In_977);
nand U2957 (N_2957,In_403,In_499);
nand U2958 (N_2958,In_870,In_222);
nor U2959 (N_2959,In_916,In_231);
and U2960 (N_2960,In_636,In_258);
nor U2961 (N_2961,In_950,In_336);
and U2962 (N_2962,In_958,In_546);
nor U2963 (N_2963,In_967,In_401);
nor U2964 (N_2964,In_457,In_108);
and U2965 (N_2965,In_427,In_261);
or U2966 (N_2966,In_540,In_823);
or U2967 (N_2967,In_866,In_882);
and U2968 (N_2968,In_146,In_355);
and U2969 (N_2969,In_879,In_690);
nor U2970 (N_2970,In_356,In_945);
and U2971 (N_2971,In_202,In_775);
nand U2972 (N_2972,In_442,In_193);
and U2973 (N_2973,In_571,In_725);
and U2974 (N_2974,In_534,In_168);
nand U2975 (N_2975,In_182,In_531);
and U2976 (N_2976,In_504,In_373);
nor U2977 (N_2977,In_836,In_200);
nand U2978 (N_2978,In_101,In_21);
and U2979 (N_2979,In_21,In_158);
nand U2980 (N_2980,In_205,In_806);
or U2981 (N_2981,In_941,In_240);
nor U2982 (N_2982,In_48,In_140);
and U2983 (N_2983,In_553,In_546);
and U2984 (N_2984,In_797,In_396);
and U2985 (N_2985,In_875,In_891);
nor U2986 (N_2986,In_155,In_882);
nor U2987 (N_2987,In_793,In_601);
and U2988 (N_2988,In_733,In_743);
and U2989 (N_2989,In_610,In_966);
and U2990 (N_2990,In_795,In_840);
or U2991 (N_2991,In_172,In_828);
or U2992 (N_2992,In_424,In_650);
nand U2993 (N_2993,In_51,In_336);
nor U2994 (N_2994,In_145,In_705);
and U2995 (N_2995,In_865,In_914);
or U2996 (N_2996,In_959,In_986);
nand U2997 (N_2997,In_200,In_326);
nor U2998 (N_2998,In_736,In_243);
and U2999 (N_2999,In_678,In_636);
nor U3000 (N_3000,In_13,In_71);
and U3001 (N_3001,In_513,In_627);
nand U3002 (N_3002,In_340,In_634);
and U3003 (N_3003,In_386,In_302);
and U3004 (N_3004,In_933,In_782);
and U3005 (N_3005,In_38,In_599);
or U3006 (N_3006,In_511,In_49);
nand U3007 (N_3007,In_124,In_247);
nand U3008 (N_3008,In_876,In_481);
nand U3009 (N_3009,In_296,In_357);
nor U3010 (N_3010,In_221,In_950);
and U3011 (N_3011,In_861,In_568);
and U3012 (N_3012,In_855,In_179);
nor U3013 (N_3013,In_106,In_979);
or U3014 (N_3014,In_737,In_120);
xnor U3015 (N_3015,In_431,In_74);
nor U3016 (N_3016,In_730,In_718);
and U3017 (N_3017,In_978,In_103);
and U3018 (N_3018,In_487,In_220);
and U3019 (N_3019,In_641,In_114);
and U3020 (N_3020,In_730,In_158);
nor U3021 (N_3021,In_81,In_397);
nand U3022 (N_3022,In_323,In_548);
nand U3023 (N_3023,In_361,In_392);
nor U3024 (N_3024,In_957,In_801);
and U3025 (N_3025,In_765,In_211);
or U3026 (N_3026,In_177,In_929);
or U3027 (N_3027,In_826,In_829);
nand U3028 (N_3028,In_185,In_201);
or U3029 (N_3029,In_274,In_985);
nor U3030 (N_3030,In_96,In_210);
or U3031 (N_3031,In_152,In_50);
or U3032 (N_3032,In_18,In_173);
or U3033 (N_3033,In_464,In_381);
and U3034 (N_3034,In_459,In_82);
nand U3035 (N_3035,In_856,In_694);
or U3036 (N_3036,In_340,In_141);
nand U3037 (N_3037,In_425,In_575);
nor U3038 (N_3038,In_275,In_999);
or U3039 (N_3039,In_180,In_731);
nor U3040 (N_3040,In_602,In_848);
or U3041 (N_3041,In_469,In_776);
and U3042 (N_3042,In_420,In_520);
and U3043 (N_3043,In_124,In_411);
nand U3044 (N_3044,In_447,In_973);
nor U3045 (N_3045,In_491,In_300);
nor U3046 (N_3046,In_368,In_559);
nor U3047 (N_3047,In_78,In_423);
and U3048 (N_3048,In_636,In_395);
or U3049 (N_3049,In_142,In_982);
nand U3050 (N_3050,In_910,In_41);
or U3051 (N_3051,In_708,In_209);
or U3052 (N_3052,In_942,In_869);
nor U3053 (N_3053,In_970,In_552);
nor U3054 (N_3054,In_481,In_248);
or U3055 (N_3055,In_107,In_655);
nand U3056 (N_3056,In_987,In_588);
and U3057 (N_3057,In_520,In_829);
and U3058 (N_3058,In_869,In_332);
and U3059 (N_3059,In_402,In_589);
or U3060 (N_3060,In_370,In_856);
nor U3061 (N_3061,In_469,In_555);
nor U3062 (N_3062,In_118,In_99);
nand U3063 (N_3063,In_666,In_694);
nand U3064 (N_3064,In_557,In_914);
nand U3065 (N_3065,In_37,In_588);
nand U3066 (N_3066,In_794,In_939);
or U3067 (N_3067,In_12,In_718);
or U3068 (N_3068,In_13,In_618);
nand U3069 (N_3069,In_970,In_5);
nand U3070 (N_3070,In_86,In_101);
nand U3071 (N_3071,In_67,In_166);
or U3072 (N_3072,In_927,In_755);
or U3073 (N_3073,In_65,In_468);
nand U3074 (N_3074,In_429,In_731);
nand U3075 (N_3075,In_179,In_977);
nand U3076 (N_3076,In_307,In_589);
nor U3077 (N_3077,In_590,In_813);
or U3078 (N_3078,In_204,In_189);
nor U3079 (N_3079,In_294,In_448);
nor U3080 (N_3080,In_575,In_419);
xor U3081 (N_3081,In_760,In_106);
and U3082 (N_3082,In_32,In_980);
nor U3083 (N_3083,In_507,In_570);
nor U3084 (N_3084,In_498,In_973);
nand U3085 (N_3085,In_829,In_142);
nand U3086 (N_3086,In_820,In_423);
nand U3087 (N_3087,In_419,In_734);
nor U3088 (N_3088,In_739,In_758);
or U3089 (N_3089,In_249,In_411);
nand U3090 (N_3090,In_814,In_242);
nand U3091 (N_3091,In_478,In_426);
or U3092 (N_3092,In_256,In_745);
or U3093 (N_3093,In_354,In_901);
nor U3094 (N_3094,In_207,In_307);
or U3095 (N_3095,In_554,In_133);
nand U3096 (N_3096,In_200,In_39);
nor U3097 (N_3097,In_982,In_782);
and U3098 (N_3098,In_218,In_338);
or U3099 (N_3099,In_92,In_610);
and U3100 (N_3100,In_966,In_190);
nor U3101 (N_3101,In_772,In_313);
nand U3102 (N_3102,In_704,In_233);
and U3103 (N_3103,In_152,In_734);
nand U3104 (N_3104,In_141,In_922);
and U3105 (N_3105,In_842,In_345);
nor U3106 (N_3106,In_542,In_787);
nand U3107 (N_3107,In_942,In_200);
and U3108 (N_3108,In_495,In_4);
and U3109 (N_3109,In_496,In_306);
nand U3110 (N_3110,In_317,In_894);
nor U3111 (N_3111,In_44,In_247);
or U3112 (N_3112,In_822,In_751);
nand U3113 (N_3113,In_837,In_391);
or U3114 (N_3114,In_782,In_292);
and U3115 (N_3115,In_547,In_741);
nor U3116 (N_3116,In_905,In_227);
or U3117 (N_3117,In_831,In_129);
nor U3118 (N_3118,In_56,In_772);
nand U3119 (N_3119,In_390,In_43);
nand U3120 (N_3120,In_330,In_997);
or U3121 (N_3121,In_594,In_465);
or U3122 (N_3122,In_858,In_516);
and U3123 (N_3123,In_541,In_302);
or U3124 (N_3124,In_976,In_967);
and U3125 (N_3125,In_766,In_228);
nand U3126 (N_3126,In_419,In_814);
nand U3127 (N_3127,In_792,In_513);
or U3128 (N_3128,In_432,In_228);
and U3129 (N_3129,In_928,In_373);
or U3130 (N_3130,In_47,In_688);
or U3131 (N_3131,In_942,In_11);
nor U3132 (N_3132,In_829,In_559);
nor U3133 (N_3133,In_182,In_218);
nand U3134 (N_3134,In_778,In_3);
nor U3135 (N_3135,In_446,In_21);
or U3136 (N_3136,In_88,In_898);
nand U3137 (N_3137,In_897,In_255);
xor U3138 (N_3138,In_369,In_582);
and U3139 (N_3139,In_182,In_590);
xnor U3140 (N_3140,In_105,In_241);
or U3141 (N_3141,In_900,In_140);
nand U3142 (N_3142,In_369,In_555);
nand U3143 (N_3143,In_469,In_90);
and U3144 (N_3144,In_609,In_40);
nor U3145 (N_3145,In_692,In_301);
nand U3146 (N_3146,In_765,In_981);
nor U3147 (N_3147,In_485,In_102);
nor U3148 (N_3148,In_271,In_452);
nor U3149 (N_3149,In_107,In_737);
nand U3150 (N_3150,In_857,In_322);
nand U3151 (N_3151,In_2,In_604);
or U3152 (N_3152,In_972,In_597);
and U3153 (N_3153,In_833,In_914);
nor U3154 (N_3154,In_166,In_395);
or U3155 (N_3155,In_860,In_218);
or U3156 (N_3156,In_154,In_507);
and U3157 (N_3157,In_259,In_995);
or U3158 (N_3158,In_465,In_740);
nor U3159 (N_3159,In_310,In_6);
or U3160 (N_3160,In_291,In_59);
and U3161 (N_3161,In_275,In_519);
nor U3162 (N_3162,In_899,In_303);
nor U3163 (N_3163,In_427,In_229);
nor U3164 (N_3164,In_957,In_391);
and U3165 (N_3165,In_498,In_804);
nand U3166 (N_3166,In_123,In_664);
nor U3167 (N_3167,In_568,In_569);
nand U3168 (N_3168,In_645,In_63);
nand U3169 (N_3169,In_769,In_877);
or U3170 (N_3170,In_2,In_239);
or U3171 (N_3171,In_794,In_897);
or U3172 (N_3172,In_910,In_261);
and U3173 (N_3173,In_55,In_19);
and U3174 (N_3174,In_843,In_685);
or U3175 (N_3175,In_126,In_811);
and U3176 (N_3176,In_911,In_320);
and U3177 (N_3177,In_661,In_176);
nor U3178 (N_3178,In_708,In_766);
or U3179 (N_3179,In_734,In_105);
nand U3180 (N_3180,In_213,In_954);
nor U3181 (N_3181,In_323,In_802);
nand U3182 (N_3182,In_753,In_767);
nor U3183 (N_3183,In_815,In_237);
nor U3184 (N_3184,In_850,In_77);
nand U3185 (N_3185,In_324,In_728);
and U3186 (N_3186,In_289,In_696);
nor U3187 (N_3187,In_609,In_170);
or U3188 (N_3188,In_544,In_868);
nand U3189 (N_3189,In_262,In_969);
nand U3190 (N_3190,In_980,In_725);
nand U3191 (N_3191,In_83,In_829);
nand U3192 (N_3192,In_882,In_222);
nand U3193 (N_3193,In_400,In_110);
or U3194 (N_3194,In_712,In_595);
or U3195 (N_3195,In_617,In_460);
or U3196 (N_3196,In_653,In_687);
and U3197 (N_3197,In_231,In_979);
and U3198 (N_3198,In_914,In_37);
and U3199 (N_3199,In_904,In_764);
and U3200 (N_3200,In_457,In_369);
and U3201 (N_3201,In_148,In_934);
nand U3202 (N_3202,In_771,In_395);
nand U3203 (N_3203,In_657,In_582);
nor U3204 (N_3204,In_958,In_592);
and U3205 (N_3205,In_903,In_639);
or U3206 (N_3206,In_332,In_791);
or U3207 (N_3207,In_563,In_612);
nand U3208 (N_3208,In_482,In_72);
or U3209 (N_3209,In_225,In_576);
nand U3210 (N_3210,In_298,In_155);
nor U3211 (N_3211,In_22,In_37);
or U3212 (N_3212,In_147,In_312);
nor U3213 (N_3213,In_276,In_628);
nand U3214 (N_3214,In_235,In_765);
nor U3215 (N_3215,In_773,In_407);
nor U3216 (N_3216,In_678,In_419);
and U3217 (N_3217,In_518,In_615);
or U3218 (N_3218,In_5,In_653);
and U3219 (N_3219,In_646,In_531);
and U3220 (N_3220,In_557,In_946);
nand U3221 (N_3221,In_365,In_614);
and U3222 (N_3222,In_316,In_143);
nand U3223 (N_3223,In_65,In_315);
or U3224 (N_3224,In_93,In_645);
nand U3225 (N_3225,In_507,In_435);
and U3226 (N_3226,In_642,In_550);
nor U3227 (N_3227,In_875,In_141);
or U3228 (N_3228,In_841,In_21);
nor U3229 (N_3229,In_921,In_425);
and U3230 (N_3230,In_313,In_430);
nor U3231 (N_3231,In_455,In_33);
nor U3232 (N_3232,In_998,In_720);
nor U3233 (N_3233,In_548,In_142);
nor U3234 (N_3234,In_900,In_264);
or U3235 (N_3235,In_5,In_26);
nor U3236 (N_3236,In_649,In_8);
or U3237 (N_3237,In_119,In_621);
or U3238 (N_3238,In_183,In_656);
and U3239 (N_3239,In_604,In_435);
nor U3240 (N_3240,In_146,In_329);
nor U3241 (N_3241,In_609,In_112);
nor U3242 (N_3242,In_254,In_617);
or U3243 (N_3243,In_264,In_412);
nand U3244 (N_3244,In_93,In_974);
and U3245 (N_3245,In_299,In_765);
xnor U3246 (N_3246,In_735,In_475);
nor U3247 (N_3247,In_908,In_569);
and U3248 (N_3248,In_504,In_453);
or U3249 (N_3249,In_317,In_78);
nand U3250 (N_3250,In_535,In_126);
and U3251 (N_3251,In_201,In_116);
nor U3252 (N_3252,In_959,In_660);
nor U3253 (N_3253,In_661,In_331);
or U3254 (N_3254,In_345,In_380);
or U3255 (N_3255,In_347,In_744);
or U3256 (N_3256,In_23,In_523);
nand U3257 (N_3257,In_384,In_2);
nand U3258 (N_3258,In_925,In_197);
nor U3259 (N_3259,In_624,In_498);
nor U3260 (N_3260,In_485,In_783);
nor U3261 (N_3261,In_513,In_447);
nor U3262 (N_3262,In_521,In_826);
nor U3263 (N_3263,In_911,In_640);
nand U3264 (N_3264,In_939,In_542);
and U3265 (N_3265,In_491,In_75);
and U3266 (N_3266,In_207,In_417);
nand U3267 (N_3267,In_509,In_591);
and U3268 (N_3268,In_339,In_408);
nor U3269 (N_3269,In_159,In_152);
or U3270 (N_3270,In_223,In_206);
nor U3271 (N_3271,In_377,In_987);
and U3272 (N_3272,In_384,In_123);
or U3273 (N_3273,In_925,In_80);
nand U3274 (N_3274,In_191,In_285);
and U3275 (N_3275,In_849,In_92);
nor U3276 (N_3276,In_194,In_709);
or U3277 (N_3277,In_697,In_634);
nand U3278 (N_3278,In_586,In_73);
nand U3279 (N_3279,In_754,In_714);
or U3280 (N_3280,In_896,In_66);
nand U3281 (N_3281,In_896,In_933);
or U3282 (N_3282,In_314,In_30);
nor U3283 (N_3283,In_688,In_60);
and U3284 (N_3284,In_851,In_254);
or U3285 (N_3285,In_84,In_629);
or U3286 (N_3286,In_194,In_377);
nor U3287 (N_3287,In_367,In_526);
or U3288 (N_3288,In_132,In_99);
nor U3289 (N_3289,In_551,In_467);
or U3290 (N_3290,In_461,In_670);
and U3291 (N_3291,In_345,In_230);
nand U3292 (N_3292,In_750,In_956);
or U3293 (N_3293,In_551,In_65);
nor U3294 (N_3294,In_221,In_422);
nand U3295 (N_3295,In_517,In_823);
or U3296 (N_3296,In_701,In_891);
nor U3297 (N_3297,In_38,In_809);
nand U3298 (N_3298,In_461,In_950);
or U3299 (N_3299,In_933,In_349);
and U3300 (N_3300,In_648,In_664);
nand U3301 (N_3301,In_320,In_831);
or U3302 (N_3302,In_434,In_382);
nor U3303 (N_3303,In_354,In_158);
nor U3304 (N_3304,In_198,In_517);
nand U3305 (N_3305,In_672,In_380);
nand U3306 (N_3306,In_530,In_268);
nand U3307 (N_3307,In_688,In_628);
or U3308 (N_3308,In_524,In_338);
nor U3309 (N_3309,In_79,In_987);
or U3310 (N_3310,In_862,In_713);
or U3311 (N_3311,In_166,In_312);
or U3312 (N_3312,In_799,In_435);
and U3313 (N_3313,In_641,In_182);
nor U3314 (N_3314,In_678,In_151);
or U3315 (N_3315,In_24,In_116);
and U3316 (N_3316,In_117,In_376);
or U3317 (N_3317,In_170,In_151);
nor U3318 (N_3318,In_731,In_777);
or U3319 (N_3319,In_467,In_12);
nor U3320 (N_3320,In_266,In_917);
and U3321 (N_3321,In_495,In_152);
and U3322 (N_3322,In_505,In_238);
nand U3323 (N_3323,In_751,In_824);
nand U3324 (N_3324,In_556,In_429);
or U3325 (N_3325,In_656,In_343);
nor U3326 (N_3326,In_620,In_878);
nor U3327 (N_3327,In_775,In_227);
and U3328 (N_3328,In_636,In_312);
nand U3329 (N_3329,In_970,In_312);
xor U3330 (N_3330,In_769,In_402);
and U3331 (N_3331,In_80,In_806);
or U3332 (N_3332,In_785,In_458);
nand U3333 (N_3333,In_742,In_488);
nor U3334 (N_3334,In_486,In_40);
or U3335 (N_3335,In_105,In_869);
nand U3336 (N_3336,In_39,In_543);
or U3337 (N_3337,In_701,In_271);
xor U3338 (N_3338,In_794,In_300);
nor U3339 (N_3339,In_806,In_173);
or U3340 (N_3340,In_472,In_610);
nor U3341 (N_3341,In_190,In_754);
or U3342 (N_3342,In_182,In_337);
or U3343 (N_3343,In_154,In_93);
nor U3344 (N_3344,In_795,In_692);
nand U3345 (N_3345,In_193,In_962);
xor U3346 (N_3346,In_481,In_759);
and U3347 (N_3347,In_686,In_279);
nand U3348 (N_3348,In_770,In_867);
and U3349 (N_3349,In_320,In_841);
and U3350 (N_3350,In_801,In_736);
or U3351 (N_3351,In_518,In_429);
nor U3352 (N_3352,In_809,In_883);
or U3353 (N_3353,In_848,In_551);
nand U3354 (N_3354,In_513,In_418);
nand U3355 (N_3355,In_960,In_361);
or U3356 (N_3356,In_947,In_8);
nand U3357 (N_3357,In_900,In_903);
or U3358 (N_3358,In_696,In_399);
nand U3359 (N_3359,In_735,In_246);
and U3360 (N_3360,In_306,In_100);
and U3361 (N_3361,In_878,In_224);
or U3362 (N_3362,In_789,In_668);
nand U3363 (N_3363,In_526,In_253);
or U3364 (N_3364,In_381,In_685);
nor U3365 (N_3365,In_729,In_955);
nor U3366 (N_3366,In_615,In_102);
nand U3367 (N_3367,In_151,In_214);
nand U3368 (N_3368,In_692,In_905);
or U3369 (N_3369,In_471,In_993);
and U3370 (N_3370,In_350,In_37);
or U3371 (N_3371,In_476,In_385);
nand U3372 (N_3372,In_830,In_972);
nand U3373 (N_3373,In_956,In_197);
nand U3374 (N_3374,In_966,In_113);
nand U3375 (N_3375,In_349,In_390);
nor U3376 (N_3376,In_616,In_62);
nor U3377 (N_3377,In_160,In_342);
and U3378 (N_3378,In_6,In_597);
and U3379 (N_3379,In_637,In_579);
and U3380 (N_3380,In_514,In_698);
nor U3381 (N_3381,In_865,In_195);
nand U3382 (N_3382,In_66,In_166);
nor U3383 (N_3383,In_740,In_1);
nor U3384 (N_3384,In_820,In_453);
nand U3385 (N_3385,In_616,In_625);
or U3386 (N_3386,In_548,In_340);
and U3387 (N_3387,In_885,In_998);
nor U3388 (N_3388,In_140,In_768);
nand U3389 (N_3389,In_57,In_408);
and U3390 (N_3390,In_287,In_513);
and U3391 (N_3391,In_553,In_882);
and U3392 (N_3392,In_950,In_651);
nand U3393 (N_3393,In_613,In_412);
and U3394 (N_3394,In_937,In_292);
nor U3395 (N_3395,In_136,In_836);
or U3396 (N_3396,In_631,In_84);
or U3397 (N_3397,In_734,In_737);
nand U3398 (N_3398,In_630,In_969);
and U3399 (N_3399,In_495,In_379);
and U3400 (N_3400,In_806,In_269);
or U3401 (N_3401,In_133,In_64);
nor U3402 (N_3402,In_838,In_569);
nor U3403 (N_3403,In_873,In_262);
nor U3404 (N_3404,In_289,In_510);
nand U3405 (N_3405,In_495,In_973);
nand U3406 (N_3406,In_184,In_159);
nand U3407 (N_3407,In_253,In_519);
and U3408 (N_3408,In_391,In_626);
xnor U3409 (N_3409,In_387,In_36);
and U3410 (N_3410,In_312,In_226);
and U3411 (N_3411,In_174,In_164);
nand U3412 (N_3412,In_995,In_872);
or U3413 (N_3413,In_334,In_971);
nor U3414 (N_3414,In_731,In_646);
or U3415 (N_3415,In_936,In_971);
and U3416 (N_3416,In_924,In_732);
or U3417 (N_3417,In_571,In_158);
nor U3418 (N_3418,In_128,In_322);
nor U3419 (N_3419,In_325,In_976);
and U3420 (N_3420,In_128,In_139);
nand U3421 (N_3421,In_941,In_162);
nand U3422 (N_3422,In_645,In_592);
nor U3423 (N_3423,In_855,In_154);
or U3424 (N_3424,In_28,In_343);
and U3425 (N_3425,In_759,In_527);
or U3426 (N_3426,In_585,In_48);
nor U3427 (N_3427,In_650,In_614);
or U3428 (N_3428,In_835,In_584);
nor U3429 (N_3429,In_184,In_894);
and U3430 (N_3430,In_320,In_757);
or U3431 (N_3431,In_934,In_720);
or U3432 (N_3432,In_800,In_700);
or U3433 (N_3433,In_941,In_148);
nand U3434 (N_3434,In_27,In_742);
nand U3435 (N_3435,In_967,In_292);
nor U3436 (N_3436,In_22,In_447);
nand U3437 (N_3437,In_840,In_188);
or U3438 (N_3438,In_908,In_384);
and U3439 (N_3439,In_214,In_686);
nor U3440 (N_3440,In_395,In_742);
nor U3441 (N_3441,In_942,In_9);
nor U3442 (N_3442,In_777,In_937);
and U3443 (N_3443,In_417,In_389);
nand U3444 (N_3444,In_756,In_4);
nor U3445 (N_3445,In_193,In_537);
nand U3446 (N_3446,In_35,In_412);
or U3447 (N_3447,In_379,In_323);
and U3448 (N_3448,In_317,In_756);
nor U3449 (N_3449,In_227,In_718);
nand U3450 (N_3450,In_264,In_598);
nand U3451 (N_3451,In_618,In_956);
and U3452 (N_3452,In_794,In_271);
nor U3453 (N_3453,In_374,In_248);
or U3454 (N_3454,In_51,In_713);
nor U3455 (N_3455,In_102,In_994);
nand U3456 (N_3456,In_95,In_887);
and U3457 (N_3457,In_194,In_299);
nand U3458 (N_3458,In_915,In_404);
or U3459 (N_3459,In_547,In_876);
nor U3460 (N_3460,In_269,In_892);
nand U3461 (N_3461,In_213,In_394);
or U3462 (N_3462,In_367,In_685);
nor U3463 (N_3463,In_929,In_544);
and U3464 (N_3464,In_435,In_142);
nor U3465 (N_3465,In_628,In_906);
nand U3466 (N_3466,In_747,In_532);
nor U3467 (N_3467,In_505,In_363);
nor U3468 (N_3468,In_434,In_874);
nor U3469 (N_3469,In_976,In_21);
and U3470 (N_3470,In_194,In_98);
or U3471 (N_3471,In_355,In_528);
nor U3472 (N_3472,In_885,In_12);
nor U3473 (N_3473,In_21,In_725);
nor U3474 (N_3474,In_865,In_327);
nand U3475 (N_3475,In_156,In_539);
nand U3476 (N_3476,In_735,In_963);
nor U3477 (N_3477,In_989,In_559);
and U3478 (N_3478,In_68,In_314);
nor U3479 (N_3479,In_691,In_531);
or U3480 (N_3480,In_181,In_406);
xor U3481 (N_3481,In_692,In_531);
nor U3482 (N_3482,In_438,In_157);
nor U3483 (N_3483,In_880,In_700);
nor U3484 (N_3484,In_833,In_292);
nor U3485 (N_3485,In_631,In_853);
nand U3486 (N_3486,In_148,In_317);
nor U3487 (N_3487,In_384,In_729);
nand U3488 (N_3488,In_239,In_770);
nor U3489 (N_3489,In_905,In_417);
or U3490 (N_3490,In_324,In_794);
and U3491 (N_3491,In_83,In_7);
nand U3492 (N_3492,In_136,In_508);
nor U3493 (N_3493,In_402,In_673);
or U3494 (N_3494,In_312,In_254);
nor U3495 (N_3495,In_395,In_174);
nor U3496 (N_3496,In_760,In_242);
nor U3497 (N_3497,In_607,In_430);
and U3498 (N_3498,In_526,In_984);
and U3499 (N_3499,In_978,In_232);
nand U3500 (N_3500,In_651,In_333);
nand U3501 (N_3501,In_904,In_359);
or U3502 (N_3502,In_665,In_973);
or U3503 (N_3503,In_811,In_41);
or U3504 (N_3504,In_898,In_187);
and U3505 (N_3505,In_255,In_708);
or U3506 (N_3506,In_796,In_346);
nand U3507 (N_3507,In_879,In_672);
nor U3508 (N_3508,In_808,In_679);
or U3509 (N_3509,In_99,In_494);
or U3510 (N_3510,In_561,In_528);
nor U3511 (N_3511,In_467,In_697);
or U3512 (N_3512,In_161,In_250);
nor U3513 (N_3513,In_208,In_33);
or U3514 (N_3514,In_926,In_671);
or U3515 (N_3515,In_251,In_422);
and U3516 (N_3516,In_344,In_796);
nor U3517 (N_3517,In_807,In_56);
nand U3518 (N_3518,In_702,In_994);
and U3519 (N_3519,In_439,In_352);
and U3520 (N_3520,In_140,In_491);
and U3521 (N_3521,In_333,In_425);
nand U3522 (N_3522,In_168,In_38);
nor U3523 (N_3523,In_159,In_503);
nand U3524 (N_3524,In_888,In_543);
nand U3525 (N_3525,In_759,In_932);
and U3526 (N_3526,In_473,In_931);
nor U3527 (N_3527,In_107,In_608);
nor U3528 (N_3528,In_172,In_318);
and U3529 (N_3529,In_743,In_934);
and U3530 (N_3530,In_580,In_907);
and U3531 (N_3531,In_210,In_170);
nor U3532 (N_3532,In_911,In_375);
or U3533 (N_3533,In_366,In_456);
nor U3534 (N_3534,In_234,In_414);
or U3535 (N_3535,In_682,In_381);
nor U3536 (N_3536,In_934,In_520);
nor U3537 (N_3537,In_96,In_436);
and U3538 (N_3538,In_733,In_334);
or U3539 (N_3539,In_210,In_731);
nor U3540 (N_3540,In_896,In_291);
nand U3541 (N_3541,In_298,In_870);
nand U3542 (N_3542,In_993,In_906);
nor U3543 (N_3543,In_438,In_730);
and U3544 (N_3544,In_905,In_877);
nand U3545 (N_3545,In_327,In_589);
or U3546 (N_3546,In_777,In_166);
nor U3547 (N_3547,In_464,In_463);
nor U3548 (N_3548,In_651,In_341);
or U3549 (N_3549,In_864,In_544);
and U3550 (N_3550,In_501,In_523);
nor U3551 (N_3551,In_427,In_706);
nor U3552 (N_3552,In_939,In_642);
and U3553 (N_3553,In_643,In_508);
or U3554 (N_3554,In_713,In_503);
nand U3555 (N_3555,In_74,In_504);
nand U3556 (N_3556,In_16,In_612);
nand U3557 (N_3557,In_581,In_567);
or U3558 (N_3558,In_800,In_993);
or U3559 (N_3559,In_72,In_392);
and U3560 (N_3560,In_291,In_507);
nand U3561 (N_3561,In_990,In_796);
nor U3562 (N_3562,In_950,In_814);
and U3563 (N_3563,In_985,In_192);
nor U3564 (N_3564,In_970,In_883);
nor U3565 (N_3565,In_379,In_198);
nor U3566 (N_3566,In_52,In_597);
or U3567 (N_3567,In_164,In_348);
nor U3568 (N_3568,In_361,In_651);
nand U3569 (N_3569,In_514,In_731);
nor U3570 (N_3570,In_935,In_963);
nor U3571 (N_3571,In_417,In_738);
or U3572 (N_3572,In_796,In_805);
and U3573 (N_3573,In_501,In_685);
nand U3574 (N_3574,In_579,In_400);
nor U3575 (N_3575,In_598,In_702);
and U3576 (N_3576,In_149,In_37);
nor U3577 (N_3577,In_326,In_963);
nor U3578 (N_3578,In_446,In_900);
nand U3579 (N_3579,In_645,In_35);
nand U3580 (N_3580,In_45,In_357);
nor U3581 (N_3581,In_31,In_426);
or U3582 (N_3582,In_220,In_384);
nor U3583 (N_3583,In_710,In_247);
or U3584 (N_3584,In_741,In_216);
or U3585 (N_3585,In_723,In_571);
and U3586 (N_3586,In_236,In_655);
and U3587 (N_3587,In_813,In_634);
and U3588 (N_3588,In_170,In_605);
and U3589 (N_3589,In_5,In_561);
xnor U3590 (N_3590,In_261,In_383);
nor U3591 (N_3591,In_853,In_333);
nor U3592 (N_3592,In_384,In_3);
or U3593 (N_3593,In_408,In_581);
or U3594 (N_3594,In_943,In_976);
nand U3595 (N_3595,In_773,In_998);
and U3596 (N_3596,In_484,In_588);
nand U3597 (N_3597,In_684,In_56);
nand U3598 (N_3598,In_990,In_448);
nor U3599 (N_3599,In_774,In_644);
nor U3600 (N_3600,In_345,In_666);
nand U3601 (N_3601,In_474,In_344);
nand U3602 (N_3602,In_560,In_11);
or U3603 (N_3603,In_797,In_18);
and U3604 (N_3604,In_451,In_421);
and U3605 (N_3605,In_868,In_962);
or U3606 (N_3606,In_332,In_54);
nor U3607 (N_3607,In_12,In_407);
or U3608 (N_3608,In_82,In_63);
or U3609 (N_3609,In_835,In_562);
nand U3610 (N_3610,In_288,In_493);
and U3611 (N_3611,In_831,In_217);
nor U3612 (N_3612,In_844,In_557);
and U3613 (N_3613,In_726,In_937);
and U3614 (N_3614,In_367,In_315);
nor U3615 (N_3615,In_278,In_268);
or U3616 (N_3616,In_981,In_576);
nor U3617 (N_3617,In_298,In_453);
nand U3618 (N_3618,In_486,In_987);
and U3619 (N_3619,In_471,In_41);
nor U3620 (N_3620,In_77,In_845);
nand U3621 (N_3621,In_440,In_240);
nor U3622 (N_3622,In_793,In_114);
nor U3623 (N_3623,In_45,In_881);
nand U3624 (N_3624,In_488,In_26);
and U3625 (N_3625,In_478,In_556);
or U3626 (N_3626,In_57,In_111);
and U3627 (N_3627,In_406,In_212);
nor U3628 (N_3628,In_412,In_97);
or U3629 (N_3629,In_601,In_676);
or U3630 (N_3630,In_414,In_49);
nor U3631 (N_3631,In_245,In_172);
nor U3632 (N_3632,In_579,In_449);
or U3633 (N_3633,In_990,In_668);
nor U3634 (N_3634,In_60,In_488);
or U3635 (N_3635,In_157,In_679);
nand U3636 (N_3636,In_619,In_967);
nand U3637 (N_3637,In_335,In_421);
or U3638 (N_3638,In_205,In_229);
or U3639 (N_3639,In_172,In_296);
nor U3640 (N_3640,In_596,In_907);
nand U3641 (N_3641,In_253,In_305);
nor U3642 (N_3642,In_509,In_639);
and U3643 (N_3643,In_766,In_929);
and U3644 (N_3644,In_22,In_878);
nor U3645 (N_3645,In_136,In_14);
and U3646 (N_3646,In_994,In_184);
nand U3647 (N_3647,In_92,In_709);
or U3648 (N_3648,In_734,In_269);
nor U3649 (N_3649,In_413,In_652);
or U3650 (N_3650,In_979,In_936);
or U3651 (N_3651,In_304,In_72);
or U3652 (N_3652,In_422,In_331);
nor U3653 (N_3653,In_77,In_385);
nor U3654 (N_3654,In_517,In_241);
or U3655 (N_3655,In_808,In_587);
or U3656 (N_3656,In_237,In_529);
nor U3657 (N_3657,In_23,In_85);
or U3658 (N_3658,In_970,In_917);
and U3659 (N_3659,In_437,In_822);
nand U3660 (N_3660,In_951,In_989);
nor U3661 (N_3661,In_189,In_871);
nor U3662 (N_3662,In_437,In_976);
and U3663 (N_3663,In_705,In_937);
and U3664 (N_3664,In_75,In_813);
and U3665 (N_3665,In_102,In_804);
nor U3666 (N_3666,In_497,In_485);
and U3667 (N_3667,In_338,In_759);
or U3668 (N_3668,In_501,In_296);
or U3669 (N_3669,In_881,In_895);
and U3670 (N_3670,In_96,In_820);
nor U3671 (N_3671,In_575,In_605);
or U3672 (N_3672,In_806,In_691);
or U3673 (N_3673,In_474,In_972);
and U3674 (N_3674,In_166,In_44);
and U3675 (N_3675,In_689,In_123);
and U3676 (N_3676,In_187,In_275);
nor U3677 (N_3677,In_646,In_793);
nand U3678 (N_3678,In_332,In_174);
nand U3679 (N_3679,In_194,In_85);
or U3680 (N_3680,In_29,In_327);
nor U3681 (N_3681,In_909,In_695);
nor U3682 (N_3682,In_595,In_75);
nand U3683 (N_3683,In_738,In_177);
and U3684 (N_3684,In_844,In_977);
nand U3685 (N_3685,In_868,In_854);
nor U3686 (N_3686,In_561,In_811);
or U3687 (N_3687,In_299,In_957);
nor U3688 (N_3688,In_327,In_829);
nand U3689 (N_3689,In_705,In_150);
or U3690 (N_3690,In_503,In_272);
nand U3691 (N_3691,In_522,In_685);
xor U3692 (N_3692,In_573,In_138);
or U3693 (N_3693,In_314,In_570);
nand U3694 (N_3694,In_72,In_411);
and U3695 (N_3695,In_499,In_687);
nand U3696 (N_3696,In_930,In_17);
nor U3697 (N_3697,In_685,In_243);
nor U3698 (N_3698,In_401,In_365);
nand U3699 (N_3699,In_695,In_239);
or U3700 (N_3700,In_327,In_364);
or U3701 (N_3701,In_378,In_407);
or U3702 (N_3702,In_405,In_684);
or U3703 (N_3703,In_756,In_95);
or U3704 (N_3704,In_790,In_581);
and U3705 (N_3705,In_495,In_53);
and U3706 (N_3706,In_653,In_30);
nor U3707 (N_3707,In_831,In_821);
nand U3708 (N_3708,In_93,In_303);
nand U3709 (N_3709,In_404,In_225);
and U3710 (N_3710,In_185,In_524);
nor U3711 (N_3711,In_587,In_541);
nand U3712 (N_3712,In_436,In_216);
or U3713 (N_3713,In_223,In_76);
nor U3714 (N_3714,In_805,In_665);
or U3715 (N_3715,In_654,In_768);
nor U3716 (N_3716,In_91,In_369);
or U3717 (N_3717,In_38,In_455);
nand U3718 (N_3718,In_578,In_129);
or U3719 (N_3719,In_275,In_11);
nand U3720 (N_3720,In_653,In_161);
nor U3721 (N_3721,In_236,In_992);
nor U3722 (N_3722,In_554,In_61);
and U3723 (N_3723,In_647,In_65);
nand U3724 (N_3724,In_755,In_863);
nand U3725 (N_3725,In_603,In_908);
nor U3726 (N_3726,In_627,In_438);
or U3727 (N_3727,In_664,In_183);
nand U3728 (N_3728,In_774,In_557);
nor U3729 (N_3729,In_563,In_370);
and U3730 (N_3730,In_855,In_691);
or U3731 (N_3731,In_868,In_122);
nand U3732 (N_3732,In_208,In_739);
nor U3733 (N_3733,In_920,In_402);
and U3734 (N_3734,In_504,In_857);
nand U3735 (N_3735,In_715,In_604);
or U3736 (N_3736,In_566,In_240);
nor U3737 (N_3737,In_426,In_29);
nand U3738 (N_3738,In_880,In_12);
or U3739 (N_3739,In_121,In_890);
or U3740 (N_3740,In_257,In_563);
xnor U3741 (N_3741,In_15,In_379);
or U3742 (N_3742,In_242,In_530);
or U3743 (N_3743,In_173,In_205);
and U3744 (N_3744,In_519,In_830);
nand U3745 (N_3745,In_850,In_119);
or U3746 (N_3746,In_190,In_664);
nor U3747 (N_3747,In_586,In_160);
or U3748 (N_3748,In_339,In_463);
or U3749 (N_3749,In_856,In_725);
or U3750 (N_3750,In_816,In_675);
or U3751 (N_3751,In_361,In_444);
and U3752 (N_3752,In_0,In_368);
and U3753 (N_3753,In_977,In_687);
nor U3754 (N_3754,In_606,In_417);
and U3755 (N_3755,In_835,In_208);
or U3756 (N_3756,In_956,In_811);
nand U3757 (N_3757,In_477,In_254);
nor U3758 (N_3758,In_34,In_937);
nor U3759 (N_3759,In_306,In_719);
nor U3760 (N_3760,In_356,In_230);
nor U3761 (N_3761,In_470,In_413);
nand U3762 (N_3762,In_360,In_750);
and U3763 (N_3763,In_444,In_330);
nor U3764 (N_3764,In_103,In_663);
or U3765 (N_3765,In_606,In_967);
nand U3766 (N_3766,In_577,In_104);
nor U3767 (N_3767,In_249,In_693);
nor U3768 (N_3768,In_715,In_256);
nor U3769 (N_3769,In_317,In_57);
and U3770 (N_3770,In_792,In_156);
and U3771 (N_3771,In_735,In_791);
and U3772 (N_3772,In_453,In_736);
and U3773 (N_3773,In_405,In_629);
or U3774 (N_3774,In_689,In_757);
nand U3775 (N_3775,In_893,In_987);
or U3776 (N_3776,In_95,In_972);
nand U3777 (N_3777,In_401,In_804);
and U3778 (N_3778,In_314,In_572);
nor U3779 (N_3779,In_215,In_227);
nand U3780 (N_3780,In_637,In_114);
or U3781 (N_3781,In_559,In_58);
and U3782 (N_3782,In_557,In_653);
and U3783 (N_3783,In_457,In_763);
or U3784 (N_3784,In_218,In_162);
nor U3785 (N_3785,In_585,In_400);
or U3786 (N_3786,In_819,In_984);
nor U3787 (N_3787,In_207,In_47);
and U3788 (N_3788,In_963,In_942);
and U3789 (N_3789,In_640,In_355);
and U3790 (N_3790,In_605,In_463);
nand U3791 (N_3791,In_474,In_856);
and U3792 (N_3792,In_334,In_897);
nor U3793 (N_3793,In_279,In_960);
or U3794 (N_3794,In_571,In_576);
nand U3795 (N_3795,In_621,In_758);
or U3796 (N_3796,In_986,In_900);
nand U3797 (N_3797,In_392,In_421);
nand U3798 (N_3798,In_839,In_603);
or U3799 (N_3799,In_873,In_864);
or U3800 (N_3800,In_879,In_137);
or U3801 (N_3801,In_50,In_508);
and U3802 (N_3802,In_989,In_432);
and U3803 (N_3803,In_92,In_800);
nor U3804 (N_3804,In_765,In_97);
or U3805 (N_3805,In_499,In_500);
nor U3806 (N_3806,In_843,In_733);
nor U3807 (N_3807,In_34,In_135);
nor U3808 (N_3808,In_717,In_508);
xor U3809 (N_3809,In_524,In_800);
nand U3810 (N_3810,In_710,In_27);
or U3811 (N_3811,In_131,In_934);
or U3812 (N_3812,In_724,In_878);
nand U3813 (N_3813,In_983,In_51);
and U3814 (N_3814,In_821,In_648);
or U3815 (N_3815,In_393,In_465);
and U3816 (N_3816,In_25,In_98);
nor U3817 (N_3817,In_27,In_951);
or U3818 (N_3818,In_700,In_28);
nor U3819 (N_3819,In_897,In_875);
and U3820 (N_3820,In_166,In_960);
nor U3821 (N_3821,In_427,In_220);
nor U3822 (N_3822,In_434,In_641);
and U3823 (N_3823,In_486,In_216);
or U3824 (N_3824,In_87,In_301);
or U3825 (N_3825,In_542,In_978);
nand U3826 (N_3826,In_890,In_746);
nand U3827 (N_3827,In_808,In_807);
nor U3828 (N_3828,In_31,In_294);
xor U3829 (N_3829,In_433,In_512);
and U3830 (N_3830,In_706,In_535);
nand U3831 (N_3831,In_729,In_920);
nand U3832 (N_3832,In_727,In_84);
nand U3833 (N_3833,In_552,In_170);
nor U3834 (N_3834,In_73,In_965);
nor U3835 (N_3835,In_509,In_596);
nand U3836 (N_3836,In_738,In_295);
nand U3837 (N_3837,In_201,In_365);
nor U3838 (N_3838,In_591,In_401);
nor U3839 (N_3839,In_326,In_865);
and U3840 (N_3840,In_379,In_349);
nor U3841 (N_3841,In_737,In_192);
nand U3842 (N_3842,In_756,In_50);
nand U3843 (N_3843,In_124,In_526);
and U3844 (N_3844,In_241,In_249);
or U3845 (N_3845,In_850,In_279);
nor U3846 (N_3846,In_513,In_870);
nand U3847 (N_3847,In_884,In_96);
nand U3848 (N_3848,In_344,In_27);
nand U3849 (N_3849,In_629,In_585);
and U3850 (N_3850,In_59,In_876);
and U3851 (N_3851,In_297,In_229);
or U3852 (N_3852,In_190,In_851);
and U3853 (N_3853,In_649,In_944);
nand U3854 (N_3854,In_158,In_145);
and U3855 (N_3855,In_494,In_453);
or U3856 (N_3856,In_986,In_951);
or U3857 (N_3857,In_425,In_748);
and U3858 (N_3858,In_866,In_326);
nand U3859 (N_3859,In_10,In_699);
or U3860 (N_3860,In_936,In_734);
or U3861 (N_3861,In_935,In_537);
nor U3862 (N_3862,In_145,In_898);
nand U3863 (N_3863,In_413,In_635);
nor U3864 (N_3864,In_363,In_358);
nor U3865 (N_3865,In_934,In_609);
or U3866 (N_3866,In_982,In_370);
or U3867 (N_3867,In_740,In_516);
nand U3868 (N_3868,In_18,In_858);
or U3869 (N_3869,In_695,In_592);
nand U3870 (N_3870,In_382,In_88);
and U3871 (N_3871,In_876,In_296);
or U3872 (N_3872,In_557,In_135);
nand U3873 (N_3873,In_264,In_406);
nand U3874 (N_3874,In_786,In_803);
or U3875 (N_3875,In_963,In_580);
and U3876 (N_3876,In_587,In_971);
and U3877 (N_3877,In_514,In_893);
nor U3878 (N_3878,In_71,In_897);
nand U3879 (N_3879,In_863,In_603);
nor U3880 (N_3880,In_416,In_435);
nand U3881 (N_3881,In_706,In_437);
or U3882 (N_3882,In_770,In_190);
or U3883 (N_3883,In_994,In_392);
nor U3884 (N_3884,In_914,In_769);
or U3885 (N_3885,In_647,In_430);
or U3886 (N_3886,In_732,In_27);
and U3887 (N_3887,In_934,In_528);
nand U3888 (N_3888,In_965,In_286);
nor U3889 (N_3889,In_398,In_107);
or U3890 (N_3890,In_822,In_584);
nand U3891 (N_3891,In_326,In_217);
nand U3892 (N_3892,In_406,In_745);
nor U3893 (N_3893,In_115,In_757);
and U3894 (N_3894,In_83,In_123);
nand U3895 (N_3895,In_341,In_649);
nand U3896 (N_3896,In_825,In_937);
nand U3897 (N_3897,In_10,In_629);
or U3898 (N_3898,In_193,In_618);
or U3899 (N_3899,In_121,In_876);
and U3900 (N_3900,In_742,In_329);
or U3901 (N_3901,In_113,In_702);
nor U3902 (N_3902,In_959,In_985);
and U3903 (N_3903,In_377,In_656);
nor U3904 (N_3904,In_718,In_368);
and U3905 (N_3905,In_300,In_641);
nand U3906 (N_3906,In_266,In_402);
or U3907 (N_3907,In_216,In_215);
nand U3908 (N_3908,In_617,In_623);
and U3909 (N_3909,In_464,In_701);
and U3910 (N_3910,In_791,In_535);
nand U3911 (N_3911,In_864,In_721);
or U3912 (N_3912,In_970,In_423);
or U3913 (N_3913,In_255,In_2);
and U3914 (N_3914,In_200,In_812);
and U3915 (N_3915,In_245,In_101);
and U3916 (N_3916,In_112,In_596);
or U3917 (N_3917,In_67,In_110);
nand U3918 (N_3918,In_512,In_486);
or U3919 (N_3919,In_537,In_391);
nand U3920 (N_3920,In_762,In_858);
and U3921 (N_3921,In_278,In_768);
and U3922 (N_3922,In_8,In_804);
nor U3923 (N_3923,In_191,In_91);
nand U3924 (N_3924,In_568,In_87);
nand U3925 (N_3925,In_160,In_531);
nor U3926 (N_3926,In_812,In_396);
or U3927 (N_3927,In_208,In_666);
nor U3928 (N_3928,In_209,In_966);
nor U3929 (N_3929,In_445,In_67);
nor U3930 (N_3930,In_595,In_0);
and U3931 (N_3931,In_508,In_886);
and U3932 (N_3932,In_522,In_210);
and U3933 (N_3933,In_431,In_522);
and U3934 (N_3934,In_866,In_514);
or U3935 (N_3935,In_30,In_529);
and U3936 (N_3936,In_67,In_126);
and U3937 (N_3937,In_584,In_206);
nand U3938 (N_3938,In_231,In_598);
or U3939 (N_3939,In_241,In_452);
nand U3940 (N_3940,In_851,In_145);
nor U3941 (N_3941,In_557,In_229);
nand U3942 (N_3942,In_169,In_516);
or U3943 (N_3943,In_154,In_647);
and U3944 (N_3944,In_399,In_570);
or U3945 (N_3945,In_951,In_540);
or U3946 (N_3946,In_922,In_274);
or U3947 (N_3947,In_862,In_984);
and U3948 (N_3948,In_13,In_113);
nor U3949 (N_3949,In_780,In_821);
and U3950 (N_3950,In_11,In_589);
nand U3951 (N_3951,In_654,In_471);
nand U3952 (N_3952,In_626,In_1);
or U3953 (N_3953,In_880,In_604);
or U3954 (N_3954,In_955,In_105);
nor U3955 (N_3955,In_305,In_598);
and U3956 (N_3956,In_283,In_529);
nor U3957 (N_3957,In_492,In_387);
nand U3958 (N_3958,In_71,In_899);
and U3959 (N_3959,In_548,In_621);
nor U3960 (N_3960,In_278,In_732);
and U3961 (N_3961,In_595,In_47);
and U3962 (N_3962,In_433,In_851);
nand U3963 (N_3963,In_354,In_895);
nand U3964 (N_3964,In_353,In_65);
or U3965 (N_3965,In_296,In_570);
or U3966 (N_3966,In_32,In_433);
nor U3967 (N_3967,In_974,In_144);
nor U3968 (N_3968,In_805,In_225);
nand U3969 (N_3969,In_731,In_540);
nand U3970 (N_3970,In_368,In_376);
and U3971 (N_3971,In_299,In_780);
and U3972 (N_3972,In_500,In_52);
nor U3973 (N_3973,In_467,In_212);
nand U3974 (N_3974,In_353,In_2);
nand U3975 (N_3975,In_91,In_197);
xor U3976 (N_3976,In_26,In_381);
nor U3977 (N_3977,In_527,In_677);
nor U3978 (N_3978,In_469,In_242);
and U3979 (N_3979,In_994,In_738);
and U3980 (N_3980,In_105,In_872);
and U3981 (N_3981,In_266,In_813);
or U3982 (N_3982,In_399,In_576);
nand U3983 (N_3983,In_948,In_514);
nor U3984 (N_3984,In_849,In_802);
or U3985 (N_3985,In_529,In_978);
nand U3986 (N_3986,In_910,In_339);
or U3987 (N_3987,In_412,In_254);
nor U3988 (N_3988,In_115,In_588);
or U3989 (N_3989,In_943,In_701);
nor U3990 (N_3990,In_146,In_500);
nand U3991 (N_3991,In_568,In_617);
and U3992 (N_3992,In_175,In_707);
or U3993 (N_3993,In_163,In_223);
and U3994 (N_3994,In_187,In_169);
or U3995 (N_3995,In_766,In_500);
or U3996 (N_3996,In_114,In_623);
nand U3997 (N_3997,In_960,In_72);
xnor U3998 (N_3998,In_174,In_595);
nor U3999 (N_3999,In_513,In_297);
or U4000 (N_4000,In_426,In_970);
and U4001 (N_4001,In_636,In_866);
nand U4002 (N_4002,In_908,In_653);
or U4003 (N_4003,In_894,In_281);
or U4004 (N_4004,In_943,In_627);
and U4005 (N_4005,In_268,In_697);
and U4006 (N_4006,In_558,In_815);
nor U4007 (N_4007,In_218,In_105);
and U4008 (N_4008,In_845,In_895);
and U4009 (N_4009,In_246,In_552);
nand U4010 (N_4010,In_132,In_540);
or U4011 (N_4011,In_143,In_821);
nand U4012 (N_4012,In_433,In_838);
and U4013 (N_4013,In_314,In_64);
nor U4014 (N_4014,In_126,In_558);
or U4015 (N_4015,In_972,In_532);
and U4016 (N_4016,In_161,In_530);
or U4017 (N_4017,In_256,In_341);
and U4018 (N_4018,In_673,In_820);
xor U4019 (N_4019,In_139,In_730);
and U4020 (N_4020,In_757,In_729);
and U4021 (N_4021,In_405,In_291);
nand U4022 (N_4022,In_516,In_987);
or U4023 (N_4023,In_782,In_444);
nor U4024 (N_4024,In_254,In_684);
and U4025 (N_4025,In_942,In_111);
nand U4026 (N_4026,In_560,In_901);
and U4027 (N_4027,In_592,In_867);
and U4028 (N_4028,In_898,In_289);
nand U4029 (N_4029,In_431,In_826);
nor U4030 (N_4030,In_335,In_165);
nand U4031 (N_4031,In_146,In_681);
and U4032 (N_4032,In_3,In_64);
or U4033 (N_4033,In_139,In_157);
nor U4034 (N_4034,In_290,In_934);
nand U4035 (N_4035,In_635,In_201);
or U4036 (N_4036,In_349,In_545);
nand U4037 (N_4037,In_630,In_662);
and U4038 (N_4038,In_417,In_847);
nand U4039 (N_4039,In_384,In_132);
nand U4040 (N_4040,In_4,In_767);
nand U4041 (N_4041,In_927,In_226);
or U4042 (N_4042,In_764,In_146);
xor U4043 (N_4043,In_691,In_606);
nor U4044 (N_4044,In_252,In_152);
or U4045 (N_4045,In_378,In_953);
or U4046 (N_4046,In_571,In_103);
nor U4047 (N_4047,In_194,In_203);
nor U4048 (N_4048,In_293,In_225);
or U4049 (N_4049,In_986,In_451);
and U4050 (N_4050,In_621,In_622);
or U4051 (N_4051,In_505,In_181);
nand U4052 (N_4052,In_942,In_446);
or U4053 (N_4053,In_299,In_903);
and U4054 (N_4054,In_618,In_952);
and U4055 (N_4055,In_376,In_651);
and U4056 (N_4056,In_215,In_567);
nor U4057 (N_4057,In_727,In_48);
nand U4058 (N_4058,In_838,In_605);
nand U4059 (N_4059,In_348,In_645);
or U4060 (N_4060,In_486,In_976);
nand U4061 (N_4061,In_506,In_527);
nor U4062 (N_4062,In_421,In_309);
and U4063 (N_4063,In_993,In_228);
nand U4064 (N_4064,In_268,In_628);
or U4065 (N_4065,In_198,In_930);
nand U4066 (N_4066,In_34,In_148);
and U4067 (N_4067,In_338,In_852);
and U4068 (N_4068,In_329,In_765);
and U4069 (N_4069,In_404,In_58);
and U4070 (N_4070,In_298,In_34);
and U4071 (N_4071,In_862,In_341);
nand U4072 (N_4072,In_446,In_142);
nor U4073 (N_4073,In_413,In_927);
or U4074 (N_4074,In_767,In_181);
nor U4075 (N_4075,In_417,In_684);
and U4076 (N_4076,In_484,In_475);
nand U4077 (N_4077,In_348,In_792);
or U4078 (N_4078,In_891,In_254);
or U4079 (N_4079,In_856,In_872);
and U4080 (N_4080,In_541,In_52);
and U4081 (N_4081,In_192,In_856);
nor U4082 (N_4082,In_449,In_221);
and U4083 (N_4083,In_704,In_639);
and U4084 (N_4084,In_123,In_502);
and U4085 (N_4085,In_634,In_51);
nor U4086 (N_4086,In_220,In_609);
nand U4087 (N_4087,In_262,In_694);
nor U4088 (N_4088,In_34,In_95);
or U4089 (N_4089,In_831,In_550);
nor U4090 (N_4090,In_293,In_344);
nand U4091 (N_4091,In_805,In_356);
nor U4092 (N_4092,In_578,In_865);
nand U4093 (N_4093,In_629,In_334);
nand U4094 (N_4094,In_349,In_664);
and U4095 (N_4095,In_965,In_49);
or U4096 (N_4096,In_60,In_309);
nand U4097 (N_4097,In_376,In_372);
nor U4098 (N_4098,In_614,In_589);
nand U4099 (N_4099,In_356,In_943);
nand U4100 (N_4100,In_9,In_98);
nand U4101 (N_4101,In_281,In_306);
or U4102 (N_4102,In_906,In_753);
or U4103 (N_4103,In_874,In_298);
or U4104 (N_4104,In_373,In_150);
and U4105 (N_4105,In_976,In_960);
nor U4106 (N_4106,In_128,In_754);
xor U4107 (N_4107,In_640,In_834);
or U4108 (N_4108,In_807,In_442);
and U4109 (N_4109,In_310,In_298);
nand U4110 (N_4110,In_373,In_48);
nor U4111 (N_4111,In_755,In_104);
and U4112 (N_4112,In_638,In_807);
or U4113 (N_4113,In_312,In_791);
xnor U4114 (N_4114,In_845,In_966);
nand U4115 (N_4115,In_70,In_506);
or U4116 (N_4116,In_142,In_827);
nand U4117 (N_4117,In_739,In_748);
and U4118 (N_4118,In_519,In_264);
or U4119 (N_4119,In_729,In_470);
nand U4120 (N_4120,In_133,In_21);
xnor U4121 (N_4121,In_910,In_523);
nor U4122 (N_4122,In_480,In_472);
and U4123 (N_4123,In_863,In_943);
and U4124 (N_4124,In_305,In_242);
and U4125 (N_4125,In_294,In_355);
nor U4126 (N_4126,In_270,In_212);
nor U4127 (N_4127,In_509,In_75);
or U4128 (N_4128,In_224,In_729);
and U4129 (N_4129,In_129,In_332);
nand U4130 (N_4130,In_785,In_378);
nor U4131 (N_4131,In_924,In_138);
and U4132 (N_4132,In_26,In_147);
nand U4133 (N_4133,In_310,In_972);
nand U4134 (N_4134,In_496,In_145);
nand U4135 (N_4135,In_489,In_116);
and U4136 (N_4136,In_880,In_465);
nor U4137 (N_4137,In_443,In_57);
nor U4138 (N_4138,In_944,In_408);
nand U4139 (N_4139,In_907,In_113);
and U4140 (N_4140,In_502,In_949);
and U4141 (N_4141,In_584,In_269);
nand U4142 (N_4142,In_116,In_189);
or U4143 (N_4143,In_19,In_186);
and U4144 (N_4144,In_550,In_702);
nor U4145 (N_4145,In_287,In_347);
and U4146 (N_4146,In_474,In_844);
and U4147 (N_4147,In_432,In_263);
nor U4148 (N_4148,In_108,In_96);
and U4149 (N_4149,In_654,In_269);
nor U4150 (N_4150,In_504,In_299);
xor U4151 (N_4151,In_409,In_879);
nor U4152 (N_4152,In_20,In_656);
and U4153 (N_4153,In_245,In_521);
nor U4154 (N_4154,In_146,In_519);
nand U4155 (N_4155,In_552,In_461);
or U4156 (N_4156,In_597,In_687);
or U4157 (N_4157,In_914,In_321);
and U4158 (N_4158,In_551,In_863);
and U4159 (N_4159,In_607,In_611);
or U4160 (N_4160,In_360,In_499);
nand U4161 (N_4161,In_641,In_193);
and U4162 (N_4162,In_547,In_327);
and U4163 (N_4163,In_909,In_622);
and U4164 (N_4164,In_213,In_273);
or U4165 (N_4165,In_413,In_869);
nand U4166 (N_4166,In_581,In_420);
or U4167 (N_4167,In_496,In_421);
and U4168 (N_4168,In_617,In_588);
nor U4169 (N_4169,In_933,In_729);
nor U4170 (N_4170,In_658,In_720);
or U4171 (N_4171,In_392,In_659);
and U4172 (N_4172,In_444,In_722);
or U4173 (N_4173,In_125,In_649);
or U4174 (N_4174,In_237,In_999);
nand U4175 (N_4175,In_54,In_95);
and U4176 (N_4176,In_310,In_102);
nand U4177 (N_4177,In_867,In_70);
and U4178 (N_4178,In_408,In_589);
nand U4179 (N_4179,In_663,In_598);
and U4180 (N_4180,In_762,In_52);
nor U4181 (N_4181,In_330,In_687);
nand U4182 (N_4182,In_636,In_756);
nand U4183 (N_4183,In_733,In_864);
nor U4184 (N_4184,In_112,In_746);
nand U4185 (N_4185,In_606,In_451);
nand U4186 (N_4186,In_138,In_85);
and U4187 (N_4187,In_732,In_415);
nor U4188 (N_4188,In_389,In_324);
and U4189 (N_4189,In_653,In_902);
or U4190 (N_4190,In_483,In_861);
and U4191 (N_4191,In_814,In_170);
and U4192 (N_4192,In_149,In_614);
and U4193 (N_4193,In_98,In_474);
and U4194 (N_4194,In_835,In_726);
or U4195 (N_4195,In_732,In_952);
or U4196 (N_4196,In_330,In_463);
nand U4197 (N_4197,In_484,In_151);
and U4198 (N_4198,In_699,In_898);
nand U4199 (N_4199,In_171,In_195);
or U4200 (N_4200,In_250,In_86);
nand U4201 (N_4201,In_417,In_789);
and U4202 (N_4202,In_249,In_463);
nand U4203 (N_4203,In_193,In_538);
nor U4204 (N_4204,In_309,In_785);
and U4205 (N_4205,In_64,In_455);
or U4206 (N_4206,In_559,In_284);
nand U4207 (N_4207,In_607,In_509);
and U4208 (N_4208,In_935,In_848);
nor U4209 (N_4209,In_439,In_74);
or U4210 (N_4210,In_40,In_726);
nand U4211 (N_4211,In_693,In_114);
or U4212 (N_4212,In_466,In_687);
and U4213 (N_4213,In_250,In_910);
and U4214 (N_4214,In_352,In_778);
nand U4215 (N_4215,In_843,In_32);
or U4216 (N_4216,In_579,In_859);
or U4217 (N_4217,In_848,In_985);
and U4218 (N_4218,In_70,In_341);
and U4219 (N_4219,In_434,In_640);
or U4220 (N_4220,In_98,In_759);
or U4221 (N_4221,In_206,In_2);
or U4222 (N_4222,In_641,In_123);
nand U4223 (N_4223,In_155,In_43);
or U4224 (N_4224,In_168,In_365);
nor U4225 (N_4225,In_847,In_574);
or U4226 (N_4226,In_285,In_959);
nand U4227 (N_4227,In_15,In_199);
or U4228 (N_4228,In_764,In_189);
nand U4229 (N_4229,In_249,In_143);
nand U4230 (N_4230,In_382,In_113);
and U4231 (N_4231,In_321,In_127);
and U4232 (N_4232,In_259,In_570);
nor U4233 (N_4233,In_823,In_694);
and U4234 (N_4234,In_894,In_38);
nand U4235 (N_4235,In_26,In_180);
nand U4236 (N_4236,In_382,In_822);
nand U4237 (N_4237,In_939,In_921);
xnor U4238 (N_4238,In_92,In_367);
and U4239 (N_4239,In_497,In_715);
nor U4240 (N_4240,In_490,In_807);
nor U4241 (N_4241,In_978,In_819);
and U4242 (N_4242,In_707,In_880);
or U4243 (N_4243,In_156,In_489);
nor U4244 (N_4244,In_147,In_105);
nand U4245 (N_4245,In_246,In_564);
and U4246 (N_4246,In_96,In_535);
nor U4247 (N_4247,In_424,In_493);
or U4248 (N_4248,In_660,In_820);
nor U4249 (N_4249,In_786,In_485);
or U4250 (N_4250,In_4,In_85);
or U4251 (N_4251,In_665,In_526);
and U4252 (N_4252,In_435,In_308);
nand U4253 (N_4253,In_548,In_285);
nor U4254 (N_4254,In_896,In_158);
and U4255 (N_4255,In_667,In_146);
nand U4256 (N_4256,In_306,In_88);
and U4257 (N_4257,In_337,In_449);
and U4258 (N_4258,In_837,In_470);
and U4259 (N_4259,In_453,In_497);
and U4260 (N_4260,In_987,In_780);
xnor U4261 (N_4261,In_134,In_14);
nor U4262 (N_4262,In_588,In_7);
nand U4263 (N_4263,In_710,In_622);
nor U4264 (N_4264,In_882,In_891);
and U4265 (N_4265,In_849,In_130);
and U4266 (N_4266,In_123,In_706);
or U4267 (N_4267,In_967,In_344);
or U4268 (N_4268,In_220,In_224);
and U4269 (N_4269,In_909,In_336);
or U4270 (N_4270,In_832,In_62);
nand U4271 (N_4271,In_638,In_68);
nor U4272 (N_4272,In_465,In_822);
nor U4273 (N_4273,In_721,In_546);
or U4274 (N_4274,In_728,In_659);
and U4275 (N_4275,In_608,In_785);
or U4276 (N_4276,In_500,In_969);
or U4277 (N_4277,In_470,In_617);
nor U4278 (N_4278,In_408,In_824);
nor U4279 (N_4279,In_285,In_500);
or U4280 (N_4280,In_455,In_708);
or U4281 (N_4281,In_953,In_252);
nor U4282 (N_4282,In_50,In_599);
nor U4283 (N_4283,In_18,In_656);
nand U4284 (N_4284,In_987,In_935);
nor U4285 (N_4285,In_852,In_74);
and U4286 (N_4286,In_287,In_232);
and U4287 (N_4287,In_270,In_643);
and U4288 (N_4288,In_182,In_825);
nor U4289 (N_4289,In_269,In_554);
and U4290 (N_4290,In_436,In_618);
and U4291 (N_4291,In_147,In_726);
and U4292 (N_4292,In_643,In_254);
or U4293 (N_4293,In_653,In_531);
nand U4294 (N_4294,In_894,In_249);
or U4295 (N_4295,In_31,In_516);
nand U4296 (N_4296,In_861,In_860);
nor U4297 (N_4297,In_590,In_192);
nor U4298 (N_4298,In_325,In_511);
nand U4299 (N_4299,In_257,In_55);
and U4300 (N_4300,In_593,In_113);
and U4301 (N_4301,In_625,In_594);
and U4302 (N_4302,In_713,In_497);
or U4303 (N_4303,In_732,In_609);
nand U4304 (N_4304,In_474,In_847);
and U4305 (N_4305,In_370,In_653);
or U4306 (N_4306,In_432,In_444);
or U4307 (N_4307,In_523,In_110);
and U4308 (N_4308,In_446,In_733);
nand U4309 (N_4309,In_616,In_622);
nand U4310 (N_4310,In_687,In_769);
or U4311 (N_4311,In_40,In_94);
nand U4312 (N_4312,In_359,In_895);
and U4313 (N_4313,In_500,In_415);
nand U4314 (N_4314,In_574,In_266);
and U4315 (N_4315,In_783,In_943);
and U4316 (N_4316,In_62,In_135);
and U4317 (N_4317,In_195,In_994);
nor U4318 (N_4318,In_127,In_265);
and U4319 (N_4319,In_638,In_432);
nand U4320 (N_4320,In_317,In_269);
or U4321 (N_4321,In_876,In_367);
or U4322 (N_4322,In_928,In_272);
or U4323 (N_4323,In_741,In_385);
or U4324 (N_4324,In_274,In_1);
nand U4325 (N_4325,In_563,In_800);
or U4326 (N_4326,In_431,In_229);
nand U4327 (N_4327,In_9,In_106);
and U4328 (N_4328,In_389,In_151);
and U4329 (N_4329,In_374,In_142);
and U4330 (N_4330,In_351,In_770);
nor U4331 (N_4331,In_549,In_91);
nand U4332 (N_4332,In_536,In_59);
or U4333 (N_4333,In_733,In_695);
and U4334 (N_4334,In_482,In_118);
or U4335 (N_4335,In_351,In_272);
nor U4336 (N_4336,In_73,In_293);
or U4337 (N_4337,In_805,In_650);
nor U4338 (N_4338,In_54,In_563);
nand U4339 (N_4339,In_547,In_129);
nand U4340 (N_4340,In_283,In_296);
or U4341 (N_4341,In_870,In_120);
and U4342 (N_4342,In_291,In_830);
nand U4343 (N_4343,In_536,In_368);
or U4344 (N_4344,In_741,In_517);
or U4345 (N_4345,In_798,In_929);
nand U4346 (N_4346,In_781,In_207);
nand U4347 (N_4347,In_781,In_984);
or U4348 (N_4348,In_695,In_469);
or U4349 (N_4349,In_938,In_566);
or U4350 (N_4350,In_382,In_524);
or U4351 (N_4351,In_528,In_193);
or U4352 (N_4352,In_876,In_730);
nand U4353 (N_4353,In_325,In_199);
and U4354 (N_4354,In_985,In_301);
nand U4355 (N_4355,In_449,In_218);
and U4356 (N_4356,In_720,In_983);
xnor U4357 (N_4357,In_592,In_197);
nand U4358 (N_4358,In_774,In_426);
nor U4359 (N_4359,In_270,In_304);
and U4360 (N_4360,In_587,In_792);
nand U4361 (N_4361,In_149,In_32);
nor U4362 (N_4362,In_379,In_940);
nor U4363 (N_4363,In_793,In_326);
and U4364 (N_4364,In_984,In_267);
and U4365 (N_4365,In_697,In_514);
nand U4366 (N_4366,In_926,In_8);
and U4367 (N_4367,In_627,In_265);
nand U4368 (N_4368,In_488,In_956);
nor U4369 (N_4369,In_146,In_126);
nand U4370 (N_4370,In_882,In_844);
xor U4371 (N_4371,In_208,In_32);
nand U4372 (N_4372,In_677,In_817);
or U4373 (N_4373,In_217,In_420);
nand U4374 (N_4374,In_746,In_300);
xor U4375 (N_4375,In_40,In_30);
or U4376 (N_4376,In_358,In_230);
nand U4377 (N_4377,In_496,In_168);
nor U4378 (N_4378,In_523,In_114);
nand U4379 (N_4379,In_385,In_372);
xor U4380 (N_4380,In_115,In_576);
nor U4381 (N_4381,In_766,In_503);
xor U4382 (N_4382,In_324,In_844);
nor U4383 (N_4383,In_384,In_321);
and U4384 (N_4384,In_864,In_892);
nor U4385 (N_4385,In_43,In_625);
and U4386 (N_4386,In_743,In_689);
or U4387 (N_4387,In_307,In_971);
or U4388 (N_4388,In_187,In_33);
nand U4389 (N_4389,In_365,In_785);
nand U4390 (N_4390,In_555,In_129);
xnor U4391 (N_4391,In_231,In_210);
or U4392 (N_4392,In_763,In_606);
nand U4393 (N_4393,In_81,In_417);
and U4394 (N_4394,In_485,In_586);
and U4395 (N_4395,In_134,In_557);
nor U4396 (N_4396,In_288,In_478);
xnor U4397 (N_4397,In_725,In_164);
nor U4398 (N_4398,In_963,In_34);
and U4399 (N_4399,In_273,In_486);
or U4400 (N_4400,In_77,In_92);
nand U4401 (N_4401,In_859,In_406);
and U4402 (N_4402,In_880,In_489);
or U4403 (N_4403,In_248,In_319);
xnor U4404 (N_4404,In_798,In_484);
or U4405 (N_4405,In_994,In_782);
nor U4406 (N_4406,In_33,In_671);
nand U4407 (N_4407,In_354,In_984);
nor U4408 (N_4408,In_329,In_13);
nand U4409 (N_4409,In_585,In_88);
nand U4410 (N_4410,In_450,In_259);
and U4411 (N_4411,In_68,In_344);
nor U4412 (N_4412,In_766,In_373);
or U4413 (N_4413,In_640,In_598);
nor U4414 (N_4414,In_947,In_67);
and U4415 (N_4415,In_107,In_77);
nor U4416 (N_4416,In_536,In_339);
and U4417 (N_4417,In_375,In_360);
xor U4418 (N_4418,In_388,In_530);
or U4419 (N_4419,In_369,In_341);
and U4420 (N_4420,In_824,In_688);
and U4421 (N_4421,In_90,In_105);
and U4422 (N_4422,In_59,In_383);
nor U4423 (N_4423,In_229,In_166);
nand U4424 (N_4424,In_211,In_22);
nand U4425 (N_4425,In_656,In_45);
nand U4426 (N_4426,In_589,In_600);
and U4427 (N_4427,In_651,In_475);
and U4428 (N_4428,In_498,In_773);
and U4429 (N_4429,In_190,In_498);
and U4430 (N_4430,In_720,In_580);
and U4431 (N_4431,In_214,In_252);
and U4432 (N_4432,In_825,In_378);
or U4433 (N_4433,In_365,In_926);
and U4434 (N_4434,In_57,In_592);
or U4435 (N_4435,In_113,In_361);
or U4436 (N_4436,In_817,In_211);
and U4437 (N_4437,In_804,In_95);
nor U4438 (N_4438,In_822,In_210);
nand U4439 (N_4439,In_136,In_567);
nor U4440 (N_4440,In_616,In_238);
nor U4441 (N_4441,In_649,In_807);
nor U4442 (N_4442,In_650,In_202);
nand U4443 (N_4443,In_538,In_463);
or U4444 (N_4444,In_47,In_320);
nand U4445 (N_4445,In_207,In_954);
xnor U4446 (N_4446,In_511,In_105);
or U4447 (N_4447,In_447,In_40);
nand U4448 (N_4448,In_918,In_827);
and U4449 (N_4449,In_176,In_429);
or U4450 (N_4450,In_876,In_653);
nor U4451 (N_4451,In_251,In_6);
nor U4452 (N_4452,In_265,In_763);
nor U4453 (N_4453,In_443,In_881);
nor U4454 (N_4454,In_770,In_140);
nor U4455 (N_4455,In_308,In_238);
and U4456 (N_4456,In_180,In_258);
nor U4457 (N_4457,In_574,In_180);
nor U4458 (N_4458,In_616,In_188);
nand U4459 (N_4459,In_193,In_364);
or U4460 (N_4460,In_717,In_264);
nor U4461 (N_4461,In_325,In_197);
and U4462 (N_4462,In_322,In_811);
and U4463 (N_4463,In_35,In_88);
and U4464 (N_4464,In_700,In_156);
and U4465 (N_4465,In_826,In_777);
nor U4466 (N_4466,In_945,In_616);
nand U4467 (N_4467,In_429,In_966);
and U4468 (N_4468,In_955,In_592);
nand U4469 (N_4469,In_884,In_291);
and U4470 (N_4470,In_438,In_728);
nand U4471 (N_4471,In_610,In_754);
and U4472 (N_4472,In_722,In_829);
or U4473 (N_4473,In_951,In_930);
and U4474 (N_4474,In_77,In_545);
or U4475 (N_4475,In_952,In_5);
nor U4476 (N_4476,In_628,In_466);
or U4477 (N_4477,In_527,In_691);
nor U4478 (N_4478,In_581,In_20);
or U4479 (N_4479,In_392,In_688);
and U4480 (N_4480,In_332,In_243);
nand U4481 (N_4481,In_518,In_702);
nand U4482 (N_4482,In_294,In_686);
or U4483 (N_4483,In_429,In_446);
and U4484 (N_4484,In_51,In_452);
nor U4485 (N_4485,In_704,In_356);
nand U4486 (N_4486,In_154,In_524);
or U4487 (N_4487,In_242,In_741);
nand U4488 (N_4488,In_347,In_692);
and U4489 (N_4489,In_326,In_718);
and U4490 (N_4490,In_696,In_52);
xor U4491 (N_4491,In_116,In_496);
nand U4492 (N_4492,In_31,In_949);
nand U4493 (N_4493,In_946,In_907);
xnor U4494 (N_4494,In_102,In_182);
nor U4495 (N_4495,In_958,In_549);
nand U4496 (N_4496,In_290,In_350);
or U4497 (N_4497,In_670,In_677);
nor U4498 (N_4498,In_580,In_793);
and U4499 (N_4499,In_201,In_35);
nand U4500 (N_4500,In_650,In_851);
nor U4501 (N_4501,In_558,In_834);
or U4502 (N_4502,In_673,In_912);
or U4503 (N_4503,In_750,In_727);
or U4504 (N_4504,In_676,In_56);
or U4505 (N_4505,In_17,In_946);
and U4506 (N_4506,In_232,In_337);
nand U4507 (N_4507,In_662,In_611);
and U4508 (N_4508,In_670,In_264);
and U4509 (N_4509,In_96,In_419);
and U4510 (N_4510,In_975,In_158);
or U4511 (N_4511,In_446,In_997);
and U4512 (N_4512,In_49,In_837);
nand U4513 (N_4513,In_600,In_495);
or U4514 (N_4514,In_178,In_537);
or U4515 (N_4515,In_390,In_396);
nor U4516 (N_4516,In_183,In_272);
or U4517 (N_4517,In_183,In_479);
and U4518 (N_4518,In_83,In_519);
nand U4519 (N_4519,In_543,In_121);
nor U4520 (N_4520,In_529,In_368);
or U4521 (N_4521,In_570,In_875);
or U4522 (N_4522,In_627,In_509);
nor U4523 (N_4523,In_737,In_795);
nand U4524 (N_4524,In_382,In_149);
nor U4525 (N_4525,In_612,In_204);
nor U4526 (N_4526,In_374,In_376);
and U4527 (N_4527,In_434,In_632);
nand U4528 (N_4528,In_167,In_847);
nand U4529 (N_4529,In_271,In_900);
or U4530 (N_4530,In_438,In_231);
nand U4531 (N_4531,In_446,In_219);
nand U4532 (N_4532,In_299,In_147);
nand U4533 (N_4533,In_761,In_309);
or U4534 (N_4534,In_391,In_953);
nor U4535 (N_4535,In_969,In_340);
nand U4536 (N_4536,In_337,In_135);
and U4537 (N_4537,In_596,In_833);
and U4538 (N_4538,In_666,In_68);
nor U4539 (N_4539,In_11,In_146);
nor U4540 (N_4540,In_102,In_988);
nor U4541 (N_4541,In_625,In_689);
or U4542 (N_4542,In_185,In_392);
or U4543 (N_4543,In_131,In_772);
or U4544 (N_4544,In_246,In_474);
nand U4545 (N_4545,In_142,In_472);
nor U4546 (N_4546,In_840,In_704);
nand U4547 (N_4547,In_183,In_898);
and U4548 (N_4548,In_781,In_798);
or U4549 (N_4549,In_267,In_299);
nand U4550 (N_4550,In_116,In_726);
or U4551 (N_4551,In_44,In_825);
nor U4552 (N_4552,In_598,In_619);
nand U4553 (N_4553,In_913,In_975);
or U4554 (N_4554,In_973,In_19);
nand U4555 (N_4555,In_926,In_912);
or U4556 (N_4556,In_333,In_286);
and U4557 (N_4557,In_728,In_683);
nand U4558 (N_4558,In_433,In_192);
nand U4559 (N_4559,In_500,In_296);
nand U4560 (N_4560,In_197,In_944);
or U4561 (N_4561,In_563,In_721);
nand U4562 (N_4562,In_181,In_135);
nor U4563 (N_4563,In_445,In_371);
nand U4564 (N_4564,In_197,In_179);
and U4565 (N_4565,In_708,In_671);
nand U4566 (N_4566,In_919,In_990);
nand U4567 (N_4567,In_474,In_67);
and U4568 (N_4568,In_383,In_636);
and U4569 (N_4569,In_638,In_237);
nand U4570 (N_4570,In_521,In_604);
or U4571 (N_4571,In_220,In_180);
nand U4572 (N_4572,In_931,In_641);
nand U4573 (N_4573,In_907,In_57);
or U4574 (N_4574,In_692,In_109);
xor U4575 (N_4575,In_262,In_236);
nand U4576 (N_4576,In_874,In_602);
and U4577 (N_4577,In_512,In_947);
and U4578 (N_4578,In_991,In_687);
or U4579 (N_4579,In_587,In_725);
and U4580 (N_4580,In_860,In_963);
and U4581 (N_4581,In_665,In_109);
nor U4582 (N_4582,In_939,In_159);
and U4583 (N_4583,In_855,In_680);
or U4584 (N_4584,In_132,In_146);
or U4585 (N_4585,In_947,In_465);
nand U4586 (N_4586,In_363,In_189);
nand U4587 (N_4587,In_541,In_821);
or U4588 (N_4588,In_427,In_882);
or U4589 (N_4589,In_227,In_6);
nand U4590 (N_4590,In_340,In_846);
nand U4591 (N_4591,In_784,In_664);
and U4592 (N_4592,In_954,In_245);
or U4593 (N_4593,In_170,In_57);
nand U4594 (N_4594,In_320,In_376);
nor U4595 (N_4595,In_961,In_328);
and U4596 (N_4596,In_962,In_23);
nor U4597 (N_4597,In_312,In_211);
and U4598 (N_4598,In_94,In_318);
nand U4599 (N_4599,In_404,In_79);
nor U4600 (N_4600,In_676,In_489);
and U4601 (N_4601,In_880,In_398);
or U4602 (N_4602,In_156,In_880);
nand U4603 (N_4603,In_787,In_632);
or U4604 (N_4604,In_269,In_848);
nand U4605 (N_4605,In_10,In_566);
and U4606 (N_4606,In_38,In_447);
nand U4607 (N_4607,In_312,In_372);
or U4608 (N_4608,In_168,In_328);
nor U4609 (N_4609,In_955,In_238);
or U4610 (N_4610,In_808,In_30);
nor U4611 (N_4611,In_426,In_902);
and U4612 (N_4612,In_293,In_162);
or U4613 (N_4613,In_413,In_171);
nor U4614 (N_4614,In_962,In_561);
or U4615 (N_4615,In_140,In_686);
nor U4616 (N_4616,In_383,In_492);
and U4617 (N_4617,In_981,In_551);
or U4618 (N_4618,In_206,In_891);
nand U4619 (N_4619,In_629,In_389);
nand U4620 (N_4620,In_650,In_228);
nand U4621 (N_4621,In_832,In_909);
and U4622 (N_4622,In_529,In_61);
or U4623 (N_4623,In_287,In_17);
or U4624 (N_4624,In_876,In_797);
or U4625 (N_4625,In_520,In_665);
and U4626 (N_4626,In_62,In_533);
and U4627 (N_4627,In_120,In_942);
nand U4628 (N_4628,In_364,In_541);
nand U4629 (N_4629,In_880,In_396);
and U4630 (N_4630,In_426,In_679);
nor U4631 (N_4631,In_607,In_485);
and U4632 (N_4632,In_171,In_567);
nor U4633 (N_4633,In_929,In_243);
nor U4634 (N_4634,In_381,In_127);
and U4635 (N_4635,In_729,In_139);
nor U4636 (N_4636,In_391,In_49);
nand U4637 (N_4637,In_299,In_157);
or U4638 (N_4638,In_676,In_274);
or U4639 (N_4639,In_926,In_665);
nand U4640 (N_4640,In_430,In_896);
nand U4641 (N_4641,In_78,In_824);
and U4642 (N_4642,In_860,In_581);
or U4643 (N_4643,In_605,In_198);
or U4644 (N_4644,In_29,In_215);
nand U4645 (N_4645,In_523,In_408);
or U4646 (N_4646,In_871,In_453);
or U4647 (N_4647,In_922,In_616);
nand U4648 (N_4648,In_192,In_818);
nor U4649 (N_4649,In_28,In_245);
or U4650 (N_4650,In_78,In_904);
nand U4651 (N_4651,In_501,In_336);
or U4652 (N_4652,In_308,In_475);
or U4653 (N_4653,In_842,In_458);
or U4654 (N_4654,In_450,In_753);
and U4655 (N_4655,In_187,In_573);
nor U4656 (N_4656,In_45,In_804);
nand U4657 (N_4657,In_96,In_531);
or U4658 (N_4658,In_186,In_150);
nor U4659 (N_4659,In_281,In_670);
and U4660 (N_4660,In_619,In_552);
nor U4661 (N_4661,In_213,In_327);
or U4662 (N_4662,In_978,In_760);
and U4663 (N_4663,In_486,In_943);
and U4664 (N_4664,In_33,In_566);
and U4665 (N_4665,In_143,In_720);
nand U4666 (N_4666,In_428,In_131);
nand U4667 (N_4667,In_939,In_746);
nor U4668 (N_4668,In_55,In_178);
nor U4669 (N_4669,In_980,In_978);
xor U4670 (N_4670,In_561,In_474);
or U4671 (N_4671,In_375,In_578);
nor U4672 (N_4672,In_777,In_628);
nor U4673 (N_4673,In_933,In_887);
nor U4674 (N_4674,In_748,In_572);
nor U4675 (N_4675,In_507,In_528);
and U4676 (N_4676,In_480,In_800);
nand U4677 (N_4677,In_449,In_25);
and U4678 (N_4678,In_453,In_383);
nand U4679 (N_4679,In_183,In_357);
nand U4680 (N_4680,In_355,In_631);
or U4681 (N_4681,In_610,In_890);
nor U4682 (N_4682,In_340,In_751);
nor U4683 (N_4683,In_792,In_530);
or U4684 (N_4684,In_785,In_819);
and U4685 (N_4685,In_349,In_492);
nor U4686 (N_4686,In_102,In_963);
and U4687 (N_4687,In_465,In_655);
nand U4688 (N_4688,In_362,In_961);
nand U4689 (N_4689,In_529,In_331);
or U4690 (N_4690,In_935,In_909);
nor U4691 (N_4691,In_363,In_466);
nor U4692 (N_4692,In_366,In_344);
and U4693 (N_4693,In_329,In_722);
or U4694 (N_4694,In_867,In_858);
nand U4695 (N_4695,In_796,In_389);
and U4696 (N_4696,In_950,In_674);
nand U4697 (N_4697,In_194,In_708);
or U4698 (N_4698,In_249,In_396);
or U4699 (N_4699,In_429,In_45);
and U4700 (N_4700,In_311,In_5);
and U4701 (N_4701,In_496,In_230);
and U4702 (N_4702,In_974,In_277);
nand U4703 (N_4703,In_474,In_228);
or U4704 (N_4704,In_619,In_850);
nor U4705 (N_4705,In_423,In_273);
and U4706 (N_4706,In_271,In_882);
nor U4707 (N_4707,In_67,In_398);
nor U4708 (N_4708,In_339,In_431);
and U4709 (N_4709,In_597,In_18);
nor U4710 (N_4710,In_71,In_331);
or U4711 (N_4711,In_459,In_828);
nor U4712 (N_4712,In_337,In_51);
nor U4713 (N_4713,In_312,In_24);
nor U4714 (N_4714,In_751,In_399);
xor U4715 (N_4715,In_25,In_276);
nor U4716 (N_4716,In_763,In_544);
or U4717 (N_4717,In_948,In_979);
and U4718 (N_4718,In_595,In_505);
nand U4719 (N_4719,In_647,In_893);
or U4720 (N_4720,In_370,In_839);
nand U4721 (N_4721,In_546,In_988);
nor U4722 (N_4722,In_462,In_280);
nand U4723 (N_4723,In_841,In_859);
nand U4724 (N_4724,In_433,In_582);
or U4725 (N_4725,In_812,In_150);
nor U4726 (N_4726,In_927,In_313);
nor U4727 (N_4727,In_522,In_949);
nand U4728 (N_4728,In_254,In_0);
or U4729 (N_4729,In_403,In_254);
nand U4730 (N_4730,In_335,In_473);
and U4731 (N_4731,In_413,In_755);
and U4732 (N_4732,In_772,In_988);
nor U4733 (N_4733,In_643,In_179);
nand U4734 (N_4734,In_490,In_663);
and U4735 (N_4735,In_733,In_646);
or U4736 (N_4736,In_396,In_176);
and U4737 (N_4737,In_154,In_220);
nor U4738 (N_4738,In_47,In_478);
nor U4739 (N_4739,In_264,In_764);
and U4740 (N_4740,In_569,In_785);
nand U4741 (N_4741,In_998,In_192);
nor U4742 (N_4742,In_99,In_600);
nor U4743 (N_4743,In_12,In_273);
or U4744 (N_4744,In_796,In_193);
nor U4745 (N_4745,In_388,In_864);
nor U4746 (N_4746,In_129,In_735);
or U4747 (N_4747,In_193,In_100);
nor U4748 (N_4748,In_847,In_531);
or U4749 (N_4749,In_572,In_207);
or U4750 (N_4750,In_795,In_698);
or U4751 (N_4751,In_609,In_955);
nor U4752 (N_4752,In_536,In_728);
nor U4753 (N_4753,In_434,In_346);
or U4754 (N_4754,In_71,In_74);
nand U4755 (N_4755,In_147,In_790);
or U4756 (N_4756,In_873,In_508);
nor U4757 (N_4757,In_950,In_548);
or U4758 (N_4758,In_765,In_161);
nand U4759 (N_4759,In_619,In_12);
nor U4760 (N_4760,In_215,In_578);
or U4761 (N_4761,In_723,In_296);
and U4762 (N_4762,In_997,In_389);
nand U4763 (N_4763,In_589,In_466);
and U4764 (N_4764,In_465,In_438);
nand U4765 (N_4765,In_303,In_32);
nor U4766 (N_4766,In_426,In_998);
or U4767 (N_4767,In_922,In_33);
and U4768 (N_4768,In_435,In_821);
nor U4769 (N_4769,In_163,In_939);
and U4770 (N_4770,In_607,In_256);
or U4771 (N_4771,In_105,In_917);
nor U4772 (N_4772,In_438,In_202);
or U4773 (N_4773,In_422,In_342);
or U4774 (N_4774,In_257,In_811);
nand U4775 (N_4775,In_226,In_840);
and U4776 (N_4776,In_976,In_59);
nor U4777 (N_4777,In_871,In_185);
nor U4778 (N_4778,In_830,In_645);
or U4779 (N_4779,In_378,In_359);
or U4780 (N_4780,In_490,In_803);
or U4781 (N_4781,In_984,In_679);
or U4782 (N_4782,In_275,In_796);
or U4783 (N_4783,In_220,In_870);
and U4784 (N_4784,In_90,In_742);
nor U4785 (N_4785,In_301,In_991);
xnor U4786 (N_4786,In_49,In_656);
nor U4787 (N_4787,In_109,In_288);
and U4788 (N_4788,In_565,In_583);
nand U4789 (N_4789,In_484,In_209);
or U4790 (N_4790,In_905,In_105);
nand U4791 (N_4791,In_507,In_634);
nand U4792 (N_4792,In_533,In_631);
nand U4793 (N_4793,In_798,In_845);
nand U4794 (N_4794,In_608,In_557);
and U4795 (N_4795,In_66,In_609);
nand U4796 (N_4796,In_265,In_187);
or U4797 (N_4797,In_854,In_634);
nor U4798 (N_4798,In_254,In_552);
and U4799 (N_4799,In_609,In_893);
or U4800 (N_4800,In_970,In_744);
and U4801 (N_4801,In_603,In_352);
nor U4802 (N_4802,In_252,In_581);
or U4803 (N_4803,In_694,In_292);
nand U4804 (N_4804,In_313,In_539);
and U4805 (N_4805,In_204,In_575);
nand U4806 (N_4806,In_714,In_184);
nor U4807 (N_4807,In_670,In_528);
nand U4808 (N_4808,In_55,In_561);
nor U4809 (N_4809,In_425,In_90);
and U4810 (N_4810,In_591,In_11);
nor U4811 (N_4811,In_826,In_678);
or U4812 (N_4812,In_480,In_609);
or U4813 (N_4813,In_698,In_375);
and U4814 (N_4814,In_909,In_496);
or U4815 (N_4815,In_748,In_543);
nor U4816 (N_4816,In_860,In_441);
and U4817 (N_4817,In_515,In_982);
nand U4818 (N_4818,In_828,In_270);
and U4819 (N_4819,In_873,In_577);
and U4820 (N_4820,In_139,In_389);
nor U4821 (N_4821,In_429,In_364);
nand U4822 (N_4822,In_835,In_330);
xnor U4823 (N_4823,In_406,In_561);
nand U4824 (N_4824,In_706,In_425);
or U4825 (N_4825,In_879,In_396);
nand U4826 (N_4826,In_669,In_394);
and U4827 (N_4827,In_469,In_552);
or U4828 (N_4828,In_848,In_928);
nor U4829 (N_4829,In_551,In_315);
or U4830 (N_4830,In_319,In_98);
and U4831 (N_4831,In_416,In_716);
nor U4832 (N_4832,In_910,In_711);
nand U4833 (N_4833,In_46,In_111);
or U4834 (N_4834,In_435,In_516);
nand U4835 (N_4835,In_648,In_86);
or U4836 (N_4836,In_295,In_164);
and U4837 (N_4837,In_534,In_538);
nand U4838 (N_4838,In_614,In_689);
or U4839 (N_4839,In_571,In_685);
and U4840 (N_4840,In_250,In_97);
nand U4841 (N_4841,In_683,In_352);
nor U4842 (N_4842,In_127,In_122);
nand U4843 (N_4843,In_690,In_215);
and U4844 (N_4844,In_639,In_609);
and U4845 (N_4845,In_629,In_171);
nor U4846 (N_4846,In_408,In_990);
and U4847 (N_4847,In_830,In_225);
nor U4848 (N_4848,In_611,In_363);
or U4849 (N_4849,In_260,In_590);
xor U4850 (N_4850,In_979,In_555);
nand U4851 (N_4851,In_997,In_158);
nand U4852 (N_4852,In_515,In_421);
or U4853 (N_4853,In_932,In_829);
and U4854 (N_4854,In_777,In_191);
nand U4855 (N_4855,In_980,In_663);
and U4856 (N_4856,In_921,In_75);
nor U4857 (N_4857,In_742,In_110);
nand U4858 (N_4858,In_826,In_370);
nor U4859 (N_4859,In_710,In_176);
nand U4860 (N_4860,In_455,In_865);
nor U4861 (N_4861,In_686,In_889);
and U4862 (N_4862,In_697,In_17);
nor U4863 (N_4863,In_15,In_818);
nand U4864 (N_4864,In_199,In_36);
and U4865 (N_4865,In_432,In_173);
nor U4866 (N_4866,In_576,In_122);
nor U4867 (N_4867,In_645,In_759);
or U4868 (N_4868,In_365,In_227);
nand U4869 (N_4869,In_215,In_46);
or U4870 (N_4870,In_0,In_197);
and U4871 (N_4871,In_237,In_380);
nand U4872 (N_4872,In_423,In_275);
nand U4873 (N_4873,In_791,In_190);
or U4874 (N_4874,In_510,In_555);
and U4875 (N_4875,In_35,In_491);
and U4876 (N_4876,In_649,In_384);
and U4877 (N_4877,In_600,In_222);
nand U4878 (N_4878,In_489,In_521);
and U4879 (N_4879,In_999,In_331);
or U4880 (N_4880,In_603,In_732);
nor U4881 (N_4881,In_353,In_847);
nand U4882 (N_4882,In_875,In_432);
nand U4883 (N_4883,In_486,In_476);
nor U4884 (N_4884,In_230,In_165);
nand U4885 (N_4885,In_957,In_828);
nand U4886 (N_4886,In_747,In_799);
nand U4887 (N_4887,In_334,In_102);
nand U4888 (N_4888,In_642,In_388);
nor U4889 (N_4889,In_636,In_404);
and U4890 (N_4890,In_301,In_386);
nor U4891 (N_4891,In_386,In_983);
nand U4892 (N_4892,In_45,In_539);
nand U4893 (N_4893,In_951,In_749);
nand U4894 (N_4894,In_169,In_517);
nor U4895 (N_4895,In_840,In_992);
nand U4896 (N_4896,In_9,In_994);
nand U4897 (N_4897,In_298,In_412);
xor U4898 (N_4898,In_951,In_352);
or U4899 (N_4899,In_917,In_58);
nor U4900 (N_4900,In_305,In_609);
nor U4901 (N_4901,In_252,In_133);
nand U4902 (N_4902,In_634,In_259);
and U4903 (N_4903,In_162,In_732);
nor U4904 (N_4904,In_250,In_904);
or U4905 (N_4905,In_438,In_143);
and U4906 (N_4906,In_207,In_897);
or U4907 (N_4907,In_21,In_794);
or U4908 (N_4908,In_12,In_846);
or U4909 (N_4909,In_686,In_676);
nand U4910 (N_4910,In_403,In_570);
nor U4911 (N_4911,In_754,In_187);
nand U4912 (N_4912,In_532,In_579);
nand U4913 (N_4913,In_823,In_717);
and U4914 (N_4914,In_259,In_672);
or U4915 (N_4915,In_723,In_412);
nor U4916 (N_4916,In_335,In_532);
or U4917 (N_4917,In_840,In_455);
nand U4918 (N_4918,In_763,In_229);
nand U4919 (N_4919,In_855,In_235);
or U4920 (N_4920,In_98,In_866);
or U4921 (N_4921,In_432,In_648);
or U4922 (N_4922,In_693,In_652);
or U4923 (N_4923,In_754,In_216);
or U4924 (N_4924,In_996,In_552);
nor U4925 (N_4925,In_610,In_118);
and U4926 (N_4926,In_926,In_443);
or U4927 (N_4927,In_300,In_562);
nor U4928 (N_4928,In_78,In_410);
or U4929 (N_4929,In_275,In_799);
and U4930 (N_4930,In_179,In_42);
nand U4931 (N_4931,In_353,In_948);
nor U4932 (N_4932,In_798,In_150);
nor U4933 (N_4933,In_885,In_528);
nand U4934 (N_4934,In_165,In_705);
nand U4935 (N_4935,In_777,In_993);
nand U4936 (N_4936,In_562,In_29);
and U4937 (N_4937,In_278,In_800);
nand U4938 (N_4938,In_562,In_841);
nand U4939 (N_4939,In_37,In_483);
or U4940 (N_4940,In_273,In_917);
nand U4941 (N_4941,In_77,In_827);
and U4942 (N_4942,In_784,In_21);
nor U4943 (N_4943,In_72,In_894);
nand U4944 (N_4944,In_928,In_346);
nor U4945 (N_4945,In_738,In_374);
or U4946 (N_4946,In_532,In_855);
nand U4947 (N_4947,In_334,In_435);
nand U4948 (N_4948,In_311,In_892);
or U4949 (N_4949,In_149,In_543);
nor U4950 (N_4950,In_684,In_444);
nand U4951 (N_4951,In_482,In_44);
nor U4952 (N_4952,In_169,In_580);
and U4953 (N_4953,In_682,In_999);
nand U4954 (N_4954,In_121,In_771);
or U4955 (N_4955,In_254,In_682);
nand U4956 (N_4956,In_47,In_336);
nor U4957 (N_4957,In_222,In_383);
nand U4958 (N_4958,In_329,In_835);
nor U4959 (N_4959,In_817,In_827);
or U4960 (N_4960,In_182,In_494);
nand U4961 (N_4961,In_67,In_293);
and U4962 (N_4962,In_927,In_81);
nor U4963 (N_4963,In_220,In_775);
nor U4964 (N_4964,In_234,In_671);
and U4965 (N_4965,In_148,In_459);
and U4966 (N_4966,In_96,In_68);
nand U4967 (N_4967,In_189,In_933);
nand U4968 (N_4968,In_81,In_342);
and U4969 (N_4969,In_760,In_36);
and U4970 (N_4970,In_799,In_37);
and U4971 (N_4971,In_866,In_540);
or U4972 (N_4972,In_667,In_42);
nand U4973 (N_4973,In_181,In_396);
and U4974 (N_4974,In_301,In_291);
or U4975 (N_4975,In_276,In_473);
and U4976 (N_4976,In_631,In_930);
or U4977 (N_4977,In_907,In_500);
and U4978 (N_4978,In_324,In_762);
and U4979 (N_4979,In_176,In_860);
or U4980 (N_4980,In_232,In_244);
nor U4981 (N_4981,In_510,In_659);
nor U4982 (N_4982,In_39,In_177);
and U4983 (N_4983,In_556,In_188);
and U4984 (N_4984,In_711,In_417);
or U4985 (N_4985,In_751,In_623);
nand U4986 (N_4986,In_368,In_992);
and U4987 (N_4987,In_652,In_985);
xor U4988 (N_4988,In_211,In_119);
nand U4989 (N_4989,In_788,In_115);
nand U4990 (N_4990,In_232,In_804);
or U4991 (N_4991,In_517,In_590);
nor U4992 (N_4992,In_468,In_455);
nor U4993 (N_4993,In_853,In_121);
nor U4994 (N_4994,In_542,In_912);
nand U4995 (N_4995,In_706,In_346);
nand U4996 (N_4996,In_74,In_460);
nor U4997 (N_4997,In_247,In_965);
and U4998 (N_4998,In_38,In_219);
nor U4999 (N_4999,In_216,In_202);
nor U5000 (N_5000,N_1903,N_3246);
or U5001 (N_5001,N_1931,N_1361);
nor U5002 (N_5002,N_89,N_2284);
nor U5003 (N_5003,N_1441,N_1249);
nand U5004 (N_5004,N_2881,N_3131);
nor U5005 (N_5005,N_240,N_3224);
or U5006 (N_5006,N_787,N_1723);
nand U5007 (N_5007,N_3718,N_1474);
nor U5008 (N_5008,N_2750,N_3440);
nand U5009 (N_5009,N_4436,N_4019);
or U5010 (N_5010,N_1707,N_4013);
nor U5011 (N_5011,N_2829,N_2594);
and U5012 (N_5012,N_863,N_3400);
or U5013 (N_5013,N_4171,N_2591);
and U5014 (N_5014,N_1025,N_2158);
or U5015 (N_5015,N_3782,N_188);
nor U5016 (N_5016,N_1711,N_1468);
nor U5017 (N_5017,N_231,N_1447);
or U5018 (N_5018,N_1505,N_2491);
nor U5019 (N_5019,N_1771,N_2804);
or U5020 (N_5020,N_4094,N_3203);
or U5021 (N_5021,N_3880,N_3466);
or U5022 (N_5022,N_1504,N_3682);
and U5023 (N_5023,N_3204,N_3567);
and U5024 (N_5024,N_4916,N_879);
or U5025 (N_5025,N_4023,N_2508);
and U5026 (N_5026,N_1416,N_1498);
nand U5027 (N_5027,N_207,N_3458);
or U5028 (N_5028,N_1642,N_2730);
or U5029 (N_5029,N_3256,N_2724);
nor U5030 (N_5030,N_1794,N_2552);
nor U5031 (N_5031,N_294,N_4361);
nor U5032 (N_5032,N_410,N_3617);
nand U5033 (N_5033,N_4294,N_2494);
nor U5034 (N_5034,N_1158,N_2350);
nor U5035 (N_5035,N_336,N_3735);
nand U5036 (N_5036,N_1252,N_2646);
nand U5037 (N_5037,N_4342,N_4708);
nand U5038 (N_5038,N_1657,N_4351);
nor U5039 (N_5039,N_4851,N_219);
or U5040 (N_5040,N_1420,N_3401);
or U5041 (N_5041,N_4163,N_4051);
nor U5042 (N_5042,N_461,N_1896);
nor U5043 (N_5043,N_160,N_2949);
nand U5044 (N_5044,N_1933,N_4880);
nor U5045 (N_5045,N_2420,N_109);
nand U5046 (N_5046,N_407,N_1424);
or U5047 (N_5047,N_3768,N_1005);
nand U5048 (N_5048,N_1448,N_3081);
nor U5049 (N_5049,N_4096,N_1189);
nor U5050 (N_5050,N_2150,N_1577);
nor U5051 (N_5051,N_2537,N_3904);
nand U5052 (N_5052,N_2713,N_4742);
and U5053 (N_5053,N_1269,N_1180);
or U5054 (N_5054,N_419,N_3226);
nor U5055 (N_5055,N_2422,N_674);
or U5056 (N_5056,N_2014,N_1442);
nor U5057 (N_5057,N_2083,N_229);
nor U5058 (N_5058,N_3283,N_3221);
and U5059 (N_5059,N_2579,N_227);
and U5060 (N_5060,N_115,N_803);
or U5061 (N_5061,N_1899,N_596);
or U5062 (N_5062,N_4828,N_871);
nand U5063 (N_5063,N_3158,N_3824);
or U5064 (N_5064,N_4634,N_712);
nor U5065 (N_5065,N_217,N_4568);
or U5066 (N_5066,N_2868,N_127);
nand U5067 (N_5067,N_466,N_1321);
nand U5068 (N_5068,N_3045,N_1220);
nand U5069 (N_5069,N_4554,N_2462);
nand U5070 (N_5070,N_59,N_2186);
nand U5071 (N_5071,N_4795,N_4335);
or U5072 (N_5072,N_134,N_3233);
nand U5073 (N_5073,N_626,N_800);
and U5074 (N_5074,N_3909,N_3223);
and U5075 (N_5075,N_282,N_1678);
nand U5076 (N_5076,N_4036,N_1060);
nor U5077 (N_5077,N_4228,N_1592);
and U5078 (N_5078,N_86,N_4856);
or U5079 (N_5079,N_776,N_4319);
and U5080 (N_5080,N_356,N_431);
or U5081 (N_5081,N_85,N_4355);
nand U5082 (N_5082,N_3004,N_1847);
nand U5083 (N_5083,N_4627,N_301);
and U5084 (N_5084,N_1417,N_1966);
or U5085 (N_5085,N_4133,N_2662);
nor U5086 (N_5086,N_4901,N_2453);
or U5087 (N_5087,N_3635,N_1101);
nor U5088 (N_5088,N_1013,N_4989);
or U5089 (N_5089,N_1664,N_2139);
nand U5090 (N_5090,N_3054,N_4276);
and U5091 (N_5091,N_2020,N_2529);
and U5092 (N_5092,N_3157,N_167);
nand U5093 (N_5093,N_1273,N_4960);
nand U5094 (N_5094,N_3385,N_4605);
and U5095 (N_5095,N_3842,N_84);
and U5096 (N_5096,N_1431,N_324);
or U5097 (N_5097,N_3036,N_4267);
and U5098 (N_5098,N_4101,N_1079);
nor U5099 (N_5099,N_3310,N_525);
or U5100 (N_5100,N_2893,N_1725);
or U5101 (N_5101,N_552,N_2262);
and U5102 (N_5102,N_4273,N_572);
and U5103 (N_5103,N_1936,N_4058);
nor U5104 (N_5104,N_2137,N_2919);
nor U5105 (N_5105,N_2401,N_2482);
and U5106 (N_5106,N_2866,N_1405);
or U5107 (N_5107,N_4277,N_715);
or U5108 (N_5108,N_3423,N_3738);
or U5109 (N_5109,N_3926,N_4701);
and U5110 (N_5110,N_1579,N_2228);
and U5111 (N_5111,N_3701,N_4069);
nand U5112 (N_5112,N_4486,N_2709);
and U5113 (N_5113,N_1885,N_3882);
nand U5114 (N_5114,N_3492,N_1700);
nor U5115 (N_5115,N_4813,N_4849);
and U5116 (N_5116,N_930,N_2680);
or U5117 (N_5117,N_112,N_1716);
or U5118 (N_5118,N_4656,N_2564);
and U5119 (N_5119,N_2864,N_3832);
nor U5120 (N_5120,N_2530,N_1715);
or U5121 (N_5121,N_2695,N_4295);
and U5122 (N_5122,N_295,N_145);
nand U5123 (N_5123,N_3202,N_1280);
nor U5124 (N_5124,N_1258,N_4979);
or U5125 (N_5125,N_429,N_97);
nor U5126 (N_5126,N_178,N_424);
nand U5127 (N_5127,N_1726,N_328);
nand U5128 (N_5128,N_4384,N_3912);
nor U5129 (N_5129,N_3424,N_1375);
nand U5130 (N_5130,N_548,N_1257);
nor U5131 (N_5131,N_3756,N_184);
nand U5132 (N_5132,N_4289,N_1337);
nand U5133 (N_5133,N_1821,N_1752);
nor U5134 (N_5134,N_508,N_4819);
nand U5135 (N_5135,N_2025,N_1215);
nor U5136 (N_5136,N_281,N_3497);
or U5137 (N_5137,N_1502,N_2369);
and U5138 (N_5138,N_447,N_1155);
or U5139 (N_5139,N_3811,N_3176);
nor U5140 (N_5140,N_3116,N_1322);
and U5141 (N_5141,N_981,N_1962);
and U5142 (N_5142,N_3625,N_3931);
xor U5143 (N_5143,N_4688,N_4877);
or U5144 (N_5144,N_2792,N_4549);
or U5145 (N_5145,N_4443,N_2843);
nand U5146 (N_5146,N_107,N_4553);
or U5147 (N_5147,N_2555,N_1440);
nor U5148 (N_5148,N_4952,N_4760);
nand U5149 (N_5149,N_1113,N_4496);
or U5150 (N_5150,N_3080,N_609);
or U5151 (N_5151,N_3667,N_3935);
and U5152 (N_5152,N_1069,N_1747);
nor U5153 (N_5153,N_259,N_4662);
nand U5154 (N_5154,N_3582,N_1225);
or U5155 (N_5155,N_3925,N_1839);
nand U5156 (N_5156,N_1953,N_149);
or U5157 (N_5157,N_619,N_2069);
nor U5158 (N_5158,N_4946,N_4690);
nand U5159 (N_5159,N_4420,N_1412);
or U5160 (N_5160,N_3345,N_1232);
and U5161 (N_5161,N_397,N_4558);
nor U5162 (N_5162,N_755,N_116);
nor U5163 (N_5163,N_1944,N_1500);
and U5164 (N_5164,N_2965,N_658);
or U5165 (N_5165,N_1414,N_3971);
and U5166 (N_5166,N_2712,N_1218);
nand U5167 (N_5167,N_4056,N_213);
nor U5168 (N_5168,N_2610,N_278);
and U5169 (N_5169,N_1951,N_3094);
or U5170 (N_5170,N_3957,N_3329);
or U5171 (N_5171,N_1087,N_4640);
nor U5172 (N_5172,N_2970,N_4291);
and U5173 (N_5173,N_2585,N_1516);
or U5174 (N_5174,N_2549,N_1928);
nand U5175 (N_5175,N_2280,N_2227);
nor U5176 (N_5176,N_40,N_3941);
nor U5177 (N_5177,N_4279,N_1179);
nand U5178 (N_5178,N_2683,N_214);
or U5179 (N_5179,N_3416,N_1669);
and U5180 (N_5180,N_1539,N_3337);
and U5181 (N_5181,N_2716,N_1254);
or U5182 (N_5182,N_2012,N_2523);
nand U5183 (N_5183,N_1305,N_4249);
or U5184 (N_5184,N_2539,N_1476);
and U5185 (N_5185,N_762,N_2272);
nand U5186 (N_5186,N_2909,N_2456);
nand U5187 (N_5187,N_2455,N_2982);
nand U5188 (N_5188,N_3343,N_3247);
and U5189 (N_5189,N_3560,N_2116);
and U5190 (N_5190,N_4261,N_3676);
and U5191 (N_5191,N_4073,N_4933);
or U5192 (N_5192,N_2247,N_81);
nor U5193 (N_5193,N_2106,N_3733);
nor U5194 (N_5194,N_3829,N_962);
or U5195 (N_5195,N_3243,N_3408);
nand U5196 (N_5196,N_4323,N_3496);
nor U5197 (N_5197,N_2432,N_2659);
and U5198 (N_5198,N_15,N_4868);
nor U5199 (N_5199,N_669,N_2205);
and U5200 (N_5200,N_943,N_4812);
or U5201 (N_5201,N_665,N_1120);
nand U5202 (N_5202,N_2723,N_1331);
nor U5203 (N_5203,N_2480,N_2830);
and U5204 (N_5204,N_2583,N_4292);
and U5205 (N_5205,N_4244,N_1996);
and U5206 (N_5206,N_3927,N_858);
nor U5207 (N_5207,N_492,N_2254);
and U5208 (N_5208,N_2080,N_4610);
or U5209 (N_5209,N_3579,N_1051);
nor U5210 (N_5210,N_443,N_2055);
and U5211 (N_5211,N_1908,N_2711);
nor U5212 (N_5212,N_2404,N_1840);
and U5213 (N_5213,N_1346,N_1197);
and U5214 (N_5214,N_262,N_4922);
and U5215 (N_5215,N_2923,N_1365);
or U5216 (N_5216,N_521,N_3569);
and U5217 (N_5217,N_242,N_2620);
or U5218 (N_5218,N_960,N_2877);
and U5219 (N_5219,N_3818,N_3961);
and U5220 (N_5220,N_4334,N_361);
nand U5221 (N_5221,N_3198,N_2327);
nand U5222 (N_5222,N_1981,N_4108);
nor U5223 (N_5223,N_460,N_1595);
or U5224 (N_5224,N_1522,N_1226);
or U5225 (N_5225,N_523,N_733);
nor U5226 (N_5226,N_877,N_4955);
or U5227 (N_5227,N_3553,N_1391);
nor U5228 (N_5228,N_3786,N_2112);
and U5229 (N_5229,N_604,N_2439);
nand U5230 (N_5230,N_1047,N_4571);
or U5231 (N_5231,N_2990,N_95);
nor U5232 (N_5232,N_4214,N_1682);
nor U5233 (N_5233,N_1761,N_1278);
nor U5234 (N_5234,N_4798,N_2486);
nor U5235 (N_5235,N_567,N_4042);
nand U5236 (N_5236,N_3373,N_3140);
xnor U5237 (N_5237,N_4944,N_352);
or U5238 (N_5238,N_2047,N_865);
and U5239 (N_5239,N_854,N_4521);
nand U5240 (N_5240,N_285,N_3041);
or U5241 (N_5241,N_2999,N_1401);
nand U5242 (N_5242,N_4642,N_1755);
and U5243 (N_5243,N_4879,N_3911);
or U5244 (N_5244,N_1181,N_3259);
nand U5245 (N_5245,N_847,N_3231);
or U5246 (N_5246,N_3845,N_2136);
or U5247 (N_5247,N_1541,N_2110);
nor U5248 (N_5248,N_3788,N_3673);
nand U5249 (N_5249,N_3210,N_3420);
and U5250 (N_5250,N_4647,N_4839);
and U5251 (N_5251,N_4583,N_4387);
nand U5252 (N_5252,N_2461,N_351);
and U5253 (N_5253,N_1061,N_4200);
xnor U5254 (N_5254,N_4009,N_885);
and U5255 (N_5255,N_2253,N_4744);
and U5256 (N_5256,N_3550,N_4485);
and U5257 (N_5257,N_3196,N_3264);
nand U5258 (N_5258,N_1817,N_1709);
or U5259 (N_5259,N_1778,N_897);
and U5260 (N_5260,N_3775,N_3908);
nor U5261 (N_5261,N_946,N_4413);
and U5262 (N_5262,N_4587,N_3009);
nor U5263 (N_5263,N_3532,N_3901);
nor U5264 (N_5264,N_2140,N_3294);
nand U5265 (N_5265,N_3787,N_2478);
nor U5266 (N_5266,N_103,N_1708);
xor U5267 (N_5267,N_4692,N_4951);
and U5268 (N_5268,N_1014,N_717);
and U5269 (N_5269,N_914,N_264);
nand U5270 (N_5270,N_1684,N_1666);
nand U5271 (N_5271,N_4272,N_354);
nand U5272 (N_5272,N_1146,N_2890);
nor U5273 (N_5273,N_3891,N_114);
nor U5274 (N_5274,N_21,N_2785);
and U5275 (N_5275,N_2364,N_2251);
or U5276 (N_5276,N_4242,N_3557);
nand U5277 (N_5277,N_1785,N_4259);
nor U5278 (N_5278,N_1187,N_3598);
and U5279 (N_5279,N_3657,N_3519);
and U5280 (N_5280,N_26,N_3742);
and U5281 (N_5281,N_1939,N_688);
nand U5282 (N_5282,N_2650,N_3924);
nand U5283 (N_5283,N_4841,N_3499);
nand U5284 (N_5284,N_3887,N_4691);
nand U5285 (N_5285,N_2633,N_3942);
xor U5286 (N_5286,N_158,N_775);
nand U5287 (N_5287,N_2958,N_826);
or U5288 (N_5288,N_3150,N_372);
and U5289 (N_5289,N_4893,N_613);
and U5290 (N_5290,N_1395,N_4569);
or U5291 (N_5291,N_3190,N_4821);
nand U5292 (N_5292,N_317,N_3178);
and U5293 (N_5293,N_1192,N_1358);
and U5294 (N_5294,N_4198,N_1982);
nand U5295 (N_5295,N_4626,N_2943);
nand U5296 (N_5296,N_4472,N_403);
nor U5297 (N_5297,N_1970,N_248);
or U5298 (N_5298,N_866,N_2221);
nor U5299 (N_5299,N_2600,N_4546);
nor U5300 (N_5300,N_412,N_1185);
or U5301 (N_5301,N_1535,N_859);
or U5302 (N_5302,N_1864,N_3334);
nand U5303 (N_5303,N_1978,N_1347);
or U5304 (N_5304,N_1411,N_1404);
and U5305 (N_5305,N_4135,N_2840);
nand U5306 (N_5306,N_1355,N_1626);
or U5307 (N_5307,N_323,N_4537);
and U5308 (N_5308,N_3921,N_1807);
nor U5309 (N_5309,N_3252,N_4547);
and U5310 (N_5310,N_3736,N_1960);
nor U5311 (N_5311,N_3282,N_2941);
or U5312 (N_5312,N_3271,N_709);
nand U5313 (N_5313,N_3121,N_2189);
or U5314 (N_5314,N_540,N_3559);
or U5315 (N_5315,N_143,N_599);
or U5316 (N_5316,N_4739,N_3652);
nand U5317 (N_5317,N_4445,N_4687);
nand U5318 (N_5318,N_4527,N_3354);
or U5319 (N_5319,N_273,N_1388);
nand U5320 (N_5320,N_4217,N_4344);
or U5321 (N_5321,N_3197,N_2337);
nand U5322 (N_5322,N_4825,N_4697);
and U5323 (N_5323,N_901,N_3762);
xor U5324 (N_5324,N_3254,N_4914);
nor U5325 (N_5325,N_1268,N_1057);
or U5326 (N_5326,N_135,N_949);
or U5327 (N_5327,N_2073,N_1310);
nand U5328 (N_5328,N_3285,N_3843);
nor U5329 (N_5329,N_1788,N_1428);
or U5330 (N_5330,N_100,N_4463);
nor U5331 (N_5331,N_2431,N_3867);
and U5332 (N_5332,N_3300,N_74);
nand U5333 (N_5333,N_4307,N_4514);
or U5334 (N_5334,N_2770,N_1233);
or U5335 (N_5335,N_3500,N_2312);
and U5336 (N_5336,N_1491,N_3035);
xnor U5337 (N_5337,N_4572,N_698);
and U5338 (N_5338,N_1834,N_4968);
nor U5339 (N_5339,N_4929,N_2479);
nand U5340 (N_5340,N_3633,N_2126);
or U5341 (N_5341,N_3397,N_1720);
nor U5342 (N_5342,N_627,N_1103);
or U5343 (N_5343,N_1425,N_0);
and U5344 (N_5344,N_1082,N_4453);
or U5345 (N_5345,N_4047,N_4579);
nand U5346 (N_5346,N_4790,N_697);
nand U5347 (N_5347,N_3093,N_2378);
nor U5348 (N_5348,N_2527,N_1674);
and U5349 (N_5349,N_759,N_844);
xor U5350 (N_5350,N_3851,N_2971);
and U5351 (N_5351,N_1703,N_2097);
nand U5352 (N_5352,N_4462,N_2295);
and U5353 (N_5353,N_504,N_3255);
and U5354 (N_5354,N_4151,N_2519);
nand U5355 (N_5355,N_1352,N_3820);
nand U5356 (N_5356,N_1067,N_764);
nor U5357 (N_5357,N_2740,N_4491);
and U5358 (N_5358,N_1940,N_4618);
or U5359 (N_5359,N_2484,N_2181);
or U5360 (N_5360,N_1887,N_802);
nand U5361 (N_5361,N_772,N_3677);
nor U5362 (N_5362,N_3215,N_4280);
nor U5363 (N_5363,N_1660,N_316);
or U5364 (N_5364,N_4076,N_3893);
and U5365 (N_5365,N_4709,N_2641);
nor U5366 (N_5366,N_3744,N_2862);
nor U5367 (N_5367,N_2836,N_3720);
nor U5368 (N_5368,N_161,N_3853);
nor U5369 (N_5369,N_1157,N_4726);
or U5370 (N_5370,N_3071,N_1315);
nand U5371 (N_5371,N_4037,N_4495);
and U5372 (N_5372,N_1594,N_3539);
or U5373 (N_5373,N_4706,N_3741);
and U5374 (N_5374,N_2123,N_3973);
and U5375 (N_5375,N_157,N_4216);
nor U5376 (N_5376,N_3881,N_2162);
nor U5377 (N_5377,N_4488,N_2744);
nor U5378 (N_5378,N_1547,N_2976);
nor U5379 (N_5379,N_4129,N_1478);
and U5380 (N_5380,N_83,N_2467);
or U5381 (N_5381,N_1991,N_984);
or U5382 (N_5382,N_3207,N_4003);
and U5383 (N_5383,N_747,N_1644);
and U5384 (N_5384,N_4220,N_1170);
and U5385 (N_5385,N_4949,N_2927);
and U5386 (N_5386,N_367,N_1556);
and U5387 (N_5387,N_524,N_441);
nand U5388 (N_5388,N_510,N_322);
and U5389 (N_5389,N_1208,N_770);
or U5390 (N_5390,N_1638,N_2997);
or U5391 (N_5391,N_2167,N_2034);
xor U5392 (N_5392,N_2753,N_4963);
and U5393 (N_5393,N_1177,N_656);
nand U5394 (N_5394,N_1891,N_3573);
or U5395 (N_5395,N_3449,N_4932);
nand U5396 (N_5396,N_2743,N_3534);
or U5397 (N_5397,N_3051,N_142);
or U5398 (N_5398,N_2901,N_1126);
nor U5399 (N_5399,N_1342,N_994);
or U5400 (N_5400,N_378,N_4007);
nand U5401 (N_5401,N_2225,N_2232);
and U5402 (N_5402,N_290,N_842);
nor U5403 (N_5403,N_138,N_2437);
or U5404 (N_5404,N_668,N_4562);
nor U5405 (N_5405,N_3603,N_1695);
nand U5406 (N_5406,N_4507,N_4021);
nor U5407 (N_5407,N_4847,N_2818);
nand U5408 (N_5408,N_2558,N_4753);
or U5409 (N_5409,N_4966,N_3076);
nor U5410 (N_5410,N_2627,N_1950);
nor U5411 (N_5411,N_1551,N_4196);
or U5412 (N_5412,N_4722,N_1266);
and U5413 (N_5413,N_1918,N_4550);
nand U5414 (N_5414,N_2791,N_2983);
nand U5415 (N_5415,N_4834,N_2894);
nor U5416 (N_5416,N_2592,N_4718);
nand U5417 (N_5417,N_838,N_2476);
and U5418 (N_5418,N_3444,N_2954);
and U5419 (N_5419,N_2218,N_2301);
nand U5420 (N_5420,N_695,N_4713);
and U5421 (N_5421,N_4698,N_4984);
or U5422 (N_5422,N_4000,N_4112);
or U5423 (N_5423,N_3399,N_3162);
nor U5424 (N_5424,N_833,N_1920);
nor U5425 (N_5425,N_1795,N_1035);
or U5426 (N_5426,N_4830,N_2384);
or U5427 (N_5427,N_3552,N_3570);
or U5428 (N_5428,N_58,N_700);
and U5429 (N_5429,N_1572,N_128);
nor U5430 (N_5430,N_1670,N_677);
nand U5431 (N_5431,N_3126,N_3984);
nor U5432 (N_5432,N_177,N_2386);
or U5433 (N_5433,N_1650,N_333);
nand U5434 (N_5434,N_3377,N_2967);
nor U5435 (N_5435,N_2664,N_4417);
nor U5436 (N_5436,N_3689,N_3546);
or U5437 (N_5437,N_4663,N_2155);
nor U5438 (N_5438,N_55,N_2147);
nand U5439 (N_5439,N_2538,N_202);
nand U5440 (N_5440,N_2,N_181);
nand U5441 (N_5441,N_2813,N_848);
nand U5442 (N_5442,N_3755,N_1446);
nor U5443 (N_5443,N_4365,N_4065);
and U5444 (N_5444,N_2336,N_487);
nand U5445 (N_5445,N_4325,N_3043);
or U5446 (N_5446,N_3623,N_4150);
or U5447 (N_5447,N_4318,N_4137);
or U5448 (N_5448,N_1086,N_3186);
or U5449 (N_5449,N_3459,N_1729);
or U5450 (N_5450,N_3413,N_3425);
xor U5451 (N_5451,N_4937,N_3543);
nand U5452 (N_5452,N_2371,N_2669);
nor U5453 (N_5453,N_851,N_2059);
and U5454 (N_5454,N_1130,N_4777);
xnor U5455 (N_5455,N_1152,N_1032);
nand U5456 (N_5456,N_3305,N_2939);
nand U5457 (N_5457,N_1493,N_4449);
nand U5458 (N_5458,N_3075,N_4107);
and U5459 (N_5459,N_391,N_4719);
nor U5460 (N_5460,N_4016,N_3236);
nand U5461 (N_5461,N_3312,N_4349);
and U5462 (N_5462,N_4039,N_2636);
nor U5463 (N_5463,N_3019,N_4589);
or U5464 (N_5464,N_1314,N_2255);
nor U5465 (N_5465,N_3618,N_4014);
or U5466 (N_5466,N_2062,N_1076);
nor U5467 (N_5467,N_4404,N_902);
nand U5468 (N_5468,N_3751,N_2267);
nor U5469 (N_5469,N_4981,N_2790);
or U5470 (N_5470,N_2496,N_512);
nand U5471 (N_5471,N_3794,N_3042);
nand U5472 (N_5472,N_2729,N_603);
nor U5473 (N_5473,N_3947,N_4164);
or U5474 (N_5474,N_3350,N_2768);
and U5475 (N_5475,N_1031,N_1290);
and U5476 (N_5476,N_2512,N_2417);
nand U5477 (N_5477,N_254,N_2865);
nor U5478 (N_5478,N_1183,N_4664);
and U5479 (N_5479,N_4985,N_435);
nand U5480 (N_5480,N_3149,N_276);
or U5481 (N_5481,N_279,N_452);
nand U5482 (N_5482,N_434,N_1073);
nand U5483 (N_5483,N_3873,N_225);
or U5484 (N_5484,N_31,N_1160);
and U5485 (N_5485,N_4675,N_3778);
or U5486 (N_5486,N_2407,N_3658);
nand U5487 (N_5487,N_1880,N_2859);
nand U5488 (N_5488,N_3545,N_910);
and U5489 (N_5489,N_988,N_3316);
and U5490 (N_5490,N_4755,N_2427);
nand U5491 (N_5491,N_2075,N_3722);
or U5492 (N_5492,N_4820,N_1721);
nor U5493 (N_5493,N_4805,N_3711);
or U5494 (N_5494,N_190,N_1033);
and U5495 (N_5495,N_2929,N_60);
or U5496 (N_5496,N_4155,N_4165);
nor U5497 (N_5497,N_1117,N_4874);
and U5498 (N_5498,N_1780,N_2634);
nor U5499 (N_5499,N_4103,N_2978);
nor U5500 (N_5500,N_3273,N_1520);
and U5501 (N_5501,N_4211,N_1270);
or U5502 (N_5502,N_195,N_267);
and U5503 (N_5503,N_88,N_2194);
nor U5504 (N_5504,N_2614,N_4157);
nor U5505 (N_5505,N_3206,N_3478);
and U5506 (N_5506,N_4237,N_1833);
nand U5507 (N_5507,N_1050,N_3796);
nand U5508 (N_5508,N_3592,N_2143);
or U5509 (N_5509,N_1814,N_1599);
and U5510 (N_5510,N_1873,N_2067);
and U5511 (N_5511,N_2060,N_3781);
nor U5512 (N_5512,N_3367,N_2164);
or U5513 (N_5513,N_1770,N_3322);
and U5514 (N_5514,N_825,N_2044);
nand U5515 (N_5515,N_4850,N_2951);
or U5516 (N_5516,N_2756,N_3584);
or U5517 (N_5517,N_1932,N_30);
nor U5518 (N_5518,N_1749,N_1859);
and U5519 (N_5519,N_986,N_870);
or U5520 (N_5520,N_3209,N_2819);
or U5521 (N_5521,N_3078,N_2847);
nand U5522 (N_5522,N_2735,N_2325);
nand U5523 (N_5523,N_1010,N_1161);
or U5524 (N_5524,N_3072,N_773);
nor U5525 (N_5525,N_4764,N_691);
nor U5526 (N_5526,N_163,N_1867);
or U5527 (N_5527,N_1636,N_1277);
and U5528 (N_5528,N_4831,N_3130);
nand U5529 (N_5529,N_1433,N_1717);
and U5530 (N_5530,N_1980,N_535);
or U5531 (N_5531,N_1109,N_4622);
nand U5532 (N_5532,N_482,N_2749);
nor U5533 (N_5533,N_2236,N_3089);
nand U5534 (N_5534,N_1396,N_3813);
or U5535 (N_5535,N_3619,N_1300);
and U5536 (N_5536,N_2320,N_1680);
or U5537 (N_5537,N_907,N_805);
and U5538 (N_5538,N_4077,N_4184);
and U5539 (N_5539,N_4078,N_2617);
nand U5540 (N_5540,N_1421,N_1345);
nor U5541 (N_5541,N_444,N_671);
nand U5542 (N_5542,N_221,N_2795);
or U5543 (N_5543,N_1967,N_784);
and U5544 (N_5544,N_222,N_514);
nand U5545 (N_5545,N_53,N_1376);
nor U5546 (N_5546,N_678,N_1540);
or U5547 (N_5547,N_605,N_4275);
nor U5548 (N_5548,N_211,N_1524);
nor U5549 (N_5549,N_2030,N_3378);
or U5550 (N_5550,N_4611,N_824);
nor U5551 (N_5551,N_4964,N_2430);
and U5552 (N_5552,N_152,N_1965);
or U5553 (N_5553,N_1250,N_1325);
nand U5554 (N_5554,N_1194,N_4167);
nor U5555 (N_5555,N_1746,N_3142);
nand U5556 (N_5556,N_4700,N_2065);
or U5557 (N_5557,N_1924,N_2454);
or U5558 (N_5558,N_2095,N_168);
nor U5559 (N_5559,N_1934,N_4950);
and U5560 (N_5560,N_4134,N_2979);
nor U5561 (N_5561,N_2352,N_1422);
or U5562 (N_5562,N_2245,N_3950);
and U5563 (N_5563,N_171,N_4401);
and U5564 (N_5564,N_3222,N_3684);
and U5565 (N_5565,N_2741,N_4432);
and U5566 (N_5566,N_4465,N_3366);
nor U5567 (N_5567,N_1151,N_1945);
nand U5568 (N_5568,N_740,N_331);
and U5569 (N_5569,N_4766,N_815);
or U5570 (N_5570,N_1862,N_3491);
and U5571 (N_5571,N_2809,N_2169);
nand U5572 (N_5572,N_1292,N_684);
nor U5573 (N_5573,N_4619,N_4727);
and U5574 (N_5574,N_591,N_2098);
and U5575 (N_5575,N_1870,N_734);
or U5576 (N_5576,N_4192,N_3715);
or U5577 (N_5577,N_2517,N_600);
nor U5578 (N_5578,N_886,N_4888);
nor U5579 (N_5579,N_3877,N_4450);
and U5580 (N_5580,N_4288,N_2446);
nand U5581 (N_5581,N_2996,N_2074);
nor U5582 (N_5582,N_2761,N_4505);
or U5583 (N_5583,N_1779,N_456);
nand U5584 (N_5584,N_1044,N_1374);
and U5585 (N_5585,N_312,N_442);
nor U5586 (N_5586,N_1510,N_828);
and U5587 (N_5587,N_186,N_2005);
or U5588 (N_5588,N_4494,N_4541);
nor U5589 (N_5589,N_2400,N_680);
or U5590 (N_5590,N_4132,N_4227);
nor U5591 (N_5591,N_1383,N_4652);
nor U5592 (N_5592,N_3737,N_2250);
or U5593 (N_5593,N_3549,N_1886);
or U5594 (N_5594,N_1209,N_3518);
nor U5595 (N_5595,N_622,N_2302);
or U5596 (N_5596,N_3361,N_131);
and U5597 (N_5597,N_2057,N_2058);
and U5598 (N_5598,N_1029,N_2751);
nor U5599 (N_5599,N_1272,N_2922);
nand U5600 (N_5600,N_2192,N_1135);
nand U5601 (N_5601,N_2497,N_884);
or U5602 (N_5602,N_2645,N_616);
nor U5603 (N_5603,N_104,N_1370);
and U5604 (N_5604,N_1646,N_1773);
nor U5605 (N_5605,N_2879,N_807);
nand U5606 (N_5606,N_2915,N_2666);
or U5607 (N_5607,N_33,N_4908);
nand U5608 (N_5608,N_4230,N_1141);
nor U5609 (N_5609,N_3407,N_1850);
and U5610 (N_5610,N_1977,N_2416);
and U5611 (N_5611,N_845,N_3763);
nand U5612 (N_5612,N_1675,N_4738);
nor U5613 (N_5613,N_857,N_1904);
and U5614 (N_5614,N_3410,N_2850);
and U5615 (N_5615,N_1016,N_3728);
nand U5616 (N_5616,N_2481,N_2219);
nand U5617 (N_5617,N_3564,N_730);
or U5618 (N_5618,N_4428,N_980);
nor U5619 (N_5619,N_1584,N_4614);
and U5620 (N_5620,N_4975,N_1494);
and U5621 (N_5621,N_4180,N_3212);
nand U5622 (N_5622,N_3159,N_714);
or U5623 (N_5623,N_2925,N_1175);
and U5624 (N_5624,N_2317,N_3461);
and U5625 (N_5625,N_1012,N_518);
nor U5626 (N_5626,N_944,N_3302);
xor U5627 (N_5627,N_6,N_1210);
nand U5628 (N_5628,N_91,N_1947);
and U5629 (N_5629,N_2947,N_1608);
xor U5630 (N_5630,N_4487,N_406);
and U5631 (N_5631,N_1762,N_4767);
or U5632 (N_5632,N_2360,N_4679);
or U5633 (N_5633,N_620,N_4341);
and U5634 (N_5634,N_4683,N_1243);
or U5635 (N_5635,N_556,N_2041);
nor U5636 (N_5636,N_4858,N_4264);
or U5637 (N_5637,N_2152,N_2354);
or U5638 (N_5638,N_4079,N_153);
nor U5639 (N_5639,N_4775,N_2027);
nor U5640 (N_5640,N_2504,N_265);
nand U5641 (N_5641,N_20,N_2955);
or U5642 (N_5642,N_1635,N_2570);
or U5643 (N_5643,N_2321,N_4591);
nand U5644 (N_5644,N_1806,N_1955);
and U5645 (N_5645,N_797,N_438);
and U5646 (N_5646,N_4584,N_1637);
or U5647 (N_5647,N_4884,N_1523);
or U5648 (N_5648,N_3562,N_3022);
or U5649 (N_5649,N_822,N_1786);
or U5650 (N_5650,N_2931,N_2385);
nor U5651 (N_5651,N_1593,N_3327);
and U5652 (N_5652,N_1943,N_2580);
and U5653 (N_5653,N_625,N_931);
and U5654 (N_5654,N_3804,N_1495);
and U5655 (N_5655,N_4680,N_1938);
and U5656 (N_5656,N_4747,N_4084);
nor U5657 (N_5657,N_4875,N_2101);
and U5658 (N_5658,N_3238,N_1339);
or U5659 (N_5659,N_1195,N_2546);
nand U5660 (N_5660,N_191,N_3520);
or U5661 (N_5661,N_1214,N_3583);
or U5662 (N_5662,N_809,N_3516);
or U5663 (N_5663,N_1201,N_1211);
or U5664 (N_5664,N_1895,N_4458);
nand U5665 (N_5665,N_1893,N_889);
nor U5666 (N_5666,N_1451,N_782);
nor U5667 (N_5667,N_4248,N_283);
nor U5668 (N_5668,N_602,N_3091);
or U5669 (N_5669,N_2373,N_1316);
or U5670 (N_5670,N_2458,N_2387);
nand U5671 (N_5671,N_2609,N_111);
nor U5672 (N_5672,N_1815,N_2764);
nand U5673 (N_5673,N_1676,N_2393);
or U5674 (N_5674,N_3148,N_2798);
or U5675 (N_5675,N_2771,N_49);
or U5676 (N_5676,N_1098,N_417);
nor U5677 (N_5677,N_1203,N_2193);
nand U5678 (N_5678,N_3138,N_4086);
nand U5679 (N_5679,N_1108,N_255);
or U5680 (N_5680,N_3063,N_366);
nand U5681 (N_5681,N_3958,N_1271);
or U5682 (N_5682,N_1742,N_2992);
and U5683 (N_5683,N_4117,N_1402);
or U5684 (N_5684,N_451,N_315);
nand U5685 (N_5685,N_2260,N_4250);
nand U5686 (N_5686,N_1810,N_3869);
nor U5687 (N_5687,N_2989,N_1731);
or U5688 (N_5688,N_4306,N_2428);
nor U5689 (N_5689,N_1216,N_3112);
and U5690 (N_5690,N_1760,N_959);
nand U5691 (N_5691,N_4873,N_405);
and U5692 (N_5692,N_3275,N_3240);
or U5693 (N_5693,N_3136,N_723);
or U5694 (N_5694,N_3338,N_3745);
or U5695 (N_5695,N_4421,N_3265);
and U5696 (N_5696,N_4185,N_3772);
nand U5697 (N_5697,N_1925,N_979);
nor U5698 (N_5698,N_2129,N_2548);
nor U5699 (N_5699,N_4269,N_3303);
nor U5700 (N_5700,N_2376,N_1546);
nand U5701 (N_5701,N_27,N_2490);
or U5702 (N_5702,N_93,N_4818);
or U5703 (N_5703,N_3484,N_1658);
and U5704 (N_5704,N_1281,N_1380);
xor U5705 (N_5705,N_1393,N_1679);
or U5706 (N_5706,N_4433,N_1915);
or U5707 (N_5707,N_3120,N_1497);
and U5708 (N_5708,N_4190,N_2937);
and U5709 (N_5709,N_4515,N_3324);
or U5710 (N_5710,N_3280,N_2367);
nor U5711 (N_5711,N_2986,N_998);
nand U5712 (N_5712,N_3691,N_377);
and U5713 (N_5713,N_1574,N_2516);
nor U5714 (N_5714,N_913,N_4232);
nor U5715 (N_5715,N_1112,N_4986);
nand U5716 (N_5716,N_2111,N_4193);
nand U5717 (N_5717,N_4221,N_1902);
and U5718 (N_5718,N_1408,N_1390);
or U5719 (N_5719,N_3645,N_3088);
nand U5720 (N_5720,N_1397,N_2535);
or U5721 (N_5721,N_1999,N_4582);
or U5722 (N_5722,N_724,N_4370);
nor U5723 (N_5723,N_120,N_3433);
or U5724 (N_5724,N_226,N_3057);
and U5725 (N_5725,N_3290,N_1059);
nand U5726 (N_5726,N_2708,N_3690);
or U5727 (N_5727,N_570,N_271);
or U5728 (N_5728,N_3237,N_908);
and U5729 (N_5729,N_3277,N_4054);
nor U5730 (N_5730,N_2545,N_993);
nor U5731 (N_5731,N_3430,N_3913);
nand U5732 (N_5732,N_4632,N_1338);
nand U5733 (N_5733,N_1323,N_4064);
nand U5734 (N_5734,N_3602,N_4513);
nand U5735 (N_5735,N_4695,N_2757);
nor U5736 (N_5736,N_810,N_3802);
nor U5737 (N_5737,N_2576,N_544);
nor U5738 (N_5738,N_4492,N_2144);
or U5739 (N_5739,N_1528,N_1557);
nor U5740 (N_5740,N_1485,N_2657);
nand U5741 (N_5741,N_2493,N_1186);
nand U5742 (N_5742,N_1048,N_1472);
or U5743 (N_5743,N_812,N_3132);
or U5744 (N_5744,N_373,N_1824);
and U5745 (N_5745,N_470,N_4506);
nor U5746 (N_5746,N_2358,N_2307);
and U5747 (N_5747,N_2805,N_2622);
and U5748 (N_5748,N_4714,N_3987);
or U5749 (N_5749,N_3010,N_4241);
nor U5750 (N_5750,N_4635,N_4089);
and U5751 (N_5751,N_4454,N_4347);
nand U5752 (N_5752,N_2213,N_2183);
and U5753 (N_5753,N_2217,N_2444);
nor U5754 (N_5754,N_615,N_804);
nand U5755 (N_5755,N_3122,N_2993);
nand U5756 (N_5756,N_1301,N_575);
or U5757 (N_5757,N_3234,N_2088);
nor U5758 (N_5758,N_2566,N_3115);
nor U5759 (N_5759,N_1812,N_3216);
or U5760 (N_5760,N_4254,N_1733);
nand U5761 (N_5761,N_3943,N_2767);
or U5762 (N_5762,N_3503,N_3328);
or U5763 (N_5763,N_3419,N_4239);
or U5764 (N_5764,N_432,N_3746);
nor U5765 (N_5765,N_2429,N_2418);
nor U5766 (N_5766,N_4312,N_1598);
nor U5767 (N_5767,N_274,N_47);
or U5768 (N_5768,N_2308,N_4397);
nor U5769 (N_5769,N_2109,N_4980);
and U5770 (N_5770,N_703,N_2839);
nand U5771 (N_5771,N_1283,N_496);
or U5772 (N_5772,N_1923,N_4577);
nand U5773 (N_5773,N_247,N_1758);
and U5774 (N_5774,N_1137,N_4862);
xor U5775 (N_5775,N_1131,N_831);
nor U5776 (N_5776,N_4114,N_3596);
nor U5777 (N_5777,N_2353,N_4682);
nor U5778 (N_5778,N_3800,N_4382);
or U5779 (N_5779,N_3951,N_2895);
or U5780 (N_5780,N_234,N_1607);
and U5781 (N_5781,N_4285,N_3760);
nand U5782 (N_5782,N_368,N_3565);
or U5783 (N_5783,N_4711,N_3490);
nor U5784 (N_5784,N_2424,N_2016);
nor U5785 (N_5785,N_243,N_1874);
nand U5786 (N_5786,N_1367,N_479);
or U5787 (N_5787,N_4500,N_2817);
nand U5788 (N_5788,N_2962,N_2104);
nor U5789 (N_5789,N_4969,N_1089);
or U5790 (N_5790,N_495,N_3403);
nor U5791 (N_5791,N_1144,N_2291);
and U5792 (N_5792,N_3291,N_541);
or U5793 (N_5793,N_1531,N_4997);
nand U5794 (N_5794,N_4897,N_4430);
and U5795 (N_5795,N_1602,N_3467);
and U5796 (N_5796,N_3245,N_3257);
or U5797 (N_5797,N_4765,N_3685);
nor U5798 (N_5798,N_428,N_756);
nand U5799 (N_5799,N_3026,N_2503);
nand U5800 (N_5800,N_349,N_4460);
nor U5801 (N_5801,N_3703,N_3241);
nor U5802 (N_5802,N_1163,N_4143);
and U5803 (N_5803,N_2351,N_2032);
nand U5804 (N_5804,N_1205,N_4809);
or U5805 (N_5805,N_1916,N_4917);
nand U5806 (N_5806,N_3020,N_3070);
or U5807 (N_5807,N_630,N_77);
nand U5808 (N_5808,N_559,N_3730);
nor U5809 (N_5809,N_1819,N_987);
nand U5810 (N_5810,N_1976,N_2861);
and U5811 (N_5811,N_2998,N_2381);
nor U5812 (N_5812,N_2639,N_3021);
nand U5813 (N_5813,N_2362,N_2489);
nand U5814 (N_5814,N_4048,N_1881);
and U5815 (N_5815,N_1884,N_2203);
nor U5816 (N_5816,N_2956,N_464);
nand U5817 (N_5817,N_3331,N_624);
xor U5818 (N_5818,N_2390,N_4033);
and U5819 (N_5819,N_2007,N_4785);
nor U5820 (N_5820,N_892,N_2263);
nor U5821 (N_5821,N_1651,N_3889);
or U5822 (N_5822,N_306,N_2343);
and U5823 (N_5823,N_758,N_2175);
nand U5824 (N_5824,N_2640,N_2878);
nand U5825 (N_5825,N_3653,N_302);
and U5826 (N_5826,N_3404,N_4072);
and U5827 (N_5827,N_343,N_4213);
nor U5828 (N_5828,N_1133,N_4467);
nand U5829 (N_5829,N_1826,N_2133);
or U5830 (N_5830,N_3008,N_655);
or U5831 (N_5831,N_2802,N_1110);
or U5832 (N_5832,N_963,N_1671);
nand U5833 (N_5833,N_1011,N_3453);
nor U5834 (N_5834,N_1114,N_4194);
nor U5835 (N_5835,N_2938,N_539);
or U5836 (N_5836,N_3669,N_1470);
nor U5837 (N_5837,N_4532,N_1849);
and U5838 (N_5838,N_4904,N_3886);
and U5839 (N_5839,N_1713,N_2737);
and U5840 (N_5840,N_2397,N_2487);
or U5841 (N_5841,N_633,N_1164);
nor U5842 (N_5842,N_2719,N_1058);
or U5843 (N_5843,N_3106,N_560);
nor U5844 (N_5844,N_1517,N_500);
nand U5845 (N_5845,N_4282,N_1348);
nor U5846 (N_5846,N_38,N_4395);
nor U5847 (N_5847,N_3229,N_2049);
or U5848 (N_5848,N_3875,N_54);
or U5849 (N_5849,N_4580,N_1212);
nor U5850 (N_5850,N_3504,N_4791);
nand U5851 (N_5851,N_3164,N_1410);
nor U5852 (N_5852,N_340,N_3489);
nand U5853 (N_5853,N_4773,N_4970);
xnor U5854 (N_5854,N_4005,N_3048);
nor U5855 (N_5855,N_4474,N_2807);
and U5856 (N_5856,N_1855,N_3952);
or U5857 (N_5857,N_3454,N_4669);
nor U5858 (N_5858,N_3512,N_2151);
and U5859 (N_5859,N_4455,N_2963);
nand U5860 (N_5860,N_1610,N_2984);
and U5861 (N_5861,N_2436,N_566);
nand U5862 (N_5862,N_3287,N_2726);
or U5863 (N_5863,N_1279,N_3960);
or U5864 (N_5864,N_4787,N_3641);
nand U5865 (N_5865,N_2347,N_3642);
and U5866 (N_5866,N_1865,N_4153);
or U5867 (N_5867,N_472,N_79);
or U5868 (N_5868,N_1901,N_1379);
or U5869 (N_5869,N_4864,N_4545);
nand U5870 (N_5870,N_3714,N_3090);
nand U5871 (N_5871,N_4032,N_4156);
and U5872 (N_5872,N_1818,N_1781);
or U5873 (N_5873,N_239,N_4377);
nand U5874 (N_5874,N_682,N_4734);
nand U5875 (N_5875,N_645,N_2421);
nor U5876 (N_5876,N_1378,N_3015);
nor U5877 (N_5877,N_3332,N_982);
or U5878 (N_5878,N_766,N_174);
and U5879 (N_5879,N_22,N_4919);
or U5880 (N_5880,N_2009,N_1844);
nor U5881 (N_5881,N_1816,N_486);
nor U5882 (N_5882,N_1332,N_2465);
nand U5883 (N_5883,N_4759,N_3776);
or U5884 (N_5884,N_4320,N_1443);
or U5885 (N_5885,N_3340,N_1184);
nor U5886 (N_5886,N_2202,N_307);
or U5887 (N_5887,N_2698,N_4728);
nand U5888 (N_5888,N_2584,N_1479);
nor U5889 (N_5889,N_2120,N_2011);
and U5890 (N_5890,N_611,N_2209);
nand U5891 (N_5891,N_2157,N_1656);
or U5892 (N_5892,N_584,N_1853);
nor U5893 (N_5893,N_2135,N_1972);
nor U5894 (N_5894,N_4310,N_1457);
nand U5895 (N_5895,N_997,N_3103);
nand U5896 (N_5896,N_3692,N_1753);
nand U5897 (N_5897,N_4721,N_2596);
nor U5898 (N_5898,N_1740,N_3477);
or U5899 (N_5899,N_3764,N_2766);
or U5900 (N_5900,N_4823,N_899);
nor U5901 (N_5901,N_4121,N_1869);
and U5902 (N_5902,N_4464,N_3095);
nor U5903 (N_5903,N_3335,N_25);
nor U5904 (N_5904,N_201,N_2611);
and U5905 (N_5905,N_3415,N_3759);
and U5906 (N_5906,N_4556,N_1905);
or U5907 (N_5907,N_4348,N_3510);
or U5908 (N_5908,N_4456,N_2134);
or U5909 (N_5909,N_1369,N_3705);
and U5910 (N_5910,N_744,N_4746);
and U5911 (N_5911,N_2099,N_66);
or U5912 (N_5912,N_1389,N_4476);
and U5913 (N_5913,N_3589,N_1949);
or U5914 (N_5914,N_4044,N_1148);
and U5915 (N_5915,N_4381,N_164);
xnor U5916 (N_5916,N_4575,N_1028);
and U5917 (N_5917,N_1191,N_3325);
or U5918 (N_5918,N_2013,N_4902);
nor U5919 (N_5919,N_533,N_1027);
nor U5920 (N_5920,N_4479,N_3170);
nor U5921 (N_5921,N_3387,N_1845);
and U5922 (N_5922,N_1772,N_1307);
nand U5923 (N_5923,N_4563,N_1018);
nand U5924 (N_5924,N_4539,N_426);
nand U5925 (N_5925,N_3086,N_3480);
or U5926 (N_5926,N_3429,N_2344);
or U5927 (N_5927,N_3627,N_339);
nor U5928 (N_5928,N_4299,N_3606);
and U5929 (N_5929,N_2084,N_3292);
nor U5930 (N_5930,N_2038,N_388);
nand U5931 (N_5931,N_2107,N_1668);
and U5932 (N_5932,N_1705,N_2775);
and U5933 (N_5933,N_3754,N_2469);
or U5934 (N_5934,N_1544,N_1576);
nor U5935 (N_5935,N_1957,N_1330);
or U5936 (N_5936,N_3997,N_2206);
and U5937 (N_5937,N_1661,N_1554);
and U5938 (N_5938,N_3307,N_3524);
nor U5939 (N_5939,N_244,N_2616);
nand U5940 (N_5940,N_3888,N_2184);
nor U5941 (N_5941,N_4617,N_2533);
nor U5942 (N_5942,N_4090,N_98);
nand U5943 (N_5943,N_3349,N_2902);
nor U5944 (N_5944,N_2704,N_2113);
nor U5945 (N_5945,N_402,N_3228);
nand U5946 (N_5946,N_3432,N_1935);
nor U5947 (N_5947,N_1231,N_2085);
or U5948 (N_5948,N_3846,N_3268);
nand U5949 (N_5949,N_2349,N_3341);
and U5950 (N_5950,N_1655,N_577);
nand U5951 (N_5951,N_878,N_3628);
or U5952 (N_5952,N_4251,N_1324);
nand U5953 (N_5953,N_4304,N_1034);
and U5954 (N_5954,N_4045,N_2039);
nor U5955 (N_5955,N_2691,N_1304);
and U5956 (N_5956,N_1492,N_12);
and U5957 (N_5957,N_2092,N_4350);
nor U5958 (N_5958,N_375,N_4311);
nor U5959 (N_5959,N_4006,N_1973);
nor U5960 (N_5960,N_4082,N_1046);
and U5961 (N_5961,N_2391,N_780);
or U5962 (N_5962,N_4974,N_291);
or U5963 (N_5963,N_2772,N_3239);
nand U5964 (N_5964,N_4391,N_2648);
nand U5965 (N_5965,N_1419,N_868);
nor U5966 (N_5966,N_1769,N_4290);
nand U5967 (N_5967,N_4811,N_1096);
xor U5968 (N_5968,N_1435,N_1293);
or U5969 (N_5969,N_3600,N_923);
or U5970 (N_5970,N_2867,N_4340);
nand U5971 (N_5971,N_1490,N_517);
nor U5972 (N_5972,N_4106,N_939);
and U5973 (N_5973,N_2515,N_2900);
nand U5974 (N_5974,N_3648,N_4252);
and U5975 (N_5975,N_4998,N_666);
nor U5976 (N_5976,N_3348,N_3414);
nor U5977 (N_5977,N_3666,N_3482);
and U5978 (N_5978,N_4570,N_1357);
or U5979 (N_5979,N_3468,N_252);
and U5980 (N_5980,N_4369,N_293);
and U5981 (N_5981,N_741,N_4136);
nand U5982 (N_5982,N_1003,N_2438);
or U5983 (N_5983,N_641,N_977);
and U5984 (N_5984,N_501,N_1842);
or U5985 (N_5985,N_685,N_3525);
or U5986 (N_5986,N_3102,N_4160);
nor U5987 (N_5987,N_2562,N_148);
or U5988 (N_5988,N_2587,N_125);
nor U5989 (N_5989,N_1828,N_3621);
or U5990 (N_5990,N_4987,N_99);
xor U5991 (N_5991,N_896,N_1097);
or U5992 (N_5992,N_1392,N_4357);
and U5993 (N_5993,N_4912,N_2035);
and U5994 (N_5994,N_3758,N_4113);
nand U5995 (N_5995,N_4145,N_1437);
xnor U5996 (N_5996,N_3725,N_3982);
xor U5997 (N_5997,N_1825,N_2168);
nor U5998 (N_5998,N_2889,N_4991);
and U5999 (N_5999,N_401,N_618);
and U6000 (N_6000,N_4175,N_3182);
nand U6001 (N_6001,N_4994,N_2624);
or U6002 (N_6002,N_4782,N_3656);
or U6003 (N_6003,N_4689,N_1536);
or U6004 (N_6004,N_3296,N_2017);
or U6005 (N_6005,N_4712,N_3526);
and U6006 (N_6006,N_1783,N_3066);
and U6007 (N_6007,N_3969,N_1585);
and U6008 (N_6008,N_1169,N_326);
nor U6009 (N_6009,N_4806,N_672);
nor U6010 (N_6010,N_4976,N_4945);
nand U6011 (N_6011,N_2725,N_1549);
nand U6012 (N_6012,N_37,N_2886);
and U6013 (N_6013,N_1351,N_3156);
or U6014 (N_6014,N_4238,N_2329);
or U6015 (N_6015,N_2848,N_2885);
or U6016 (N_6016,N_3470,N_3805);
and U6017 (N_6017,N_4859,N_947);
nor U6018 (N_6018,N_2899,N_3841);
nand U6019 (N_6019,N_1159,N_2911);
or U6020 (N_6020,N_4087,N_3808);
nor U6021 (N_6021,N_3266,N_2077);
nor U6022 (N_6022,N_2722,N_595);
and U6023 (N_6023,N_2146,N_3288);
nor U6024 (N_6024,N_1868,N_549);
or U6025 (N_6025,N_3165,N_454);
and U6026 (N_6026,N_3065,N_4882);
xnor U6027 (N_6027,N_2082,N_1080);
and U6028 (N_6028,N_2226,N_2363);
or U6029 (N_6029,N_3994,N_4305);
nand U6030 (N_6030,N_3297,N_2924);
or U6031 (N_6031,N_3837,N_3595);
and U6032 (N_6032,N_505,N_4601);
and U6033 (N_6033,N_2554,N_1919);
and U6034 (N_6034,N_1162,N_2286);
nor U6035 (N_6035,N_3001,N_531);
or U6036 (N_6036,N_743,N_1063);
or U6037 (N_6037,N_4707,N_3915);
or U6038 (N_6038,N_1056,N_2638);
nor U6039 (N_6039,N_2676,N_4434);
nand U6040 (N_6040,N_3590,N_19);
nand U6041 (N_6041,N_1418,N_4598);
or U6042 (N_6042,N_704,N_1455);
and U6043 (N_6043,N_1724,N_3826);
nor U6044 (N_6044,N_948,N_3897);
or U6045 (N_6045,N_4829,N_2488);
nand U6046 (N_6046,N_4894,N_781);
and U6047 (N_6047,N_1766,N_4231);
nor U6048 (N_6048,N_2064,N_346);
and U6049 (N_6049,N_3098,N_1054);
nand U6050 (N_6050,N_4824,N_711);
nor U6051 (N_6051,N_3067,N_1006);
or U6052 (N_6052,N_2276,N_3261);
or U6053 (N_6053,N_350,N_439);
or U6054 (N_6054,N_228,N_1890);
or U6055 (N_6055,N_2742,N_494);
nand U6056 (N_6056,N_3320,N_2834);
and U6057 (N_6057,N_4195,N_681);
or U6058 (N_6058,N_2355,N_70);
or U6059 (N_6059,N_4148,N_4995);
nor U6060 (N_6060,N_3687,N_4287);
or U6061 (N_6061,N_365,N_4780);
and U6062 (N_6062,N_3955,N_550);
or U6063 (N_6063,N_543,N_392);
nor U6064 (N_6064,N_1481,N_3622);
nor U6065 (N_6065,N_3967,N_4437);
nand U6066 (N_6066,N_793,N_3773);
or U6067 (N_6067,N_2759,N_4704);
or U6068 (N_6068,N_2396,N_150);
nor U6069 (N_6069,N_2522,N_2637);
nand U6070 (N_6070,N_4438,N_2783);
and U6071 (N_6071,N_4534,N_1465);
nor U6072 (N_6072,N_1036,N_2803);
nor U6073 (N_6073,N_2511,N_2714);
or U6074 (N_6074,N_1583,N_3517);
and U6075 (N_6075,N_1260,N_869);
or U6076 (N_6076,N_754,N_3883);
and U6077 (N_6077,N_3494,N_4543);
and U6078 (N_6078,N_245,N_1987);
xnor U6079 (N_6079,N_1686,N_4883);
nor U6080 (N_6080,N_4978,N_3866);
nand U6081 (N_6081,N_2243,N_3096);
and U6082 (N_6082,N_1264,N_4131);
nand U6083 (N_6083,N_2912,N_2820);
nor U6084 (N_6084,N_2460,N_4204);
nand U6085 (N_6085,N_900,N_2409);
or U6086 (N_6086,N_996,N_771);
and U6087 (N_6087,N_1199,N_3286);
and U6088 (N_6088,N_894,N_404);
nand U6089 (N_6089,N_3858,N_4366);
or U6090 (N_6090,N_455,N_2808);
nor U6091 (N_6091,N_2568,N_2271);
and U6092 (N_6092,N_2731,N_893);
or U6093 (N_6093,N_2153,N_4972);
nand U6094 (N_6094,N_4781,N_639);
or U6095 (N_6095,N_4126,N_2934);
and U6096 (N_6096,N_3105,N_1078);
and U6097 (N_6097,N_3037,N_449);
and U6098 (N_6098,N_895,N_2128);
or U6099 (N_6099,N_2578,N_2655);
or U6100 (N_6100,N_1519,N_3304);
and U6101 (N_6101,N_1565,N_1882);
nand U6102 (N_6102,N_3538,N_938);
nand U6103 (N_6103,N_509,N_1538);
nand U6104 (N_6104,N_4609,N_867);
and U6105 (N_6105,N_3405,N_4293);
nand U6106 (N_6106,N_122,N_2628);
and U6107 (N_6107,N_3922,N_1597);
and U6108 (N_6108,N_3299,N_905);
or U6109 (N_6109,N_817,N_1286);
and U6110 (N_6110,N_1095,N_1946);
or U6111 (N_6111,N_659,N_2200);
nor U6112 (N_6112,N_101,N_3448);
and U6113 (N_6113,N_2828,N_183);
and U6114 (N_6114,N_475,N_299);
nand U6115 (N_6115,N_4581,N_2440);
and U6116 (N_6116,N_3946,N_393);
and U6117 (N_6117,N_529,N_3605);
nand U6118 (N_6118,N_3502,N_1466);
nand U6119 (N_6119,N_2268,N_2037);
and U6120 (N_6120,N_4124,N_1986);
nand U6121 (N_6121,N_1838,N_2547);
nand U6122 (N_6122,N_4095,N_2448);
and U6123 (N_6123,N_2797,N_2670);
and U6124 (N_6124,N_4938,N_1632);
nand U6125 (N_6125,N_3726,N_1464);
and U6126 (N_6126,N_3445,N_3522);
or U6127 (N_6127,N_2466,N_4199);
nand U6128 (N_6128,N_4012,N_1373);
nand U6129 (N_6129,N_1791,N_3928);
nand U6130 (N_6130,N_4258,N_87);
nor U6131 (N_6131,N_463,N_4338);
nand U6132 (N_6132,N_2520,N_1318);
nand U6133 (N_6133,N_4959,N_4219);
xor U6134 (N_6134,N_3314,N_2697);
nor U6135 (N_6135,N_4333,N_3932);
nand U6136 (N_6136,N_4085,N_3929);
or U6137 (N_6137,N_2412,N_2656);
or U6138 (N_6138,N_4240,N_4552);
or U6139 (N_6139,N_2053,N_673);
and U6140 (N_6140,N_1306,N_4317);
xnor U6141 (N_6141,N_4774,N_1956);
nand U6142 (N_6142,N_1040,N_1017);
nand U6143 (N_6143,N_1230,N_3953);
nand U6144 (N_6144,N_2215,N_4186);
or U6145 (N_6145,N_1229,N_1150);
nor U6146 (N_6146,N_1427,N_1193);
and U6147 (N_6147,N_928,N_904);
nand U6148 (N_6148,N_3472,N_3747);
or U6149 (N_6149,N_9,N_3232);
and U6150 (N_6150,N_4763,N_1429);
nand U6151 (N_6151,N_4352,N_2070);
or U6152 (N_6152,N_4659,N_4118);
and U6153 (N_6153,N_1889,N_3055);
or U6154 (N_6154,N_1105,N_1702);
nand U6155 (N_6155,N_4918,N_4419);
nor U6156 (N_6156,N_2571,N_4608);
and U6157 (N_6157,N_1372,N_2015);
xnor U6158 (N_6158,N_4891,N_2241);
nand U6159 (N_6159,N_1247,N_4665);
nor U6160 (N_6160,N_537,N_1763);
and U6161 (N_6161,N_3388,N_3632);
or U6162 (N_6162,N_1856,N_2290);
nor U6163 (N_6163,N_1077,N_2572);
nand U6164 (N_6164,N_3707,N_147);
nand U6165 (N_6165,N_3281,N_4807);
nand U6166 (N_6166,N_598,N_2668);
or U6167 (N_6167,N_2598,N_2589);
nor U6168 (N_6168,N_4876,N_1732);
or U6169 (N_6169,N_4745,N_975);
or U6170 (N_6170,N_82,N_3360);
nor U6171 (N_6171,N_1537,N_4826);
or U6172 (N_6172,N_2896,N_2004);
nand U6173 (N_6173,N_1072,N_4263);
nand U6174 (N_6174,N_2869,N_4957);
and U6175 (N_6175,N_4383,N_1641);
and U6176 (N_6176,N_3230,N_3801);
nor U6177 (N_6177,N_2880,N_4621);
nor U6178 (N_6178,N_3018,N_1100);
or U6179 (N_6179,N_4741,N_820);
nor U6180 (N_6180,N_3117,N_648);
or U6181 (N_6181,N_2739,N_4246);
nand U6182 (N_6182,N_589,N_2090);
or U6183 (N_6183,N_4324,N_3113);
nor U6184 (N_6184,N_4800,N_4846);
nor U6185 (N_6185,N_4226,N_1327);
or U6186 (N_6186,N_2928,N_423);
nand U6187 (N_6187,N_705,N_4967);
or U6188 (N_6188,N_3860,N_2115);
or U6189 (N_6189,N_608,N_1093);
or U6190 (N_6190,N_2826,N_310);
nor U6191 (N_6191,N_1692,N_832);
nor U6192 (N_6192,N_3217,N_3983);
nor U6193 (N_6193,N_4817,N_386);
or U6194 (N_6194,N_2608,N_2748);
xor U6195 (N_6195,N_1496,N_3092);
nand U6196 (N_6196,N_4378,N_4845);
and U6197 (N_6197,N_3631,N_130);
nand U6198 (N_6198,N_1213,N_3907);
nand U6199 (N_6199,N_2615,N_751);
nor U6200 (N_6200,N_3810,N_4181);
nor U6201 (N_6201,N_1964,N_3879);
nand U6202 (N_6202,N_4367,N_3311);
nor U6203 (N_6203,N_3900,N_1041);
and U6204 (N_6204,N_1913,N_4548);
or U6205 (N_6205,N_1852,N_1460);
or U6206 (N_6206,N_297,N_3079);
or U6207 (N_6207,N_493,N_2851);
or U6208 (N_6208,N_4594,N_4840);
nor U6209 (N_6209,N_2066,N_720);
or U6210 (N_6210,N_4061,N_2019);
and U6211 (N_6211,N_4860,N_2796);
nor U6212 (N_6212,N_1628,N_1319);
and U6213 (N_6213,N_2884,N_3547);
nand U6214 (N_6214,N_4606,N_4940);
and U6215 (N_6215,N_1426,N_576);
and U6216 (N_6216,N_4100,N_1);
nor U6217 (N_6217,N_3456,N_3464);
nor U6218 (N_6218,N_1068,N_3514);
nand U6219 (N_6219,N_2023,N_1569);
or U6220 (N_6220,N_891,N_311);
nor U6221 (N_6221,N_2913,N_3521);
or U6222 (N_6222,N_1990,N_732);
nand U6223 (N_6223,N_3859,N_4948);
nor U6224 (N_6224,N_3171,N_3774);
and U6225 (N_6225,N_4169,N_532);
and U6226 (N_6226,N_4729,N_2747);
or U6227 (N_6227,N_3769,N_3431);
xor U6228 (N_6228,N_4943,N_1616);
nor U6229 (N_6229,N_777,N_2605);
and U6230 (N_6230,N_3675,N_4362);
nand U6231 (N_6231,N_199,N_2506);
nor U6232 (N_6232,N_3200,N_2040);
and U6233 (N_6233,N_4607,N_2612);
xnor U6234 (N_6234,N_2304,N_3840);
and U6235 (N_6235,N_2472,N_2935);
nor U6236 (N_6236,N_4098,N_2375);
nand U6237 (N_6237,N_2374,N_2685);
nand U6238 (N_6238,N_2699,N_1328);
or U6239 (N_6239,N_4017,N_65);
nor U6240 (N_6240,N_4425,N_1640);
nor U6241 (N_6241,N_1515,N_473);
or U6242 (N_6242,N_2464,N_4468);
nor U6243 (N_6243,N_418,N_3380);
xnor U6244 (N_6244,N_498,N_1176);
or U6245 (N_6245,N_3878,N_3854);
or U6246 (N_6246,N_2882,N_35);
or U6247 (N_6247,N_4770,N_2148);
nor U6248 (N_6248,N_2403,N_4838);
nor U6249 (N_6249,N_995,N_3823);
or U6250 (N_6250,N_4906,N_4224);
and U6251 (N_6251,N_2590,N_3100);
and U6252 (N_6252,N_1434,N_737);
or U6253 (N_6253,N_951,N_5);
and U6254 (N_6254,N_3383,N_2536);
nand U6255 (N_6255,N_1722,N_2345);
nand U6256 (N_6256,N_179,N_3604);
and U6257 (N_6257,N_3578,N_2814);
and U6258 (N_6258,N_3034,N_1603);
or U6259 (N_6259,N_3127,N_4406);
and U6260 (N_6260,N_818,N_3452);
and U6261 (N_6261,N_853,N_2994);
or U6262 (N_6262,N_1929,N_4613);
or U6263 (N_6263,N_430,N_1071);
or U6264 (N_6264,N_763,N_2833);
nand U6265 (N_6265,N_2299,N_735);
and U6266 (N_6266,N_1296,N_3274);
nor U6267 (N_6267,N_2588,N_4490);
nor U6268 (N_6268,N_912,N_3693);
nor U6269 (N_6269,N_1797,N_1153);
or U6270 (N_6270,N_4363,N_1444);
and U6271 (N_6271,N_3649,N_2799);
and U6272 (N_6272,N_3847,N_3087);
nor U6273 (N_6273,N_1803,N_4920);
xor U6274 (N_6274,N_3073,N_3789);
or U6275 (N_6275,N_1364,N_3660);
and U6276 (N_6276,N_2176,N_4815);
nor U6277 (N_6277,N_3359,N_1605);
nor U6278 (N_6278,N_3319,N_3363);
nor U6279 (N_6279,N_4412,N_4452);
or U6280 (N_6280,N_767,N_4961);
or U6281 (N_6281,N_2758,N_1299);
nor U6282 (N_6282,N_2459,N_2423);
nand U6283 (N_6283,N_334,N_4423);
or U6284 (N_6284,N_4769,N_159);
nand U6285 (N_6285,N_3119,N_2447);
or U6286 (N_6286,N_3540,N_4936);
and U6287 (N_6287,N_1288,N_3743);
and U6288 (N_6288,N_594,N_3963);
or U6289 (N_6289,N_3771,N_1683);
and U6290 (N_6290,N_3861,N_4992);
or U6291 (N_6291,N_2684,N_4593);
xor U6292 (N_6292,N_3,N_137);
and U6293 (N_6293,N_2553,N_2907);
or U6294 (N_6294,N_2710,N_3371);
and U6295 (N_6295,N_4636,N_719);
nand U6296 (N_6296,N_968,N_1623);
and U6297 (N_6297,N_4053,N_3825);
and U6298 (N_6298,N_4390,N_840);
or U6299 (N_6299,N_2024,N_4386);
and U6300 (N_6300,N_769,N_2359);
and U6301 (N_6301,N_2824,N_2854);
nor U6302 (N_6302,N_4332,N_4737);
nand U6303 (N_6303,N_749,N_4388);
nand U6304 (N_6304,N_3462,N_4046);
nand U6305 (N_6305,N_2942,N_3379);
xor U6306 (N_6306,N_679,N_3678);
nor U6307 (N_6307,N_3551,N_3047);
and U6308 (N_6308,N_2838,N_2298);
and U6309 (N_6309,N_4166,N_1975);
nand U6310 (N_6310,N_3976,N_829);
or U6311 (N_6311,N_4561,N_2392);
and U6312 (N_6312,N_2720,N_2222);
nor U6313 (N_6313,N_4439,N_1143);
nor U6314 (N_6314,N_440,N_1065);
nor U6315 (N_6315,N_4502,N_4717);
or U6316 (N_6316,N_2738,N_3663);
and U6317 (N_6317,N_3143,N_690);
nand U6318 (N_6318,N_1792,N_296);
or U6319 (N_6319,N_1622,N_675);
nand U6320 (N_6320,N_1774,N_4639);
nor U6321 (N_6321,N_644,N_4266);
nand U6322 (N_6322,N_4376,N_3375);
nor U6323 (N_6323,N_4628,N_3688);
nor U6324 (N_6324,N_3981,N_746);
nor U6325 (N_6325,N_628,N_2653);
nand U6326 (N_6326,N_872,N_2959);
nand U6327 (N_6327,N_3708,N_4327);
nand U6328 (N_6328,N_1789,N_1793);
and U6329 (N_6329,N_3013,N_1961);
nor U6330 (N_6330,N_4776,N_3062);
nand U6331 (N_6331,N_568,N_1228);
and U6332 (N_6332,N_796,N_3293);
and U6333 (N_6333,N_4138,N_4501);
nand U6334 (N_6334,N_4127,N_2237);
and U6335 (N_6335,N_2593,N_1712);
nand U6336 (N_6336,N_2727,N_2837);
nand U6337 (N_6337,N_2930,N_3876);
nand U6338 (N_6338,N_2196,N_3262);
or U6339 (N_6339,N_3169,N_64);
nor U6340 (N_6340,N_1748,N_651);
nor U6341 (N_6341,N_268,N_2981);
nand U6342 (N_6342,N_1329,N_3479);
nor U6343 (N_6343,N_3219,N_728);
nand U6344 (N_6344,N_2214,N_2042);
and U6345 (N_6345,N_4392,N_1617);
nor U6346 (N_6346,N_1127,N_4574);
nor U6347 (N_6347,N_3850,N_2366);
and U6348 (N_6348,N_2340,N_3394);
xnor U6349 (N_6349,N_2199,N_4303);
nor U6350 (N_6350,N_3734,N_223);
nor U6351 (N_6351,N_24,N_729);
and U6352 (N_6352,N_1064,N_3139);
nor U6353 (N_6353,N_2658,N_3626);
nand U6354 (N_6354,N_2988,N_4380);
nor U6355 (N_6355,N_144,N_945);
nand U6356 (N_6356,N_4364,N_3783);
and U6357 (N_6357,N_2632,N_17);
nor U6358 (N_6358,N_2577,N_2816);
nand U6359 (N_6359,N_3108,N_808);
nor U6360 (N_6360,N_4560,N_3439);
or U6361 (N_6361,N_3914,N_3289);
nor U6362 (N_6362,N_3934,N_4522);
or U6363 (N_6363,N_436,N_936);
and U6364 (N_6364,N_3177,N_4080);
and U6365 (N_6365,N_1581,N_2524);
nand U6366 (N_6366,N_1168,N_329);
and U6367 (N_6367,N_2948,N_3060);
or U6368 (N_6368,N_3816,N_390);
and U6369 (N_6369,N_4854,N_2502);
nand U6370 (N_6370,N_3033,N_1037);
or U6371 (N_6371,N_1439,N_2297);
nand U6372 (N_6372,N_2356,N_839);
nand U6373 (N_6373,N_1652,N_4725);
nand U6374 (N_6374,N_1256,N_3699);
and U6375 (N_6375,N_4612,N_2264);
nand U6376 (N_6376,N_3214,N_2567);
and U6377 (N_6377,N_241,N_4623);
or U6378 (N_6378,N_757,N_3709);
and U6379 (N_6379,N_4010,N_3141);
nand U6380 (N_6380,N_477,N_4694);
nor U6381 (N_6381,N_193,N_4794);
or U6382 (N_6382,N_1998,N_4557);
or U6383 (N_6383,N_925,N_1930);
nor U6384 (N_6384,N_2036,N_1477);
nand U6385 (N_6385,N_3263,N_816);
or U6386 (N_6386,N_2908,N_3382);
or U6387 (N_6387,N_1759,N_1094);
and U6388 (N_6388,N_4630,N_860);
or U6389 (N_6389,N_3949,N_3362);
nor U6390 (N_6390,N_3392,N_2746);
or U6391 (N_6391,N_4566,N_4643);
nor U6392 (N_6392,N_4212,N_488);
nand U6393 (N_6393,N_1564,N_1469);
and U6394 (N_6394,N_1062,N_1488);
nor U6395 (N_6395,N_2198,N_1088);
or U6396 (N_6396,N_2477,N_1863);
nand U6397 (N_6397,N_3032,N_1349);
nand U6398 (N_6398,N_3260,N_1081);
and U6399 (N_6399,N_593,N_4035);
nor U6400 (N_6400,N_205,N_280);
nor U6401 (N_6401,N_2277,N_3856);
and U6402 (N_6402,N_4724,N_2573);
nor U6403 (N_6403,N_4678,N_4399);
or U6404 (N_6404,N_1685,N_80);
nor U6405 (N_6405,N_3166,N_1223);
nor U6406 (N_6406,N_3134,N_976);
or U6407 (N_6407,N_4004,N_3731);
and U6408 (N_6408,N_3784,N_4099);
and U6409 (N_6409,N_4315,N_2339);
nand U6410 (N_6410,N_2873,N_4424);
and U6411 (N_6411,N_2224,N_2810);
nor U6412 (N_6412,N_414,N_2473);
nor U6413 (N_6413,N_919,N_3326);
and U6414 (N_6414,N_4147,N_1689);
nand U6415 (N_6415,N_448,N_4034);
nand U6416 (N_6416,N_453,N_4516);
nor U6417 (N_6417,N_480,N_2045);
nand U6418 (N_6418,N_462,N_3014);
and U6419 (N_6419,N_2705,N_3485);
and U6420 (N_6420,N_935,N_1875);
and U6421 (N_6421,N_1877,N_3487);
nor U6422 (N_6422,N_4855,N_200);
and U6423 (N_6423,N_2871,N_1236);
or U6424 (N_6424,N_4808,N_2599);
nand U6425 (N_6425,N_2883,N_1561);
nor U6426 (N_6426,N_3330,N_1997);
nand U6427 (N_6427,N_3892,N_364);
nand U6428 (N_6428,N_3803,N_3721);
and U6429 (N_6429,N_118,N_4907);
nor U6430 (N_6430,N_3025,N_647);
or U6431 (N_6431,N_1860,N_2159);
and U6432 (N_6432,N_4092,N_1503);
nor U6433 (N_6433,N_4483,N_1507);
nor U6434 (N_6434,N_1699,N_1407);
or U6435 (N_6435,N_63,N_476);
nand U6436 (N_6436,N_3752,N_811);
nand U6437 (N_6437,N_3761,N_657);
nor U6438 (N_6438,N_926,N_4603);
or U6439 (N_6439,N_355,N_1846);
nand U6440 (N_6440,N_1883,N_3056);
and U6441 (N_6441,N_2309,N_1587);
nand U6442 (N_6442,N_3996,N_3739);
and U6443 (N_6443,N_4123,N_953);
nand U6444 (N_6444,N_2187,N_2654);
nor U6445 (N_6445,N_3809,N_4599);
nor U6446 (N_6446,N_1366,N_1992);
nor U6447 (N_6447,N_888,N_2774);
nand U6448 (N_6448,N_661,N_4743);
or U6449 (N_6449,N_1026,N_2368);
nand U6450 (N_6450,N_3785,N_3529);
nor U6451 (N_6451,N_3591,N_4751);
nand U6452 (N_6452,N_4191,N_133);
nor U6453 (N_6453,N_3372,N_4928);
nor U6454 (N_6454,N_1611,N_2647);
nor U6455 (N_6455,N_3563,N_2849);
and U6456 (N_6456,N_3665,N_2402);
or U6457 (N_6457,N_4038,N_258);
nor U6458 (N_6458,N_3039,N_1645);
nand U6459 (N_6459,N_3395,N_4596);
or U6460 (N_6460,N_3220,N_1196);
and U6461 (N_6461,N_3599,N_2238);
nor U6462 (N_6462,N_1518,N_2507);
and U6463 (N_6463,N_1070,N_738);
nor U6464 (N_6464,N_3133,N_3919);
nand U6465 (N_6465,N_3607,N_4158);
nor U6466 (N_6466,N_4827,N_2435);
and U6467 (N_6467,N_2643,N_380);
or U6468 (N_6468,N_2468,N_39);
nand U6469 (N_6469,N_400,N_4146);
nand U6470 (N_6470,N_4661,N_3639);
nor U6471 (N_6471,N_4921,N_3985);
or U6472 (N_6472,N_2540,N_3757);
and U6473 (N_6473,N_335,N_649);
nand U6474 (N_6474,N_2383,N_140);
or U6475 (N_6475,N_1525,N_238);
or U6476 (N_6476,N_4426,N_224);
nor U6477 (N_6477,N_1979,N_204);
and U6478 (N_6478,N_4551,N_45);
and U6479 (N_6479,N_2173,N_3174);
nor U6480 (N_6480,N_1284,N_941);
nor U6481 (N_6481,N_4493,N_4732);
or U6482 (N_6482,N_4837,N_3183);
or U6483 (N_6483,N_3704,N_3972);
nand U6484 (N_6484,N_1432,N_1436);
nor U6485 (N_6485,N_1706,N_3189);
nor U6486 (N_6486,N_2521,N_3988);
and U6487 (N_6487,N_875,N_2117);
or U6488 (N_6488,N_1294,N_4536);
nor U6489 (N_6489,N_972,N_852);
or U6490 (N_6490,N_2328,N_3713);
nor U6491 (N_6491,N_2665,N_3792);
nand U6492 (N_6492,N_4926,N_4336);
or U6493 (N_6493,N_4924,N_1403);
and U6494 (N_6494,N_445,N_3548);
and U6495 (N_6495,N_4658,N_166);
and U6496 (N_6496,N_883,N_2127);
nor U6497 (N_6497,N_3187,N_2072);
or U6498 (N_6498,N_2754,N_580);
nand U6499 (N_6499,N_3000,N_1295);
nor U6500 (N_6500,N_1312,N_903);
nand U6501 (N_6501,N_3258,N_2105);
or U6502 (N_6502,N_4203,N_394);
or U6503 (N_6503,N_3937,N_3839);
nand U6504 (N_6504,N_374,N_1892);
and U6505 (N_6505,N_3040,N_2875);
nor U6506 (N_6506,N_123,N_4510);
or U6507 (N_6507,N_2619,N_3993);
nor U6508 (N_6508,N_565,N_2171);
nor U6509 (N_6509,N_1533,N_156);
nand U6510 (N_6510,N_1489,N_2001);
or U6511 (N_6511,N_4620,N_3029);
and U6512 (N_6512,N_1287,N_235);
or U6513 (N_6513,N_2991,N_197);
nand U6514 (N_6514,N_2161,N_2474);
nor U6515 (N_6515,N_1182,N_3028);
nand U6516 (N_6516,N_304,N_1362);
or U6517 (N_6517,N_2335,N_882);
nor U6518 (N_6518,N_4528,N_990);
nand U6519 (N_6519,N_2811,N_469);
and U6520 (N_6520,N_985,N_2234);
nand U6521 (N_6521,N_1341,N_792);
nor U6522 (N_6522,N_795,N_4471);
and U6523 (N_6523,N_1527,N_3005);
nor U6524 (N_6524,N_3455,N_4511);
and U6525 (N_6525,N_4188,N_1333);
and U6526 (N_6526,N_650,N_3554);
nand U6527 (N_6527,N_2463,N_2876);
or U6528 (N_6528,N_3698,N_3990);
nand U6529 (N_6529,N_2966,N_1009);
nand U6530 (N_6530,N_4075,N_4857);
or U6531 (N_6531,N_3059,N_2208);
and U6532 (N_6532,N_4509,N_3791);
xnor U6533 (N_6533,N_2888,N_3474);
or U6534 (N_6534,N_73,N_3513);
nor U6535 (N_6535,N_4431,N_3447);
nand U6536 (N_6536,N_3417,N_4116);
nor U6537 (N_6537,N_2300,N_3422);
and U6538 (N_6538,N_4177,N_4469);
nand U6539 (N_6539,N_1604,N_4284);
nor U6540 (N_6540,N_3706,N_4498);
and U6541 (N_6541,N_4531,N_4062);
or U6542 (N_6542,N_1106,N_4517);
or U6543 (N_6543,N_2542,N_119);
or U6544 (N_6544,N_506,N_3833);
and U6545 (N_6545,N_3427,N_2204);
nand U6546 (N_6546,N_4189,N_105);
nand U6547 (N_6547,N_3696,N_3838);
or U6548 (N_6548,N_629,N_1618);
nor U6549 (N_6549,N_3995,N_44);
and U6550 (N_6550,N_2801,N_2372);
or U6551 (N_6551,N_2845,N_2625);
and U6552 (N_6552,N_383,N_1823);
nor U6553 (N_6553,N_1907,N_1508);
nand U6554 (N_6554,N_92,N_3975);
and U6555 (N_6555,N_4504,N_2244);
nand U6556 (N_6556,N_1007,N_1529);
nand U6557 (N_6557,N_3179,N_1334);
nor U6558 (N_6558,N_2745,N_3664);
or U6559 (N_6559,N_954,N_4300);
nand U6560 (N_6560,N_4942,N_1200);
and U6561 (N_6561,N_1730,N_2717);
and U6562 (N_6562,N_2425,N_4247);
or U6563 (N_6563,N_1326,N_2426);
or U6564 (N_6564,N_411,N_4881);
nand U6565 (N_6565,N_750,N_3834);
and U6566 (N_6566,N_3898,N_185);
nor U6567 (N_6567,N_4757,N_357);
or U6568 (N_6568,N_4052,N_3765);
and U6569 (N_6569,N_819,N_2827);
or U6570 (N_6570,N_3460,N_4049);
nand U6571 (N_6571,N_2905,N_261);
nor U6572 (N_6572,N_1343,N_4833);
nand U6573 (N_6573,N_3301,N_2331);
nand U6574 (N_6574,N_1751,N_528);
and U6575 (N_6575,N_2334,N_4654);
or U6576 (N_6576,N_1667,N_3333);
xnor U6577 (N_6577,N_3411,N_4567);
and U6578 (N_6578,N_4368,N_3697);
and U6579 (N_6579,N_4899,N_545);
nand U6580 (N_6580,N_2316,N_2629);
nand U6581 (N_6581,N_2679,N_3568);
or U6582 (N_6582,N_2952,N_2388);
nor U6583 (N_6583,N_3964,N_1590);
and U6584 (N_6584,N_4346,N_489);
nor U6585 (N_6585,N_4733,N_1897);
or U6586 (N_6586,N_465,N_433);
nand U6587 (N_6587,N_3668,N_2528);
nand U6588 (N_6588,N_3085,N_1693);
nor U6589 (N_6589,N_1142,N_2974);
nor U6590 (N_6590,N_67,N_3597);
and U6591 (N_6591,N_3147,N_4616);
or U6592 (N_6592,N_194,N_2289);
xnor U6593 (N_6593,N_4245,N_4710);
or U6594 (N_6594,N_1567,N_2786);
xnor U6595 (N_6595,N_4909,N_3201);
or U6596 (N_6596,N_823,N_3936);
nor U6597 (N_6597,N_1483,N_1776);
nor U6598 (N_6598,N_513,N_2165);
nor U6599 (N_6599,N_3777,N_4105);
or U6600 (N_6600,N_874,N_4671);
nor U6601 (N_6601,N_1104,N_1917);
and U6602 (N_6602,N_4520,N_4296);
and U6603 (N_6603,N_2470,N_379);
or U6604 (N_6604,N_4257,N_2141);
nor U6605 (N_6605,N_1573,N_1514);
nand U6606 (N_6606,N_582,N_332);
and U6607 (N_6607,N_2229,N_4895);
and U6608 (N_6608,N_4176,N_2945);
nor U6609 (N_6609,N_1344,N_2380);
and U6610 (N_6610,N_3974,N_3457);
or U6611 (N_6611,N_991,N_1910);
nor U6612 (N_6612,N_578,N_4326);
or U6613 (N_6613,N_2855,N_551);
nor U6614 (N_6614,N_753,N_4754);
or U6615 (N_6615,N_2056,N_2760);
nand U6616 (N_6616,N_4638,N_1222);
or U6617 (N_6617,N_2788,N_4018);
nand U6618 (N_6618,N_706,N_2995);
or U6619 (N_6619,N_4578,N_485);
and U6620 (N_6620,N_1262,N_4863);
nor U6621 (N_6621,N_4201,N_4174);
nand U6622 (N_6622,N_3836,N_640);
nor U6623 (N_6623,N_1083,N_3601);
nor U6624 (N_6624,N_292,N_3770);
and U6625 (N_6625,N_922,N_4197);
nor U6626 (N_6626,N_4525,N_3654);
nand U6627 (N_6627,N_3930,N_2185);
nor U6628 (N_6628,N_3558,N_2787);
or U6629 (N_6629,N_165,N_16);
and U6630 (N_6630,N_3807,N_2230);
and U6631 (N_6631,N_4372,N_2212);
and U6632 (N_6632,N_3979,N_3038);
and U6633 (N_6633,N_1801,N_3917);
or U6634 (N_6634,N_783,N_2028);
and U6635 (N_6635,N_2220,N_527);
nand U6636 (N_6636,N_4861,N_1045);
nand U6637 (N_6637,N_220,N_631);
or U6638 (N_6638,N_2089,N_3865);
or U6639 (N_6639,N_2149,N_967);
and U6640 (N_6640,N_2006,N_409);
nor U6641 (N_6641,N_2483,N_3295);
nand U6642 (N_6642,N_4648,N_1983);
and U6643 (N_6643,N_909,N_1066);
or U6644 (N_6644,N_642,N_3225);
nor U6645 (N_6645,N_4761,N_4448);
nor U6646 (N_6646,N_667,N_2216);
or U6647 (N_6647,N_3694,N_3218);
nand U6648 (N_6648,N_3655,N_2946);
xnor U6649 (N_6649,N_4886,N_2414);
nor U6650 (N_6650,N_1298,N_696);
and U6651 (N_6651,N_1091,N_881);
nand U6652 (N_6652,N_2972,N_1459);
and U6653 (N_6653,N_2776,N_1521);
and U6654 (N_6654,N_2950,N_4408);
and U6655 (N_6655,N_2781,N_344);
and U6656 (N_6656,N_4461,N_3890);
and U6657 (N_6657,N_1121,N_3428);
or U6658 (N_6658,N_467,N_1475);
and U6659 (N_6659,N_2906,N_739);
or U6660 (N_6660,N_3276,N_4752);
and U6661 (N_6661,N_269,N_3647);
or U6662 (N_6662,N_4954,N_2269);
and U6663 (N_6663,N_3577,N_1084);
or U6664 (N_6664,N_507,N_1454);
or U6665 (N_6665,N_3451,N_4600);
and U6666 (N_6666,N_961,N_4283);
or U6667 (N_6667,N_4371,N_212);
nand U6668 (N_6668,N_3269,N_4385);
nor U6669 (N_6669,N_237,N_4497);
and U6670 (N_6670,N_3315,N_4784);
or U6671 (N_6671,N_4778,N_1501);
and U6672 (N_6672,N_3608,N_4925);
and U6673 (N_6673,N_1118,N_534);
nand U6674 (N_6674,N_3046,N_4564);
and U6675 (N_6675,N_1718,N_1055);
xor U6676 (N_6676,N_2904,N_4802);
nand U6677 (N_6677,N_4771,N_2550);
nor U6678 (N_6678,N_2285,N_3101);
nor U6679 (N_6679,N_2093,N_2259);
nor U6680 (N_6680,N_864,N_3355);
or U6681 (N_6681,N_2408,N_2433);
nor U6682 (N_6682,N_2172,N_1458);
or U6683 (N_6683,N_2382,N_2283);
and U6684 (N_6684,N_942,N_4996);
nor U6685 (N_6685,N_4024,N_2492);
nor U6686 (N_6686,N_563,N_4870);
nor U6687 (N_6687,N_2449,N_1317);
or U6688 (N_6688,N_3347,N_62);
nor U6689 (N_6689,N_3346,N_4057);
nand U6690 (N_6690,N_415,N_4789);
nand U6691 (N_6691,N_3483,N_3194);
nor U6692 (N_6692,N_4792,N_1509);
or U6693 (N_6693,N_1350,N_3852);
nand U6694 (N_6694,N_2287,N_4526);
and U6695 (N_6695,N_1202,N_94);
xor U6696 (N_6696,N_3978,N_4442);
and U6697 (N_6697,N_4379,N_3536);
or U6698 (N_6698,N_3193,N_3446);
nand U6699 (N_6699,N_1394,N_1129);
nor U6700 (N_6700,N_362,N_713);
or U6701 (N_6701,N_2728,N_4872);
or U6702 (N_6702,N_3790,N_2319);
nor U6703 (N_6703,N_2415,N_2863);
nor U6704 (N_6704,N_4533,N_3581);
and U6705 (N_6705,N_2644,N_917);
nand U6706 (N_6706,N_4001,N_2509);
or U6707 (N_6707,N_2252,N_2601);
nor U6708 (N_6708,N_2495,N_210);
or U6709 (N_6709,N_3817,N_382);
and U6710 (N_6710,N_1111,N_2673);
nor U6711 (N_6711,N_1790,N_2677);
and U6712 (N_6712,N_3279,N_4653);
nand U6713 (N_6713,N_3885,N_940);
or U6714 (N_6714,N_3391,N_3192);
or U6715 (N_6715,N_3390,N_4793);
nor U6716 (N_6716,N_3610,N_1830);
nand U6717 (N_6717,N_637,N_1482);
nand U6718 (N_6718,N_289,N_4783);
or U6719 (N_6719,N_1134,N_3966);
or U6720 (N_6720,N_416,N_1526);
or U6721 (N_6721,N_2701,N_50);
or U6722 (N_6722,N_957,N_1308);
and U6723 (N_6723,N_2046,N_573);
and U6724 (N_6724,N_2917,N_3270);
or U6725 (N_6725,N_7,N_1276);
or U6726 (N_6726,N_3750,N_973);
nor U6727 (N_6727,N_3030,N_653);
nor U6728 (N_6728,N_522,N_4260);
nand U6729 (N_6729,N_459,N_547);
or U6730 (N_6730,N_3278,N_4667);
and U6731 (N_6731,N_1952,N_4693);
and U6732 (N_6732,N_2916,N_3052);
and U6733 (N_6733,N_3172,N_1768);
or U6734 (N_6734,N_1649,N_555);
nor U6735 (N_6735,N_1124,N_2933);
nor U6736 (N_6736,N_3587,N_2734);
or U6737 (N_6737,N_4223,N_3695);
nor U6738 (N_6738,N_3012,N_3368);
and U6739 (N_6739,N_4586,N_4067);
or U6740 (N_6740,N_1123,N_2079);
nand U6741 (N_6741,N_1589,N_3650);
nand U6742 (N_6742,N_916,N_1132);
or U6743 (N_6743,N_4672,N_303);
nand U6744 (N_6744,N_4286,N_3748);
or U6745 (N_6745,N_3672,N_4649);
nand U6746 (N_6746,N_2514,N_1543);
or U6747 (N_6747,N_398,N_3857);
and U6748 (N_6748,N_2765,N_1586);
or U6749 (N_6749,N_2108,N_363);
and U6750 (N_6750,N_4179,N_3144);
nand U6751 (N_6751,N_360,N_4576);
nand U6752 (N_6752,N_2233,N_2142);
nor U6753 (N_6753,N_4674,N_3068);
and U6754 (N_6754,N_2518,N_4026);
or U6755 (N_6755,N_1971,N_2607);
nand U6756 (N_6756,N_43,N_3173);
nor U6757 (N_6757,N_1004,N_4645);
nand U6758 (N_6758,N_3163,N_68);
or U6759 (N_6759,N_3155,N_4588);
and U6760 (N_6760,N_3181,N_155);
nor U6761 (N_6761,N_1461,N_1750);
or U6762 (N_6762,N_3069,N_4411);
and U6763 (N_6763,N_2920,N_4524);
and U6764 (N_6764,N_4911,N_3624);
nand U6765 (N_6765,N_1092,N_3129);
and U6766 (N_6766,N_1837,N_2022);
nand U6767 (N_6767,N_3306,N_3620);
and U6768 (N_6768,N_4339,N_4892);
nor U6769 (N_6769,N_4168,N_3084);
nor U6770 (N_6770,N_471,N_1878);
nand U6771 (N_6771,N_3006,N_1204);
nor U6772 (N_6772,N_1968,N_3636);
or U6773 (N_6773,N_2557,N_606);
and U6774 (N_6774,N_1799,N_52);
and U6775 (N_6775,N_2613,N_1994);
nor U6776 (N_6776,N_396,N_189);
and U6777 (N_6777,N_3393,N_3412);
nor U6778 (N_6778,N_3965,N_915);
and U6779 (N_6779,N_2389,N_1238);
nand U6780 (N_6780,N_4396,N_3242);
nand U6781 (N_6781,N_3402,N_1506);
nor U6782 (N_6782,N_121,N_3205);
nor U6783 (N_6783,N_3465,N_4301);
nand U6784 (N_6784,N_4529,N_3611);
nor U6785 (N_6785,N_1813,N_2690);
nor U6786 (N_6786,N_314,N_4270);
or U6787 (N_6787,N_1145,N_446);
nand U6788 (N_6788,N_1647,N_1398);
nor U6789 (N_6789,N_14,N_3441);
nor U6790 (N_6790,N_1805,N_4958);
xnor U6791 (N_6791,N_557,N_1809);
and U6792 (N_6792,N_1619,N_1728);
or U6793 (N_6793,N_4977,N_4173);
nand U6794 (N_6794,N_4218,N_4573);
or U6795 (N_6795,N_4629,N_2333);
and U6796 (N_6796,N_898,N_2242);
nand U6797 (N_6797,N_2348,N_8);
nand U6798 (N_6798,N_662,N_2763);
or U6799 (N_6799,N_2311,N_1452);
nand U6800 (N_6800,N_1090,N_2026);
and U6801 (N_6801,N_1985,N_1588);
xnor U6802 (N_6802,N_4779,N_2635);
and U6803 (N_6803,N_3894,N_1615);
nand U6804 (N_6804,N_1174,N_634);
nor U6805 (N_6805,N_4402,N_4965);
nor U6806 (N_6806,N_4400,N_233);
nor U6807 (N_6807,N_1244,N_3812);
or U6808 (N_6808,N_1267,N_632);
and U6809 (N_6809,N_3835,N_1912);
or U6810 (N_6810,N_837,N_1116);
nand U6811 (N_6811,N_2071,N_4585);
or U6812 (N_6812,N_1021,N_4927);
nand U6813 (N_6813,N_3831,N_2858);
and U6814 (N_6814,N_3213,N_4542);
and U6815 (N_6815,N_2973,N_3421);
nor U6816 (N_6816,N_1550,N_2926);
or U6817 (N_6817,N_2145,N_1023);
nor U6818 (N_6818,N_721,N_4209);
nor U6819 (N_6819,N_660,N_1008);
and U6820 (N_6820,N_2732,N_1136);
nor U6821 (N_6821,N_246,N_484);
nand U6822 (N_6822,N_218,N_4298);
nor U6823 (N_6823,N_1255,N_2154);
or U6824 (N_6824,N_2156,N_151);
nand U6825 (N_6825,N_587,N_4202);
nor U6826 (N_6826,N_3386,N_1552);
and U6827 (N_6827,N_4015,N_4842);
and U6828 (N_6828,N_18,N_4170);
or U6829 (N_6829,N_2231,N_2812);
nand U6830 (N_6830,N_880,N_4555);
nand U6831 (N_6831,N_4595,N_592);
and U6832 (N_6832,N_843,N_3481);
nand U6833 (N_6833,N_1653,N_3175);
or U6834 (N_6834,N_1782,N_1714);
nor U6835 (N_6835,N_2543,N_319);
or U6836 (N_6836,N_3511,N_2857);
or U6837 (N_6837,N_389,N_4008);
and U6838 (N_6838,N_2021,N_707);
or U6839 (N_6839,N_2563,N_288);
xnor U6840 (N_6840,N_325,N_2191);
or U6841 (N_6841,N_1756,N_3541);
and U6842 (N_6842,N_686,N_3053);
nor U6843 (N_6843,N_2779,N_57);
and U6844 (N_6844,N_1843,N_924);
or U6845 (N_6845,N_1415,N_2054);
nand U6846 (N_6846,N_1922,N_337);
and U6847 (N_6847,N_3710,N_4480);
and U6848 (N_6848,N_4375,N_1804);
and U6849 (N_6849,N_3002,N_3638);
nor U6850 (N_6850,N_71,N_4111);
or U6851 (N_6851,N_1861,N_129);
or U6852 (N_6852,N_1851,N_2270);
or U6853 (N_6853,N_2442,N_718);
or U6854 (N_6854,N_2832,N_1719);
and U6855 (N_6855,N_132,N_1866);
nand U6856 (N_6856,N_2103,N_1737);
or U6857 (N_6857,N_798,N_4604);
and U6858 (N_6858,N_2003,N_369);
nor U6859 (N_6859,N_1171,N_4222);
nand U6860 (N_6860,N_4988,N_3145);
nand U6861 (N_6861,N_2282,N_2706);
or U6862 (N_6862,N_4360,N_745);
nand U6863 (N_6863,N_4256,N_3531);
nor U6864 (N_6864,N_260,N_1673);
and U6865 (N_6865,N_1289,N_3555);
or U6866 (N_6866,N_3999,N_731);
and U6867 (N_6867,N_4059,N_3493);
and U6868 (N_6868,N_1612,N_786);
or U6869 (N_6869,N_4083,N_1580);
nor U6870 (N_6870,N_1969,N_3473);
or U6871 (N_6871,N_799,N_1377);
or U6872 (N_6872,N_4071,N_4696);
or U6873 (N_6873,N_806,N_511);
xor U6874 (N_6874,N_2898,N_1798);
nor U6875 (N_6875,N_3729,N_1052);
and U6876 (N_6876,N_3313,N_1020);
and U6877 (N_6877,N_2207,N_1297);
and U6878 (N_6878,N_251,N_1165);
or U6879 (N_6879,N_1198,N_1613);
nor U6880 (N_6880,N_491,N_4715);
and U6881 (N_6881,N_1206,N_4025);
and U6882 (N_6882,N_2841,N_1024);
or U6883 (N_6883,N_4796,N_2281);
nand U6884 (N_6884,N_4070,N_4205);
nor U6885 (N_6885,N_4142,N_4440);
xor U6886 (N_6886,N_42,N_385);
or U6887 (N_6887,N_727,N_4040);
or U6888 (N_6888,N_4592,N_4930);
or U6889 (N_6889,N_4398,N_4208);
or U6890 (N_6890,N_2526,N_890);
nor U6891 (N_6891,N_2957,N_2086);
or U6892 (N_6892,N_3118,N_4788);
and U6893 (N_6893,N_2248,N_3844);
nor U6894 (N_6894,N_841,N_2166);
nor U6895 (N_6895,N_3819,N_3180);
nor U6896 (N_6896,N_3646,N_4740);
and U6897 (N_6897,N_710,N_1085);
or U6898 (N_6898,N_821,N_1237);
or U6899 (N_6899,N_1438,N_1430);
nor U6900 (N_6900,N_4120,N_3896);
or U6901 (N_6901,N_3848,N_4268);
or U6902 (N_6902,N_3923,N_1119);
and U6903 (N_6903,N_1074,N_3195);
and U6904 (N_6904,N_4519,N_270);
nand U6905 (N_6905,N_1942,N_3249);
nor U6906 (N_6906,N_4178,N_2257);
or U6907 (N_6907,N_1371,N_3128);
nor U6908 (N_6908,N_2874,N_2987);
and U6909 (N_6909,N_663,N_313);
nor U6910 (N_6910,N_2569,N_4756);
nor U6911 (N_6911,N_3396,N_2160);
nor U6912 (N_6912,N_450,N_4748);
nor U6913 (N_6913,N_256,N_29);
xor U6914 (N_6914,N_3680,N_3321);
or U6915 (N_6915,N_1687,N_3561);
nand U6916 (N_6916,N_483,N_2002);
and U6917 (N_6917,N_2256,N_3716);
nand U6918 (N_6918,N_320,N_1857);
and U6919 (N_6919,N_1354,N_3253);
nand U6920 (N_6920,N_1219,N_2696);
or U6921 (N_6921,N_617,N_2326);
nand U6922 (N_6922,N_2755,N_2621);
xnor U6923 (N_6923,N_196,N_2969);
and U6924 (N_6924,N_4668,N_1542);
or U6925 (N_6925,N_3323,N_3109);
nor U6926 (N_6926,N_2932,N_2210);
and U6927 (N_6927,N_927,N_516);
and U6928 (N_6928,N_1449,N_76);
nor U6929 (N_6929,N_1513,N_3505);
nor U6930 (N_6930,N_2773,N_2310);
or U6931 (N_6931,N_4470,N_2910);
and U6932 (N_6932,N_1775,N_4597);
nor U6933 (N_6933,N_28,N_3740);
nor U6934 (N_6934,N_4646,N_542);
nand U6935 (N_6935,N_236,N_4122);
or U6936 (N_6936,N_3077,N_3064);
nor U6937 (N_6937,N_4002,N_102);
nand U6938 (N_6938,N_175,N_1677);
and U6939 (N_6939,N_1989,N_4029);
nand U6940 (N_6940,N_1235,N_614);
or U6941 (N_6941,N_4703,N_2398);
and U6942 (N_6942,N_3797,N_370);
nor U6943 (N_6943,N_4030,N_2551);
and U6944 (N_6944,N_4590,N_2078);
and U6945 (N_6945,N_4723,N_1221);
nor U6946 (N_6946,N_4422,N_4359);
nor U6947 (N_6947,N_3849,N_2960);
nand U6948 (N_6948,N_4913,N_4415);
nand U6949 (N_6949,N_3398,N_4447);
and U6950 (N_6950,N_272,N_3903);
nor U6951 (N_6951,N_4637,N_3434);
nand U6952 (N_6952,N_4931,N_321);
and U6953 (N_6953,N_359,N_610);
nor U6954 (N_6954,N_1335,N_2618);
nor U6955 (N_6955,N_579,N_4481);
nand U6956 (N_6956,N_2434,N_78);
or U6957 (N_6957,N_2687,N_1629);
nand U6958 (N_6958,N_4990,N_3630);
nand U6959 (N_6959,N_4354,N_4389);
or U6960 (N_6960,N_2332,N_169);
and U6961 (N_6961,N_4206,N_3640);
nor U6962 (N_6962,N_1242,N_1563);
nor U6963 (N_6963,N_2379,N_4229);
nor U6964 (N_6964,N_4939,N_1659);
nor U6965 (N_6965,N_4043,N_1311);
and U6966 (N_6966,N_230,N_2821);
nor U6967 (N_6967,N_1224,N_929);
nand U6968 (N_6968,N_3609,N_1115);
nor U6969 (N_6969,N_2122,N_2944);
nand U6970 (N_6970,N_3767,N_846);
nor U6971 (N_6971,N_3027,N_1368);
and U6972 (N_6972,N_2275,N_2330);
nand U6973 (N_6973,N_3107,N_4602);
nand U6974 (N_6974,N_277,N_1102);
nand U6975 (N_6975,N_2853,N_989);
and U6976 (N_6976,N_4265,N_2306);
or U6977 (N_6977,N_481,N_4655);
nor U6978 (N_6978,N_699,N_2891);
and U6979 (N_6979,N_347,N_3309);
nor U6980 (N_6980,N_1609,N_2703);
or U6981 (N_6981,N_2846,N_4660);
nand U6982 (N_6982,N_4934,N_437);
or U6983 (N_6983,N_3318,N_538);
nand U6984 (N_6984,N_3933,N_4115);
and U6985 (N_6985,N_1777,N_2125);
nand U6986 (N_6986,N_722,N_670);
or U6987 (N_6987,N_1259,N_1166);
nor U6988 (N_6988,N_2239,N_1423);
nor U6989 (N_6989,N_3384,N_36);
nand U6990 (N_6990,N_1741,N_4478);
or U6991 (N_6991,N_2063,N_1282);
nand U6992 (N_6992,N_2102,N_381);
nor U6993 (N_6993,N_2651,N_399);
and U6994 (N_6994,N_2499,N_2531);
and U6995 (N_6995,N_585,N_2961);
nor U6996 (N_6996,N_3727,N_1735);
nor U6997 (N_6997,N_353,N_4418);
nor U6998 (N_6998,N_4215,N_2784);
and U6999 (N_6999,N_3989,N_4835);
nand U7000 (N_7000,N_554,N_1848);
or U7001 (N_7001,N_4088,N_2096);
nor U7002 (N_7002,N_209,N_216);
and U7003 (N_7003,N_1639,N_187);
nand U7004 (N_7004,N_1463,N_4686);
and U7005 (N_7005,N_3184,N_1387);
or U7006 (N_7006,N_502,N_790);
and U7007 (N_7007,N_2174,N_2100);
and U7008 (N_7008,N_569,N_3827);
nor U7009 (N_7009,N_4144,N_4518);
nand U7010 (N_7010,N_4705,N_3671);
or U7011 (N_7011,N_3023,N_4801);
nand U7012 (N_7012,N_3779,N_2223);
or U7013 (N_7013,N_855,N_2510);
or U7014 (N_7014,N_13,N_4322);
nand U7015 (N_7015,N_4321,N_736);
and U7016 (N_7016,N_141,N_683);
nor U7017 (N_7017,N_2292,N_4393);
and U7018 (N_7018,N_876,N_3016);
and U7019 (N_7019,N_1662,N_1876);
nor U7020 (N_7020,N_3659,N_2338);
or U7021 (N_7021,N_3662,N_1854);
nand U7022 (N_7022,N_2370,N_1019);
and U7023 (N_7023,N_3571,N_1879);
or U7024 (N_7024,N_4330,N_3616);
and U7025 (N_7025,N_1285,N_3125);
or U7026 (N_7026,N_2029,N_4444);
and U7027 (N_7027,N_4535,N_742);
and U7028 (N_7028,N_3556,N_4022);
and U7029 (N_7029,N_1796,N_4405);
nor U7030 (N_7030,N_4915,N_3940);
nand U7031 (N_7031,N_338,N_4750);
nand U7032 (N_7032,N_4128,N_249);
nand U7033 (N_7033,N_3991,N_3267);
xnor U7034 (N_7034,N_4441,N_1532);
nor U7035 (N_7035,N_1099,N_4313);
or U7036 (N_7036,N_1954,N_182);
or U7037 (N_7037,N_3476,N_3544);
nand U7038 (N_7038,N_4409,N_1696);
or U7039 (N_7039,N_3572,N_4316);
nand U7040 (N_7040,N_564,N_3211);
nor U7041 (N_7041,N_2780,N_2815);
nor U7042 (N_7042,N_2733,N_2642);
and U7043 (N_7043,N_72,N_1643);
nor U7044 (N_7044,N_1627,N_4810);
or U7045 (N_7045,N_906,N_154);
or U7046 (N_7046,N_2138,N_3509);
nand U7047 (N_7047,N_3868,N_2541);
or U7048 (N_7048,N_474,N_387);
nand U7049 (N_7049,N_3498,N_956);
or U7050 (N_7050,N_2324,N_1156);
and U7051 (N_7051,N_4890,N_3612);
and U7052 (N_7052,N_2121,N_3099);
or U7053 (N_7053,N_2700,N_774);
nand U7054 (N_7054,N_203,N_3899);
nand U7055 (N_7055,N_4540,N_3864);
and U7056 (N_7056,N_1511,N_4832);
nor U7057 (N_7057,N_2842,N_308);
or U7058 (N_7058,N_2500,N_4848);
nand U7059 (N_7059,N_3199,N_1471);
nor U7060 (N_7060,N_4799,N_3863);
nor U7061 (N_7061,N_1251,N_1941);
and U7062 (N_7062,N_2413,N_4499);
or U7063 (N_7063,N_2177,N_2777);
xnor U7064 (N_7064,N_4503,N_2303);
nor U7065 (N_7065,N_3717,N_4278);
and U7066 (N_7066,N_4843,N_2667);
nand U7067 (N_7067,N_969,N_2736);
nor U7068 (N_7068,N_2694,N_4345);
nand U7069 (N_7069,N_801,N_4508);
nand U7070 (N_7070,N_1245,N_4104);
nor U7071 (N_7071,N_3956,N_2195);
nor U7072 (N_7072,N_2561,N_3154);
and U7073 (N_7073,N_2831,N_2794);
or U7074 (N_7074,N_3244,N_2953);
and U7075 (N_7075,N_2190,N_3227);
and U7076 (N_7076,N_3011,N_425);
and U7077 (N_7077,N_1911,N_4473);
and U7078 (N_7078,N_4187,N_2560);
nor U7079 (N_7079,N_2661,N_4271);
and U7080 (N_7080,N_1927,N_4482);
or U7081 (N_7081,N_932,N_3097);
nor U7082 (N_7082,N_2010,N_408);
and U7083 (N_7083,N_2163,N_4055);
nor U7084 (N_7084,N_3523,N_2188);
and U7085 (N_7085,N_126,N_1263);
nor U7086 (N_7086,N_4867,N_601);
nor U7087 (N_7087,N_965,N_286);
nor U7088 (N_7088,N_1313,N_1499);
nand U7089 (N_7089,N_3535,N_1049);
nand U7090 (N_7090,N_2052,N_117);
and U7091 (N_7091,N_788,N_4797);
nor U7092 (N_7092,N_4878,N_2179);
nand U7093 (N_7093,N_4394,N_3643);
or U7094 (N_7094,N_4736,N_3679);
nand U7095 (N_7095,N_3124,N_3438);
and U7096 (N_7096,N_3977,N_2689);
nor U7097 (N_7097,N_1015,N_597);
nand U7098 (N_7098,N_3370,N_3471);
nand U7099 (N_7099,N_4274,N_4530);
nor U7100 (N_7100,N_4403,N_3389);
nor U7101 (N_7101,N_3369,N_3970);
and U7102 (N_7102,N_4699,N_3629);
and U7103 (N_7103,N_4852,N_46);
or U7104 (N_7104,N_2525,N_4110);
nand U7105 (N_7105,N_2131,N_2485);
nand U7106 (N_7106,N_3049,N_298);
or U7107 (N_7107,N_2769,N_1467);
and U7108 (N_7108,N_2365,N_526);
or U7109 (N_7109,N_933,N_1030);
nand U7110 (N_7110,N_4982,N_3862);
nor U7111 (N_7111,N_3814,N_34);
nor U7112 (N_7112,N_4956,N_3475);
nor U7113 (N_7113,N_1309,N_4141);
nor U7114 (N_7114,N_3418,N_3168);
nand U7115 (N_7115,N_3110,N_4941);
nand U7116 (N_7116,N_3828,N_1450);
nor U7117 (N_7117,N_198,N_1075);
nor U7118 (N_7118,N_2399,N_3357);
and U7119 (N_7119,N_2261,N_376);
nor U7120 (N_7120,N_2565,N_1984);
nor U7121 (N_7121,N_4657,N_146);
or U7122 (N_7122,N_3566,N_1562);
or U7123 (N_7123,N_2721,N_1400);
nand U7124 (N_7124,N_1633,N_1253);
nand U7125 (N_7125,N_1698,N_2872);
nand U7126 (N_7126,N_1039,N_1871);
nand U7127 (N_7127,N_4538,N_3317);
and U7128 (N_7128,N_1399,N_4641);
nand U7129 (N_7129,N_4973,N_3542);
and U7130 (N_7130,N_701,N_546);
nor U7131 (N_7131,N_4459,N_1784);
nand U7132 (N_7132,N_1487,N_583);
nor U7133 (N_7133,N_2921,N_2452);
or U7134 (N_7134,N_3527,N_2505);
and U7135 (N_7135,N_2043,N_1909);
or U7136 (N_7136,N_2197,N_4896);
nand U7137 (N_7137,N_1386,N_3916);
or U7138 (N_7138,N_490,N_2778);
nor U7139 (N_7139,N_48,N_3576);
nand U7140 (N_7140,N_162,N_607);
or U7141 (N_7141,N_3007,N_2681);
nand U7142 (N_7142,N_768,N_3374);
nand U7143 (N_7143,N_2682,N_3651);
and U7144 (N_7144,N_3406,N_4685);
and U7145 (N_7145,N_3574,N_3780);
or U7146 (N_7146,N_4063,N_2692);
and U7147 (N_7147,N_4853,N_4302);
nand U7148 (N_7148,N_1835,N_421);
or U7149 (N_7149,N_173,N_3336);
and U7150 (N_7150,N_2892,N_562);
nand U7151 (N_7151,N_3822,N_646);
or U7152 (N_7152,N_1690,N_830);
nand U7153 (N_7153,N_3530,N_1665);
nand U7154 (N_7154,N_708,N_4869);
and U7155 (N_7155,N_3437,N_2180);
and U7156 (N_7156,N_1320,N_1559);
and U7157 (N_7157,N_348,N_2806);
nand U7158 (N_7158,N_1738,N_621);
or U7159 (N_7159,N_638,N_1125);
nand U7160 (N_7160,N_1974,N_4050);
nor U7161 (N_7161,N_4822,N_4262);
nand U7162 (N_7162,N_3506,N_4993);
and U7163 (N_7163,N_2631,N_206);
nand U7164 (N_7164,N_1993,N_2377);
and U7165 (N_7165,N_3161,N_1701);
and U7166 (N_7166,N_1900,N_752);
or U7167 (N_7167,N_1739,N_3533);
nor U7168 (N_7168,N_3593,N_4027);
nor U7169 (N_7169,N_4253,N_4730);
and U7170 (N_7170,N_862,N_2870);
or U7171 (N_7171,N_309,N_4161);
nor U7172 (N_7172,N_726,N_3152);
or U7173 (N_7173,N_4353,N_4871);
nor U7174 (N_7174,N_2273,N_1122);
and U7175 (N_7175,N_2574,N_3634);
and U7176 (N_7176,N_536,N_3031);
or U7177 (N_7177,N_1764,N_3855);
or U7178 (N_7178,N_2606,N_2322);
nor U7179 (N_7179,N_1743,N_4373);
nand U7180 (N_7180,N_4624,N_4768);
nor U7181 (N_7181,N_3615,N_2033);
and U7182 (N_7182,N_2050,N_911);
nor U7183 (N_7183,N_2936,N_4172);
or U7184 (N_7184,N_4328,N_10);
or U7185 (N_7185,N_4130,N_920);
or U7186 (N_7186,N_1704,N_4644);
nand U7187 (N_7187,N_253,N_3436);
and U7188 (N_7188,N_3954,N_1921);
or U7189 (N_7189,N_1043,N_4068);
or U7190 (N_7190,N_4,N_1217);
nand U7191 (N_7191,N_1800,N_1591);
and U7192 (N_7192,N_1620,N_3793);
xnor U7193 (N_7193,N_23,N_2626);
and U7194 (N_7194,N_1601,N_1820);
nor U7195 (N_7195,N_3895,N_779);
nor U7196 (N_7196,N_2675,N_2752);
or U7197 (N_7197,N_2581,N_2361);
nand U7198 (N_7198,N_623,N_2031);
and U7199 (N_7199,N_3353,N_4898);
nand U7200 (N_7200,N_4243,N_2649);
nand U7201 (N_7201,N_2451,N_1575);
nand U7202 (N_7202,N_1248,N_4702);
nand U7203 (N_7203,N_921,N_3114);
and U7204 (N_7204,N_4905,N_1631);
nand U7205 (N_7205,N_4182,N_856);
and U7206 (N_7206,N_2341,N_2296);
nand U7207 (N_7207,N_3450,N_2980);
and U7208 (N_7208,N_3137,N_1530);
or U7209 (N_7209,N_2293,N_4615);
or U7210 (N_7210,N_1744,N_1512);
nor U7211 (N_7211,N_4308,N_2441);
and U7212 (N_7212,N_1038,N_2498);
nor U7213 (N_7213,N_3167,N_918);
and U7214 (N_7214,N_172,N_1691);
nand U7215 (N_7215,N_1340,N_4633);
and U7216 (N_7216,N_3356,N_950);
or U7217 (N_7217,N_3719,N_3515);
nand U7218 (N_7218,N_1596,N_1246);
and U7219 (N_7219,N_3661,N_1154);
and U7220 (N_7220,N_1558,N_1555);
nor U7221 (N_7221,N_4953,N_4414);
and U7222 (N_7222,N_4720,N_1042);
nand U7223 (N_7223,N_1621,N_3248);
or U7224 (N_7224,N_1841,N_1606);
or U7225 (N_7225,N_1614,N_1937);
nand U7226 (N_7226,N_964,N_3495);
or U7227 (N_7227,N_2835,N_3017);
and U7228 (N_7228,N_1291,N_2258);
nor U7229 (N_7229,N_1178,N_3250);
nor U7230 (N_7230,N_4081,N_4983);
or U7231 (N_7231,N_3938,N_3381);
or U7232 (N_7232,N_2178,N_1406);
and U7233 (N_7233,N_2603,N_1275);
nand U7234 (N_7234,N_2081,N_664);
and U7235 (N_7235,N_139,N_3151);
or U7236 (N_7236,N_2825,N_3501);
and U7237 (N_7237,N_1566,N_3050);
or U7238 (N_7238,N_873,N_3732);
nand U7239 (N_7239,N_1190,N_3586);
and U7240 (N_7240,N_342,N_3724);
or U7241 (N_7241,N_3351,N_4735);
and U7242 (N_7242,N_3918,N_836);
nand U7243 (N_7243,N_4803,N_4407);
xor U7244 (N_7244,N_4236,N_2534);
or U7245 (N_7245,N_2411,N_2235);
or U7246 (N_7246,N_4309,N_395);
and U7247 (N_7247,N_2602,N_1486);
nand U7248 (N_7248,N_1053,N_789);
nand U7249 (N_7249,N_2688,N_999);
nor U7250 (N_7250,N_2000,N_341);
or U7251 (N_7251,N_4762,N_75);
and U7252 (N_7252,N_3061,N_1811);
nand U7253 (N_7253,N_3910,N_4149);
nand U7254 (N_7254,N_170,N_3948);
or U7255 (N_7255,N_345,N_574);
or U7256 (N_7256,N_2274,N_3488);
nand U7257 (N_7257,N_1240,N_861);
nand U7258 (N_7258,N_760,N_4140);
and U7259 (N_7259,N_3585,N_586);
nor U7260 (N_7260,N_2471,N_2597);
or U7261 (N_7261,N_4020,N_4772);
nor U7262 (N_7262,N_4343,N_2678);
and U7263 (N_7263,N_588,N_1553);
or U7264 (N_7264,N_478,N_687);
or U7265 (N_7265,N_4677,N_4625);
nor U7266 (N_7266,N_3082,N_3146);
and U7267 (N_7267,N_3537,N_305);
nand U7268 (N_7268,N_955,N_1274);
and U7269 (N_7269,N_2718,N_2124);
and U7270 (N_7270,N_2556,N_300);
nand U7271 (N_7271,N_1727,N_748);
and U7272 (N_7272,N_3753,N_4041);
xor U7273 (N_7273,N_937,N_2887);
and U7274 (N_7274,N_330,N_4429);
nor U7275 (N_7275,N_2313,N_952);
nand U7276 (N_7276,N_384,N_2457);
and U7277 (N_7277,N_2278,N_2132);
or U7278 (N_7278,N_3798,N_3874);
nand U7279 (N_7279,N_2762,N_1872);
nor U7280 (N_7280,N_1002,N_2501);
or U7281 (N_7281,N_2652,N_3251);
nand U7282 (N_7282,N_2305,N_427);
nand U7283 (N_7283,N_2686,N_3902);
and U7284 (N_7284,N_1453,N_652);
nand U7285 (N_7285,N_702,N_468);
or U7286 (N_7286,N_1894,N_636);
or U7287 (N_7287,N_4457,N_1959);
nor U7288 (N_7288,N_3135,N_3920);
nand U7289 (N_7289,N_2068,N_4066);
nor U7290 (N_7290,N_2406,N_2968);
and U7291 (N_7291,N_3003,N_1302);
or U7292 (N_7292,N_3058,N_3644);
nor U7293 (N_7293,N_2559,N_3575);
xor U7294 (N_7294,N_1898,N_3637);
nand U7295 (N_7295,N_2964,N_2674);
nor U7296 (N_7296,N_3580,N_1382);
nor U7297 (N_7297,N_3700,N_232);
nor U7298 (N_7298,N_761,N_2844);
nand U7299 (N_7299,N_90,N_4999);
nand U7300 (N_7300,N_978,N_4314);
nor U7301 (N_7301,N_4865,N_1147);
nor U7302 (N_7302,N_2800,N_581);
nand U7303 (N_7303,N_1462,N_1734);
nor U7304 (N_7304,N_2087,N_1000);
nor U7305 (N_7305,N_2314,N_612);
nor U7306 (N_7306,N_3185,N_4559);
nor U7307 (N_7307,N_3884,N_318);
xor U7308 (N_7308,N_136,N_813);
nand U7309 (N_7309,N_2394,N_2130);
nor U7310 (N_7310,N_3376,N_3342);
and U7311 (N_7311,N_2118,N_1480);
and U7312 (N_7312,N_3208,N_56);
or U7313 (N_7313,N_794,N_1239);
or U7314 (N_7314,N_4109,N_515);
nand U7315 (N_7315,N_2903,N_1832);
nor U7316 (N_7316,N_4544,N_327);
nor U7317 (N_7317,N_2532,N_1149);
nand U7318 (N_7318,N_1139,N_2450);
or U7319 (N_7319,N_2793,N_1694);
nand U7320 (N_7320,N_635,N_778);
nor U7321 (N_7321,N_2342,N_4631);
nor U7322 (N_7322,N_4233,N_2279);
or U7323 (N_7323,N_1600,N_4885);
or U7324 (N_7324,N_1234,N_41);
or U7325 (N_7325,N_2008,N_4119);
nand U7326 (N_7326,N_2595,N_4670);
nand U7327 (N_7327,N_1167,N_3998);
nand U7328 (N_7328,N_4074,N_3426);
and U7329 (N_7329,N_2114,N_1353);
or U7330 (N_7330,N_180,N_1227);
nand U7331 (N_7331,N_1754,N_834);
and U7332 (N_7332,N_2249,N_3364);
nand U7333 (N_7333,N_2357,N_215);
nor U7334 (N_7334,N_176,N_4093);
and U7335 (N_7335,N_1409,N_676);
nor U7336 (N_7336,N_827,N_51);
nand U7337 (N_7337,N_2318,N_1822);
nand U7338 (N_7338,N_3358,N_1022);
nand U7339 (N_7339,N_1827,N_2246);
and U7340 (N_7340,N_4866,N_3723);
nor U7341 (N_7341,N_371,N_1745);
and U7342 (N_7342,N_850,N_3962);
and U7343 (N_7343,N_61,N_2395);
or U7344 (N_7344,N_4139,N_1570);
nor U7345 (N_7345,N_3160,N_1188);
nand U7346 (N_7346,N_420,N_983);
and U7347 (N_7347,N_2852,N_4971);
nand U7348 (N_7348,N_2823,N_4512);
and U7349 (N_7349,N_4297,N_3674);
or U7350 (N_7350,N_1802,N_520);
nor U7351 (N_7351,N_2443,N_2315);
or U7352 (N_7352,N_2265,N_32);
and U7353 (N_7353,N_2822,N_716);
nor U7354 (N_7354,N_4681,N_2977);
and U7355 (N_7355,N_1385,N_1625);
or U7356 (N_7356,N_4416,N_4255);
or U7357 (N_7357,N_2266,N_3463);
nor U7358 (N_7358,N_3906,N_643);
or U7359 (N_7359,N_2918,N_4183);
nor U7360 (N_7360,N_3712,N_2940);
nand U7361 (N_7361,N_275,N_3308);
and U7362 (N_7362,N_2445,N_2323);
or U7363 (N_7363,N_2201,N_3344);
nor U7364 (N_7364,N_3123,N_2575);
and U7365 (N_7365,N_3795,N_1634);
nand U7366 (N_7366,N_4650,N_2702);
or U7367 (N_7367,N_4097,N_1906);
and U7368 (N_7368,N_1445,N_1128);
and U7369 (N_7369,N_2975,N_457);
and U7370 (N_7370,N_2630,N_4235);
and U7371 (N_7371,N_3104,N_499);
or U7372 (N_7372,N_4225,N_992);
nor U7373 (N_7373,N_1363,N_1545);
nand U7374 (N_7374,N_4060,N_4836);
nor U7375 (N_7375,N_4234,N_11);
or U7376 (N_7376,N_4749,N_4331);
or U7377 (N_7377,N_287,N_3872);
nor U7378 (N_7378,N_2294,N_2475);
nor U7379 (N_7379,N_4475,N_3702);
and U7380 (N_7380,N_693,N_1624);
nor U7381 (N_7381,N_814,N_4887);
nor U7382 (N_7382,N_3235,N_69);
nor U7383 (N_7383,N_558,N_3613);
or U7384 (N_7384,N_2582,N_4102);
and U7385 (N_7385,N_2860,N_694);
xnor U7386 (N_7386,N_2170,N_3074);
nand U7387 (N_7387,N_1456,N_2513);
nand U7388 (N_7388,N_1988,N_257);
or U7389 (N_7389,N_4489,N_1261);
or U7390 (N_7390,N_250,N_1484);
and U7391 (N_7391,N_849,N_4451);
and U7392 (N_7392,N_1710,N_1697);
or U7393 (N_7393,N_358,N_1672);
nand U7394 (N_7394,N_4903,N_966);
or U7395 (N_7395,N_4814,N_4281);
and U7396 (N_7396,N_4816,N_3442);
nand U7397 (N_7397,N_3044,N_2018);
nand U7398 (N_7398,N_4935,N_2782);
nand U7399 (N_7399,N_3614,N_2119);
nand U7400 (N_7400,N_3024,N_4684);
or U7401 (N_7401,N_1303,N_3409);
or U7402 (N_7402,N_1995,N_1336);
nor U7403 (N_7403,N_1582,N_1140);
nor U7404 (N_7404,N_2660,N_2897);
nor U7405 (N_7405,N_1359,N_4651);
and U7406 (N_7406,N_1107,N_422);
or U7407 (N_7407,N_1765,N_4466);
or U7408 (N_7408,N_1548,N_4565);
nand U7409 (N_7409,N_3528,N_3588);
or U7410 (N_7410,N_96,N_4523);
and U7411 (N_7411,N_1534,N_4477);
or U7412 (N_7412,N_3191,N_1681);
nor U7413 (N_7413,N_3945,N_2914);
or U7414 (N_7414,N_689,N_3766);
nand U7415 (N_7415,N_2544,N_4427);
or U7416 (N_7416,N_192,N_971);
and U7417 (N_7417,N_887,N_1829);
or U7418 (N_7418,N_1173,N_1914);
or U7419 (N_7419,N_3469,N_3968);
nor U7420 (N_7420,N_3992,N_835);
nor U7421 (N_7421,N_4947,N_2586);
and U7422 (N_7422,N_3986,N_1413);
nand U7423 (N_7423,N_970,N_1265);
nand U7424 (N_7424,N_4923,N_2604);
and U7425 (N_7425,N_553,N_4900);
and U7426 (N_7426,N_3944,N_2856);
or U7427 (N_7427,N_561,N_3980);
or U7428 (N_7428,N_4804,N_2671);
and U7429 (N_7429,N_1630,N_1001);
or U7430 (N_7430,N_1787,N_3594);
nor U7431 (N_7431,N_530,N_590);
nor U7432 (N_7432,N_4484,N_108);
nand U7433 (N_7433,N_284,N_2076);
and U7434 (N_7434,N_503,N_1571);
or U7435 (N_7435,N_2061,N_4962);
nand U7436 (N_7436,N_3905,N_113);
or U7437 (N_7437,N_2623,N_3830);
or U7438 (N_7438,N_654,N_1356);
nand U7439 (N_7439,N_1207,N_4159);
nand U7440 (N_7440,N_1578,N_3670);
nand U7441 (N_7441,N_3272,N_1381);
and U7442 (N_7442,N_4329,N_1648);
and U7443 (N_7443,N_1384,N_3284);
or U7444 (N_7444,N_2789,N_2663);
nand U7445 (N_7445,N_3352,N_3871);
nand U7446 (N_7446,N_4210,N_4889);
nor U7447 (N_7447,N_1688,N_110);
or U7448 (N_7448,N_4125,N_2419);
nor U7449 (N_7449,N_1808,N_4844);
nor U7450 (N_7450,N_3815,N_2091);
nor U7451 (N_7451,N_3339,N_1568);
or U7452 (N_7452,N_3298,N_519);
nand U7453 (N_7453,N_3486,N_2405);
nand U7454 (N_7454,N_3870,N_3959);
xor U7455 (N_7455,N_4356,N_1757);
nand U7456 (N_7456,N_4786,N_785);
nand U7457 (N_7457,N_692,N_4666);
nand U7458 (N_7458,N_2693,N_4435);
and U7459 (N_7459,N_266,N_3443);
nand U7460 (N_7460,N_1836,N_4031);
nand U7461 (N_7461,N_2048,N_1888);
or U7462 (N_7462,N_1560,N_3435);
nor U7463 (N_7463,N_1241,N_208);
or U7464 (N_7464,N_2346,N_934);
nor U7465 (N_7465,N_4011,N_4162);
and U7466 (N_7466,N_1360,N_1831);
or U7467 (N_7467,N_1963,N_1654);
and U7468 (N_7468,N_1736,N_124);
nor U7469 (N_7469,N_3111,N_2240);
nor U7470 (N_7470,N_3821,N_3799);
nand U7471 (N_7471,N_4152,N_3508);
and U7472 (N_7472,N_4446,N_497);
and U7473 (N_7473,N_2288,N_2051);
or U7474 (N_7474,N_571,N_974);
nand U7475 (N_7475,N_1767,N_4028);
nor U7476 (N_7476,N_4731,N_3681);
nand U7477 (N_7477,N_1473,N_3683);
or U7478 (N_7478,N_2094,N_3365);
or U7479 (N_7479,N_3188,N_1858);
and U7480 (N_7480,N_725,N_4673);
nand U7481 (N_7481,N_4091,N_2672);
nand U7482 (N_7482,N_4758,N_958);
and U7483 (N_7483,N_106,N_1172);
or U7484 (N_7484,N_1926,N_3507);
and U7485 (N_7485,N_4374,N_1663);
nor U7486 (N_7486,N_4358,N_2985);
or U7487 (N_7487,N_413,N_3153);
or U7488 (N_7488,N_791,N_2211);
nand U7489 (N_7489,N_3749,N_1138);
nand U7490 (N_7490,N_2410,N_4207);
nor U7491 (N_7491,N_458,N_2182);
nand U7492 (N_7492,N_4410,N_2707);
and U7493 (N_7493,N_4154,N_4910);
nor U7494 (N_7494,N_3939,N_3686);
nand U7495 (N_7495,N_3806,N_4676);
nand U7496 (N_7496,N_4716,N_1958);
nand U7497 (N_7497,N_2715,N_765);
nand U7498 (N_7498,N_4337,N_3083);
nand U7499 (N_7499,N_263,N_1948);
or U7500 (N_7500,N_4446,N_1029);
nand U7501 (N_7501,N_652,N_3763);
nor U7502 (N_7502,N_2609,N_2301);
or U7503 (N_7503,N_511,N_3601);
nor U7504 (N_7504,N_4885,N_4389);
nor U7505 (N_7505,N_3684,N_3437);
nor U7506 (N_7506,N_1493,N_2093);
nand U7507 (N_7507,N_345,N_3678);
nand U7508 (N_7508,N_1090,N_4050);
nor U7509 (N_7509,N_2828,N_4417);
or U7510 (N_7510,N_4906,N_623);
nand U7511 (N_7511,N_588,N_1588);
and U7512 (N_7512,N_1371,N_1229);
and U7513 (N_7513,N_369,N_3147);
nor U7514 (N_7514,N_3008,N_436);
or U7515 (N_7515,N_3796,N_3651);
and U7516 (N_7516,N_159,N_296);
nor U7517 (N_7517,N_356,N_4967);
or U7518 (N_7518,N_2401,N_4952);
and U7519 (N_7519,N_696,N_1442);
nor U7520 (N_7520,N_1990,N_3412);
and U7521 (N_7521,N_2735,N_1047);
nand U7522 (N_7522,N_53,N_580);
or U7523 (N_7523,N_1786,N_4089);
nor U7524 (N_7524,N_4483,N_2457);
and U7525 (N_7525,N_931,N_4097);
nand U7526 (N_7526,N_4952,N_3745);
nor U7527 (N_7527,N_3385,N_2459);
nand U7528 (N_7528,N_4655,N_2324);
nand U7529 (N_7529,N_2829,N_4643);
nand U7530 (N_7530,N_584,N_2420);
nor U7531 (N_7531,N_935,N_1580);
nor U7532 (N_7532,N_2688,N_4924);
or U7533 (N_7533,N_4013,N_59);
nand U7534 (N_7534,N_2812,N_3627);
nor U7535 (N_7535,N_358,N_750);
nor U7536 (N_7536,N_3667,N_2419);
and U7537 (N_7537,N_2862,N_4667);
and U7538 (N_7538,N_1950,N_437);
or U7539 (N_7539,N_3574,N_1011);
nand U7540 (N_7540,N_3479,N_208);
nand U7541 (N_7541,N_2492,N_1448);
nor U7542 (N_7542,N_2592,N_4104);
nand U7543 (N_7543,N_3246,N_2586);
or U7544 (N_7544,N_1628,N_3511);
or U7545 (N_7545,N_3001,N_4127);
and U7546 (N_7546,N_1603,N_1724);
and U7547 (N_7547,N_2969,N_548);
nor U7548 (N_7548,N_655,N_4275);
or U7549 (N_7549,N_2239,N_488);
nand U7550 (N_7550,N_2914,N_591);
or U7551 (N_7551,N_1732,N_4591);
xnor U7552 (N_7552,N_1034,N_35);
nand U7553 (N_7553,N_4353,N_4562);
and U7554 (N_7554,N_3688,N_3336);
nor U7555 (N_7555,N_4266,N_1328);
nand U7556 (N_7556,N_1839,N_2546);
nor U7557 (N_7557,N_4178,N_4980);
nor U7558 (N_7558,N_2629,N_3692);
nor U7559 (N_7559,N_2268,N_1395);
nor U7560 (N_7560,N_4235,N_952);
nor U7561 (N_7561,N_4053,N_2610);
nand U7562 (N_7562,N_1968,N_837);
and U7563 (N_7563,N_3069,N_3371);
and U7564 (N_7564,N_3569,N_3511);
and U7565 (N_7565,N_3377,N_1839);
and U7566 (N_7566,N_3759,N_1884);
nor U7567 (N_7567,N_3554,N_1614);
nor U7568 (N_7568,N_1914,N_3490);
and U7569 (N_7569,N_4906,N_1667);
nor U7570 (N_7570,N_272,N_3624);
nand U7571 (N_7571,N_2575,N_1801);
nor U7572 (N_7572,N_172,N_4277);
or U7573 (N_7573,N_2197,N_3704);
and U7574 (N_7574,N_3520,N_1961);
nand U7575 (N_7575,N_4644,N_2315);
or U7576 (N_7576,N_805,N_4290);
or U7577 (N_7577,N_4742,N_211);
nand U7578 (N_7578,N_1131,N_1023);
nand U7579 (N_7579,N_1790,N_4044);
nand U7580 (N_7580,N_3635,N_799);
nand U7581 (N_7581,N_1484,N_2244);
nor U7582 (N_7582,N_2625,N_2651);
and U7583 (N_7583,N_1787,N_4264);
and U7584 (N_7584,N_3636,N_906);
or U7585 (N_7585,N_2621,N_3098);
and U7586 (N_7586,N_4116,N_2078);
nand U7587 (N_7587,N_1999,N_569);
and U7588 (N_7588,N_777,N_4670);
and U7589 (N_7589,N_2384,N_4788);
nor U7590 (N_7590,N_4441,N_668);
or U7591 (N_7591,N_1956,N_3790);
nor U7592 (N_7592,N_3270,N_4427);
nor U7593 (N_7593,N_2618,N_2820);
or U7594 (N_7594,N_718,N_4249);
and U7595 (N_7595,N_2142,N_4673);
or U7596 (N_7596,N_4860,N_62);
and U7597 (N_7597,N_1833,N_3564);
or U7598 (N_7598,N_3905,N_431);
or U7599 (N_7599,N_3948,N_3078);
nand U7600 (N_7600,N_4711,N_634);
nand U7601 (N_7601,N_2114,N_3105);
nor U7602 (N_7602,N_2379,N_657);
nand U7603 (N_7603,N_4970,N_430);
or U7604 (N_7604,N_4379,N_485);
nand U7605 (N_7605,N_453,N_469);
or U7606 (N_7606,N_3028,N_4994);
nand U7607 (N_7607,N_2231,N_231);
nand U7608 (N_7608,N_766,N_872);
or U7609 (N_7609,N_2288,N_4507);
or U7610 (N_7610,N_1723,N_898);
or U7611 (N_7611,N_1265,N_4888);
nor U7612 (N_7612,N_4872,N_504);
or U7613 (N_7613,N_4313,N_4452);
nor U7614 (N_7614,N_578,N_2265);
and U7615 (N_7615,N_834,N_2146);
nand U7616 (N_7616,N_4714,N_488);
and U7617 (N_7617,N_761,N_300);
and U7618 (N_7618,N_2427,N_710);
and U7619 (N_7619,N_2047,N_4298);
and U7620 (N_7620,N_3081,N_1013);
nor U7621 (N_7621,N_797,N_273);
or U7622 (N_7622,N_4615,N_2450);
and U7623 (N_7623,N_1201,N_2234);
nor U7624 (N_7624,N_1774,N_838);
or U7625 (N_7625,N_2572,N_1853);
xor U7626 (N_7626,N_1842,N_2408);
nor U7627 (N_7627,N_2335,N_3329);
and U7628 (N_7628,N_1850,N_3749);
nor U7629 (N_7629,N_2847,N_3136);
and U7630 (N_7630,N_1111,N_940);
and U7631 (N_7631,N_3178,N_2294);
nand U7632 (N_7632,N_330,N_2690);
and U7633 (N_7633,N_2916,N_3124);
nor U7634 (N_7634,N_749,N_3897);
and U7635 (N_7635,N_1985,N_2428);
or U7636 (N_7636,N_4458,N_4961);
nor U7637 (N_7637,N_2855,N_1718);
or U7638 (N_7638,N_3054,N_3784);
and U7639 (N_7639,N_3324,N_528);
and U7640 (N_7640,N_4587,N_2315);
nor U7641 (N_7641,N_3708,N_3259);
nand U7642 (N_7642,N_87,N_2931);
and U7643 (N_7643,N_1884,N_351);
nand U7644 (N_7644,N_236,N_1938);
nand U7645 (N_7645,N_2639,N_3988);
and U7646 (N_7646,N_3174,N_2715);
and U7647 (N_7647,N_2347,N_1078);
nand U7648 (N_7648,N_1437,N_1667);
nand U7649 (N_7649,N_1336,N_3866);
nor U7650 (N_7650,N_1238,N_2107);
or U7651 (N_7651,N_3918,N_4463);
nor U7652 (N_7652,N_3844,N_1633);
and U7653 (N_7653,N_1280,N_1651);
or U7654 (N_7654,N_1854,N_4723);
nand U7655 (N_7655,N_2331,N_4823);
or U7656 (N_7656,N_2534,N_39);
nand U7657 (N_7657,N_2024,N_1249);
nand U7658 (N_7658,N_579,N_586);
or U7659 (N_7659,N_1858,N_404);
and U7660 (N_7660,N_400,N_4881);
nand U7661 (N_7661,N_3780,N_2989);
or U7662 (N_7662,N_2668,N_3922);
and U7663 (N_7663,N_1789,N_4876);
nor U7664 (N_7664,N_988,N_4674);
and U7665 (N_7665,N_24,N_4510);
nand U7666 (N_7666,N_4195,N_2943);
or U7667 (N_7667,N_1691,N_4586);
or U7668 (N_7668,N_176,N_4425);
or U7669 (N_7669,N_2491,N_3926);
and U7670 (N_7670,N_788,N_2352);
and U7671 (N_7671,N_1602,N_1782);
or U7672 (N_7672,N_3562,N_4421);
nand U7673 (N_7673,N_157,N_4738);
or U7674 (N_7674,N_236,N_2177);
or U7675 (N_7675,N_2472,N_4981);
or U7676 (N_7676,N_761,N_3185);
and U7677 (N_7677,N_1811,N_4184);
or U7678 (N_7678,N_347,N_4526);
and U7679 (N_7679,N_2859,N_1406);
and U7680 (N_7680,N_321,N_1759);
nor U7681 (N_7681,N_4483,N_2779);
or U7682 (N_7682,N_4140,N_2413);
and U7683 (N_7683,N_1008,N_4825);
nor U7684 (N_7684,N_622,N_3594);
and U7685 (N_7685,N_4986,N_1748);
or U7686 (N_7686,N_2376,N_2473);
or U7687 (N_7687,N_4983,N_3926);
nand U7688 (N_7688,N_4029,N_3275);
nor U7689 (N_7689,N_3548,N_4911);
and U7690 (N_7690,N_1024,N_2078);
or U7691 (N_7691,N_3054,N_2005);
and U7692 (N_7692,N_3116,N_4438);
nor U7693 (N_7693,N_2982,N_948);
nand U7694 (N_7694,N_1766,N_4824);
and U7695 (N_7695,N_1687,N_990);
and U7696 (N_7696,N_621,N_3224);
nand U7697 (N_7697,N_3638,N_2173);
nor U7698 (N_7698,N_4008,N_264);
and U7699 (N_7699,N_2933,N_796);
and U7700 (N_7700,N_4702,N_3004);
nor U7701 (N_7701,N_4800,N_3045);
nor U7702 (N_7702,N_642,N_3539);
and U7703 (N_7703,N_2284,N_4970);
nor U7704 (N_7704,N_2061,N_4394);
or U7705 (N_7705,N_1477,N_4436);
nor U7706 (N_7706,N_4729,N_4173);
or U7707 (N_7707,N_1250,N_4652);
or U7708 (N_7708,N_1907,N_4268);
or U7709 (N_7709,N_3767,N_1555);
or U7710 (N_7710,N_4844,N_1877);
or U7711 (N_7711,N_1847,N_3021);
or U7712 (N_7712,N_2760,N_3278);
and U7713 (N_7713,N_3082,N_1100);
nor U7714 (N_7714,N_8,N_779);
nor U7715 (N_7715,N_1045,N_548);
nor U7716 (N_7716,N_4738,N_816);
and U7717 (N_7717,N_3594,N_4859);
or U7718 (N_7718,N_4077,N_4932);
nor U7719 (N_7719,N_3778,N_624);
nand U7720 (N_7720,N_3971,N_3870);
or U7721 (N_7721,N_1821,N_3991);
nor U7722 (N_7722,N_4932,N_4451);
nor U7723 (N_7723,N_187,N_1307);
and U7724 (N_7724,N_2163,N_4362);
and U7725 (N_7725,N_2173,N_4982);
nor U7726 (N_7726,N_150,N_3435);
and U7727 (N_7727,N_1366,N_4048);
and U7728 (N_7728,N_4544,N_3058);
or U7729 (N_7729,N_1154,N_2266);
xor U7730 (N_7730,N_2768,N_4215);
nor U7731 (N_7731,N_240,N_1479);
and U7732 (N_7732,N_1633,N_2343);
nand U7733 (N_7733,N_3918,N_1866);
nand U7734 (N_7734,N_683,N_2926);
or U7735 (N_7735,N_967,N_4257);
nand U7736 (N_7736,N_520,N_1113);
or U7737 (N_7737,N_4938,N_1379);
and U7738 (N_7738,N_1232,N_4941);
or U7739 (N_7739,N_279,N_4377);
and U7740 (N_7740,N_2291,N_4693);
and U7741 (N_7741,N_2128,N_3414);
and U7742 (N_7742,N_3208,N_3007);
nor U7743 (N_7743,N_770,N_2480);
nand U7744 (N_7744,N_4479,N_4221);
or U7745 (N_7745,N_2930,N_2693);
and U7746 (N_7746,N_1987,N_2314);
nand U7747 (N_7747,N_4818,N_234);
and U7748 (N_7748,N_2878,N_3758);
or U7749 (N_7749,N_4681,N_1297);
nor U7750 (N_7750,N_2493,N_2108);
and U7751 (N_7751,N_2086,N_2895);
and U7752 (N_7752,N_792,N_3605);
and U7753 (N_7753,N_1633,N_2039);
or U7754 (N_7754,N_341,N_2653);
and U7755 (N_7755,N_1521,N_2777);
nand U7756 (N_7756,N_145,N_1151);
nor U7757 (N_7757,N_613,N_2627);
or U7758 (N_7758,N_3126,N_304);
nor U7759 (N_7759,N_3398,N_1454);
nand U7760 (N_7760,N_184,N_2215);
and U7761 (N_7761,N_1839,N_4323);
nor U7762 (N_7762,N_3707,N_2693);
and U7763 (N_7763,N_4235,N_1934);
nand U7764 (N_7764,N_2993,N_3498);
and U7765 (N_7765,N_343,N_101);
or U7766 (N_7766,N_3508,N_2350);
and U7767 (N_7767,N_506,N_4428);
nor U7768 (N_7768,N_1862,N_4067);
or U7769 (N_7769,N_2422,N_736);
and U7770 (N_7770,N_1670,N_4864);
nor U7771 (N_7771,N_1103,N_4911);
and U7772 (N_7772,N_802,N_877);
nor U7773 (N_7773,N_3809,N_2419);
and U7774 (N_7774,N_4798,N_1141);
or U7775 (N_7775,N_4914,N_2060);
nand U7776 (N_7776,N_2949,N_3033);
nor U7777 (N_7777,N_3780,N_4648);
nand U7778 (N_7778,N_3899,N_3623);
or U7779 (N_7779,N_1525,N_2305);
and U7780 (N_7780,N_1701,N_839);
or U7781 (N_7781,N_2374,N_1165);
and U7782 (N_7782,N_705,N_1562);
and U7783 (N_7783,N_1124,N_4581);
nand U7784 (N_7784,N_4972,N_2168);
nor U7785 (N_7785,N_3118,N_406);
and U7786 (N_7786,N_3201,N_1980);
nor U7787 (N_7787,N_3843,N_4144);
and U7788 (N_7788,N_3824,N_1933);
and U7789 (N_7789,N_950,N_611);
and U7790 (N_7790,N_3612,N_428);
nand U7791 (N_7791,N_1597,N_963);
nor U7792 (N_7792,N_4669,N_3632);
and U7793 (N_7793,N_4008,N_592);
and U7794 (N_7794,N_632,N_1682);
or U7795 (N_7795,N_2919,N_4763);
and U7796 (N_7796,N_256,N_982);
and U7797 (N_7797,N_4122,N_3093);
or U7798 (N_7798,N_2962,N_2864);
and U7799 (N_7799,N_2299,N_682);
nor U7800 (N_7800,N_930,N_1159);
nand U7801 (N_7801,N_1052,N_1851);
nand U7802 (N_7802,N_710,N_1531);
and U7803 (N_7803,N_1511,N_848);
nand U7804 (N_7804,N_2458,N_1448);
or U7805 (N_7805,N_4188,N_1403);
xor U7806 (N_7806,N_128,N_1438);
nand U7807 (N_7807,N_4148,N_3992);
and U7808 (N_7808,N_1444,N_1924);
nand U7809 (N_7809,N_1116,N_2727);
nor U7810 (N_7810,N_3656,N_1383);
nand U7811 (N_7811,N_23,N_1226);
or U7812 (N_7812,N_4323,N_4755);
nand U7813 (N_7813,N_2451,N_2205);
nor U7814 (N_7814,N_4430,N_3954);
nor U7815 (N_7815,N_3058,N_4701);
xnor U7816 (N_7816,N_3426,N_2833);
nand U7817 (N_7817,N_1088,N_3834);
or U7818 (N_7818,N_343,N_4610);
and U7819 (N_7819,N_3781,N_4495);
nand U7820 (N_7820,N_2337,N_1989);
and U7821 (N_7821,N_771,N_2168);
or U7822 (N_7822,N_1431,N_1290);
or U7823 (N_7823,N_2628,N_1245);
or U7824 (N_7824,N_1222,N_4909);
nand U7825 (N_7825,N_1130,N_1059);
and U7826 (N_7826,N_464,N_2748);
nand U7827 (N_7827,N_3738,N_4671);
nor U7828 (N_7828,N_4163,N_4854);
and U7829 (N_7829,N_441,N_1651);
or U7830 (N_7830,N_811,N_1404);
or U7831 (N_7831,N_1381,N_2451);
nand U7832 (N_7832,N_2,N_1268);
and U7833 (N_7833,N_3565,N_327);
or U7834 (N_7834,N_1572,N_4344);
nor U7835 (N_7835,N_1245,N_1288);
nand U7836 (N_7836,N_2266,N_910);
nor U7837 (N_7837,N_146,N_179);
nand U7838 (N_7838,N_1733,N_2629);
nor U7839 (N_7839,N_3087,N_2005);
nor U7840 (N_7840,N_2472,N_4796);
nor U7841 (N_7841,N_78,N_3343);
and U7842 (N_7842,N_1366,N_3663);
and U7843 (N_7843,N_4143,N_2893);
and U7844 (N_7844,N_2868,N_940);
nand U7845 (N_7845,N_1062,N_1587);
nor U7846 (N_7846,N_2336,N_1924);
or U7847 (N_7847,N_789,N_4473);
or U7848 (N_7848,N_1579,N_2132);
and U7849 (N_7849,N_2666,N_3581);
nand U7850 (N_7850,N_1686,N_2044);
nor U7851 (N_7851,N_4079,N_2080);
or U7852 (N_7852,N_3091,N_910);
or U7853 (N_7853,N_1430,N_3815);
and U7854 (N_7854,N_1100,N_1489);
nor U7855 (N_7855,N_1736,N_3019);
and U7856 (N_7856,N_2010,N_752);
and U7857 (N_7857,N_3196,N_4803);
and U7858 (N_7858,N_4365,N_1232);
nand U7859 (N_7859,N_202,N_3593);
nor U7860 (N_7860,N_2455,N_2512);
nor U7861 (N_7861,N_2123,N_2134);
nor U7862 (N_7862,N_1865,N_2471);
or U7863 (N_7863,N_597,N_2697);
or U7864 (N_7864,N_165,N_2880);
or U7865 (N_7865,N_3474,N_4499);
nand U7866 (N_7866,N_190,N_2086);
nand U7867 (N_7867,N_3451,N_4605);
nand U7868 (N_7868,N_1784,N_169);
nand U7869 (N_7869,N_4992,N_717);
and U7870 (N_7870,N_982,N_1391);
nand U7871 (N_7871,N_2864,N_102);
nor U7872 (N_7872,N_181,N_4240);
nor U7873 (N_7873,N_1377,N_1107);
nand U7874 (N_7874,N_1107,N_4891);
and U7875 (N_7875,N_751,N_1518);
nor U7876 (N_7876,N_1833,N_2666);
nand U7877 (N_7877,N_1452,N_257);
nor U7878 (N_7878,N_4525,N_3299);
or U7879 (N_7879,N_1753,N_2851);
and U7880 (N_7880,N_1969,N_3550);
or U7881 (N_7881,N_17,N_2870);
nor U7882 (N_7882,N_413,N_3871);
nor U7883 (N_7883,N_4294,N_2128);
nor U7884 (N_7884,N_2643,N_1508);
nand U7885 (N_7885,N_2734,N_3464);
nand U7886 (N_7886,N_685,N_1639);
nor U7887 (N_7887,N_1991,N_3957);
and U7888 (N_7888,N_4316,N_783);
xnor U7889 (N_7889,N_334,N_927);
nor U7890 (N_7890,N_3019,N_1485);
nor U7891 (N_7891,N_2759,N_2032);
nand U7892 (N_7892,N_1507,N_2009);
and U7893 (N_7893,N_3689,N_3359);
nand U7894 (N_7894,N_4010,N_4608);
nand U7895 (N_7895,N_2376,N_4185);
nand U7896 (N_7896,N_2598,N_4999);
nor U7897 (N_7897,N_4445,N_3420);
and U7898 (N_7898,N_2863,N_429);
nor U7899 (N_7899,N_3605,N_2307);
nor U7900 (N_7900,N_513,N_4893);
and U7901 (N_7901,N_612,N_937);
and U7902 (N_7902,N_1807,N_409);
xnor U7903 (N_7903,N_1338,N_3896);
or U7904 (N_7904,N_3848,N_4623);
and U7905 (N_7905,N_3936,N_2068);
nor U7906 (N_7906,N_4235,N_50);
or U7907 (N_7907,N_1965,N_2560);
nand U7908 (N_7908,N_2179,N_4253);
and U7909 (N_7909,N_2127,N_3696);
or U7910 (N_7910,N_3,N_1906);
and U7911 (N_7911,N_949,N_3937);
and U7912 (N_7912,N_2488,N_95);
nor U7913 (N_7913,N_1833,N_805);
nor U7914 (N_7914,N_4095,N_1235);
or U7915 (N_7915,N_3113,N_2588);
or U7916 (N_7916,N_448,N_3943);
nor U7917 (N_7917,N_2974,N_4337);
or U7918 (N_7918,N_3927,N_3126);
or U7919 (N_7919,N_2006,N_4540);
nor U7920 (N_7920,N_726,N_801);
and U7921 (N_7921,N_700,N_3412);
or U7922 (N_7922,N_1879,N_1898);
nand U7923 (N_7923,N_4520,N_4208);
nor U7924 (N_7924,N_4396,N_2048);
nor U7925 (N_7925,N_3317,N_4265);
nor U7926 (N_7926,N_3095,N_385);
nand U7927 (N_7927,N_1904,N_306);
nand U7928 (N_7928,N_1493,N_1418);
nand U7929 (N_7929,N_1254,N_4265);
xor U7930 (N_7930,N_641,N_2505);
nand U7931 (N_7931,N_3770,N_3691);
nor U7932 (N_7932,N_223,N_4906);
nand U7933 (N_7933,N_687,N_761);
and U7934 (N_7934,N_4925,N_4306);
or U7935 (N_7935,N_2441,N_2214);
or U7936 (N_7936,N_1403,N_2281);
or U7937 (N_7937,N_3272,N_3584);
nor U7938 (N_7938,N_3267,N_283);
and U7939 (N_7939,N_2340,N_2618);
and U7940 (N_7940,N_666,N_4101);
nor U7941 (N_7941,N_2624,N_1801);
nor U7942 (N_7942,N_3805,N_2915);
nor U7943 (N_7943,N_3970,N_1403);
nand U7944 (N_7944,N_2062,N_2533);
and U7945 (N_7945,N_933,N_16);
nand U7946 (N_7946,N_1275,N_2329);
or U7947 (N_7947,N_1334,N_4405);
or U7948 (N_7948,N_2428,N_925);
xor U7949 (N_7949,N_4851,N_399);
nor U7950 (N_7950,N_1688,N_57);
nand U7951 (N_7951,N_428,N_2096);
or U7952 (N_7952,N_3314,N_49);
and U7953 (N_7953,N_3623,N_3036);
nand U7954 (N_7954,N_4103,N_4166);
nand U7955 (N_7955,N_2099,N_3141);
and U7956 (N_7956,N_3899,N_761);
nor U7957 (N_7957,N_1151,N_4455);
nor U7958 (N_7958,N_4562,N_3306);
nand U7959 (N_7959,N_4224,N_1215);
and U7960 (N_7960,N_1982,N_1000);
or U7961 (N_7961,N_3695,N_1905);
or U7962 (N_7962,N_556,N_939);
nor U7963 (N_7963,N_992,N_1136);
nor U7964 (N_7964,N_911,N_1231);
nor U7965 (N_7965,N_4762,N_4213);
and U7966 (N_7966,N_618,N_1943);
or U7967 (N_7967,N_1003,N_2682);
and U7968 (N_7968,N_271,N_400);
and U7969 (N_7969,N_2836,N_3032);
and U7970 (N_7970,N_3387,N_4841);
nor U7971 (N_7971,N_532,N_1622);
nor U7972 (N_7972,N_1795,N_1574);
and U7973 (N_7973,N_2154,N_4380);
nor U7974 (N_7974,N_2642,N_774);
or U7975 (N_7975,N_140,N_4012);
and U7976 (N_7976,N_4090,N_3627);
and U7977 (N_7977,N_310,N_1164);
nor U7978 (N_7978,N_4371,N_3932);
nand U7979 (N_7979,N_2775,N_1301);
or U7980 (N_7980,N_1933,N_1454);
or U7981 (N_7981,N_3963,N_4304);
or U7982 (N_7982,N_785,N_2992);
and U7983 (N_7983,N_251,N_2784);
or U7984 (N_7984,N_3347,N_1192);
nand U7985 (N_7985,N_2971,N_2752);
nand U7986 (N_7986,N_51,N_3143);
and U7987 (N_7987,N_1475,N_746);
or U7988 (N_7988,N_1761,N_1751);
and U7989 (N_7989,N_814,N_4732);
nor U7990 (N_7990,N_1141,N_2584);
or U7991 (N_7991,N_477,N_640);
and U7992 (N_7992,N_4465,N_3114);
or U7993 (N_7993,N_1480,N_800);
nand U7994 (N_7994,N_3158,N_4917);
and U7995 (N_7995,N_2578,N_4250);
or U7996 (N_7996,N_922,N_3474);
and U7997 (N_7997,N_2193,N_2549);
and U7998 (N_7998,N_3367,N_4989);
and U7999 (N_7999,N_3490,N_3161);
nand U8000 (N_8000,N_3572,N_2485);
nor U8001 (N_8001,N_4756,N_937);
nor U8002 (N_8002,N_2252,N_4686);
nor U8003 (N_8003,N_1830,N_3041);
nor U8004 (N_8004,N_1384,N_3888);
nor U8005 (N_8005,N_1410,N_812);
or U8006 (N_8006,N_82,N_4563);
or U8007 (N_8007,N_2524,N_3026);
nor U8008 (N_8008,N_3386,N_4586);
nor U8009 (N_8009,N_3372,N_2655);
and U8010 (N_8010,N_4713,N_302);
or U8011 (N_8011,N_2538,N_4752);
nand U8012 (N_8012,N_792,N_2492);
nor U8013 (N_8013,N_3423,N_932);
or U8014 (N_8014,N_1239,N_2681);
nor U8015 (N_8015,N_1349,N_1195);
nor U8016 (N_8016,N_457,N_1759);
nor U8017 (N_8017,N_4167,N_404);
nor U8018 (N_8018,N_4589,N_2806);
and U8019 (N_8019,N_1572,N_3091);
or U8020 (N_8020,N_435,N_1595);
or U8021 (N_8021,N_1201,N_2612);
and U8022 (N_8022,N_706,N_3177);
nand U8023 (N_8023,N_1142,N_553);
nand U8024 (N_8024,N_4521,N_538);
and U8025 (N_8025,N_1214,N_973);
nor U8026 (N_8026,N_4093,N_1094);
nand U8027 (N_8027,N_2019,N_759);
and U8028 (N_8028,N_4906,N_187);
and U8029 (N_8029,N_2233,N_1318);
nand U8030 (N_8030,N_1222,N_4599);
nand U8031 (N_8031,N_4596,N_480);
nand U8032 (N_8032,N_2893,N_1918);
nor U8033 (N_8033,N_4505,N_3275);
nor U8034 (N_8034,N_1476,N_905);
nand U8035 (N_8035,N_2021,N_2694);
nor U8036 (N_8036,N_185,N_3387);
xor U8037 (N_8037,N_3518,N_1500);
nand U8038 (N_8038,N_885,N_53);
nor U8039 (N_8039,N_2669,N_935);
and U8040 (N_8040,N_2670,N_1570);
nand U8041 (N_8041,N_2773,N_3365);
nor U8042 (N_8042,N_3660,N_281);
or U8043 (N_8043,N_2201,N_3657);
and U8044 (N_8044,N_3807,N_3129);
nor U8045 (N_8045,N_1908,N_4351);
nor U8046 (N_8046,N_2725,N_1168);
and U8047 (N_8047,N_106,N_1836);
and U8048 (N_8048,N_3108,N_4038);
xnor U8049 (N_8049,N_1587,N_681);
and U8050 (N_8050,N_3862,N_1867);
or U8051 (N_8051,N_2083,N_4549);
or U8052 (N_8052,N_268,N_4460);
or U8053 (N_8053,N_1228,N_4470);
nand U8054 (N_8054,N_3190,N_4209);
nor U8055 (N_8055,N_2418,N_4056);
or U8056 (N_8056,N_1898,N_334);
nor U8057 (N_8057,N_3598,N_3476);
nor U8058 (N_8058,N_3494,N_2355);
nand U8059 (N_8059,N_2511,N_348);
nor U8060 (N_8060,N_3295,N_2544);
and U8061 (N_8061,N_1101,N_4576);
and U8062 (N_8062,N_3727,N_1707);
and U8063 (N_8063,N_4110,N_4596);
and U8064 (N_8064,N_2760,N_2527);
nor U8065 (N_8065,N_710,N_4459);
nor U8066 (N_8066,N_4320,N_2020);
or U8067 (N_8067,N_4788,N_2116);
and U8068 (N_8068,N_3402,N_609);
and U8069 (N_8069,N_1109,N_1487);
and U8070 (N_8070,N_1832,N_26);
nand U8071 (N_8071,N_148,N_1089);
and U8072 (N_8072,N_2689,N_4963);
nor U8073 (N_8073,N_90,N_3944);
or U8074 (N_8074,N_2596,N_1273);
and U8075 (N_8075,N_892,N_1526);
and U8076 (N_8076,N_2947,N_3542);
nor U8077 (N_8077,N_4413,N_1559);
nor U8078 (N_8078,N_2188,N_1839);
and U8079 (N_8079,N_4487,N_1094);
nor U8080 (N_8080,N_2293,N_2953);
nand U8081 (N_8081,N_321,N_4227);
nand U8082 (N_8082,N_2139,N_1644);
nand U8083 (N_8083,N_2900,N_4544);
nand U8084 (N_8084,N_688,N_3723);
nor U8085 (N_8085,N_3567,N_137);
and U8086 (N_8086,N_4684,N_681);
nand U8087 (N_8087,N_4576,N_1190);
nor U8088 (N_8088,N_2527,N_962);
nand U8089 (N_8089,N_3008,N_3429);
and U8090 (N_8090,N_1044,N_4504);
nor U8091 (N_8091,N_4317,N_1815);
and U8092 (N_8092,N_2146,N_3902);
or U8093 (N_8093,N_3833,N_1927);
and U8094 (N_8094,N_1813,N_1940);
and U8095 (N_8095,N_377,N_1032);
and U8096 (N_8096,N_1976,N_603);
and U8097 (N_8097,N_3514,N_1464);
nor U8098 (N_8098,N_722,N_3893);
nand U8099 (N_8099,N_2551,N_1249);
or U8100 (N_8100,N_2794,N_2842);
nor U8101 (N_8101,N_748,N_1933);
nand U8102 (N_8102,N_3108,N_1423);
nor U8103 (N_8103,N_4614,N_4887);
or U8104 (N_8104,N_1843,N_1645);
nand U8105 (N_8105,N_636,N_4208);
or U8106 (N_8106,N_1459,N_2000);
and U8107 (N_8107,N_3990,N_1071);
nor U8108 (N_8108,N_1067,N_2040);
and U8109 (N_8109,N_3501,N_2522);
or U8110 (N_8110,N_3981,N_825);
nand U8111 (N_8111,N_3291,N_4220);
or U8112 (N_8112,N_2957,N_4067);
and U8113 (N_8113,N_4256,N_451);
nor U8114 (N_8114,N_561,N_420);
and U8115 (N_8115,N_469,N_501);
or U8116 (N_8116,N_2440,N_4073);
xor U8117 (N_8117,N_4800,N_4207);
nand U8118 (N_8118,N_1126,N_2413);
nor U8119 (N_8119,N_2561,N_4415);
or U8120 (N_8120,N_1062,N_2245);
nor U8121 (N_8121,N_3365,N_1360);
nor U8122 (N_8122,N_635,N_4595);
nor U8123 (N_8123,N_1772,N_1852);
or U8124 (N_8124,N_4361,N_3152);
nor U8125 (N_8125,N_1776,N_126);
nand U8126 (N_8126,N_4033,N_1463);
nand U8127 (N_8127,N_4651,N_552);
or U8128 (N_8128,N_2998,N_408);
or U8129 (N_8129,N_1498,N_890);
nor U8130 (N_8130,N_2931,N_3764);
nor U8131 (N_8131,N_4325,N_2107);
nand U8132 (N_8132,N_2956,N_4096);
nand U8133 (N_8133,N_317,N_876);
nor U8134 (N_8134,N_4356,N_2306);
or U8135 (N_8135,N_3397,N_2495);
nor U8136 (N_8136,N_1069,N_1175);
or U8137 (N_8137,N_4215,N_1052);
and U8138 (N_8138,N_3936,N_2096);
nor U8139 (N_8139,N_3082,N_501);
nor U8140 (N_8140,N_3298,N_1611);
and U8141 (N_8141,N_1058,N_993);
nor U8142 (N_8142,N_54,N_1519);
and U8143 (N_8143,N_2573,N_4234);
or U8144 (N_8144,N_711,N_3788);
or U8145 (N_8145,N_115,N_4635);
nand U8146 (N_8146,N_2112,N_2185);
and U8147 (N_8147,N_1549,N_4762);
nand U8148 (N_8148,N_4813,N_182);
or U8149 (N_8149,N_3274,N_311);
xor U8150 (N_8150,N_2775,N_4139);
and U8151 (N_8151,N_3127,N_267);
and U8152 (N_8152,N_339,N_1647);
or U8153 (N_8153,N_4197,N_3274);
nand U8154 (N_8154,N_3072,N_3970);
nor U8155 (N_8155,N_189,N_658);
and U8156 (N_8156,N_2911,N_3292);
nand U8157 (N_8157,N_4742,N_1649);
nand U8158 (N_8158,N_3182,N_2225);
and U8159 (N_8159,N_954,N_1466);
nor U8160 (N_8160,N_4774,N_4614);
nor U8161 (N_8161,N_2600,N_921);
xnor U8162 (N_8162,N_4623,N_1723);
nand U8163 (N_8163,N_412,N_2668);
nand U8164 (N_8164,N_3940,N_2230);
and U8165 (N_8165,N_1643,N_3108);
or U8166 (N_8166,N_1250,N_3655);
and U8167 (N_8167,N_765,N_957);
nor U8168 (N_8168,N_2336,N_3769);
nor U8169 (N_8169,N_3435,N_3922);
or U8170 (N_8170,N_1055,N_460);
and U8171 (N_8171,N_2992,N_2596);
nor U8172 (N_8172,N_526,N_2876);
and U8173 (N_8173,N_3302,N_2482);
nor U8174 (N_8174,N_1010,N_161);
and U8175 (N_8175,N_3827,N_3442);
nand U8176 (N_8176,N_2947,N_595);
nor U8177 (N_8177,N_21,N_4131);
nand U8178 (N_8178,N_2974,N_4960);
or U8179 (N_8179,N_2360,N_3648);
nor U8180 (N_8180,N_2006,N_2749);
and U8181 (N_8181,N_1362,N_1745);
nand U8182 (N_8182,N_1599,N_3539);
nand U8183 (N_8183,N_107,N_4456);
nand U8184 (N_8184,N_4568,N_3565);
nand U8185 (N_8185,N_4718,N_108);
nand U8186 (N_8186,N_3492,N_1793);
and U8187 (N_8187,N_869,N_1576);
or U8188 (N_8188,N_1313,N_4870);
nor U8189 (N_8189,N_4602,N_4324);
and U8190 (N_8190,N_265,N_3398);
nand U8191 (N_8191,N_4817,N_113);
nor U8192 (N_8192,N_4320,N_3397);
or U8193 (N_8193,N_1434,N_3895);
and U8194 (N_8194,N_3955,N_1307);
nand U8195 (N_8195,N_1350,N_3684);
and U8196 (N_8196,N_3076,N_345);
nand U8197 (N_8197,N_2502,N_981);
and U8198 (N_8198,N_1231,N_3856);
and U8199 (N_8199,N_1314,N_3124);
nand U8200 (N_8200,N_4606,N_572);
nor U8201 (N_8201,N_3808,N_2615);
and U8202 (N_8202,N_1437,N_2773);
nor U8203 (N_8203,N_2669,N_3313);
xnor U8204 (N_8204,N_0,N_3867);
nand U8205 (N_8205,N_283,N_646);
xnor U8206 (N_8206,N_238,N_2906);
nand U8207 (N_8207,N_890,N_4440);
nand U8208 (N_8208,N_2645,N_3690);
nor U8209 (N_8209,N_948,N_4595);
and U8210 (N_8210,N_1042,N_983);
and U8211 (N_8211,N_1145,N_4299);
nand U8212 (N_8212,N_1981,N_3209);
or U8213 (N_8213,N_598,N_1813);
xnor U8214 (N_8214,N_267,N_4289);
nor U8215 (N_8215,N_4369,N_4801);
or U8216 (N_8216,N_397,N_2967);
and U8217 (N_8217,N_413,N_4879);
nor U8218 (N_8218,N_1326,N_2878);
or U8219 (N_8219,N_2271,N_4757);
and U8220 (N_8220,N_3253,N_616);
nand U8221 (N_8221,N_1424,N_2944);
and U8222 (N_8222,N_759,N_2989);
or U8223 (N_8223,N_3213,N_2451);
and U8224 (N_8224,N_1027,N_409);
nor U8225 (N_8225,N_775,N_2712);
or U8226 (N_8226,N_3046,N_3431);
nand U8227 (N_8227,N_946,N_2000);
or U8228 (N_8228,N_3885,N_2556);
nand U8229 (N_8229,N_4947,N_4453);
or U8230 (N_8230,N_394,N_3141);
nor U8231 (N_8231,N_1966,N_1497);
nand U8232 (N_8232,N_3275,N_2537);
or U8233 (N_8233,N_3496,N_1388);
nor U8234 (N_8234,N_4438,N_60);
or U8235 (N_8235,N_2426,N_3210);
and U8236 (N_8236,N_1527,N_891);
nand U8237 (N_8237,N_4855,N_2127);
nand U8238 (N_8238,N_3622,N_1221);
nand U8239 (N_8239,N_4951,N_4193);
nand U8240 (N_8240,N_2434,N_2521);
nand U8241 (N_8241,N_1710,N_2101);
or U8242 (N_8242,N_1252,N_3789);
and U8243 (N_8243,N_1383,N_3951);
nand U8244 (N_8244,N_242,N_3276);
or U8245 (N_8245,N_610,N_2671);
or U8246 (N_8246,N_4772,N_2851);
and U8247 (N_8247,N_2514,N_4806);
or U8248 (N_8248,N_4773,N_2936);
nand U8249 (N_8249,N_4036,N_1783);
nand U8250 (N_8250,N_112,N_921);
nor U8251 (N_8251,N_2197,N_1924);
or U8252 (N_8252,N_4778,N_4652);
and U8253 (N_8253,N_1533,N_1961);
and U8254 (N_8254,N_3951,N_4609);
nor U8255 (N_8255,N_3509,N_3495);
or U8256 (N_8256,N_4386,N_4538);
and U8257 (N_8257,N_2411,N_2758);
or U8258 (N_8258,N_302,N_1928);
nand U8259 (N_8259,N_4190,N_614);
or U8260 (N_8260,N_207,N_3076);
nor U8261 (N_8261,N_4930,N_2905);
or U8262 (N_8262,N_1840,N_3271);
or U8263 (N_8263,N_3039,N_1400);
or U8264 (N_8264,N_1723,N_1777);
nor U8265 (N_8265,N_217,N_1148);
or U8266 (N_8266,N_1104,N_2611);
and U8267 (N_8267,N_3369,N_397);
and U8268 (N_8268,N_4010,N_3729);
nor U8269 (N_8269,N_315,N_4276);
or U8270 (N_8270,N_4767,N_1447);
and U8271 (N_8271,N_569,N_4341);
or U8272 (N_8272,N_73,N_1162);
nand U8273 (N_8273,N_2948,N_4609);
nand U8274 (N_8274,N_2045,N_451);
nor U8275 (N_8275,N_4070,N_1717);
nor U8276 (N_8276,N_4797,N_3176);
nand U8277 (N_8277,N_3918,N_2614);
and U8278 (N_8278,N_3000,N_2919);
nor U8279 (N_8279,N_3078,N_216);
and U8280 (N_8280,N_2587,N_2187);
and U8281 (N_8281,N_3769,N_3757);
nand U8282 (N_8282,N_2009,N_3475);
nor U8283 (N_8283,N_2194,N_359);
nand U8284 (N_8284,N_3606,N_2436);
or U8285 (N_8285,N_3242,N_265);
and U8286 (N_8286,N_1109,N_2978);
or U8287 (N_8287,N_1658,N_1974);
nor U8288 (N_8288,N_149,N_3867);
or U8289 (N_8289,N_3963,N_1682);
nor U8290 (N_8290,N_4170,N_1009);
nand U8291 (N_8291,N_856,N_4119);
and U8292 (N_8292,N_4421,N_1188);
and U8293 (N_8293,N_1404,N_2512);
nor U8294 (N_8294,N_4799,N_1747);
nor U8295 (N_8295,N_2281,N_3301);
and U8296 (N_8296,N_322,N_1071);
nor U8297 (N_8297,N_4700,N_707);
or U8298 (N_8298,N_4827,N_283);
nand U8299 (N_8299,N_2630,N_3112);
nand U8300 (N_8300,N_314,N_4344);
xnor U8301 (N_8301,N_4862,N_1233);
nor U8302 (N_8302,N_3378,N_3323);
nand U8303 (N_8303,N_5,N_1693);
or U8304 (N_8304,N_2958,N_1348);
nand U8305 (N_8305,N_383,N_1344);
xnor U8306 (N_8306,N_24,N_527);
nor U8307 (N_8307,N_2505,N_1965);
nor U8308 (N_8308,N_682,N_889);
or U8309 (N_8309,N_3787,N_4132);
nand U8310 (N_8310,N_660,N_797);
and U8311 (N_8311,N_4043,N_691);
and U8312 (N_8312,N_722,N_1792);
nor U8313 (N_8313,N_4142,N_4605);
and U8314 (N_8314,N_3026,N_4755);
and U8315 (N_8315,N_3116,N_4705);
and U8316 (N_8316,N_1297,N_4261);
nor U8317 (N_8317,N_868,N_332);
nand U8318 (N_8318,N_2027,N_4103);
or U8319 (N_8319,N_1962,N_3045);
nand U8320 (N_8320,N_1735,N_3914);
nand U8321 (N_8321,N_659,N_2096);
and U8322 (N_8322,N_1594,N_1024);
nor U8323 (N_8323,N_3998,N_2757);
and U8324 (N_8324,N_3179,N_3162);
and U8325 (N_8325,N_364,N_1405);
or U8326 (N_8326,N_4720,N_820);
nor U8327 (N_8327,N_2226,N_2359);
nor U8328 (N_8328,N_4939,N_4143);
and U8329 (N_8329,N_2163,N_3295);
nor U8330 (N_8330,N_3984,N_2175);
nand U8331 (N_8331,N_194,N_2034);
nor U8332 (N_8332,N_2200,N_3117);
and U8333 (N_8333,N_557,N_4385);
or U8334 (N_8334,N_209,N_1932);
nor U8335 (N_8335,N_3160,N_1427);
nor U8336 (N_8336,N_4103,N_4503);
nand U8337 (N_8337,N_2380,N_780);
nand U8338 (N_8338,N_4699,N_4065);
nand U8339 (N_8339,N_1249,N_1316);
nand U8340 (N_8340,N_99,N_2939);
and U8341 (N_8341,N_4405,N_3647);
and U8342 (N_8342,N_1021,N_2155);
nand U8343 (N_8343,N_1023,N_501);
nand U8344 (N_8344,N_309,N_2704);
nor U8345 (N_8345,N_1865,N_608);
nor U8346 (N_8346,N_1105,N_1480);
or U8347 (N_8347,N_2060,N_3387);
or U8348 (N_8348,N_3668,N_936);
or U8349 (N_8349,N_1610,N_760);
and U8350 (N_8350,N_2486,N_2071);
or U8351 (N_8351,N_2741,N_4557);
and U8352 (N_8352,N_2199,N_3371);
nor U8353 (N_8353,N_344,N_1391);
nand U8354 (N_8354,N_4105,N_1803);
and U8355 (N_8355,N_254,N_2227);
and U8356 (N_8356,N_1506,N_3942);
nor U8357 (N_8357,N_3439,N_4009);
or U8358 (N_8358,N_1289,N_4777);
nand U8359 (N_8359,N_4673,N_4137);
nand U8360 (N_8360,N_67,N_2226);
nand U8361 (N_8361,N_1787,N_4851);
or U8362 (N_8362,N_3766,N_26);
and U8363 (N_8363,N_962,N_3737);
and U8364 (N_8364,N_65,N_474);
nor U8365 (N_8365,N_1509,N_1988);
or U8366 (N_8366,N_2898,N_3118);
nand U8367 (N_8367,N_807,N_4853);
nand U8368 (N_8368,N_4903,N_3503);
nand U8369 (N_8369,N_1493,N_4613);
and U8370 (N_8370,N_1289,N_551);
and U8371 (N_8371,N_1023,N_2863);
and U8372 (N_8372,N_325,N_861);
nor U8373 (N_8373,N_4801,N_2715);
nor U8374 (N_8374,N_2755,N_4117);
nor U8375 (N_8375,N_2481,N_3009);
nor U8376 (N_8376,N_317,N_2444);
or U8377 (N_8377,N_1939,N_406);
nor U8378 (N_8378,N_2136,N_3084);
or U8379 (N_8379,N_2612,N_2590);
nor U8380 (N_8380,N_2301,N_4136);
and U8381 (N_8381,N_2933,N_3784);
nand U8382 (N_8382,N_4937,N_3247);
and U8383 (N_8383,N_2182,N_1745);
nand U8384 (N_8384,N_1392,N_563);
nor U8385 (N_8385,N_1398,N_1489);
nand U8386 (N_8386,N_1155,N_3908);
or U8387 (N_8387,N_3020,N_1933);
nand U8388 (N_8388,N_708,N_583);
nand U8389 (N_8389,N_2176,N_4313);
and U8390 (N_8390,N_1825,N_3720);
nor U8391 (N_8391,N_3281,N_707);
and U8392 (N_8392,N_1068,N_391);
nand U8393 (N_8393,N_245,N_1887);
or U8394 (N_8394,N_4463,N_3128);
and U8395 (N_8395,N_1926,N_4978);
nor U8396 (N_8396,N_2639,N_2535);
nor U8397 (N_8397,N_1677,N_1892);
nor U8398 (N_8398,N_2935,N_210);
nand U8399 (N_8399,N_1278,N_1334);
nor U8400 (N_8400,N_4931,N_4099);
nand U8401 (N_8401,N_4512,N_4267);
nor U8402 (N_8402,N_3410,N_3659);
or U8403 (N_8403,N_2646,N_3192);
nand U8404 (N_8404,N_2363,N_2588);
and U8405 (N_8405,N_271,N_2990);
and U8406 (N_8406,N_1245,N_4991);
xnor U8407 (N_8407,N_4573,N_235);
and U8408 (N_8408,N_2563,N_3201);
nor U8409 (N_8409,N_1268,N_1574);
and U8410 (N_8410,N_545,N_4725);
nand U8411 (N_8411,N_4845,N_3403);
and U8412 (N_8412,N_2092,N_1553);
or U8413 (N_8413,N_1863,N_1703);
nand U8414 (N_8414,N_2410,N_1005);
nand U8415 (N_8415,N_1129,N_3308);
nand U8416 (N_8416,N_468,N_4741);
or U8417 (N_8417,N_2336,N_4341);
nand U8418 (N_8418,N_1446,N_2591);
and U8419 (N_8419,N_4161,N_669);
nor U8420 (N_8420,N_352,N_2008);
nor U8421 (N_8421,N_1798,N_2062);
nand U8422 (N_8422,N_415,N_3880);
or U8423 (N_8423,N_1664,N_1755);
nand U8424 (N_8424,N_2166,N_2153);
nand U8425 (N_8425,N_1909,N_2576);
or U8426 (N_8426,N_4393,N_3098);
and U8427 (N_8427,N_2057,N_479);
nand U8428 (N_8428,N_3367,N_1944);
or U8429 (N_8429,N_916,N_4788);
nand U8430 (N_8430,N_1828,N_4414);
nor U8431 (N_8431,N_1509,N_341);
nor U8432 (N_8432,N_2037,N_3591);
or U8433 (N_8433,N_4210,N_4691);
nor U8434 (N_8434,N_3179,N_4626);
and U8435 (N_8435,N_2396,N_954);
nand U8436 (N_8436,N_4301,N_1528);
nand U8437 (N_8437,N_2480,N_430);
nand U8438 (N_8438,N_551,N_4758);
nand U8439 (N_8439,N_4799,N_3845);
or U8440 (N_8440,N_4888,N_3596);
nor U8441 (N_8441,N_2722,N_2973);
nand U8442 (N_8442,N_3809,N_1535);
nand U8443 (N_8443,N_3052,N_2424);
and U8444 (N_8444,N_4620,N_4228);
and U8445 (N_8445,N_2751,N_1249);
or U8446 (N_8446,N_2850,N_4630);
or U8447 (N_8447,N_4145,N_2170);
nor U8448 (N_8448,N_3553,N_282);
nor U8449 (N_8449,N_1128,N_1221);
or U8450 (N_8450,N_1335,N_4999);
nand U8451 (N_8451,N_510,N_1843);
nor U8452 (N_8452,N_4493,N_1087);
nor U8453 (N_8453,N_3338,N_983);
nor U8454 (N_8454,N_4989,N_3349);
or U8455 (N_8455,N_3015,N_4765);
and U8456 (N_8456,N_1042,N_4102);
or U8457 (N_8457,N_2830,N_4026);
and U8458 (N_8458,N_501,N_1861);
nand U8459 (N_8459,N_2322,N_2439);
nor U8460 (N_8460,N_3209,N_2568);
or U8461 (N_8461,N_442,N_3314);
or U8462 (N_8462,N_1516,N_3222);
or U8463 (N_8463,N_1918,N_3609);
nor U8464 (N_8464,N_4419,N_3971);
nor U8465 (N_8465,N_3956,N_2136);
or U8466 (N_8466,N_1833,N_1967);
nand U8467 (N_8467,N_2412,N_1773);
or U8468 (N_8468,N_3953,N_3455);
nand U8469 (N_8469,N_3584,N_1587);
nand U8470 (N_8470,N_107,N_2675);
nor U8471 (N_8471,N_97,N_1598);
nand U8472 (N_8472,N_4200,N_90);
nand U8473 (N_8473,N_759,N_2205);
or U8474 (N_8474,N_2297,N_3968);
and U8475 (N_8475,N_4938,N_3876);
nor U8476 (N_8476,N_2940,N_4095);
nor U8477 (N_8477,N_56,N_4393);
nor U8478 (N_8478,N_1490,N_1990);
nand U8479 (N_8479,N_2496,N_4150);
and U8480 (N_8480,N_1574,N_4377);
and U8481 (N_8481,N_3807,N_4351);
nand U8482 (N_8482,N_2542,N_4042);
and U8483 (N_8483,N_2458,N_4272);
and U8484 (N_8484,N_3445,N_3187);
or U8485 (N_8485,N_119,N_2560);
and U8486 (N_8486,N_3307,N_385);
nand U8487 (N_8487,N_3075,N_1435);
nand U8488 (N_8488,N_2247,N_3717);
and U8489 (N_8489,N_3164,N_4332);
nand U8490 (N_8490,N_4495,N_2720);
nand U8491 (N_8491,N_1261,N_210);
nand U8492 (N_8492,N_400,N_721);
or U8493 (N_8493,N_4412,N_1431);
nand U8494 (N_8494,N_4713,N_3597);
nand U8495 (N_8495,N_4466,N_2751);
nor U8496 (N_8496,N_4847,N_1271);
or U8497 (N_8497,N_598,N_1048);
or U8498 (N_8498,N_4929,N_4126);
and U8499 (N_8499,N_1748,N_185);
or U8500 (N_8500,N_3815,N_955);
nor U8501 (N_8501,N_807,N_120);
nand U8502 (N_8502,N_4460,N_2977);
nor U8503 (N_8503,N_19,N_3762);
nand U8504 (N_8504,N_1978,N_4573);
nand U8505 (N_8505,N_3903,N_3415);
or U8506 (N_8506,N_4924,N_2673);
nand U8507 (N_8507,N_855,N_4748);
or U8508 (N_8508,N_4601,N_2044);
and U8509 (N_8509,N_2144,N_2041);
nand U8510 (N_8510,N_692,N_4475);
nand U8511 (N_8511,N_327,N_2550);
nor U8512 (N_8512,N_2454,N_4743);
nor U8513 (N_8513,N_3310,N_2303);
nor U8514 (N_8514,N_2072,N_1415);
nor U8515 (N_8515,N_4647,N_900);
nand U8516 (N_8516,N_697,N_1769);
and U8517 (N_8517,N_1594,N_4134);
or U8518 (N_8518,N_139,N_1397);
or U8519 (N_8519,N_3318,N_1882);
nor U8520 (N_8520,N_1925,N_3002);
nor U8521 (N_8521,N_4009,N_4528);
nor U8522 (N_8522,N_1361,N_592);
nand U8523 (N_8523,N_2080,N_2738);
or U8524 (N_8524,N_4908,N_647);
or U8525 (N_8525,N_3373,N_4715);
and U8526 (N_8526,N_278,N_951);
nor U8527 (N_8527,N_1522,N_3009);
nor U8528 (N_8528,N_363,N_3337);
or U8529 (N_8529,N_3156,N_3199);
nand U8530 (N_8530,N_77,N_3334);
nand U8531 (N_8531,N_4991,N_957);
nor U8532 (N_8532,N_767,N_4102);
and U8533 (N_8533,N_53,N_2646);
nand U8534 (N_8534,N_358,N_1916);
and U8535 (N_8535,N_3930,N_1182);
or U8536 (N_8536,N_1655,N_2179);
nor U8537 (N_8537,N_178,N_4760);
or U8538 (N_8538,N_3459,N_2966);
nor U8539 (N_8539,N_2681,N_923);
nand U8540 (N_8540,N_1007,N_70);
nor U8541 (N_8541,N_1473,N_1327);
and U8542 (N_8542,N_3405,N_2685);
or U8543 (N_8543,N_723,N_3564);
or U8544 (N_8544,N_457,N_844);
or U8545 (N_8545,N_4848,N_1283);
and U8546 (N_8546,N_1897,N_638);
xnor U8547 (N_8547,N_2133,N_4635);
nor U8548 (N_8548,N_263,N_4706);
or U8549 (N_8549,N_2258,N_1164);
or U8550 (N_8550,N_2446,N_3965);
and U8551 (N_8551,N_4407,N_4205);
and U8552 (N_8552,N_4207,N_2577);
and U8553 (N_8553,N_3257,N_719);
and U8554 (N_8554,N_4629,N_1463);
nor U8555 (N_8555,N_3411,N_2482);
nand U8556 (N_8556,N_1449,N_2054);
nor U8557 (N_8557,N_4094,N_2051);
and U8558 (N_8558,N_4356,N_3125);
and U8559 (N_8559,N_74,N_1508);
and U8560 (N_8560,N_2114,N_1315);
nand U8561 (N_8561,N_4241,N_1915);
nand U8562 (N_8562,N_1448,N_2443);
nor U8563 (N_8563,N_4608,N_2779);
and U8564 (N_8564,N_4021,N_3463);
nand U8565 (N_8565,N_4903,N_3095);
nand U8566 (N_8566,N_1338,N_4318);
nor U8567 (N_8567,N_54,N_3018);
and U8568 (N_8568,N_4583,N_2084);
or U8569 (N_8569,N_2114,N_1400);
xnor U8570 (N_8570,N_1516,N_4138);
nor U8571 (N_8571,N_3684,N_1589);
nand U8572 (N_8572,N_63,N_4001);
and U8573 (N_8573,N_4853,N_148);
and U8574 (N_8574,N_1133,N_3506);
and U8575 (N_8575,N_575,N_3862);
nor U8576 (N_8576,N_2494,N_1264);
and U8577 (N_8577,N_3341,N_1807);
nand U8578 (N_8578,N_3934,N_878);
nor U8579 (N_8579,N_4745,N_944);
or U8580 (N_8580,N_4450,N_3192);
and U8581 (N_8581,N_3604,N_162);
nand U8582 (N_8582,N_4545,N_1609);
xnor U8583 (N_8583,N_393,N_161);
nor U8584 (N_8584,N_1460,N_1903);
or U8585 (N_8585,N_4514,N_1624);
nand U8586 (N_8586,N_4171,N_2670);
nor U8587 (N_8587,N_4751,N_1896);
and U8588 (N_8588,N_1528,N_1380);
nor U8589 (N_8589,N_1543,N_467);
nand U8590 (N_8590,N_1887,N_4216);
or U8591 (N_8591,N_3873,N_3259);
nor U8592 (N_8592,N_4137,N_4860);
nand U8593 (N_8593,N_2570,N_2591);
or U8594 (N_8594,N_1745,N_1585);
and U8595 (N_8595,N_4056,N_1576);
nand U8596 (N_8596,N_4321,N_2121);
nand U8597 (N_8597,N_2278,N_2725);
nand U8598 (N_8598,N_2034,N_798);
or U8599 (N_8599,N_3144,N_2541);
and U8600 (N_8600,N_107,N_4596);
nand U8601 (N_8601,N_4114,N_4107);
or U8602 (N_8602,N_2710,N_1482);
and U8603 (N_8603,N_2622,N_2265);
nor U8604 (N_8604,N_1680,N_1374);
or U8605 (N_8605,N_1693,N_239);
or U8606 (N_8606,N_2047,N_3586);
or U8607 (N_8607,N_462,N_1268);
nor U8608 (N_8608,N_253,N_4008);
nor U8609 (N_8609,N_3301,N_1784);
or U8610 (N_8610,N_4103,N_2697);
and U8611 (N_8611,N_4093,N_3435);
or U8612 (N_8612,N_4703,N_616);
or U8613 (N_8613,N_572,N_2339);
nand U8614 (N_8614,N_760,N_1457);
nor U8615 (N_8615,N_1095,N_4522);
and U8616 (N_8616,N_1508,N_2256);
nand U8617 (N_8617,N_1001,N_3882);
nand U8618 (N_8618,N_2131,N_3905);
nor U8619 (N_8619,N_3570,N_262);
and U8620 (N_8620,N_1620,N_1763);
nor U8621 (N_8621,N_366,N_1460);
nand U8622 (N_8622,N_142,N_1035);
nor U8623 (N_8623,N_2285,N_1798);
or U8624 (N_8624,N_4190,N_1425);
nor U8625 (N_8625,N_3929,N_3851);
or U8626 (N_8626,N_4112,N_3027);
nand U8627 (N_8627,N_1306,N_2167);
and U8628 (N_8628,N_2652,N_345);
or U8629 (N_8629,N_851,N_1970);
and U8630 (N_8630,N_4860,N_3202);
nand U8631 (N_8631,N_4504,N_1667);
or U8632 (N_8632,N_3922,N_621);
or U8633 (N_8633,N_1599,N_4405);
or U8634 (N_8634,N_4391,N_3679);
or U8635 (N_8635,N_4598,N_805);
and U8636 (N_8636,N_4329,N_1794);
or U8637 (N_8637,N_88,N_2486);
or U8638 (N_8638,N_2531,N_1853);
nor U8639 (N_8639,N_1865,N_1720);
nand U8640 (N_8640,N_1087,N_1416);
and U8641 (N_8641,N_365,N_2085);
nand U8642 (N_8642,N_4403,N_3711);
xnor U8643 (N_8643,N_358,N_4024);
xnor U8644 (N_8644,N_357,N_1773);
or U8645 (N_8645,N_2185,N_1907);
nand U8646 (N_8646,N_507,N_1064);
nor U8647 (N_8647,N_1586,N_2326);
and U8648 (N_8648,N_2000,N_1237);
nand U8649 (N_8649,N_3676,N_894);
or U8650 (N_8650,N_4581,N_3787);
nor U8651 (N_8651,N_1550,N_3453);
nand U8652 (N_8652,N_3348,N_4674);
and U8653 (N_8653,N_4170,N_4153);
nand U8654 (N_8654,N_1297,N_939);
or U8655 (N_8655,N_3977,N_3990);
nor U8656 (N_8656,N_3079,N_3128);
nand U8657 (N_8657,N_3216,N_1433);
nor U8658 (N_8658,N_1314,N_1943);
and U8659 (N_8659,N_2675,N_89);
and U8660 (N_8660,N_3815,N_1862);
and U8661 (N_8661,N_2867,N_2618);
nand U8662 (N_8662,N_2844,N_1729);
nor U8663 (N_8663,N_4228,N_1023);
nand U8664 (N_8664,N_1202,N_4068);
nand U8665 (N_8665,N_564,N_4248);
nor U8666 (N_8666,N_1624,N_3245);
and U8667 (N_8667,N_117,N_1531);
nand U8668 (N_8668,N_3294,N_2520);
nand U8669 (N_8669,N_2215,N_4630);
or U8670 (N_8670,N_942,N_2642);
or U8671 (N_8671,N_467,N_3174);
and U8672 (N_8672,N_1034,N_1770);
nand U8673 (N_8673,N_3441,N_184);
or U8674 (N_8674,N_4177,N_2148);
and U8675 (N_8675,N_1833,N_1745);
nand U8676 (N_8676,N_2930,N_1368);
xnor U8677 (N_8677,N_3929,N_4966);
and U8678 (N_8678,N_1462,N_3345);
or U8679 (N_8679,N_796,N_626);
or U8680 (N_8680,N_1678,N_2682);
nand U8681 (N_8681,N_4062,N_1047);
and U8682 (N_8682,N_4427,N_2370);
nor U8683 (N_8683,N_2159,N_3342);
nand U8684 (N_8684,N_3303,N_302);
and U8685 (N_8685,N_3478,N_1051);
nor U8686 (N_8686,N_1929,N_4667);
nand U8687 (N_8687,N_2129,N_4255);
or U8688 (N_8688,N_2835,N_764);
nor U8689 (N_8689,N_4381,N_1704);
nand U8690 (N_8690,N_1359,N_3892);
or U8691 (N_8691,N_3439,N_2543);
and U8692 (N_8692,N_1304,N_4779);
and U8693 (N_8693,N_4755,N_4315);
and U8694 (N_8694,N_3642,N_1348);
nand U8695 (N_8695,N_1037,N_4897);
or U8696 (N_8696,N_2970,N_4326);
nor U8697 (N_8697,N_4370,N_3012);
or U8698 (N_8698,N_4849,N_4054);
nand U8699 (N_8699,N_1699,N_4400);
nand U8700 (N_8700,N_1333,N_4140);
nor U8701 (N_8701,N_1731,N_4048);
xnor U8702 (N_8702,N_1113,N_1914);
nor U8703 (N_8703,N_3987,N_2125);
or U8704 (N_8704,N_1478,N_3389);
or U8705 (N_8705,N_3839,N_2500);
and U8706 (N_8706,N_567,N_2187);
nor U8707 (N_8707,N_1874,N_4630);
and U8708 (N_8708,N_2717,N_1714);
nand U8709 (N_8709,N_2239,N_4990);
or U8710 (N_8710,N_4363,N_1134);
nand U8711 (N_8711,N_2077,N_1469);
nor U8712 (N_8712,N_858,N_4071);
nor U8713 (N_8713,N_2642,N_2950);
nand U8714 (N_8714,N_397,N_3172);
nand U8715 (N_8715,N_1677,N_1931);
or U8716 (N_8716,N_375,N_2412);
and U8717 (N_8717,N_529,N_2891);
and U8718 (N_8718,N_674,N_3150);
or U8719 (N_8719,N_2821,N_34);
and U8720 (N_8720,N_134,N_4529);
nand U8721 (N_8721,N_4757,N_821);
and U8722 (N_8722,N_2567,N_711);
and U8723 (N_8723,N_1088,N_4579);
and U8724 (N_8724,N_3335,N_2910);
nor U8725 (N_8725,N_564,N_3960);
or U8726 (N_8726,N_3399,N_4297);
and U8727 (N_8727,N_3857,N_3861);
or U8728 (N_8728,N_2363,N_4703);
nor U8729 (N_8729,N_2735,N_3712);
or U8730 (N_8730,N_962,N_856);
and U8731 (N_8731,N_3674,N_1881);
and U8732 (N_8732,N_3535,N_3216);
and U8733 (N_8733,N_1376,N_3149);
nor U8734 (N_8734,N_1726,N_2128);
or U8735 (N_8735,N_2311,N_4940);
nand U8736 (N_8736,N_2320,N_1634);
nor U8737 (N_8737,N_4090,N_4287);
nor U8738 (N_8738,N_1260,N_3911);
or U8739 (N_8739,N_3038,N_3719);
and U8740 (N_8740,N_1466,N_2376);
nor U8741 (N_8741,N_1718,N_3475);
and U8742 (N_8742,N_2866,N_136);
nor U8743 (N_8743,N_2614,N_3217);
and U8744 (N_8744,N_83,N_741);
nand U8745 (N_8745,N_4423,N_3059);
nor U8746 (N_8746,N_932,N_858);
or U8747 (N_8747,N_4456,N_2182);
and U8748 (N_8748,N_74,N_4815);
nand U8749 (N_8749,N_2428,N_4309);
nor U8750 (N_8750,N_3075,N_3122);
and U8751 (N_8751,N_3320,N_1911);
and U8752 (N_8752,N_1042,N_3755);
nor U8753 (N_8753,N_1467,N_2923);
nor U8754 (N_8754,N_3027,N_2722);
and U8755 (N_8755,N_2482,N_3506);
nor U8756 (N_8756,N_3458,N_984);
nand U8757 (N_8757,N_1429,N_1866);
nand U8758 (N_8758,N_2018,N_4093);
or U8759 (N_8759,N_4998,N_2044);
and U8760 (N_8760,N_4245,N_2651);
and U8761 (N_8761,N_664,N_439);
nor U8762 (N_8762,N_2897,N_3419);
nand U8763 (N_8763,N_1155,N_2335);
nand U8764 (N_8764,N_4688,N_2291);
nor U8765 (N_8765,N_2861,N_2605);
nand U8766 (N_8766,N_4442,N_2164);
and U8767 (N_8767,N_82,N_1470);
nand U8768 (N_8768,N_843,N_3593);
or U8769 (N_8769,N_3247,N_2550);
nor U8770 (N_8770,N_2908,N_164);
and U8771 (N_8771,N_3973,N_4439);
nor U8772 (N_8772,N_3719,N_1232);
nand U8773 (N_8773,N_2193,N_4038);
nand U8774 (N_8774,N_2727,N_4005);
nand U8775 (N_8775,N_4137,N_4222);
nand U8776 (N_8776,N_670,N_321);
nand U8777 (N_8777,N_4112,N_950);
and U8778 (N_8778,N_637,N_2029);
nand U8779 (N_8779,N_4147,N_4888);
nor U8780 (N_8780,N_753,N_4956);
nor U8781 (N_8781,N_2496,N_2570);
and U8782 (N_8782,N_718,N_3731);
and U8783 (N_8783,N_325,N_377);
or U8784 (N_8784,N_4847,N_1302);
or U8785 (N_8785,N_1470,N_289);
and U8786 (N_8786,N_4287,N_2175);
nand U8787 (N_8787,N_3204,N_3471);
and U8788 (N_8788,N_4444,N_3471);
nor U8789 (N_8789,N_1828,N_4802);
or U8790 (N_8790,N_4631,N_1640);
nor U8791 (N_8791,N_1504,N_3897);
nand U8792 (N_8792,N_1506,N_970);
and U8793 (N_8793,N_2551,N_392);
or U8794 (N_8794,N_1234,N_3778);
nor U8795 (N_8795,N_4677,N_218);
nor U8796 (N_8796,N_2749,N_1957);
and U8797 (N_8797,N_4496,N_2100);
nand U8798 (N_8798,N_2959,N_2041);
nor U8799 (N_8799,N_4865,N_4008);
nand U8800 (N_8800,N_3653,N_1198);
nor U8801 (N_8801,N_1688,N_333);
nor U8802 (N_8802,N_212,N_4050);
nor U8803 (N_8803,N_1594,N_884);
nand U8804 (N_8804,N_2669,N_745);
nor U8805 (N_8805,N_3526,N_4851);
nor U8806 (N_8806,N_3272,N_4945);
nand U8807 (N_8807,N_2366,N_3115);
nand U8808 (N_8808,N_3540,N_3691);
nor U8809 (N_8809,N_1974,N_1373);
and U8810 (N_8810,N_1001,N_4481);
or U8811 (N_8811,N_1501,N_2513);
nor U8812 (N_8812,N_3047,N_3227);
nor U8813 (N_8813,N_592,N_1620);
xnor U8814 (N_8814,N_169,N_1925);
nand U8815 (N_8815,N_2693,N_3532);
nand U8816 (N_8816,N_995,N_741);
or U8817 (N_8817,N_3257,N_889);
nand U8818 (N_8818,N_4173,N_917);
or U8819 (N_8819,N_3788,N_1077);
and U8820 (N_8820,N_3982,N_2018);
nor U8821 (N_8821,N_2314,N_3503);
nor U8822 (N_8822,N_1526,N_4606);
nand U8823 (N_8823,N_390,N_0);
or U8824 (N_8824,N_2098,N_4187);
nand U8825 (N_8825,N_443,N_445);
nand U8826 (N_8826,N_2803,N_976);
nor U8827 (N_8827,N_1678,N_2403);
nand U8828 (N_8828,N_4279,N_4412);
nor U8829 (N_8829,N_4764,N_3728);
and U8830 (N_8830,N_466,N_4339);
or U8831 (N_8831,N_2810,N_4902);
or U8832 (N_8832,N_243,N_4988);
nand U8833 (N_8833,N_4750,N_4134);
or U8834 (N_8834,N_1951,N_4119);
nor U8835 (N_8835,N_725,N_4877);
nand U8836 (N_8836,N_1729,N_264);
or U8837 (N_8837,N_1550,N_2346);
or U8838 (N_8838,N_2165,N_1866);
and U8839 (N_8839,N_4934,N_1836);
nand U8840 (N_8840,N_2822,N_3322);
or U8841 (N_8841,N_599,N_2476);
nor U8842 (N_8842,N_2678,N_2708);
or U8843 (N_8843,N_1782,N_4791);
and U8844 (N_8844,N_3820,N_3179);
and U8845 (N_8845,N_925,N_4677);
nand U8846 (N_8846,N_2144,N_2231);
and U8847 (N_8847,N_1025,N_4965);
nand U8848 (N_8848,N_3131,N_2854);
and U8849 (N_8849,N_4636,N_4308);
or U8850 (N_8850,N_3341,N_4683);
and U8851 (N_8851,N_3699,N_3220);
and U8852 (N_8852,N_3972,N_2926);
nor U8853 (N_8853,N_1890,N_2775);
and U8854 (N_8854,N_2664,N_3801);
nand U8855 (N_8855,N_3761,N_1467);
and U8856 (N_8856,N_4255,N_1595);
nand U8857 (N_8857,N_1084,N_356);
xor U8858 (N_8858,N_3368,N_837);
nand U8859 (N_8859,N_2492,N_6);
nand U8860 (N_8860,N_1035,N_1648);
or U8861 (N_8861,N_3155,N_271);
or U8862 (N_8862,N_2338,N_229);
nor U8863 (N_8863,N_4903,N_3953);
nand U8864 (N_8864,N_4615,N_1482);
nor U8865 (N_8865,N_3570,N_598);
and U8866 (N_8866,N_1498,N_3524);
and U8867 (N_8867,N_3986,N_1144);
nor U8868 (N_8868,N_4548,N_1080);
and U8869 (N_8869,N_252,N_2833);
nor U8870 (N_8870,N_3742,N_1503);
nor U8871 (N_8871,N_3172,N_530);
nor U8872 (N_8872,N_4366,N_679);
and U8873 (N_8873,N_4251,N_4656);
nor U8874 (N_8874,N_722,N_3645);
and U8875 (N_8875,N_1266,N_2300);
nor U8876 (N_8876,N_433,N_611);
nand U8877 (N_8877,N_3348,N_3209);
or U8878 (N_8878,N_1556,N_4382);
nand U8879 (N_8879,N_3571,N_3811);
and U8880 (N_8880,N_533,N_3594);
nand U8881 (N_8881,N_3527,N_2092);
nor U8882 (N_8882,N_1836,N_2624);
nand U8883 (N_8883,N_3257,N_4573);
nand U8884 (N_8884,N_1790,N_10);
and U8885 (N_8885,N_1219,N_1640);
and U8886 (N_8886,N_2070,N_3037);
nand U8887 (N_8887,N_2552,N_3360);
nor U8888 (N_8888,N_2602,N_4573);
nand U8889 (N_8889,N_3161,N_2256);
nand U8890 (N_8890,N_4239,N_383);
nand U8891 (N_8891,N_3575,N_654);
nand U8892 (N_8892,N_2028,N_56);
nand U8893 (N_8893,N_930,N_2941);
and U8894 (N_8894,N_789,N_1193);
nand U8895 (N_8895,N_2718,N_4767);
or U8896 (N_8896,N_4955,N_4809);
and U8897 (N_8897,N_4158,N_2108);
and U8898 (N_8898,N_3300,N_3001);
nor U8899 (N_8899,N_3427,N_4589);
nand U8900 (N_8900,N_2119,N_1223);
nor U8901 (N_8901,N_1441,N_3929);
or U8902 (N_8902,N_2070,N_2981);
and U8903 (N_8903,N_3682,N_2032);
and U8904 (N_8904,N_3810,N_1357);
nand U8905 (N_8905,N_1827,N_1775);
and U8906 (N_8906,N_4334,N_3511);
nand U8907 (N_8907,N_1478,N_4380);
or U8908 (N_8908,N_2533,N_914);
nor U8909 (N_8909,N_3540,N_3095);
or U8910 (N_8910,N_2067,N_2265);
and U8911 (N_8911,N_1263,N_2240);
nand U8912 (N_8912,N_437,N_2272);
xnor U8913 (N_8913,N_1842,N_4244);
and U8914 (N_8914,N_4334,N_2564);
and U8915 (N_8915,N_3900,N_4137);
or U8916 (N_8916,N_3088,N_2857);
and U8917 (N_8917,N_3578,N_2597);
nor U8918 (N_8918,N_4086,N_3341);
nor U8919 (N_8919,N_2443,N_2580);
or U8920 (N_8920,N_1848,N_1594);
nor U8921 (N_8921,N_4008,N_1388);
xnor U8922 (N_8922,N_1270,N_3321);
and U8923 (N_8923,N_4716,N_594);
nor U8924 (N_8924,N_3445,N_2598);
nor U8925 (N_8925,N_3880,N_2203);
and U8926 (N_8926,N_3321,N_3005);
and U8927 (N_8927,N_1535,N_1555);
nor U8928 (N_8928,N_4660,N_1308);
nor U8929 (N_8929,N_596,N_2359);
or U8930 (N_8930,N_1836,N_2260);
nor U8931 (N_8931,N_4734,N_2798);
and U8932 (N_8932,N_1597,N_125);
and U8933 (N_8933,N_2885,N_1203);
nand U8934 (N_8934,N_498,N_264);
or U8935 (N_8935,N_3143,N_709);
or U8936 (N_8936,N_2999,N_663);
or U8937 (N_8937,N_2861,N_3401);
or U8938 (N_8938,N_432,N_3881);
nor U8939 (N_8939,N_3962,N_371);
nor U8940 (N_8940,N_4723,N_498);
nand U8941 (N_8941,N_3924,N_872);
and U8942 (N_8942,N_1652,N_1241);
and U8943 (N_8943,N_3872,N_470);
and U8944 (N_8944,N_1675,N_3039);
or U8945 (N_8945,N_618,N_495);
or U8946 (N_8946,N_3177,N_2426);
nor U8947 (N_8947,N_3128,N_3206);
or U8948 (N_8948,N_1366,N_3754);
nand U8949 (N_8949,N_1156,N_2099);
or U8950 (N_8950,N_2390,N_2451);
nor U8951 (N_8951,N_1674,N_2657);
nand U8952 (N_8952,N_2149,N_2648);
nor U8953 (N_8953,N_4241,N_1047);
nand U8954 (N_8954,N_748,N_2823);
nor U8955 (N_8955,N_3105,N_1038);
or U8956 (N_8956,N_384,N_464);
or U8957 (N_8957,N_1141,N_2323);
nor U8958 (N_8958,N_581,N_821);
or U8959 (N_8959,N_34,N_771);
nand U8960 (N_8960,N_3065,N_2937);
nand U8961 (N_8961,N_3301,N_4679);
nand U8962 (N_8962,N_1595,N_3203);
nand U8963 (N_8963,N_1581,N_4012);
and U8964 (N_8964,N_4171,N_2707);
nor U8965 (N_8965,N_4690,N_3851);
or U8966 (N_8966,N_2594,N_2185);
nand U8967 (N_8967,N_3994,N_2430);
or U8968 (N_8968,N_986,N_416);
and U8969 (N_8969,N_800,N_4366);
and U8970 (N_8970,N_271,N_3749);
and U8971 (N_8971,N_15,N_3666);
nand U8972 (N_8972,N_2841,N_3506);
nand U8973 (N_8973,N_52,N_2558);
and U8974 (N_8974,N_978,N_4658);
nor U8975 (N_8975,N_537,N_3757);
nor U8976 (N_8976,N_711,N_3576);
nor U8977 (N_8977,N_1183,N_3271);
and U8978 (N_8978,N_4609,N_4675);
xor U8979 (N_8979,N_2676,N_677);
and U8980 (N_8980,N_682,N_3924);
and U8981 (N_8981,N_1498,N_1231);
nor U8982 (N_8982,N_2263,N_3121);
nor U8983 (N_8983,N_3667,N_1276);
nand U8984 (N_8984,N_3006,N_3012);
and U8985 (N_8985,N_2332,N_296);
or U8986 (N_8986,N_1094,N_3558);
nor U8987 (N_8987,N_948,N_3392);
and U8988 (N_8988,N_3765,N_1331);
and U8989 (N_8989,N_648,N_368);
and U8990 (N_8990,N_4714,N_571);
or U8991 (N_8991,N_4912,N_4067);
nand U8992 (N_8992,N_3423,N_3722);
or U8993 (N_8993,N_898,N_4569);
and U8994 (N_8994,N_2979,N_2214);
nand U8995 (N_8995,N_4122,N_1368);
nand U8996 (N_8996,N_4971,N_4132);
and U8997 (N_8997,N_1618,N_1036);
or U8998 (N_8998,N_1453,N_2796);
xor U8999 (N_8999,N_3844,N_3809);
nor U9000 (N_9000,N_800,N_3734);
nor U9001 (N_9001,N_2726,N_1394);
nor U9002 (N_9002,N_4770,N_1040);
or U9003 (N_9003,N_2753,N_4717);
and U9004 (N_9004,N_2519,N_4020);
or U9005 (N_9005,N_3073,N_2908);
and U9006 (N_9006,N_4615,N_1445);
and U9007 (N_9007,N_2512,N_2933);
or U9008 (N_9008,N_2342,N_277);
nor U9009 (N_9009,N_2356,N_2832);
nand U9010 (N_9010,N_3669,N_2298);
nand U9011 (N_9011,N_583,N_314);
or U9012 (N_9012,N_276,N_2309);
nand U9013 (N_9013,N_636,N_2933);
nand U9014 (N_9014,N_3511,N_3773);
nand U9015 (N_9015,N_3716,N_2286);
nand U9016 (N_9016,N_2041,N_3579);
nor U9017 (N_9017,N_4259,N_3914);
nor U9018 (N_9018,N_4361,N_1155);
nand U9019 (N_9019,N_1780,N_1911);
nor U9020 (N_9020,N_1216,N_373);
and U9021 (N_9021,N_581,N_1907);
or U9022 (N_9022,N_1486,N_1165);
nor U9023 (N_9023,N_250,N_1924);
and U9024 (N_9024,N_4087,N_1716);
and U9025 (N_9025,N_317,N_541);
and U9026 (N_9026,N_3700,N_3567);
and U9027 (N_9027,N_1115,N_328);
and U9028 (N_9028,N_1879,N_4163);
nand U9029 (N_9029,N_4109,N_3224);
nand U9030 (N_9030,N_3045,N_4132);
nand U9031 (N_9031,N_4540,N_2706);
nor U9032 (N_9032,N_3258,N_764);
nor U9033 (N_9033,N_3186,N_3747);
nand U9034 (N_9034,N_995,N_2136);
or U9035 (N_9035,N_1708,N_3370);
and U9036 (N_9036,N_3635,N_996);
or U9037 (N_9037,N_645,N_2590);
and U9038 (N_9038,N_3085,N_4416);
or U9039 (N_9039,N_3799,N_2045);
or U9040 (N_9040,N_4867,N_4035);
and U9041 (N_9041,N_2064,N_3127);
nand U9042 (N_9042,N_2773,N_270);
and U9043 (N_9043,N_2954,N_2377);
and U9044 (N_9044,N_1446,N_4574);
nand U9045 (N_9045,N_4928,N_3435);
or U9046 (N_9046,N_1502,N_1839);
nand U9047 (N_9047,N_2920,N_1326);
and U9048 (N_9048,N_1233,N_1192);
nand U9049 (N_9049,N_1538,N_725);
nor U9050 (N_9050,N_2121,N_4420);
nand U9051 (N_9051,N_1887,N_3688);
nand U9052 (N_9052,N_2662,N_770);
or U9053 (N_9053,N_1852,N_845);
nor U9054 (N_9054,N_2718,N_540);
nand U9055 (N_9055,N_4817,N_2276);
nor U9056 (N_9056,N_3269,N_2163);
or U9057 (N_9057,N_3876,N_1003);
and U9058 (N_9058,N_762,N_2096);
and U9059 (N_9059,N_1380,N_2341);
and U9060 (N_9060,N_2649,N_4357);
and U9061 (N_9061,N_4677,N_3741);
and U9062 (N_9062,N_4637,N_3328);
or U9063 (N_9063,N_1153,N_399);
and U9064 (N_9064,N_2395,N_3936);
nor U9065 (N_9065,N_1647,N_4823);
nand U9066 (N_9066,N_1242,N_1695);
and U9067 (N_9067,N_3614,N_3121);
and U9068 (N_9068,N_1041,N_3349);
nand U9069 (N_9069,N_2615,N_2129);
and U9070 (N_9070,N_1484,N_3279);
nand U9071 (N_9071,N_1674,N_2662);
nor U9072 (N_9072,N_2075,N_1889);
and U9073 (N_9073,N_1901,N_4014);
nand U9074 (N_9074,N_1696,N_2954);
or U9075 (N_9075,N_2324,N_608);
nand U9076 (N_9076,N_4638,N_536);
nand U9077 (N_9077,N_1149,N_3045);
nand U9078 (N_9078,N_1721,N_2178);
nor U9079 (N_9079,N_2413,N_3462);
and U9080 (N_9080,N_549,N_889);
and U9081 (N_9081,N_632,N_3782);
and U9082 (N_9082,N_2037,N_346);
or U9083 (N_9083,N_1737,N_2093);
nand U9084 (N_9084,N_4475,N_3114);
nand U9085 (N_9085,N_2308,N_3788);
nand U9086 (N_9086,N_742,N_3063);
or U9087 (N_9087,N_2475,N_4696);
and U9088 (N_9088,N_2617,N_2615);
and U9089 (N_9089,N_3945,N_1529);
nor U9090 (N_9090,N_3929,N_4493);
nand U9091 (N_9091,N_1234,N_4650);
and U9092 (N_9092,N_273,N_3162);
nand U9093 (N_9093,N_472,N_4165);
nand U9094 (N_9094,N_2078,N_2267);
nand U9095 (N_9095,N_1143,N_3499);
nor U9096 (N_9096,N_3998,N_288);
or U9097 (N_9097,N_1968,N_1167);
nor U9098 (N_9098,N_3629,N_2584);
nand U9099 (N_9099,N_1840,N_397);
nand U9100 (N_9100,N_894,N_4713);
and U9101 (N_9101,N_1719,N_2015);
nor U9102 (N_9102,N_1083,N_162);
nor U9103 (N_9103,N_3117,N_3434);
nand U9104 (N_9104,N_3060,N_4192);
and U9105 (N_9105,N_4933,N_2691);
and U9106 (N_9106,N_4282,N_1442);
nand U9107 (N_9107,N_3579,N_3251);
or U9108 (N_9108,N_249,N_2449);
nand U9109 (N_9109,N_3850,N_2845);
nand U9110 (N_9110,N_3766,N_2000);
nor U9111 (N_9111,N_3195,N_1842);
nor U9112 (N_9112,N_527,N_1211);
and U9113 (N_9113,N_371,N_604);
nor U9114 (N_9114,N_3242,N_162);
or U9115 (N_9115,N_4508,N_3014);
or U9116 (N_9116,N_1398,N_3125);
nor U9117 (N_9117,N_2808,N_1814);
nand U9118 (N_9118,N_1585,N_4501);
and U9119 (N_9119,N_4503,N_4295);
nand U9120 (N_9120,N_2926,N_2187);
or U9121 (N_9121,N_1213,N_2500);
or U9122 (N_9122,N_4925,N_3730);
nand U9123 (N_9123,N_1662,N_2574);
nor U9124 (N_9124,N_3925,N_2229);
or U9125 (N_9125,N_1330,N_3325);
nor U9126 (N_9126,N_2682,N_805);
or U9127 (N_9127,N_64,N_3720);
and U9128 (N_9128,N_2029,N_1056);
nand U9129 (N_9129,N_1375,N_3748);
and U9130 (N_9130,N_2988,N_2186);
and U9131 (N_9131,N_2735,N_2738);
nand U9132 (N_9132,N_4121,N_2836);
nand U9133 (N_9133,N_3443,N_4643);
and U9134 (N_9134,N_1279,N_2481);
nor U9135 (N_9135,N_1491,N_2062);
or U9136 (N_9136,N_4859,N_1904);
nand U9137 (N_9137,N_1920,N_3477);
xor U9138 (N_9138,N_4699,N_165);
and U9139 (N_9139,N_242,N_2461);
or U9140 (N_9140,N_3973,N_1296);
nor U9141 (N_9141,N_2136,N_4565);
nor U9142 (N_9142,N_4249,N_4746);
nand U9143 (N_9143,N_2775,N_1034);
and U9144 (N_9144,N_675,N_4805);
or U9145 (N_9145,N_1735,N_2083);
nand U9146 (N_9146,N_3841,N_2256);
nor U9147 (N_9147,N_1897,N_1439);
nor U9148 (N_9148,N_497,N_1711);
nor U9149 (N_9149,N_40,N_3843);
nand U9150 (N_9150,N_1417,N_4751);
or U9151 (N_9151,N_2120,N_976);
or U9152 (N_9152,N_782,N_3496);
or U9153 (N_9153,N_3195,N_502);
or U9154 (N_9154,N_3640,N_4831);
nor U9155 (N_9155,N_3665,N_4701);
nand U9156 (N_9156,N_1245,N_4617);
nand U9157 (N_9157,N_2314,N_867);
or U9158 (N_9158,N_1900,N_867);
nor U9159 (N_9159,N_1517,N_2708);
nor U9160 (N_9160,N_3905,N_1164);
or U9161 (N_9161,N_1314,N_2608);
nand U9162 (N_9162,N_4745,N_1258);
and U9163 (N_9163,N_4851,N_2072);
nand U9164 (N_9164,N_1611,N_1734);
or U9165 (N_9165,N_3855,N_3044);
nand U9166 (N_9166,N_777,N_502);
xnor U9167 (N_9167,N_3684,N_3746);
nand U9168 (N_9168,N_4363,N_3187);
nor U9169 (N_9169,N_3388,N_1773);
nand U9170 (N_9170,N_3843,N_1704);
or U9171 (N_9171,N_4196,N_159);
and U9172 (N_9172,N_4063,N_2431);
nor U9173 (N_9173,N_3851,N_2267);
nand U9174 (N_9174,N_4327,N_2803);
and U9175 (N_9175,N_4394,N_882);
nand U9176 (N_9176,N_1486,N_2276);
nand U9177 (N_9177,N_874,N_4893);
nand U9178 (N_9178,N_2741,N_1209);
or U9179 (N_9179,N_4194,N_3165);
and U9180 (N_9180,N_4781,N_4442);
or U9181 (N_9181,N_3914,N_1853);
or U9182 (N_9182,N_860,N_2717);
nand U9183 (N_9183,N_2168,N_1647);
or U9184 (N_9184,N_3724,N_3217);
and U9185 (N_9185,N_2795,N_2851);
and U9186 (N_9186,N_2776,N_3254);
and U9187 (N_9187,N_4387,N_2448);
and U9188 (N_9188,N_207,N_4936);
and U9189 (N_9189,N_4311,N_1119);
and U9190 (N_9190,N_356,N_3753);
nand U9191 (N_9191,N_1911,N_1024);
or U9192 (N_9192,N_464,N_293);
nor U9193 (N_9193,N_1517,N_3795);
nor U9194 (N_9194,N_4798,N_75);
nor U9195 (N_9195,N_2890,N_4567);
nand U9196 (N_9196,N_4004,N_1025);
and U9197 (N_9197,N_1412,N_574);
or U9198 (N_9198,N_4458,N_1434);
nand U9199 (N_9199,N_1003,N_1476);
and U9200 (N_9200,N_1899,N_2169);
nor U9201 (N_9201,N_1606,N_3971);
nor U9202 (N_9202,N_1404,N_4878);
or U9203 (N_9203,N_4636,N_3871);
or U9204 (N_9204,N_4280,N_2676);
and U9205 (N_9205,N_3355,N_2957);
nor U9206 (N_9206,N_4536,N_2241);
or U9207 (N_9207,N_2415,N_2497);
or U9208 (N_9208,N_2809,N_4299);
nand U9209 (N_9209,N_4024,N_4815);
and U9210 (N_9210,N_450,N_1828);
or U9211 (N_9211,N_3746,N_1767);
and U9212 (N_9212,N_3182,N_4014);
nor U9213 (N_9213,N_185,N_1659);
nand U9214 (N_9214,N_829,N_1649);
nand U9215 (N_9215,N_3682,N_703);
or U9216 (N_9216,N_4550,N_211);
nand U9217 (N_9217,N_3830,N_2374);
nor U9218 (N_9218,N_1903,N_3881);
or U9219 (N_9219,N_273,N_1547);
or U9220 (N_9220,N_4242,N_1033);
nand U9221 (N_9221,N_3288,N_4172);
and U9222 (N_9222,N_1789,N_2518);
or U9223 (N_9223,N_4103,N_4496);
nor U9224 (N_9224,N_3392,N_133);
and U9225 (N_9225,N_470,N_70);
and U9226 (N_9226,N_2323,N_1117);
nand U9227 (N_9227,N_1648,N_373);
or U9228 (N_9228,N_4175,N_3940);
and U9229 (N_9229,N_4642,N_2383);
and U9230 (N_9230,N_3365,N_1754);
or U9231 (N_9231,N_489,N_4946);
and U9232 (N_9232,N_667,N_1782);
nand U9233 (N_9233,N_902,N_2936);
nand U9234 (N_9234,N_4334,N_2279);
or U9235 (N_9235,N_2527,N_928);
nor U9236 (N_9236,N_2955,N_3568);
and U9237 (N_9237,N_3917,N_3906);
and U9238 (N_9238,N_2994,N_2507);
nor U9239 (N_9239,N_3398,N_3248);
nor U9240 (N_9240,N_3932,N_4011);
or U9241 (N_9241,N_832,N_2736);
nand U9242 (N_9242,N_1144,N_3651);
and U9243 (N_9243,N_4149,N_3814);
or U9244 (N_9244,N_4104,N_27);
nor U9245 (N_9245,N_1644,N_4029);
or U9246 (N_9246,N_4748,N_1454);
nor U9247 (N_9247,N_1793,N_4559);
or U9248 (N_9248,N_4103,N_4877);
nor U9249 (N_9249,N_329,N_3239);
nand U9250 (N_9250,N_3440,N_4571);
nor U9251 (N_9251,N_2987,N_260);
nor U9252 (N_9252,N_2972,N_1499);
nand U9253 (N_9253,N_4217,N_4883);
nor U9254 (N_9254,N_2458,N_2638);
nor U9255 (N_9255,N_3163,N_1263);
nand U9256 (N_9256,N_2019,N_904);
and U9257 (N_9257,N_3301,N_4117);
and U9258 (N_9258,N_1704,N_4224);
nor U9259 (N_9259,N_1564,N_424);
nor U9260 (N_9260,N_3722,N_4634);
nor U9261 (N_9261,N_1825,N_1681);
or U9262 (N_9262,N_1194,N_3609);
nand U9263 (N_9263,N_3547,N_828);
and U9264 (N_9264,N_0,N_2343);
or U9265 (N_9265,N_3851,N_3111);
and U9266 (N_9266,N_4497,N_4260);
and U9267 (N_9267,N_4146,N_1854);
nor U9268 (N_9268,N_2705,N_796);
and U9269 (N_9269,N_3741,N_2670);
nor U9270 (N_9270,N_2164,N_4684);
and U9271 (N_9271,N_937,N_692);
and U9272 (N_9272,N_1794,N_537);
nand U9273 (N_9273,N_839,N_3177);
or U9274 (N_9274,N_425,N_4968);
and U9275 (N_9275,N_238,N_4969);
and U9276 (N_9276,N_883,N_2842);
nor U9277 (N_9277,N_2695,N_361);
or U9278 (N_9278,N_1658,N_3520);
nand U9279 (N_9279,N_3762,N_4896);
nor U9280 (N_9280,N_1259,N_1584);
and U9281 (N_9281,N_364,N_35);
nor U9282 (N_9282,N_2353,N_3453);
nand U9283 (N_9283,N_3784,N_1805);
nand U9284 (N_9284,N_1817,N_206);
or U9285 (N_9285,N_3667,N_4038);
nor U9286 (N_9286,N_55,N_2159);
nand U9287 (N_9287,N_1763,N_161);
or U9288 (N_9288,N_95,N_2655);
or U9289 (N_9289,N_2962,N_533);
nor U9290 (N_9290,N_4425,N_3017);
nor U9291 (N_9291,N_3727,N_4897);
and U9292 (N_9292,N_108,N_1200);
nand U9293 (N_9293,N_4721,N_3088);
and U9294 (N_9294,N_2754,N_4214);
and U9295 (N_9295,N_840,N_2881);
nor U9296 (N_9296,N_2426,N_4225);
nor U9297 (N_9297,N_689,N_3557);
or U9298 (N_9298,N_4879,N_2569);
or U9299 (N_9299,N_3589,N_2853);
nand U9300 (N_9300,N_4228,N_467);
or U9301 (N_9301,N_1002,N_944);
nor U9302 (N_9302,N_4675,N_626);
or U9303 (N_9303,N_1710,N_4199);
nor U9304 (N_9304,N_3251,N_1402);
and U9305 (N_9305,N_2435,N_4226);
nor U9306 (N_9306,N_4870,N_2941);
and U9307 (N_9307,N_3091,N_1267);
nand U9308 (N_9308,N_4460,N_2576);
nor U9309 (N_9309,N_998,N_3798);
and U9310 (N_9310,N_1097,N_4739);
nand U9311 (N_9311,N_849,N_2958);
or U9312 (N_9312,N_2452,N_4564);
or U9313 (N_9313,N_3127,N_3075);
nand U9314 (N_9314,N_3632,N_246);
nand U9315 (N_9315,N_3084,N_2612);
nor U9316 (N_9316,N_572,N_1806);
nand U9317 (N_9317,N_559,N_482);
xnor U9318 (N_9318,N_3888,N_815);
nand U9319 (N_9319,N_4283,N_4300);
and U9320 (N_9320,N_132,N_3700);
and U9321 (N_9321,N_475,N_3209);
nand U9322 (N_9322,N_2350,N_1594);
and U9323 (N_9323,N_1029,N_3549);
or U9324 (N_9324,N_2987,N_1017);
nor U9325 (N_9325,N_2011,N_724);
nor U9326 (N_9326,N_299,N_4206);
nor U9327 (N_9327,N_3914,N_564);
and U9328 (N_9328,N_824,N_2030);
and U9329 (N_9329,N_1406,N_2858);
or U9330 (N_9330,N_1515,N_1498);
and U9331 (N_9331,N_86,N_2159);
and U9332 (N_9332,N_2016,N_1572);
and U9333 (N_9333,N_438,N_4129);
nand U9334 (N_9334,N_2080,N_3938);
nand U9335 (N_9335,N_1625,N_820);
and U9336 (N_9336,N_1904,N_4411);
nand U9337 (N_9337,N_2043,N_951);
nor U9338 (N_9338,N_2837,N_4722);
nor U9339 (N_9339,N_1155,N_1445);
or U9340 (N_9340,N_887,N_1965);
nand U9341 (N_9341,N_3649,N_985);
or U9342 (N_9342,N_3201,N_2616);
or U9343 (N_9343,N_3601,N_4245);
and U9344 (N_9344,N_3938,N_165);
and U9345 (N_9345,N_4064,N_2942);
nor U9346 (N_9346,N_2365,N_987);
nand U9347 (N_9347,N_2337,N_224);
and U9348 (N_9348,N_4552,N_1477);
or U9349 (N_9349,N_1441,N_632);
or U9350 (N_9350,N_3589,N_4092);
nand U9351 (N_9351,N_2571,N_2606);
and U9352 (N_9352,N_423,N_4044);
and U9353 (N_9353,N_241,N_1108);
nand U9354 (N_9354,N_612,N_323);
nor U9355 (N_9355,N_1317,N_4403);
or U9356 (N_9356,N_2043,N_3991);
nand U9357 (N_9357,N_972,N_332);
nand U9358 (N_9358,N_4424,N_2774);
and U9359 (N_9359,N_2663,N_2174);
nand U9360 (N_9360,N_3817,N_4845);
and U9361 (N_9361,N_3805,N_4099);
nand U9362 (N_9362,N_3439,N_2517);
nor U9363 (N_9363,N_2100,N_1505);
and U9364 (N_9364,N_4345,N_4097);
and U9365 (N_9365,N_3645,N_1358);
nand U9366 (N_9366,N_3177,N_4107);
nor U9367 (N_9367,N_3530,N_3463);
nor U9368 (N_9368,N_2612,N_4806);
nor U9369 (N_9369,N_4182,N_4927);
or U9370 (N_9370,N_2288,N_1783);
nand U9371 (N_9371,N_4183,N_4907);
nor U9372 (N_9372,N_3129,N_260);
nor U9373 (N_9373,N_4741,N_4609);
and U9374 (N_9374,N_2820,N_3517);
nor U9375 (N_9375,N_3851,N_1778);
or U9376 (N_9376,N_4674,N_4850);
nor U9377 (N_9377,N_457,N_3381);
nand U9378 (N_9378,N_21,N_685);
and U9379 (N_9379,N_4127,N_458);
nor U9380 (N_9380,N_192,N_3907);
or U9381 (N_9381,N_3811,N_951);
and U9382 (N_9382,N_285,N_2918);
nor U9383 (N_9383,N_3604,N_1352);
xor U9384 (N_9384,N_3149,N_651);
xnor U9385 (N_9385,N_3568,N_1615);
nand U9386 (N_9386,N_145,N_4341);
nor U9387 (N_9387,N_4223,N_2320);
or U9388 (N_9388,N_3463,N_2026);
nor U9389 (N_9389,N_2703,N_698);
or U9390 (N_9390,N_1529,N_759);
nor U9391 (N_9391,N_532,N_1210);
or U9392 (N_9392,N_4248,N_483);
and U9393 (N_9393,N_3221,N_3286);
nor U9394 (N_9394,N_3513,N_4996);
nand U9395 (N_9395,N_108,N_1979);
nand U9396 (N_9396,N_4764,N_2112);
nor U9397 (N_9397,N_290,N_4412);
or U9398 (N_9398,N_3580,N_4490);
nor U9399 (N_9399,N_180,N_444);
nand U9400 (N_9400,N_1105,N_2294);
nand U9401 (N_9401,N_2418,N_682);
or U9402 (N_9402,N_2815,N_2388);
and U9403 (N_9403,N_4263,N_661);
nor U9404 (N_9404,N_2450,N_2077);
nor U9405 (N_9405,N_729,N_2137);
nand U9406 (N_9406,N_3740,N_1418);
nor U9407 (N_9407,N_2215,N_1037);
xor U9408 (N_9408,N_4047,N_2734);
or U9409 (N_9409,N_4935,N_105);
or U9410 (N_9410,N_4468,N_186);
or U9411 (N_9411,N_619,N_1977);
and U9412 (N_9412,N_1257,N_4062);
and U9413 (N_9413,N_3886,N_645);
nand U9414 (N_9414,N_3292,N_3367);
or U9415 (N_9415,N_2591,N_1549);
nand U9416 (N_9416,N_2097,N_1816);
nand U9417 (N_9417,N_3080,N_882);
nand U9418 (N_9418,N_3397,N_620);
and U9419 (N_9419,N_2330,N_1352);
nor U9420 (N_9420,N_2947,N_1465);
and U9421 (N_9421,N_2997,N_1518);
or U9422 (N_9422,N_3814,N_4899);
or U9423 (N_9423,N_985,N_1878);
nor U9424 (N_9424,N_2166,N_2938);
and U9425 (N_9425,N_2243,N_125);
and U9426 (N_9426,N_3806,N_201);
and U9427 (N_9427,N_2721,N_1774);
or U9428 (N_9428,N_3202,N_4064);
nand U9429 (N_9429,N_3927,N_407);
nor U9430 (N_9430,N_998,N_972);
and U9431 (N_9431,N_4786,N_2567);
and U9432 (N_9432,N_4985,N_4176);
xor U9433 (N_9433,N_1048,N_3958);
or U9434 (N_9434,N_2801,N_1702);
nor U9435 (N_9435,N_689,N_4704);
and U9436 (N_9436,N_214,N_2553);
nand U9437 (N_9437,N_2438,N_2436);
xnor U9438 (N_9438,N_221,N_1623);
and U9439 (N_9439,N_3794,N_628);
nor U9440 (N_9440,N_4425,N_4184);
nand U9441 (N_9441,N_1294,N_1365);
or U9442 (N_9442,N_2069,N_3626);
and U9443 (N_9443,N_3955,N_2527);
nor U9444 (N_9444,N_3703,N_2559);
or U9445 (N_9445,N_1821,N_1154);
and U9446 (N_9446,N_3165,N_2668);
nand U9447 (N_9447,N_1164,N_4156);
and U9448 (N_9448,N_4399,N_3001);
and U9449 (N_9449,N_3286,N_3012);
and U9450 (N_9450,N_4614,N_2914);
and U9451 (N_9451,N_3727,N_4625);
or U9452 (N_9452,N_2550,N_1742);
nor U9453 (N_9453,N_3556,N_4409);
xor U9454 (N_9454,N_2015,N_192);
nand U9455 (N_9455,N_2156,N_3510);
nand U9456 (N_9456,N_3823,N_1551);
or U9457 (N_9457,N_2113,N_3369);
nand U9458 (N_9458,N_4452,N_725);
nand U9459 (N_9459,N_2017,N_2949);
or U9460 (N_9460,N_4310,N_3913);
nand U9461 (N_9461,N_3939,N_3100);
nand U9462 (N_9462,N_3555,N_189);
nand U9463 (N_9463,N_661,N_3263);
or U9464 (N_9464,N_1526,N_3483);
and U9465 (N_9465,N_649,N_684);
xor U9466 (N_9466,N_1655,N_896);
nand U9467 (N_9467,N_4706,N_3293);
nand U9468 (N_9468,N_815,N_1563);
nand U9469 (N_9469,N_3883,N_1056);
nor U9470 (N_9470,N_2216,N_2379);
nor U9471 (N_9471,N_167,N_898);
or U9472 (N_9472,N_4679,N_1084);
or U9473 (N_9473,N_2539,N_152);
or U9474 (N_9474,N_1331,N_1788);
and U9475 (N_9475,N_3027,N_1021);
or U9476 (N_9476,N_238,N_1318);
and U9477 (N_9477,N_4311,N_3089);
and U9478 (N_9478,N_2177,N_3063);
nor U9479 (N_9479,N_3459,N_2567);
or U9480 (N_9480,N_3240,N_1849);
and U9481 (N_9481,N_1159,N_1692);
nor U9482 (N_9482,N_2004,N_4754);
and U9483 (N_9483,N_1950,N_1194);
nor U9484 (N_9484,N_4608,N_4043);
nor U9485 (N_9485,N_1019,N_4888);
and U9486 (N_9486,N_1498,N_1746);
nor U9487 (N_9487,N_2285,N_1992);
nand U9488 (N_9488,N_4325,N_705);
nor U9489 (N_9489,N_3972,N_3747);
nand U9490 (N_9490,N_3900,N_2428);
nand U9491 (N_9491,N_2215,N_1475);
or U9492 (N_9492,N_3472,N_1216);
or U9493 (N_9493,N_195,N_3967);
or U9494 (N_9494,N_1182,N_4699);
nor U9495 (N_9495,N_1778,N_1598);
nor U9496 (N_9496,N_4088,N_1349);
nor U9497 (N_9497,N_4951,N_3642);
and U9498 (N_9498,N_2433,N_3971);
nand U9499 (N_9499,N_2752,N_3948);
and U9500 (N_9500,N_1156,N_1790);
nand U9501 (N_9501,N_3961,N_4309);
nor U9502 (N_9502,N_3170,N_4749);
nand U9503 (N_9503,N_3013,N_201);
or U9504 (N_9504,N_3905,N_16);
nor U9505 (N_9505,N_989,N_4305);
nand U9506 (N_9506,N_168,N_190);
and U9507 (N_9507,N_4921,N_1845);
nor U9508 (N_9508,N_3994,N_4639);
and U9509 (N_9509,N_4513,N_2323);
nor U9510 (N_9510,N_3742,N_4278);
nor U9511 (N_9511,N_274,N_316);
and U9512 (N_9512,N_4891,N_4478);
and U9513 (N_9513,N_1669,N_1033);
xor U9514 (N_9514,N_4935,N_3138);
nand U9515 (N_9515,N_1357,N_3513);
and U9516 (N_9516,N_3532,N_3782);
and U9517 (N_9517,N_3258,N_4954);
nand U9518 (N_9518,N_2929,N_3359);
nand U9519 (N_9519,N_2764,N_1873);
or U9520 (N_9520,N_289,N_765);
nor U9521 (N_9521,N_2627,N_1733);
nand U9522 (N_9522,N_2578,N_36);
or U9523 (N_9523,N_3974,N_1019);
nand U9524 (N_9524,N_4935,N_531);
or U9525 (N_9525,N_2018,N_3666);
nand U9526 (N_9526,N_3085,N_738);
nor U9527 (N_9527,N_4699,N_2652);
nand U9528 (N_9528,N_308,N_61);
or U9529 (N_9529,N_2180,N_3351);
nand U9530 (N_9530,N_3335,N_4054);
nor U9531 (N_9531,N_2165,N_2891);
and U9532 (N_9532,N_1401,N_1764);
nand U9533 (N_9533,N_2815,N_694);
and U9534 (N_9534,N_649,N_4212);
nor U9535 (N_9535,N_3886,N_2341);
and U9536 (N_9536,N_1064,N_4840);
nand U9537 (N_9537,N_1949,N_755);
nand U9538 (N_9538,N_4269,N_1263);
nor U9539 (N_9539,N_2157,N_2000);
or U9540 (N_9540,N_2068,N_4983);
nand U9541 (N_9541,N_2262,N_1375);
or U9542 (N_9542,N_4921,N_303);
or U9543 (N_9543,N_4662,N_3810);
or U9544 (N_9544,N_3191,N_951);
xnor U9545 (N_9545,N_3665,N_4028);
nor U9546 (N_9546,N_3915,N_1180);
nor U9547 (N_9547,N_4015,N_1204);
nand U9548 (N_9548,N_1625,N_2055);
and U9549 (N_9549,N_2244,N_4512);
nand U9550 (N_9550,N_3650,N_2493);
and U9551 (N_9551,N_4034,N_2531);
and U9552 (N_9552,N_1688,N_1213);
and U9553 (N_9553,N_3289,N_2773);
nand U9554 (N_9554,N_2779,N_4158);
and U9555 (N_9555,N_2214,N_1874);
nor U9556 (N_9556,N_4474,N_1999);
or U9557 (N_9557,N_4007,N_4336);
and U9558 (N_9558,N_2923,N_665);
nor U9559 (N_9559,N_4759,N_3058);
or U9560 (N_9560,N_3012,N_3283);
and U9561 (N_9561,N_4464,N_176);
nand U9562 (N_9562,N_1246,N_2976);
and U9563 (N_9563,N_2275,N_4520);
nand U9564 (N_9564,N_620,N_1710);
and U9565 (N_9565,N_3171,N_376);
nand U9566 (N_9566,N_2217,N_3334);
and U9567 (N_9567,N_2120,N_2583);
nand U9568 (N_9568,N_3234,N_490);
and U9569 (N_9569,N_3643,N_2004);
or U9570 (N_9570,N_719,N_4688);
nor U9571 (N_9571,N_3783,N_4868);
and U9572 (N_9572,N_2201,N_4279);
nor U9573 (N_9573,N_2980,N_496);
nand U9574 (N_9574,N_2027,N_111);
or U9575 (N_9575,N_4302,N_1457);
nor U9576 (N_9576,N_4747,N_1732);
nor U9577 (N_9577,N_784,N_1907);
nor U9578 (N_9578,N_3952,N_4715);
nor U9579 (N_9579,N_3039,N_4907);
nand U9580 (N_9580,N_854,N_4519);
and U9581 (N_9581,N_3773,N_4257);
nand U9582 (N_9582,N_4619,N_2977);
nor U9583 (N_9583,N_3467,N_2559);
nand U9584 (N_9584,N_3842,N_2693);
or U9585 (N_9585,N_610,N_1682);
nor U9586 (N_9586,N_4251,N_2438);
or U9587 (N_9587,N_3430,N_4944);
nand U9588 (N_9588,N_1072,N_3165);
and U9589 (N_9589,N_3797,N_4352);
nor U9590 (N_9590,N_1971,N_4979);
nand U9591 (N_9591,N_3976,N_2165);
or U9592 (N_9592,N_2256,N_4536);
nand U9593 (N_9593,N_150,N_4016);
and U9594 (N_9594,N_2866,N_2898);
or U9595 (N_9595,N_4114,N_1472);
nor U9596 (N_9596,N_1890,N_307);
nand U9597 (N_9597,N_4924,N_2569);
or U9598 (N_9598,N_3230,N_3416);
or U9599 (N_9599,N_2725,N_3154);
and U9600 (N_9600,N_409,N_192);
nor U9601 (N_9601,N_1493,N_4414);
nor U9602 (N_9602,N_4958,N_2472);
or U9603 (N_9603,N_1177,N_3064);
nand U9604 (N_9604,N_2612,N_723);
nand U9605 (N_9605,N_3767,N_1397);
nor U9606 (N_9606,N_2314,N_3089);
or U9607 (N_9607,N_1558,N_587);
and U9608 (N_9608,N_2354,N_280);
or U9609 (N_9609,N_4695,N_3250);
nand U9610 (N_9610,N_3175,N_4704);
nand U9611 (N_9611,N_1844,N_1428);
and U9612 (N_9612,N_85,N_936);
nand U9613 (N_9613,N_4935,N_2798);
nor U9614 (N_9614,N_3407,N_2917);
or U9615 (N_9615,N_4544,N_4432);
and U9616 (N_9616,N_1223,N_4552);
or U9617 (N_9617,N_2810,N_610);
nand U9618 (N_9618,N_3425,N_2424);
and U9619 (N_9619,N_4163,N_3347);
nor U9620 (N_9620,N_844,N_3669);
nor U9621 (N_9621,N_2165,N_812);
and U9622 (N_9622,N_3466,N_842);
nand U9623 (N_9623,N_4930,N_4180);
nor U9624 (N_9624,N_4190,N_1848);
or U9625 (N_9625,N_2450,N_4543);
nor U9626 (N_9626,N_2527,N_2621);
and U9627 (N_9627,N_3201,N_1357);
nor U9628 (N_9628,N_2181,N_2469);
xnor U9629 (N_9629,N_2320,N_581);
or U9630 (N_9630,N_2208,N_2006);
nand U9631 (N_9631,N_1606,N_1482);
and U9632 (N_9632,N_3139,N_1403);
or U9633 (N_9633,N_1265,N_1079);
and U9634 (N_9634,N_796,N_3538);
nor U9635 (N_9635,N_3227,N_10);
nor U9636 (N_9636,N_3592,N_3359);
nand U9637 (N_9637,N_2127,N_1560);
nor U9638 (N_9638,N_2246,N_3616);
nand U9639 (N_9639,N_388,N_4869);
or U9640 (N_9640,N_223,N_4522);
or U9641 (N_9641,N_4566,N_3960);
nor U9642 (N_9642,N_3199,N_2648);
or U9643 (N_9643,N_1012,N_275);
nand U9644 (N_9644,N_1084,N_1031);
and U9645 (N_9645,N_4390,N_4612);
or U9646 (N_9646,N_1050,N_1600);
and U9647 (N_9647,N_864,N_4850);
nand U9648 (N_9648,N_153,N_4608);
or U9649 (N_9649,N_1168,N_1289);
nand U9650 (N_9650,N_4146,N_4855);
and U9651 (N_9651,N_2202,N_1099);
nor U9652 (N_9652,N_4736,N_2487);
nand U9653 (N_9653,N_3738,N_262);
and U9654 (N_9654,N_2814,N_783);
or U9655 (N_9655,N_1117,N_4381);
nor U9656 (N_9656,N_1274,N_425);
nor U9657 (N_9657,N_1600,N_1518);
or U9658 (N_9658,N_3106,N_2687);
nand U9659 (N_9659,N_1777,N_2461);
and U9660 (N_9660,N_184,N_1755);
nor U9661 (N_9661,N_499,N_3499);
nor U9662 (N_9662,N_2783,N_2050);
nor U9663 (N_9663,N_3307,N_2858);
nand U9664 (N_9664,N_4636,N_1452);
nand U9665 (N_9665,N_3566,N_2764);
nor U9666 (N_9666,N_4617,N_4961);
or U9667 (N_9667,N_1258,N_1874);
or U9668 (N_9668,N_4097,N_734);
or U9669 (N_9669,N_1280,N_4394);
nor U9670 (N_9670,N_835,N_1939);
nor U9671 (N_9671,N_1122,N_4712);
nand U9672 (N_9672,N_3855,N_4905);
nor U9673 (N_9673,N_3752,N_377);
or U9674 (N_9674,N_537,N_4776);
and U9675 (N_9675,N_2461,N_1162);
or U9676 (N_9676,N_886,N_3824);
or U9677 (N_9677,N_2829,N_3351);
or U9678 (N_9678,N_3927,N_4705);
or U9679 (N_9679,N_3214,N_2699);
and U9680 (N_9680,N_2995,N_4025);
nand U9681 (N_9681,N_1465,N_1108);
nand U9682 (N_9682,N_119,N_2153);
nor U9683 (N_9683,N_2126,N_4594);
nand U9684 (N_9684,N_1288,N_1036);
nor U9685 (N_9685,N_3531,N_2201);
nand U9686 (N_9686,N_4372,N_2229);
nand U9687 (N_9687,N_1189,N_1626);
nor U9688 (N_9688,N_3119,N_4166);
nand U9689 (N_9689,N_4759,N_156);
and U9690 (N_9690,N_1248,N_2009);
nand U9691 (N_9691,N_312,N_4612);
or U9692 (N_9692,N_3810,N_4033);
and U9693 (N_9693,N_2627,N_2874);
or U9694 (N_9694,N_2869,N_3506);
and U9695 (N_9695,N_3002,N_2862);
nand U9696 (N_9696,N_2776,N_1194);
and U9697 (N_9697,N_4368,N_1279);
or U9698 (N_9698,N_4878,N_1027);
or U9699 (N_9699,N_1351,N_248);
nor U9700 (N_9700,N_3892,N_1357);
nand U9701 (N_9701,N_3432,N_2943);
nor U9702 (N_9702,N_2027,N_340);
or U9703 (N_9703,N_4551,N_3188);
and U9704 (N_9704,N_4476,N_4128);
nor U9705 (N_9705,N_446,N_13);
nor U9706 (N_9706,N_3917,N_641);
and U9707 (N_9707,N_4084,N_4428);
and U9708 (N_9708,N_932,N_2777);
nand U9709 (N_9709,N_4455,N_571);
nor U9710 (N_9710,N_3825,N_2845);
nand U9711 (N_9711,N_3899,N_2879);
and U9712 (N_9712,N_3066,N_3083);
and U9713 (N_9713,N_862,N_278);
or U9714 (N_9714,N_4506,N_3259);
or U9715 (N_9715,N_1466,N_808);
and U9716 (N_9716,N_1381,N_3818);
nand U9717 (N_9717,N_2103,N_1309);
nor U9718 (N_9718,N_4410,N_4720);
nand U9719 (N_9719,N_3851,N_4317);
or U9720 (N_9720,N_4695,N_306);
nand U9721 (N_9721,N_2195,N_3424);
nand U9722 (N_9722,N_3189,N_2337);
nor U9723 (N_9723,N_3028,N_2698);
and U9724 (N_9724,N_1575,N_4852);
and U9725 (N_9725,N_1409,N_4711);
or U9726 (N_9726,N_1237,N_2167);
nor U9727 (N_9727,N_429,N_1599);
nor U9728 (N_9728,N_2494,N_2642);
nor U9729 (N_9729,N_3858,N_4668);
and U9730 (N_9730,N_4075,N_2387);
and U9731 (N_9731,N_3929,N_3515);
or U9732 (N_9732,N_2682,N_2064);
and U9733 (N_9733,N_4612,N_3129);
and U9734 (N_9734,N_2641,N_3018);
nand U9735 (N_9735,N_3453,N_1520);
and U9736 (N_9736,N_2392,N_2192);
and U9737 (N_9737,N_3678,N_2047);
nand U9738 (N_9738,N_1034,N_1537);
and U9739 (N_9739,N_1914,N_1181);
nand U9740 (N_9740,N_3037,N_2135);
or U9741 (N_9741,N_4700,N_2395);
nand U9742 (N_9742,N_4677,N_1625);
or U9743 (N_9743,N_3170,N_2362);
or U9744 (N_9744,N_4968,N_2370);
nand U9745 (N_9745,N_3836,N_4503);
nor U9746 (N_9746,N_4629,N_656);
nand U9747 (N_9747,N_1548,N_1873);
and U9748 (N_9748,N_818,N_3260);
nand U9749 (N_9749,N_4801,N_4655);
or U9750 (N_9750,N_1121,N_996);
nand U9751 (N_9751,N_1995,N_2026);
nand U9752 (N_9752,N_2260,N_4555);
and U9753 (N_9753,N_1775,N_1986);
nand U9754 (N_9754,N_3657,N_4760);
or U9755 (N_9755,N_1231,N_925);
nor U9756 (N_9756,N_4559,N_4363);
or U9757 (N_9757,N_462,N_4317);
or U9758 (N_9758,N_980,N_468);
or U9759 (N_9759,N_2255,N_4113);
nand U9760 (N_9760,N_1800,N_4330);
or U9761 (N_9761,N_4532,N_4957);
nand U9762 (N_9762,N_2614,N_2821);
and U9763 (N_9763,N_3241,N_2714);
nand U9764 (N_9764,N_4221,N_1022);
and U9765 (N_9765,N_3821,N_973);
nand U9766 (N_9766,N_3689,N_1471);
nand U9767 (N_9767,N_266,N_4368);
or U9768 (N_9768,N_3083,N_2725);
nor U9769 (N_9769,N_4478,N_2388);
and U9770 (N_9770,N_2371,N_2015);
and U9771 (N_9771,N_3997,N_2515);
and U9772 (N_9772,N_1087,N_3466);
or U9773 (N_9773,N_2723,N_540);
nor U9774 (N_9774,N_1346,N_875);
xnor U9775 (N_9775,N_1699,N_488);
nor U9776 (N_9776,N_1223,N_3492);
or U9777 (N_9777,N_4996,N_1256);
and U9778 (N_9778,N_4834,N_1871);
nor U9779 (N_9779,N_1854,N_3450);
nand U9780 (N_9780,N_3212,N_4720);
and U9781 (N_9781,N_1119,N_1172);
nand U9782 (N_9782,N_1422,N_1110);
nand U9783 (N_9783,N_4272,N_1798);
nor U9784 (N_9784,N_2114,N_3499);
nor U9785 (N_9785,N_885,N_2084);
and U9786 (N_9786,N_1118,N_2861);
and U9787 (N_9787,N_3535,N_2082);
or U9788 (N_9788,N_1520,N_4786);
or U9789 (N_9789,N_4408,N_386);
nor U9790 (N_9790,N_3832,N_1592);
and U9791 (N_9791,N_1551,N_3223);
nand U9792 (N_9792,N_4969,N_2622);
or U9793 (N_9793,N_767,N_4211);
nor U9794 (N_9794,N_2591,N_1842);
and U9795 (N_9795,N_1640,N_2993);
nor U9796 (N_9796,N_2198,N_1897);
nand U9797 (N_9797,N_3387,N_3473);
or U9798 (N_9798,N_3070,N_3039);
nand U9799 (N_9799,N_2934,N_1116);
or U9800 (N_9800,N_2540,N_4752);
nor U9801 (N_9801,N_2982,N_708);
nand U9802 (N_9802,N_776,N_1811);
or U9803 (N_9803,N_2848,N_677);
nand U9804 (N_9804,N_1313,N_2258);
and U9805 (N_9805,N_1878,N_3249);
nand U9806 (N_9806,N_1845,N_1950);
or U9807 (N_9807,N_4631,N_1178);
and U9808 (N_9808,N_275,N_3921);
or U9809 (N_9809,N_2493,N_4100);
and U9810 (N_9810,N_599,N_1901);
or U9811 (N_9811,N_246,N_4054);
or U9812 (N_9812,N_3667,N_1313);
nand U9813 (N_9813,N_2539,N_3852);
nand U9814 (N_9814,N_3484,N_3848);
and U9815 (N_9815,N_1287,N_1544);
and U9816 (N_9816,N_2650,N_522);
nand U9817 (N_9817,N_1424,N_2411);
nand U9818 (N_9818,N_2951,N_998);
nor U9819 (N_9819,N_2462,N_2755);
or U9820 (N_9820,N_1943,N_2030);
or U9821 (N_9821,N_1190,N_747);
or U9822 (N_9822,N_4107,N_4286);
and U9823 (N_9823,N_3856,N_497);
nand U9824 (N_9824,N_1985,N_4214);
nor U9825 (N_9825,N_3230,N_2127);
and U9826 (N_9826,N_448,N_4804);
nand U9827 (N_9827,N_516,N_3835);
nand U9828 (N_9828,N_1690,N_2543);
nand U9829 (N_9829,N_2062,N_3681);
nor U9830 (N_9830,N_3616,N_2298);
or U9831 (N_9831,N_2866,N_1398);
xnor U9832 (N_9832,N_4242,N_4553);
nor U9833 (N_9833,N_2240,N_4367);
nand U9834 (N_9834,N_3709,N_1493);
or U9835 (N_9835,N_385,N_3918);
or U9836 (N_9836,N_3199,N_4623);
and U9837 (N_9837,N_1520,N_1434);
and U9838 (N_9838,N_3732,N_1258);
or U9839 (N_9839,N_1756,N_3248);
nor U9840 (N_9840,N_3339,N_2917);
nor U9841 (N_9841,N_4261,N_4238);
and U9842 (N_9842,N_1753,N_1542);
and U9843 (N_9843,N_2166,N_3155);
and U9844 (N_9844,N_2787,N_1135);
and U9845 (N_9845,N_3282,N_2928);
nand U9846 (N_9846,N_2500,N_167);
or U9847 (N_9847,N_3515,N_799);
nand U9848 (N_9848,N_3477,N_4876);
xor U9849 (N_9849,N_997,N_817);
nor U9850 (N_9850,N_2962,N_2968);
nor U9851 (N_9851,N_2122,N_2142);
nand U9852 (N_9852,N_2493,N_3775);
and U9853 (N_9853,N_3730,N_2723);
nor U9854 (N_9854,N_967,N_1642);
nand U9855 (N_9855,N_2044,N_221);
nand U9856 (N_9856,N_3331,N_2109);
or U9857 (N_9857,N_4123,N_2780);
and U9858 (N_9858,N_3655,N_3275);
nand U9859 (N_9859,N_3907,N_2203);
nand U9860 (N_9860,N_101,N_3237);
nand U9861 (N_9861,N_2716,N_2234);
or U9862 (N_9862,N_3972,N_1106);
nand U9863 (N_9863,N_3807,N_1841);
and U9864 (N_9864,N_4437,N_2275);
nand U9865 (N_9865,N_227,N_3110);
or U9866 (N_9866,N_2598,N_4436);
or U9867 (N_9867,N_126,N_349);
or U9868 (N_9868,N_4477,N_4236);
nand U9869 (N_9869,N_1669,N_1516);
nand U9870 (N_9870,N_777,N_977);
or U9871 (N_9871,N_2466,N_781);
nand U9872 (N_9872,N_4736,N_561);
nand U9873 (N_9873,N_4704,N_4211);
and U9874 (N_9874,N_1559,N_2669);
nor U9875 (N_9875,N_208,N_4147);
nor U9876 (N_9876,N_4595,N_3572);
nand U9877 (N_9877,N_3262,N_4909);
or U9878 (N_9878,N_4547,N_4636);
and U9879 (N_9879,N_1954,N_4850);
nor U9880 (N_9880,N_1889,N_527);
nor U9881 (N_9881,N_877,N_1175);
or U9882 (N_9882,N_2386,N_221);
and U9883 (N_9883,N_1125,N_3690);
nor U9884 (N_9884,N_3068,N_179);
nand U9885 (N_9885,N_509,N_2978);
nor U9886 (N_9886,N_37,N_4379);
nor U9887 (N_9887,N_3064,N_649);
or U9888 (N_9888,N_3982,N_2975);
nor U9889 (N_9889,N_127,N_2938);
or U9890 (N_9890,N_3492,N_1949);
and U9891 (N_9891,N_2484,N_2734);
and U9892 (N_9892,N_2862,N_4468);
nand U9893 (N_9893,N_2324,N_2989);
and U9894 (N_9894,N_4307,N_900);
and U9895 (N_9895,N_4423,N_2753);
nor U9896 (N_9896,N_3065,N_2443);
or U9897 (N_9897,N_3189,N_3123);
nand U9898 (N_9898,N_1785,N_1813);
nor U9899 (N_9899,N_4637,N_2441);
nand U9900 (N_9900,N_1514,N_3469);
and U9901 (N_9901,N_4005,N_55);
and U9902 (N_9902,N_405,N_914);
nand U9903 (N_9903,N_2872,N_2517);
or U9904 (N_9904,N_860,N_388);
nor U9905 (N_9905,N_65,N_937);
nor U9906 (N_9906,N_699,N_3652);
nor U9907 (N_9907,N_927,N_3414);
and U9908 (N_9908,N_3346,N_1055);
nor U9909 (N_9909,N_4134,N_3071);
nor U9910 (N_9910,N_4314,N_2192);
and U9911 (N_9911,N_4056,N_2355);
nand U9912 (N_9912,N_4480,N_483);
or U9913 (N_9913,N_4072,N_2624);
nand U9914 (N_9914,N_877,N_113);
nand U9915 (N_9915,N_3440,N_4257);
nand U9916 (N_9916,N_2279,N_3869);
nand U9917 (N_9917,N_2253,N_2847);
and U9918 (N_9918,N_1359,N_3565);
nor U9919 (N_9919,N_433,N_1726);
or U9920 (N_9920,N_632,N_3071);
or U9921 (N_9921,N_4244,N_4);
nor U9922 (N_9922,N_894,N_916);
and U9923 (N_9923,N_3107,N_361);
or U9924 (N_9924,N_2319,N_2504);
and U9925 (N_9925,N_2392,N_2775);
or U9926 (N_9926,N_3507,N_2810);
xor U9927 (N_9927,N_3416,N_4201);
xor U9928 (N_9928,N_3783,N_2988);
or U9929 (N_9929,N_2530,N_1537);
or U9930 (N_9930,N_55,N_361);
nand U9931 (N_9931,N_935,N_1084);
or U9932 (N_9932,N_530,N_2994);
and U9933 (N_9933,N_1245,N_1677);
nand U9934 (N_9934,N_3742,N_2139);
or U9935 (N_9935,N_1852,N_2002);
or U9936 (N_9936,N_3533,N_294);
nand U9937 (N_9937,N_3185,N_2625);
nor U9938 (N_9938,N_2782,N_82);
nor U9939 (N_9939,N_2272,N_1319);
nand U9940 (N_9940,N_1690,N_1017);
nor U9941 (N_9941,N_4707,N_4590);
nand U9942 (N_9942,N_703,N_2462);
or U9943 (N_9943,N_1219,N_1027);
or U9944 (N_9944,N_1260,N_4211);
or U9945 (N_9945,N_3547,N_2836);
or U9946 (N_9946,N_2975,N_1821);
and U9947 (N_9947,N_2772,N_4348);
nand U9948 (N_9948,N_4388,N_3913);
nand U9949 (N_9949,N_2178,N_4713);
nor U9950 (N_9950,N_2732,N_631);
and U9951 (N_9951,N_3483,N_1931);
nand U9952 (N_9952,N_2321,N_2424);
and U9953 (N_9953,N_711,N_4048);
or U9954 (N_9954,N_2842,N_4009);
nand U9955 (N_9955,N_4400,N_185);
nand U9956 (N_9956,N_4178,N_2071);
nand U9957 (N_9957,N_186,N_2913);
nor U9958 (N_9958,N_950,N_1158);
nor U9959 (N_9959,N_1764,N_4891);
nand U9960 (N_9960,N_698,N_1369);
and U9961 (N_9961,N_3052,N_4480);
nor U9962 (N_9962,N_4919,N_2857);
or U9963 (N_9963,N_3672,N_1436);
nor U9964 (N_9964,N_3928,N_2841);
and U9965 (N_9965,N_1685,N_1103);
and U9966 (N_9966,N_3026,N_2469);
and U9967 (N_9967,N_3916,N_93);
nand U9968 (N_9968,N_2831,N_595);
nand U9969 (N_9969,N_3310,N_4097);
and U9970 (N_9970,N_4237,N_3899);
nor U9971 (N_9971,N_742,N_377);
nand U9972 (N_9972,N_1533,N_3533);
nand U9973 (N_9973,N_3225,N_2822);
nand U9974 (N_9974,N_1981,N_3881);
nand U9975 (N_9975,N_439,N_2827);
or U9976 (N_9976,N_1884,N_2042);
nor U9977 (N_9977,N_2318,N_3984);
nand U9978 (N_9978,N_2940,N_1948);
nor U9979 (N_9979,N_152,N_715);
and U9980 (N_9980,N_4154,N_3766);
nand U9981 (N_9981,N_2075,N_3095);
or U9982 (N_9982,N_2670,N_3189);
nand U9983 (N_9983,N_4535,N_1883);
or U9984 (N_9984,N_659,N_2808);
and U9985 (N_9985,N_3765,N_4948);
or U9986 (N_9986,N_4047,N_856);
or U9987 (N_9987,N_3734,N_3415);
nand U9988 (N_9988,N_3539,N_4469);
and U9989 (N_9989,N_4056,N_3268);
or U9990 (N_9990,N_63,N_883);
or U9991 (N_9991,N_1593,N_455);
nand U9992 (N_9992,N_542,N_1792);
or U9993 (N_9993,N_34,N_1384);
nor U9994 (N_9994,N_333,N_128);
and U9995 (N_9995,N_2598,N_3995);
nand U9996 (N_9996,N_4028,N_612);
nor U9997 (N_9997,N_1583,N_4999);
xor U9998 (N_9998,N_3466,N_3268);
nand U9999 (N_9999,N_2152,N_2141);
and UO_0 (O_0,N_9771,N_9577);
or UO_1 (O_1,N_6903,N_5930);
and UO_2 (O_2,N_5067,N_8959);
and UO_3 (O_3,N_6193,N_8808);
xnor UO_4 (O_4,N_6948,N_6357);
and UO_5 (O_5,N_7384,N_6319);
nor UO_6 (O_6,N_7174,N_6028);
nand UO_7 (O_7,N_5761,N_9756);
nor UO_8 (O_8,N_5918,N_5404);
nand UO_9 (O_9,N_6512,N_7774);
and UO_10 (O_10,N_6770,N_5876);
and UO_11 (O_11,N_8750,N_9229);
nand UO_12 (O_12,N_9420,N_8668);
nor UO_13 (O_13,N_9408,N_6789);
or UO_14 (O_14,N_5383,N_6934);
and UO_15 (O_15,N_6620,N_7622);
nand UO_16 (O_16,N_5784,N_6020);
and UO_17 (O_17,N_7363,N_9601);
nor UO_18 (O_18,N_6187,N_6264);
and UO_19 (O_19,N_5965,N_5433);
and UO_20 (O_20,N_8924,N_8384);
nand UO_21 (O_21,N_6541,N_6091);
and UO_22 (O_22,N_5599,N_9707);
or UO_23 (O_23,N_7080,N_5622);
nor UO_24 (O_24,N_9659,N_6731);
or UO_25 (O_25,N_8089,N_5739);
nor UO_26 (O_26,N_8921,N_7752);
and UO_27 (O_27,N_5580,N_5139);
nor UO_28 (O_28,N_6073,N_5280);
or UO_29 (O_29,N_6261,N_7579);
nor UO_30 (O_30,N_5571,N_9445);
nand UO_31 (O_31,N_7568,N_8457);
and UO_32 (O_32,N_9563,N_8938);
or UO_33 (O_33,N_7414,N_8615);
nor UO_34 (O_34,N_5933,N_8854);
nand UO_35 (O_35,N_6463,N_8720);
or UO_36 (O_36,N_9073,N_6806);
nor UO_37 (O_37,N_9672,N_8942);
and UO_38 (O_38,N_7743,N_7625);
and UO_39 (O_39,N_9622,N_5665);
nand UO_40 (O_40,N_9608,N_6672);
nor UO_41 (O_41,N_8125,N_9815);
nand UO_42 (O_42,N_7633,N_7137);
or UO_43 (O_43,N_5693,N_9744);
or UO_44 (O_44,N_6895,N_8161);
nor UO_45 (O_45,N_8440,N_8989);
and UO_46 (O_46,N_8629,N_8986);
nor UO_47 (O_47,N_6059,N_8988);
nand UO_48 (O_48,N_5824,N_8110);
nor UO_49 (O_49,N_6314,N_5012);
nor UO_50 (O_50,N_9027,N_8180);
or UO_51 (O_51,N_9400,N_7531);
nand UO_52 (O_52,N_7772,N_8920);
nor UO_53 (O_53,N_8168,N_6348);
or UO_54 (O_54,N_8639,N_8330);
and UO_55 (O_55,N_7157,N_8607);
nand UO_56 (O_56,N_5114,N_6669);
and UO_57 (O_57,N_8548,N_8382);
nor UO_58 (O_58,N_8796,N_8401);
nand UO_59 (O_59,N_9728,N_7381);
and UO_60 (O_60,N_5407,N_9307);
nor UO_61 (O_61,N_9240,N_5745);
nor UO_62 (O_62,N_9721,N_7515);
and UO_63 (O_63,N_7972,N_5578);
and UO_64 (O_64,N_6009,N_7527);
or UO_65 (O_65,N_6554,N_5830);
or UO_66 (O_66,N_5440,N_6379);
nand UO_67 (O_67,N_6698,N_6859);
or UO_68 (O_68,N_5983,N_8383);
and UO_69 (O_69,N_6837,N_8503);
nand UO_70 (O_70,N_8289,N_7204);
and UO_71 (O_71,N_6253,N_8293);
or UO_72 (O_72,N_7061,N_8357);
or UO_73 (O_73,N_8941,N_9546);
nor UO_74 (O_74,N_6579,N_9607);
and UO_75 (O_75,N_7053,N_8380);
and UO_76 (O_76,N_7993,N_8890);
nor UO_77 (O_77,N_5333,N_9545);
nand UO_78 (O_78,N_5191,N_5102);
xnor UO_79 (O_79,N_7698,N_8037);
and UO_80 (O_80,N_9138,N_7407);
nand UO_81 (O_81,N_5699,N_7911);
nand UO_82 (O_82,N_5397,N_7702);
nor UO_83 (O_83,N_8041,N_9317);
or UO_84 (O_84,N_7282,N_8431);
nor UO_85 (O_85,N_8079,N_5766);
or UO_86 (O_86,N_8265,N_5522);
nor UO_87 (O_87,N_7941,N_9414);
nand UO_88 (O_88,N_6492,N_7055);
and UO_89 (O_89,N_7188,N_9915);
and UO_90 (O_90,N_8246,N_9781);
nand UO_91 (O_91,N_5121,N_5332);
and UO_92 (O_92,N_9191,N_9823);
and UO_93 (O_93,N_7025,N_5411);
nand UO_94 (O_94,N_6323,N_5301);
or UO_95 (O_95,N_9626,N_7769);
or UO_96 (O_96,N_7651,N_7899);
or UO_97 (O_97,N_7646,N_6537);
or UO_98 (O_98,N_7992,N_9597);
nand UO_99 (O_99,N_7526,N_6234);
or UO_100 (O_100,N_6000,N_9247);
and UO_101 (O_101,N_6795,N_7467);
nand UO_102 (O_102,N_9740,N_9000);
or UO_103 (O_103,N_5452,N_8755);
and UO_104 (O_104,N_9074,N_7555);
nor UO_105 (O_105,N_7288,N_6036);
nand UO_106 (O_106,N_5620,N_5006);
and UO_107 (O_107,N_6787,N_5808);
nor UO_108 (O_108,N_6912,N_7541);
nand UO_109 (O_109,N_6160,N_9984);
nand UO_110 (O_110,N_7585,N_7222);
or UO_111 (O_111,N_7105,N_7889);
nor UO_112 (O_112,N_6128,N_5753);
and UO_113 (O_113,N_8785,N_5449);
nor UO_114 (O_114,N_9853,N_5386);
nor UO_115 (O_115,N_6729,N_8099);
nand UO_116 (O_116,N_5773,N_5828);
or UO_117 (O_117,N_8622,N_8308);
nor UO_118 (O_118,N_6716,N_5178);
nor UO_119 (O_119,N_5291,N_5647);
and UO_120 (O_120,N_9471,N_5169);
and UO_121 (O_121,N_5970,N_8351);
or UO_122 (O_122,N_7897,N_5678);
or UO_123 (O_123,N_9560,N_8956);
or UO_124 (O_124,N_8208,N_5216);
nand UO_125 (O_125,N_5335,N_9557);
or UO_126 (O_126,N_5323,N_9169);
or UO_127 (O_127,N_6515,N_6227);
nor UO_128 (O_128,N_6797,N_8459);
nand UO_129 (O_129,N_7716,N_6821);
and UO_130 (O_130,N_6500,N_6468);
nor UO_131 (O_131,N_8723,N_7162);
nand UO_132 (O_132,N_8582,N_9200);
and UO_133 (O_133,N_6016,N_8837);
or UO_134 (O_134,N_7424,N_8331);
nor UO_135 (O_135,N_5330,N_7106);
nor UO_136 (O_136,N_5023,N_8297);
nand UO_137 (O_137,N_7655,N_7130);
or UO_138 (O_138,N_5146,N_8193);
and UO_139 (O_139,N_5909,N_5130);
nand UO_140 (O_140,N_6351,N_8824);
nor UO_141 (O_141,N_5061,N_7054);
nand UO_142 (O_142,N_8427,N_8029);
or UO_143 (O_143,N_6218,N_5062);
nand UO_144 (O_144,N_5629,N_6131);
and UO_145 (O_145,N_5305,N_9023);
and UO_146 (O_146,N_5233,N_8196);
and UO_147 (O_147,N_6876,N_7310);
nand UO_148 (O_148,N_7375,N_6400);
or UO_149 (O_149,N_9924,N_9848);
nand UO_150 (O_150,N_5314,N_8525);
or UO_151 (O_151,N_7994,N_8329);
and UO_152 (O_152,N_6423,N_5247);
and UO_153 (O_153,N_9393,N_8189);
or UO_154 (O_154,N_5715,N_8939);
and UO_155 (O_155,N_8157,N_7015);
and UO_156 (O_156,N_6265,N_9437);
nor UO_157 (O_157,N_8368,N_6947);
nor UO_158 (O_158,N_9183,N_8577);
nand UO_159 (O_159,N_7160,N_7408);
nand UO_160 (O_160,N_9215,N_6258);
nand UO_161 (O_161,N_9892,N_9035);
nor UO_162 (O_162,N_8150,N_8520);
and UO_163 (O_163,N_8226,N_6842);
nor UO_164 (O_164,N_9658,N_9602);
nand UO_165 (O_165,N_8913,N_9660);
and UO_166 (O_166,N_8828,N_7166);
nand UO_167 (O_167,N_9613,N_7165);
and UO_168 (O_168,N_7864,N_6869);
nand UO_169 (O_169,N_8515,N_7668);
nor UO_170 (O_170,N_5357,N_9012);
and UO_171 (O_171,N_6014,N_5221);
nand UO_172 (O_172,N_9682,N_6219);
nor UO_173 (O_173,N_5765,N_6018);
and UO_174 (O_174,N_8376,N_6827);
and UO_175 (O_175,N_7938,N_6157);
and UO_176 (O_176,N_7001,N_9795);
and UO_177 (O_177,N_5995,N_8145);
and UO_178 (O_178,N_9278,N_5757);
nand UO_179 (O_179,N_7308,N_6437);
and UO_180 (O_180,N_7559,N_8983);
and UO_181 (O_181,N_8230,N_8809);
nand UO_182 (O_182,N_9401,N_5858);
nor UO_183 (O_183,N_9446,N_9640);
and UO_184 (O_184,N_5657,N_9881);
nor UO_185 (O_185,N_7194,N_6617);
nor UO_186 (O_186,N_7476,N_6360);
nand UO_187 (O_187,N_5512,N_5103);
nand UO_188 (O_188,N_8497,N_5189);
nand UO_189 (O_189,N_8963,N_5519);
nand UO_190 (O_190,N_9389,N_7692);
nand UO_191 (O_191,N_7558,N_5829);
and UO_192 (O_192,N_5166,N_7886);
and UO_193 (O_193,N_8218,N_5896);
nor UO_194 (O_194,N_8812,N_7244);
and UO_195 (O_195,N_5531,N_5489);
nand UO_196 (O_196,N_9411,N_6387);
nor UO_197 (O_197,N_5800,N_9113);
nand UO_198 (O_198,N_5934,N_9912);
and UO_199 (O_199,N_5977,N_5959);
or UO_200 (O_200,N_6170,N_6373);
nand UO_201 (O_201,N_5374,N_6655);
and UO_202 (O_202,N_6419,N_9678);
nor UO_203 (O_203,N_5298,N_7287);
and UO_204 (O_204,N_9165,N_9211);
and UO_205 (O_205,N_7047,N_7656);
nand UO_206 (O_206,N_6803,N_8852);
or UO_207 (O_207,N_7828,N_7529);
nand UO_208 (O_208,N_6352,N_8543);
xnor UO_209 (O_209,N_6650,N_8999);
or UO_210 (O_210,N_7564,N_9048);
and UO_211 (O_211,N_9859,N_5226);
or UO_212 (O_212,N_7754,N_7936);
nand UO_213 (O_213,N_8892,N_7950);
or UO_214 (O_214,N_8019,N_9754);
or UO_215 (O_215,N_9811,N_5202);
and UO_216 (O_216,N_8735,N_7708);
nor UO_217 (O_217,N_6823,N_8231);
or UO_218 (O_218,N_9468,N_6539);
and UO_219 (O_219,N_5395,N_6317);
or UO_220 (O_220,N_9619,N_5295);
and UO_221 (O_221,N_6935,N_5082);
nor UO_222 (O_222,N_8372,N_8700);
nor UO_223 (O_223,N_6915,N_6956);
and UO_224 (O_224,N_6094,N_9464);
and UO_225 (O_225,N_7271,N_5837);
or UO_226 (O_226,N_9675,N_5867);
nand UO_227 (O_227,N_8940,N_6232);
and UO_228 (O_228,N_7836,N_6674);
or UO_229 (O_229,N_8815,N_7300);
nor UO_230 (O_230,N_6205,N_5484);
nand UO_231 (O_231,N_7850,N_5050);
and UO_232 (O_232,N_8990,N_5453);
and UO_233 (O_233,N_6761,N_7535);
nor UO_234 (O_234,N_9220,N_7470);
nand UO_235 (O_235,N_8491,N_5016);
and UO_236 (O_236,N_9809,N_7482);
or UO_237 (O_237,N_7248,N_5642);
nor UO_238 (O_238,N_9382,N_6773);
and UO_239 (O_239,N_5385,N_6484);
or UO_240 (O_240,N_5596,N_7815);
nand UO_241 (O_241,N_8754,N_7067);
nand UO_242 (O_242,N_5913,N_7514);
and UO_243 (O_243,N_5211,N_9574);
nand UO_244 (O_244,N_6883,N_6231);
or UO_245 (O_245,N_9348,N_6248);
or UO_246 (O_246,N_6355,N_5463);
and UO_247 (O_247,N_7892,N_6964);
or UO_248 (O_248,N_9784,N_9407);
and UO_249 (O_249,N_8429,N_9070);
and UO_250 (O_250,N_9555,N_7352);
nor UO_251 (O_251,N_8091,N_5749);
nor UO_252 (O_252,N_7219,N_8165);
nor UO_253 (O_253,N_8298,N_9126);
or UO_254 (O_254,N_9775,N_8620);
nor UO_255 (O_255,N_8239,N_6172);
or UO_256 (O_256,N_5505,N_9803);
nand UO_257 (O_257,N_6004,N_7978);
and UO_258 (O_258,N_7620,N_9441);
nor UO_259 (O_259,N_9131,N_6431);
nand UO_260 (O_260,N_9397,N_8124);
nand UO_261 (O_261,N_9482,N_8618);
nor UO_262 (O_262,N_6350,N_9919);
nor UO_263 (O_263,N_6051,N_8279);
and UO_264 (O_264,N_6905,N_8316);
and UO_265 (O_265,N_5071,N_5841);
nand UO_266 (O_266,N_7662,N_9891);
or UO_267 (O_267,N_6140,N_9145);
nor UO_268 (O_268,N_9989,N_9531);
nand UO_269 (O_269,N_7332,N_6755);
nor UO_270 (O_270,N_7979,N_6450);
and UO_271 (O_271,N_5601,N_6631);
nand UO_272 (O_272,N_9294,N_5785);
or UO_273 (O_273,N_5272,N_9703);
nor UO_274 (O_274,N_6724,N_6334);
nor UO_275 (O_275,N_6712,N_5863);
or UO_276 (O_276,N_5112,N_6572);
nor UO_277 (O_277,N_8778,N_6588);
xor UO_278 (O_278,N_7861,N_8234);
nor UO_279 (O_279,N_6275,N_5241);
and UO_280 (O_280,N_5008,N_8562);
and UO_281 (O_281,N_5975,N_9599);
nand UO_282 (O_282,N_7091,N_8593);
nor UO_283 (O_283,N_8862,N_5238);
and UO_284 (O_284,N_9743,N_6462);
nand UO_285 (O_285,N_9173,N_9295);
and UO_286 (O_286,N_7933,N_7723);
and UO_287 (O_287,N_8553,N_5420);
and UO_288 (O_288,N_8428,N_8743);
and UO_289 (O_289,N_6690,N_8807);
nand UO_290 (O_290,N_8822,N_5853);
and UO_291 (O_291,N_8385,N_5005);
nand UO_292 (O_292,N_6138,N_5821);
or UO_293 (O_293,N_6678,N_6955);
nand UO_294 (O_294,N_9333,N_7755);
and UO_295 (O_295,N_5587,N_7904);
and UO_296 (O_296,N_7885,N_5470);
or UO_297 (O_297,N_8447,N_9772);
nor UO_298 (O_298,N_6095,N_9605);
and UO_299 (O_299,N_7240,N_7614);
nor UO_300 (O_300,N_7851,N_5827);
nor UO_301 (O_301,N_8679,N_9536);
nand UO_302 (O_302,N_8613,N_8024);
and UO_303 (O_303,N_6296,N_6118);
or UO_304 (O_304,N_5992,N_9208);
nor UO_305 (O_305,N_5171,N_8001);
or UO_306 (O_306,N_9983,N_7198);
or UO_307 (O_307,N_5706,N_6695);
nor UO_308 (O_308,N_9630,N_7366);
nand UO_309 (O_309,N_7502,N_5261);
nand UO_310 (O_310,N_8415,N_5145);
nor UO_311 (O_311,N_6836,N_7506);
nor UO_312 (O_312,N_8064,N_7036);
or UO_313 (O_313,N_6144,N_9716);
nand UO_314 (O_314,N_6881,N_5412);
nand UO_315 (O_315,N_6046,N_8819);
xor UO_316 (O_316,N_9872,N_7425);
and UO_317 (O_317,N_8569,N_8972);
and UO_318 (O_318,N_6173,N_9284);
or UO_319 (O_319,N_7314,N_7849);
nor UO_320 (O_320,N_8387,N_5836);
nand UO_321 (O_321,N_7301,N_5986);
or UO_322 (O_322,N_8136,N_9436);
or UO_323 (O_323,N_7202,N_6852);
nor UO_324 (O_324,N_7169,N_6483);
and UO_325 (O_325,N_8360,N_6306);
and UO_326 (O_326,N_9049,N_6993);
nor UO_327 (O_327,N_5514,N_7883);
or UO_328 (O_328,N_8531,N_6839);
nand UO_329 (O_329,N_5344,N_7675);
nand UO_330 (O_330,N_9897,N_8564);
nand UO_331 (O_331,N_5328,N_6485);
and UO_332 (O_332,N_9293,N_8379);
nor UO_333 (O_333,N_7016,N_9477);
or UO_334 (O_334,N_8419,N_7684);
or UO_335 (O_335,N_9046,N_7814);
or UO_336 (O_336,N_9806,N_6177);
nor UO_337 (O_337,N_5899,N_7534);
nor UO_338 (O_338,N_6713,N_6333);
and UO_339 (O_339,N_9033,N_9904);
and UO_340 (O_340,N_7447,N_6949);
and UO_341 (O_341,N_6079,N_9620);
and UO_342 (O_342,N_6607,N_7812);
or UO_343 (O_343,N_7109,N_6403);
nor UO_344 (O_344,N_9755,N_6705);
and UO_345 (O_345,N_9082,N_6377);
nand UO_346 (O_346,N_9971,N_7421);
and UO_347 (O_347,N_5160,N_8597);
nor UO_348 (O_348,N_6771,N_6486);
and UO_349 (O_349,N_9738,N_6080);
nand UO_350 (O_350,N_5123,N_5214);
nor UO_351 (O_351,N_7676,N_8434);
nand UO_352 (O_352,N_5161,N_9075);
or UO_353 (O_353,N_7082,N_9518);
or UO_354 (O_354,N_6612,N_9857);
and UO_355 (O_355,N_6222,N_8104);
nor UO_356 (O_356,N_7365,N_9769);
nand UO_357 (O_357,N_8727,N_5560);
or UO_358 (O_358,N_6584,N_9258);
nor UO_359 (O_359,N_7090,N_8530);
nor UO_360 (O_360,N_9162,N_6656);
nor UO_361 (O_361,N_8121,N_9592);
and UO_362 (O_362,N_9926,N_7838);
and UO_363 (O_363,N_9019,N_8652);
nand UO_364 (O_364,N_8529,N_5010);
and UO_365 (O_365,N_6075,N_8690);
nor UO_366 (O_366,N_5777,N_5334);
or UO_367 (O_367,N_8045,N_7030);
and UO_368 (O_368,N_9923,N_5499);
nand UO_369 (O_369,N_6371,N_8737);
or UO_370 (O_370,N_6208,N_6101);
or UO_371 (O_371,N_8444,N_5738);
and UO_372 (O_372,N_5477,N_6608);
nor UO_373 (O_373,N_9717,N_6410);
nand UO_374 (O_374,N_8393,N_8332);
or UO_375 (O_375,N_7413,N_7013);
or UO_376 (O_376,N_5310,N_6929);
nand UO_377 (O_377,N_6860,N_7139);
nand UO_378 (O_378,N_8685,N_9103);
nand UO_379 (O_379,N_5721,N_9720);
nor UO_380 (O_380,N_7356,N_6359);
nand UO_381 (O_381,N_7613,N_5228);
or UO_382 (O_382,N_8187,N_6078);
and UO_383 (O_383,N_8965,N_7273);
nand UO_384 (O_384,N_6963,N_7749);
and UO_385 (O_385,N_8952,N_6042);
nand UO_386 (O_386,N_9190,N_6039);
and UO_387 (O_387,N_6610,N_5763);
and UO_388 (O_388,N_6420,N_7325);
nor UO_389 (O_389,N_9326,N_7419);
nor UO_390 (O_390,N_9729,N_9324);
and UO_391 (O_391,N_9451,N_7298);
nor UO_392 (O_392,N_8506,N_5403);
or UO_393 (O_393,N_6439,N_7491);
nor UO_394 (O_394,N_8845,N_8449);
nand UO_395 (O_395,N_6105,N_5901);
nand UO_396 (O_396,N_8314,N_8736);
nand UO_397 (O_397,N_7435,N_5686);
nand UO_398 (O_398,N_5375,N_7557);
nand UO_399 (O_399,N_7385,N_5609);
nand UO_400 (O_400,N_6611,N_7512);
and UO_401 (O_401,N_8896,N_6427);
and UO_402 (O_402,N_7295,N_8834);
nand UO_403 (O_403,N_9055,N_7417);
and UO_404 (O_404,N_8069,N_9080);
or UO_405 (O_405,N_5060,N_5313);
nand UO_406 (O_406,N_9948,N_6343);
nand UO_407 (O_407,N_6076,N_6808);
nor UO_408 (O_408,N_8404,N_7234);
nor UO_409 (O_409,N_7856,N_6730);
nor UO_410 (O_410,N_8311,N_9203);
nor UO_411 (O_411,N_5022,N_8070);
and UO_412 (O_412,N_5900,N_7017);
nor UO_413 (O_413,N_6970,N_9473);
or UO_414 (O_414,N_5026,N_7533);
or UO_415 (O_415,N_7480,N_9136);
nand UO_416 (O_416,N_8366,N_8937);
or UO_417 (O_417,N_5373,N_9489);
or UO_418 (O_418,N_9936,N_6805);
nand UO_419 (O_419,N_6077,N_7056);
or UO_420 (O_420,N_9645,N_8855);
xnor UO_421 (O_421,N_5217,N_9487);
and UO_422 (O_422,N_9802,N_8062);
nand UO_423 (O_423,N_8695,N_9346);
and UO_424 (O_424,N_6299,N_5653);
and UO_425 (O_425,N_7628,N_8585);
nor UO_426 (O_426,N_9016,N_7928);
or UO_427 (O_427,N_6050,N_8842);
or UO_428 (O_428,N_6374,N_9874);
or UO_429 (O_429,N_5859,N_6582);
and UO_430 (O_430,N_7397,N_5898);
and UO_431 (O_431,N_9362,N_5340);
nand UO_432 (O_432,N_7832,N_9519);
nor UO_433 (O_433,N_5890,N_7286);
and UO_434 (O_434,N_9665,N_6098);
nand UO_435 (O_435,N_8637,N_5302);
nand UO_436 (O_436,N_7426,N_7642);
or UO_437 (O_437,N_7276,N_9888);
nor UO_438 (O_438,N_8733,N_9951);
and UO_439 (O_439,N_5300,N_7083);
nor UO_440 (O_440,N_5823,N_5209);
nor UO_441 (O_441,N_7780,N_6295);
nand UO_442 (O_442,N_7536,N_6938);
nor UO_443 (O_443,N_6184,N_9292);
or UO_444 (O_444,N_5475,N_6542);
or UO_445 (O_445,N_9793,N_7768);
nand UO_446 (O_446,N_7507,N_6775);
nor UO_447 (O_447,N_6943,N_9336);
and UO_448 (O_448,N_6467,N_9522);
and UO_449 (O_449,N_5183,N_9986);
and UO_450 (O_450,N_6100,N_7953);
nor UO_451 (O_451,N_6958,N_7919);
xor UO_452 (O_452,N_8634,N_8420);
nor UO_453 (O_453,N_5154,N_8934);
nand UO_454 (O_454,N_6532,N_7415);
nand UO_455 (O_455,N_6549,N_5090);
and UO_456 (O_456,N_7974,N_6473);
nor UO_457 (O_457,N_9373,N_8836);
nor UO_458 (O_458,N_8967,N_9641);
nand UO_459 (O_459,N_7667,N_7862);
nand UO_460 (O_460,N_6507,N_8228);
and UO_461 (O_461,N_8933,N_8347);
nor UO_462 (O_462,N_9496,N_8077);
nor UO_463 (O_463,N_7672,N_7649);
and UO_464 (O_464,N_8766,N_7177);
and UO_465 (O_465,N_5447,N_6124);
nor UO_466 (O_466,N_6302,N_9540);
nor UO_467 (O_467,N_9332,N_9011);
nand UO_468 (O_468,N_5274,N_6376);
nand UO_469 (O_469,N_9866,N_6973);
or UO_470 (O_470,N_5058,N_8378);
nand UO_471 (O_471,N_8867,N_5928);
nand UO_472 (O_472,N_8839,N_6506);
nor UO_473 (O_473,N_8038,N_5521);
nand UO_474 (O_474,N_6968,N_9520);
and UO_475 (O_475,N_9862,N_5915);
and UO_476 (O_476,N_6282,N_9251);
nand UO_477 (O_477,N_7767,N_8878);
nor UO_478 (O_478,N_9791,N_6591);
or UO_479 (O_479,N_8726,N_7220);
or UO_480 (O_480,N_9943,N_7623);
and UO_481 (O_481,N_9523,N_9340);
nand UO_482 (O_482,N_5633,N_7060);
or UO_483 (O_483,N_5164,N_8900);
nand UO_484 (O_484,N_7147,N_5450);
and UO_485 (O_485,N_5709,N_7734);
and UO_486 (O_486,N_9182,N_7762);
nor UO_487 (O_487,N_5905,N_6576);
or UO_488 (O_488,N_8350,N_8021);
and UO_489 (O_489,N_8884,N_5728);
nor UO_490 (O_490,N_8795,N_5287);
nor UO_491 (O_491,N_7239,N_5619);
nand UO_492 (O_492,N_5188,N_5535);
nand UO_493 (O_493,N_9217,N_7086);
or UO_494 (O_494,N_8793,N_9179);
or UO_495 (O_495,N_5133,N_9731);
nand UO_496 (O_496,N_9349,N_9038);
or UO_497 (O_497,N_5409,N_8566);
and UO_498 (O_498,N_7010,N_9455);
and UO_499 (O_499,N_6313,N_6918);
nand UO_500 (O_500,N_8752,N_7664);
and UO_501 (O_501,N_6767,N_6939);
nor UO_502 (O_502,N_9379,N_9821);
and UO_503 (O_503,N_9202,N_7283);
nor UO_504 (O_504,N_6119,N_8876);
and UO_505 (O_505,N_5394,N_5249);
nor UO_506 (O_506,N_8528,N_6201);
nor UO_507 (O_507,N_7110,N_7921);
or UO_508 (O_508,N_7678,N_6475);
nor UO_509 (O_509,N_7377,N_7800);
nand UO_510 (O_510,N_9910,N_5074);
or UO_511 (O_511,N_7250,N_8522);
or UO_512 (O_512,N_9495,N_7445);
nand UO_513 (O_513,N_6324,N_5520);
nand UO_514 (O_514,N_5718,N_7589);
nor UO_515 (O_515,N_9141,N_9752);
or UO_516 (O_516,N_5916,N_6758);
and UO_517 (O_517,N_6395,N_9914);
or UO_518 (O_518,N_5526,N_8375);
and UO_519 (O_519,N_9045,N_8948);
or UO_520 (O_520,N_9363,N_7657);
nor UO_521 (O_521,N_8799,N_5931);
nor UO_522 (O_522,N_9558,N_5680);
and UO_523 (O_523,N_5396,N_9515);
nand UO_524 (O_524,N_8605,N_7517);
and UO_525 (O_525,N_6067,N_9861);
nor UO_526 (O_526,N_5410,N_5754);
nand UO_527 (O_527,N_8954,N_8711);
nor UO_528 (O_528,N_5246,N_9656);
nand UO_529 (O_529,N_9314,N_9993);
and UO_530 (O_530,N_5972,N_6783);
and UO_531 (O_531,N_5834,N_5077);
nand UO_532 (O_532,N_5982,N_9172);
or UO_533 (O_533,N_9008,N_5689);
nor UO_534 (O_534,N_5919,N_8040);
nor UO_535 (O_535,N_6849,N_6969);
and UO_536 (O_536,N_7376,N_8840);
or UO_537 (O_537,N_9328,N_8468);
or UO_538 (O_538,N_6472,N_5894);
nor UO_539 (O_539,N_6877,N_5494);
or UO_540 (O_540,N_6936,N_8757);
nand UO_541 (O_541,N_6072,N_5129);
or UO_542 (O_542,N_8753,N_6441);
nand UO_543 (O_543,N_9820,N_5617);
nand UO_544 (O_544,N_5762,N_9100);
and UO_545 (O_545,N_6482,N_7989);
nand UO_546 (O_546,N_5380,N_5632);
or UO_547 (O_547,N_6525,N_9123);
nand UO_548 (O_548,N_9824,N_7094);
nor UO_549 (O_549,N_6156,N_7808);
nor UO_550 (O_550,N_7947,N_9634);
or UO_551 (O_551,N_7439,N_5028);
nor UO_552 (O_552,N_9702,N_5377);
nand UO_553 (O_553,N_5885,N_5879);
nand UO_554 (O_554,N_8320,N_7538);
or UO_555 (O_555,N_7218,N_5117);
and UO_556 (O_556,N_8838,N_7607);
nand UO_557 (O_557,N_5575,N_9969);
or UO_558 (O_558,N_6848,N_9273);
nor UO_559 (O_559,N_9153,N_8864);
or UO_560 (O_560,N_7519,N_8746);
nor UO_561 (O_561,N_6278,N_6049);
nand UO_562 (O_562,N_9837,N_7677);
nor UO_563 (O_563,N_5729,N_5388);
or UO_564 (O_564,N_5068,N_7545);
nand UO_565 (O_565,N_6638,N_6202);
or UO_566 (O_566,N_5254,N_7869);
nor UO_567 (O_567,N_6738,N_9007);
or UO_568 (O_568,N_7315,N_7870);
and UO_569 (O_569,N_6727,N_9654);
nand UO_570 (O_570,N_5767,N_8744);
and UO_571 (O_571,N_8406,N_8433);
nor UO_572 (O_572,N_9689,N_5529);
nor UO_573 (O_573,N_7180,N_8782);
nand UO_574 (O_574,N_7809,N_8825);
nand UO_575 (O_575,N_6345,N_9152);
nand UO_576 (O_576,N_6762,N_5845);
nand UO_577 (O_577,N_6759,N_8523);
nor UO_578 (O_578,N_6086,N_6854);
nand UO_579 (O_579,N_7057,N_9488);
nor UO_580 (O_580,N_5849,N_9958);
and UO_581 (O_581,N_9053,N_5850);
or UO_582 (O_582,N_5359,N_5273);
and UO_583 (O_583,N_5093,N_7371);
and UO_584 (O_584,N_9167,N_7146);
nor UO_585 (O_585,N_7392,N_7145);
and UO_586 (O_586,N_5507,N_6747);
or UO_587 (O_587,N_8266,N_7996);
and UO_588 (O_588,N_9741,N_9513);
or UO_589 (O_589,N_8699,N_5487);
nand UO_590 (O_590,N_9564,N_7187);
and UO_591 (O_591,N_8490,N_9883);
or UO_592 (O_592,N_9072,N_7679);
nor UO_593 (O_593,N_7252,N_7499);
nor UO_594 (O_594,N_5270,N_8355);
nor UO_595 (O_595,N_7292,N_8424);
or UO_596 (O_596,N_5712,N_7437);
nor UO_597 (O_597,N_7835,N_8255);
nand UO_598 (O_598,N_6857,N_8565);
or UO_599 (O_599,N_6106,N_6459);
and UO_600 (O_600,N_6390,N_6633);
nor UO_601 (O_601,N_7469,N_8646);
nor UO_602 (O_602,N_5843,N_6581);
or UO_603 (O_603,N_7128,N_6432);
nand UO_604 (O_604,N_7882,N_5110);
nor UO_605 (O_605,N_9681,N_5636);
or UO_606 (O_606,N_7150,N_7964);
nor UO_607 (O_607,N_8056,N_5402);
nor UO_608 (O_608,N_6417,N_9614);
and UO_609 (O_609,N_8325,N_6752);
and UO_610 (O_610,N_7874,N_8830);
nand UO_611 (O_611,N_5251,N_5131);
nand UO_612 (O_612,N_8499,N_9937);
nor UO_613 (O_613,N_7720,N_7750);
nand UO_614 (O_614,N_9409,N_7804);
nor UO_615 (O_615,N_6634,N_9934);
nand UO_616 (O_616,N_8075,N_8321);
and UO_617 (O_617,N_5423,N_7370);
or UO_618 (O_618,N_9422,N_6155);
or UO_619 (O_619,N_8953,N_7000);
nor UO_620 (O_620,N_8771,N_8638);
or UO_621 (O_621,N_5541,N_5585);
or UO_622 (O_622,N_5549,N_6625);
and UO_623 (O_623,N_9684,N_7685);
nand UO_624 (O_624,N_6691,N_9481);
or UO_625 (O_625,N_6288,N_6602);
or UO_626 (O_626,N_5539,N_5413);
and UO_627 (O_627,N_6801,N_6799);
nand UO_628 (O_628,N_6375,N_6151);
nand UO_629 (O_629,N_9034,N_7508);
or UO_630 (O_630,N_5366,N_9938);
nor UO_631 (O_631,N_8643,N_6658);
nor UO_632 (O_632,N_6740,N_9289);
or UO_633 (O_633,N_9788,N_9071);
or UO_634 (O_634,N_6224,N_5259);
nand UO_635 (O_635,N_7647,N_5358);
or UO_636 (O_636,N_6765,N_8443);
nand UO_637 (O_637,N_5182,N_7305);
or UO_638 (O_638,N_9134,N_8402);
nor UO_639 (O_639,N_5736,N_7309);
or UO_640 (O_640,N_5153,N_8621);
and UO_641 (O_641,N_8147,N_9633);
or UO_642 (O_642,N_8511,N_6543);
and UO_643 (O_643,N_5128,N_7361);
nor UO_644 (O_644,N_6725,N_8059);
and UO_645 (O_645,N_7394,N_8536);
nor UO_646 (O_646,N_7550,N_8504);
or UO_647 (O_647,N_5156,N_5798);
and UO_648 (O_648,N_9297,N_5725);
and UO_649 (O_649,N_6340,N_8510);
and UO_650 (O_650,N_8252,N_7224);
and UO_651 (O_651,N_7826,N_9219);
nor UO_652 (O_652,N_9076,N_9920);
nand UO_653 (O_653,N_5072,N_7304);
or UO_654 (O_654,N_7232,N_7316);
nor UO_655 (O_655,N_6241,N_9427);
and UO_656 (O_656,N_8719,N_8964);
nand UO_657 (O_657,N_7383,N_9968);
or UO_658 (O_658,N_5318,N_7019);
and UO_659 (O_659,N_8268,N_8759);
and UO_660 (O_660,N_6824,N_8879);
nand UO_661 (O_661,N_7488,N_5746);
nor UO_662 (O_662,N_7940,N_8686);
xnor UO_663 (O_663,N_7207,N_6262);
xnor UO_664 (O_664,N_7777,N_5844);
nand UO_665 (O_665,N_5815,N_7127);
and UO_666 (O_666,N_7605,N_5219);
or UO_667 (O_667,N_8335,N_5355);
nand UO_668 (O_668,N_8694,N_7032);
and UO_669 (O_669,N_8903,N_8273);
and UO_670 (O_670,N_7236,N_7511);
and UO_671 (O_671,N_7446,N_6292);
nand UO_672 (O_672,N_6268,N_7050);
or UO_673 (O_673,N_6888,N_7877);
and UO_674 (O_674,N_8507,N_6835);
nor UO_675 (O_675,N_6338,N_8893);
and UO_676 (O_676,N_5778,N_7341);
nand UO_677 (O_677,N_5860,N_6425);
and UO_678 (O_678,N_8392,N_6293);
and UO_679 (O_679,N_7489,N_5176);
or UO_680 (O_680,N_5064,N_7072);
nand UO_681 (O_681,N_6195,N_9737);
nor UO_682 (O_682,N_5020,N_7063);
nor UO_683 (O_683,N_8882,N_7626);
or UO_684 (O_684,N_7441,N_8692);
nor UO_685 (O_685,N_6382,N_6815);
nor UO_686 (O_686,N_6648,N_6979);
nand UO_687 (O_687,N_9843,N_8557);
nor UO_688 (O_688,N_5664,N_6272);
nand UO_689 (O_689,N_7879,N_7690);
or UO_690 (O_690,N_5697,N_7659);
nand UO_691 (O_691,N_6697,N_6793);
nor UO_692 (O_692,N_7552,N_7624);
and UO_693 (O_693,N_7713,N_5196);
or UO_694 (O_694,N_9358,N_9125);
nand UO_695 (O_695,N_9856,N_8140);
nand UO_696 (O_696,N_9644,N_6365);
or UO_697 (O_697,N_7709,N_7631);
nand UO_698 (O_698,N_8789,N_7200);
xnor UO_699 (O_699,N_7088,N_5878);
or UO_700 (O_700,N_7797,N_6239);
nor UO_701 (O_701,N_7759,N_7806);
nor UO_702 (O_702,N_8777,N_9975);
and UO_703 (O_703,N_9988,N_5184);
or UO_704 (O_704,N_9591,N_5925);
and UO_705 (O_705,N_9079,N_7455);
nand UO_706 (O_706,N_5115,N_8917);
and UO_707 (O_707,N_6412,N_8333);
nand UO_708 (O_708,N_6448,N_6381);
nand UO_709 (O_709,N_7773,N_6197);
nor UO_710 (O_710,N_8932,N_9808);
and UO_711 (O_711,N_6781,N_8814);
nand UO_712 (O_712,N_9460,N_6550);
or UO_713 (O_713,N_6396,N_6802);
nand UO_714 (O_714,N_8391,N_9879);
and UO_715 (O_715,N_5120,N_8614);
or UO_716 (O_716,N_5125,N_9024);
or UO_717 (O_717,N_7186,N_5946);
nand UO_718 (O_718,N_7751,N_6181);
nor UO_719 (O_719,N_6782,N_6346);
nand UO_720 (O_720,N_8734,N_8439);
and UO_721 (O_721,N_5369,N_8101);
nand UO_722 (O_722,N_5051,N_8563);
nor UO_723 (O_723,N_9003,N_6788);
or UO_724 (O_724,N_5600,N_5927);
nand UO_725 (O_725,N_8797,N_8470);
or UO_726 (O_726,N_5495,N_7694);
or UO_727 (O_727,N_9525,N_5271);
or UO_728 (O_728,N_9275,N_8550);
nand UO_729 (O_729,N_5581,N_7460);
nor UO_730 (O_730,N_9554,N_9262);
and UO_731 (O_731,N_6885,N_6865);
and UO_732 (O_732,N_7172,N_5205);
or UO_733 (O_733,N_5324,N_9085);
or UO_734 (O_734,N_7427,N_7982);
nand UO_735 (O_735,N_8142,N_9476);
or UO_736 (O_736,N_7093,N_5755);
nor UO_737 (O_737,N_5109,N_6048);
nand UO_738 (O_738,N_7722,N_8790);
nor UO_739 (O_739,N_9304,N_6477);
or UO_740 (O_740,N_8192,N_5956);
nand UO_741 (O_741,N_6520,N_6356);
nor UO_742 (O_742,N_5704,N_5460);
and UO_743 (O_743,N_6772,N_5265);
or UO_744 (O_744,N_6284,N_6959);
or UO_745 (O_745,N_7687,N_8826);
nor UO_746 (O_746,N_8086,N_7209);
nand UO_747 (O_747,N_9760,N_7498);
and UO_748 (O_748,N_6983,N_8076);
nand UO_749 (O_749,N_8349,N_8642);
or UO_750 (O_750,N_5462,N_6413);
and UO_751 (O_751,N_6245,N_8714);
nand UO_752 (O_752,N_8509,N_8792);
or UO_753 (O_753,N_9444,N_9337);
nor UO_754 (O_754,N_8898,N_7700);
and UO_755 (O_755,N_8027,N_9858);
nand UO_756 (O_756,N_7420,N_5167);
nand UO_757 (O_757,N_6455,N_7142);
and UO_758 (O_758,N_8107,N_6126);
or UO_759 (O_759,N_8975,N_5311);
nand UO_760 (O_760,N_7650,N_8657);
nor UO_761 (O_761,N_5149,N_9285);
and UO_762 (O_762,N_7952,N_7245);
xor UO_763 (O_763,N_5623,N_7887);
nor UO_764 (O_764,N_7438,N_5759);
or UO_765 (O_765,N_7942,N_5857);
nand UO_766 (O_766,N_6142,N_7452);
nor UO_767 (O_767,N_7496,N_5835);
nand UO_768 (O_768,N_8633,N_9352);
and UO_769 (O_769,N_6978,N_7779);
nor UO_770 (O_770,N_9902,N_8122);
and UO_771 (O_771,N_9017,N_5748);
and UO_772 (O_772,N_5190,N_6415);
or UO_773 (O_773,N_6190,N_9051);
nor UO_774 (O_774,N_6902,N_7103);
nor UO_775 (O_775,N_9147,N_7249);
nand UO_776 (O_776,N_6213,N_5574);
nand UO_777 (O_777,N_9221,N_8644);
nor UO_778 (O_778,N_7891,N_9241);
nor UO_779 (O_779,N_9995,N_8927);
or UO_780 (O_780,N_5174,N_8946);
or UO_781 (O_781,N_5923,N_5339);
nor UO_782 (O_782,N_9090,N_9345);
or UO_783 (O_783,N_8857,N_8236);
nand UO_784 (O_784,N_8661,N_7963);
nand UO_785 (O_785,N_6774,N_5424);
or UO_786 (O_786,N_8595,N_9341);
nand UO_787 (O_787,N_6952,N_8598);
nor UO_788 (O_788,N_7571,N_8177);
or UO_789 (O_789,N_8327,N_5553);
nor UO_790 (O_790,N_6706,N_6430);
and UO_791 (O_791,N_7881,N_6113);
or UO_792 (O_792,N_8418,N_9706);
nor UO_793 (O_793,N_5895,N_9742);
nor UO_794 (O_794,N_6629,N_8768);
or UO_795 (O_795,N_7578,N_6212);
nor UO_796 (O_796,N_5244,N_8725);
nor UO_797 (O_797,N_7432,N_9484);
nand UO_798 (O_798,N_5348,N_8012);
or UO_799 (O_799,N_8035,N_5771);
nand UO_800 (O_800,N_7320,N_6675);
nor UO_801 (O_801,N_9600,N_5086);
nor UO_802 (O_802,N_6344,N_9266);
and UO_803 (O_803,N_5116,N_7844);
and UO_804 (O_804,N_6909,N_6493);
nand UO_805 (O_805,N_9226,N_5338);
nor UO_806 (O_806,N_7618,N_6897);
and UO_807 (O_807,N_9365,N_5471);
or UO_808 (O_808,N_5831,N_6397);
or UO_809 (O_809,N_6811,N_6137);
nand UO_810 (O_810,N_8494,N_7640);
nor UO_811 (O_811,N_5181,N_5625);
and UO_812 (O_812,N_8015,N_5782);
nand UO_813 (O_813,N_5935,N_8801);
and UO_814 (O_814,N_5892,N_9233);
and UO_815 (O_815,N_9181,N_5379);
nor UO_816 (O_816,N_8370,N_6930);
nand UO_817 (O_817,N_6604,N_6025);
or UO_818 (O_818,N_9299,N_8374);
nand UO_819 (O_819,N_5558,N_6107);
or UO_820 (O_820,N_8126,N_7573);
and UO_821 (O_821,N_9529,N_6103);
nand UO_822 (O_822,N_8043,N_8962);
nand UO_823 (O_823,N_7382,N_5260);
or UO_824 (O_824,N_8786,N_6027);
nand UO_825 (O_825,N_6052,N_6800);
or UO_826 (O_826,N_6874,N_9148);
or UO_827 (O_827,N_7263,N_7695);
or UO_828 (O_828,N_8591,N_7711);
nand UO_829 (O_829,N_7018,N_8205);
nand UO_830 (O_830,N_8926,N_6501);
nor UO_831 (O_831,N_5588,N_7900);
and UO_832 (O_832,N_7598,N_6822);
nand UO_833 (O_833,N_6358,N_5756);
nor UO_834 (O_834,N_8943,N_7121);
nand UO_835 (O_835,N_9705,N_9320);
nand UO_836 (O_836,N_5907,N_6872);
nand UO_837 (O_837,N_6898,N_8602);
nor UO_838 (O_838,N_9816,N_5532);
nor UO_839 (O_839,N_9551,N_9256);
nand UO_840 (O_840,N_9311,N_9492);
and UO_841 (O_841,N_8816,N_6702);
or UO_842 (O_842,N_6555,N_5920);
xnor UO_843 (O_843,N_9508,N_9255);
and UO_844 (O_844,N_9121,N_7680);
nor UO_845 (O_845,N_5803,N_8315);
nand UO_846 (O_846,N_7327,N_8508);
or UO_847 (O_847,N_8286,N_8158);
nor UO_848 (O_848,N_5152,N_6438);
nand UO_849 (O_849,N_8261,N_7453);
and UO_850 (O_850,N_7334,N_9454);
nor UO_851 (O_851,N_8334,N_7112);
nand UO_852 (O_852,N_5941,N_6779);
nand UO_853 (O_853,N_8571,N_5138);
nand UO_854 (O_854,N_6560,N_9096);
nor UO_855 (O_855,N_7463,N_5141);
and UO_856 (O_856,N_8178,N_5530);
nand UO_857 (O_857,N_9650,N_8486);
nand UO_858 (O_858,N_9418,N_9732);
or UO_859 (O_859,N_5105,N_5838);
and UO_860 (O_860,N_9018,N_5590);
nor UO_861 (O_861,N_7006,N_5737);
nand UO_862 (O_862,N_6364,N_6583);
or UO_863 (O_863,N_5603,N_5942);
nand UO_864 (O_864,N_9161,N_8740);
or UO_865 (O_865,N_6033,N_6628);
nand UO_866 (O_866,N_5897,N_8031);
or UO_867 (O_867,N_6528,N_9896);
nor UO_868 (O_868,N_6911,N_7931);
nand UO_869 (O_869,N_9099,N_7122);
and UO_870 (O_870,N_9442,N_9590);
nand UO_871 (O_871,N_8235,N_6928);
nand UO_872 (O_872,N_8251,N_8919);
or UO_873 (O_873,N_5586,N_9384);
or UO_874 (O_874,N_8594,N_5608);
or UO_875 (O_875,N_9237,N_9394);
nor UO_876 (O_876,N_9606,N_5218);
or UO_877 (O_877,N_6309,N_8253);
or UO_878 (O_878,N_6130,N_8033);
nor UO_879 (O_879,N_9061,N_6444);
nor UO_880 (O_880,N_9447,N_6065);
or UO_881 (O_881,N_5059,N_9005);
and UO_882 (O_882,N_7411,N_5990);
nor UO_883 (O_883,N_9589,N_9244);
nand UO_884 (O_884,N_5637,N_5097);
nor UO_885 (O_885,N_5312,N_5873);
nor UO_886 (O_886,N_5872,N_8345);
nand UO_887 (O_887,N_6392,N_8250);
nand UO_888 (O_888,N_5971,N_7242);
nand UO_889 (O_889,N_5910,N_6884);
and UO_890 (O_890,N_6692,N_5780);
and UO_891 (O_891,N_7213,N_6920);
nor UO_892 (O_892,N_5014,N_8951);
and UO_893 (O_893,N_8827,N_5382);
nor UO_894 (O_894,N_6720,N_9714);
nand UO_895 (O_895,N_9457,N_7661);
nand UO_896 (O_896,N_9963,N_8017);
and UO_897 (O_897,N_8272,N_8659);
nand UO_898 (O_898,N_8013,N_6174);
and UO_899 (O_899,N_7399,N_9521);
and UO_900 (O_900,N_7357,N_5877);
nor UO_901 (O_901,N_6090,N_5989);
nand UO_902 (O_902,N_7600,N_8312);
or UO_903 (O_903,N_7903,N_6249);
and UO_904 (O_904,N_8745,N_5618);
and UO_905 (O_905,N_7537,N_9159);
and UO_906 (O_906,N_7995,N_8044);
and UO_907 (O_907,N_8495,N_9327);
and UO_908 (O_908,N_5820,N_8820);
nand UO_909 (O_909,N_9370,N_5092);
or UO_910 (O_910,N_9787,N_8950);
and UO_911 (O_911,N_9693,N_7611);
or UO_912 (O_912,N_6850,N_6598);
nand UO_913 (O_913,N_7183,N_5914);
or UO_914 (O_914,N_7771,N_9351);
nand UO_915 (O_915,N_7932,N_8861);
nand UO_916 (O_916,N_6901,N_7161);
or UO_917 (O_917,N_9087,N_9566);
nor UO_918 (O_918,N_5263,N_6251);
or UO_919 (O_919,N_8606,N_5794);
and UO_920 (O_920,N_5732,N_7229);
nor UO_921 (O_921,N_6516,N_8873);
or UO_922 (O_922,N_7065,N_9376);
nand UO_923 (O_923,N_8010,N_9850);
or UO_924 (O_924,N_5887,N_9434);
and UO_925 (O_925,N_6556,N_9973);
nand UO_926 (O_926,N_6817,N_5964);
and UO_927 (O_927,N_5534,N_7189);
nor UO_928 (O_928,N_8578,N_7038);
or UO_929 (O_929,N_8144,N_9325);
nor UO_930 (O_930,N_8767,N_8899);
nand UO_931 (O_931,N_6709,N_8880);
nor UO_932 (O_932,N_9830,N_6982);
nor UO_933 (O_933,N_6117,N_5096);
nand UO_934 (O_934,N_6831,N_8991);
xnor UO_935 (O_935,N_6487,N_8860);
nor UO_936 (O_936,N_5315,N_6164);
or UO_937 (O_937,N_6665,N_6337);
nand UO_938 (O_938,N_8575,N_6421);
or UO_939 (O_939,N_7044,N_6074);
or UO_940 (O_940,N_5151,N_5528);
nor UO_941 (O_941,N_6559,N_7197);
and UO_942 (O_942,N_6192,N_6726);
nor UO_943 (O_943,N_8961,N_7264);
nor UO_944 (O_944,N_5387,N_7652);
nor UO_945 (O_945,N_8677,N_5650);
nor UO_946 (O_946,N_8201,N_7348);
and UO_947 (O_947,N_7275,N_5078);
nand UO_948 (O_948,N_8596,N_9399);
or UO_949 (O_949,N_7523,N_9786);
or UO_950 (O_950,N_7966,N_5517);
or UO_951 (O_951,N_8835,N_5589);
nand UO_952 (O_952,N_5687,N_7596);
nor UO_953 (O_953,N_6651,N_9204);
or UO_954 (O_954,N_6913,N_9347);
nand UO_955 (O_955,N_8540,N_5908);
or UO_956 (O_956,N_5702,N_7002);
nand UO_957 (O_957,N_8364,N_8541);
nand UO_958 (O_958,N_5107,N_6777);
xor UO_959 (O_959,N_5296,N_5070);
nand UO_960 (O_960,N_6587,N_9242);
and UO_961 (O_961,N_6434,N_7457);
or UO_962 (O_962,N_9403,N_8474);
nor UO_963 (O_963,N_7868,N_9412);
and UO_964 (O_964,N_7306,N_8025);
and UO_965 (O_965,N_7379,N_5200);
and UO_966 (O_966,N_8324,N_9223);
or UO_967 (O_967,N_8191,N_8220);
or UO_968 (O_968,N_7216,N_9041);
nand UO_969 (O_969,N_5790,N_6508);
and UO_970 (O_970,N_7343,N_5414);
nor UO_971 (O_971,N_5768,N_7297);
or UO_972 (O_972,N_6163,N_8996);
and UO_973 (O_973,N_5789,N_5904);
or UO_974 (O_974,N_6780,N_6906);
and UO_975 (O_975,N_6723,N_5685);
and UO_976 (O_976,N_7681,N_9063);
nor UO_977 (O_977,N_9171,N_7654);
nor UO_978 (O_978,N_9282,N_8718);
nand UO_979 (O_979,N_7465,N_5540);
or UO_980 (O_980,N_6259,N_8749);
or UO_981 (O_981,N_6136,N_5676);
nand UO_982 (O_982,N_9974,N_5572);
xor UO_983 (O_983,N_7818,N_8242);
or UO_984 (O_984,N_5478,N_9617);
nor UO_985 (O_985,N_6880,N_9359);
nor UO_986 (O_986,N_6739,N_6624);
and UO_987 (O_987,N_9170,N_7725);
nor UO_988 (O_988,N_8426,N_9069);
xnor UO_989 (O_989,N_5673,N_6303);
and UO_990 (O_990,N_7580,N_6491);
nand UO_991 (O_991,N_7390,N_9032);
nor UO_992 (O_992,N_9847,N_9908);
and UO_993 (O_993,N_8048,N_8254);
and UO_994 (O_994,N_9548,N_7311);
nor UO_995 (O_995,N_6989,N_9750);
nand UO_996 (O_996,N_8513,N_7442);
nand UO_997 (O_997,N_6402,N_5993);
nor UO_998 (O_998,N_6139,N_6260);
nand UO_999 (O_999,N_7185,N_9834);
and UO_1000 (O_1000,N_5839,N_5118);
and UO_1001 (O_1001,N_5019,N_9648);
or UO_1002 (O_1002,N_5669,N_9748);
and UO_1003 (O_1003,N_8304,N_6545);
and UO_1004 (O_1004,N_5179,N_5947);
and UO_1005 (O_1005,N_9774,N_7785);
or UO_1006 (O_1006,N_8115,N_9670);
nor UO_1007 (O_1007,N_9835,N_6404);
and UO_1008 (O_1008,N_7373,N_6593);
or UO_1009 (O_1009,N_7079,N_6096);
or UO_1010 (O_1010,N_6825,N_6289);
and UO_1011 (O_1011,N_7487,N_5258);
nand UO_1012 (O_1012,N_5286,N_8410);
and UO_1013 (O_1013,N_6647,N_9851);
nand UO_1014 (O_1014,N_5654,N_5099);
or UO_1015 (O_1015,N_9206,N_8281);
or UO_1016 (O_1016,N_6517,N_7666);
nand UO_1017 (O_1017,N_7205,N_6998);
and UO_1018 (O_1018,N_7155,N_6246);
and UO_1019 (O_1019,N_7569,N_8535);
and UO_1020 (O_1020,N_5041,N_9078);
nor UO_1021 (O_1021,N_5613,N_5569);
nor UO_1022 (O_1022,N_9882,N_9727);
nand UO_1023 (O_1023,N_8610,N_8295);
nand UO_1024 (O_1024,N_6887,N_7521);
and UO_1025 (O_1025,N_8061,N_5698);
or UO_1026 (O_1026,N_6242,N_7360);
or UO_1027 (O_1027,N_7026,N_9967);
nand UO_1028 (O_1028,N_7969,N_7075);
and UO_1029 (O_1029,N_9780,N_5716);
nand UO_1030 (O_1030,N_8200,N_8050);
nand UO_1031 (O_1031,N_7143,N_8448);
nand UO_1032 (O_1032,N_9921,N_9947);
or UO_1033 (O_1033,N_9330,N_8701);
nor UO_1034 (O_1034,N_7203,N_5978);
nand UO_1035 (O_1035,N_7329,N_6122);
nor UO_1036 (O_1036,N_6223,N_7645);
and UO_1037 (O_1037,N_5370,N_8993);
or UO_1038 (O_1038,N_7744,N_7410);
nor UO_1039 (O_1039,N_6250,N_7331);
and UO_1040 (O_1040,N_5646,N_9056);
nor UO_1041 (O_1041,N_9699,N_6161);
nand UO_1042 (O_1042,N_6380,N_5634);
or UO_1043 (O_1043,N_8803,N_9691);
and UO_1044 (O_1044,N_7549,N_9686);
or UO_1045 (O_1045,N_7733,N_6996);
nor UO_1046 (O_1046,N_9711,N_6892);
xnor UO_1047 (O_1047,N_9318,N_5955);
nor UO_1048 (O_1048,N_9192,N_6683);
nand UO_1049 (O_1049,N_7840,N_6917);
nand UO_1050 (O_1050,N_9207,N_9396);
and UO_1051 (O_1051,N_8442,N_9091);
and UO_1052 (O_1052,N_9067,N_9150);
nor UO_1053 (O_1053,N_8224,N_7369);
nand UO_1054 (O_1054,N_8832,N_8326);
nand UO_1055 (O_1055,N_6315,N_5461);
nor UO_1056 (O_1056,N_8113,N_6866);
nand UO_1057 (O_1057,N_6256,N_6503);
nor UO_1058 (O_1058,N_8313,N_6644);
nand UO_1059 (O_1059,N_7988,N_5772);
or UO_1060 (O_1060,N_8039,N_7111);
or UO_1061 (O_1061,N_6370,N_7865);
nor UO_1062 (O_1062,N_7970,N_9688);
and UO_1063 (O_1063,N_8000,N_9849);
or UO_1064 (O_1064,N_8465,N_7278);
nor UO_1065 (O_1065,N_7669,N_8527);
or UO_1066 (O_1066,N_6029,N_7290);
nor UO_1067 (O_1067,N_9291,N_6894);
and UO_1068 (O_1068,N_9885,N_6411);
and UO_1069 (O_1069,N_5501,N_7846);
nor UO_1070 (O_1070,N_5741,N_7326);
or UO_1071 (O_1071,N_6654,N_5027);
and UO_1072 (O_1072,N_7269,N_5822);
nand UO_1073 (O_1073,N_6810,N_5425);
and UO_1074 (O_1074,N_9263,N_8570);
or UO_1075 (O_1075,N_9636,N_6209);
or UO_1076 (O_1076,N_6062,N_8092);
or UO_1077 (O_1077,N_8663,N_6199);
and UO_1078 (O_1078,N_6274,N_7860);
or UO_1079 (O_1079,N_5658,N_5162);
nand UO_1080 (O_1080,N_8478,N_7459);
or UO_1081 (O_1081,N_8885,N_5733);
nor UO_1082 (O_1082,N_8063,N_6855);
or UO_1083 (O_1083,N_9386,N_9671);
or UO_1084 (O_1084,N_6418,N_6237);
and UO_1085 (O_1085,N_7393,N_6024);
or UO_1086 (O_1086,N_8060,N_8708);
nand UO_1087 (O_1087,N_8787,N_7977);
nor UO_1088 (O_1088,N_8875,N_9305);
or UO_1089 (O_1089,N_6856,N_8054);
nor UO_1090 (O_1090,N_9433,N_9163);
or UO_1091 (O_1091,N_8455,N_5726);
nand UO_1092 (O_1092,N_8118,N_5994);
nand UO_1093 (O_1093,N_6603,N_7567);
nor UO_1094 (O_1094,N_6927,N_6907);
nand UO_1095 (O_1095,N_5401,N_5158);
and UO_1096 (O_1096,N_8558,N_9997);
nor UO_1097 (O_1097,N_6362,N_5100);
or UO_1098 (O_1098,N_9749,N_8190);
nand UO_1099 (O_1099,N_6464,N_7347);
nand UO_1100 (O_1100,N_8367,N_7108);
and UO_1101 (O_1101,N_5155,N_9652);
nor UO_1102 (O_1102,N_8872,N_7575);
nand UO_1103 (O_1103,N_5215,N_9877);
nor UO_1104 (O_1104,N_8207,N_9801);
nor UO_1105 (O_1105,N_9118,N_8676);
and UO_1106 (O_1106,N_5469,N_6331);
or UO_1107 (O_1107,N_8603,N_8264);
nand UO_1108 (O_1108,N_9494,N_6154);
nor UO_1109 (O_1109,N_9031,N_6708);
nand UO_1110 (O_1110,N_7914,N_9981);
or UO_1111 (O_1111,N_7639,N_7509);
nor UO_1112 (O_1112,N_7214,N_8095);
nand UO_1113 (O_1113,N_6870,N_8662);
nor UO_1114 (O_1114,N_5468,N_9980);
nand UO_1115 (O_1115,N_6615,N_7581);
or UO_1116 (O_1116,N_7697,N_5492);
or UO_1117 (O_1117,N_7621,N_8475);
or UO_1118 (O_1118,N_9955,N_5331);
nor UO_1119 (O_1119,N_5770,N_9704);
and UO_1120 (O_1120,N_7530,N_6660);
nor UO_1121 (O_1121,N_9724,N_7848);
or UO_1122 (O_1122,N_5309,N_6985);
nand UO_1123 (O_1123,N_5033,N_5595);
nand UO_1124 (O_1124,N_7277,N_7144);
nand UO_1125 (O_1125,N_6010,N_8262);
nor UO_1126 (O_1126,N_7956,N_5802);
or UO_1127 (O_1127,N_9453,N_5953);
and UO_1128 (O_1128,N_7805,N_9458);
nand UO_1129 (O_1129,N_9709,N_7770);
nor UO_1130 (O_1130,N_9475,N_5527);
or UO_1131 (O_1131,N_6312,N_6999);
or UO_1132 (O_1132,N_5691,N_5688);
nor UO_1133 (O_1133,N_5880,N_5951);
nand UO_1134 (O_1134,N_5961,N_9015);
or UO_1135 (O_1135,N_9900,N_6861);
or UO_1136 (O_1136,N_9511,N_6736);
nor UO_1137 (O_1137,N_6252,N_8146);
and UO_1138 (O_1138,N_7584,N_7791);
or UO_1139 (O_1139,N_6645,N_8788);
or UO_1140 (O_1140,N_9653,N_5486);
nand UO_1141 (O_1141,N_7842,N_9283);
and UO_1142 (O_1142,N_7893,N_6561);
nor UO_1143 (O_1143,N_7682,N_9637);
and UO_1144 (O_1144,N_5856,N_8446);
or UO_1145 (O_1145,N_7317,N_9137);
and UO_1146 (O_1146,N_7544,N_9663);
nor UO_1147 (O_1147,N_9524,N_6923);
and UO_1148 (O_1148,N_5550,N_7821);
or UO_1149 (O_1149,N_7985,N_7671);
or UO_1150 (O_1150,N_9277,N_8968);
and UO_1151 (O_1151,N_5063,N_7745);
nand UO_1152 (O_1152,N_7951,N_6257);
nor UO_1153 (O_1153,N_6133,N_5132);
and UO_1154 (O_1154,N_5279,N_5173);
and UO_1155 (O_1155,N_9174,N_5707);
nor UO_1156 (O_1156,N_9160,N_8904);
xor UO_1157 (O_1157,N_5866,N_8483);
or UO_1158 (O_1158,N_6746,N_5046);
nor UO_1159 (O_1159,N_6446,N_9042);
nor UO_1160 (O_1160,N_9596,N_9998);
or UO_1161 (O_1161,N_7782,N_9763);
nor UO_1162 (O_1162,N_8761,N_6529);
nand UO_1163 (O_1163,N_7196,N_6019);
nor UO_1164 (O_1164,N_9216,N_7260);
nor UO_1165 (O_1165,N_5066,N_8032);
nor UO_1166 (O_1166,N_5040,N_8732);
and UO_1167 (O_1167,N_8704,N_8260);
nand UO_1168 (O_1168,N_8670,N_5087);
nand UO_1169 (O_1169,N_7461,N_6742);
nor UO_1170 (O_1170,N_5264,N_5256);
and UO_1171 (O_1171,N_7281,N_8923);
or UO_1172 (O_1172,N_9547,N_8871);
or UO_1173 (O_1173,N_6166,N_7801);
xor UO_1174 (O_1174,N_7004,N_8532);
nand UO_1175 (O_1175,N_8756,N_9790);
nor UO_1176 (O_1176,N_7284,N_8373);
and UO_1177 (O_1177,N_6165,N_6987);
nand UO_1178 (O_1178,N_9909,N_9587);
nand UO_1179 (O_1179,N_7274,N_5036);
or UO_1180 (O_1180,N_5106,N_7693);
or UO_1181 (O_1181,N_6456,N_7005);
and UO_1182 (O_1182,N_7946,N_6069);
and UO_1183 (O_1183,N_6526,N_5474);
nor UO_1184 (O_1184,N_9533,N_5007);
or UO_1185 (O_1185,N_5038,N_7665);
or UO_1186 (O_1186,N_8715,N_8395);
nor UO_1187 (O_1187,N_7163,N_5441);
nand UO_1188 (O_1188,N_7440,N_8219);
and UO_1189 (O_1189,N_6329,N_7939);
and UO_1190 (O_1190,N_6182,N_5577);
nor UO_1191 (O_1191,N_7730,N_9097);
or UO_1192 (O_1192,N_7475,N_6300);
and UO_1193 (O_1193,N_7689,N_6123);
nand UO_1194 (O_1194,N_6662,N_6342);
and UO_1195 (O_1195,N_5605,N_5893);
and UO_1196 (O_1196,N_9960,N_7052);
nand UO_1197 (O_1197,N_9158,N_8229);
and UO_1198 (O_1198,N_8287,N_8539);
or UO_1199 (O_1199,N_6215,N_6469);
and UO_1200 (O_1200,N_6931,N_5057);
or UO_1201 (O_1201,N_9826,N_5288);
nor UO_1202 (O_1202,N_9339,N_5000);
and UO_1203 (O_1203,N_8421,N_7924);
nand UO_1204 (O_1204,N_7402,N_5052);
or UO_1205 (O_1205,N_8702,N_5954);
nor UO_1206 (O_1206,N_7820,N_9057);
and UO_1207 (O_1207,N_8083,N_9871);
or UO_1208 (O_1208,N_7888,N_6183);
and UO_1209 (O_1209,N_7582,N_7595);
or UO_1210 (O_1210,N_6703,N_6841);
nand UO_1211 (O_1211,N_5868,N_7637);
and UO_1212 (O_1212,N_5127,N_9264);
and UO_1213 (O_1213,N_5564,N_5142);
nor UO_1214 (O_1214,N_8805,N_9674);
nor UO_1215 (O_1215,N_9323,N_8987);
or UO_1216 (O_1216,N_9733,N_7592);
nor UO_1217 (O_1217,N_5347,N_9942);
nor UO_1218 (O_1218,N_5150,N_5360);
and UO_1219 (O_1219,N_5979,N_8212);
or UO_1220 (O_1220,N_9416,N_5056);
and UO_1221 (O_1221,N_5628,N_9154);
nor UO_1222 (O_1222,N_9361,N_9679);
or UO_1223 (O_1223,N_7707,N_6230);
nand UO_1224 (O_1224,N_7524,N_5760);
or UO_1225 (O_1225,N_8887,N_9956);
nand UO_1226 (O_1226,N_7627,N_7518);
and UO_1227 (O_1227,N_8982,N_8341);
nor UO_1228 (O_1228,N_8456,N_8105);
nor UO_1229 (O_1229,N_9854,N_7522);
and UO_1230 (O_1230,N_7045,N_8303);
or UO_1231 (O_1231,N_7253,N_8907);
nand UO_1232 (O_1232,N_8716,N_5743);
nor UO_1233 (O_1233,N_9746,N_5349);
and UO_1234 (O_1234,N_5516,N_5444);
or UO_1235 (O_1235,N_6926,N_6940);
nand UO_1236 (O_1236,N_7909,N_8616);
nor UO_1237 (O_1237,N_7551,N_7975);
or UO_1238 (O_1238,N_5891,N_8748);
nand UO_1239 (O_1239,N_8302,N_7617);
nor UO_1240 (O_1240,N_9037,N_7078);
or UO_1241 (O_1241,N_6053,N_5957);
and UO_1242 (O_1242,N_7910,N_9498);
nor UO_1243 (O_1243,N_8071,N_7456);
or UO_1244 (O_1244,N_5391,N_7610);
or UO_1245 (O_1245,N_6748,N_6068);
or UO_1246 (O_1246,N_7825,N_9805);
or UO_1247 (O_1247,N_5796,N_8057);
nand UO_1248 (O_1248,N_9507,N_5675);
and UO_1249 (O_1249,N_8034,N_5543);
or UO_1250 (O_1250,N_5952,N_9270);
or UO_1251 (O_1251,N_9846,N_7495);
and UO_1252 (O_1252,N_9542,N_9064);
nor UO_1253 (O_1253,N_5917,N_5278);
or UO_1254 (O_1254,N_6125,N_8100);
nand UO_1255 (O_1255,N_8340,N_7493);
nor UO_1256 (O_1256,N_9894,N_9610);
nor UO_1257 (O_1257,N_6636,N_6451);
nand UO_1258 (O_1258,N_5464,N_8283);
nor UO_1259 (O_1259,N_9887,N_6045);
or UO_1260 (O_1260,N_8300,N_6667);
xnor UO_1261 (O_1261,N_6523,N_8072);
or UO_1262 (O_1262,N_9585,N_6814);
nor UO_1263 (O_1263,N_5735,N_7895);
nor UO_1264 (O_1264,N_5883,N_5713);
nand UO_1265 (O_1265,N_5307,N_5294);
xor UO_1266 (O_1266,N_7070,N_5807);
nand UO_1267 (O_1267,N_7051,N_8182);
and UO_1268 (O_1268,N_5616,N_6040);
or UO_1269 (O_1269,N_7227,N_7829);
nand UO_1270 (O_1270,N_9360,N_6882);
and UO_1271 (O_1271,N_7098,N_5630);
or UO_1272 (O_1272,N_5497,N_7954);
or UO_1273 (O_1273,N_7221,N_9825);
nand UO_1274 (O_1274,N_9106,N_8626);
nor UO_1275 (O_1275,N_9354,N_5336);
and UO_1276 (O_1276,N_7201,N_5362);
nand UO_1277 (O_1277,N_6965,N_7193);
and UO_1278 (O_1278,N_5417,N_5137);
or UO_1279 (O_1279,N_5734,N_8780);
or UO_1280 (O_1280,N_6693,N_8818);
and UO_1281 (O_1281,N_7466,N_7863);
or UO_1282 (O_1282,N_8197,N_6891);
or UO_1283 (O_1283,N_7778,N_8713);
and UO_1284 (O_1284,N_8844,N_8011);
and UO_1285 (O_1285,N_7076,N_9329);
nand UO_1286 (O_1286,N_7927,N_9661);
nor UO_1287 (O_1287,N_5882,N_9905);
nand UO_1288 (O_1288,N_5788,N_9449);
nor UO_1289 (O_1289,N_5945,N_7599);
or UO_1290 (O_1290,N_7401,N_9701);
nand UO_1291 (O_1291,N_7429,N_8774);
and UO_1292 (O_1292,N_7328,N_8518);
and UO_1293 (O_1293,N_9764,N_6176);
or UO_1294 (O_1294,N_9440,N_8587);
nand UO_1295 (O_1295,N_9907,N_7175);
nand UO_1296 (O_1296,N_6732,N_8773);
nand UO_1297 (O_1297,N_9300,N_5045);
nand UO_1298 (O_1298,N_7724,N_8170);
and UO_1299 (O_1299,N_9651,N_8480);
or UO_1300 (O_1300,N_7182,N_6460);
or UO_1301 (O_1301,N_9840,N_8188);
nor UO_1302 (O_1302,N_5299,N_9575);
and UO_1303 (O_1303,N_9999,N_8318);
nor UO_1304 (O_1304,N_7294,N_8706);
or UO_1305 (O_1305,N_6807,N_5135);
or UO_1306 (O_1306,N_8471,N_7062);
or UO_1307 (O_1307,N_5177,N_9267);
nor UO_1308 (O_1308,N_7813,N_7404);
or UO_1309 (O_1309,N_8971,N_6186);
nor UO_1310 (O_1310,N_7338,N_5985);
and UO_1311 (O_1311,N_9538,N_5795);
or UO_1312 (O_1312,N_6443,N_8831);
nand UO_1313 (O_1313,N_7739,N_6637);
nand UO_1314 (O_1314,N_5371,N_5384);
and UO_1315 (O_1315,N_7961,N_8305);
nand UO_1316 (O_1316,N_5055,N_8970);
nor UO_1317 (O_1317,N_6893,N_5165);
and UO_1318 (O_1318,N_5399,N_8436);
and UO_1319 (O_1319,N_5912,N_6924);
nor UO_1320 (O_1320,N_8829,N_8775);
nand UO_1321 (O_1321,N_9715,N_8625);
nand UO_1322 (O_1322,N_6868,N_9259);
nor UO_1323 (O_1323,N_9696,N_6369);
nand UO_1324 (O_1324,N_5234,N_9356);
or UO_1325 (O_1325,N_5926,N_8109);
nor UO_1326 (O_1326,N_5742,N_6700);
nand UO_1327 (O_1327,N_5283,N_7683);
or UO_1328 (O_1328,N_6031,N_6766);
and UO_1329 (O_1329,N_7096,N_7500);
and UO_1330 (O_1330,N_7984,N_5752);
or UO_1331 (O_1331,N_8680,N_9101);
nor UO_1332 (O_1332,N_7313,N_6514);
nand UO_1333 (O_1333,N_9766,N_7412);
or UO_1334 (O_1334,N_9884,N_5053);
or UO_1335 (O_1335,N_9687,N_9274);
and UO_1336 (O_1336,N_7758,N_5024);
nand UO_1337 (O_1337,N_5198,N_5523);
nand UO_1338 (O_1338,N_8886,N_8974);
nor UO_1339 (O_1339,N_5075,N_8361);
and UO_1340 (O_1340,N_6626,N_8269);
and UO_1341 (O_1341,N_7020,N_5237);
or UO_1342 (O_1342,N_7878,N_7706);
nand UO_1343 (O_1343,N_9526,N_6643);
nand UO_1344 (O_1344,N_8883,N_8194);
and UO_1345 (O_1345,N_6057,N_6980);
or UO_1346 (O_1346,N_8084,N_7034);
or UO_1347 (O_1347,N_8342,N_8310);
nand UO_1348 (O_1348,N_7138,N_8588);
and UO_1349 (O_1349,N_7179,N_5865);
nand UO_1350 (O_1350,N_7884,N_9095);
and UO_1351 (O_1351,N_5597,N_9343);
and UO_1352 (O_1352,N_6332,N_7591);
nor UO_1353 (O_1353,N_7391,N_8055);
and UO_1354 (O_1354,N_5175,N_9039);
nand UO_1355 (O_1355,N_8400,N_5363);
or UO_1356 (O_1356,N_7210,N_8028);
and UO_1357 (O_1357,N_5536,N_6567);
xnor UO_1358 (O_1358,N_7462,N_8542);
or UO_1359 (O_1359,N_5779,N_6552);
nand UO_1360 (O_1360,N_7212,N_9010);
or UO_1361 (O_1361,N_9839,N_7434);
nor UO_1362 (O_1362,N_9429,N_6185);
nand UO_1363 (O_1363,N_9212,N_5242);
or UO_1364 (O_1364,N_9534,N_7593);
and UO_1365 (O_1365,N_8658,N_9669);
nor UO_1366 (O_1366,N_8517,N_7159);
nor UO_1367 (O_1367,N_5513,N_6680);
nand UO_1368 (O_1368,N_9378,N_5091);
xnor UO_1369 (O_1369,N_7428,N_5722);
and UO_1370 (O_1370,N_8106,N_7876);
and UO_1371 (O_1371,N_6089,N_7937);
nand UO_1372 (O_1372,N_7450,N_6325);
nand UO_1373 (O_1373,N_9426,N_8278);
nand UO_1374 (O_1374,N_5269,N_6204);
and UO_1375 (O_1375,N_9257,N_5562);
nor UO_1376 (O_1376,N_5806,N_6809);
nand UO_1377 (O_1377,N_7319,N_5751);
or UO_1378 (O_1378,N_5253,N_8184);
and UO_1379 (O_1379,N_7644,N_9470);
and UO_1380 (O_1380,N_7494,N_9209);
or UO_1381 (O_1381,N_5967,N_6150);
or UO_1382 (O_1382,N_6210,N_9954);
nor UO_1383 (O_1383,N_8487,N_8275);
and UO_1384 (O_1384,N_9252,N_7866);
and UO_1385 (O_1385,N_6844,N_5694);
and UO_1386 (O_1386,N_8849,N_8466);
or UO_1387 (O_1387,N_5938,N_9799);
nor UO_1388 (O_1388,N_5076,N_9104);
and UO_1389 (O_1389,N_8739,N_5466);
nor UO_1390 (O_1390,N_6435,N_7532);
or UO_1391 (O_1391,N_9246,N_7089);
and UO_1392 (O_1392,N_5224,N_9210);
xor UO_1393 (O_1393,N_5570,N_6326);
nand UO_1394 (O_1394,N_5906,N_5551);
nor UO_1395 (O_1395,N_5791,N_7117);
or UO_1396 (O_1396,N_9164,N_8721);
nor UO_1397 (O_1397,N_8181,N_9201);
and UO_1398 (O_1398,N_7258,N_5833);
or UO_1399 (O_1399,N_7748,N_7431);
nor UO_1400 (O_1400,N_6828,N_5515);
or UO_1401 (O_1401,N_6580,N_8233);
and UO_1402 (O_1402,N_9030,N_7737);
and UO_1403 (O_1403,N_8905,N_6933);
or UO_1404 (O_1404,N_8267,N_7520);
nand UO_1405 (O_1405,N_6562,N_9828);
and UO_1406 (O_1406,N_9377,N_6422);
nor UO_1407 (O_1407,N_7238,N_8074);
or UO_1408 (O_1408,N_5871,N_6673);
or UO_1409 (O_1409,N_8102,N_9419);
and UO_1410 (O_1410,N_5436,N_7616);
or UO_1411 (O_1411,N_5537,N_9903);
or UO_1412 (O_1412,N_9243,N_8492);
nand UO_1413 (O_1413,N_8263,N_7472);
or UO_1414 (O_1414,N_7894,N_7880);
and UO_1415 (O_1415,N_5319,N_8722);
nand UO_1416 (O_1416,N_8453,N_5591);
nor UO_1417 (O_1417,N_6499,N_5243);
or UO_1418 (O_1418,N_6007,N_9559);
nand UO_1419 (O_1419,N_9757,N_8238);
and UO_1420 (O_1420,N_9088,N_6696);
nand UO_1421 (O_1421,N_7763,N_9941);
nor UO_1422 (O_1422,N_7126,N_5604);
or UO_1423 (O_1423,N_8985,N_6478);
or UO_1424 (O_1424,N_7418,N_7560);
or UO_1425 (O_1425,N_5415,N_5607);
nand UO_1426 (O_1426,N_9086,N_9611);
nor UO_1427 (O_1427,N_8023,N_5262);
nand UO_1428 (O_1428,N_8501,N_9500);
or UO_1429 (O_1429,N_8546,N_8450);
and UO_1430 (O_1430,N_8258,N_5206);
or UO_1431 (O_1431,N_7323,N_6889);
nand UO_1432 (O_1432,N_5974,N_6769);
and UO_1433 (O_1433,N_9962,N_8270);
nand UO_1434 (O_1434,N_5949,N_6718);
nor UO_1435 (O_1435,N_7158,N_6524);
or UO_1436 (O_1436,N_8005,N_5017);
nand UO_1437 (O_1437,N_8665,N_9556);
or UO_1438 (O_1438,N_6530,N_6058);
or UO_1439 (O_1439,N_7816,N_6504);
and UO_1440 (O_1440,N_6914,N_7170);
or UO_1441 (O_1441,N_5434,N_5643);
and UO_1442 (O_1442,N_7674,N_7291);
nor UO_1443 (O_1443,N_6169,N_8847);
or UO_1444 (O_1444,N_7254,N_9338);
or UO_1445 (O_1445,N_7699,N_6819);
or UO_1446 (O_1446,N_8274,N_5073);
and UO_1447 (O_1447,N_6391,N_6820);
or UO_1448 (O_1448,N_6668,N_7873);
nor UO_1449 (O_1449,N_5612,N_5740);
nand UO_1450 (O_1450,N_8171,N_9271);
and UO_1451 (O_1451,N_7064,N_5508);
and UO_1452 (O_1452,N_5459,N_9759);
or UO_1453 (O_1453,N_6471,N_6235);
nand UO_1454 (O_1454,N_7024,N_5438);
and UO_1455 (O_1455,N_6167,N_5476);
and UO_1456 (O_1456,N_6035,N_6280);
nor UO_1457 (O_1457,N_8460,N_8346);
and UO_1458 (O_1458,N_9505,N_8798);
and UO_1459 (O_1459,N_8895,N_8167);
nand UO_1460 (O_1460,N_7351,N_9443);
and UO_1461 (O_1461,N_6757,N_6203);
or UO_1462 (O_1462,N_9994,N_9657);
or UO_1463 (O_1463,N_8560,N_7854);
nand UO_1464 (O_1464,N_8337,N_8888);
nand UO_1465 (O_1465,N_7602,N_6778);
or UO_1466 (O_1466,N_7468,N_8359);
or UO_1467 (O_1467,N_6088,N_7742);
nand UO_1468 (O_1468,N_6606,N_8691);
nand UO_1469 (O_1469,N_5252,N_8493);
and UO_1470 (O_1470,N_5185,N_8206);
or UO_1471 (O_1471,N_5048,N_7346);
or UO_1472 (O_1472,N_7228,N_7436);
nor UO_1473 (O_1473,N_6565,N_5888);
nand UO_1474 (O_1474,N_7014,N_7406);
and UO_1475 (O_1475,N_5503,N_8244);
nor UO_1476 (O_1476,N_7890,N_8123);
or UO_1477 (O_1477,N_6495,N_5457);
nand UO_1478 (O_1478,N_6108,N_5884);
or UO_1479 (O_1479,N_6960,N_5862);
or UO_1480 (O_1480,N_9301,N_9248);
nor UO_1481 (O_1481,N_7594,N_9553);
nand UO_1482 (O_1482,N_9875,N_5997);
nor UO_1483 (O_1483,N_6694,N_9726);
or UO_1484 (O_1484,N_8696,N_9116);
or UO_1485 (O_1485,N_8707,N_6474);
nor UO_1486 (O_1486,N_6254,N_7307);
nor UO_1487 (O_1487,N_5980,N_7980);
xor UO_1488 (O_1488,N_6497,N_9013);
and UO_1489 (O_1489,N_7852,N_6022);
nand UO_1490 (O_1490,N_8552,N_7349);
nor UO_1491 (O_1491,N_9719,N_7795);
nor UO_1492 (O_1492,N_9667,N_5792);
and UO_1493 (O_1493,N_7853,N_9767);
or UO_1494 (O_1494,N_9949,N_8132);
nor UO_1495 (O_1495,N_8584,N_9965);
and UO_1496 (O_1496,N_9646,N_8869);
nor UO_1497 (O_1497,N_6619,N_6341);
nor UO_1498 (O_1498,N_9119,N_8472);
nor UO_1499 (O_1499,N_6578,N_8417);
endmodule