module basic_750_5000_1000_5_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nor U0 (N_0,In_57,In_374);
nand U1 (N_1,In_289,In_120);
and U2 (N_2,In_128,In_108);
nand U3 (N_3,In_551,In_574);
nor U4 (N_4,In_645,In_256);
nor U5 (N_5,In_548,In_745);
xnor U6 (N_6,In_169,In_598);
or U7 (N_7,In_36,In_64);
nand U8 (N_8,In_189,In_436);
and U9 (N_9,In_718,In_504);
or U10 (N_10,In_243,In_335);
nor U11 (N_11,In_382,In_121);
nor U12 (N_12,In_300,In_539);
nand U13 (N_13,In_449,In_587);
nand U14 (N_14,In_650,In_725);
nand U15 (N_15,In_403,In_80);
xor U16 (N_16,In_383,In_495);
nor U17 (N_17,In_547,In_63);
and U18 (N_18,In_558,In_740);
xnor U19 (N_19,In_688,In_59);
nand U20 (N_20,In_507,In_174);
and U21 (N_21,In_171,In_513);
and U22 (N_22,In_224,In_451);
and U23 (N_23,In_514,In_331);
xor U24 (N_24,In_311,In_32);
or U25 (N_25,In_409,In_392);
and U26 (N_26,In_413,In_143);
or U27 (N_27,In_453,In_590);
xnor U28 (N_28,In_86,In_31);
xnor U29 (N_29,In_434,In_417);
nand U30 (N_30,In_217,In_597);
nand U31 (N_31,In_540,In_589);
xnor U32 (N_32,In_167,In_466);
and U33 (N_33,In_103,In_237);
or U34 (N_34,In_160,In_441);
and U35 (N_35,In_663,In_435);
nand U36 (N_36,In_502,In_527);
xnor U37 (N_37,In_588,In_673);
and U38 (N_38,In_235,In_329);
and U39 (N_39,In_135,In_90);
nand U40 (N_40,In_675,In_586);
nand U41 (N_41,In_117,In_584);
xnor U42 (N_42,In_198,In_68);
or U43 (N_43,In_608,In_572);
or U44 (N_44,In_689,In_708);
nand U45 (N_45,In_272,In_467);
xor U46 (N_46,In_294,In_488);
xor U47 (N_47,In_376,In_313);
and U48 (N_48,In_686,In_385);
nor U49 (N_49,In_278,In_369);
nand U50 (N_50,In_429,In_210);
nor U51 (N_51,In_620,In_398);
and U52 (N_52,In_671,In_119);
nand U53 (N_53,In_552,In_746);
and U54 (N_54,In_430,In_685);
and U55 (N_55,In_79,In_297);
nor U56 (N_56,In_270,In_405);
nand U57 (N_57,In_88,In_11);
nand U58 (N_58,In_260,In_643);
and U59 (N_59,In_394,In_658);
or U60 (N_60,In_332,In_164);
nand U61 (N_61,In_646,In_660);
and U62 (N_62,In_125,In_105);
or U63 (N_63,In_357,In_697);
xor U64 (N_64,In_437,In_498);
or U65 (N_65,In_720,In_264);
nand U66 (N_66,In_209,In_271);
or U67 (N_67,In_98,In_230);
nand U68 (N_68,In_499,In_211);
nand U69 (N_69,In_265,In_705);
nor U70 (N_70,In_95,In_529);
xnor U71 (N_71,In_338,In_74);
xor U72 (N_72,In_472,In_606);
nor U73 (N_73,In_622,In_581);
or U74 (N_74,In_518,In_291);
nand U75 (N_75,In_418,In_460);
nor U76 (N_76,In_13,In_516);
xnor U77 (N_77,In_431,In_35);
and U78 (N_78,In_456,In_591);
xor U79 (N_79,In_533,In_503);
or U80 (N_80,In_474,In_344);
xor U81 (N_81,In_468,In_323);
nand U82 (N_82,In_139,In_531);
nor U83 (N_83,In_293,In_333);
nor U84 (N_84,In_25,In_185);
nand U85 (N_85,In_423,In_215);
nand U86 (N_86,In_681,In_568);
nand U87 (N_87,In_562,In_47);
nor U88 (N_88,In_316,In_604);
nand U89 (N_89,In_384,In_223);
xor U90 (N_90,In_303,In_616);
xor U91 (N_91,In_283,In_302);
nor U92 (N_92,In_480,In_690);
nor U93 (N_93,In_360,In_255);
and U94 (N_94,In_582,In_266);
and U95 (N_95,In_583,In_627);
nand U96 (N_96,In_678,In_595);
nor U97 (N_97,In_107,In_654);
nand U98 (N_98,In_359,In_680);
nand U99 (N_99,In_182,In_482);
nor U100 (N_100,In_530,In_142);
nor U101 (N_101,In_393,In_132);
nor U102 (N_102,In_258,In_555);
or U103 (N_103,In_236,In_487);
nor U104 (N_104,In_240,In_82);
nand U105 (N_105,In_306,In_150);
xor U106 (N_106,In_375,In_228);
xnor U107 (N_107,In_284,In_470);
xor U108 (N_108,In_29,In_118);
nor U109 (N_109,In_162,In_477);
or U110 (N_110,In_613,In_484);
nand U111 (N_111,In_734,In_286);
nand U112 (N_112,In_700,In_567);
and U113 (N_113,In_231,In_173);
nor U114 (N_114,In_483,In_501);
or U115 (N_115,In_250,In_263);
xor U116 (N_116,In_3,In_137);
or U117 (N_117,In_239,In_199);
xnor U118 (N_118,In_695,In_87);
or U119 (N_119,In_140,In_546);
nand U120 (N_120,In_556,In_717);
xnor U121 (N_121,In_448,In_43);
or U122 (N_122,In_402,In_455);
or U123 (N_123,In_274,In_148);
nand U124 (N_124,In_349,In_577);
or U125 (N_125,In_330,In_261);
xnor U126 (N_126,In_309,In_112);
nand U127 (N_127,In_412,In_519);
nand U128 (N_128,In_78,In_386);
xor U129 (N_129,In_42,In_600);
and U130 (N_130,In_351,In_92);
nand U131 (N_131,In_565,In_337);
nand U132 (N_132,In_341,In_522);
or U133 (N_133,In_670,In_226);
or U134 (N_134,In_75,In_447);
nand U135 (N_135,In_644,In_355);
and U136 (N_136,In_267,In_299);
or U137 (N_137,In_15,In_296);
nor U138 (N_138,In_542,In_242);
and U139 (N_139,In_244,In_268);
or U140 (N_140,In_102,In_561);
nor U141 (N_141,In_679,In_343);
or U142 (N_142,In_181,In_677);
xnor U143 (N_143,In_67,In_462);
nand U144 (N_144,In_599,In_742);
nor U145 (N_145,In_94,In_634);
nor U146 (N_146,In_439,In_326);
nor U147 (N_147,In_560,In_44);
or U148 (N_148,In_629,In_636);
or U149 (N_149,In_592,In_668);
or U150 (N_150,In_141,In_69);
xor U151 (N_151,In_649,In_563);
and U152 (N_152,In_41,In_486);
and U153 (N_153,In_307,In_14);
or U154 (N_154,In_706,In_640);
xor U155 (N_155,In_346,In_505);
or U156 (N_156,In_106,In_364);
xnor U157 (N_157,In_535,In_459);
nand U158 (N_158,In_334,In_372);
and U159 (N_159,In_452,In_471);
xnor U160 (N_160,In_183,In_17);
nor U161 (N_161,In_152,In_731);
or U162 (N_162,In_692,In_191);
nor U163 (N_163,In_73,In_596);
xor U164 (N_164,In_353,In_659);
nor U165 (N_165,In_401,In_342);
nor U166 (N_166,In_515,In_602);
xnor U167 (N_167,In_373,In_218);
and U168 (N_168,In_221,In_469);
and U169 (N_169,In_525,In_425);
xor U170 (N_170,In_485,In_411);
nor U171 (N_171,In_40,In_532);
nor U172 (N_172,In_524,In_0);
nand U173 (N_173,In_238,In_179);
or U174 (N_174,In_53,In_348);
xnor U175 (N_175,In_509,In_497);
and U176 (N_176,In_396,In_716);
nand U177 (N_177,In_5,In_65);
xnor U178 (N_178,In_192,In_736);
xor U179 (N_179,In_26,In_553);
xor U180 (N_180,In_155,In_20);
nor U181 (N_181,In_696,In_245);
or U182 (N_182,In_664,In_214);
xnor U183 (N_183,In_726,In_83);
or U184 (N_184,In_336,In_698);
xnor U185 (N_185,In_433,In_631);
xnor U186 (N_186,In_156,In_728);
and U187 (N_187,In_633,In_197);
and U188 (N_188,In_724,In_637);
and U189 (N_189,In_432,In_166);
and U190 (N_190,In_420,In_168);
or U191 (N_191,In_395,In_543);
nor U192 (N_192,In_8,In_149);
or U193 (N_193,In_269,In_730);
xnor U194 (N_194,In_715,In_76);
or U195 (N_195,In_450,In_699);
nor U196 (N_196,In_279,In_234);
xnor U197 (N_197,In_314,In_207);
nor U198 (N_198,In_632,In_512);
nor U199 (N_199,In_573,In_30);
xor U200 (N_200,In_557,In_22);
or U201 (N_201,In_665,In_248);
and U202 (N_202,In_259,In_356);
nor U203 (N_203,In_612,In_446);
and U204 (N_204,In_414,In_693);
or U205 (N_205,In_661,In_415);
and U206 (N_206,In_749,In_281);
or U207 (N_207,In_609,In_319);
or U208 (N_208,In_380,In_400);
or U209 (N_209,In_157,In_454);
nand U210 (N_210,In_172,In_554);
xor U211 (N_211,In_287,In_714);
nor U212 (N_212,In_111,In_408);
or U213 (N_213,In_427,In_290);
and U214 (N_214,In_615,In_370);
nor U215 (N_215,In_748,In_571);
nand U216 (N_216,In_365,In_397);
nand U217 (N_217,In_492,In_147);
and U218 (N_218,In_196,In_362);
nor U219 (N_219,In_711,In_12);
or U220 (N_220,In_672,In_301);
nor U221 (N_221,In_225,In_144);
and U222 (N_222,In_479,In_352);
and U223 (N_223,In_647,In_491);
nor U224 (N_224,In_619,In_276);
nand U225 (N_225,In_37,In_23);
xnor U226 (N_226,In_461,In_445);
nand U227 (N_227,In_428,In_4);
nor U228 (N_228,In_626,In_607);
nor U229 (N_229,In_361,In_703);
nor U230 (N_230,In_324,In_579);
nor U231 (N_231,In_438,In_426);
xnor U232 (N_232,In_146,In_617);
nor U233 (N_233,In_123,In_521);
nand U234 (N_234,In_623,In_457);
xnor U235 (N_235,In_721,In_131);
and U236 (N_236,In_478,In_494);
or U237 (N_237,In_594,In_101);
nor U238 (N_238,In_404,In_97);
nand U239 (N_239,In_545,In_158);
nand U240 (N_240,In_463,In_292);
xor U241 (N_241,In_136,In_58);
nand U242 (N_242,In_202,In_630);
or U243 (N_243,In_683,In_241);
xor U244 (N_244,In_378,In_130);
xnor U245 (N_245,In_339,In_687);
and U246 (N_246,In_684,In_126);
nor U247 (N_247,In_628,In_305);
or U248 (N_248,In_249,In_735);
nor U249 (N_249,In_739,In_614);
or U250 (N_250,In_419,In_641);
nor U251 (N_251,In_744,In_399);
or U252 (N_252,In_710,In_246);
xnor U253 (N_253,In_662,In_325);
nor U254 (N_254,In_89,In_618);
and U255 (N_255,In_318,In_712);
xor U256 (N_256,In_388,In_345);
nor U257 (N_257,In_70,In_421);
nor U258 (N_258,In_251,In_327);
nand U259 (N_259,In_46,In_322);
xnor U260 (N_260,In_190,In_741);
nor U261 (N_261,In_85,In_50);
or U262 (N_262,In_213,In_737);
and U263 (N_263,In_151,In_180);
nand U264 (N_264,In_526,In_458);
nor U265 (N_265,In_549,In_10);
xnor U266 (N_266,In_187,In_115);
or U267 (N_267,In_253,In_216);
xor U268 (N_268,In_298,In_377);
nand U269 (N_269,In_71,In_277);
or U270 (N_270,In_18,In_55);
and U271 (N_271,In_667,In_537);
xor U272 (N_272,In_391,In_295);
xnor U273 (N_273,In_328,In_27);
or U274 (N_274,In_367,In_91);
or U275 (N_275,In_177,In_593);
and U276 (N_276,In_340,In_416);
nor U277 (N_277,In_77,In_363);
nand U278 (N_278,In_489,In_127);
nor U279 (N_279,In_475,In_350);
or U280 (N_280,In_347,In_273);
or U281 (N_281,In_16,In_159);
nor U282 (N_282,In_9,In_45);
nand U283 (N_283,In_676,In_536);
or U284 (N_284,In_729,In_138);
xor U285 (N_285,In_444,In_576);
xor U286 (N_286,In_575,In_114);
xnor U287 (N_287,In_368,In_694);
nor U288 (N_288,In_496,In_288);
and U289 (N_289,In_387,In_406);
or U290 (N_290,In_635,In_702);
xnor U291 (N_291,In_733,In_280);
nand U292 (N_292,In_262,In_56);
or U293 (N_293,In_204,In_490);
xnor U294 (N_294,In_66,In_61);
xor U295 (N_295,In_358,In_222);
nor U296 (N_296,In_569,In_390);
xor U297 (N_297,In_194,In_176);
nand U298 (N_298,In_219,In_603);
xnor U299 (N_299,In_638,In_282);
nand U300 (N_300,In_691,In_232);
and U301 (N_301,In_550,In_113);
nand U302 (N_302,In_621,In_585);
nand U303 (N_303,In_648,In_100);
nand U304 (N_304,In_578,In_682);
nor U305 (N_305,In_674,In_7);
nor U306 (N_306,In_559,In_354);
or U307 (N_307,In_175,In_165);
or U308 (N_308,In_528,In_161);
or U309 (N_309,In_19,In_124);
xnor U310 (N_310,In_723,In_639);
and U311 (N_311,In_233,In_727);
and U312 (N_312,In_133,In_1);
xnor U313 (N_313,In_493,In_96);
nand U314 (N_314,In_72,In_624);
nor U315 (N_315,In_379,In_62);
xor U316 (N_316,In_669,In_410);
nor U317 (N_317,In_510,In_2);
nand U318 (N_318,In_247,In_481);
and U319 (N_319,In_657,In_200);
xor U320 (N_320,In_566,In_229);
and U321 (N_321,In_719,In_304);
nor U322 (N_322,In_440,In_33);
xor U323 (N_323,In_652,In_642);
and U324 (N_324,In_544,In_500);
xor U325 (N_325,In_407,In_371);
xnor U326 (N_326,In_704,In_275);
or U327 (N_327,In_170,In_605);
xor U328 (N_328,In_747,In_227);
and U329 (N_329,In_464,In_129);
nand U330 (N_330,In_366,In_738);
nor U331 (N_331,In_611,In_580);
or U332 (N_332,In_116,In_506);
or U333 (N_333,In_320,In_722);
xnor U334 (N_334,In_321,In_186);
nor U335 (N_335,In_666,In_534);
xnor U336 (N_336,In_84,In_651);
and U337 (N_337,In_51,In_122);
nand U338 (N_338,In_570,In_465);
xnor U339 (N_339,In_424,In_655);
and U340 (N_340,In_178,In_99);
or U341 (N_341,In_707,In_442);
or U342 (N_342,In_39,In_511);
and U343 (N_343,In_34,In_110);
xor U344 (N_344,In_625,In_252);
or U345 (N_345,In_201,In_153);
nor U346 (N_346,In_713,In_205);
or U347 (N_347,In_443,In_212);
or U348 (N_348,In_381,In_701);
nor U349 (N_349,In_206,In_564);
nor U350 (N_350,In_93,In_610);
or U351 (N_351,In_203,In_52);
and U352 (N_352,In_476,In_601);
and U353 (N_353,In_517,In_732);
or U354 (N_354,In_163,In_145);
xnor U355 (N_355,In_220,In_520);
nand U356 (N_356,In_312,In_422);
and U357 (N_357,In_154,In_709);
nand U358 (N_358,In_285,In_193);
nand U359 (N_359,In_523,In_389);
and U360 (N_360,In_508,In_541);
xor U361 (N_361,In_49,In_38);
xnor U362 (N_362,In_254,In_48);
and U363 (N_363,In_656,In_24);
or U364 (N_364,In_315,In_81);
nand U365 (N_365,In_184,In_653);
xor U366 (N_366,In_21,In_257);
or U367 (N_367,In_60,In_104);
nor U368 (N_368,In_310,In_743);
nor U369 (N_369,In_208,In_28);
or U370 (N_370,In_317,In_54);
xnor U371 (N_371,In_308,In_6);
nor U372 (N_372,In_538,In_188);
and U373 (N_373,In_134,In_195);
or U374 (N_374,In_473,In_109);
or U375 (N_375,In_496,In_748);
or U376 (N_376,In_166,In_73);
and U377 (N_377,In_213,In_452);
nand U378 (N_378,In_129,In_670);
xnor U379 (N_379,In_690,In_147);
or U380 (N_380,In_516,In_283);
nor U381 (N_381,In_56,In_422);
and U382 (N_382,In_194,In_604);
nand U383 (N_383,In_502,In_279);
xnor U384 (N_384,In_407,In_723);
and U385 (N_385,In_502,In_188);
nand U386 (N_386,In_14,In_82);
nor U387 (N_387,In_534,In_745);
and U388 (N_388,In_45,In_372);
nor U389 (N_389,In_687,In_628);
nand U390 (N_390,In_575,In_325);
nand U391 (N_391,In_666,In_24);
xnor U392 (N_392,In_282,In_468);
nand U393 (N_393,In_354,In_480);
xor U394 (N_394,In_464,In_49);
nand U395 (N_395,In_298,In_201);
or U396 (N_396,In_263,In_357);
xor U397 (N_397,In_438,In_605);
xnor U398 (N_398,In_721,In_70);
nor U399 (N_399,In_343,In_66);
nor U400 (N_400,In_386,In_473);
nor U401 (N_401,In_615,In_446);
xnor U402 (N_402,In_569,In_101);
or U403 (N_403,In_439,In_120);
or U404 (N_404,In_517,In_677);
xor U405 (N_405,In_616,In_356);
and U406 (N_406,In_173,In_729);
or U407 (N_407,In_373,In_208);
xnor U408 (N_408,In_595,In_267);
and U409 (N_409,In_560,In_518);
or U410 (N_410,In_724,In_687);
or U411 (N_411,In_380,In_313);
or U412 (N_412,In_599,In_567);
or U413 (N_413,In_450,In_101);
nor U414 (N_414,In_13,In_402);
or U415 (N_415,In_271,In_403);
nand U416 (N_416,In_330,In_432);
nor U417 (N_417,In_619,In_466);
or U418 (N_418,In_572,In_684);
nand U419 (N_419,In_685,In_220);
nand U420 (N_420,In_248,In_519);
nand U421 (N_421,In_484,In_234);
nor U422 (N_422,In_486,In_635);
nor U423 (N_423,In_228,In_522);
and U424 (N_424,In_26,In_379);
xor U425 (N_425,In_455,In_136);
xor U426 (N_426,In_611,In_229);
nor U427 (N_427,In_211,In_213);
nor U428 (N_428,In_157,In_638);
nand U429 (N_429,In_133,In_35);
nor U430 (N_430,In_738,In_320);
and U431 (N_431,In_313,In_579);
xnor U432 (N_432,In_328,In_326);
xor U433 (N_433,In_117,In_23);
nor U434 (N_434,In_123,In_336);
nor U435 (N_435,In_293,In_420);
nand U436 (N_436,In_585,In_263);
xor U437 (N_437,In_91,In_715);
or U438 (N_438,In_89,In_551);
xor U439 (N_439,In_720,In_286);
and U440 (N_440,In_703,In_584);
or U441 (N_441,In_700,In_145);
or U442 (N_442,In_524,In_292);
nand U443 (N_443,In_403,In_356);
xnor U444 (N_444,In_342,In_612);
or U445 (N_445,In_466,In_61);
xnor U446 (N_446,In_366,In_325);
or U447 (N_447,In_560,In_151);
nor U448 (N_448,In_197,In_123);
xnor U449 (N_449,In_479,In_186);
and U450 (N_450,In_289,In_273);
and U451 (N_451,In_534,In_324);
xnor U452 (N_452,In_182,In_196);
or U453 (N_453,In_296,In_31);
xnor U454 (N_454,In_53,In_588);
or U455 (N_455,In_489,In_642);
or U456 (N_456,In_3,In_493);
xnor U457 (N_457,In_164,In_241);
and U458 (N_458,In_619,In_553);
or U459 (N_459,In_490,In_27);
and U460 (N_460,In_40,In_489);
and U461 (N_461,In_280,In_424);
xnor U462 (N_462,In_285,In_632);
and U463 (N_463,In_474,In_617);
and U464 (N_464,In_472,In_62);
xor U465 (N_465,In_161,In_463);
or U466 (N_466,In_475,In_139);
or U467 (N_467,In_164,In_737);
nand U468 (N_468,In_551,In_30);
xor U469 (N_469,In_589,In_663);
nand U470 (N_470,In_38,In_262);
and U471 (N_471,In_733,In_563);
and U472 (N_472,In_58,In_13);
nand U473 (N_473,In_502,In_196);
or U474 (N_474,In_345,In_262);
nand U475 (N_475,In_236,In_35);
nor U476 (N_476,In_21,In_48);
xor U477 (N_477,In_134,In_596);
nand U478 (N_478,In_612,In_346);
and U479 (N_479,In_632,In_537);
and U480 (N_480,In_71,In_560);
or U481 (N_481,In_52,In_563);
or U482 (N_482,In_99,In_68);
nor U483 (N_483,In_681,In_500);
xor U484 (N_484,In_461,In_593);
nand U485 (N_485,In_33,In_81);
and U486 (N_486,In_485,In_358);
nand U487 (N_487,In_725,In_454);
xnor U488 (N_488,In_148,In_572);
nand U489 (N_489,In_536,In_451);
or U490 (N_490,In_459,In_212);
nor U491 (N_491,In_498,In_260);
xnor U492 (N_492,In_370,In_572);
or U493 (N_493,In_238,In_91);
nor U494 (N_494,In_612,In_178);
nor U495 (N_495,In_276,In_345);
and U496 (N_496,In_616,In_359);
or U497 (N_497,In_32,In_121);
or U498 (N_498,In_38,In_96);
nand U499 (N_499,In_214,In_743);
nor U500 (N_500,In_71,In_340);
or U501 (N_501,In_473,In_703);
and U502 (N_502,In_673,In_408);
xnor U503 (N_503,In_518,In_417);
nand U504 (N_504,In_415,In_225);
nor U505 (N_505,In_741,In_438);
xnor U506 (N_506,In_514,In_253);
or U507 (N_507,In_178,In_455);
nand U508 (N_508,In_319,In_437);
nor U509 (N_509,In_240,In_80);
and U510 (N_510,In_149,In_706);
xnor U511 (N_511,In_129,In_700);
xor U512 (N_512,In_708,In_173);
nand U513 (N_513,In_742,In_42);
nor U514 (N_514,In_494,In_534);
and U515 (N_515,In_350,In_29);
nor U516 (N_516,In_121,In_223);
and U517 (N_517,In_177,In_596);
xor U518 (N_518,In_204,In_747);
or U519 (N_519,In_588,In_529);
or U520 (N_520,In_208,In_56);
or U521 (N_521,In_497,In_73);
and U522 (N_522,In_612,In_547);
xnor U523 (N_523,In_320,In_41);
and U524 (N_524,In_157,In_422);
nor U525 (N_525,In_201,In_71);
nor U526 (N_526,In_371,In_80);
xnor U527 (N_527,In_662,In_417);
or U528 (N_528,In_445,In_332);
nand U529 (N_529,In_83,In_602);
nor U530 (N_530,In_182,In_705);
nand U531 (N_531,In_488,In_570);
nor U532 (N_532,In_139,In_144);
or U533 (N_533,In_225,In_409);
nor U534 (N_534,In_25,In_522);
or U535 (N_535,In_620,In_253);
or U536 (N_536,In_40,In_171);
xnor U537 (N_537,In_574,In_534);
nor U538 (N_538,In_461,In_170);
nor U539 (N_539,In_356,In_270);
nor U540 (N_540,In_2,In_155);
and U541 (N_541,In_320,In_282);
and U542 (N_542,In_497,In_166);
and U543 (N_543,In_655,In_403);
nor U544 (N_544,In_150,In_517);
and U545 (N_545,In_425,In_716);
or U546 (N_546,In_494,In_337);
nand U547 (N_547,In_390,In_392);
nand U548 (N_548,In_22,In_501);
xnor U549 (N_549,In_363,In_58);
nor U550 (N_550,In_643,In_30);
or U551 (N_551,In_745,In_376);
or U552 (N_552,In_326,In_178);
and U553 (N_553,In_617,In_365);
and U554 (N_554,In_154,In_49);
and U555 (N_555,In_672,In_550);
or U556 (N_556,In_270,In_390);
nor U557 (N_557,In_495,In_68);
nor U558 (N_558,In_714,In_261);
or U559 (N_559,In_71,In_255);
nor U560 (N_560,In_345,In_613);
or U561 (N_561,In_223,In_105);
and U562 (N_562,In_585,In_635);
xor U563 (N_563,In_446,In_493);
or U564 (N_564,In_10,In_656);
nand U565 (N_565,In_661,In_43);
and U566 (N_566,In_421,In_502);
or U567 (N_567,In_512,In_423);
nor U568 (N_568,In_22,In_35);
and U569 (N_569,In_703,In_26);
or U570 (N_570,In_95,In_428);
nand U571 (N_571,In_417,In_561);
xnor U572 (N_572,In_21,In_252);
nor U573 (N_573,In_727,In_564);
nor U574 (N_574,In_439,In_549);
nand U575 (N_575,In_628,In_49);
or U576 (N_576,In_165,In_652);
and U577 (N_577,In_305,In_669);
or U578 (N_578,In_350,In_168);
or U579 (N_579,In_730,In_175);
or U580 (N_580,In_268,In_370);
xnor U581 (N_581,In_676,In_421);
and U582 (N_582,In_406,In_301);
nand U583 (N_583,In_414,In_512);
or U584 (N_584,In_425,In_235);
nor U585 (N_585,In_274,In_382);
nand U586 (N_586,In_483,In_221);
nand U587 (N_587,In_146,In_531);
nor U588 (N_588,In_375,In_361);
nor U589 (N_589,In_384,In_150);
and U590 (N_590,In_685,In_262);
or U591 (N_591,In_676,In_81);
and U592 (N_592,In_353,In_115);
nor U593 (N_593,In_277,In_592);
or U594 (N_594,In_44,In_59);
and U595 (N_595,In_138,In_691);
xnor U596 (N_596,In_647,In_198);
nor U597 (N_597,In_405,In_721);
nand U598 (N_598,In_243,In_540);
nand U599 (N_599,In_565,In_65);
nor U600 (N_600,In_15,In_152);
nor U601 (N_601,In_298,In_515);
and U602 (N_602,In_417,In_313);
and U603 (N_603,In_144,In_584);
and U604 (N_604,In_556,In_482);
or U605 (N_605,In_72,In_555);
xnor U606 (N_606,In_466,In_648);
or U607 (N_607,In_257,In_266);
nand U608 (N_608,In_302,In_276);
nor U609 (N_609,In_466,In_364);
and U610 (N_610,In_322,In_309);
or U611 (N_611,In_480,In_640);
or U612 (N_612,In_75,In_715);
nor U613 (N_613,In_739,In_144);
and U614 (N_614,In_467,In_698);
xnor U615 (N_615,In_34,In_194);
or U616 (N_616,In_85,In_319);
nor U617 (N_617,In_193,In_478);
and U618 (N_618,In_0,In_380);
or U619 (N_619,In_481,In_724);
or U620 (N_620,In_2,In_468);
xnor U621 (N_621,In_210,In_161);
nor U622 (N_622,In_138,In_719);
xor U623 (N_623,In_446,In_575);
xnor U624 (N_624,In_401,In_692);
nor U625 (N_625,In_167,In_453);
xor U626 (N_626,In_351,In_512);
xnor U627 (N_627,In_120,In_351);
nor U628 (N_628,In_307,In_676);
nor U629 (N_629,In_701,In_333);
nand U630 (N_630,In_215,In_131);
xor U631 (N_631,In_375,In_100);
nand U632 (N_632,In_438,In_581);
and U633 (N_633,In_67,In_694);
nand U634 (N_634,In_624,In_594);
nand U635 (N_635,In_87,In_221);
nor U636 (N_636,In_342,In_80);
nand U637 (N_637,In_583,In_475);
nand U638 (N_638,In_220,In_584);
and U639 (N_639,In_514,In_208);
or U640 (N_640,In_746,In_728);
nor U641 (N_641,In_710,In_127);
and U642 (N_642,In_604,In_142);
xor U643 (N_643,In_23,In_483);
or U644 (N_644,In_109,In_704);
xnor U645 (N_645,In_619,In_570);
nand U646 (N_646,In_700,In_368);
or U647 (N_647,In_408,In_565);
and U648 (N_648,In_120,In_496);
nor U649 (N_649,In_435,In_632);
or U650 (N_650,In_253,In_599);
and U651 (N_651,In_739,In_145);
nand U652 (N_652,In_223,In_554);
or U653 (N_653,In_121,In_677);
nor U654 (N_654,In_199,In_75);
or U655 (N_655,In_18,In_714);
nor U656 (N_656,In_102,In_524);
or U657 (N_657,In_694,In_616);
and U658 (N_658,In_324,In_350);
and U659 (N_659,In_299,In_428);
and U660 (N_660,In_743,In_530);
or U661 (N_661,In_469,In_62);
nand U662 (N_662,In_437,In_614);
and U663 (N_663,In_393,In_169);
and U664 (N_664,In_53,In_332);
xor U665 (N_665,In_478,In_241);
nand U666 (N_666,In_142,In_666);
nor U667 (N_667,In_322,In_487);
nor U668 (N_668,In_722,In_685);
or U669 (N_669,In_88,In_93);
xnor U670 (N_670,In_547,In_366);
or U671 (N_671,In_385,In_553);
and U672 (N_672,In_162,In_407);
nand U673 (N_673,In_119,In_145);
or U674 (N_674,In_366,In_657);
nor U675 (N_675,In_340,In_493);
or U676 (N_676,In_646,In_512);
and U677 (N_677,In_591,In_162);
and U678 (N_678,In_591,In_365);
or U679 (N_679,In_235,In_47);
nor U680 (N_680,In_96,In_13);
xor U681 (N_681,In_99,In_193);
xor U682 (N_682,In_388,In_443);
and U683 (N_683,In_746,In_710);
xnor U684 (N_684,In_438,In_43);
and U685 (N_685,In_409,In_68);
xnor U686 (N_686,In_675,In_692);
xor U687 (N_687,In_372,In_695);
nor U688 (N_688,In_230,In_406);
or U689 (N_689,In_333,In_698);
nand U690 (N_690,In_166,In_703);
nor U691 (N_691,In_615,In_206);
or U692 (N_692,In_411,In_314);
nor U693 (N_693,In_327,In_214);
nand U694 (N_694,In_437,In_538);
nand U695 (N_695,In_626,In_525);
nor U696 (N_696,In_260,In_400);
nand U697 (N_697,In_393,In_182);
nor U698 (N_698,In_116,In_709);
nor U699 (N_699,In_174,In_410);
and U700 (N_700,In_600,In_199);
nand U701 (N_701,In_394,In_307);
or U702 (N_702,In_205,In_623);
xor U703 (N_703,In_364,In_275);
nand U704 (N_704,In_723,In_257);
xor U705 (N_705,In_38,In_92);
and U706 (N_706,In_96,In_733);
nand U707 (N_707,In_169,In_625);
or U708 (N_708,In_59,In_480);
nor U709 (N_709,In_318,In_334);
nor U710 (N_710,In_421,In_383);
xor U711 (N_711,In_540,In_494);
or U712 (N_712,In_74,In_3);
xnor U713 (N_713,In_658,In_3);
or U714 (N_714,In_435,In_101);
or U715 (N_715,In_296,In_702);
and U716 (N_716,In_143,In_409);
or U717 (N_717,In_193,In_415);
xor U718 (N_718,In_141,In_338);
nand U719 (N_719,In_236,In_712);
and U720 (N_720,In_628,In_239);
nand U721 (N_721,In_375,In_435);
xor U722 (N_722,In_706,In_135);
xor U723 (N_723,In_61,In_731);
nor U724 (N_724,In_297,In_638);
nand U725 (N_725,In_233,In_105);
or U726 (N_726,In_675,In_656);
nor U727 (N_727,In_252,In_639);
and U728 (N_728,In_677,In_237);
nor U729 (N_729,In_533,In_146);
or U730 (N_730,In_169,In_44);
or U731 (N_731,In_601,In_51);
or U732 (N_732,In_543,In_647);
and U733 (N_733,In_445,In_412);
and U734 (N_734,In_671,In_575);
nor U735 (N_735,In_673,In_624);
and U736 (N_736,In_385,In_159);
nor U737 (N_737,In_545,In_245);
nor U738 (N_738,In_616,In_182);
or U739 (N_739,In_459,In_730);
nand U740 (N_740,In_572,In_614);
nor U741 (N_741,In_111,In_411);
nor U742 (N_742,In_561,In_559);
xor U743 (N_743,In_711,In_119);
xnor U744 (N_744,In_15,In_437);
nand U745 (N_745,In_140,In_615);
nor U746 (N_746,In_243,In_487);
nor U747 (N_747,In_535,In_679);
xor U748 (N_748,In_201,In_707);
nand U749 (N_749,In_392,In_408);
and U750 (N_750,In_568,In_284);
xnor U751 (N_751,In_135,In_328);
nand U752 (N_752,In_368,In_109);
xor U753 (N_753,In_71,In_159);
and U754 (N_754,In_636,In_228);
xor U755 (N_755,In_341,In_710);
nand U756 (N_756,In_673,In_170);
nor U757 (N_757,In_234,In_254);
and U758 (N_758,In_161,In_642);
or U759 (N_759,In_318,In_257);
nor U760 (N_760,In_522,In_394);
nor U761 (N_761,In_247,In_49);
or U762 (N_762,In_302,In_66);
or U763 (N_763,In_333,In_291);
nand U764 (N_764,In_394,In_326);
nor U765 (N_765,In_304,In_337);
nand U766 (N_766,In_372,In_43);
xnor U767 (N_767,In_683,In_551);
nor U768 (N_768,In_610,In_71);
or U769 (N_769,In_115,In_123);
xnor U770 (N_770,In_491,In_355);
xnor U771 (N_771,In_50,In_692);
or U772 (N_772,In_407,In_79);
nand U773 (N_773,In_292,In_137);
nand U774 (N_774,In_94,In_9);
and U775 (N_775,In_525,In_44);
and U776 (N_776,In_715,In_533);
or U777 (N_777,In_334,In_170);
or U778 (N_778,In_558,In_685);
nand U779 (N_779,In_668,In_363);
or U780 (N_780,In_461,In_101);
or U781 (N_781,In_426,In_185);
nand U782 (N_782,In_296,In_180);
nand U783 (N_783,In_385,In_638);
or U784 (N_784,In_215,In_180);
nor U785 (N_785,In_736,In_245);
xnor U786 (N_786,In_689,In_666);
and U787 (N_787,In_661,In_679);
nand U788 (N_788,In_484,In_673);
nand U789 (N_789,In_271,In_496);
nand U790 (N_790,In_733,In_488);
or U791 (N_791,In_2,In_455);
nor U792 (N_792,In_134,In_440);
nand U793 (N_793,In_327,In_164);
nand U794 (N_794,In_8,In_567);
xnor U795 (N_795,In_580,In_167);
or U796 (N_796,In_376,In_585);
nor U797 (N_797,In_362,In_556);
or U798 (N_798,In_689,In_391);
or U799 (N_799,In_644,In_559);
and U800 (N_800,In_0,In_99);
nand U801 (N_801,In_686,In_205);
xor U802 (N_802,In_557,In_744);
xnor U803 (N_803,In_652,In_565);
and U804 (N_804,In_320,In_622);
nand U805 (N_805,In_536,In_708);
and U806 (N_806,In_473,In_596);
or U807 (N_807,In_169,In_541);
or U808 (N_808,In_245,In_173);
nor U809 (N_809,In_144,In_195);
nand U810 (N_810,In_395,In_384);
nor U811 (N_811,In_659,In_140);
nor U812 (N_812,In_305,In_75);
xnor U813 (N_813,In_54,In_541);
and U814 (N_814,In_148,In_541);
nand U815 (N_815,In_399,In_58);
or U816 (N_816,In_346,In_515);
nand U817 (N_817,In_181,In_508);
xnor U818 (N_818,In_451,In_204);
and U819 (N_819,In_377,In_380);
and U820 (N_820,In_148,In_573);
nand U821 (N_821,In_589,In_409);
or U822 (N_822,In_252,In_498);
xnor U823 (N_823,In_694,In_640);
and U824 (N_824,In_210,In_219);
nor U825 (N_825,In_641,In_414);
and U826 (N_826,In_365,In_603);
nand U827 (N_827,In_319,In_405);
nor U828 (N_828,In_229,In_509);
nor U829 (N_829,In_296,In_365);
xor U830 (N_830,In_235,In_21);
nor U831 (N_831,In_478,In_104);
and U832 (N_832,In_474,In_54);
xnor U833 (N_833,In_673,In_366);
xor U834 (N_834,In_487,In_3);
xnor U835 (N_835,In_422,In_720);
xnor U836 (N_836,In_591,In_53);
nand U837 (N_837,In_721,In_733);
xor U838 (N_838,In_227,In_701);
nand U839 (N_839,In_110,In_188);
nand U840 (N_840,In_445,In_13);
or U841 (N_841,In_153,In_610);
and U842 (N_842,In_195,In_428);
or U843 (N_843,In_50,In_558);
and U844 (N_844,In_736,In_613);
or U845 (N_845,In_199,In_655);
xnor U846 (N_846,In_226,In_343);
nand U847 (N_847,In_613,In_623);
and U848 (N_848,In_13,In_429);
xor U849 (N_849,In_383,In_279);
nand U850 (N_850,In_287,In_506);
xor U851 (N_851,In_153,In_381);
nand U852 (N_852,In_278,In_531);
nor U853 (N_853,In_170,In_313);
nand U854 (N_854,In_101,In_301);
nand U855 (N_855,In_313,In_460);
xor U856 (N_856,In_551,In_12);
and U857 (N_857,In_12,In_637);
nor U858 (N_858,In_526,In_244);
or U859 (N_859,In_613,In_121);
and U860 (N_860,In_485,In_210);
and U861 (N_861,In_93,In_691);
nand U862 (N_862,In_517,In_491);
and U863 (N_863,In_644,In_142);
and U864 (N_864,In_307,In_362);
xnor U865 (N_865,In_297,In_285);
nor U866 (N_866,In_180,In_92);
or U867 (N_867,In_717,In_400);
and U868 (N_868,In_239,In_450);
and U869 (N_869,In_528,In_239);
nand U870 (N_870,In_682,In_730);
or U871 (N_871,In_60,In_644);
xor U872 (N_872,In_561,In_54);
or U873 (N_873,In_349,In_541);
nand U874 (N_874,In_487,In_670);
or U875 (N_875,In_481,In_411);
and U876 (N_876,In_15,In_46);
and U877 (N_877,In_628,In_304);
nor U878 (N_878,In_681,In_310);
nand U879 (N_879,In_477,In_371);
xnor U880 (N_880,In_462,In_654);
nor U881 (N_881,In_127,In_496);
or U882 (N_882,In_567,In_506);
xnor U883 (N_883,In_17,In_93);
xnor U884 (N_884,In_124,In_554);
xor U885 (N_885,In_364,In_345);
nand U886 (N_886,In_504,In_23);
nor U887 (N_887,In_639,In_619);
and U888 (N_888,In_709,In_463);
nor U889 (N_889,In_338,In_732);
xor U890 (N_890,In_493,In_253);
xor U891 (N_891,In_607,In_698);
xor U892 (N_892,In_194,In_143);
or U893 (N_893,In_361,In_27);
nand U894 (N_894,In_158,In_25);
nor U895 (N_895,In_243,In_467);
xor U896 (N_896,In_223,In_334);
nand U897 (N_897,In_13,In_611);
nand U898 (N_898,In_535,In_224);
and U899 (N_899,In_261,In_622);
and U900 (N_900,In_315,In_661);
xnor U901 (N_901,In_312,In_279);
nand U902 (N_902,In_504,In_291);
and U903 (N_903,In_25,In_624);
nand U904 (N_904,In_450,In_169);
nand U905 (N_905,In_513,In_255);
and U906 (N_906,In_84,In_417);
and U907 (N_907,In_446,In_494);
or U908 (N_908,In_350,In_68);
xor U909 (N_909,In_66,In_472);
nand U910 (N_910,In_390,In_293);
nand U911 (N_911,In_130,In_259);
or U912 (N_912,In_301,In_100);
nor U913 (N_913,In_486,In_619);
or U914 (N_914,In_668,In_416);
or U915 (N_915,In_610,In_717);
nand U916 (N_916,In_633,In_9);
xnor U917 (N_917,In_144,In_241);
and U918 (N_918,In_385,In_656);
and U919 (N_919,In_667,In_201);
and U920 (N_920,In_109,In_536);
nor U921 (N_921,In_737,In_744);
nor U922 (N_922,In_328,In_79);
nand U923 (N_923,In_8,In_238);
or U924 (N_924,In_223,In_100);
xor U925 (N_925,In_48,In_235);
xor U926 (N_926,In_284,In_282);
xor U927 (N_927,In_588,In_27);
and U928 (N_928,In_400,In_627);
or U929 (N_929,In_174,In_461);
nor U930 (N_930,In_487,In_171);
or U931 (N_931,In_629,In_503);
nor U932 (N_932,In_302,In_207);
and U933 (N_933,In_397,In_387);
or U934 (N_934,In_578,In_144);
nand U935 (N_935,In_348,In_707);
and U936 (N_936,In_342,In_350);
and U937 (N_937,In_673,In_571);
nor U938 (N_938,In_339,In_200);
nor U939 (N_939,In_495,In_61);
and U940 (N_940,In_205,In_343);
or U941 (N_941,In_685,In_348);
xnor U942 (N_942,In_99,In_110);
nand U943 (N_943,In_474,In_33);
and U944 (N_944,In_381,In_59);
and U945 (N_945,In_247,In_91);
xnor U946 (N_946,In_85,In_686);
and U947 (N_947,In_152,In_663);
xnor U948 (N_948,In_606,In_162);
nand U949 (N_949,In_380,In_730);
xor U950 (N_950,In_481,In_93);
or U951 (N_951,In_417,In_0);
nor U952 (N_952,In_325,In_709);
or U953 (N_953,In_218,In_614);
nand U954 (N_954,In_591,In_10);
xnor U955 (N_955,In_474,In_212);
and U956 (N_956,In_73,In_416);
and U957 (N_957,In_129,In_588);
xnor U958 (N_958,In_362,In_598);
xnor U959 (N_959,In_216,In_412);
nor U960 (N_960,In_629,In_540);
xnor U961 (N_961,In_275,In_436);
nor U962 (N_962,In_361,In_491);
nand U963 (N_963,In_466,In_439);
and U964 (N_964,In_247,In_141);
nor U965 (N_965,In_165,In_29);
nor U966 (N_966,In_127,In_284);
nand U967 (N_967,In_240,In_399);
and U968 (N_968,In_281,In_321);
or U969 (N_969,In_538,In_260);
nor U970 (N_970,In_50,In_167);
nor U971 (N_971,In_92,In_476);
nand U972 (N_972,In_483,In_50);
nor U973 (N_973,In_420,In_556);
nand U974 (N_974,In_563,In_94);
or U975 (N_975,In_371,In_417);
nor U976 (N_976,In_247,In_686);
or U977 (N_977,In_329,In_686);
xor U978 (N_978,In_281,In_501);
xnor U979 (N_979,In_133,In_249);
nor U980 (N_980,In_317,In_70);
and U981 (N_981,In_730,In_191);
or U982 (N_982,In_299,In_580);
nor U983 (N_983,In_227,In_430);
or U984 (N_984,In_480,In_717);
and U985 (N_985,In_720,In_201);
and U986 (N_986,In_693,In_204);
xor U987 (N_987,In_395,In_482);
nand U988 (N_988,In_404,In_290);
nor U989 (N_989,In_270,In_242);
or U990 (N_990,In_372,In_11);
nor U991 (N_991,In_688,In_214);
nor U992 (N_992,In_623,In_147);
or U993 (N_993,In_97,In_74);
nor U994 (N_994,In_92,In_623);
nor U995 (N_995,In_322,In_445);
nand U996 (N_996,In_232,In_704);
xor U997 (N_997,In_141,In_383);
and U998 (N_998,In_76,In_428);
or U999 (N_999,In_125,In_294);
nor U1000 (N_1000,N_303,N_738);
and U1001 (N_1001,N_789,N_235);
nor U1002 (N_1002,N_253,N_262);
or U1003 (N_1003,N_974,N_514);
and U1004 (N_1004,N_9,N_424);
nand U1005 (N_1005,N_243,N_746);
nand U1006 (N_1006,N_241,N_747);
xor U1007 (N_1007,N_247,N_300);
and U1008 (N_1008,N_357,N_242);
xor U1009 (N_1009,N_511,N_146);
or U1010 (N_1010,N_491,N_804);
nand U1011 (N_1011,N_376,N_682);
nand U1012 (N_1012,N_256,N_35);
xnor U1013 (N_1013,N_634,N_895);
or U1014 (N_1014,N_506,N_745);
xor U1015 (N_1015,N_344,N_609);
and U1016 (N_1016,N_957,N_86);
nand U1017 (N_1017,N_662,N_369);
nand U1018 (N_1018,N_655,N_2);
and U1019 (N_1019,N_534,N_388);
nand U1020 (N_1020,N_59,N_148);
xor U1021 (N_1021,N_577,N_210);
nor U1022 (N_1022,N_890,N_525);
and U1023 (N_1023,N_352,N_96);
and U1024 (N_1024,N_781,N_374);
xor U1025 (N_1025,N_685,N_674);
and U1026 (N_1026,N_765,N_283);
and U1027 (N_1027,N_702,N_697);
and U1028 (N_1028,N_778,N_908);
xnor U1029 (N_1029,N_666,N_350);
and U1030 (N_1030,N_589,N_153);
nand U1031 (N_1031,N_271,N_735);
nor U1032 (N_1032,N_751,N_251);
and U1033 (N_1033,N_721,N_232);
nand U1034 (N_1034,N_569,N_434);
xnor U1035 (N_1035,N_901,N_415);
nor U1036 (N_1036,N_503,N_586);
nand U1037 (N_1037,N_293,N_310);
and U1038 (N_1038,N_630,N_842);
xnor U1039 (N_1039,N_969,N_370);
and U1040 (N_1040,N_522,N_888);
nand U1041 (N_1041,N_692,N_460);
xor U1042 (N_1042,N_759,N_383);
nand U1043 (N_1043,N_177,N_298);
xor U1044 (N_1044,N_85,N_476);
and U1045 (N_1045,N_474,N_638);
xnor U1046 (N_1046,N_632,N_339);
and U1047 (N_1047,N_275,N_433);
or U1048 (N_1048,N_504,N_902);
nand U1049 (N_1049,N_80,N_653);
or U1050 (N_1050,N_933,N_118);
nor U1051 (N_1051,N_62,N_590);
xnor U1052 (N_1052,N_190,N_757);
or U1053 (N_1053,N_158,N_714);
nand U1054 (N_1054,N_451,N_749);
nor U1055 (N_1055,N_207,N_616);
and U1056 (N_1056,N_122,N_169);
and U1057 (N_1057,N_612,N_165);
nand U1058 (N_1058,N_677,N_250);
or U1059 (N_1059,N_464,N_830);
and U1060 (N_1060,N_209,N_940);
nand U1061 (N_1061,N_964,N_400);
nor U1062 (N_1062,N_429,N_663);
xnor U1063 (N_1063,N_208,N_260);
xor U1064 (N_1064,N_281,N_454);
and U1065 (N_1065,N_582,N_566);
xor U1066 (N_1066,N_646,N_156);
nand U1067 (N_1067,N_681,N_455);
xor U1068 (N_1068,N_294,N_659);
nor U1069 (N_1069,N_224,N_588);
nand U1070 (N_1070,N_91,N_529);
or U1071 (N_1071,N_617,N_696);
nor U1072 (N_1072,N_758,N_54);
nand U1073 (N_1073,N_73,N_136);
xnor U1074 (N_1074,N_314,N_564);
and U1075 (N_1075,N_329,N_572);
xnor U1076 (N_1076,N_23,N_623);
nand U1077 (N_1077,N_510,N_457);
or U1078 (N_1078,N_594,N_140);
and U1079 (N_1079,N_528,N_484);
nand U1080 (N_1080,N_462,N_797);
and U1081 (N_1081,N_8,N_337);
or U1082 (N_1082,N_186,N_205);
xor U1083 (N_1083,N_25,N_280);
or U1084 (N_1084,N_611,N_905);
nor U1085 (N_1085,N_29,N_107);
xor U1086 (N_1086,N_924,N_315);
xor U1087 (N_1087,N_548,N_166);
and U1088 (N_1088,N_785,N_768);
and U1089 (N_1089,N_371,N_626);
nor U1090 (N_1090,N_105,N_356);
and U1091 (N_1091,N_248,N_953);
and U1092 (N_1092,N_816,N_296);
and U1093 (N_1093,N_954,N_642);
xnor U1094 (N_1094,N_869,N_812);
xnor U1095 (N_1095,N_173,N_951);
and U1096 (N_1096,N_864,N_563);
nand U1097 (N_1097,N_643,N_212);
and U1098 (N_1098,N_762,N_414);
nand U1099 (N_1099,N_716,N_944);
or U1100 (N_1100,N_903,N_375);
or U1101 (N_1101,N_921,N_641);
xor U1102 (N_1102,N_992,N_684);
or U1103 (N_1103,N_852,N_79);
or U1104 (N_1104,N_958,N_809);
and U1105 (N_1105,N_95,N_452);
nor U1106 (N_1106,N_541,N_149);
or U1107 (N_1107,N_573,N_89);
nor U1108 (N_1108,N_81,N_167);
nor U1109 (N_1109,N_48,N_245);
nor U1110 (N_1110,N_907,N_627);
and U1111 (N_1111,N_889,N_448);
nand U1112 (N_1112,N_43,N_976);
xnor U1113 (N_1113,N_559,N_172);
nor U1114 (N_1114,N_238,N_555);
nand U1115 (N_1115,N_575,N_814);
xnor U1116 (N_1116,N_854,N_318);
or U1117 (N_1117,N_776,N_366);
nor U1118 (N_1118,N_328,N_479);
nor U1119 (N_1119,N_618,N_526);
or U1120 (N_1120,N_741,N_143);
xor U1121 (N_1121,N_792,N_710);
xor U1122 (N_1122,N_391,N_187);
nand U1123 (N_1123,N_636,N_715);
nor U1124 (N_1124,N_628,N_218);
nand U1125 (N_1125,N_267,N_996);
nand U1126 (N_1126,N_282,N_904);
and U1127 (N_1127,N_425,N_891);
xor U1128 (N_1128,N_977,N_246);
and U1129 (N_1129,N_19,N_911);
or U1130 (N_1130,N_341,N_1);
nor U1131 (N_1131,N_828,N_919);
xor U1132 (N_1132,N_377,N_740);
or U1133 (N_1133,N_703,N_881);
and U1134 (N_1134,N_239,N_693);
and U1135 (N_1135,N_113,N_130);
and U1136 (N_1136,N_335,N_614);
nand U1137 (N_1137,N_288,N_756);
nand U1138 (N_1138,N_423,N_732);
and U1139 (N_1139,N_116,N_955);
xnor U1140 (N_1140,N_578,N_39);
nand U1141 (N_1141,N_915,N_297);
and U1142 (N_1142,N_553,N_547);
nor U1143 (N_1143,N_446,N_126);
nor U1144 (N_1144,N_860,N_412);
nand U1145 (N_1145,N_321,N_517);
nor U1146 (N_1146,N_821,N_712);
nand U1147 (N_1147,N_603,N_203);
xor U1148 (N_1148,N_426,N_538);
xnor U1149 (N_1149,N_468,N_707);
or U1150 (N_1150,N_98,N_348);
nand U1151 (N_1151,N_824,N_191);
xnor U1152 (N_1152,N_66,N_754);
nand U1153 (N_1153,N_863,N_583);
and U1154 (N_1154,N_316,N_742);
nor U1155 (N_1155,N_57,N_93);
or U1156 (N_1156,N_979,N_436);
nor U1157 (N_1157,N_445,N_355);
xnor U1158 (N_1158,N_305,N_875);
and U1159 (N_1159,N_439,N_989);
nor U1160 (N_1160,N_309,N_160);
nand U1161 (N_1161,N_111,N_103);
and U1162 (N_1162,N_420,N_900);
or U1163 (N_1163,N_161,N_438);
nand U1164 (N_1164,N_61,N_92);
nand U1165 (N_1165,N_482,N_437);
nor U1166 (N_1166,N_380,N_11);
nand U1167 (N_1167,N_913,N_967);
nand U1168 (N_1168,N_724,N_497);
and U1169 (N_1169,N_13,N_711);
nand U1170 (N_1170,N_151,N_988);
xnor U1171 (N_1171,N_385,N_810);
xnor U1172 (N_1172,N_660,N_163);
nor U1173 (N_1173,N_58,N_894);
nor U1174 (N_1174,N_308,N_928);
or U1175 (N_1175,N_960,N_233);
nor U1176 (N_1176,N_815,N_923);
or U1177 (N_1177,N_651,N_405);
nor U1178 (N_1178,N_699,N_593);
and U1179 (N_1179,N_195,N_77);
or U1180 (N_1180,N_453,N_121);
xnor U1181 (N_1181,N_325,N_878);
nand U1182 (N_1182,N_304,N_544);
xnor U1183 (N_1183,N_200,N_927);
xor U1184 (N_1184,N_868,N_115);
nand U1185 (N_1185,N_847,N_899);
and U1186 (N_1186,N_40,N_270);
xnor U1187 (N_1187,N_222,N_197);
nand U1188 (N_1188,N_700,N_607);
or U1189 (N_1189,N_667,N_470);
nand U1190 (N_1190,N_65,N_500);
or U1191 (N_1191,N_384,N_273);
or U1192 (N_1192,N_560,N_463);
nand U1193 (N_1193,N_717,N_192);
nand U1194 (N_1194,N_787,N_272);
or U1195 (N_1195,N_42,N_83);
and U1196 (N_1196,N_132,N_520);
or U1197 (N_1197,N_961,N_743);
nand U1198 (N_1198,N_22,N_221);
xor U1199 (N_1199,N_543,N_202);
or U1200 (N_1200,N_893,N_109);
and U1201 (N_1201,N_21,N_284);
nand U1202 (N_1202,N_990,N_264);
and U1203 (N_1203,N_521,N_379);
or U1204 (N_1204,N_128,N_803);
and U1205 (N_1205,N_605,N_896);
nor U1206 (N_1206,N_856,N_258);
xnor U1207 (N_1207,N_606,N_88);
nor U1208 (N_1208,N_502,N_70);
and U1209 (N_1209,N_129,N_608);
nor U1210 (N_1210,N_817,N_972);
or U1211 (N_1211,N_211,N_495);
or U1212 (N_1212,N_596,N_786);
xor U1213 (N_1213,N_635,N_485);
nand U1214 (N_1214,N_276,N_155);
xnor U1215 (N_1215,N_885,N_935);
nor U1216 (N_1216,N_162,N_585);
nor U1217 (N_1217,N_650,N_368);
nor U1218 (N_1218,N_469,N_669);
xor U1219 (N_1219,N_975,N_41);
and U1220 (N_1220,N_857,N_230);
or U1221 (N_1221,N_215,N_392);
nor U1222 (N_1222,N_932,N_886);
nor U1223 (N_1223,N_999,N_862);
nor U1224 (N_1224,N_505,N_565);
nand U1225 (N_1225,N_189,N_458);
xor U1226 (N_1226,N_610,N_326);
and U1227 (N_1227,N_139,N_141);
and U1228 (N_1228,N_849,N_995);
or U1229 (N_1229,N_311,N_289);
and U1230 (N_1230,N_595,N_84);
xnor U1231 (N_1231,N_219,N_686);
nand U1232 (N_1232,N_841,N_154);
nor U1233 (N_1233,N_982,N_673);
and U1234 (N_1234,N_515,N_934);
xor U1235 (N_1235,N_265,N_447);
nor U1236 (N_1236,N_561,N_164);
xnor U1237 (N_1237,N_866,N_259);
or U1238 (N_1238,N_867,N_394);
or U1239 (N_1239,N_533,N_798);
nand U1240 (N_1240,N_488,N_680);
or U1241 (N_1241,N_125,N_225);
or U1242 (N_1242,N_10,N_748);
or U1243 (N_1243,N_340,N_55);
or U1244 (N_1244,N_973,N_509);
or U1245 (N_1245,N_45,N_362);
nor U1246 (N_1246,N_3,N_654);
nor U1247 (N_1247,N_584,N_184);
or U1248 (N_1248,N_939,N_552);
nand U1249 (N_1249,N_472,N_37);
or U1250 (N_1250,N_372,N_364);
xor U1251 (N_1251,N_591,N_941);
or U1252 (N_1252,N_327,N_870);
nand U1253 (N_1253,N_227,N_946);
nand U1254 (N_1254,N_317,N_771);
xor U1255 (N_1255,N_175,N_734);
and U1256 (N_1256,N_286,N_620);
nand U1257 (N_1257,N_373,N_807);
and U1258 (N_1258,N_631,N_966);
or U1259 (N_1259,N_825,N_475);
and U1260 (N_1260,N_604,N_997);
and U1261 (N_1261,N_850,N_938);
and U1262 (N_1262,N_4,N_645);
nand U1263 (N_1263,N_619,N_652);
xnor U1264 (N_1264,N_929,N_664);
and U1265 (N_1265,N_312,N_467);
xor U1266 (N_1266,N_461,N_358);
xor U1267 (N_1267,N_333,N_621);
xor U1268 (N_1268,N_535,N_237);
nand U1269 (N_1269,N_772,N_656);
xor U1270 (N_1270,N_450,N_912);
and U1271 (N_1271,N_922,N_382);
nand U1272 (N_1272,N_695,N_794);
nand U1273 (N_1273,N_257,N_287);
or U1274 (N_1274,N_401,N_806);
and U1275 (N_1275,N_49,N_948);
nor U1276 (N_1276,N_725,N_20);
or U1277 (N_1277,N_629,N_775);
or U1278 (N_1278,N_110,N_492);
or U1279 (N_1279,N_719,N_127);
and U1280 (N_1280,N_861,N_501);
and U1281 (N_1281,N_567,N_827);
or U1282 (N_1282,N_539,N_570);
nor U1283 (N_1283,N_959,N_324);
xor U1284 (N_1284,N_278,N_483);
xnor U1285 (N_1285,N_926,N_694);
nor U1286 (N_1286,N_32,N_490);
or U1287 (N_1287,N_234,N_920);
nor U1288 (N_1288,N_430,N_120);
or U1289 (N_1289,N_114,N_625);
xnor U1290 (N_1290,N_551,N_853);
or U1291 (N_1291,N_100,N_240);
xnor U1292 (N_1292,N_788,N_834);
xnor U1293 (N_1293,N_102,N_837);
or U1294 (N_1294,N_602,N_507);
nand U1295 (N_1295,N_887,N_813);
nor U1296 (N_1296,N_183,N_170);
xor U1297 (N_1297,N_942,N_678);
nor U1298 (N_1298,N_945,N_763);
nor U1299 (N_1299,N_213,N_831);
nor U1300 (N_1300,N_811,N_936);
xor U1301 (N_1301,N_440,N_581);
or U1302 (N_1302,N_550,N_131);
or U1303 (N_1303,N_925,N_87);
nand U1304 (N_1304,N_343,N_832);
nand U1305 (N_1305,N_793,N_365);
and U1306 (N_1306,N_637,N_349);
xor U1307 (N_1307,N_307,N_418);
and U1308 (N_1308,N_730,N_194);
xor U1309 (N_1309,N_351,N_963);
xnor U1310 (N_1310,N_723,N_579);
xnor U1311 (N_1311,N_68,N_268);
nand U1312 (N_1312,N_780,N_930);
nand U1313 (N_1313,N_897,N_252);
xnor U1314 (N_1314,N_112,N_640);
nor U1315 (N_1315,N_872,N_159);
and U1316 (N_1316,N_493,N_918);
and U1317 (N_1317,N_513,N_443);
nor U1318 (N_1318,N_404,N_279);
xnor U1319 (N_1319,N_135,N_877);
nor U1320 (N_1320,N_106,N_835);
nor U1321 (N_1321,N_519,N_459);
nor U1322 (N_1322,N_882,N_687);
and U1323 (N_1323,N_0,N_104);
and U1324 (N_1324,N_180,N_668);
nor U1325 (N_1325,N_683,N_367);
nand U1326 (N_1326,N_33,N_7);
nor U1327 (N_1327,N_399,N_398);
xor U1328 (N_1328,N_15,N_152);
nor U1329 (N_1329,N_389,N_644);
nor U1330 (N_1330,N_845,N_728);
or U1331 (N_1331,N_331,N_422);
nand U1332 (N_1332,N_592,N_465);
and U1333 (N_1333,N_226,N_193);
nor U1334 (N_1334,N_524,N_980);
xnor U1335 (N_1335,N_108,N_196);
nand U1336 (N_1336,N_123,N_790);
and U1337 (N_1337,N_839,N_873);
nor U1338 (N_1338,N_580,N_14);
nor U1339 (N_1339,N_556,N_983);
nand U1340 (N_1340,N_843,N_292);
and U1341 (N_1341,N_767,N_421);
or U1342 (N_1342,N_613,N_799);
nor U1343 (N_1343,N_576,N_508);
xor U1344 (N_1344,N_498,N_290);
xnor U1345 (N_1345,N_26,N_117);
or U1346 (N_1346,N_378,N_481);
nand U1347 (N_1347,N_171,N_532);
xor U1348 (N_1348,N_657,N_540);
and U1349 (N_1349,N_858,N_987);
nor U1350 (N_1350,N_204,N_546);
nor U1351 (N_1351,N_622,N_220);
and U1352 (N_1352,N_542,N_848);
and U1353 (N_1353,N_181,N_701);
xnor U1354 (N_1354,N_56,N_417);
nand U1355 (N_1355,N_16,N_427);
and U1356 (N_1356,N_338,N_442);
and U1357 (N_1357,N_261,N_456);
or U1358 (N_1358,N_536,N_319);
nor U1359 (N_1359,N_214,N_615);
and U1360 (N_1360,N_52,N_336);
xnor U1361 (N_1361,N_706,N_487);
nor U1362 (N_1362,N_855,N_523);
nand U1363 (N_1363,N_345,N_665);
or U1364 (N_1364,N_216,N_884);
or U1365 (N_1365,N_836,N_50);
nor U1366 (N_1366,N_883,N_347);
xor U1367 (N_1367,N_968,N_597);
nor U1368 (N_1368,N_598,N_601);
or U1369 (N_1369,N_914,N_994);
xor U1370 (N_1370,N_64,N_779);
or U1371 (N_1371,N_477,N_133);
nand U1372 (N_1372,N_931,N_28);
nor U1373 (N_1373,N_819,N_851);
xor U1374 (N_1374,N_299,N_393);
xor U1375 (N_1375,N_688,N_733);
xor U1376 (N_1376,N_431,N_244);
xor U1377 (N_1377,N_332,N_409);
nand U1378 (N_1378,N_182,N_138);
nor U1379 (N_1379,N_496,N_829);
nand U1380 (N_1380,N_600,N_231);
nand U1381 (N_1381,N_846,N_71);
nor U1382 (N_1382,N_60,N_78);
or U1383 (N_1383,N_722,N_647);
nand U1384 (N_1384,N_361,N_97);
xor U1385 (N_1385,N_142,N_6);
or U1386 (N_1386,N_24,N_63);
xnor U1387 (N_1387,N_998,N_47);
nor U1388 (N_1388,N_38,N_263);
nor U1389 (N_1389,N_744,N_174);
or U1390 (N_1390,N_970,N_134);
and U1391 (N_1391,N_549,N_770);
nor U1392 (N_1392,N_783,N_879);
and U1393 (N_1393,N_844,N_545);
nand U1394 (N_1394,N_334,N_124);
nand U1395 (N_1395,N_90,N_396);
nor U1396 (N_1396,N_826,N_360);
and U1397 (N_1397,N_822,N_962);
and U1398 (N_1398,N_704,N_760);
xor U1399 (N_1399,N_512,N_587);
or U1400 (N_1400,N_859,N_249);
nor U1401 (N_1401,N_554,N_568);
nand U1402 (N_1402,N_906,N_471);
xnor U1403 (N_1403,N_18,N_150);
and U1404 (N_1404,N_624,N_909);
and U1405 (N_1405,N_777,N_408);
or U1406 (N_1406,N_823,N_255);
nor U1407 (N_1407,N_670,N_675);
nand U1408 (N_1408,N_943,N_274);
and U1409 (N_1409,N_708,N_51);
xor U1410 (N_1410,N_69,N_689);
nor U1411 (N_1411,N_949,N_838);
or U1412 (N_1412,N_381,N_473);
nand U1413 (N_1413,N_435,N_737);
xnor U1414 (N_1414,N_397,N_705);
and U1415 (N_1415,N_910,N_984);
and U1416 (N_1416,N_478,N_416);
nor U1417 (N_1417,N_833,N_36);
or U1418 (N_1418,N_527,N_801);
xor U1419 (N_1419,N_185,N_75);
xnor U1420 (N_1420,N_137,N_764);
nand U1421 (N_1421,N_698,N_229);
nand U1422 (N_1422,N_769,N_99);
xnor U1423 (N_1423,N_727,N_277);
or U1424 (N_1424,N_486,N_363);
xnor U1425 (N_1425,N_649,N_880);
xor U1426 (N_1426,N_752,N_947);
or U1427 (N_1427,N_46,N_731);
nand U1428 (N_1428,N_346,N_386);
and U1429 (N_1429,N_661,N_753);
xnor U1430 (N_1430,N_516,N_217);
xnor U1431 (N_1431,N_729,N_648);
xor U1432 (N_1432,N_406,N_27);
nand U1433 (N_1433,N_726,N_444);
nor U1434 (N_1434,N_796,N_411);
nor U1435 (N_1435,N_199,N_269);
nor U1436 (N_1436,N_993,N_74);
nor U1437 (N_1437,N_53,N_201);
or U1438 (N_1438,N_971,N_639);
or U1439 (N_1439,N_94,N_320);
xor U1440 (N_1440,N_494,N_782);
or U1441 (N_1441,N_188,N_395);
or U1442 (N_1442,N_840,N_17);
and U1443 (N_1443,N_802,N_390);
and U1444 (N_1444,N_176,N_254);
and U1445 (N_1445,N_387,N_419);
nor U1446 (N_1446,N_354,N_795);
nand U1447 (N_1447,N_978,N_557);
and U1448 (N_1448,N_876,N_72);
nand U1449 (N_1449,N_295,N_691);
and U1450 (N_1450,N_428,N_671);
nor U1451 (N_1451,N_808,N_537);
nand U1452 (N_1452,N_518,N_755);
and U1453 (N_1453,N_410,N_917);
and U1454 (N_1454,N_736,N_266);
nor U1455 (N_1455,N_76,N_353);
or U1456 (N_1456,N_898,N_157);
nor U1457 (N_1457,N_530,N_403);
xor U1458 (N_1458,N_739,N_818);
and U1459 (N_1459,N_820,N_291);
nand U1460 (N_1460,N_5,N_489);
xnor U1461 (N_1461,N_871,N_228);
nand U1462 (N_1462,N_67,N_101);
or U1463 (N_1463,N_223,N_986);
or U1464 (N_1464,N_449,N_402);
nand U1465 (N_1465,N_147,N_679);
nand U1466 (N_1466,N_690,N_413);
nand U1467 (N_1467,N_892,N_773);
nand U1468 (N_1468,N_44,N_991);
or U1469 (N_1469,N_31,N_30);
nand U1470 (N_1470,N_168,N_145);
and U1471 (N_1471,N_432,N_672);
nor U1472 (N_1472,N_774,N_599);
or U1473 (N_1473,N_937,N_633);
nand U1474 (N_1474,N_407,N_709);
nor U1475 (N_1475,N_342,N_805);
nand U1476 (N_1476,N_558,N_12);
xnor U1477 (N_1477,N_562,N_178);
xnor U1478 (N_1478,N_800,N_499);
and U1479 (N_1479,N_206,N_119);
or U1480 (N_1480,N_236,N_965);
xnor U1481 (N_1481,N_323,N_865);
nor U1482 (N_1482,N_750,N_784);
xor U1483 (N_1483,N_302,N_301);
nand U1484 (N_1484,N_874,N_718);
and U1485 (N_1485,N_34,N_956);
nor U1486 (N_1486,N_916,N_179);
or U1487 (N_1487,N_574,N_359);
and U1488 (N_1488,N_480,N_441);
xnor U1489 (N_1489,N_198,N_791);
nand U1490 (N_1490,N_985,N_144);
and U1491 (N_1491,N_306,N_531);
or U1492 (N_1492,N_571,N_82);
nor U1493 (N_1493,N_761,N_466);
xnor U1494 (N_1494,N_285,N_981);
and U1495 (N_1495,N_950,N_676);
xnor U1496 (N_1496,N_658,N_330);
or U1497 (N_1497,N_322,N_313);
or U1498 (N_1498,N_952,N_713);
and U1499 (N_1499,N_766,N_720);
or U1500 (N_1500,N_613,N_158);
or U1501 (N_1501,N_503,N_674);
nor U1502 (N_1502,N_241,N_162);
or U1503 (N_1503,N_604,N_695);
and U1504 (N_1504,N_600,N_229);
and U1505 (N_1505,N_591,N_108);
nor U1506 (N_1506,N_419,N_311);
or U1507 (N_1507,N_430,N_948);
xnor U1508 (N_1508,N_321,N_849);
xnor U1509 (N_1509,N_167,N_773);
and U1510 (N_1510,N_835,N_362);
or U1511 (N_1511,N_504,N_845);
nand U1512 (N_1512,N_815,N_609);
or U1513 (N_1513,N_623,N_763);
nor U1514 (N_1514,N_172,N_75);
or U1515 (N_1515,N_249,N_585);
xnor U1516 (N_1516,N_301,N_258);
or U1517 (N_1517,N_558,N_234);
xor U1518 (N_1518,N_777,N_699);
nor U1519 (N_1519,N_656,N_207);
nand U1520 (N_1520,N_11,N_511);
xor U1521 (N_1521,N_465,N_754);
or U1522 (N_1522,N_611,N_560);
or U1523 (N_1523,N_633,N_314);
and U1524 (N_1524,N_469,N_921);
nor U1525 (N_1525,N_328,N_81);
nand U1526 (N_1526,N_818,N_812);
xnor U1527 (N_1527,N_602,N_448);
xor U1528 (N_1528,N_918,N_799);
or U1529 (N_1529,N_45,N_570);
and U1530 (N_1530,N_902,N_20);
and U1531 (N_1531,N_979,N_693);
or U1532 (N_1532,N_549,N_8);
or U1533 (N_1533,N_353,N_395);
and U1534 (N_1534,N_152,N_494);
xnor U1535 (N_1535,N_998,N_748);
nand U1536 (N_1536,N_561,N_871);
and U1537 (N_1537,N_948,N_311);
and U1538 (N_1538,N_560,N_962);
xor U1539 (N_1539,N_330,N_689);
nor U1540 (N_1540,N_558,N_899);
and U1541 (N_1541,N_949,N_674);
nor U1542 (N_1542,N_516,N_446);
and U1543 (N_1543,N_87,N_239);
nand U1544 (N_1544,N_919,N_440);
nor U1545 (N_1545,N_314,N_813);
nor U1546 (N_1546,N_786,N_316);
nand U1547 (N_1547,N_182,N_443);
and U1548 (N_1548,N_586,N_599);
xor U1549 (N_1549,N_721,N_94);
xnor U1550 (N_1550,N_31,N_334);
or U1551 (N_1551,N_493,N_8);
nor U1552 (N_1552,N_240,N_651);
nor U1553 (N_1553,N_4,N_660);
or U1554 (N_1554,N_704,N_712);
xor U1555 (N_1555,N_728,N_913);
xor U1556 (N_1556,N_32,N_208);
or U1557 (N_1557,N_843,N_245);
or U1558 (N_1558,N_197,N_238);
xnor U1559 (N_1559,N_193,N_211);
nor U1560 (N_1560,N_385,N_458);
or U1561 (N_1561,N_298,N_702);
xnor U1562 (N_1562,N_404,N_952);
and U1563 (N_1563,N_447,N_398);
and U1564 (N_1564,N_150,N_900);
nand U1565 (N_1565,N_674,N_683);
and U1566 (N_1566,N_979,N_351);
or U1567 (N_1567,N_213,N_707);
xnor U1568 (N_1568,N_122,N_90);
xor U1569 (N_1569,N_146,N_735);
and U1570 (N_1570,N_763,N_427);
nor U1571 (N_1571,N_400,N_99);
and U1572 (N_1572,N_258,N_814);
nand U1573 (N_1573,N_324,N_492);
nand U1574 (N_1574,N_59,N_567);
nand U1575 (N_1575,N_10,N_290);
nor U1576 (N_1576,N_486,N_385);
or U1577 (N_1577,N_886,N_138);
or U1578 (N_1578,N_672,N_359);
nand U1579 (N_1579,N_847,N_969);
or U1580 (N_1580,N_595,N_270);
and U1581 (N_1581,N_407,N_103);
nor U1582 (N_1582,N_77,N_377);
or U1583 (N_1583,N_386,N_20);
or U1584 (N_1584,N_196,N_749);
and U1585 (N_1585,N_437,N_54);
nand U1586 (N_1586,N_551,N_721);
nor U1587 (N_1587,N_240,N_266);
xor U1588 (N_1588,N_77,N_266);
or U1589 (N_1589,N_40,N_548);
and U1590 (N_1590,N_466,N_647);
or U1591 (N_1591,N_572,N_111);
xnor U1592 (N_1592,N_806,N_307);
nand U1593 (N_1593,N_951,N_8);
or U1594 (N_1594,N_194,N_478);
nand U1595 (N_1595,N_905,N_32);
xnor U1596 (N_1596,N_557,N_597);
xor U1597 (N_1597,N_357,N_195);
xor U1598 (N_1598,N_82,N_721);
nand U1599 (N_1599,N_502,N_879);
xor U1600 (N_1600,N_838,N_725);
xor U1601 (N_1601,N_797,N_866);
xor U1602 (N_1602,N_806,N_575);
nand U1603 (N_1603,N_946,N_12);
or U1604 (N_1604,N_951,N_997);
or U1605 (N_1605,N_915,N_637);
and U1606 (N_1606,N_362,N_817);
xor U1607 (N_1607,N_885,N_920);
xnor U1608 (N_1608,N_864,N_620);
or U1609 (N_1609,N_343,N_445);
nor U1610 (N_1610,N_354,N_412);
or U1611 (N_1611,N_898,N_944);
xor U1612 (N_1612,N_446,N_969);
or U1613 (N_1613,N_923,N_767);
xor U1614 (N_1614,N_173,N_847);
nor U1615 (N_1615,N_665,N_528);
or U1616 (N_1616,N_3,N_197);
and U1617 (N_1617,N_758,N_241);
nand U1618 (N_1618,N_591,N_59);
xnor U1619 (N_1619,N_106,N_613);
nand U1620 (N_1620,N_413,N_777);
and U1621 (N_1621,N_72,N_983);
and U1622 (N_1622,N_561,N_825);
and U1623 (N_1623,N_336,N_5);
or U1624 (N_1624,N_243,N_49);
xor U1625 (N_1625,N_764,N_578);
xor U1626 (N_1626,N_415,N_649);
nand U1627 (N_1627,N_446,N_46);
xor U1628 (N_1628,N_703,N_715);
or U1629 (N_1629,N_392,N_155);
nor U1630 (N_1630,N_536,N_743);
xor U1631 (N_1631,N_640,N_805);
or U1632 (N_1632,N_35,N_394);
nor U1633 (N_1633,N_499,N_3);
and U1634 (N_1634,N_832,N_631);
xnor U1635 (N_1635,N_447,N_590);
and U1636 (N_1636,N_65,N_542);
nor U1637 (N_1637,N_922,N_826);
xnor U1638 (N_1638,N_305,N_29);
and U1639 (N_1639,N_942,N_675);
nor U1640 (N_1640,N_299,N_948);
nor U1641 (N_1641,N_163,N_78);
or U1642 (N_1642,N_303,N_943);
xnor U1643 (N_1643,N_926,N_82);
nand U1644 (N_1644,N_267,N_976);
nand U1645 (N_1645,N_341,N_307);
xnor U1646 (N_1646,N_212,N_7);
nand U1647 (N_1647,N_832,N_608);
nand U1648 (N_1648,N_937,N_635);
nand U1649 (N_1649,N_183,N_914);
xnor U1650 (N_1650,N_72,N_858);
and U1651 (N_1651,N_454,N_143);
nor U1652 (N_1652,N_252,N_258);
xnor U1653 (N_1653,N_729,N_831);
xor U1654 (N_1654,N_632,N_114);
xor U1655 (N_1655,N_0,N_167);
nor U1656 (N_1656,N_802,N_164);
nor U1657 (N_1657,N_369,N_487);
or U1658 (N_1658,N_441,N_596);
and U1659 (N_1659,N_482,N_110);
nand U1660 (N_1660,N_507,N_389);
or U1661 (N_1661,N_76,N_20);
xor U1662 (N_1662,N_847,N_323);
nand U1663 (N_1663,N_991,N_878);
nand U1664 (N_1664,N_258,N_57);
nand U1665 (N_1665,N_211,N_110);
nand U1666 (N_1666,N_745,N_520);
nor U1667 (N_1667,N_271,N_869);
nand U1668 (N_1668,N_907,N_178);
xor U1669 (N_1669,N_324,N_305);
and U1670 (N_1670,N_905,N_83);
xnor U1671 (N_1671,N_126,N_26);
or U1672 (N_1672,N_138,N_153);
nor U1673 (N_1673,N_950,N_994);
and U1674 (N_1674,N_757,N_539);
and U1675 (N_1675,N_843,N_502);
xor U1676 (N_1676,N_843,N_875);
nor U1677 (N_1677,N_305,N_489);
nor U1678 (N_1678,N_926,N_560);
nor U1679 (N_1679,N_838,N_717);
nor U1680 (N_1680,N_236,N_814);
or U1681 (N_1681,N_979,N_339);
or U1682 (N_1682,N_231,N_815);
nor U1683 (N_1683,N_338,N_404);
nor U1684 (N_1684,N_637,N_362);
nor U1685 (N_1685,N_307,N_591);
nor U1686 (N_1686,N_771,N_849);
nand U1687 (N_1687,N_927,N_224);
and U1688 (N_1688,N_57,N_948);
or U1689 (N_1689,N_789,N_953);
nand U1690 (N_1690,N_631,N_206);
or U1691 (N_1691,N_296,N_539);
and U1692 (N_1692,N_949,N_870);
and U1693 (N_1693,N_105,N_89);
or U1694 (N_1694,N_22,N_820);
or U1695 (N_1695,N_616,N_398);
xor U1696 (N_1696,N_810,N_671);
and U1697 (N_1697,N_745,N_823);
nand U1698 (N_1698,N_709,N_430);
nor U1699 (N_1699,N_5,N_688);
and U1700 (N_1700,N_184,N_575);
nor U1701 (N_1701,N_640,N_8);
nor U1702 (N_1702,N_622,N_659);
nor U1703 (N_1703,N_221,N_906);
nor U1704 (N_1704,N_928,N_450);
or U1705 (N_1705,N_12,N_734);
or U1706 (N_1706,N_811,N_851);
or U1707 (N_1707,N_87,N_253);
nor U1708 (N_1708,N_254,N_612);
and U1709 (N_1709,N_410,N_670);
nor U1710 (N_1710,N_537,N_609);
xor U1711 (N_1711,N_301,N_943);
nor U1712 (N_1712,N_99,N_868);
or U1713 (N_1713,N_268,N_934);
xnor U1714 (N_1714,N_138,N_3);
or U1715 (N_1715,N_685,N_720);
or U1716 (N_1716,N_852,N_956);
and U1717 (N_1717,N_31,N_578);
nor U1718 (N_1718,N_842,N_406);
nand U1719 (N_1719,N_543,N_640);
xor U1720 (N_1720,N_816,N_347);
xor U1721 (N_1721,N_808,N_452);
and U1722 (N_1722,N_39,N_248);
or U1723 (N_1723,N_728,N_313);
or U1724 (N_1724,N_406,N_185);
nor U1725 (N_1725,N_150,N_351);
and U1726 (N_1726,N_67,N_292);
nand U1727 (N_1727,N_909,N_259);
xor U1728 (N_1728,N_572,N_381);
nor U1729 (N_1729,N_528,N_551);
nand U1730 (N_1730,N_645,N_58);
and U1731 (N_1731,N_867,N_890);
nor U1732 (N_1732,N_527,N_224);
and U1733 (N_1733,N_503,N_284);
xor U1734 (N_1734,N_249,N_573);
nor U1735 (N_1735,N_601,N_561);
nand U1736 (N_1736,N_62,N_562);
nor U1737 (N_1737,N_382,N_95);
nand U1738 (N_1738,N_619,N_705);
or U1739 (N_1739,N_828,N_504);
and U1740 (N_1740,N_268,N_970);
nand U1741 (N_1741,N_612,N_155);
nor U1742 (N_1742,N_498,N_653);
nand U1743 (N_1743,N_573,N_986);
xnor U1744 (N_1744,N_236,N_784);
nor U1745 (N_1745,N_135,N_26);
xnor U1746 (N_1746,N_363,N_196);
nand U1747 (N_1747,N_545,N_579);
and U1748 (N_1748,N_848,N_512);
or U1749 (N_1749,N_589,N_301);
and U1750 (N_1750,N_450,N_383);
nor U1751 (N_1751,N_948,N_136);
and U1752 (N_1752,N_267,N_16);
xnor U1753 (N_1753,N_711,N_566);
xor U1754 (N_1754,N_272,N_399);
nor U1755 (N_1755,N_249,N_840);
xnor U1756 (N_1756,N_278,N_986);
and U1757 (N_1757,N_283,N_684);
or U1758 (N_1758,N_495,N_872);
or U1759 (N_1759,N_343,N_545);
and U1760 (N_1760,N_642,N_785);
nand U1761 (N_1761,N_87,N_86);
or U1762 (N_1762,N_915,N_590);
xor U1763 (N_1763,N_463,N_339);
and U1764 (N_1764,N_32,N_631);
or U1765 (N_1765,N_430,N_781);
nor U1766 (N_1766,N_316,N_194);
xnor U1767 (N_1767,N_83,N_490);
xnor U1768 (N_1768,N_63,N_458);
or U1769 (N_1769,N_149,N_952);
and U1770 (N_1770,N_99,N_877);
and U1771 (N_1771,N_655,N_605);
and U1772 (N_1772,N_208,N_705);
nor U1773 (N_1773,N_394,N_211);
xnor U1774 (N_1774,N_302,N_663);
or U1775 (N_1775,N_190,N_794);
or U1776 (N_1776,N_947,N_618);
or U1777 (N_1777,N_155,N_551);
xnor U1778 (N_1778,N_468,N_1);
nor U1779 (N_1779,N_47,N_175);
xor U1780 (N_1780,N_224,N_566);
nor U1781 (N_1781,N_895,N_611);
xnor U1782 (N_1782,N_270,N_300);
nor U1783 (N_1783,N_858,N_964);
or U1784 (N_1784,N_594,N_925);
nor U1785 (N_1785,N_887,N_685);
or U1786 (N_1786,N_573,N_667);
xor U1787 (N_1787,N_294,N_700);
nand U1788 (N_1788,N_484,N_82);
or U1789 (N_1789,N_78,N_668);
or U1790 (N_1790,N_51,N_105);
xor U1791 (N_1791,N_562,N_565);
and U1792 (N_1792,N_408,N_920);
nor U1793 (N_1793,N_466,N_343);
and U1794 (N_1794,N_828,N_238);
nor U1795 (N_1795,N_775,N_616);
and U1796 (N_1796,N_190,N_750);
or U1797 (N_1797,N_281,N_812);
nand U1798 (N_1798,N_685,N_919);
or U1799 (N_1799,N_112,N_495);
and U1800 (N_1800,N_356,N_924);
nand U1801 (N_1801,N_371,N_424);
xor U1802 (N_1802,N_593,N_3);
and U1803 (N_1803,N_484,N_778);
nand U1804 (N_1804,N_177,N_741);
xnor U1805 (N_1805,N_89,N_557);
nor U1806 (N_1806,N_610,N_808);
nor U1807 (N_1807,N_493,N_836);
xnor U1808 (N_1808,N_473,N_890);
xnor U1809 (N_1809,N_561,N_793);
nor U1810 (N_1810,N_357,N_259);
and U1811 (N_1811,N_685,N_35);
nand U1812 (N_1812,N_676,N_607);
and U1813 (N_1813,N_760,N_505);
and U1814 (N_1814,N_485,N_136);
nor U1815 (N_1815,N_609,N_380);
xnor U1816 (N_1816,N_82,N_599);
and U1817 (N_1817,N_759,N_935);
and U1818 (N_1818,N_890,N_309);
or U1819 (N_1819,N_787,N_634);
and U1820 (N_1820,N_480,N_216);
nand U1821 (N_1821,N_723,N_305);
nand U1822 (N_1822,N_271,N_555);
nor U1823 (N_1823,N_915,N_887);
and U1824 (N_1824,N_790,N_602);
or U1825 (N_1825,N_248,N_93);
xnor U1826 (N_1826,N_463,N_616);
nor U1827 (N_1827,N_197,N_585);
xnor U1828 (N_1828,N_345,N_947);
or U1829 (N_1829,N_222,N_445);
xor U1830 (N_1830,N_416,N_846);
nor U1831 (N_1831,N_788,N_391);
or U1832 (N_1832,N_161,N_455);
nor U1833 (N_1833,N_48,N_151);
nand U1834 (N_1834,N_202,N_540);
and U1835 (N_1835,N_106,N_808);
nor U1836 (N_1836,N_703,N_594);
xor U1837 (N_1837,N_350,N_310);
xor U1838 (N_1838,N_52,N_395);
nand U1839 (N_1839,N_806,N_511);
xor U1840 (N_1840,N_325,N_131);
nand U1841 (N_1841,N_469,N_567);
and U1842 (N_1842,N_911,N_767);
nand U1843 (N_1843,N_333,N_820);
and U1844 (N_1844,N_860,N_732);
and U1845 (N_1845,N_91,N_601);
nand U1846 (N_1846,N_371,N_647);
nand U1847 (N_1847,N_319,N_232);
xor U1848 (N_1848,N_390,N_651);
or U1849 (N_1849,N_225,N_691);
nor U1850 (N_1850,N_535,N_965);
or U1851 (N_1851,N_174,N_473);
or U1852 (N_1852,N_477,N_422);
nor U1853 (N_1853,N_687,N_559);
xnor U1854 (N_1854,N_312,N_872);
nor U1855 (N_1855,N_711,N_422);
and U1856 (N_1856,N_828,N_195);
or U1857 (N_1857,N_753,N_866);
or U1858 (N_1858,N_331,N_754);
nand U1859 (N_1859,N_300,N_870);
or U1860 (N_1860,N_288,N_280);
and U1861 (N_1861,N_960,N_927);
nand U1862 (N_1862,N_780,N_628);
and U1863 (N_1863,N_451,N_676);
or U1864 (N_1864,N_273,N_595);
nand U1865 (N_1865,N_358,N_997);
or U1866 (N_1866,N_724,N_977);
or U1867 (N_1867,N_65,N_336);
and U1868 (N_1868,N_995,N_696);
or U1869 (N_1869,N_352,N_224);
xor U1870 (N_1870,N_225,N_72);
or U1871 (N_1871,N_954,N_577);
xor U1872 (N_1872,N_514,N_795);
or U1873 (N_1873,N_880,N_559);
xor U1874 (N_1874,N_82,N_300);
xor U1875 (N_1875,N_267,N_925);
nor U1876 (N_1876,N_626,N_344);
and U1877 (N_1877,N_518,N_995);
and U1878 (N_1878,N_839,N_369);
and U1879 (N_1879,N_141,N_987);
xor U1880 (N_1880,N_522,N_44);
xnor U1881 (N_1881,N_282,N_410);
nand U1882 (N_1882,N_840,N_627);
xnor U1883 (N_1883,N_807,N_281);
or U1884 (N_1884,N_238,N_254);
nor U1885 (N_1885,N_649,N_130);
and U1886 (N_1886,N_70,N_235);
or U1887 (N_1887,N_372,N_354);
nor U1888 (N_1888,N_935,N_891);
nand U1889 (N_1889,N_895,N_239);
or U1890 (N_1890,N_775,N_588);
xnor U1891 (N_1891,N_25,N_502);
nor U1892 (N_1892,N_620,N_970);
nor U1893 (N_1893,N_917,N_135);
nand U1894 (N_1894,N_105,N_500);
xor U1895 (N_1895,N_832,N_852);
nor U1896 (N_1896,N_787,N_196);
or U1897 (N_1897,N_671,N_175);
xnor U1898 (N_1898,N_274,N_937);
xnor U1899 (N_1899,N_536,N_15);
xor U1900 (N_1900,N_842,N_474);
nand U1901 (N_1901,N_70,N_926);
or U1902 (N_1902,N_667,N_78);
or U1903 (N_1903,N_757,N_100);
or U1904 (N_1904,N_506,N_5);
nand U1905 (N_1905,N_395,N_298);
nor U1906 (N_1906,N_287,N_193);
nor U1907 (N_1907,N_887,N_657);
and U1908 (N_1908,N_875,N_851);
and U1909 (N_1909,N_780,N_253);
and U1910 (N_1910,N_644,N_559);
nand U1911 (N_1911,N_528,N_967);
nor U1912 (N_1912,N_499,N_331);
nor U1913 (N_1913,N_275,N_371);
nand U1914 (N_1914,N_674,N_417);
nor U1915 (N_1915,N_518,N_289);
xor U1916 (N_1916,N_461,N_611);
nand U1917 (N_1917,N_968,N_351);
or U1918 (N_1918,N_486,N_362);
or U1919 (N_1919,N_818,N_724);
nor U1920 (N_1920,N_330,N_47);
and U1921 (N_1921,N_381,N_485);
and U1922 (N_1922,N_784,N_163);
and U1923 (N_1923,N_176,N_117);
and U1924 (N_1924,N_808,N_436);
nand U1925 (N_1925,N_71,N_799);
nor U1926 (N_1926,N_561,N_762);
or U1927 (N_1927,N_501,N_841);
nand U1928 (N_1928,N_266,N_714);
nor U1929 (N_1929,N_269,N_967);
nor U1930 (N_1930,N_845,N_443);
or U1931 (N_1931,N_385,N_464);
or U1932 (N_1932,N_51,N_974);
xnor U1933 (N_1933,N_886,N_28);
nand U1934 (N_1934,N_204,N_811);
nor U1935 (N_1935,N_457,N_256);
nand U1936 (N_1936,N_739,N_245);
and U1937 (N_1937,N_946,N_299);
and U1938 (N_1938,N_216,N_683);
and U1939 (N_1939,N_715,N_372);
nand U1940 (N_1940,N_462,N_335);
xor U1941 (N_1941,N_912,N_436);
and U1942 (N_1942,N_447,N_43);
xor U1943 (N_1943,N_625,N_865);
and U1944 (N_1944,N_110,N_264);
or U1945 (N_1945,N_825,N_685);
xnor U1946 (N_1946,N_442,N_113);
nand U1947 (N_1947,N_256,N_948);
nand U1948 (N_1948,N_913,N_684);
and U1949 (N_1949,N_502,N_362);
xnor U1950 (N_1950,N_661,N_160);
or U1951 (N_1951,N_851,N_768);
and U1952 (N_1952,N_536,N_520);
nor U1953 (N_1953,N_274,N_858);
or U1954 (N_1954,N_695,N_747);
and U1955 (N_1955,N_838,N_208);
nor U1956 (N_1956,N_779,N_30);
xnor U1957 (N_1957,N_936,N_509);
nor U1958 (N_1958,N_539,N_4);
or U1959 (N_1959,N_745,N_123);
or U1960 (N_1960,N_678,N_403);
and U1961 (N_1961,N_887,N_965);
or U1962 (N_1962,N_663,N_93);
nand U1963 (N_1963,N_867,N_955);
nor U1964 (N_1964,N_196,N_235);
nand U1965 (N_1965,N_556,N_741);
nand U1966 (N_1966,N_483,N_906);
and U1967 (N_1967,N_604,N_123);
or U1968 (N_1968,N_76,N_425);
nor U1969 (N_1969,N_827,N_991);
nor U1970 (N_1970,N_993,N_301);
or U1971 (N_1971,N_59,N_484);
nor U1972 (N_1972,N_629,N_574);
and U1973 (N_1973,N_851,N_434);
nor U1974 (N_1974,N_355,N_335);
nor U1975 (N_1975,N_881,N_555);
nand U1976 (N_1976,N_466,N_311);
and U1977 (N_1977,N_525,N_137);
nor U1978 (N_1978,N_874,N_521);
xor U1979 (N_1979,N_712,N_499);
nand U1980 (N_1980,N_335,N_406);
and U1981 (N_1981,N_938,N_410);
and U1982 (N_1982,N_968,N_53);
nand U1983 (N_1983,N_153,N_980);
xor U1984 (N_1984,N_895,N_131);
or U1985 (N_1985,N_861,N_759);
and U1986 (N_1986,N_520,N_0);
and U1987 (N_1987,N_437,N_881);
xnor U1988 (N_1988,N_926,N_752);
nor U1989 (N_1989,N_34,N_787);
or U1990 (N_1990,N_2,N_270);
and U1991 (N_1991,N_100,N_863);
or U1992 (N_1992,N_984,N_774);
nor U1993 (N_1993,N_376,N_5);
nand U1994 (N_1994,N_407,N_554);
nor U1995 (N_1995,N_175,N_321);
xnor U1996 (N_1996,N_709,N_644);
and U1997 (N_1997,N_585,N_44);
and U1998 (N_1998,N_972,N_204);
or U1999 (N_1999,N_262,N_987);
xor U2000 (N_2000,N_1393,N_1143);
nand U2001 (N_2001,N_1302,N_1010);
nand U2002 (N_2002,N_1792,N_1111);
xnor U2003 (N_2003,N_1548,N_1445);
and U2004 (N_2004,N_1529,N_1171);
and U2005 (N_2005,N_1704,N_1468);
nor U2006 (N_2006,N_1084,N_1401);
xnor U2007 (N_2007,N_1581,N_1169);
xor U2008 (N_2008,N_1956,N_1073);
xnor U2009 (N_2009,N_1103,N_1141);
nor U2010 (N_2010,N_1561,N_1244);
and U2011 (N_2011,N_1379,N_1504);
or U2012 (N_2012,N_1148,N_1885);
xnor U2013 (N_2013,N_1672,N_1368);
nor U2014 (N_2014,N_1353,N_1452);
or U2015 (N_2015,N_1791,N_1205);
nand U2016 (N_2016,N_1824,N_1714);
nor U2017 (N_2017,N_1499,N_1950);
xnor U2018 (N_2018,N_1895,N_1695);
xnor U2019 (N_2019,N_1182,N_1159);
nand U2020 (N_2020,N_1338,N_1803);
and U2021 (N_2021,N_1640,N_1936);
xor U2022 (N_2022,N_1115,N_1594);
or U2023 (N_2023,N_1264,N_1736);
xor U2024 (N_2024,N_1013,N_1218);
nand U2025 (N_2025,N_1390,N_1252);
nor U2026 (N_2026,N_1707,N_1836);
nor U2027 (N_2027,N_1643,N_1727);
nor U2028 (N_2028,N_1217,N_1523);
xnor U2029 (N_2029,N_1380,N_1577);
nand U2030 (N_2030,N_1710,N_1097);
nor U2031 (N_2031,N_1224,N_1023);
nor U2032 (N_2032,N_1914,N_1237);
nand U2033 (N_2033,N_1630,N_1460);
and U2034 (N_2034,N_1133,N_1656);
xnor U2035 (N_2035,N_1383,N_1279);
or U2036 (N_2036,N_1170,N_1689);
or U2037 (N_2037,N_1278,N_1729);
and U2038 (N_2038,N_1344,N_1832);
and U2039 (N_2039,N_1785,N_1453);
nand U2040 (N_2040,N_1846,N_1022);
nor U2041 (N_2041,N_1873,N_1860);
xor U2042 (N_2042,N_1810,N_1038);
nor U2043 (N_2043,N_1705,N_1905);
or U2044 (N_2044,N_1116,N_1228);
nand U2045 (N_2045,N_1417,N_1756);
or U2046 (N_2046,N_1029,N_1996);
nand U2047 (N_2047,N_1871,N_1197);
xor U2048 (N_2048,N_1564,N_1247);
nand U2049 (N_2049,N_1907,N_1476);
nand U2050 (N_2050,N_1855,N_1250);
xor U2051 (N_2051,N_1935,N_1575);
nand U2052 (N_2052,N_1555,N_1212);
nand U2053 (N_2053,N_1176,N_1489);
or U2054 (N_2054,N_1520,N_1089);
or U2055 (N_2055,N_1969,N_1915);
and U2056 (N_2056,N_1110,N_1214);
nor U2057 (N_2057,N_1139,N_1168);
and U2058 (N_2058,N_1323,N_1617);
or U2059 (N_2059,N_1986,N_1373);
and U2060 (N_2060,N_1844,N_1501);
xnor U2061 (N_2061,N_1590,N_1028);
and U2062 (N_2062,N_1075,N_1574);
nor U2063 (N_2063,N_1222,N_1475);
nor U2064 (N_2064,N_1778,N_1507);
or U2065 (N_2065,N_1641,N_1067);
or U2066 (N_2066,N_1734,N_1570);
nor U2067 (N_2067,N_1632,N_1653);
or U2068 (N_2068,N_1544,N_1709);
and U2069 (N_2069,N_1271,N_1203);
nor U2070 (N_2070,N_1195,N_1358);
and U2071 (N_2071,N_1891,N_1443);
and U2072 (N_2072,N_1510,N_1807);
or U2073 (N_2073,N_1400,N_1151);
and U2074 (N_2074,N_1137,N_1883);
nand U2075 (N_2075,N_1684,N_1955);
and U2076 (N_2076,N_1953,N_1193);
nor U2077 (N_2077,N_1863,N_1861);
nor U2078 (N_2078,N_1668,N_1306);
and U2079 (N_2079,N_1127,N_1649);
or U2080 (N_2080,N_1455,N_1093);
nor U2081 (N_2081,N_1335,N_1738);
or U2082 (N_2082,N_1864,N_1790);
nor U2083 (N_2083,N_1675,N_1341);
or U2084 (N_2084,N_1181,N_1773);
or U2085 (N_2085,N_1291,N_1673);
and U2086 (N_2086,N_1929,N_1776);
nand U2087 (N_2087,N_1389,N_1300);
and U2088 (N_2088,N_1613,N_1866);
nor U2089 (N_2089,N_1669,N_1635);
or U2090 (N_2090,N_1772,N_1098);
xor U2091 (N_2091,N_1842,N_1664);
and U2092 (N_2092,N_1311,N_1216);
and U2093 (N_2093,N_1678,N_1850);
and U2094 (N_2094,N_1579,N_1814);
or U2095 (N_2095,N_1048,N_1627);
or U2096 (N_2096,N_1622,N_1392);
nand U2097 (N_2097,N_1735,N_1294);
xnor U2098 (N_2098,N_1328,N_1078);
or U2099 (N_2099,N_1830,N_1977);
nor U2100 (N_2100,N_1811,N_1715);
or U2101 (N_2101,N_1530,N_1015);
nand U2102 (N_2102,N_1270,N_1615);
or U2103 (N_2103,N_1545,N_1638);
nand U2104 (N_2104,N_1718,N_1509);
and U2105 (N_2105,N_1888,N_1265);
xnor U2106 (N_2106,N_1085,N_1500);
or U2107 (N_2107,N_1961,N_1055);
or U2108 (N_2108,N_1558,N_1998);
xor U2109 (N_2109,N_1881,N_1488);
and U2110 (N_2110,N_1976,N_1021);
xor U2111 (N_2111,N_1113,N_1798);
xnor U2112 (N_2112,N_1648,N_1207);
and U2113 (N_2113,N_1326,N_1823);
xor U2114 (N_2114,N_1248,N_1070);
xnor U2115 (N_2115,N_1962,N_1919);
nand U2116 (N_2116,N_1610,N_1629);
nand U2117 (N_2117,N_1336,N_1502);
nand U2118 (N_2118,N_1251,N_1342);
xor U2119 (N_2119,N_1471,N_1107);
xnor U2120 (N_2120,N_1087,N_1145);
and U2121 (N_2121,N_1525,N_1533);
nor U2122 (N_2122,N_1833,N_1659);
nand U2123 (N_2123,N_1835,N_1019);
nor U2124 (N_2124,N_1063,N_1982);
nand U2125 (N_2125,N_1598,N_1543);
or U2126 (N_2126,N_1122,N_1517);
and U2127 (N_2127,N_1035,N_1356);
xnor U2128 (N_2128,N_1020,N_1050);
nand U2129 (N_2129,N_1876,N_1540);
nand U2130 (N_2130,N_1424,N_1674);
or U2131 (N_2131,N_1481,N_1354);
nand U2132 (N_2132,N_1566,N_1438);
xnor U2133 (N_2133,N_1650,N_1394);
nand U2134 (N_2134,N_1849,N_1210);
nand U2135 (N_2135,N_1806,N_1219);
xnor U2136 (N_2136,N_1370,N_1762);
nand U2137 (N_2137,N_1140,N_1769);
and U2138 (N_2138,N_1421,N_1550);
nor U2139 (N_2139,N_1005,N_1194);
nor U2140 (N_2140,N_1596,N_1202);
or U2141 (N_2141,N_1920,N_1902);
or U2142 (N_2142,N_1966,N_1295);
nor U2143 (N_2143,N_1293,N_1817);
or U2144 (N_2144,N_1828,N_1747);
xnor U2145 (N_2145,N_1765,N_1428);
nor U2146 (N_2146,N_1211,N_1446);
nand U2147 (N_2147,N_1376,N_1466);
xnor U2148 (N_2148,N_1227,N_1016);
xnor U2149 (N_2149,N_1166,N_1246);
xor U2150 (N_2150,N_1869,N_1486);
nand U2151 (N_2151,N_1425,N_1694);
or U2152 (N_2152,N_1126,N_1427);
nand U2153 (N_2153,N_1268,N_1411);
xor U2154 (N_2154,N_1625,N_1988);
nand U2155 (N_2155,N_1973,N_1741);
and U2156 (N_2156,N_1034,N_1031);
nand U2157 (N_2157,N_1174,N_1853);
and U2158 (N_2158,N_1101,N_1436);
or U2159 (N_2159,N_1681,N_1737);
and U2160 (N_2160,N_1721,N_1775);
xnor U2161 (N_2161,N_1809,N_1144);
nor U2162 (N_2162,N_1926,N_1584);
nand U2163 (N_2163,N_1442,N_1928);
nand U2164 (N_2164,N_1794,N_1275);
nand U2165 (N_2165,N_1467,N_1758);
nor U2166 (N_2166,N_1535,N_1118);
nand U2167 (N_2167,N_1386,N_1628);
nand U2168 (N_2168,N_1944,N_1801);
nor U2169 (N_2169,N_1997,N_1167);
and U2170 (N_2170,N_1760,N_1770);
and U2171 (N_2171,N_1404,N_1521);
xnor U2172 (N_2172,N_1751,N_1150);
xor U2173 (N_2173,N_1355,N_1951);
xnor U2174 (N_2174,N_1670,N_1877);
and U2175 (N_2175,N_1420,N_1135);
or U2176 (N_2176,N_1130,N_1041);
and U2177 (N_2177,N_1164,N_1831);
nor U2178 (N_2178,N_1706,N_1387);
and U2179 (N_2179,N_1585,N_1560);
or U2180 (N_2180,N_1633,N_1946);
and U2181 (N_2181,N_1125,N_1325);
and U2182 (N_2182,N_1190,N_1789);
and U2183 (N_2183,N_1094,N_1539);
nor U2184 (N_2184,N_1066,N_1698);
and U2185 (N_2185,N_1708,N_1027);
nand U2186 (N_2186,N_1221,N_1730);
and U2187 (N_2187,N_1273,N_1337);
nand U2188 (N_2188,N_1634,N_1463);
nor U2189 (N_2189,N_1030,N_1645);
nor U2190 (N_2190,N_1567,N_1006);
or U2191 (N_2191,N_1316,N_1423);
xnor U2192 (N_2192,N_1360,N_1091);
and U2193 (N_2193,N_1851,N_1260);
xor U2194 (N_2194,N_1124,N_1080);
and U2195 (N_2195,N_1981,N_1683);
nor U2196 (N_2196,N_1037,N_1954);
nor U2197 (N_2197,N_1026,N_1152);
nor U2198 (N_2198,N_1192,N_1686);
nand U2199 (N_2199,N_1435,N_1395);
or U2200 (N_2200,N_1315,N_1723);
xor U2201 (N_2201,N_1253,N_1477);
nor U2202 (N_2202,N_1661,N_1082);
nor U2203 (N_2203,N_1987,N_1254);
nand U2204 (N_2204,N_1366,N_1682);
or U2205 (N_2205,N_1991,N_1972);
or U2206 (N_2206,N_1465,N_1215);
nand U2207 (N_2207,N_1515,N_1652);
nand U2208 (N_2208,N_1478,N_1878);
nand U2209 (N_2209,N_1099,N_1267);
or U2210 (N_2210,N_1587,N_1909);
nor U2211 (N_2211,N_1918,N_1018);
nor U2212 (N_2212,N_1680,N_1974);
nand U2213 (N_2213,N_1292,N_1937);
nor U2214 (N_2214,N_1095,N_1288);
nand U2215 (N_2215,N_1198,N_1565);
or U2216 (N_2216,N_1511,N_1434);
xnor U2217 (N_2217,N_1474,N_1017);
and U2218 (N_2218,N_1940,N_1984);
and U2219 (N_2219,N_1872,N_1603);
or U2220 (N_2220,N_1262,N_1939);
nor U2221 (N_2221,N_1583,N_1179);
and U2222 (N_2222,N_1884,N_1609);
nor U2223 (N_2223,N_1599,N_1802);
nand U2224 (N_2224,N_1359,N_1241);
nor U2225 (N_2225,N_1547,N_1999);
xnor U2226 (N_2226,N_1989,N_1514);
or U2227 (N_2227,N_1748,N_1155);
nand U2228 (N_2228,N_1952,N_1405);
or U2229 (N_2229,N_1052,N_1549);
or U2230 (N_2230,N_1679,N_1600);
nand U2231 (N_2231,N_1572,N_1597);
nor U2232 (N_2232,N_1757,N_1464);
and U2233 (N_2233,N_1391,N_1303);
xor U2234 (N_2234,N_1009,N_1636);
xnor U2235 (N_2235,N_1403,N_1595);
nor U2236 (N_2236,N_1007,N_1922);
nor U2237 (N_2237,N_1322,N_1942);
nand U2238 (N_2238,N_1556,N_1384);
xor U2239 (N_2239,N_1308,N_1120);
or U2240 (N_2240,N_1283,N_1978);
nand U2241 (N_2241,N_1943,N_1722);
nand U2242 (N_2242,N_1196,N_1257);
nor U2243 (N_2243,N_1361,N_1690);
xor U2244 (N_2244,N_1903,N_1496);
xor U2245 (N_2245,N_1908,N_1519);
nand U2246 (N_2246,N_1346,N_1559);
xor U2247 (N_2247,N_1582,N_1104);
and U2248 (N_2248,N_1898,N_1739);
nand U2249 (N_2249,N_1818,N_1297);
nor U2250 (N_2250,N_1750,N_1534);
or U2251 (N_2251,N_1693,N_1239);
nor U2252 (N_2252,N_1081,N_1284);
and U2253 (N_2253,N_1890,N_1378);
nand U2254 (N_2254,N_1651,N_1456);
xnor U2255 (N_2255,N_1971,N_1777);
xor U2256 (N_2256,N_1287,N_1604);
nor U2257 (N_2257,N_1588,N_1230);
nor U2258 (N_2258,N_1994,N_1829);
nor U2259 (N_2259,N_1123,N_1495);
nand U2260 (N_2260,N_1518,N_1183);
or U2261 (N_2261,N_1317,N_1800);
nor U2262 (N_2262,N_1282,N_1749);
nor U2263 (N_2263,N_1385,N_1377);
and U2264 (N_2264,N_1350,N_1397);
and U2265 (N_2265,N_1313,N_1779);
nand U2266 (N_2266,N_1119,N_1362);
nand U2267 (N_2267,N_1068,N_1764);
nor U2268 (N_2268,N_1774,N_1677);
and U2269 (N_2269,N_1444,N_1056);
nand U2270 (N_2270,N_1932,N_1357);
or U2271 (N_2271,N_1812,N_1508);
nor U2272 (N_2272,N_1147,N_1437);
nor U2273 (N_2273,N_1834,N_1001);
nand U2274 (N_2274,N_1837,N_1112);
nand U2275 (N_2275,N_1036,N_1004);
nor U2276 (N_2276,N_1225,N_1223);
nor U2277 (N_2277,N_1503,N_1605);
and U2278 (N_2278,N_1199,N_1146);
or U2279 (N_2279,N_1069,N_1970);
or U2280 (N_2280,N_1745,N_1963);
nor U2281 (N_2281,N_1793,N_1980);
xnor U2282 (N_2282,N_1422,N_1746);
and U2283 (N_2283,N_1771,N_1624);
nor U2284 (N_2284,N_1149,N_1431);
xnor U2285 (N_2285,N_1923,N_1458);
or U2286 (N_2286,N_1235,N_1343);
and U2287 (N_2287,N_1426,N_1957);
nand U2288 (N_2288,N_1057,N_1375);
and U2289 (N_2289,N_1204,N_1412);
xnor U2290 (N_2290,N_1717,N_1162);
nor U2291 (N_2291,N_1701,N_1720);
and U2292 (N_2292,N_1912,N_1485);
or U2293 (N_2293,N_1046,N_1059);
and U2294 (N_2294,N_1138,N_1573);
nor U2295 (N_2295,N_1945,N_1430);
xor U2296 (N_2296,N_1896,N_1025);
and U2297 (N_2297,N_1882,N_1347);
nor U2298 (N_2298,N_1177,N_1134);
and U2299 (N_2299,N_1541,N_1381);
xor U2300 (N_2300,N_1666,N_1079);
and U2301 (N_2301,N_1186,N_1924);
and U2302 (N_2302,N_1941,N_1416);
xnor U2303 (N_2303,N_1290,N_1409);
and U2304 (N_2304,N_1374,N_1839);
nor U2305 (N_2305,N_1506,N_1040);
and U2306 (N_2306,N_1843,N_1011);
and U2307 (N_2307,N_1894,N_1537);
xor U2308 (N_2308,N_1470,N_1880);
and U2309 (N_2309,N_1242,N_1327);
or U2310 (N_2310,N_1526,N_1191);
and U2311 (N_2311,N_1848,N_1983);
or U2312 (N_2312,N_1528,N_1187);
or U2313 (N_2313,N_1838,N_1305);
nor U2314 (N_2314,N_1563,N_1889);
and U2315 (N_2315,N_1178,N_1238);
and U2316 (N_2316,N_1484,N_1531);
nor U2317 (N_2317,N_1274,N_1269);
or U2318 (N_2318,N_1200,N_1554);
nand U2319 (N_2319,N_1333,N_1568);
nand U2320 (N_2320,N_1696,N_1208);
xor U2321 (N_2321,N_1105,N_1618);
or U2322 (N_2322,N_1473,N_1711);
xor U2323 (N_2323,N_1784,N_1688);
xor U2324 (N_2324,N_1213,N_1345);
xnor U2325 (N_2325,N_1616,N_1921);
and U2326 (N_2326,N_1142,N_1856);
and U2327 (N_2327,N_1813,N_1136);
nand U2328 (N_2328,N_1916,N_1296);
nand U2329 (N_2329,N_1712,N_1259);
nand U2330 (N_2330,N_1348,N_1805);
xor U2331 (N_2331,N_1157,N_1959);
nor U2332 (N_2332,N_1781,N_1388);
nand U2333 (N_2333,N_1049,N_1289);
xor U2334 (N_2334,N_1449,N_1642);
nand U2335 (N_2335,N_1447,N_1092);
xnor U2336 (N_2336,N_1867,N_1612);
and U2337 (N_2337,N_1911,N_1490);
xor U2338 (N_2338,N_1538,N_1163);
nor U2339 (N_2339,N_1900,N_1782);
or U2340 (N_2340,N_1154,N_1286);
xor U2341 (N_2341,N_1947,N_1285);
nor U2342 (N_2342,N_1255,N_1448);
xnor U2343 (N_2343,N_1700,N_1826);
xnor U2344 (N_2344,N_1979,N_1591);
nand U2345 (N_2345,N_1062,N_1402);
and U2346 (N_2346,N_1086,N_1546);
or U2347 (N_2347,N_1396,N_1655);
or U2348 (N_2348,N_1188,N_1121);
xnor U2349 (N_2349,N_1433,N_1958);
nand U2350 (N_2350,N_1408,N_1637);
xnor U2351 (N_2351,N_1862,N_1440);
nand U2352 (N_2352,N_1044,N_1457);
and U2353 (N_2353,N_1053,N_1744);
and U2354 (N_2354,N_1459,N_1369);
and U2355 (N_2355,N_1058,N_1886);
and U2356 (N_2356,N_1608,N_1281);
and U2357 (N_2357,N_1324,N_1074);
or U2358 (N_2358,N_1184,N_1816);
xor U2359 (N_2359,N_1352,N_1060);
or U2360 (N_2360,N_1505,N_1258);
xor U2361 (N_2361,N_1948,N_1318);
or U2362 (N_2362,N_1524,N_1586);
xor U2363 (N_2363,N_1562,N_1263);
nor U2364 (N_2364,N_1312,N_1232);
nand U2365 (N_2365,N_1450,N_1047);
xnor U2366 (N_2366,N_1407,N_1868);
xor U2367 (N_2367,N_1787,N_1160);
nor U2368 (N_2368,N_1461,N_1331);
nand U2369 (N_2369,N_1780,N_1854);
or U2370 (N_2370,N_1619,N_1304);
nor U2371 (N_2371,N_1913,N_1930);
xor U2372 (N_2372,N_1233,N_1611);
and U2373 (N_2373,N_1665,N_1899);
xor U2374 (N_2374,N_1761,N_1752);
or U2375 (N_2375,N_1858,N_1754);
and U2376 (N_2376,N_1076,N_1161);
nor U2377 (N_2377,N_1189,N_1875);
nand U2378 (N_2378,N_1569,N_1910);
or U2379 (N_2379,N_1330,N_1593);
and U2380 (N_2380,N_1716,N_1702);
xnor U2381 (N_2381,N_1879,N_1256);
nor U2382 (N_2382,N_1692,N_1931);
or U2383 (N_2383,N_1580,N_1236);
xnor U2384 (N_2384,N_1892,N_1786);
nor U2385 (N_2385,N_1512,N_1731);
and U2386 (N_2386,N_1493,N_1578);
and U2387 (N_2387,N_1601,N_1516);
or U2388 (N_2388,N_1719,N_1307);
nor U2389 (N_2389,N_1299,N_1483);
or U2390 (N_2390,N_1117,N_1220);
and U2391 (N_2391,N_1887,N_1697);
nor U2392 (N_2392,N_1454,N_1000);
or U2393 (N_2393,N_1660,N_1349);
nor U2394 (N_2394,N_1685,N_1657);
xor U2395 (N_2395,N_1960,N_1042);
or U2396 (N_2396,N_1280,N_1231);
or U2397 (N_2397,N_1226,N_1158);
nor U2398 (N_2398,N_1414,N_1100);
nor U2399 (N_2399,N_1819,N_1024);
and U2400 (N_2400,N_1536,N_1925);
nand U2401 (N_2401,N_1180,N_1309);
xor U2402 (N_2402,N_1229,N_1571);
nor U2403 (N_2403,N_1276,N_1106);
or U2404 (N_2404,N_1243,N_1607);
or U2405 (N_2405,N_1795,N_1399);
or U2406 (N_2406,N_1492,N_1874);
nor U2407 (N_2407,N_1072,N_1993);
nand U2408 (N_2408,N_1901,N_1763);
and U2409 (N_2409,N_1852,N_1432);
xor U2410 (N_2410,N_1382,N_1339);
and U2411 (N_2411,N_1728,N_1209);
xnor U2412 (N_2412,N_1033,N_1441);
nand U2413 (N_2413,N_1491,N_1003);
nand U2414 (N_2414,N_1687,N_1906);
nand U2415 (N_2415,N_1310,N_1201);
or U2416 (N_2416,N_1410,N_1451);
xor U2417 (N_2417,N_1240,N_1245);
and U2418 (N_2418,N_1090,N_1319);
xor U2419 (N_2419,N_1132,N_1626);
nand U2420 (N_2420,N_1614,N_1415);
and U2421 (N_2421,N_1808,N_1043);
xor U2422 (N_2422,N_1153,N_1743);
xnor U2423 (N_2423,N_1732,N_1742);
nand U2424 (N_2424,N_1277,N_1128);
xnor U2425 (N_2425,N_1788,N_1320);
nor U2426 (N_2426,N_1482,N_1799);
and U2427 (N_2427,N_1553,N_1663);
nand U2428 (N_2428,N_1002,N_1825);
nor U2429 (N_2429,N_1933,N_1606);
and U2430 (N_2430,N_1967,N_1185);
xnor U2431 (N_2431,N_1841,N_1479);
nor U2432 (N_2432,N_1429,N_1494);
nor U2433 (N_2433,N_1975,N_1592);
nor U2434 (N_2434,N_1175,N_1298);
nand U2435 (N_2435,N_1755,N_1797);
or U2436 (N_2436,N_1321,N_1840);
nor U2437 (N_2437,N_1542,N_1497);
nor U2438 (N_2438,N_1740,N_1406);
or U2439 (N_2439,N_1968,N_1012);
xnor U2440 (N_2440,N_1796,N_1893);
nand U2441 (N_2441,N_1261,N_1551);
or U2442 (N_2442,N_1753,N_1859);
nand U2443 (N_2443,N_1904,N_1418);
or U2444 (N_2444,N_1364,N_1114);
and U2445 (N_2445,N_1065,N_1847);
xor U2446 (N_2446,N_1367,N_1472);
nor U2447 (N_2447,N_1857,N_1045);
nand U2448 (N_2448,N_1096,N_1108);
xnor U2449 (N_2449,N_1365,N_1513);
nand U2450 (N_2450,N_1667,N_1662);
or U2451 (N_2451,N_1897,N_1703);
or U2452 (N_2452,N_1234,N_1639);
and U2453 (N_2453,N_1372,N_1815);
nor U2454 (N_2454,N_1172,N_1644);
or U2455 (N_2455,N_1699,N_1822);
or U2456 (N_2456,N_1398,N_1314);
nor U2457 (N_2457,N_1845,N_1064);
nor U2458 (N_2458,N_1301,N_1934);
and U2459 (N_2459,N_1083,N_1552);
nand U2460 (N_2460,N_1759,N_1654);
or U2461 (N_2461,N_1039,N_1165);
xor U2462 (N_2462,N_1206,N_1766);
nor U2463 (N_2463,N_1768,N_1995);
xnor U2464 (N_2464,N_1480,N_1827);
nor U2465 (N_2465,N_1557,N_1820);
nor U2466 (N_2466,N_1462,N_1266);
and U2467 (N_2467,N_1071,N_1949);
nand U2468 (N_2468,N_1602,N_1724);
xor U2469 (N_2469,N_1992,N_1938);
nand U2470 (N_2470,N_1102,N_1713);
xor U2471 (N_2471,N_1129,N_1054);
nor U2472 (N_2472,N_1990,N_1733);
nand U2473 (N_2473,N_1927,N_1109);
xnor U2474 (N_2474,N_1620,N_1419);
or U2475 (N_2475,N_1725,N_1646);
or U2476 (N_2476,N_1088,N_1658);
xor U2477 (N_2477,N_1865,N_1917);
xnor U2478 (N_2478,N_1334,N_1576);
and U2479 (N_2479,N_1413,N_1783);
nor U2480 (N_2480,N_1332,N_1329);
and U2481 (N_2481,N_1767,N_1623);
and U2482 (N_2482,N_1532,N_1051);
nand U2483 (N_2483,N_1249,N_1870);
xor U2484 (N_2484,N_1077,N_1156);
and U2485 (N_2485,N_1351,N_1985);
and U2486 (N_2486,N_1173,N_1363);
xnor U2487 (N_2487,N_1671,N_1621);
xnor U2488 (N_2488,N_1691,N_1340);
and U2489 (N_2489,N_1676,N_1965);
and U2490 (N_2490,N_1032,N_1589);
nand U2491 (N_2491,N_1964,N_1008);
or U2492 (N_2492,N_1631,N_1522);
nor U2493 (N_2493,N_1061,N_1439);
nand U2494 (N_2494,N_1272,N_1804);
and U2495 (N_2495,N_1469,N_1487);
nand U2496 (N_2496,N_1131,N_1647);
or U2497 (N_2497,N_1371,N_1498);
and U2498 (N_2498,N_1527,N_1726);
and U2499 (N_2499,N_1014,N_1821);
nand U2500 (N_2500,N_1314,N_1762);
or U2501 (N_2501,N_1474,N_1129);
or U2502 (N_2502,N_1747,N_1129);
and U2503 (N_2503,N_1153,N_1943);
nor U2504 (N_2504,N_1774,N_1952);
nand U2505 (N_2505,N_1403,N_1384);
nor U2506 (N_2506,N_1109,N_1372);
xnor U2507 (N_2507,N_1566,N_1755);
nor U2508 (N_2508,N_1585,N_1679);
xnor U2509 (N_2509,N_1315,N_1545);
xnor U2510 (N_2510,N_1107,N_1781);
and U2511 (N_2511,N_1862,N_1512);
nor U2512 (N_2512,N_1213,N_1401);
nand U2513 (N_2513,N_1819,N_1499);
nand U2514 (N_2514,N_1901,N_1716);
and U2515 (N_2515,N_1638,N_1446);
xnor U2516 (N_2516,N_1058,N_1613);
nand U2517 (N_2517,N_1623,N_1515);
nand U2518 (N_2518,N_1096,N_1251);
nor U2519 (N_2519,N_1125,N_1533);
or U2520 (N_2520,N_1257,N_1268);
or U2521 (N_2521,N_1321,N_1667);
nor U2522 (N_2522,N_1551,N_1631);
or U2523 (N_2523,N_1911,N_1235);
or U2524 (N_2524,N_1322,N_1439);
and U2525 (N_2525,N_1656,N_1324);
xor U2526 (N_2526,N_1451,N_1270);
or U2527 (N_2527,N_1961,N_1745);
xnor U2528 (N_2528,N_1508,N_1200);
xnor U2529 (N_2529,N_1257,N_1314);
or U2530 (N_2530,N_1877,N_1342);
xnor U2531 (N_2531,N_1497,N_1071);
or U2532 (N_2532,N_1701,N_1323);
xor U2533 (N_2533,N_1755,N_1713);
nand U2534 (N_2534,N_1230,N_1291);
or U2535 (N_2535,N_1829,N_1197);
xor U2536 (N_2536,N_1096,N_1870);
nand U2537 (N_2537,N_1993,N_1466);
nand U2538 (N_2538,N_1447,N_1431);
nand U2539 (N_2539,N_1376,N_1143);
and U2540 (N_2540,N_1046,N_1387);
or U2541 (N_2541,N_1433,N_1878);
and U2542 (N_2542,N_1771,N_1953);
xnor U2543 (N_2543,N_1151,N_1814);
and U2544 (N_2544,N_1003,N_1256);
nand U2545 (N_2545,N_1792,N_1324);
or U2546 (N_2546,N_1785,N_1868);
xor U2547 (N_2547,N_1628,N_1645);
and U2548 (N_2548,N_1466,N_1559);
nand U2549 (N_2549,N_1250,N_1762);
nand U2550 (N_2550,N_1547,N_1797);
or U2551 (N_2551,N_1186,N_1922);
xor U2552 (N_2552,N_1177,N_1474);
nor U2553 (N_2553,N_1188,N_1816);
nor U2554 (N_2554,N_1937,N_1161);
xor U2555 (N_2555,N_1719,N_1371);
and U2556 (N_2556,N_1280,N_1805);
and U2557 (N_2557,N_1332,N_1290);
nand U2558 (N_2558,N_1711,N_1567);
or U2559 (N_2559,N_1755,N_1526);
nand U2560 (N_2560,N_1461,N_1032);
nand U2561 (N_2561,N_1763,N_1565);
nand U2562 (N_2562,N_1080,N_1981);
nand U2563 (N_2563,N_1630,N_1494);
and U2564 (N_2564,N_1897,N_1695);
or U2565 (N_2565,N_1085,N_1270);
and U2566 (N_2566,N_1818,N_1244);
nor U2567 (N_2567,N_1281,N_1609);
or U2568 (N_2568,N_1613,N_1566);
xnor U2569 (N_2569,N_1441,N_1297);
nor U2570 (N_2570,N_1328,N_1049);
nand U2571 (N_2571,N_1998,N_1905);
and U2572 (N_2572,N_1378,N_1823);
nand U2573 (N_2573,N_1349,N_1526);
and U2574 (N_2574,N_1898,N_1585);
xnor U2575 (N_2575,N_1981,N_1267);
nand U2576 (N_2576,N_1177,N_1702);
nand U2577 (N_2577,N_1089,N_1682);
nor U2578 (N_2578,N_1511,N_1973);
nand U2579 (N_2579,N_1343,N_1138);
and U2580 (N_2580,N_1354,N_1737);
nor U2581 (N_2581,N_1174,N_1373);
or U2582 (N_2582,N_1967,N_1437);
nand U2583 (N_2583,N_1560,N_1596);
nand U2584 (N_2584,N_1159,N_1912);
or U2585 (N_2585,N_1857,N_1195);
and U2586 (N_2586,N_1353,N_1278);
nor U2587 (N_2587,N_1324,N_1759);
xor U2588 (N_2588,N_1548,N_1260);
nor U2589 (N_2589,N_1465,N_1801);
nor U2590 (N_2590,N_1496,N_1776);
or U2591 (N_2591,N_1348,N_1255);
and U2592 (N_2592,N_1467,N_1956);
nand U2593 (N_2593,N_1147,N_1228);
nand U2594 (N_2594,N_1067,N_1276);
and U2595 (N_2595,N_1178,N_1564);
and U2596 (N_2596,N_1111,N_1485);
or U2597 (N_2597,N_1974,N_1830);
and U2598 (N_2598,N_1185,N_1082);
nand U2599 (N_2599,N_1735,N_1259);
nor U2600 (N_2600,N_1443,N_1100);
and U2601 (N_2601,N_1717,N_1912);
nand U2602 (N_2602,N_1136,N_1147);
nor U2603 (N_2603,N_1373,N_1470);
nor U2604 (N_2604,N_1650,N_1236);
nor U2605 (N_2605,N_1555,N_1301);
nand U2606 (N_2606,N_1200,N_1627);
xnor U2607 (N_2607,N_1650,N_1497);
or U2608 (N_2608,N_1880,N_1153);
nand U2609 (N_2609,N_1695,N_1928);
nor U2610 (N_2610,N_1914,N_1557);
or U2611 (N_2611,N_1742,N_1698);
nand U2612 (N_2612,N_1497,N_1151);
nand U2613 (N_2613,N_1172,N_1119);
or U2614 (N_2614,N_1383,N_1967);
and U2615 (N_2615,N_1218,N_1635);
nand U2616 (N_2616,N_1646,N_1827);
nor U2617 (N_2617,N_1219,N_1159);
nand U2618 (N_2618,N_1632,N_1374);
nor U2619 (N_2619,N_1275,N_1227);
or U2620 (N_2620,N_1862,N_1200);
or U2621 (N_2621,N_1463,N_1095);
nand U2622 (N_2622,N_1691,N_1236);
or U2623 (N_2623,N_1111,N_1009);
and U2624 (N_2624,N_1119,N_1019);
or U2625 (N_2625,N_1009,N_1586);
or U2626 (N_2626,N_1059,N_1523);
nor U2627 (N_2627,N_1563,N_1930);
and U2628 (N_2628,N_1353,N_1654);
or U2629 (N_2629,N_1641,N_1406);
nor U2630 (N_2630,N_1426,N_1208);
xnor U2631 (N_2631,N_1550,N_1152);
or U2632 (N_2632,N_1046,N_1579);
xnor U2633 (N_2633,N_1010,N_1420);
and U2634 (N_2634,N_1626,N_1745);
nor U2635 (N_2635,N_1449,N_1007);
or U2636 (N_2636,N_1536,N_1302);
xor U2637 (N_2637,N_1982,N_1837);
nand U2638 (N_2638,N_1809,N_1580);
or U2639 (N_2639,N_1856,N_1740);
and U2640 (N_2640,N_1709,N_1537);
nand U2641 (N_2641,N_1248,N_1175);
nor U2642 (N_2642,N_1045,N_1102);
nor U2643 (N_2643,N_1342,N_1125);
xor U2644 (N_2644,N_1128,N_1777);
nor U2645 (N_2645,N_1411,N_1012);
nor U2646 (N_2646,N_1125,N_1002);
or U2647 (N_2647,N_1661,N_1330);
or U2648 (N_2648,N_1432,N_1014);
nand U2649 (N_2649,N_1509,N_1875);
nor U2650 (N_2650,N_1734,N_1262);
nor U2651 (N_2651,N_1714,N_1389);
nor U2652 (N_2652,N_1937,N_1963);
nand U2653 (N_2653,N_1406,N_1927);
xor U2654 (N_2654,N_1892,N_1535);
nor U2655 (N_2655,N_1832,N_1906);
or U2656 (N_2656,N_1780,N_1788);
nor U2657 (N_2657,N_1692,N_1278);
xor U2658 (N_2658,N_1686,N_1363);
and U2659 (N_2659,N_1694,N_1554);
and U2660 (N_2660,N_1254,N_1759);
nor U2661 (N_2661,N_1991,N_1732);
or U2662 (N_2662,N_1685,N_1941);
and U2663 (N_2663,N_1885,N_1525);
xnor U2664 (N_2664,N_1820,N_1482);
nand U2665 (N_2665,N_1992,N_1538);
nor U2666 (N_2666,N_1451,N_1379);
or U2667 (N_2667,N_1147,N_1964);
and U2668 (N_2668,N_1899,N_1121);
nand U2669 (N_2669,N_1621,N_1609);
nand U2670 (N_2670,N_1973,N_1542);
xor U2671 (N_2671,N_1044,N_1040);
or U2672 (N_2672,N_1949,N_1207);
and U2673 (N_2673,N_1811,N_1939);
and U2674 (N_2674,N_1834,N_1888);
xnor U2675 (N_2675,N_1582,N_1734);
nand U2676 (N_2676,N_1498,N_1292);
or U2677 (N_2677,N_1504,N_1466);
nand U2678 (N_2678,N_1883,N_1354);
nor U2679 (N_2679,N_1612,N_1649);
nor U2680 (N_2680,N_1894,N_1375);
or U2681 (N_2681,N_1792,N_1395);
nor U2682 (N_2682,N_1250,N_1969);
nand U2683 (N_2683,N_1510,N_1119);
nand U2684 (N_2684,N_1423,N_1637);
or U2685 (N_2685,N_1325,N_1097);
nor U2686 (N_2686,N_1033,N_1261);
xor U2687 (N_2687,N_1749,N_1878);
nor U2688 (N_2688,N_1016,N_1590);
and U2689 (N_2689,N_1318,N_1525);
or U2690 (N_2690,N_1860,N_1486);
xnor U2691 (N_2691,N_1814,N_1613);
nor U2692 (N_2692,N_1001,N_1579);
xnor U2693 (N_2693,N_1619,N_1073);
or U2694 (N_2694,N_1918,N_1082);
nor U2695 (N_2695,N_1465,N_1278);
xnor U2696 (N_2696,N_1138,N_1699);
nand U2697 (N_2697,N_1971,N_1021);
nand U2698 (N_2698,N_1574,N_1889);
or U2699 (N_2699,N_1395,N_1827);
nor U2700 (N_2700,N_1580,N_1149);
xnor U2701 (N_2701,N_1138,N_1971);
and U2702 (N_2702,N_1733,N_1735);
and U2703 (N_2703,N_1078,N_1314);
nand U2704 (N_2704,N_1858,N_1390);
nor U2705 (N_2705,N_1725,N_1811);
nand U2706 (N_2706,N_1002,N_1588);
nor U2707 (N_2707,N_1183,N_1656);
nand U2708 (N_2708,N_1161,N_1528);
nand U2709 (N_2709,N_1757,N_1459);
and U2710 (N_2710,N_1983,N_1404);
xor U2711 (N_2711,N_1492,N_1604);
nor U2712 (N_2712,N_1037,N_1805);
nor U2713 (N_2713,N_1168,N_1155);
xnor U2714 (N_2714,N_1746,N_1273);
and U2715 (N_2715,N_1191,N_1555);
nor U2716 (N_2716,N_1673,N_1005);
and U2717 (N_2717,N_1536,N_1350);
nand U2718 (N_2718,N_1694,N_1195);
and U2719 (N_2719,N_1435,N_1198);
or U2720 (N_2720,N_1043,N_1611);
nand U2721 (N_2721,N_1511,N_1397);
nor U2722 (N_2722,N_1071,N_1207);
nor U2723 (N_2723,N_1070,N_1378);
and U2724 (N_2724,N_1518,N_1466);
nand U2725 (N_2725,N_1207,N_1048);
or U2726 (N_2726,N_1098,N_1609);
nand U2727 (N_2727,N_1807,N_1547);
xor U2728 (N_2728,N_1130,N_1553);
nand U2729 (N_2729,N_1426,N_1920);
or U2730 (N_2730,N_1422,N_1671);
xor U2731 (N_2731,N_1522,N_1271);
and U2732 (N_2732,N_1759,N_1148);
and U2733 (N_2733,N_1771,N_1975);
nand U2734 (N_2734,N_1557,N_1246);
xor U2735 (N_2735,N_1434,N_1911);
xor U2736 (N_2736,N_1798,N_1667);
nand U2737 (N_2737,N_1710,N_1972);
nor U2738 (N_2738,N_1937,N_1593);
nor U2739 (N_2739,N_1883,N_1161);
or U2740 (N_2740,N_1039,N_1465);
nor U2741 (N_2741,N_1168,N_1336);
or U2742 (N_2742,N_1382,N_1777);
nand U2743 (N_2743,N_1205,N_1287);
nor U2744 (N_2744,N_1547,N_1022);
xnor U2745 (N_2745,N_1346,N_1820);
xnor U2746 (N_2746,N_1039,N_1607);
nand U2747 (N_2747,N_1317,N_1003);
nand U2748 (N_2748,N_1259,N_1410);
nor U2749 (N_2749,N_1240,N_1084);
or U2750 (N_2750,N_1917,N_1673);
nand U2751 (N_2751,N_1189,N_1459);
or U2752 (N_2752,N_1718,N_1692);
nor U2753 (N_2753,N_1434,N_1861);
and U2754 (N_2754,N_1413,N_1375);
or U2755 (N_2755,N_1309,N_1175);
nor U2756 (N_2756,N_1541,N_1621);
nand U2757 (N_2757,N_1206,N_1411);
and U2758 (N_2758,N_1482,N_1617);
and U2759 (N_2759,N_1822,N_1932);
nand U2760 (N_2760,N_1406,N_1717);
and U2761 (N_2761,N_1647,N_1758);
nand U2762 (N_2762,N_1971,N_1712);
or U2763 (N_2763,N_1888,N_1096);
or U2764 (N_2764,N_1890,N_1501);
nor U2765 (N_2765,N_1927,N_1130);
xor U2766 (N_2766,N_1709,N_1873);
nor U2767 (N_2767,N_1351,N_1651);
xnor U2768 (N_2768,N_1442,N_1822);
and U2769 (N_2769,N_1607,N_1236);
or U2770 (N_2770,N_1507,N_1123);
and U2771 (N_2771,N_1369,N_1030);
xor U2772 (N_2772,N_1465,N_1844);
nand U2773 (N_2773,N_1605,N_1463);
or U2774 (N_2774,N_1941,N_1254);
xnor U2775 (N_2775,N_1530,N_1693);
nor U2776 (N_2776,N_1082,N_1752);
and U2777 (N_2777,N_1188,N_1679);
and U2778 (N_2778,N_1195,N_1054);
or U2779 (N_2779,N_1412,N_1974);
xnor U2780 (N_2780,N_1385,N_1522);
or U2781 (N_2781,N_1486,N_1626);
nor U2782 (N_2782,N_1368,N_1857);
nand U2783 (N_2783,N_1383,N_1416);
or U2784 (N_2784,N_1031,N_1878);
nand U2785 (N_2785,N_1091,N_1571);
and U2786 (N_2786,N_1807,N_1863);
or U2787 (N_2787,N_1146,N_1282);
or U2788 (N_2788,N_1594,N_1705);
and U2789 (N_2789,N_1729,N_1654);
nor U2790 (N_2790,N_1223,N_1986);
and U2791 (N_2791,N_1224,N_1356);
nor U2792 (N_2792,N_1431,N_1947);
xnor U2793 (N_2793,N_1125,N_1670);
nand U2794 (N_2794,N_1234,N_1460);
and U2795 (N_2795,N_1146,N_1231);
or U2796 (N_2796,N_1971,N_1136);
nand U2797 (N_2797,N_1213,N_1025);
nor U2798 (N_2798,N_1081,N_1970);
and U2799 (N_2799,N_1931,N_1081);
nand U2800 (N_2800,N_1410,N_1272);
nand U2801 (N_2801,N_1072,N_1938);
nor U2802 (N_2802,N_1577,N_1100);
nand U2803 (N_2803,N_1622,N_1542);
nand U2804 (N_2804,N_1567,N_1629);
xnor U2805 (N_2805,N_1013,N_1602);
nand U2806 (N_2806,N_1283,N_1361);
and U2807 (N_2807,N_1111,N_1294);
xor U2808 (N_2808,N_1902,N_1734);
and U2809 (N_2809,N_1501,N_1608);
and U2810 (N_2810,N_1838,N_1324);
xnor U2811 (N_2811,N_1715,N_1565);
nand U2812 (N_2812,N_1722,N_1028);
nor U2813 (N_2813,N_1951,N_1400);
nor U2814 (N_2814,N_1535,N_1456);
and U2815 (N_2815,N_1528,N_1020);
nand U2816 (N_2816,N_1385,N_1357);
xor U2817 (N_2817,N_1513,N_1643);
nand U2818 (N_2818,N_1477,N_1252);
or U2819 (N_2819,N_1477,N_1804);
nand U2820 (N_2820,N_1185,N_1958);
or U2821 (N_2821,N_1200,N_1923);
and U2822 (N_2822,N_1582,N_1636);
and U2823 (N_2823,N_1007,N_1422);
nor U2824 (N_2824,N_1270,N_1088);
and U2825 (N_2825,N_1135,N_1667);
and U2826 (N_2826,N_1232,N_1635);
or U2827 (N_2827,N_1189,N_1873);
nand U2828 (N_2828,N_1259,N_1175);
nor U2829 (N_2829,N_1453,N_1411);
or U2830 (N_2830,N_1596,N_1715);
or U2831 (N_2831,N_1824,N_1275);
nor U2832 (N_2832,N_1410,N_1056);
nor U2833 (N_2833,N_1192,N_1491);
nor U2834 (N_2834,N_1357,N_1840);
nand U2835 (N_2835,N_1181,N_1985);
and U2836 (N_2836,N_1201,N_1659);
nor U2837 (N_2837,N_1980,N_1201);
nor U2838 (N_2838,N_1845,N_1052);
nand U2839 (N_2839,N_1558,N_1415);
nor U2840 (N_2840,N_1238,N_1711);
and U2841 (N_2841,N_1974,N_1846);
xnor U2842 (N_2842,N_1789,N_1131);
xor U2843 (N_2843,N_1424,N_1553);
nor U2844 (N_2844,N_1899,N_1760);
nand U2845 (N_2845,N_1523,N_1898);
and U2846 (N_2846,N_1365,N_1674);
nor U2847 (N_2847,N_1234,N_1200);
nor U2848 (N_2848,N_1503,N_1447);
or U2849 (N_2849,N_1873,N_1702);
or U2850 (N_2850,N_1858,N_1585);
and U2851 (N_2851,N_1080,N_1785);
nor U2852 (N_2852,N_1120,N_1424);
nor U2853 (N_2853,N_1124,N_1787);
or U2854 (N_2854,N_1305,N_1454);
and U2855 (N_2855,N_1384,N_1800);
nor U2856 (N_2856,N_1461,N_1104);
and U2857 (N_2857,N_1913,N_1662);
or U2858 (N_2858,N_1807,N_1251);
nand U2859 (N_2859,N_1059,N_1153);
nor U2860 (N_2860,N_1789,N_1924);
xnor U2861 (N_2861,N_1479,N_1760);
nor U2862 (N_2862,N_1856,N_1477);
or U2863 (N_2863,N_1277,N_1611);
xnor U2864 (N_2864,N_1287,N_1452);
and U2865 (N_2865,N_1379,N_1415);
and U2866 (N_2866,N_1826,N_1416);
nor U2867 (N_2867,N_1906,N_1239);
and U2868 (N_2868,N_1374,N_1854);
nand U2869 (N_2869,N_1704,N_1622);
xnor U2870 (N_2870,N_1193,N_1489);
nand U2871 (N_2871,N_1056,N_1822);
and U2872 (N_2872,N_1281,N_1634);
nand U2873 (N_2873,N_1647,N_1249);
nand U2874 (N_2874,N_1060,N_1091);
nor U2875 (N_2875,N_1733,N_1616);
or U2876 (N_2876,N_1472,N_1106);
nand U2877 (N_2877,N_1120,N_1026);
nor U2878 (N_2878,N_1955,N_1245);
nor U2879 (N_2879,N_1630,N_1326);
nor U2880 (N_2880,N_1257,N_1925);
xnor U2881 (N_2881,N_1790,N_1222);
nor U2882 (N_2882,N_1615,N_1243);
or U2883 (N_2883,N_1099,N_1063);
or U2884 (N_2884,N_1940,N_1922);
nand U2885 (N_2885,N_1327,N_1989);
xnor U2886 (N_2886,N_1062,N_1193);
and U2887 (N_2887,N_1071,N_1083);
nand U2888 (N_2888,N_1632,N_1578);
and U2889 (N_2889,N_1236,N_1422);
nand U2890 (N_2890,N_1563,N_1461);
nand U2891 (N_2891,N_1703,N_1494);
or U2892 (N_2892,N_1381,N_1156);
nand U2893 (N_2893,N_1402,N_1450);
nor U2894 (N_2894,N_1824,N_1960);
and U2895 (N_2895,N_1558,N_1621);
and U2896 (N_2896,N_1730,N_1759);
nor U2897 (N_2897,N_1685,N_1210);
nor U2898 (N_2898,N_1810,N_1661);
and U2899 (N_2899,N_1110,N_1958);
and U2900 (N_2900,N_1227,N_1191);
nor U2901 (N_2901,N_1775,N_1643);
nand U2902 (N_2902,N_1456,N_1014);
or U2903 (N_2903,N_1295,N_1110);
xnor U2904 (N_2904,N_1308,N_1410);
nor U2905 (N_2905,N_1593,N_1457);
and U2906 (N_2906,N_1290,N_1122);
nand U2907 (N_2907,N_1850,N_1428);
or U2908 (N_2908,N_1548,N_1526);
nand U2909 (N_2909,N_1152,N_1005);
nor U2910 (N_2910,N_1746,N_1978);
or U2911 (N_2911,N_1040,N_1037);
nand U2912 (N_2912,N_1845,N_1126);
nand U2913 (N_2913,N_1626,N_1298);
xor U2914 (N_2914,N_1185,N_1974);
and U2915 (N_2915,N_1947,N_1421);
nand U2916 (N_2916,N_1827,N_1772);
nor U2917 (N_2917,N_1465,N_1175);
or U2918 (N_2918,N_1975,N_1509);
nor U2919 (N_2919,N_1480,N_1382);
nor U2920 (N_2920,N_1027,N_1433);
nor U2921 (N_2921,N_1145,N_1398);
and U2922 (N_2922,N_1408,N_1130);
or U2923 (N_2923,N_1932,N_1189);
or U2924 (N_2924,N_1090,N_1376);
nor U2925 (N_2925,N_1065,N_1344);
xnor U2926 (N_2926,N_1791,N_1283);
and U2927 (N_2927,N_1750,N_1338);
xor U2928 (N_2928,N_1888,N_1728);
xnor U2929 (N_2929,N_1204,N_1529);
and U2930 (N_2930,N_1256,N_1031);
nand U2931 (N_2931,N_1798,N_1934);
xnor U2932 (N_2932,N_1476,N_1948);
nor U2933 (N_2933,N_1685,N_1377);
nand U2934 (N_2934,N_1137,N_1126);
or U2935 (N_2935,N_1441,N_1160);
xnor U2936 (N_2936,N_1183,N_1590);
xnor U2937 (N_2937,N_1525,N_1373);
xor U2938 (N_2938,N_1018,N_1249);
nand U2939 (N_2939,N_1595,N_1571);
nor U2940 (N_2940,N_1277,N_1325);
or U2941 (N_2941,N_1128,N_1288);
and U2942 (N_2942,N_1688,N_1586);
and U2943 (N_2943,N_1109,N_1284);
nor U2944 (N_2944,N_1111,N_1185);
xnor U2945 (N_2945,N_1629,N_1733);
nand U2946 (N_2946,N_1227,N_1682);
xor U2947 (N_2947,N_1681,N_1016);
nor U2948 (N_2948,N_1961,N_1602);
nor U2949 (N_2949,N_1098,N_1090);
nand U2950 (N_2950,N_1251,N_1280);
or U2951 (N_2951,N_1202,N_1501);
or U2952 (N_2952,N_1868,N_1935);
nor U2953 (N_2953,N_1911,N_1699);
and U2954 (N_2954,N_1202,N_1326);
or U2955 (N_2955,N_1432,N_1331);
and U2956 (N_2956,N_1507,N_1806);
nor U2957 (N_2957,N_1148,N_1898);
nor U2958 (N_2958,N_1262,N_1762);
or U2959 (N_2959,N_1474,N_1134);
and U2960 (N_2960,N_1885,N_1998);
xnor U2961 (N_2961,N_1766,N_1467);
and U2962 (N_2962,N_1069,N_1058);
nor U2963 (N_2963,N_1659,N_1102);
and U2964 (N_2964,N_1097,N_1180);
xor U2965 (N_2965,N_1250,N_1579);
xnor U2966 (N_2966,N_1818,N_1091);
nor U2967 (N_2967,N_1295,N_1972);
xor U2968 (N_2968,N_1693,N_1245);
or U2969 (N_2969,N_1692,N_1706);
nand U2970 (N_2970,N_1827,N_1453);
or U2971 (N_2971,N_1483,N_1335);
or U2972 (N_2972,N_1644,N_1308);
nand U2973 (N_2973,N_1907,N_1695);
or U2974 (N_2974,N_1015,N_1344);
nor U2975 (N_2975,N_1619,N_1248);
nand U2976 (N_2976,N_1490,N_1386);
nand U2977 (N_2977,N_1462,N_1632);
and U2978 (N_2978,N_1276,N_1717);
or U2979 (N_2979,N_1988,N_1141);
or U2980 (N_2980,N_1250,N_1887);
or U2981 (N_2981,N_1896,N_1685);
nor U2982 (N_2982,N_1856,N_1669);
and U2983 (N_2983,N_1161,N_1040);
nor U2984 (N_2984,N_1634,N_1365);
and U2985 (N_2985,N_1277,N_1561);
or U2986 (N_2986,N_1207,N_1900);
nand U2987 (N_2987,N_1540,N_1848);
and U2988 (N_2988,N_1954,N_1205);
xnor U2989 (N_2989,N_1070,N_1236);
nand U2990 (N_2990,N_1026,N_1775);
and U2991 (N_2991,N_1586,N_1308);
and U2992 (N_2992,N_1769,N_1915);
xor U2993 (N_2993,N_1526,N_1978);
or U2994 (N_2994,N_1601,N_1664);
or U2995 (N_2995,N_1514,N_1200);
nand U2996 (N_2996,N_1338,N_1769);
nor U2997 (N_2997,N_1176,N_1221);
or U2998 (N_2998,N_1819,N_1368);
or U2999 (N_2999,N_1478,N_1763);
nand U3000 (N_3000,N_2970,N_2334);
nor U3001 (N_3001,N_2679,N_2883);
xor U3002 (N_3002,N_2676,N_2780);
nor U3003 (N_3003,N_2398,N_2107);
or U3004 (N_3004,N_2853,N_2683);
and U3005 (N_3005,N_2375,N_2696);
nor U3006 (N_3006,N_2370,N_2618);
or U3007 (N_3007,N_2663,N_2130);
or U3008 (N_3008,N_2723,N_2388);
nand U3009 (N_3009,N_2118,N_2405);
xnor U3010 (N_3010,N_2368,N_2600);
and U3011 (N_3011,N_2743,N_2478);
or U3012 (N_3012,N_2872,N_2981);
nand U3013 (N_3013,N_2055,N_2886);
nand U3014 (N_3014,N_2201,N_2988);
and U3015 (N_3015,N_2897,N_2814);
and U3016 (N_3016,N_2012,N_2690);
or U3017 (N_3017,N_2215,N_2893);
xor U3018 (N_3018,N_2868,N_2717);
nor U3019 (N_3019,N_2638,N_2374);
or U3020 (N_3020,N_2385,N_2255);
nor U3021 (N_3021,N_2654,N_2603);
and U3022 (N_3022,N_2517,N_2644);
nand U3023 (N_3023,N_2411,N_2154);
nor U3024 (N_3024,N_2680,N_2533);
nand U3025 (N_3025,N_2586,N_2347);
nor U3026 (N_3026,N_2104,N_2731);
and U3027 (N_3027,N_2135,N_2168);
nor U3028 (N_3028,N_2386,N_2394);
and U3029 (N_3029,N_2968,N_2448);
and U3030 (N_3030,N_2636,N_2254);
nand U3031 (N_3031,N_2585,N_2826);
nor U3032 (N_3032,N_2068,N_2187);
or U3033 (N_3033,N_2662,N_2619);
nand U3034 (N_3034,N_2082,N_2206);
and U3035 (N_3035,N_2588,N_2271);
or U3036 (N_3036,N_2026,N_2319);
nor U3037 (N_3037,N_2125,N_2818);
or U3038 (N_3038,N_2174,N_2983);
nor U3039 (N_3039,N_2067,N_2220);
or U3040 (N_3040,N_2734,N_2544);
nand U3041 (N_3041,N_2178,N_2891);
nor U3042 (N_3042,N_2545,N_2350);
nor U3043 (N_3043,N_2955,N_2623);
nand U3044 (N_3044,N_2035,N_2439);
nor U3045 (N_3045,N_2356,N_2828);
nand U3046 (N_3046,N_2102,N_2904);
nor U3047 (N_3047,N_2792,N_2087);
or U3048 (N_3048,N_2906,N_2628);
nand U3049 (N_3049,N_2438,N_2530);
nor U3050 (N_3050,N_2274,N_2519);
and U3051 (N_3051,N_2236,N_2835);
and U3052 (N_3052,N_2971,N_2993);
and U3053 (N_3053,N_2708,N_2015);
xnor U3054 (N_3054,N_2304,N_2963);
and U3055 (N_3055,N_2570,N_2624);
nor U3056 (N_3056,N_2475,N_2937);
or U3057 (N_3057,N_2337,N_2443);
or U3058 (N_3058,N_2806,N_2090);
nor U3059 (N_3059,N_2435,N_2568);
and U3060 (N_3060,N_2006,N_2101);
nor U3061 (N_3061,N_2562,N_2115);
nor U3062 (N_3062,N_2693,N_2023);
or U3063 (N_3063,N_2414,N_2521);
nand U3064 (N_3064,N_2277,N_2177);
or U3065 (N_3065,N_2343,N_2653);
nand U3066 (N_3066,N_2310,N_2261);
nand U3067 (N_3067,N_2445,N_2563);
xor U3068 (N_3068,N_2045,N_2524);
or U3069 (N_3069,N_2852,N_2161);
nor U3070 (N_3070,N_2273,N_2484);
nor U3071 (N_3071,N_2540,N_2434);
or U3072 (N_3072,N_2040,N_2338);
or U3073 (N_3073,N_2071,N_2634);
nor U3074 (N_3074,N_2013,N_2776);
nand U3075 (N_3075,N_2739,N_2060);
or U3076 (N_3076,N_2997,N_2204);
nand U3077 (N_3077,N_2751,N_2749);
xnor U3078 (N_3078,N_2722,N_2011);
xnor U3079 (N_3079,N_2899,N_2353);
nand U3080 (N_3080,N_2326,N_2831);
or U3081 (N_3081,N_2873,N_2054);
xor U3082 (N_3082,N_2639,N_2557);
nand U3083 (N_3083,N_2805,N_2876);
nand U3084 (N_3084,N_2073,N_2939);
or U3085 (N_3085,N_2487,N_2740);
nor U3086 (N_3086,N_2268,N_2413);
nand U3087 (N_3087,N_2670,N_2964);
nor U3088 (N_3088,N_2660,N_2622);
xnor U3089 (N_3089,N_2454,N_2596);
and U3090 (N_3090,N_2667,N_2311);
nor U3091 (N_3091,N_2492,N_2599);
nand U3092 (N_3092,N_2033,N_2844);
or U3093 (N_3093,N_2216,N_2437);
nor U3094 (N_3094,N_2895,N_2147);
or U3095 (N_3095,N_2296,N_2635);
nor U3096 (N_3096,N_2941,N_2127);
or U3097 (N_3097,N_2822,N_2610);
xor U3098 (N_3098,N_2851,N_2834);
and U3099 (N_3099,N_2764,N_2905);
nor U3100 (N_3100,N_2214,N_2179);
xor U3101 (N_3101,N_2138,N_2203);
and U3102 (N_3102,N_2701,N_2167);
xor U3103 (N_3103,N_2756,N_2998);
nor U3104 (N_3104,N_2601,N_2213);
nand U3105 (N_3105,N_2205,N_2547);
and U3106 (N_3106,N_2485,N_2777);
or U3107 (N_3107,N_2200,N_2894);
nor U3108 (N_3108,N_2244,N_2004);
nor U3109 (N_3109,N_2666,N_2348);
and U3110 (N_3110,N_2452,N_2755);
and U3111 (N_3111,N_2808,N_2164);
and U3112 (N_3112,N_2075,N_2856);
xnor U3113 (N_3113,N_2473,N_2387);
xnor U3114 (N_3114,N_2565,N_2199);
xor U3115 (N_3115,N_2037,N_2265);
nand U3116 (N_3116,N_2264,N_2005);
nor U3117 (N_3117,N_2317,N_2744);
nand U3118 (N_3118,N_2202,N_2057);
nand U3119 (N_3119,N_2043,N_2661);
nor U3120 (N_3120,N_2501,N_2312);
nand U3121 (N_3121,N_2916,N_2909);
nor U3122 (N_3122,N_2280,N_2198);
or U3123 (N_3123,N_2572,N_2742);
and U3124 (N_3124,N_2640,N_2694);
nor U3125 (N_3125,N_2827,N_2787);
nand U3126 (N_3126,N_2675,N_2995);
nand U3127 (N_3127,N_2299,N_2745);
xor U3128 (N_3128,N_2417,N_2463);
or U3129 (N_3129,N_2382,N_2260);
or U3130 (N_3130,N_2173,N_2929);
nor U3131 (N_3131,N_2218,N_2464);
nor U3132 (N_3132,N_2594,N_2726);
nand U3133 (N_3133,N_2323,N_2719);
nand U3134 (N_3134,N_2598,N_2207);
nor U3135 (N_3135,N_2952,N_2864);
or U3136 (N_3136,N_2817,N_2149);
or U3137 (N_3137,N_2058,N_2959);
or U3138 (N_3138,N_2537,N_2589);
nand U3139 (N_3139,N_2583,N_2773);
or U3140 (N_3140,N_2151,N_2935);
and U3141 (N_3141,N_2221,N_2921);
nand U3142 (N_3142,N_2597,N_2684);
nor U3143 (N_3143,N_2630,N_2558);
nand U3144 (N_3144,N_2290,N_2321);
or U3145 (N_3145,N_2896,N_2195);
or U3146 (N_3146,N_2812,N_2181);
and U3147 (N_3147,N_2249,N_2209);
or U3148 (N_3148,N_2720,N_2030);
nand U3149 (N_3149,N_2307,N_2924);
nor U3150 (N_3150,N_2627,N_2088);
nor U3151 (N_3151,N_2632,N_2769);
and U3152 (N_3152,N_2910,N_2930);
and U3153 (N_3153,N_2373,N_2357);
and U3154 (N_3154,N_2697,N_2625);
and U3155 (N_3155,N_2380,N_2227);
and U3156 (N_3156,N_2902,N_2928);
nor U3157 (N_3157,N_2775,N_2222);
nand U3158 (N_3158,N_2143,N_2032);
xor U3159 (N_3159,N_2943,N_2578);
and U3160 (N_3160,N_2136,N_2566);
nor U3161 (N_3161,N_2132,N_2284);
nand U3162 (N_3162,N_2108,N_2302);
nand U3163 (N_3163,N_2472,N_2303);
xnor U3164 (N_3164,N_2223,N_2591);
or U3165 (N_3165,N_2468,N_2686);
nor U3166 (N_3166,N_2316,N_2238);
nand U3167 (N_3167,N_2887,N_2110);
and U3168 (N_3168,N_2092,N_2421);
nor U3169 (N_3169,N_2103,N_2888);
and U3170 (N_3170,N_2919,N_2066);
and U3171 (N_3171,N_2276,N_2352);
nor U3172 (N_3172,N_2183,N_2538);
nor U3173 (N_3173,N_2907,N_2849);
xnor U3174 (N_3174,N_2608,N_2460);
or U3175 (N_3175,N_2432,N_2241);
nand U3176 (N_3176,N_2516,N_2165);
and U3177 (N_3177,N_2620,N_2409);
xor U3178 (N_3178,N_2359,N_2840);
xor U3179 (N_3179,N_2763,N_2674);
or U3180 (N_3180,N_2070,N_2129);
xnor U3181 (N_3181,N_2823,N_2447);
xor U3182 (N_3182,N_2502,N_2613);
nand U3183 (N_3183,N_2954,N_2607);
xnor U3184 (N_3184,N_2306,N_2162);
xor U3185 (N_3185,N_2678,N_2875);
or U3186 (N_3186,N_2820,N_2969);
or U3187 (N_3187,N_2455,N_2837);
nand U3188 (N_3188,N_2267,N_2940);
nand U3189 (N_3189,N_2383,N_2142);
nor U3190 (N_3190,N_2677,N_2192);
xor U3191 (N_3191,N_2089,N_2692);
and U3192 (N_3192,N_2131,N_2987);
xnor U3193 (N_3193,N_2523,N_2711);
nand U3194 (N_3194,N_2890,N_2480);
nand U3195 (N_3195,N_2511,N_2091);
or U3196 (N_3196,N_2642,N_2458);
or U3197 (N_3197,N_2672,N_2766);
nor U3198 (N_3198,N_2977,N_2975);
and U3199 (N_3199,N_2390,N_2750);
and U3200 (N_3200,N_2982,N_2436);
and U3201 (N_3201,N_2514,N_2339);
xor U3202 (N_3202,N_2564,N_2291);
and U3203 (N_3203,N_2320,N_2190);
and U3204 (N_3204,N_2122,N_2522);
or U3205 (N_3205,N_2830,N_2211);
or U3206 (N_3206,N_2315,N_2470);
nor U3207 (N_3207,N_2865,N_2590);
nor U3208 (N_3208,N_2469,N_2710);
or U3209 (N_3209,N_2592,N_2543);
and U3210 (N_3210,N_2248,N_2879);
and U3211 (N_3211,N_2372,N_2245);
and U3212 (N_3212,N_2712,N_2786);
nor U3213 (N_3213,N_2424,N_2197);
xor U3214 (N_3214,N_2481,N_2504);
nor U3215 (N_3215,N_2360,N_2718);
xnor U3216 (N_3216,N_2099,N_2170);
or U3217 (N_3217,N_2846,N_2295);
nor U3218 (N_3218,N_2093,N_2908);
xnor U3219 (N_3219,N_2736,N_2498);
nand U3220 (N_3220,N_2815,N_2425);
or U3221 (N_3221,N_2239,N_2819);
nor U3222 (N_3222,N_2194,N_2735);
nor U3223 (N_3223,N_2656,N_2258);
xnor U3224 (N_3224,N_2048,N_2778);
or U3225 (N_3225,N_2546,N_2606);
nand U3226 (N_3226,N_2783,N_2933);
nor U3227 (N_3227,N_2991,N_2156);
nand U3228 (N_3228,N_2184,N_2577);
or U3229 (N_3229,N_2990,N_2560);
or U3230 (N_3230,N_2233,N_2476);
or U3231 (N_3231,N_2729,N_2673);
xnor U3232 (N_3232,N_2761,N_2477);
xor U3233 (N_3233,N_2658,N_2474);
or U3234 (N_3234,N_2376,N_2926);
xor U3235 (N_3235,N_2934,N_2003);
or U3236 (N_3236,N_2440,N_2272);
nor U3237 (N_3237,N_2451,N_2800);
nor U3238 (N_3238,N_2083,N_2422);
xor U3239 (N_3239,N_2158,N_2633);
and U3240 (N_3240,N_2467,N_2196);
nand U3241 (N_3241,N_2027,N_2361);
nor U3242 (N_3242,N_2381,N_2384);
nor U3243 (N_3243,N_2801,N_2892);
nor U3244 (N_3244,N_2554,N_2076);
nor U3245 (N_3245,N_2760,N_2240);
xor U3246 (N_3246,N_2839,N_2612);
nor U3247 (N_3247,N_2652,N_2884);
or U3248 (N_3248,N_2911,N_2486);
nand U3249 (N_3249,N_2278,N_2431);
or U3250 (N_3250,N_2141,N_2062);
nand U3251 (N_3251,N_2917,N_2681);
nor U3252 (N_3252,N_2292,N_2500);
xnor U3253 (N_3253,N_2378,N_2803);
and U3254 (N_3254,N_2269,N_2655);
xnor U3255 (N_3255,N_2746,N_2645);
nand U3256 (N_3256,N_2737,N_2938);
xnor U3257 (N_3257,N_2647,N_2858);
or U3258 (N_3258,N_2495,N_2017);
nand U3259 (N_3259,N_2410,N_2301);
xor U3260 (N_3260,N_2648,N_2086);
xnor U3261 (N_3261,N_2553,N_2309);
xor U3262 (N_3262,N_2024,N_2157);
nor U3263 (N_3263,N_2931,N_2163);
or U3264 (N_3264,N_2231,N_2541);
nor U3265 (N_3265,N_2397,N_2286);
or U3266 (N_3266,N_2914,N_2242);
nand U3267 (N_3267,N_2235,N_2246);
nor U3268 (N_3268,N_2738,N_2420);
or U3269 (N_3269,N_2113,N_2465);
and U3270 (N_3270,N_2515,N_2936);
and U3271 (N_3271,N_2080,N_2641);
or U3272 (N_3272,N_2979,N_2809);
nand U3273 (N_3273,N_2989,N_2488);
nor U3274 (N_3274,N_2009,N_2252);
xnor U3275 (N_3275,N_2428,N_2811);
nand U3276 (N_3276,N_2064,N_2377);
xor U3277 (N_3277,N_2682,N_2785);
and U3278 (N_3278,N_2918,N_2646);
and U3279 (N_3279,N_2716,N_2081);
or U3280 (N_3280,N_2243,N_2077);
xor U3281 (N_3281,N_2871,N_2889);
or U3282 (N_3282,N_2335,N_2462);
xor U3283 (N_3283,N_2687,N_2496);
nand U3284 (N_3284,N_2126,N_2580);
nand U3285 (N_3285,N_2283,N_2791);
and U3286 (N_3286,N_2691,N_2985);
xor U3287 (N_3287,N_2752,N_2419);
nand U3288 (N_3288,N_2406,N_2582);
nand U3289 (N_3289,N_2704,N_2958);
or U3290 (N_3290,N_2669,N_2724);
nor U3291 (N_3291,N_2664,N_2000);
xnor U3292 (N_3292,N_2259,N_2671);
nand U3293 (N_3293,N_2456,N_2574);
xor U3294 (N_3294,N_2789,N_2366);
or U3295 (N_3295,N_2703,N_2715);
nand U3296 (N_3296,N_2721,N_2407);
nand U3297 (N_3297,N_2945,N_2551);
or U3298 (N_3298,N_2951,N_2137);
or U3299 (N_3299,N_2604,N_2349);
nand U3300 (N_3300,N_2838,N_2539);
nor U3301 (N_3301,N_2617,N_2528);
and U3302 (N_3302,N_2059,N_2391);
xor U3303 (N_3303,N_2150,N_2327);
xnor U3304 (N_3304,N_2605,N_2257);
nand U3305 (N_3305,N_2446,N_2845);
and U3306 (N_3306,N_2867,N_2065);
or U3307 (N_3307,N_2313,N_2146);
nor U3308 (N_3308,N_2561,N_2573);
nor U3309 (N_3309,N_2340,N_2518);
nand U3310 (N_3310,N_2020,N_2507);
and U3311 (N_3311,N_2920,N_2039);
nor U3312 (N_3312,N_2595,N_2297);
or U3313 (N_3313,N_2688,N_2795);
xnor U3314 (N_3314,N_2714,N_2430);
nand U3315 (N_3315,N_2270,N_2139);
and U3316 (N_3316,N_2531,N_2025);
xor U3317 (N_3317,N_2426,N_2281);
or U3318 (N_3318,N_2796,N_2956);
xor U3319 (N_3319,N_2491,N_2813);
nor U3320 (N_3320,N_2169,N_2251);
or U3321 (N_3321,N_2322,N_2247);
nor U3322 (N_3322,N_2848,N_2946);
xor U3323 (N_3323,N_2781,N_2986);
or U3324 (N_3324,N_2289,N_2793);
and U3325 (N_3325,N_2836,N_2450);
nand U3326 (N_3326,N_2362,N_2713);
nor U3327 (N_3327,N_2224,N_2965);
nand U3328 (N_3328,N_2915,N_2877);
nand U3329 (N_3329,N_2332,N_2219);
and U3330 (N_3330,N_2569,N_2621);
and U3331 (N_3331,N_2293,N_2133);
nand U3332 (N_3332,N_2074,N_2193);
nand U3333 (N_3333,N_2482,N_2978);
nor U3334 (N_3334,N_2880,N_2626);
or U3335 (N_3335,N_2085,N_2282);
or U3336 (N_3336,N_2275,N_2782);
xor U3337 (N_3337,N_2234,N_2134);
and U3338 (N_3338,N_2847,N_2493);
or U3339 (N_3339,N_2759,N_2643);
nand U3340 (N_3340,N_2148,N_2449);
nor U3341 (N_3341,N_2525,N_2900);
and U3342 (N_3342,N_2471,N_2041);
nor U3343 (N_3343,N_2798,N_2364);
nand U3344 (N_3344,N_2651,N_2018);
and U3345 (N_3345,N_2114,N_2802);
nand U3346 (N_3346,N_2308,N_2657);
or U3347 (N_3347,N_2534,N_2427);
nor U3348 (N_3348,N_2850,N_2189);
nor U3349 (N_3349,N_2753,N_2160);
or U3350 (N_3350,N_2228,N_2459);
or U3351 (N_3351,N_2949,N_2333);
and U3352 (N_3352,N_2695,N_2416);
nor U3353 (N_3353,N_2881,N_2707);
nand U3354 (N_3354,N_2226,N_2957);
or U3355 (N_3355,N_2559,N_2874);
nand U3356 (N_3356,N_2770,N_2288);
xnor U3357 (N_3357,N_2863,N_2365);
and U3358 (N_3358,N_2393,N_2927);
or U3359 (N_3359,N_2342,N_2790);
and U3360 (N_3360,N_2549,N_2799);
nand U3361 (N_3361,N_2185,N_2318);
and U3362 (N_3362,N_2367,N_2842);
or U3363 (N_3363,N_2503,N_2078);
nand U3364 (N_3364,N_2857,N_2489);
nor U3365 (N_3365,N_2176,N_2741);
or U3366 (N_3366,N_2649,N_2556);
nand U3367 (N_3367,N_2829,N_2399);
and U3368 (N_3368,N_2974,N_2250);
nor U3369 (N_3369,N_2774,N_2014);
nand U3370 (N_3370,N_2415,N_2038);
or U3371 (N_3371,N_2191,N_2555);
or U3372 (N_3372,N_2659,N_2212);
and U3373 (N_3373,N_2001,N_2109);
nand U3374 (N_3374,N_2029,N_2237);
xnor U3375 (N_3375,N_2855,N_2144);
nor U3376 (N_3376,N_2520,N_2925);
and U3377 (N_3377,N_2768,N_2727);
nand U3378 (N_3378,N_2279,N_2112);
xor U3379 (N_3379,N_2797,N_2408);
and U3380 (N_3380,N_2121,N_2355);
xnor U3381 (N_3381,N_2111,N_2728);
nand U3382 (N_3382,N_2159,N_2441);
and U3383 (N_3383,N_2433,N_2602);
nor U3384 (N_3384,N_2097,N_2166);
nor U3385 (N_3385,N_2861,N_2765);
xnor U3386 (N_3386,N_2732,N_2096);
and U3387 (N_3387,N_2913,N_2046);
xnor U3388 (N_3388,N_2351,N_2689);
or U3389 (N_3389,N_2175,N_2825);
xor U3390 (N_3390,N_2002,N_2535);
or U3391 (N_3391,N_2287,N_2944);
xor U3392 (N_3392,N_2120,N_2358);
and U3393 (N_3393,N_2581,N_2329);
and U3394 (N_3394,N_2542,N_2567);
nor U3395 (N_3395,N_2395,N_2882);
or U3396 (N_3396,N_2637,N_2336);
nand U3397 (N_3397,N_2379,N_2866);
xor U3398 (N_3398,N_2128,N_2699);
xor U3399 (N_3399,N_2912,N_2980);
or U3400 (N_3400,N_2821,N_2841);
and U3401 (N_3401,N_2172,N_2396);
and U3402 (N_3402,N_2973,N_2984);
nand U3403 (N_3403,N_2548,N_2807);
nor U3404 (N_3404,N_2063,N_2950);
or U3405 (N_3405,N_2210,N_2631);
nor U3406 (N_3406,N_2300,N_2709);
and U3407 (N_3407,N_2152,N_2593);
or U3408 (N_3408,N_2571,N_2510);
nor U3409 (N_3409,N_2069,N_2513);
nand U3410 (N_3410,N_2922,N_2031);
nor U3411 (N_3411,N_2266,N_2754);
nand U3412 (N_3412,N_2771,N_2816);
or U3413 (N_3413,N_2843,N_2584);
nor U3414 (N_3414,N_2967,N_2529);
or U3415 (N_3415,N_2788,N_2098);
and U3416 (N_3416,N_2706,N_2007);
nor U3417 (N_3417,N_2748,N_2056);
or U3418 (N_3418,N_2429,N_2217);
and U3419 (N_3419,N_2705,N_2403);
nand U3420 (N_3420,N_2901,N_2972);
xor U3421 (N_3421,N_2047,N_2490);
nand U3422 (N_3422,N_2629,N_2942);
or U3423 (N_3423,N_2314,N_2044);
nor U3424 (N_3424,N_2832,N_2833);
xor U3425 (N_3425,N_2298,N_2423);
and U3426 (N_3426,N_2049,N_2932);
xor U3427 (N_3427,N_2053,N_2550);
or U3428 (N_3428,N_2116,N_2389);
nand U3429 (N_3429,N_2345,N_2702);
nor U3430 (N_3430,N_2106,N_2263);
and U3431 (N_3431,N_2650,N_2552);
or U3432 (N_3432,N_2155,N_2575);
and U3433 (N_3433,N_2145,N_2579);
nand U3434 (N_3434,N_2784,N_2404);
or U3435 (N_3435,N_2587,N_2665);
and U3436 (N_3436,N_2794,N_2885);
nand U3437 (N_3437,N_2225,N_2100);
nand U3438 (N_3438,N_2034,N_2061);
nor U3439 (N_3439,N_2479,N_2527);
nor U3440 (N_3440,N_2509,N_2050);
nor U3441 (N_3441,N_2700,N_2767);
or U3442 (N_3442,N_2685,N_2757);
nor U3443 (N_3443,N_2363,N_2079);
xnor U3444 (N_3444,N_2230,N_2733);
and U3445 (N_3445,N_2505,N_2117);
nor U3446 (N_3446,N_2698,N_2341);
xnor U3447 (N_3447,N_2609,N_2124);
and U3448 (N_3448,N_2966,N_2022);
and U3449 (N_3449,N_2772,N_2052);
or U3450 (N_3450,N_2140,N_2095);
nor U3451 (N_3451,N_2010,N_2953);
nor U3452 (N_3452,N_2779,N_2804);
nor U3453 (N_3453,N_2036,N_2016);
nor U3454 (N_3454,N_2344,N_2859);
or U3455 (N_3455,N_2870,N_2810);
nor U3456 (N_3456,N_2346,N_2854);
xor U3457 (N_3457,N_2758,N_2325);
and U3458 (N_3458,N_2084,N_2305);
or U3459 (N_3459,N_2354,N_2019);
xnor U3460 (N_3460,N_2418,N_2992);
xor U3461 (N_3461,N_2400,N_2903);
and U3462 (N_3462,N_2208,N_2371);
and U3463 (N_3463,N_2497,N_2042);
and U3464 (N_3464,N_2008,N_2119);
nor U3465 (N_3465,N_2668,N_2532);
nor U3466 (N_3466,N_2188,N_2453);
and U3467 (N_3467,N_2330,N_2328);
and U3468 (N_3468,N_2962,N_2294);
nand U3469 (N_3469,N_2094,N_2392);
nor U3470 (N_3470,N_2994,N_2730);
or U3471 (N_3471,N_2123,N_2869);
or U3472 (N_3472,N_2860,N_2923);
nand U3473 (N_3473,N_2028,N_2576);
xnor U3474 (N_3474,N_2747,N_2105);
nor U3475 (N_3475,N_2483,N_2512);
nor U3476 (N_3476,N_2186,N_2256);
nor U3477 (N_3477,N_2153,N_2457);
xor U3478 (N_3478,N_2536,N_2402);
nand U3479 (N_3479,N_2324,N_2999);
xnor U3480 (N_3480,N_2051,N_2615);
or U3481 (N_3481,N_2229,N_2072);
or U3482 (N_3482,N_2444,N_2171);
or U3483 (N_3483,N_2947,N_2898);
nor U3484 (N_3484,N_2262,N_2466);
nor U3485 (N_3485,N_2762,N_2494);
or U3486 (N_3486,N_2412,N_2021);
and U3487 (N_3487,N_2180,N_2616);
or U3488 (N_3488,N_2961,N_2499);
nor U3489 (N_3489,N_2960,N_2976);
xor U3490 (N_3490,N_2996,N_2611);
and U3491 (N_3491,N_2253,N_2369);
or U3492 (N_3492,N_2526,N_2725);
or U3493 (N_3493,N_2948,N_2442);
xor U3494 (N_3494,N_2614,N_2285);
nand U3495 (N_3495,N_2824,N_2182);
and U3496 (N_3496,N_2878,N_2506);
and U3497 (N_3497,N_2862,N_2331);
or U3498 (N_3498,N_2508,N_2401);
or U3499 (N_3499,N_2232,N_2461);
and U3500 (N_3500,N_2592,N_2030);
nand U3501 (N_3501,N_2125,N_2925);
nand U3502 (N_3502,N_2834,N_2586);
xor U3503 (N_3503,N_2746,N_2177);
xor U3504 (N_3504,N_2272,N_2354);
xor U3505 (N_3505,N_2309,N_2295);
xor U3506 (N_3506,N_2257,N_2715);
xor U3507 (N_3507,N_2438,N_2783);
and U3508 (N_3508,N_2387,N_2194);
xnor U3509 (N_3509,N_2099,N_2726);
nor U3510 (N_3510,N_2183,N_2142);
xnor U3511 (N_3511,N_2629,N_2994);
nand U3512 (N_3512,N_2576,N_2946);
xor U3513 (N_3513,N_2712,N_2744);
nor U3514 (N_3514,N_2365,N_2477);
nor U3515 (N_3515,N_2681,N_2729);
and U3516 (N_3516,N_2365,N_2669);
xor U3517 (N_3517,N_2112,N_2091);
xor U3518 (N_3518,N_2592,N_2399);
nand U3519 (N_3519,N_2702,N_2163);
xnor U3520 (N_3520,N_2152,N_2312);
nor U3521 (N_3521,N_2403,N_2593);
or U3522 (N_3522,N_2198,N_2973);
xnor U3523 (N_3523,N_2929,N_2190);
xnor U3524 (N_3524,N_2507,N_2161);
nand U3525 (N_3525,N_2981,N_2760);
xnor U3526 (N_3526,N_2245,N_2688);
nand U3527 (N_3527,N_2338,N_2947);
xnor U3528 (N_3528,N_2017,N_2795);
nand U3529 (N_3529,N_2146,N_2151);
nand U3530 (N_3530,N_2310,N_2452);
nor U3531 (N_3531,N_2575,N_2164);
xor U3532 (N_3532,N_2698,N_2441);
nand U3533 (N_3533,N_2618,N_2132);
nand U3534 (N_3534,N_2685,N_2424);
nand U3535 (N_3535,N_2949,N_2676);
nand U3536 (N_3536,N_2212,N_2251);
or U3537 (N_3537,N_2371,N_2166);
nand U3538 (N_3538,N_2678,N_2608);
xnor U3539 (N_3539,N_2441,N_2648);
nand U3540 (N_3540,N_2247,N_2139);
or U3541 (N_3541,N_2172,N_2497);
nand U3542 (N_3542,N_2632,N_2648);
nand U3543 (N_3543,N_2537,N_2949);
or U3544 (N_3544,N_2569,N_2349);
nand U3545 (N_3545,N_2740,N_2405);
and U3546 (N_3546,N_2183,N_2064);
and U3547 (N_3547,N_2328,N_2912);
and U3548 (N_3548,N_2290,N_2606);
xnor U3549 (N_3549,N_2696,N_2405);
xor U3550 (N_3550,N_2070,N_2999);
nor U3551 (N_3551,N_2774,N_2274);
nand U3552 (N_3552,N_2199,N_2730);
nand U3553 (N_3553,N_2827,N_2889);
xor U3554 (N_3554,N_2968,N_2867);
xor U3555 (N_3555,N_2425,N_2350);
or U3556 (N_3556,N_2947,N_2047);
nand U3557 (N_3557,N_2697,N_2867);
or U3558 (N_3558,N_2659,N_2225);
xor U3559 (N_3559,N_2536,N_2803);
nand U3560 (N_3560,N_2619,N_2509);
nand U3561 (N_3561,N_2336,N_2650);
or U3562 (N_3562,N_2066,N_2446);
xor U3563 (N_3563,N_2455,N_2443);
or U3564 (N_3564,N_2947,N_2896);
or U3565 (N_3565,N_2500,N_2502);
or U3566 (N_3566,N_2709,N_2435);
and U3567 (N_3567,N_2257,N_2533);
nor U3568 (N_3568,N_2871,N_2747);
xor U3569 (N_3569,N_2391,N_2450);
xor U3570 (N_3570,N_2015,N_2728);
nand U3571 (N_3571,N_2283,N_2018);
nor U3572 (N_3572,N_2098,N_2087);
nand U3573 (N_3573,N_2973,N_2582);
nand U3574 (N_3574,N_2987,N_2655);
and U3575 (N_3575,N_2108,N_2921);
xnor U3576 (N_3576,N_2476,N_2722);
and U3577 (N_3577,N_2201,N_2631);
and U3578 (N_3578,N_2842,N_2575);
xor U3579 (N_3579,N_2766,N_2178);
xnor U3580 (N_3580,N_2637,N_2096);
and U3581 (N_3581,N_2812,N_2057);
and U3582 (N_3582,N_2280,N_2701);
nand U3583 (N_3583,N_2462,N_2338);
or U3584 (N_3584,N_2497,N_2438);
and U3585 (N_3585,N_2201,N_2610);
and U3586 (N_3586,N_2569,N_2233);
nor U3587 (N_3587,N_2217,N_2381);
xnor U3588 (N_3588,N_2365,N_2857);
nor U3589 (N_3589,N_2779,N_2144);
xor U3590 (N_3590,N_2833,N_2479);
nor U3591 (N_3591,N_2750,N_2970);
nor U3592 (N_3592,N_2575,N_2914);
xnor U3593 (N_3593,N_2410,N_2390);
or U3594 (N_3594,N_2215,N_2221);
or U3595 (N_3595,N_2049,N_2666);
xor U3596 (N_3596,N_2693,N_2511);
nor U3597 (N_3597,N_2280,N_2929);
nand U3598 (N_3598,N_2887,N_2857);
and U3599 (N_3599,N_2157,N_2499);
or U3600 (N_3600,N_2912,N_2302);
and U3601 (N_3601,N_2307,N_2218);
xor U3602 (N_3602,N_2075,N_2895);
nor U3603 (N_3603,N_2114,N_2209);
nor U3604 (N_3604,N_2349,N_2828);
nor U3605 (N_3605,N_2969,N_2594);
and U3606 (N_3606,N_2615,N_2589);
xnor U3607 (N_3607,N_2935,N_2522);
xor U3608 (N_3608,N_2463,N_2026);
nand U3609 (N_3609,N_2597,N_2781);
and U3610 (N_3610,N_2814,N_2827);
nand U3611 (N_3611,N_2751,N_2944);
nand U3612 (N_3612,N_2238,N_2331);
nor U3613 (N_3613,N_2317,N_2162);
and U3614 (N_3614,N_2998,N_2439);
xnor U3615 (N_3615,N_2911,N_2035);
or U3616 (N_3616,N_2147,N_2891);
or U3617 (N_3617,N_2408,N_2067);
xor U3618 (N_3618,N_2118,N_2435);
and U3619 (N_3619,N_2346,N_2220);
and U3620 (N_3620,N_2171,N_2951);
nor U3621 (N_3621,N_2912,N_2139);
nand U3622 (N_3622,N_2132,N_2655);
xor U3623 (N_3623,N_2220,N_2163);
xnor U3624 (N_3624,N_2893,N_2251);
nand U3625 (N_3625,N_2822,N_2196);
or U3626 (N_3626,N_2380,N_2291);
xor U3627 (N_3627,N_2916,N_2769);
nand U3628 (N_3628,N_2570,N_2433);
or U3629 (N_3629,N_2217,N_2116);
or U3630 (N_3630,N_2941,N_2659);
nor U3631 (N_3631,N_2827,N_2763);
xnor U3632 (N_3632,N_2483,N_2566);
xnor U3633 (N_3633,N_2695,N_2315);
and U3634 (N_3634,N_2287,N_2455);
nand U3635 (N_3635,N_2074,N_2616);
nand U3636 (N_3636,N_2276,N_2380);
nor U3637 (N_3637,N_2257,N_2183);
xnor U3638 (N_3638,N_2300,N_2617);
nand U3639 (N_3639,N_2042,N_2826);
nor U3640 (N_3640,N_2055,N_2514);
and U3641 (N_3641,N_2419,N_2937);
nand U3642 (N_3642,N_2048,N_2483);
and U3643 (N_3643,N_2053,N_2797);
xor U3644 (N_3644,N_2121,N_2311);
nand U3645 (N_3645,N_2677,N_2472);
nor U3646 (N_3646,N_2114,N_2584);
nor U3647 (N_3647,N_2186,N_2253);
nand U3648 (N_3648,N_2954,N_2003);
nor U3649 (N_3649,N_2222,N_2022);
nand U3650 (N_3650,N_2126,N_2543);
or U3651 (N_3651,N_2188,N_2927);
nand U3652 (N_3652,N_2576,N_2208);
nand U3653 (N_3653,N_2928,N_2625);
or U3654 (N_3654,N_2782,N_2574);
nand U3655 (N_3655,N_2910,N_2631);
or U3656 (N_3656,N_2542,N_2660);
nand U3657 (N_3657,N_2924,N_2370);
nor U3658 (N_3658,N_2201,N_2708);
xor U3659 (N_3659,N_2876,N_2075);
or U3660 (N_3660,N_2156,N_2568);
nor U3661 (N_3661,N_2349,N_2418);
nor U3662 (N_3662,N_2005,N_2948);
nor U3663 (N_3663,N_2113,N_2391);
and U3664 (N_3664,N_2383,N_2298);
xor U3665 (N_3665,N_2215,N_2809);
nand U3666 (N_3666,N_2163,N_2915);
or U3667 (N_3667,N_2793,N_2517);
nor U3668 (N_3668,N_2514,N_2326);
or U3669 (N_3669,N_2164,N_2933);
xnor U3670 (N_3670,N_2310,N_2078);
nor U3671 (N_3671,N_2271,N_2735);
xnor U3672 (N_3672,N_2253,N_2155);
xor U3673 (N_3673,N_2607,N_2538);
or U3674 (N_3674,N_2751,N_2542);
or U3675 (N_3675,N_2624,N_2785);
or U3676 (N_3676,N_2838,N_2505);
and U3677 (N_3677,N_2420,N_2508);
nor U3678 (N_3678,N_2238,N_2764);
xor U3679 (N_3679,N_2111,N_2540);
xnor U3680 (N_3680,N_2299,N_2384);
nand U3681 (N_3681,N_2789,N_2298);
nor U3682 (N_3682,N_2117,N_2353);
or U3683 (N_3683,N_2603,N_2365);
nand U3684 (N_3684,N_2493,N_2205);
and U3685 (N_3685,N_2325,N_2114);
and U3686 (N_3686,N_2165,N_2910);
xnor U3687 (N_3687,N_2907,N_2107);
nand U3688 (N_3688,N_2634,N_2341);
xnor U3689 (N_3689,N_2838,N_2418);
or U3690 (N_3690,N_2147,N_2690);
nand U3691 (N_3691,N_2161,N_2387);
nor U3692 (N_3692,N_2588,N_2401);
xor U3693 (N_3693,N_2743,N_2719);
nor U3694 (N_3694,N_2702,N_2916);
or U3695 (N_3695,N_2211,N_2788);
or U3696 (N_3696,N_2221,N_2513);
nand U3697 (N_3697,N_2435,N_2119);
nor U3698 (N_3698,N_2582,N_2054);
and U3699 (N_3699,N_2589,N_2103);
nor U3700 (N_3700,N_2971,N_2549);
nand U3701 (N_3701,N_2288,N_2133);
and U3702 (N_3702,N_2465,N_2905);
or U3703 (N_3703,N_2654,N_2635);
and U3704 (N_3704,N_2811,N_2712);
and U3705 (N_3705,N_2974,N_2799);
xor U3706 (N_3706,N_2596,N_2573);
xor U3707 (N_3707,N_2428,N_2326);
xor U3708 (N_3708,N_2202,N_2190);
nand U3709 (N_3709,N_2792,N_2205);
xnor U3710 (N_3710,N_2602,N_2978);
nand U3711 (N_3711,N_2705,N_2542);
or U3712 (N_3712,N_2172,N_2048);
xnor U3713 (N_3713,N_2918,N_2814);
nand U3714 (N_3714,N_2774,N_2237);
and U3715 (N_3715,N_2297,N_2287);
xnor U3716 (N_3716,N_2166,N_2663);
xor U3717 (N_3717,N_2501,N_2451);
xor U3718 (N_3718,N_2788,N_2786);
nor U3719 (N_3719,N_2078,N_2956);
and U3720 (N_3720,N_2365,N_2271);
and U3721 (N_3721,N_2169,N_2913);
xor U3722 (N_3722,N_2635,N_2245);
nor U3723 (N_3723,N_2885,N_2647);
and U3724 (N_3724,N_2313,N_2559);
nand U3725 (N_3725,N_2497,N_2825);
nor U3726 (N_3726,N_2855,N_2171);
nand U3727 (N_3727,N_2724,N_2051);
nand U3728 (N_3728,N_2372,N_2948);
nor U3729 (N_3729,N_2934,N_2677);
xnor U3730 (N_3730,N_2549,N_2995);
and U3731 (N_3731,N_2063,N_2241);
nand U3732 (N_3732,N_2186,N_2323);
nand U3733 (N_3733,N_2682,N_2658);
or U3734 (N_3734,N_2631,N_2113);
xor U3735 (N_3735,N_2586,N_2856);
or U3736 (N_3736,N_2732,N_2632);
xnor U3737 (N_3737,N_2393,N_2899);
and U3738 (N_3738,N_2236,N_2346);
nor U3739 (N_3739,N_2454,N_2030);
xor U3740 (N_3740,N_2705,N_2591);
xor U3741 (N_3741,N_2884,N_2501);
nor U3742 (N_3742,N_2983,N_2284);
xnor U3743 (N_3743,N_2487,N_2953);
and U3744 (N_3744,N_2726,N_2695);
nor U3745 (N_3745,N_2471,N_2465);
xnor U3746 (N_3746,N_2031,N_2082);
nand U3747 (N_3747,N_2968,N_2860);
xor U3748 (N_3748,N_2768,N_2878);
or U3749 (N_3749,N_2909,N_2876);
and U3750 (N_3750,N_2098,N_2371);
xnor U3751 (N_3751,N_2968,N_2171);
nor U3752 (N_3752,N_2110,N_2328);
nor U3753 (N_3753,N_2230,N_2525);
or U3754 (N_3754,N_2431,N_2401);
or U3755 (N_3755,N_2383,N_2777);
or U3756 (N_3756,N_2743,N_2946);
nor U3757 (N_3757,N_2998,N_2959);
or U3758 (N_3758,N_2354,N_2042);
xnor U3759 (N_3759,N_2835,N_2778);
nor U3760 (N_3760,N_2639,N_2905);
nor U3761 (N_3761,N_2127,N_2664);
nand U3762 (N_3762,N_2753,N_2136);
nor U3763 (N_3763,N_2260,N_2563);
xor U3764 (N_3764,N_2304,N_2086);
nor U3765 (N_3765,N_2092,N_2780);
or U3766 (N_3766,N_2019,N_2494);
xor U3767 (N_3767,N_2189,N_2537);
nor U3768 (N_3768,N_2698,N_2123);
nand U3769 (N_3769,N_2016,N_2722);
nor U3770 (N_3770,N_2237,N_2299);
nor U3771 (N_3771,N_2577,N_2121);
nor U3772 (N_3772,N_2035,N_2709);
or U3773 (N_3773,N_2446,N_2492);
and U3774 (N_3774,N_2338,N_2053);
and U3775 (N_3775,N_2628,N_2886);
or U3776 (N_3776,N_2199,N_2003);
or U3777 (N_3777,N_2324,N_2861);
nor U3778 (N_3778,N_2425,N_2318);
or U3779 (N_3779,N_2608,N_2670);
xor U3780 (N_3780,N_2924,N_2115);
and U3781 (N_3781,N_2211,N_2816);
and U3782 (N_3782,N_2252,N_2717);
nor U3783 (N_3783,N_2959,N_2084);
and U3784 (N_3784,N_2052,N_2348);
and U3785 (N_3785,N_2718,N_2093);
nor U3786 (N_3786,N_2059,N_2418);
and U3787 (N_3787,N_2336,N_2831);
nand U3788 (N_3788,N_2588,N_2746);
and U3789 (N_3789,N_2662,N_2647);
or U3790 (N_3790,N_2459,N_2541);
nand U3791 (N_3791,N_2670,N_2389);
or U3792 (N_3792,N_2963,N_2389);
nor U3793 (N_3793,N_2433,N_2755);
nand U3794 (N_3794,N_2220,N_2423);
nor U3795 (N_3795,N_2744,N_2819);
nand U3796 (N_3796,N_2652,N_2075);
or U3797 (N_3797,N_2955,N_2083);
nor U3798 (N_3798,N_2709,N_2684);
nand U3799 (N_3799,N_2959,N_2601);
and U3800 (N_3800,N_2559,N_2574);
nand U3801 (N_3801,N_2048,N_2405);
and U3802 (N_3802,N_2699,N_2162);
nand U3803 (N_3803,N_2706,N_2430);
nand U3804 (N_3804,N_2653,N_2444);
and U3805 (N_3805,N_2294,N_2526);
nand U3806 (N_3806,N_2567,N_2922);
xor U3807 (N_3807,N_2633,N_2055);
xnor U3808 (N_3808,N_2363,N_2403);
and U3809 (N_3809,N_2044,N_2400);
xnor U3810 (N_3810,N_2368,N_2033);
nor U3811 (N_3811,N_2270,N_2617);
xor U3812 (N_3812,N_2326,N_2426);
or U3813 (N_3813,N_2772,N_2465);
nand U3814 (N_3814,N_2855,N_2708);
and U3815 (N_3815,N_2458,N_2199);
or U3816 (N_3816,N_2793,N_2992);
and U3817 (N_3817,N_2938,N_2827);
xnor U3818 (N_3818,N_2773,N_2842);
and U3819 (N_3819,N_2488,N_2505);
or U3820 (N_3820,N_2595,N_2500);
xnor U3821 (N_3821,N_2560,N_2941);
xor U3822 (N_3822,N_2959,N_2562);
and U3823 (N_3823,N_2023,N_2269);
and U3824 (N_3824,N_2475,N_2721);
nand U3825 (N_3825,N_2199,N_2152);
xnor U3826 (N_3826,N_2564,N_2571);
xnor U3827 (N_3827,N_2303,N_2922);
or U3828 (N_3828,N_2242,N_2637);
xnor U3829 (N_3829,N_2099,N_2596);
nor U3830 (N_3830,N_2934,N_2969);
and U3831 (N_3831,N_2954,N_2600);
xnor U3832 (N_3832,N_2889,N_2906);
or U3833 (N_3833,N_2578,N_2422);
nor U3834 (N_3834,N_2743,N_2643);
nand U3835 (N_3835,N_2391,N_2253);
xnor U3836 (N_3836,N_2366,N_2457);
nand U3837 (N_3837,N_2541,N_2321);
xnor U3838 (N_3838,N_2403,N_2199);
xor U3839 (N_3839,N_2919,N_2946);
xor U3840 (N_3840,N_2601,N_2281);
and U3841 (N_3841,N_2982,N_2087);
and U3842 (N_3842,N_2981,N_2664);
nor U3843 (N_3843,N_2369,N_2335);
nand U3844 (N_3844,N_2595,N_2184);
nor U3845 (N_3845,N_2440,N_2282);
or U3846 (N_3846,N_2448,N_2080);
nand U3847 (N_3847,N_2503,N_2001);
nand U3848 (N_3848,N_2721,N_2739);
or U3849 (N_3849,N_2915,N_2263);
or U3850 (N_3850,N_2188,N_2334);
nor U3851 (N_3851,N_2015,N_2353);
or U3852 (N_3852,N_2748,N_2348);
nor U3853 (N_3853,N_2980,N_2482);
nand U3854 (N_3854,N_2111,N_2210);
nand U3855 (N_3855,N_2007,N_2293);
nor U3856 (N_3856,N_2471,N_2125);
nor U3857 (N_3857,N_2206,N_2290);
nor U3858 (N_3858,N_2236,N_2748);
nor U3859 (N_3859,N_2460,N_2331);
nand U3860 (N_3860,N_2472,N_2154);
or U3861 (N_3861,N_2245,N_2735);
or U3862 (N_3862,N_2923,N_2422);
and U3863 (N_3863,N_2921,N_2099);
and U3864 (N_3864,N_2685,N_2596);
or U3865 (N_3865,N_2807,N_2949);
nor U3866 (N_3866,N_2431,N_2749);
and U3867 (N_3867,N_2464,N_2340);
xor U3868 (N_3868,N_2589,N_2345);
or U3869 (N_3869,N_2051,N_2462);
or U3870 (N_3870,N_2160,N_2705);
or U3871 (N_3871,N_2218,N_2148);
and U3872 (N_3872,N_2977,N_2654);
xnor U3873 (N_3873,N_2325,N_2120);
and U3874 (N_3874,N_2405,N_2552);
or U3875 (N_3875,N_2368,N_2653);
nand U3876 (N_3876,N_2163,N_2458);
and U3877 (N_3877,N_2198,N_2132);
nand U3878 (N_3878,N_2416,N_2247);
and U3879 (N_3879,N_2184,N_2640);
xor U3880 (N_3880,N_2992,N_2907);
xor U3881 (N_3881,N_2188,N_2473);
and U3882 (N_3882,N_2794,N_2820);
or U3883 (N_3883,N_2632,N_2913);
nand U3884 (N_3884,N_2402,N_2923);
and U3885 (N_3885,N_2598,N_2046);
nor U3886 (N_3886,N_2340,N_2961);
or U3887 (N_3887,N_2350,N_2819);
nand U3888 (N_3888,N_2364,N_2465);
and U3889 (N_3889,N_2233,N_2161);
nand U3890 (N_3890,N_2600,N_2836);
and U3891 (N_3891,N_2169,N_2909);
nand U3892 (N_3892,N_2384,N_2391);
nor U3893 (N_3893,N_2943,N_2238);
nor U3894 (N_3894,N_2341,N_2914);
nor U3895 (N_3895,N_2400,N_2876);
and U3896 (N_3896,N_2817,N_2229);
or U3897 (N_3897,N_2647,N_2538);
nand U3898 (N_3898,N_2501,N_2350);
or U3899 (N_3899,N_2581,N_2739);
and U3900 (N_3900,N_2454,N_2127);
and U3901 (N_3901,N_2317,N_2544);
xor U3902 (N_3902,N_2192,N_2619);
and U3903 (N_3903,N_2493,N_2480);
nor U3904 (N_3904,N_2465,N_2895);
xnor U3905 (N_3905,N_2009,N_2092);
nand U3906 (N_3906,N_2260,N_2258);
nor U3907 (N_3907,N_2757,N_2962);
xnor U3908 (N_3908,N_2161,N_2216);
nand U3909 (N_3909,N_2870,N_2180);
nand U3910 (N_3910,N_2587,N_2871);
nand U3911 (N_3911,N_2214,N_2516);
xor U3912 (N_3912,N_2385,N_2543);
and U3913 (N_3913,N_2724,N_2472);
nand U3914 (N_3914,N_2126,N_2651);
nor U3915 (N_3915,N_2475,N_2159);
nor U3916 (N_3916,N_2896,N_2246);
nor U3917 (N_3917,N_2419,N_2028);
nor U3918 (N_3918,N_2540,N_2985);
nand U3919 (N_3919,N_2660,N_2483);
nor U3920 (N_3920,N_2318,N_2910);
nand U3921 (N_3921,N_2005,N_2977);
and U3922 (N_3922,N_2098,N_2525);
nand U3923 (N_3923,N_2747,N_2062);
or U3924 (N_3924,N_2425,N_2242);
and U3925 (N_3925,N_2554,N_2130);
nand U3926 (N_3926,N_2460,N_2929);
nor U3927 (N_3927,N_2163,N_2662);
nor U3928 (N_3928,N_2280,N_2727);
or U3929 (N_3929,N_2954,N_2522);
nor U3930 (N_3930,N_2329,N_2859);
or U3931 (N_3931,N_2370,N_2425);
or U3932 (N_3932,N_2515,N_2256);
or U3933 (N_3933,N_2432,N_2820);
or U3934 (N_3934,N_2440,N_2258);
nand U3935 (N_3935,N_2255,N_2530);
nand U3936 (N_3936,N_2762,N_2818);
nor U3937 (N_3937,N_2094,N_2817);
or U3938 (N_3938,N_2295,N_2816);
nor U3939 (N_3939,N_2778,N_2542);
and U3940 (N_3940,N_2225,N_2366);
nand U3941 (N_3941,N_2165,N_2365);
xnor U3942 (N_3942,N_2042,N_2416);
nand U3943 (N_3943,N_2572,N_2741);
xor U3944 (N_3944,N_2359,N_2052);
xnor U3945 (N_3945,N_2698,N_2334);
nand U3946 (N_3946,N_2785,N_2894);
nand U3947 (N_3947,N_2740,N_2755);
nor U3948 (N_3948,N_2851,N_2397);
nor U3949 (N_3949,N_2981,N_2245);
xor U3950 (N_3950,N_2289,N_2612);
or U3951 (N_3951,N_2268,N_2489);
or U3952 (N_3952,N_2028,N_2039);
xnor U3953 (N_3953,N_2159,N_2649);
nand U3954 (N_3954,N_2820,N_2967);
or U3955 (N_3955,N_2345,N_2823);
nor U3956 (N_3956,N_2510,N_2047);
nor U3957 (N_3957,N_2866,N_2962);
and U3958 (N_3958,N_2421,N_2102);
xor U3959 (N_3959,N_2840,N_2124);
xor U3960 (N_3960,N_2564,N_2981);
nor U3961 (N_3961,N_2876,N_2762);
or U3962 (N_3962,N_2035,N_2719);
xor U3963 (N_3963,N_2210,N_2164);
xnor U3964 (N_3964,N_2582,N_2114);
nand U3965 (N_3965,N_2093,N_2551);
or U3966 (N_3966,N_2369,N_2536);
xor U3967 (N_3967,N_2481,N_2517);
xor U3968 (N_3968,N_2329,N_2723);
xor U3969 (N_3969,N_2621,N_2256);
and U3970 (N_3970,N_2485,N_2717);
or U3971 (N_3971,N_2589,N_2484);
or U3972 (N_3972,N_2243,N_2930);
and U3973 (N_3973,N_2970,N_2647);
nand U3974 (N_3974,N_2247,N_2508);
nand U3975 (N_3975,N_2039,N_2638);
xnor U3976 (N_3976,N_2552,N_2509);
xor U3977 (N_3977,N_2519,N_2480);
or U3978 (N_3978,N_2935,N_2842);
and U3979 (N_3979,N_2296,N_2373);
or U3980 (N_3980,N_2901,N_2928);
and U3981 (N_3981,N_2408,N_2822);
nor U3982 (N_3982,N_2980,N_2926);
and U3983 (N_3983,N_2178,N_2630);
nor U3984 (N_3984,N_2674,N_2573);
and U3985 (N_3985,N_2010,N_2338);
nor U3986 (N_3986,N_2413,N_2821);
nand U3987 (N_3987,N_2798,N_2226);
nor U3988 (N_3988,N_2518,N_2400);
nor U3989 (N_3989,N_2558,N_2196);
or U3990 (N_3990,N_2505,N_2136);
xnor U3991 (N_3991,N_2884,N_2106);
or U3992 (N_3992,N_2707,N_2318);
and U3993 (N_3993,N_2365,N_2823);
and U3994 (N_3994,N_2274,N_2535);
and U3995 (N_3995,N_2283,N_2401);
and U3996 (N_3996,N_2208,N_2584);
and U3997 (N_3997,N_2335,N_2734);
xor U3998 (N_3998,N_2596,N_2300);
xor U3999 (N_3999,N_2997,N_2987);
nand U4000 (N_4000,N_3848,N_3332);
and U4001 (N_4001,N_3226,N_3075);
nor U4002 (N_4002,N_3253,N_3961);
nand U4003 (N_4003,N_3880,N_3249);
xor U4004 (N_4004,N_3927,N_3658);
xor U4005 (N_4005,N_3959,N_3565);
nand U4006 (N_4006,N_3761,N_3200);
nor U4007 (N_4007,N_3909,N_3683);
xor U4008 (N_4008,N_3285,N_3214);
and U4009 (N_4009,N_3508,N_3888);
nor U4010 (N_4010,N_3279,N_3623);
xor U4011 (N_4011,N_3489,N_3059);
nor U4012 (N_4012,N_3600,N_3706);
nor U4013 (N_4013,N_3037,N_3762);
or U4014 (N_4014,N_3423,N_3187);
and U4015 (N_4015,N_3510,N_3447);
or U4016 (N_4016,N_3230,N_3188);
xor U4017 (N_4017,N_3719,N_3297);
xor U4018 (N_4018,N_3232,N_3984);
nor U4019 (N_4019,N_3399,N_3239);
or U4020 (N_4020,N_3671,N_3513);
nor U4021 (N_4021,N_3266,N_3060);
nor U4022 (N_4022,N_3550,N_3135);
or U4023 (N_4023,N_3735,N_3670);
or U4024 (N_4024,N_3713,N_3901);
and U4025 (N_4025,N_3672,N_3351);
or U4026 (N_4026,N_3331,N_3631);
or U4027 (N_4027,N_3234,N_3745);
nand U4028 (N_4028,N_3584,N_3988);
and U4029 (N_4029,N_3215,N_3580);
or U4030 (N_4030,N_3146,N_3841);
or U4031 (N_4031,N_3451,N_3291);
xor U4032 (N_4032,N_3524,N_3894);
xnor U4033 (N_4033,N_3324,N_3690);
xor U4034 (N_4034,N_3705,N_3979);
and U4035 (N_4035,N_3015,N_3852);
xor U4036 (N_4036,N_3669,N_3829);
and U4037 (N_4037,N_3117,N_3268);
nor U4038 (N_4038,N_3686,N_3620);
nor U4039 (N_4039,N_3677,N_3047);
xor U4040 (N_4040,N_3640,N_3070);
nand U4041 (N_4041,N_3098,N_3521);
nor U4042 (N_4042,N_3644,N_3471);
or U4043 (N_4043,N_3741,N_3042);
nor U4044 (N_4044,N_3664,N_3058);
or U4045 (N_4045,N_3743,N_3002);
nor U4046 (N_4046,N_3696,N_3845);
xor U4047 (N_4047,N_3595,N_3577);
and U4048 (N_4048,N_3914,N_3196);
nand U4049 (N_4049,N_3139,N_3405);
or U4050 (N_4050,N_3859,N_3803);
and U4051 (N_4051,N_3786,N_3320);
nand U4052 (N_4052,N_3081,N_3000);
nand U4053 (N_4053,N_3025,N_3121);
nor U4054 (N_4054,N_3211,N_3434);
and U4055 (N_4055,N_3474,N_3978);
nor U4056 (N_4056,N_3478,N_3290);
or U4057 (N_4057,N_3662,N_3828);
nand U4058 (N_4058,N_3906,N_3569);
nand U4059 (N_4059,N_3326,N_3077);
and U4060 (N_4060,N_3368,N_3406);
nand U4061 (N_4061,N_3892,N_3764);
and U4062 (N_4062,N_3468,N_3411);
or U4063 (N_4063,N_3364,N_3503);
xor U4064 (N_4064,N_3944,N_3744);
and U4065 (N_4065,N_3144,N_3344);
nor U4066 (N_4066,N_3821,N_3240);
nor U4067 (N_4067,N_3302,N_3907);
and U4068 (N_4068,N_3358,N_3768);
and U4069 (N_4069,N_3430,N_3955);
nor U4070 (N_4070,N_3052,N_3122);
xor U4071 (N_4071,N_3977,N_3257);
and U4072 (N_4072,N_3536,N_3053);
nand U4073 (N_4073,N_3572,N_3017);
xor U4074 (N_4074,N_3167,N_3209);
nand U4075 (N_4075,N_3023,N_3830);
and U4076 (N_4076,N_3881,N_3874);
xnor U4077 (N_4077,N_3793,N_3750);
and U4078 (N_4078,N_3490,N_3773);
and U4079 (N_4079,N_3723,N_3464);
xnor U4080 (N_4080,N_3221,N_3715);
nor U4081 (N_4081,N_3377,N_3061);
nand U4082 (N_4082,N_3816,N_3753);
nand U4083 (N_4083,N_3260,N_3805);
and U4084 (N_4084,N_3383,N_3031);
or U4085 (N_4085,N_3417,N_3124);
and U4086 (N_4086,N_3547,N_3854);
nor U4087 (N_4087,N_3030,N_3076);
nor U4088 (N_4088,N_3526,N_3137);
and U4089 (N_4089,N_3731,N_3292);
or U4090 (N_4090,N_3330,N_3783);
and U4091 (N_4091,N_3770,N_3225);
or U4092 (N_4092,N_3782,N_3428);
xnor U4093 (N_4093,N_3095,N_3817);
and U4094 (N_4094,N_3987,N_3767);
and U4095 (N_4095,N_3836,N_3827);
or U4096 (N_4096,N_3456,N_3748);
nor U4097 (N_4097,N_3610,N_3850);
and U4098 (N_4098,N_3591,N_3158);
nand U4099 (N_4099,N_3991,N_3790);
nor U4100 (N_4100,N_3376,N_3439);
nand U4101 (N_4101,N_3400,N_3995);
or U4102 (N_4102,N_3933,N_3866);
nand U4103 (N_4103,N_3651,N_3870);
or U4104 (N_4104,N_3908,N_3774);
nor U4105 (N_4105,N_3024,N_3616);
nand U4106 (N_4106,N_3523,N_3823);
nand U4107 (N_4107,N_3867,N_3804);
or U4108 (N_4108,N_3343,N_3083);
nor U4109 (N_4109,N_3420,N_3341);
nor U4110 (N_4110,N_3068,N_3375);
xnor U4111 (N_4111,N_3861,N_3974);
nand U4112 (N_4112,N_3179,N_3585);
or U4113 (N_4113,N_3262,N_3598);
and U4114 (N_4114,N_3414,N_3971);
and U4115 (N_4115,N_3578,N_3701);
nand U4116 (N_4116,N_3402,N_3919);
xor U4117 (N_4117,N_3111,N_3833);
nand U4118 (N_4118,N_3501,N_3967);
nor U4119 (N_4119,N_3448,N_3182);
nor U4120 (N_4120,N_3831,N_3877);
xnor U4121 (N_4121,N_3667,N_3599);
nor U4122 (N_4122,N_3084,N_3588);
nand U4123 (N_4123,N_3204,N_3732);
nor U4124 (N_4124,N_3635,N_3758);
nand U4125 (N_4125,N_3120,N_3647);
xnor U4126 (N_4126,N_3333,N_3717);
nand U4127 (N_4127,N_3739,N_3065);
nor U4128 (N_4128,N_3958,N_3632);
nor U4129 (N_4129,N_3655,N_3558);
and U4130 (N_4130,N_3794,N_3384);
nand U4131 (N_4131,N_3467,N_3224);
or U4132 (N_4132,N_3592,N_3033);
or U4133 (N_4133,N_3891,N_3582);
nand U4134 (N_4134,N_3756,N_3656);
nor U4135 (N_4135,N_3596,N_3528);
nor U4136 (N_4136,N_3839,N_3514);
nand U4137 (N_4137,N_3721,N_3163);
nand U4138 (N_4138,N_3294,N_3217);
xnor U4139 (N_4139,N_3286,N_3976);
xnor U4140 (N_4140,N_3601,N_3789);
or U4141 (N_4141,N_3028,N_3115);
or U4142 (N_4142,N_3304,N_3359);
or U4143 (N_4143,N_3273,N_3477);
or U4144 (N_4144,N_3872,N_3408);
or U4145 (N_4145,N_3079,N_3102);
and U4146 (N_4146,N_3488,N_3936);
and U4147 (N_4147,N_3512,N_3511);
or U4148 (N_4148,N_3010,N_3485);
and U4149 (N_4149,N_3777,N_3504);
and U4150 (N_4150,N_3493,N_3602);
xnor U4151 (N_4151,N_3825,N_3272);
or U4152 (N_4152,N_3553,N_3957);
xnor U4153 (N_4153,N_3624,N_3549);
xnor U4154 (N_4154,N_3530,N_3176);
or U4155 (N_4155,N_3155,N_3172);
or U4156 (N_4156,N_3012,N_3609);
and U4157 (N_4157,N_3818,N_3401);
nor U4158 (N_4158,N_3222,N_3537);
nand U4159 (N_4159,N_3943,N_3412);
and U4160 (N_4160,N_3787,N_3396);
nand U4161 (N_4161,N_3449,N_3245);
or U4162 (N_4162,N_3940,N_3100);
nor U4163 (N_4163,N_3844,N_3242);
nor U4164 (N_4164,N_3252,N_3022);
and U4165 (N_4165,N_3807,N_3551);
nor U4166 (N_4166,N_3150,N_3915);
and U4167 (N_4167,N_3265,N_3063);
xor U4168 (N_4168,N_3453,N_3676);
xor U4169 (N_4169,N_3295,N_3021);
nor U4170 (N_4170,N_3674,N_3785);
or U4171 (N_4171,N_3806,N_3161);
nand U4172 (N_4172,N_3563,N_3666);
nor U4173 (N_4173,N_3856,N_3296);
or U4174 (N_4174,N_3492,N_3751);
xor U4175 (N_4175,N_3173,N_3930);
nand U4176 (N_4176,N_3840,N_3973);
nand U4177 (N_4177,N_3863,N_3837);
xnor U4178 (N_4178,N_3085,N_3811);
or U4179 (N_4179,N_3244,N_3498);
xor U4180 (N_4180,N_3073,N_3246);
nand U4181 (N_4181,N_3050,N_3066);
nand U4182 (N_4182,N_3425,N_3048);
nand U4183 (N_4183,N_3939,N_3499);
nand U4184 (N_4184,N_3185,N_3890);
nand U4185 (N_4185,N_3484,N_3282);
or U4186 (N_4186,N_3847,N_3335);
and U4187 (N_4187,N_3634,N_3080);
and U4188 (N_4188,N_3727,N_3712);
xnor U4189 (N_4189,N_3328,N_3626);
nand U4190 (N_4190,N_3921,N_3308);
nor U4191 (N_4191,N_3809,N_3905);
nor U4192 (N_4192,N_3548,N_3231);
xor U4193 (N_4193,N_3878,N_3673);
or U4194 (N_4194,N_3440,N_3834);
and U4195 (N_4195,N_3757,N_3646);
nor U4196 (N_4196,N_3742,N_3795);
or U4197 (N_4197,N_3594,N_3394);
or U4198 (N_4198,N_3638,N_3057);
xor U4199 (N_4199,N_3966,N_3116);
nor U4200 (N_4200,N_3293,N_3149);
xnor U4201 (N_4201,N_3812,N_3882);
and U4202 (N_4202,N_3869,N_3665);
nor U4203 (N_4203,N_3347,N_3298);
nand U4204 (N_4204,N_3035,N_3661);
and U4205 (N_4205,N_3561,N_3926);
or U4206 (N_4206,N_3802,N_3636);
and U4207 (N_4207,N_3889,N_3051);
nor U4208 (N_4208,N_3032,N_3583);
nor U4209 (N_4209,N_3813,N_3250);
xor U4210 (N_4210,N_3317,N_3642);
and U4211 (N_4211,N_3476,N_3772);
nor U4212 (N_4212,N_3494,N_3018);
or U4213 (N_4213,N_3985,N_3645);
nor U4214 (N_4214,N_3233,N_3535);
nand U4215 (N_4215,N_3153,N_3119);
or U4216 (N_4216,N_3981,N_3996);
and U4217 (N_4217,N_3928,N_3784);
and U4218 (N_4218,N_3495,N_3746);
xor U4219 (N_4219,N_3082,N_3415);
nor U4220 (N_4220,N_3203,N_3473);
nor U4221 (N_4221,N_3067,N_3557);
or U4222 (N_4222,N_3165,N_3160);
or U4223 (N_4223,N_3339,N_3738);
nand U4224 (N_4224,N_3722,N_3127);
nor U4225 (N_4225,N_3897,N_3178);
nand U4226 (N_4226,N_3134,N_3353);
and U4227 (N_4227,N_3103,N_3615);
nor U4228 (N_4228,N_3113,N_3932);
nand U4229 (N_4229,N_3682,N_3797);
xor U4230 (N_4230,N_3539,N_3452);
and U4231 (N_4231,N_3444,N_3322);
and U4232 (N_4232,N_3952,N_3126);
or U4233 (N_4233,N_3019,N_3003);
nand U4234 (N_4234,N_3969,N_3092);
nor U4235 (N_4235,N_3641,N_3389);
or U4236 (N_4236,N_3431,N_3754);
nand U4237 (N_4237,N_3760,N_3049);
and U4238 (N_4238,N_3980,N_3518);
xor U4239 (N_4239,N_3419,N_3348);
or U4240 (N_4240,N_3532,N_3381);
or U4241 (N_4241,N_3029,N_3734);
nor U4242 (N_4242,N_3581,N_3469);
or U4243 (N_4243,N_3446,N_3154);
xor U4244 (N_4244,N_3393,N_3005);
nor U4245 (N_4245,N_3487,N_3462);
xnor U4246 (N_4246,N_3934,N_3857);
nor U4247 (N_4247,N_3574,N_3954);
or U4248 (N_4248,N_3953,N_3708);
xnor U4249 (N_4249,N_3680,N_3370);
and U4250 (N_4250,N_3109,N_3148);
xnor U4251 (N_4251,N_3258,N_3175);
xor U4252 (N_4252,N_3106,N_3107);
and U4253 (N_4253,N_3858,N_3479);
and U4254 (N_4254,N_3001,N_3788);
and U4255 (N_4255,N_3482,N_3422);
nor U4256 (N_4256,N_3710,N_3289);
and U4257 (N_4257,N_3733,N_3965);
xnor U4258 (N_4258,N_3781,N_3443);
and U4259 (N_4259,N_3895,N_3704);
nand U4260 (N_4260,N_3993,N_3612);
or U4261 (N_4261,N_3192,N_3131);
or U4262 (N_4262,N_3832,N_3517);
nand U4263 (N_4263,N_3392,N_3835);
nor U4264 (N_4264,N_3862,N_3189);
nor U4265 (N_4265,N_3929,N_3147);
nor U4266 (N_4266,N_3014,N_3949);
nand U4267 (N_4267,N_3792,N_3034);
xnor U4268 (N_4268,N_3931,N_3718);
or U4269 (N_4269,N_3303,N_3605);
nand U4270 (N_4270,N_3278,N_3055);
xnor U4271 (N_4271,N_3212,N_3086);
and U4272 (N_4272,N_3367,N_3301);
xor U4273 (N_4273,N_3455,N_3555);
or U4274 (N_4274,N_3432,N_3181);
xor U4275 (N_4275,N_3305,N_3261);
xor U4276 (N_4276,N_3218,N_3685);
nor U4277 (N_4277,N_3207,N_3737);
nand U4278 (N_4278,N_3648,N_3195);
xor U4279 (N_4279,N_3445,N_3128);
xor U4280 (N_4280,N_3300,N_3824);
or U4281 (N_4281,N_3654,N_3287);
nor U4282 (N_4282,N_3660,N_3608);
and U4283 (N_4283,N_3227,N_3194);
nand U4284 (N_4284,N_3184,N_3540);
xnor U4285 (N_4285,N_3156,N_3069);
and U4286 (N_4286,N_3164,N_3045);
nand U4287 (N_4287,N_3091,N_3639);
nand U4288 (N_4288,N_3763,N_3938);
nor U4289 (N_4289,N_3472,N_3519);
nand U4290 (N_4290,N_3433,N_3129);
or U4291 (N_4291,N_3288,N_3500);
xor U4292 (N_4292,N_3141,N_3779);
xnor U4293 (N_4293,N_3720,N_3275);
xnor U4294 (N_4294,N_3505,N_3570);
and U4295 (N_4295,N_3114,N_3791);
nand U4296 (N_4296,N_3334,N_3235);
or U4297 (N_4297,N_3459,N_3123);
nand U4298 (N_4298,N_3691,N_3403);
nor U4299 (N_4299,N_3177,N_3284);
and U4300 (N_4300,N_3887,N_3418);
and U4301 (N_4301,N_3820,N_3649);
xnor U4302 (N_4302,N_3509,N_3590);
nand U4303 (N_4303,N_3964,N_3992);
nand U4304 (N_4304,N_3314,N_3140);
and U4305 (N_4305,N_3228,N_3917);
or U4306 (N_4306,N_3559,N_3264);
nor U4307 (N_4307,N_3946,N_3798);
nand U4308 (N_4308,N_3088,N_3956);
xor U4309 (N_4309,N_3345,N_3920);
and U4310 (N_4310,N_3263,N_3810);
and U4311 (N_4311,N_3545,N_3143);
nand U4312 (N_4312,N_3404,N_3349);
nand U4313 (N_4313,N_3619,N_3999);
xor U4314 (N_4314,N_3243,N_3986);
or U4315 (N_4315,N_3714,N_3587);
or U4316 (N_4316,N_3950,N_3046);
or U4317 (N_4317,N_3759,N_3819);
nand U4318 (N_4318,N_3883,N_3573);
xor U4319 (N_4319,N_3925,N_3363);
nor U4320 (N_4320,N_3982,N_3617);
or U4321 (N_4321,N_3884,N_3520);
nor U4322 (N_4322,N_3271,N_3483);
or U4323 (N_4323,N_3313,N_3145);
and U4324 (N_4324,N_3397,N_3752);
and U4325 (N_4325,N_3766,N_3997);
or U4326 (N_4326,N_3475,N_3062);
nor U4327 (N_4327,N_3538,N_3597);
or U4328 (N_4328,N_3480,N_3277);
and U4329 (N_4329,N_3593,N_3366);
or U4330 (N_4330,N_3251,N_3998);
nor U4331 (N_4331,N_3316,N_3603);
nand U4332 (N_4332,N_3210,N_3340);
nand U4333 (N_4333,N_3096,N_3202);
nor U4334 (N_4334,N_3373,N_3637);
or U4335 (N_4335,N_3311,N_3703);
xor U4336 (N_4336,N_3778,N_3910);
nor U4337 (N_4337,N_3441,N_3390);
or U4338 (N_4338,N_3044,N_3541);
nor U4339 (N_4339,N_3369,N_3281);
nor U4340 (N_4340,N_3924,N_3942);
nor U4341 (N_4341,N_3698,N_3554);
and U4342 (N_4342,N_3438,N_3435);
xor U4343 (N_4343,N_3918,N_3410);
or U4344 (N_4344,N_3709,N_3531);
nor U4345 (N_4345,N_3579,N_3138);
nand U4346 (N_4346,N_3198,N_3653);
nor U4347 (N_4347,N_3206,N_3650);
nand U4348 (N_4348,N_3566,N_3112);
or U4349 (N_4349,N_3975,N_3372);
xnor U4350 (N_4350,N_3454,N_3516);
nor U4351 (N_4351,N_3568,N_3142);
or U4352 (N_4352,N_3157,N_3885);
nand U4353 (N_4353,N_3436,N_3913);
nor U4354 (N_4354,N_3355,N_3460);
nand U4355 (N_4355,N_3694,N_3007);
and U4356 (N_4356,N_3556,N_3534);
nand U4357 (N_4357,N_3038,N_3470);
and U4358 (N_4358,N_3151,N_3327);
xnor U4359 (N_4359,N_3219,N_3527);
xnor U4360 (N_4360,N_3507,N_3801);
nand U4361 (N_4361,N_3989,N_3255);
xor U4362 (N_4362,N_3630,N_3174);
and U4363 (N_4363,N_3357,N_3220);
and U4364 (N_4364,N_3170,N_3216);
nand U4365 (N_4365,N_3575,N_3197);
and U4366 (N_4366,N_3533,N_3416);
nor U4367 (N_4367,N_3171,N_3497);
or U4368 (N_4368,N_3016,N_3380);
or U4369 (N_4369,N_3087,N_3108);
nand U4370 (N_4370,N_3962,N_3398);
nor U4371 (N_4371,N_3097,N_3522);
or U4372 (N_4372,N_3871,N_3183);
nor U4373 (N_4373,N_3481,N_3132);
or U4374 (N_4374,N_3873,N_3385);
nor U4375 (N_4375,N_3621,N_3900);
or U4376 (N_4376,N_3702,N_3502);
xnor U4377 (N_4377,N_3688,N_3486);
nor U4378 (N_4378,N_3796,N_3697);
xnor U4379 (N_4379,N_3699,N_3089);
xnor U4380 (N_4380,N_3618,N_3090);
nor U4381 (N_4381,N_3544,N_3896);
or U4382 (N_4382,N_3983,N_3945);
and U4383 (N_4383,N_3633,N_3201);
xnor U4384 (N_4384,N_3728,N_3011);
nand U4385 (N_4385,N_3668,N_3152);
nand U4386 (N_4386,N_3379,N_3684);
nor U4387 (N_4387,N_3681,N_3749);
nand U4388 (N_4388,N_3361,N_3104);
or U4389 (N_4389,N_3315,N_3923);
and U4390 (N_4390,N_3276,N_3611);
nor U4391 (N_4391,N_3947,N_3136);
or U4392 (N_4392,N_3236,N_3564);
or U4393 (N_4393,N_3130,N_3360);
and U4394 (N_4394,N_3238,N_3094);
xor U4395 (N_4395,N_3855,N_3838);
and U4396 (N_4396,N_3338,N_3299);
and U4397 (N_4397,N_3450,N_3695);
xor U4398 (N_4398,N_3799,N_3054);
nand U4399 (N_4399,N_3237,N_3571);
or U4400 (N_4400,N_3254,N_3562);
nor U4401 (N_4401,N_3166,N_3625);
or U4402 (N_4402,N_3280,N_3409);
nand U4403 (N_4403,N_3186,N_3628);
nand U4404 (N_4404,N_3716,N_3576);
nand U4405 (N_4405,N_3711,N_3865);
nand U4406 (N_4406,N_3365,N_3849);
nor U4407 (N_4407,N_3769,N_3466);
xnor U4408 (N_4408,N_3008,N_3356);
nor U4409 (N_4409,N_3072,N_3125);
nor U4410 (N_4410,N_3162,N_3442);
or U4411 (N_4411,N_3169,N_3318);
and U4412 (N_4412,N_3529,N_3604);
nand U4413 (N_4413,N_3860,N_3110);
xnor U4414 (N_4414,N_3006,N_3378);
and U4415 (N_4415,N_3013,N_3325);
nand U4416 (N_4416,N_3004,N_3730);
nand U4417 (N_4417,N_3105,N_3729);
xnor U4418 (N_4418,N_3724,N_3319);
and U4419 (N_4419,N_3362,N_3463);
or U4420 (N_4420,N_3118,N_3627);
nor U4421 (N_4421,N_3321,N_3815);
and U4422 (N_4422,N_3643,N_3205);
xor U4423 (N_4423,N_3168,N_3851);
nand U4424 (N_4424,N_3354,N_3826);
nor U4425 (N_4425,N_3903,N_3199);
nand U4426 (N_4426,N_3413,N_3270);
or U4427 (N_4427,N_3342,N_3159);
or U4428 (N_4428,N_3458,N_3248);
nand U4429 (N_4429,N_3941,N_3267);
or U4430 (N_4430,N_3629,N_3613);
nor U4431 (N_4431,N_3968,N_3606);
nand U4432 (N_4432,N_3496,N_3960);
nand U4433 (N_4433,N_3336,N_3657);
xnor U4434 (N_4434,N_3391,N_3274);
or U4435 (N_4435,N_3241,N_3382);
nand U4436 (N_4436,N_3780,N_3622);
or U4437 (N_4437,N_3190,N_3027);
nor U4438 (N_4438,N_3309,N_3310);
or U4439 (N_4439,N_3922,N_3323);
or U4440 (N_4440,N_3026,N_3879);
or U4441 (N_4441,N_3371,N_3306);
or U4442 (N_4442,N_3071,N_3040);
nor U4443 (N_4443,N_3388,N_3427);
nor U4444 (N_4444,N_3678,N_3994);
xor U4445 (N_4445,N_3948,N_3036);
nand U4446 (N_4446,N_3064,N_3970);
and U4447 (N_4447,N_3374,N_3099);
and U4448 (N_4448,N_3679,N_3093);
nor U4449 (N_4449,N_3213,N_3307);
nor U4450 (N_4450,N_3337,N_3912);
and U4451 (N_4451,N_3771,N_3800);
nor U4452 (N_4452,N_3589,N_3614);
xnor U4453 (N_4453,N_3457,N_3972);
nand U4454 (N_4454,N_3937,N_3546);
and U4455 (N_4455,N_3853,N_3009);
xnor U4456 (N_4456,N_3726,N_3893);
and U4457 (N_4457,N_3101,N_3843);
nor U4458 (N_4458,N_3133,N_3747);
xnor U4459 (N_4459,N_3607,N_3056);
xnor U4460 (N_4460,N_3515,N_3543);
nand U4461 (N_4461,N_3350,N_3560);
nand U4462 (N_4462,N_3552,N_3041);
or U4463 (N_4463,N_3814,N_3689);
and U4464 (N_4464,N_3461,N_3765);
and U4465 (N_4465,N_3755,N_3191);
or U4466 (N_4466,N_3525,N_3386);
nor U4467 (N_4467,N_3707,N_3842);
nor U4468 (N_4468,N_3424,N_3911);
or U4469 (N_4469,N_3675,N_3346);
nor U4470 (N_4470,N_3822,N_3808);
xor U4471 (N_4471,N_3567,N_3352);
or U4472 (N_4472,N_3269,N_3687);
nand U4473 (N_4473,N_3693,N_3876);
xnor U4474 (N_4474,N_3692,N_3043);
nor U4475 (N_4475,N_3387,N_3775);
xor U4476 (N_4476,N_3899,N_3256);
nor U4477 (N_4477,N_3542,N_3990);
nor U4478 (N_4478,N_3659,N_3663);
and U4479 (N_4479,N_3465,N_3078);
nor U4480 (N_4480,N_3247,N_3963);
nor U4481 (N_4481,N_3421,N_3846);
or U4482 (N_4482,N_3736,N_3437);
and U4483 (N_4483,N_3429,N_3039);
xnor U4484 (N_4484,N_3916,N_3886);
xnor U4485 (N_4485,N_3407,N_3725);
and U4486 (N_4486,N_3491,N_3935);
nor U4487 (N_4487,N_3875,N_3864);
or U4488 (N_4488,N_3259,N_3312);
nor U4489 (N_4489,N_3898,N_3776);
nor U4490 (N_4490,N_3740,N_3223);
nor U4491 (N_4491,N_3426,N_3700);
xor U4492 (N_4492,N_3902,N_3193);
and U4493 (N_4493,N_3506,N_3329);
nor U4494 (N_4494,N_3020,N_3395);
xnor U4495 (N_4495,N_3904,N_3208);
nand U4496 (N_4496,N_3229,N_3283);
xor U4497 (N_4497,N_3652,N_3951);
and U4498 (N_4498,N_3074,N_3586);
nand U4499 (N_4499,N_3180,N_3868);
xor U4500 (N_4500,N_3233,N_3398);
nor U4501 (N_4501,N_3853,N_3814);
nor U4502 (N_4502,N_3980,N_3204);
or U4503 (N_4503,N_3016,N_3700);
nand U4504 (N_4504,N_3987,N_3682);
or U4505 (N_4505,N_3923,N_3208);
nand U4506 (N_4506,N_3039,N_3768);
and U4507 (N_4507,N_3398,N_3725);
nand U4508 (N_4508,N_3444,N_3681);
xor U4509 (N_4509,N_3944,N_3088);
or U4510 (N_4510,N_3664,N_3553);
nand U4511 (N_4511,N_3468,N_3465);
and U4512 (N_4512,N_3311,N_3590);
nor U4513 (N_4513,N_3111,N_3364);
xnor U4514 (N_4514,N_3735,N_3931);
and U4515 (N_4515,N_3549,N_3309);
nor U4516 (N_4516,N_3675,N_3900);
or U4517 (N_4517,N_3506,N_3195);
and U4518 (N_4518,N_3717,N_3944);
and U4519 (N_4519,N_3364,N_3385);
nor U4520 (N_4520,N_3117,N_3609);
nor U4521 (N_4521,N_3253,N_3430);
xnor U4522 (N_4522,N_3110,N_3415);
nand U4523 (N_4523,N_3786,N_3837);
or U4524 (N_4524,N_3382,N_3468);
and U4525 (N_4525,N_3960,N_3324);
nor U4526 (N_4526,N_3118,N_3261);
nand U4527 (N_4527,N_3939,N_3494);
and U4528 (N_4528,N_3352,N_3744);
nor U4529 (N_4529,N_3332,N_3486);
nor U4530 (N_4530,N_3933,N_3594);
and U4531 (N_4531,N_3596,N_3025);
xor U4532 (N_4532,N_3742,N_3618);
nor U4533 (N_4533,N_3431,N_3095);
xnor U4534 (N_4534,N_3741,N_3661);
and U4535 (N_4535,N_3137,N_3300);
or U4536 (N_4536,N_3338,N_3307);
or U4537 (N_4537,N_3943,N_3041);
xnor U4538 (N_4538,N_3361,N_3407);
nor U4539 (N_4539,N_3505,N_3015);
nand U4540 (N_4540,N_3536,N_3633);
xor U4541 (N_4541,N_3605,N_3841);
or U4542 (N_4542,N_3596,N_3632);
or U4543 (N_4543,N_3052,N_3528);
xnor U4544 (N_4544,N_3628,N_3716);
and U4545 (N_4545,N_3381,N_3917);
nor U4546 (N_4546,N_3864,N_3455);
nor U4547 (N_4547,N_3865,N_3874);
and U4548 (N_4548,N_3427,N_3617);
or U4549 (N_4549,N_3853,N_3298);
xor U4550 (N_4550,N_3254,N_3754);
or U4551 (N_4551,N_3910,N_3445);
xnor U4552 (N_4552,N_3024,N_3151);
nand U4553 (N_4553,N_3711,N_3274);
and U4554 (N_4554,N_3459,N_3440);
and U4555 (N_4555,N_3593,N_3725);
nor U4556 (N_4556,N_3032,N_3728);
nor U4557 (N_4557,N_3499,N_3958);
or U4558 (N_4558,N_3913,N_3019);
and U4559 (N_4559,N_3509,N_3057);
xnor U4560 (N_4560,N_3325,N_3520);
or U4561 (N_4561,N_3131,N_3992);
and U4562 (N_4562,N_3024,N_3084);
xnor U4563 (N_4563,N_3044,N_3762);
nand U4564 (N_4564,N_3244,N_3120);
nor U4565 (N_4565,N_3281,N_3225);
or U4566 (N_4566,N_3744,N_3068);
nand U4567 (N_4567,N_3166,N_3394);
nand U4568 (N_4568,N_3252,N_3444);
and U4569 (N_4569,N_3570,N_3294);
or U4570 (N_4570,N_3824,N_3183);
and U4571 (N_4571,N_3689,N_3015);
or U4572 (N_4572,N_3519,N_3395);
xnor U4573 (N_4573,N_3215,N_3376);
nor U4574 (N_4574,N_3377,N_3375);
and U4575 (N_4575,N_3308,N_3883);
nor U4576 (N_4576,N_3021,N_3679);
and U4577 (N_4577,N_3418,N_3857);
or U4578 (N_4578,N_3722,N_3427);
and U4579 (N_4579,N_3141,N_3647);
and U4580 (N_4580,N_3352,N_3817);
xnor U4581 (N_4581,N_3643,N_3369);
nand U4582 (N_4582,N_3375,N_3883);
xor U4583 (N_4583,N_3574,N_3139);
nand U4584 (N_4584,N_3064,N_3679);
or U4585 (N_4585,N_3385,N_3903);
xor U4586 (N_4586,N_3340,N_3050);
nand U4587 (N_4587,N_3854,N_3049);
nor U4588 (N_4588,N_3978,N_3499);
or U4589 (N_4589,N_3058,N_3433);
xor U4590 (N_4590,N_3579,N_3285);
or U4591 (N_4591,N_3900,N_3594);
nor U4592 (N_4592,N_3846,N_3697);
or U4593 (N_4593,N_3063,N_3832);
or U4594 (N_4594,N_3492,N_3684);
or U4595 (N_4595,N_3066,N_3016);
or U4596 (N_4596,N_3538,N_3696);
nand U4597 (N_4597,N_3038,N_3296);
xnor U4598 (N_4598,N_3225,N_3501);
nand U4599 (N_4599,N_3132,N_3960);
xor U4600 (N_4600,N_3994,N_3744);
xor U4601 (N_4601,N_3572,N_3069);
or U4602 (N_4602,N_3347,N_3148);
and U4603 (N_4603,N_3348,N_3998);
nor U4604 (N_4604,N_3865,N_3089);
and U4605 (N_4605,N_3224,N_3209);
nand U4606 (N_4606,N_3705,N_3074);
or U4607 (N_4607,N_3231,N_3431);
or U4608 (N_4608,N_3980,N_3442);
xnor U4609 (N_4609,N_3861,N_3918);
xor U4610 (N_4610,N_3786,N_3411);
nor U4611 (N_4611,N_3702,N_3048);
and U4612 (N_4612,N_3459,N_3577);
and U4613 (N_4613,N_3928,N_3630);
and U4614 (N_4614,N_3952,N_3899);
nand U4615 (N_4615,N_3858,N_3908);
or U4616 (N_4616,N_3443,N_3344);
and U4617 (N_4617,N_3139,N_3786);
and U4618 (N_4618,N_3490,N_3875);
nand U4619 (N_4619,N_3343,N_3010);
nand U4620 (N_4620,N_3086,N_3162);
and U4621 (N_4621,N_3489,N_3708);
xor U4622 (N_4622,N_3231,N_3079);
nand U4623 (N_4623,N_3306,N_3767);
or U4624 (N_4624,N_3238,N_3438);
or U4625 (N_4625,N_3322,N_3395);
nor U4626 (N_4626,N_3725,N_3238);
xnor U4627 (N_4627,N_3243,N_3526);
nand U4628 (N_4628,N_3882,N_3056);
xnor U4629 (N_4629,N_3401,N_3836);
xnor U4630 (N_4630,N_3296,N_3504);
nor U4631 (N_4631,N_3615,N_3775);
or U4632 (N_4632,N_3808,N_3395);
or U4633 (N_4633,N_3046,N_3041);
and U4634 (N_4634,N_3738,N_3884);
xor U4635 (N_4635,N_3515,N_3443);
nor U4636 (N_4636,N_3575,N_3009);
nand U4637 (N_4637,N_3572,N_3596);
nor U4638 (N_4638,N_3004,N_3487);
nand U4639 (N_4639,N_3590,N_3952);
xnor U4640 (N_4640,N_3965,N_3785);
nand U4641 (N_4641,N_3247,N_3752);
or U4642 (N_4642,N_3586,N_3452);
and U4643 (N_4643,N_3038,N_3773);
xnor U4644 (N_4644,N_3845,N_3385);
nor U4645 (N_4645,N_3979,N_3956);
nand U4646 (N_4646,N_3305,N_3866);
and U4647 (N_4647,N_3565,N_3509);
or U4648 (N_4648,N_3168,N_3816);
nand U4649 (N_4649,N_3484,N_3064);
nand U4650 (N_4650,N_3723,N_3949);
nand U4651 (N_4651,N_3970,N_3404);
or U4652 (N_4652,N_3728,N_3818);
nand U4653 (N_4653,N_3459,N_3979);
nor U4654 (N_4654,N_3889,N_3185);
and U4655 (N_4655,N_3187,N_3720);
and U4656 (N_4656,N_3906,N_3948);
nand U4657 (N_4657,N_3903,N_3667);
or U4658 (N_4658,N_3864,N_3536);
and U4659 (N_4659,N_3689,N_3428);
or U4660 (N_4660,N_3497,N_3259);
nor U4661 (N_4661,N_3160,N_3566);
xor U4662 (N_4662,N_3647,N_3770);
and U4663 (N_4663,N_3932,N_3697);
or U4664 (N_4664,N_3633,N_3695);
nor U4665 (N_4665,N_3193,N_3402);
xor U4666 (N_4666,N_3613,N_3869);
nand U4667 (N_4667,N_3479,N_3865);
nor U4668 (N_4668,N_3672,N_3741);
or U4669 (N_4669,N_3745,N_3850);
nor U4670 (N_4670,N_3195,N_3534);
and U4671 (N_4671,N_3007,N_3677);
xor U4672 (N_4672,N_3101,N_3418);
or U4673 (N_4673,N_3846,N_3406);
nand U4674 (N_4674,N_3357,N_3667);
nand U4675 (N_4675,N_3314,N_3202);
nand U4676 (N_4676,N_3687,N_3697);
or U4677 (N_4677,N_3954,N_3554);
nor U4678 (N_4678,N_3729,N_3663);
nand U4679 (N_4679,N_3072,N_3063);
nor U4680 (N_4680,N_3617,N_3666);
nor U4681 (N_4681,N_3109,N_3806);
nand U4682 (N_4682,N_3846,N_3537);
nand U4683 (N_4683,N_3568,N_3880);
nand U4684 (N_4684,N_3826,N_3887);
or U4685 (N_4685,N_3398,N_3777);
nand U4686 (N_4686,N_3849,N_3067);
xnor U4687 (N_4687,N_3753,N_3623);
xor U4688 (N_4688,N_3447,N_3921);
xnor U4689 (N_4689,N_3797,N_3002);
xnor U4690 (N_4690,N_3316,N_3946);
nor U4691 (N_4691,N_3826,N_3764);
nor U4692 (N_4692,N_3753,N_3262);
xnor U4693 (N_4693,N_3669,N_3698);
nor U4694 (N_4694,N_3381,N_3121);
and U4695 (N_4695,N_3149,N_3374);
xor U4696 (N_4696,N_3423,N_3332);
and U4697 (N_4697,N_3875,N_3838);
or U4698 (N_4698,N_3376,N_3417);
nor U4699 (N_4699,N_3298,N_3821);
xnor U4700 (N_4700,N_3364,N_3477);
nor U4701 (N_4701,N_3322,N_3172);
nor U4702 (N_4702,N_3485,N_3942);
and U4703 (N_4703,N_3715,N_3626);
nand U4704 (N_4704,N_3248,N_3666);
nor U4705 (N_4705,N_3646,N_3065);
and U4706 (N_4706,N_3145,N_3422);
nand U4707 (N_4707,N_3516,N_3044);
or U4708 (N_4708,N_3473,N_3712);
nand U4709 (N_4709,N_3281,N_3863);
nor U4710 (N_4710,N_3527,N_3456);
xnor U4711 (N_4711,N_3105,N_3053);
and U4712 (N_4712,N_3682,N_3831);
xor U4713 (N_4713,N_3781,N_3409);
nand U4714 (N_4714,N_3905,N_3082);
nor U4715 (N_4715,N_3689,N_3127);
nand U4716 (N_4716,N_3937,N_3515);
nand U4717 (N_4717,N_3012,N_3615);
xor U4718 (N_4718,N_3194,N_3829);
nand U4719 (N_4719,N_3653,N_3134);
or U4720 (N_4720,N_3084,N_3515);
and U4721 (N_4721,N_3127,N_3880);
nor U4722 (N_4722,N_3689,N_3112);
nor U4723 (N_4723,N_3779,N_3777);
nand U4724 (N_4724,N_3749,N_3459);
and U4725 (N_4725,N_3716,N_3493);
or U4726 (N_4726,N_3521,N_3216);
nor U4727 (N_4727,N_3171,N_3803);
xor U4728 (N_4728,N_3348,N_3938);
xnor U4729 (N_4729,N_3855,N_3578);
nand U4730 (N_4730,N_3574,N_3218);
nor U4731 (N_4731,N_3062,N_3102);
and U4732 (N_4732,N_3389,N_3496);
nor U4733 (N_4733,N_3246,N_3926);
and U4734 (N_4734,N_3025,N_3090);
and U4735 (N_4735,N_3423,N_3206);
or U4736 (N_4736,N_3857,N_3527);
or U4737 (N_4737,N_3576,N_3631);
and U4738 (N_4738,N_3422,N_3439);
nand U4739 (N_4739,N_3943,N_3188);
nor U4740 (N_4740,N_3799,N_3624);
or U4741 (N_4741,N_3886,N_3210);
or U4742 (N_4742,N_3370,N_3324);
nand U4743 (N_4743,N_3926,N_3500);
xor U4744 (N_4744,N_3739,N_3843);
nor U4745 (N_4745,N_3736,N_3797);
xnor U4746 (N_4746,N_3345,N_3823);
xnor U4747 (N_4747,N_3923,N_3443);
nor U4748 (N_4748,N_3538,N_3154);
nand U4749 (N_4749,N_3788,N_3148);
nor U4750 (N_4750,N_3800,N_3606);
nand U4751 (N_4751,N_3276,N_3443);
nor U4752 (N_4752,N_3516,N_3724);
nand U4753 (N_4753,N_3347,N_3348);
xnor U4754 (N_4754,N_3436,N_3996);
nand U4755 (N_4755,N_3251,N_3111);
xor U4756 (N_4756,N_3083,N_3305);
nor U4757 (N_4757,N_3742,N_3120);
or U4758 (N_4758,N_3697,N_3642);
and U4759 (N_4759,N_3694,N_3911);
nand U4760 (N_4760,N_3641,N_3681);
and U4761 (N_4761,N_3856,N_3365);
and U4762 (N_4762,N_3278,N_3283);
nand U4763 (N_4763,N_3424,N_3270);
or U4764 (N_4764,N_3982,N_3838);
or U4765 (N_4765,N_3294,N_3953);
nor U4766 (N_4766,N_3707,N_3051);
and U4767 (N_4767,N_3547,N_3257);
nor U4768 (N_4768,N_3514,N_3271);
nand U4769 (N_4769,N_3640,N_3726);
xnor U4770 (N_4770,N_3376,N_3159);
or U4771 (N_4771,N_3651,N_3489);
xor U4772 (N_4772,N_3318,N_3909);
or U4773 (N_4773,N_3579,N_3290);
xnor U4774 (N_4774,N_3663,N_3930);
or U4775 (N_4775,N_3268,N_3170);
xnor U4776 (N_4776,N_3611,N_3629);
or U4777 (N_4777,N_3965,N_3586);
and U4778 (N_4778,N_3919,N_3171);
nand U4779 (N_4779,N_3182,N_3872);
and U4780 (N_4780,N_3935,N_3431);
nor U4781 (N_4781,N_3229,N_3294);
xnor U4782 (N_4782,N_3659,N_3781);
nand U4783 (N_4783,N_3171,N_3636);
and U4784 (N_4784,N_3345,N_3424);
xor U4785 (N_4785,N_3856,N_3873);
xor U4786 (N_4786,N_3313,N_3686);
nand U4787 (N_4787,N_3707,N_3086);
nand U4788 (N_4788,N_3750,N_3807);
and U4789 (N_4789,N_3866,N_3364);
or U4790 (N_4790,N_3475,N_3435);
xor U4791 (N_4791,N_3716,N_3712);
nor U4792 (N_4792,N_3174,N_3026);
and U4793 (N_4793,N_3008,N_3524);
xnor U4794 (N_4794,N_3538,N_3203);
nand U4795 (N_4795,N_3658,N_3682);
or U4796 (N_4796,N_3238,N_3983);
xnor U4797 (N_4797,N_3642,N_3282);
xor U4798 (N_4798,N_3153,N_3641);
nor U4799 (N_4799,N_3682,N_3436);
or U4800 (N_4800,N_3300,N_3481);
nor U4801 (N_4801,N_3246,N_3123);
nor U4802 (N_4802,N_3823,N_3806);
xor U4803 (N_4803,N_3279,N_3826);
or U4804 (N_4804,N_3978,N_3727);
nor U4805 (N_4805,N_3391,N_3583);
and U4806 (N_4806,N_3396,N_3678);
or U4807 (N_4807,N_3073,N_3925);
nor U4808 (N_4808,N_3659,N_3197);
nand U4809 (N_4809,N_3351,N_3931);
xor U4810 (N_4810,N_3374,N_3429);
nor U4811 (N_4811,N_3236,N_3360);
or U4812 (N_4812,N_3872,N_3064);
and U4813 (N_4813,N_3011,N_3592);
nor U4814 (N_4814,N_3120,N_3651);
xnor U4815 (N_4815,N_3796,N_3486);
or U4816 (N_4816,N_3880,N_3166);
nor U4817 (N_4817,N_3372,N_3779);
nor U4818 (N_4818,N_3442,N_3971);
nand U4819 (N_4819,N_3461,N_3145);
nor U4820 (N_4820,N_3358,N_3867);
nor U4821 (N_4821,N_3477,N_3708);
or U4822 (N_4822,N_3687,N_3644);
and U4823 (N_4823,N_3423,N_3628);
nand U4824 (N_4824,N_3134,N_3410);
nand U4825 (N_4825,N_3623,N_3084);
and U4826 (N_4826,N_3367,N_3588);
nor U4827 (N_4827,N_3067,N_3355);
nor U4828 (N_4828,N_3260,N_3952);
nor U4829 (N_4829,N_3704,N_3451);
nand U4830 (N_4830,N_3689,N_3010);
nand U4831 (N_4831,N_3406,N_3879);
xor U4832 (N_4832,N_3496,N_3948);
nand U4833 (N_4833,N_3037,N_3538);
nor U4834 (N_4834,N_3209,N_3060);
xor U4835 (N_4835,N_3074,N_3905);
or U4836 (N_4836,N_3354,N_3394);
and U4837 (N_4837,N_3016,N_3564);
nand U4838 (N_4838,N_3306,N_3734);
nand U4839 (N_4839,N_3674,N_3693);
nand U4840 (N_4840,N_3565,N_3009);
and U4841 (N_4841,N_3905,N_3715);
or U4842 (N_4842,N_3347,N_3181);
nor U4843 (N_4843,N_3599,N_3589);
xnor U4844 (N_4844,N_3213,N_3752);
xor U4845 (N_4845,N_3367,N_3717);
nand U4846 (N_4846,N_3315,N_3595);
xor U4847 (N_4847,N_3083,N_3560);
or U4848 (N_4848,N_3129,N_3728);
or U4849 (N_4849,N_3367,N_3869);
nor U4850 (N_4850,N_3406,N_3343);
xor U4851 (N_4851,N_3387,N_3979);
or U4852 (N_4852,N_3642,N_3283);
and U4853 (N_4853,N_3086,N_3529);
or U4854 (N_4854,N_3987,N_3604);
or U4855 (N_4855,N_3389,N_3532);
xor U4856 (N_4856,N_3472,N_3658);
and U4857 (N_4857,N_3678,N_3060);
nor U4858 (N_4858,N_3170,N_3350);
nor U4859 (N_4859,N_3193,N_3029);
xor U4860 (N_4860,N_3244,N_3398);
or U4861 (N_4861,N_3387,N_3983);
nand U4862 (N_4862,N_3970,N_3589);
or U4863 (N_4863,N_3853,N_3042);
xor U4864 (N_4864,N_3766,N_3455);
or U4865 (N_4865,N_3732,N_3401);
nand U4866 (N_4866,N_3638,N_3359);
or U4867 (N_4867,N_3687,N_3931);
nor U4868 (N_4868,N_3023,N_3273);
nand U4869 (N_4869,N_3692,N_3165);
nand U4870 (N_4870,N_3088,N_3821);
nor U4871 (N_4871,N_3559,N_3938);
nor U4872 (N_4872,N_3140,N_3284);
or U4873 (N_4873,N_3222,N_3146);
nand U4874 (N_4874,N_3089,N_3229);
nand U4875 (N_4875,N_3496,N_3256);
and U4876 (N_4876,N_3297,N_3305);
nor U4877 (N_4877,N_3178,N_3780);
or U4878 (N_4878,N_3576,N_3491);
nor U4879 (N_4879,N_3303,N_3434);
xor U4880 (N_4880,N_3297,N_3541);
or U4881 (N_4881,N_3821,N_3788);
nor U4882 (N_4882,N_3089,N_3205);
or U4883 (N_4883,N_3735,N_3703);
xnor U4884 (N_4884,N_3359,N_3315);
and U4885 (N_4885,N_3317,N_3349);
xnor U4886 (N_4886,N_3886,N_3386);
xor U4887 (N_4887,N_3516,N_3224);
nor U4888 (N_4888,N_3473,N_3984);
nand U4889 (N_4889,N_3868,N_3929);
or U4890 (N_4890,N_3914,N_3351);
or U4891 (N_4891,N_3349,N_3855);
or U4892 (N_4892,N_3515,N_3705);
or U4893 (N_4893,N_3609,N_3480);
or U4894 (N_4894,N_3870,N_3945);
xor U4895 (N_4895,N_3689,N_3279);
nand U4896 (N_4896,N_3440,N_3408);
and U4897 (N_4897,N_3071,N_3924);
xor U4898 (N_4898,N_3075,N_3328);
nand U4899 (N_4899,N_3945,N_3931);
and U4900 (N_4900,N_3145,N_3025);
or U4901 (N_4901,N_3211,N_3957);
or U4902 (N_4902,N_3421,N_3997);
xor U4903 (N_4903,N_3551,N_3839);
nor U4904 (N_4904,N_3265,N_3417);
nor U4905 (N_4905,N_3832,N_3477);
nor U4906 (N_4906,N_3439,N_3614);
or U4907 (N_4907,N_3267,N_3977);
xor U4908 (N_4908,N_3919,N_3380);
and U4909 (N_4909,N_3641,N_3215);
nor U4910 (N_4910,N_3312,N_3384);
xor U4911 (N_4911,N_3455,N_3021);
xor U4912 (N_4912,N_3786,N_3517);
or U4913 (N_4913,N_3403,N_3004);
xnor U4914 (N_4914,N_3783,N_3881);
nand U4915 (N_4915,N_3023,N_3013);
and U4916 (N_4916,N_3641,N_3492);
nand U4917 (N_4917,N_3087,N_3507);
nor U4918 (N_4918,N_3582,N_3230);
or U4919 (N_4919,N_3509,N_3145);
xor U4920 (N_4920,N_3260,N_3399);
nor U4921 (N_4921,N_3635,N_3522);
or U4922 (N_4922,N_3740,N_3480);
and U4923 (N_4923,N_3827,N_3346);
xor U4924 (N_4924,N_3632,N_3120);
xnor U4925 (N_4925,N_3820,N_3392);
or U4926 (N_4926,N_3187,N_3356);
xnor U4927 (N_4927,N_3212,N_3723);
xnor U4928 (N_4928,N_3775,N_3480);
or U4929 (N_4929,N_3588,N_3695);
and U4930 (N_4930,N_3371,N_3999);
nand U4931 (N_4931,N_3196,N_3668);
or U4932 (N_4932,N_3313,N_3912);
or U4933 (N_4933,N_3789,N_3118);
xnor U4934 (N_4934,N_3923,N_3137);
xnor U4935 (N_4935,N_3506,N_3996);
nand U4936 (N_4936,N_3516,N_3264);
nor U4937 (N_4937,N_3355,N_3561);
nor U4938 (N_4938,N_3532,N_3517);
nand U4939 (N_4939,N_3024,N_3735);
or U4940 (N_4940,N_3413,N_3091);
nand U4941 (N_4941,N_3616,N_3128);
and U4942 (N_4942,N_3487,N_3578);
and U4943 (N_4943,N_3009,N_3371);
xnor U4944 (N_4944,N_3047,N_3655);
or U4945 (N_4945,N_3924,N_3130);
nand U4946 (N_4946,N_3700,N_3099);
or U4947 (N_4947,N_3597,N_3979);
and U4948 (N_4948,N_3232,N_3770);
or U4949 (N_4949,N_3684,N_3152);
nor U4950 (N_4950,N_3853,N_3135);
or U4951 (N_4951,N_3937,N_3057);
xor U4952 (N_4952,N_3802,N_3894);
or U4953 (N_4953,N_3461,N_3844);
and U4954 (N_4954,N_3402,N_3902);
and U4955 (N_4955,N_3805,N_3652);
or U4956 (N_4956,N_3171,N_3801);
nand U4957 (N_4957,N_3697,N_3624);
nor U4958 (N_4958,N_3430,N_3107);
xnor U4959 (N_4959,N_3033,N_3073);
nand U4960 (N_4960,N_3348,N_3356);
xor U4961 (N_4961,N_3757,N_3916);
or U4962 (N_4962,N_3382,N_3017);
xnor U4963 (N_4963,N_3052,N_3184);
nor U4964 (N_4964,N_3833,N_3175);
and U4965 (N_4965,N_3187,N_3958);
or U4966 (N_4966,N_3787,N_3879);
and U4967 (N_4967,N_3052,N_3068);
nand U4968 (N_4968,N_3476,N_3347);
or U4969 (N_4969,N_3089,N_3245);
or U4970 (N_4970,N_3602,N_3526);
nand U4971 (N_4971,N_3790,N_3738);
and U4972 (N_4972,N_3721,N_3169);
and U4973 (N_4973,N_3458,N_3313);
or U4974 (N_4974,N_3562,N_3434);
xnor U4975 (N_4975,N_3892,N_3034);
or U4976 (N_4976,N_3612,N_3656);
nor U4977 (N_4977,N_3161,N_3660);
nand U4978 (N_4978,N_3264,N_3037);
and U4979 (N_4979,N_3186,N_3149);
and U4980 (N_4980,N_3625,N_3146);
or U4981 (N_4981,N_3472,N_3459);
nand U4982 (N_4982,N_3680,N_3334);
nor U4983 (N_4983,N_3652,N_3806);
or U4984 (N_4984,N_3826,N_3997);
nor U4985 (N_4985,N_3654,N_3961);
xnor U4986 (N_4986,N_3602,N_3066);
and U4987 (N_4987,N_3433,N_3205);
or U4988 (N_4988,N_3681,N_3741);
and U4989 (N_4989,N_3744,N_3843);
nand U4990 (N_4990,N_3925,N_3718);
xnor U4991 (N_4991,N_3399,N_3665);
or U4992 (N_4992,N_3869,N_3104);
and U4993 (N_4993,N_3682,N_3926);
xnor U4994 (N_4994,N_3234,N_3851);
and U4995 (N_4995,N_3826,N_3014);
nand U4996 (N_4996,N_3097,N_3250);
and U4997 (N_4997,N_3877,N_3298);
nand U4998 (N_4998,N_3039,N_3811);
nor U4999 (N_4999,N_3527,N_3759);
nor UO_0 (O_0,N_4468,N_4994);
nor UO_1 (O_1,N_4946,N_4127);
xnor UO_2 (O_2,N_4721,N_4858);
nor UO_3 (O_3,N_4520,N_4637);
or UO_4 (O_4,N_4782,N_4112);
xnor UO_5 (O_5,N_4053,N_4656);
and UO_6 (O_6,N_4562,N_4786);
or UO_7 (O_7,N_4934,N_4666);
xnor UO_8 (O_8,N_4716,N_4434);
and UO_9 (O_9,N_4883,N_4373);
or UO_10 (O_10,N_4458,N_4004);
and UO_11 (O_11,N_4330,N_4884);
xnor UO_12 (O_12,N_4660,N_4857);
xor UO_13 (O_13,N_4210,N_4541);
nand UO_14 (O_14,N_4255,N_4751);
or UO_15 (O_15,N_4849,N_4524);
and UO_16 (O_16,N_4226,N_4615);
nand UO_17 (O_17,N_4225,N_4517);
nand UO_18 (O_18,N_4655,N_4794);
and UO_19 (O_19,N_4002,N_4193);
and UO_20 (O_20,N_4907,N_4737);
nor UO_21 (O_21,N_4793,N_4351);
nand UO_22 (O_22,N_4810,N_4558);
nand UO_23 (O_23,N_4145,N_4236);
nor UO_24 (O_24,N_4986,N_4771);
nor UO_25 (O_25,N_4115,N_4902);
nor UO_26 (O_26,N_4270,N_4433);
xnor UO_27 (O_27,N_4046,N_4528);
or UO_28 (O_28,N_4951,N_4886);
nor UO_29 (O_29,N_4108,N_4582);
or UO_30 (O_30,N_4387,N_4937);
nand UO_31 (O_31,N_4231,N_4530);
xnor UO_32 (O_32,N_4215,N_4241);
or UO_33 (O_33,N_4773,N_4739);
nor UO_34 (O_34,N_4459,N_4194);
and UO_35 (O_35,N_4734,N_4341);
xnor UO_36 (O_36,N_4579,N_4779);
nor UO_37 (O_37,N_4221,N_4217);
or UO_38 (O_38,N_4527,N_4532);
nor UO_39 (O_39,N_4589,N_4346);
nand UO_40 (O_40,N_4283,N_4791);
xor UO_41 (O_41,N_4321,N_4631);
nand UO_42 (O_42,N_4186,N_4168);
nand UO_43 (O_43,N_4824,N_4602);
xor UO_44 (O_44,N_4293,N_4109);
nand UO_45 (O_45,N_4161,N_4822);
or UO_46 (O_46,N_4104,N_4788);
nor UO_47 (O_47,N_4795,N_4585);
and UO_48 (O_48,N_4845,N_4633);
nor UO_49 (O_49,N_4727,N_4759);
nor UO_50 (O_50,N_4804,N_4724);
or UO_51 (O_51,N_4000,N_4890);
nand UO_52 (O_52,N_4422,N_4614);
nand UO_53 (O_53,N_4088,N_4314);
xnor UO_54 (O_54,N_4392,N_4407);
nand UO_55 (O_55,N_4509,N_4184);
xor UO_56 (O_56,N_4489,N_4204);
nand UO_57 (O_57,N_4120,N_4682);
or UO_58 (O_58,N_4467,N_4089);
nand UO_59 (O_59,N_4571,N_4006);
nor UO_60 (O_60,N_4889,N_4622);
or UO_61 (O_61,N_4877,N_4757);
or UO_62 (O_62,N_4160,N_4708);
and UO_63 (O_63,N_4235,N_4087);
xor UO_64 (O_64,N_4548,N_4691);
nand UO_65 (O_65,N_4985,N_4769);
and UO_66 (O_66,N_4428,N_4572);
or UO_67 (O_67,N_4008,N_4393);
xor UO_68 (O_68,N_4820,N_4930);
nand UO_69 (O_69,N_4480,N_4383);
nand UO_70 (O_70,N_4277,N_4167);
xor UO_71 (O_71,N_4617,N_4090);
xor UO_72 (O_72,N_4591,N_4342);
or UO_73 (O_73,N_4578,N_4675);
xnor UO_74 (O_74,N_4534,N_4550);
or UO_75 (O_75,N_4110,N_4653);
nand UO_76 (O_76,N_4745,N_4546);
or UO_77 (O_77,N_4254,N_4316);
nand UO_78 (O_78,N_4970,N_4093);
or UO_79 (O_79,N_4418,N_4893);
nand UO_80 (O_80,N_4073,N_4010);
nand UO_81 (O_81,N_4180,N_4685);
or UO_82 (O_82,N_4224,N_4466);
xnor UO_83 (O_83,N_4755,N_4308);
or UO_84 (O_84,N_4230,N_4162);
and UO_85 (O_85,N_4920,N_4057);
nor UO_86 (O_86,N_4706,N_4031);
or UO_87 (O_87,N_4540,N_4928);
and UO_88 (O_88,N_4923,N_4077);
and UO_89 (O_89,N_4697,N_4686);
or UO_90 (O_90,N_4835,N_4095);
and UO_91 (O_91,N_4752,N_4113);
nand UO_92 (O_92,N_4762,N_4324);
or UO_93 (O_93,N_4340,N_4555);
nor UO_94 (O_94,N_4575,N_4134);
nor UO_95 (O_95,N_4438,N_4958);
nor UO_96 (O_96,N_4398,N_4482);
and UO_97 (O_97,N_4083,N_4876);
xor UO_98 (O_98,N_4303,N_4574);
or UO_99 (O_99,N_4016,N_4623);
nor UO_100 (O_100,N_4065,N_4763);
and UO_101 (O_101,N_4538,N_4983);
xor UO_102 (O_102,N_4978,N_4605);
nand UO_103 (O_103,N_4462,N_4137);
and UO_104 (O_104,N_4613,N_4536);
xor UO_105 (O_105,N_4074,N_4882);
or UO_106 (O_106,N_4817,N_4750);
nor UO_107 (O_107,N_4583,N_4245);
nor UO_108 (O_108,N_4408,N_4445);
nand UO_109 (O_109,N_4441,N_4945);
nand UO_110 (O_110,N_4785,N_4586);
nor UO_111 (O_111,N_4363,N_4250);
nor UO_112 (O_112,N_4220,N_4123);
nor UO_113 (O_113,N_4331,N_4329);
and UO_114 (O_114,N_4717,N_4029);
nor UO_115 (O_115,N_4776,N_4045);
and UO_116 (O_116,N_4543,N_4508);
or UO_117 (O_117,N_4625,N_4672);
or UO_118 (O_118,N_4306,N_4126);
nand UO_119 (O_119,N_4023,N_4566);
or UO_120 (O_120,N_4696,N_4499);
or UO_121 (O_121,N_4673,N_4654);
xor UO_122 (O_122,N_4216,N_4298);
and UO_123 (O_123,N_4052,N_4659);
or UO_124 (O_124,N_4081,N_4243);
or UO_125 (O_125,N_4568,N_4909);
or UO_126 (O_126,N_4638,N_4827);
xor UO_127 (O_127,N_4967,N_4015);
or UO_128 (O_128,N_4900,N_4064);
and UO_129 (O_129,N_4311,N_4512);
nand UO_130 (O_130,N_4916,N_4878);
nand UO_131 (O_131,N_4896,N_4189);
or UO_132 (O_132,N_4292,N_4781);
xor UO_133 (O_133,N_4606,N_4357);
nand UO_134 (O_134,N_4834,N_4816);
xor UO_135 (O_135,N_4792,N_4344);
nand UO_136 (O_136,N_4670,N_4136);
nor UO_137 (O_137,N_4478,N_4417);
nand UO_138 (O_138,N_4910,N_4961);
or UO_139 (O_139,N_4688,N_4309);
or UO_140 (O_140,N_4078,N_4118);
xor UO_141 (O_141,N_4378,N_4826);
xnor UO_142 (O_142,N_4263,N_4313);
nor UO_143 (O_143,N_4275,N_4036);
or UO_144 (O_144,N_4103,N_4107);
and UO_145 (O_145,N_4232,N_4304);
nand UO_146 (O_146,N_4477,N_4828);
nand UO_147 (O_147,N_4227,N_4474);
or UO_148 (O_148,N_4476,N_4269);
or UO_149 (O_149,N_4922,N_4479);
nor UO_150 (O_150,N_4367,N_4473);
nand UO_151 (O_151,N_4680,N_4720);
or UO_152 (O_152,N_4328,N_4287);
nand UO_153 (O_153,N_4669,N_4619);
and UO_154 (O_154,N_4425,N_4322);
nor UO_155 (O_155,N_4011,N_4173);
and UO_156 (O_156,N_4833,N_4394);
xor UO_157 (O_157,N_4987,N_4362);
nor UO_158 (O_158,N_4620,N_4405);
or UO_159 (O_159,N_4264,N_4732);
or UO_160 (O_160,N_4544,N_4412);
nand UO_161 (O_161,N_4164,N_4454);
nand UO_162 (O_162,N_4690,N_4609);
nand UO_163 (O_163,N_4183,N_4797);
or UO_164 (O_164,N_4005,N_4860);
nand UO_165 (O_165,N_4977,N_4449);
and UO_166 (O_166,N_4025,N_4139);
nor UO_167 (O_167,N_4808,N_4166);
xnor UO_168 (O_168,N_4192,N_4472);
and UO_169 (O_169,N_4610,N_4068);
nand UO_170 (O_170,N_4359,N_4246);
nand UO_171 (O_171,N_4452,N_4629);
or UO_172 (O_172,N_4514,N_4396);
or UO_173 (O_173,N_4897,N_4502);
or UO_174 (O_174,N_4584,N_4879);
or UO_175 (O_175,N_4526,N_4498);
and UO_176 (O_176,N_4076,N_4624);
and UO_177 (O_177,N_4385,N_4069);
or UO_178 (O_178,N_4554,N_4969);
nor UO_179 (O_179,N_4409,N_4919);
xor UO_180 (O_180,N_4872,N_4741);
or UO_181 (O_181,N_4196,N_4059);
nand UO_182 (O_182,N_4681,N_4847);
or UO_183 (O_183,N_4040,N_4604);
xnor UO_184 (O_184,N_4297,N_4100);
nand UO_185 (O_185,N_4377,N_4097);
nand UO_186 (O_186,N_4353,N_4490);
or UO_187 (O_187,N_4481,N_4033);
xor UO_188 (O_188,N_4956,N_4121);
and UO_189 (O_189,N_4140,N_4778);
xor UO_190 (O_190,N_4101,N_4460);
and UO_191 (O_191,N_4349,N_4042);
and UO_192 (O_192,N_4178,N_4205);
nand UO_193 (O_193,N_4608,N_4705);
or UO_194 (O_194,N_4047,N_4819);
nand UO_195 (O_195,N_4372,N_4749);
nor UO_196 (O_196,N_4163,N_4895);
nor UO_197 (O_197,N_4117,N_4865);
and UO_198 (O_198,N_4701,N_4188);
nand UO_199 (O_199,N_4846,N_4950);
and UO_200 (O_200,N_4948,N_4080);
nor UO_201 (O_201,N_4809,N_4147);
nor UO_202 (O_202,N_4823,N_4856);
or UO_203 (O_203,N_4627,N_4171);
and UO_204 (O_204,N_4281,N_4726);
nand UO_205 (O_205,N_4746,N_4679);
nor UO_206 (O_206,N_4198,N_4249);
or UO_207 (O_207,N_4256,N_4949);
or UO_208 (O_208,N_4326,N_4212);
and UO_209 (O_209,N_4818,N_4457);
and UO_210 (O_210,N_4354,N_4237);
nand UO_211 (O_211,N_4487,N_4632);
nor UO_212 (O_212,N_4772,N_4401);
and UO_213 (O_213,N_4430,N_4567);
xnor UO_214 (O_214,N_4844,N_4259);
nand UO_215 (O_215,N_4456,N_4796);
and UO_216 (O_216,N_4291,N_4975);
and UO_217 (O_217,N_4825,N_4646);
and UO_218 (O_218,N_4429,N_4239);
nand UO_219 (O_219,N_4894,N_4932);
or UO_220 (O_220,N_4661,N_4348);
nor UO_221 (O_221,N_4455,N_4470);
nand UO_222 (O_222,N_4390,N_4347);
or UO_223 (O_223,N_4503,N_4335);
or UO_224 (O_224,N_4174,N_4537);
or UO_225 (O_225,N_4634,N_4294);
nand UO_226 (O_226,N_4742,N_4169);
nand UO_227 (O_227,N_4507,N_4038);
nor UO_228 (O_228,N_4301,N_4272);
and UO_229 (O_229,N_4652,N_4024);
xnor UO_230 (O_230,N_4130,N_4596);
xor UO_231 (O_231,N_4391,N_4247);
and UO_232 (O_232,N_4838,N_4873);
xor UO_233 (O_233,N_4406,N_4523);
nor UO_234 (O_234,N_4784,N_4616);
and UO_235 (O_235,N_4182,N_4718);
and UO_236 (O_236,N_4668,N_4547);
or UO_237 (O_237,N_4626,N_4775);
nand UO_238 (O_238,N_4840,N_4731);
xnor UO_239 (O_239,N_4411,N_4658);
nand UO_240 (O_240,N_4601,N_4404);
and UO_241 (O_241,N_4060,N_4942);
nand UO_242 (O_242,N_4159,N_4501);
nand UO_243 (O_243,N_4802,N_4268);
xor UO_244 (O_244,N_4261,N_4091);
xor UO_245 (O_245,N_4560,N_4175);
or UO_246 (O_246,N_4343,N_4267);
or UO_247 (O_247,N_4027,N_4993);
or UO_248 (O_248,N_4018,N_4891);
nor UO_249 (O_249,N_4648,N_4929);
nor UO_250 (O_250,N_4233,N_4228);
nand UO_251 (O_251,N_4310,N_4594);
and UO_252 (O_252,N_4244,N_4995);
and UO_253 (O_253,N_4397,N_4754);
nor UO_254 (O_254,N_4248,N_4687);
nand UO_255 (O_255,N_4419,N_4282);
nor UO_256 (O_256,N_4735,N_4700);
nor UO_257 (O_257,N_4049,N_4003);
or UO_258 (O_258,N_4063,N_4376);
xnor UO_259 (O_259,N_4102,N_4465);
nor UO_260 (O_260,N_4729,N_4370);
nor UO_261 (O_261,N_4753,N_4111);
and UO_262 (O_262,N_4152,N_4054);
xor UO_263 (O_263,N_4092,N_4319);
nor UO_264 (O_264,N_4592,N_4009);
xor UO_265 (O_265,N_4260,N_4832);
nor UO_266 (O_266,N_4071,N_4984);
or UO_267 (O_267,N_4400,N_4384);
nor UO_268 (O_268,N_4369,N_4657);
and UO_269 (O_269,N_4851,N_4019);
or UO_270 (O_270,N_4761,N_4667);
or UO_271 (O_271,N_4713,N_4295);
or UO_272 (O_272,N_4611,N_4278);
or UO_273 (O_273,N_4442,N_4725);
or UO_274 (O_274,N_4436,N_4446);
xnor UO_275 (O_275,N_4997,N_4960);
or UO_276 (O_276,N_4553,N_4240);
or UO_277 (O_277,N_4711,N_4318);
nand UO_278 (O_278,N_4219,N_4143);
or UO_279 (O_279,N_4056,N_4258);
nor UO_280 (O_280,N_4395,N_4728);
xnor UO_281 (O_281,N_4787,N_4551);
or UO_282 (O_282,N_4981,N_4513);
and UO_283 (O_283,N_4381,N_4830);
nand UO_284 (O_284,N_4821,N_4229);
nor UO_285 (O_285,N_4689,N_4423);
nand UO_286 (O_286,N_4525,N_4158);
nor UO_287 (O_287,N_4133,N_4875);
xnor UO_288 (O_288,N_4743,N_4148);
xnor UO_289 (O_289,N_4307,N_4765);
or UO_290 (O_290,N_4564,N_4070);
or UO_291 (O_291,N_4050,N_4190);
nand UO_292 (O_292,N_4976,N_4955);
xor UO_293 (O_293,N_4800,N_4837);
nand UO_294 (O_294,N_4201,N_4427);
xor UO_295 (O_295,N_4518,N_4420);
nand UO_296 (O_296,N_4736,N_4815);
nand UO_297 (O_297,N_4814,N_4475);
or UO_298 (O_298,N_4842,N_4124);
xnor UO_299 (O_299,N_4360,N_4813);
xnor UO_300 (O_300,N_4157,N_4590);
nor UO_301 (O_301,N_4315,N_4209);
nand UO_302 (O_302,N_4099,N_4971);
nor UO_303 (O_303,N_4181,N_4086);
nand UO_304 (O_304,N_4251,N_4125);
nand UO_305 (O_305,N_4048,N_4388);
nand UO_306 (O_306,N_4563,N_4663);
and UO_307 (O_307,N_4106,N_4870);
and UO_308 (O_308,N_4402,N_4361);
xnor UO_309 (O_309,N_4222,N_4767);
or UO_310 (O_310,N_4698,N_4988);
or UO_311 (O_311,N_4020,N_4839);
nand UO_312 (O_312,N_4829,N_4364);
xnor UO_313 (O_313,N_4549,N_4756);
xnor UO_314 (O_314,N_4154,N_4723);
or UO_315 (O_315,N_4671,N_4651);
nor UO_316 (O_316,N_4580,N_4067);
nand UO_317 (O_317,N_4177,N_4707);
nor UO_318 (O_318,N_4510,N_4991);
or UO_319 (O_319,N_4569,N_4545);
nor UO_320 (O_320,N_4841,N_4208);
nand UO_321 (O_321,N_4676,N_4296);
nand UO_322 (O_322,N_4386,N_4940);
nor UO_323 (O_323,N_4075,N_4740);
or UO_324 (O_324,N_4336,N_4305);
or UO_325 (O_325,N_4271,N_4904);
nor UO_326 (O_326,N_4603,N_4098);
and UO_327 (O_327,N_4665,N_4947);
xor UO_328 (O_328,N_4760,N_4021);
and UO_329 (O_329,N_4338,N_4368);
xnor UO_330 (O_330,N_4051,N_4055);
and UO_331 (O_331,N_4966,N_4469);
nor UO_332 (O_332,N_4887,N_4062);
and UO_333 (O_333,N_4079,N_4935);
nand UO_334 (O_334,N_4790,N_4030);
nand UO_335 (O_335,N_4963,N_4630);
or UO_336 (O_336,N_4013,N_4848);
nand UO_337 (O_337,N_4733,N_4214);
nor UO_338 (O_338,N_4085,N_4415);
and UO_339 (O_339,N_4612,N_4366);
and UO_340 (O_340,N_4265,N_4200);
xnor UO_341 (O_341,N_4043,N_4375);
and UO_342 (O_342,N_4628,N_4964);
nand UO_343 (O_343,N_4252,N_4938);
xor UO_344 (O_344,N_4519,N_4035);
nor UO_345 (O_345,N_4153,N_4202);
xnor UO_346 (O_346,N_4486,N_4443);
xnor UO_347 (O_347,N_4931,N_4905);
nand UO_348 (O_348,N_4061,N_4593);
nand UO_349 (O_349,N_4327,N_4644);
and UO_350 (O_350,N_4521,N_4421);
or UO_351 (O_351,N_4149,N_4650);
and UO_352 (O_352,N_4165,N_4693);
and UO_353 (O_353,N_4012,N_4439);
xor UO_354 (O_354,N_4323,N_4768);
nor UO_355 (O_355,N_4965,N_4597);
and UO_356 (O_356,N_4389,N_4944);
or UO_357 (O_357,N_4803,N_4289);
nand UO_358 (O_358,N_4722,N_4766);
and UO_359 (O_359,N_4285,N_4866);
and UO_360 (O_360,N_4119,N_4719);
or UO_361 (O_361,N_4500,N_4494);
xnor UO_362 (O_362,N_4730,N_4641);
and UO_363 (O_363,N_4587,N_4511);
or UO_364 (O_364,N_4712,N_4999);
or UO_365 (O_365,N_4864,N_4424);
and UO_366 (O_366,N_4274,N_4709);
or UO_367 (O_367,N_4643,N_4504);
nand UO_368 (O_368,N_4094,N_4176);
xnor UO_369 (O_369,N_4913,N_4379);
or UO_370 (O_370,N_4276,N_4533);
nor UO_371 (O_371,N_4715,N_4156);
and UO_372 (O_372,N_4356,N_4704);
and UO_373 (O_373,N_4032,N_4885);
nand UO_374 (O_374,N_4414,N_4805);
or UO_375 (O_375,N_4855,N_4598);
xor UO_376 (O_376,N_4852,N_4968);
or UO_377 (O_377,N_4144,N_4618);
nand UO_378 (O_378,N_4992,N_4461);
and UO_379 (O_379,N_4952,N_4432);
and UO_380 (O_380,N_4874,N_4565);
xor UO_381 (O_381,N_4863,N_4780);
xor UO_382 (O_382,N_4440,N_4072);
and UO_383 (O_383,N_4413,N_4451);
nor UO_384 (O_384,N_4677,N_4801);
nand UO_385 (O_385,N_4898,N_4556);
xnor UO_386 (O_386,N_4843,N_4096);
nand UO_387 (O_387,N_4744,N_4382);
or UO_388 (O_388,N_4933,N_4869);
and UO_389 (O_389,N_4223,N_4234);
or UO_390 (O_390,N_4426,N_4774);
nor UO_391 (O_391,N_4539,N_4084);
nor UO_392 (O_392,N_4279,N_4924);
xnor UO_393 (O_393,N_4355,N_4962);
xnor UO_394 (O_394,N_4497,N_4645);
xnor UO_395 (O_395,N_4542,N_4374);
nor UO_396 (O_396,N_4901,N_4288);
nor UO_397 (O_397,N_4936,N_4170);
xnor UO_398 (O_398,N_4570,N_4664);
and UO_399 (O_399,N_4197,N_4974);
or UO_400 (O_400,N_4262,N_4853);
nor UO_401 (O_401,N_4918,N_4317);
or UO_402 (O_402,N_4129,N_4989);
nand UO_403 (O_403,N_4151,N_4703);
nor UO_404 (O_404,N_4485,N_4595);
nand UO_405 (O_405,N_4320,N_4471);
xnor UO_406 (O_406,N_4635,N_4806);
nor UO_407 (O_407,N_4284,N_4710);
xnor UO_408 (O_408,N_4001,N_4135);
and UO_409 (O_409,N_4927,N_4082);
and UO_410 (O_410,N_4831,N_4191);
xnor UO_411 (O_411,N_4990,N_4561);
nand UO_412 (O_412,N_4812,N_4581);
or UO_413 (O_413,N_4639,N_4531);
nor UO_414 (O_414,N_4522,N_4345);
nor UO_415 (O_415,N_4647,N_4506);
xnor UO_416 (O_416,N_4954,N_4973);
and UO_417 (O_417,N_4516,N_4577);
or UO_418 (O_418,N_4380,N_4939);
xnor UO_419 (O_419,N_4290,N_4600);
or UO_420 (O_420,N_4892,N_4777);
and UO_421 (O_421,N_4836,N_4535);
xnor UO_422 (O_422,N_4496,N_4266);
or UO_423 (O_423,N_4943,N_4207);
and UO_424 (O_424,N_4206,N_4914);
and UO_425 (O_425,N_4491,N_4435);
nand UO_426 (O_426,N_4017,N_4037);
nor UO_427 (O_427,N_4495,N_4621);
xor UO_428 (O_428,N_4333,N_4399);
xor UO_429 (O_429,N_4058,N_4488);
xnor UO_430 (O_430,N_4702,N_4861);
or UO_431 (O_431,N_4447,N_4312);
xor UO_432 (O_432,N_4453,N_4437);
and UO_433 (O_433,N_4748,N_4041);
nand UO_434 (O_434,N_4915,N_4242);
nand UO_435 (O_435,N_4280,N_4926);
or UO_436 (O_436,N_4195,N_4908);
nand UO_437 (O_437,N_4747,N_4862);
xor UO_438 (O_438,N_4557,N_4695);
nor UO_439 (O_439,N_4483,N_4529);
xnor UO_440 (O_440,N_4416,N_4448);
xor UO_441 (O_441,N_4906,N_4683);
xnor UO_442 (O_442,N_4694,N_4871);
nand UO_443 (O_443,N_4559,N_4492);
nand UO_444 (O_444,N_4917,N_4789);
and UO_445 (O_445,N_4132,N_4141);
nor UO_446 (O_446,N_4758,N_4146);
nor UO_447 (O_447,N_4150,N_4187);
nand UO_448 (O_448,N_4179,N_4128);
and UO_449 (O_449,N_4365,N_4684);
or UO_450 (O_450,N_4925,N_4979);
xnor UO_451 (O_451,N_4505,N_4122);
xnor UO_452 (O_452,N_4142,N_4185);
nand UO_453 (O_453,N_4642,N_4764);
and UO_454 (O_454,N_4213,N_4921);
or UO_455 (O_455,N_4980,N_4854);
nand UO_456 (O_456,N_4028,N_4325);
or UO_457 (O_457,N_4941,N_4996);
or UO_458 (O_458,N_4273,N_4337);
nand UO_459 (O_459,N_4014,N_4982);
nor UO_460 (O_460,N_4807,N_4463);
or UO_461 (O_461,N_4850,N_4493);
and UO_462 (O_462,N_4131,N_4403);
or UO_463 (O_463,N_4211,N_4350);
nand UO_464 (O_464,N_4026,N_4116);
or UO_465 (O_465,N_4299,N_4957);
nor UO_466 (O_466,N_4770,N_4998);
and UO_467 (O_467,N_4352,N_4674);
and UO_468 (O_468,N_4253,N_4172);
or UO_469 (O_469,N_4798,N_4450);
nand UO_470 (O_470,N_4155,N_4588);
or UO_471 (O_471,N_4953,N_4358);
and UO_472 (O_472,N_4662,N_4007);
and UO_473 (O_473,N_4431,N_4332);
nor UO_474 (O_474,N_4114,N_4903);
or UO_475 (O_475,N_4783,N_4039);
nand UO_476 (O_476,N_4034,N_4859);
nand UO_477 (O_477,N_4912,N_4302);
nand UO_478 (O_478,N_4607,N_4484);
nor UO_479 (O_479,N_4199,N_4334);
nor UO_480 (O_480,N_4714,N_4880);
nor UO_481 (O_481,N_4599,N_4138);
and UO_482 (O_482,N_4203,N_4699);
xor UO_483 (O_483,N_4218,N_4105);
nor UO_484 (O_484,N_4576,N_4286);
or UO_485 (O_485,N_4888,N_4300);
nor UO_486 (O_486,N_4868,N_4238);
and UO_487 (O_487,N_4410,N_4044);
or UO_488 (O_488,N_4899,N_4738);
and UO_489 (O_489,N_4881,N_4692);
nand UO_490 (O_490,N_4649,N_4972);
and UO_491 (O_491,N_4799,N_4959);
nor UO_492 (O_492,N_4911,N_4867);
and UO_493 (O_493,N_4552,N_4464);
and UO_494 (O_494,N_4444,N_4636);
nor UO_495 (O_495,N_4515,N_4257);
and UO_496 (O_496,N_4339,N_4640);
or UO_497 (O_497,N_4371,N_4066);
xnor UO_498 (O_498,N_4678,N_4573);
xor UO_499 (O_499,N_4811,N_4022);
nor UO_500 (O_500,N_4720,N_4047);
xnor UO_501 (O_501,N_4601,N_4035);
nor UO_502 (O_502,N_4312,N_4992);
nor UO_503 (O_503,N_4458,N_4329);
xor UO_504 (O_504,N_4656,N_4830);
nor UO_505 (O_505,N_4448,N_4305);
nor UO_506 (O_506,N_4620,N_4747);
nor UO_507 (O_507,N_4031,N_4907);
or UO_508 (O_508,N_4481,N_4149);
nor UO_509 (O_509,N_4369,N_4932);
xnor UO_510 (O_510,N_4012,N_4868);
nand UO_511 (O_511,N_4161,N_4453);
or UO_512 (O_512,N_4619,N_4341);
nand UO_513 (O_513,N_4388,N_4884);
and UO_514 (O_514,N_4865,N_4686);
nor UO_515 (O_515,N_4951,N_4436);
nor UO_516 (O_516,N_4913,N_4508);
and UO_517 (O_517,N_4628,N_4249);
nor UO_518 (O_518,N_4276,N_4971);
or UO_519 (O_519,N_4301,N_4653);
xor UO_520 (O_520,N_4540,N_4404);
xor UO_521 (O_521,N_4925,N_4488);
nand UO_522 (O_522,N_4386,N_4928);
xor UO_523 (O_523,N_4526,N_4014);
nand UO_524 (O_524,N_4045,N_4423);
or UO_525 (O_525,N_4069,N_4457);
nand UO_526 (O_526,N_4804,N_4575);
xnor UO_527 (O_527,N_4899,N_4911);
or UO_528 (O_528,N_4023,N_4306);
and UO_529 (O_529,N_4654,N_4442);
xor UO_530 (O_530,N_4780,N_4442);
and UO_531 (O_531,N_4615,N_4174);
and UO_532 (O_532,N_4460,N_4275);
and UO_533 (O_533,N_4757,N_4357);
xor UO_534 (O_534,N_4602,N_4508);
nand UO_535 (O_535,N_4218,N_4718);
nand UO_536 (O_536,N_4067,N_4599);
nand UO_537 (O_537,N_4851,N_4621);
or UO_538 (O_538,N_4387,N_4201);
nand UO_539 (O_539,N_4734,N_4900);
nand UO_540 (O_540,N_4456,N_4339);
or UO_541 (O_541,N_4705,N_4765);
xor UO_542 (O_542,N_4136,N_4490);
xnor UO_543 (O_543,N_4385,N_4559);
nor UO_544 (O_544,N_4983,N_4455);
xnor UO_545 (O_545,N_4973,N_4914);
nand UO_546 (O_546,N_4902,N_4516);
or UO_547 (O_547,N_4520,N_4558);
nor UO_548 (O_548,N_4059,N_4327);
or UO_549 (O_549,N_4459,N_4001);
or UO_550 (O_550,N_4083,N_4920);
nand UO_551 (O_551,N_4071,N_4804);
nor UO_552 (O_552,N_4470,N_4229);
and UO_553 (O_553,N_4891,N_4612);
xnor UO_554 (O_554,N_4098,N_4362);
nand UO_555 (O_555,N_4780,N_4891);
nand UO_556 (O_556,N_4381,N_4239);
xnor UO_557 (O_557,N_4067,N_4405);
or UO_558 (O_558,N_4672,N_4620);
nor UO_559 (O_559,N_4339,N_4537);
xnor UO_560 (O_560,N_4269,N_4123);
nand UO_561 (O_561,N_4806,N_4147);
or UO_562 (O_562,N_4737,N_4720);
and UO_563 (O_563,N_4425,N_4206);
xor UO_564 (O_564,N_4520,N_4173);
nor UO_565 (O_565,N_4805,N_4144);
nor UO_566 (O_566,N_4160,N_4375);
or UO_567 (O_567,N_4879,N_4551);
xnor UO_568 (O_568,N_4133,N_4048);
and UO_569 (O_569,N_4813,N_4178);
nand UO_570 (O_570,N_4408,N_4090);
nand UO_571 (O_571,N_4171,N_4487);
and UO_572 (O_572,N_4884,N_4806);
nor UO_573 (O_573,N_4191,N_4766);
xnor UO_574 (O_574,N_4370,N_4731);
nand UO_575 (O_575,N_4071,N_4321);
xnor UO_576 (O_576,N_4224,N_4336);
and UO_577 (O_577,N_4322,N_4932);
nor UO_578 (O_578,N_4774,N_4379);
xnor UO_579 (O_579,N_4709,N_4190);
nand UO_580 (O_580,N_4325,N_4681);
xnor UO_581 (O_581,N_4472,N_4381);
nand UO_582 (O_582,N_4131,N_4554);
nand UO_583 (O_583,N_4449,N_4893);
xnor UO_584 (O_584,N_4284,N_4779);
xor UO_585 (O_585,N_4725,N_4396);
xnor UO_586 (O_586,N_4849,N_4252);
xor UO_587 (O_587,N_4207,N_4663);
or UO_588 (O_588,N_4385,N_4245);
or UO_589 (O_589,N_4022,N_4092);
nand UO_590 (O_590,N_4934,N_4158);
xor UO_591 (O_591,N_4547,N_4054);
nor UO_592 (O_592,N_4738,N_4263);
nor UO_593 (O_593,N_4885,N_4110);
xnor UO_594 (O_594,N_4628,N_4659);
nand UO_595 (O_595,N_4032,N_4739);
nor UO_596 (O_596,N_4127,N_4506);
and UO_597 (O_597,N_4674,N_4140);
nor UO_598 (O_598,N_4908,N_4435);
or UO_599 (O_599,N_4915,N_4481);
nor UO_600 (O_600,N_4108,N_4325);
nand UO_601 (O_601,N_4348,N_4124);
nor UO_602 (O_602,N_4222,N_4699);
xor UO_603 (O_603,N_4846,N_4788);
or UO_604 (O_604,N_4606,N_4983);
nand UO_605 (O_605,N_4523,N_4826);
xor UO_606 (O_606,N_4155,N_4403);
or UO_607 (O_607,N_4366,N_4178);
nor UO_608 (O_608,N_4567,N_4113);
and UO_609 (O_609,N_4660,N_4042);
and UO_610 (O_610,N_4668,N_4427);
or UO_611 (O_611,N_4535,N_4555);
nor UO_612 (O_612,N_4754,N_4011);
or UO_613 (O_613,N_4628,N_4965);
nor UO_614 (O_614,N_4432,N_4487);
nor UO_615 (O_615,N_4198,N_4030);
nand UO_616 (O_616,N_4102,N_4171);
xor UO_617 (O_617,N_4694,N_4361);
nand UO_618 (O_618,N_4970,N_4295);
nor UO_619 (O_619,N_4065,N_4517);
and UO_620 (O_620,N_4475,N_4139);
nand UO_621 (O_621,N_4445,N_4688);
and UO_622 (O_622,N_4134,N_4785);
nor UO_623 (O_623,N_4438,N_4466);
nor UO_624 (O_624,N_4856,N_4415);
or UO_625 (O_625,N_4950,N_4983);
and UO_626 (O_626,N_4838,N_4001);
and UO_627 (O_627,N_4146,N_4294);
or UO_628 (O_628,N_4424,N_4800);
nor UO_629 (O_629,N_4142,N_4593);
nand UO_630 (O_630,N_4379,N_4184);
xnor UO_631 (O_631,N_4874,N_4140);
or UO_632 (O_632,N_4609,N_4257);
nor UO_633 (O_633,N_4947,N_4574);
xor UO_634 (O_634,N_4748,N_4929);
or UO_635 (O_635,N_4645,N_4079);
or UO_636 (O_636,N_4014,N_4742);
nand UO_637 (O_637,N_4480,N_4677);
and UO_638 (O_638,N_4349,N_4363);
xnor UO_639 (O_639,N_4259,N_4794);
nor UO_640 (O_640,N_4061,N_4788);
xnor UO_641 (O_641,N_4445,N_4501);
and UO_642 (O_642,N_4478,N_4466);
nand UO_643 (O_643,N_4868,N_4515);
and UO_644 (O_644,N_4235,N_4908);
nor UO_645 (O_645,N_4280,N_4144);
or UO_646 (O_646,N_4580,N_4272);
nor UO_647 (O_647,N_4123,N_4547);
nand UO_648 (O_648,N_4611,N_4571);
nand UO_649 (O_649,N_4601,N_4527);
or UO_650 (O_650,N_4435,N_4838);
or UO_651 (O_651,N_4353,N_4731);
nor UO_652 (O_652,N_4058,N_4062);
or UO_653 (O_653,N_4449,N_4731);
xnor UO_654 (O_654,N_4985,N_4953);
xnor UO_655 (O_655,N_4415,N_4145);
and UO_656 (O_656,N_4474,N_4953);
xnor UO_657 (O_657,N_4497,N_4756);
nor UO_658 (O_658,N_4942,N_4499);
nor UO_659 (O_659,N_4391,N_4166);
nor UO_660 (O_660,N_4785,N_4827);
or UO_661 (O_661,N_4363,N_4671);
and UO_662 (O_662,N_4210,N_4859);
and UO_663 (O_663,N_4956,N_4909);
and UO_664 (O_664,N_4154,N_4236);
nand UO_665 (O_665,N_4097,N_4597);
xnor UO_666 (O_666,N_4768,N_4800);
nor UO_667 (O_667,N_4947,N_4886);
xor UO_668 (O_668,N_4858,N_4506);
and UO_669 (O_669,N_4831,N_4668);
xnor UO_670 (O_670,N_4648,N_4669);
xnor UO_671 (O_671,N_4172,N_4890);
xnor UO_672 (O_672,N_4306,N_4450);
nand UO_673 (O_673,N_4410,N_4009);
nor UO_674 (O_674,N_4073,N_4857);
nand UO_675 (O_675,N_4590,N_4623);
nand UO_676 (O_676,N_4889,N_4758);
xnor UO_677 (O_677,N_4432,N_4190);
nand UO_678 (O_678,N_4256,N_4986);
and UO_679 (O_679,N_4386,N_4028);
nor UO_680 (O_680,N_4463,N_4041);
nand UO_681 (O_681,N_4221,N_4307);
or UO_682 (O_682,N_4479,N_4874);
and UO_683 (O_683,N_4819,N_4592);
nor UO_684 (O_684,N_4204,N_4856);
nor UO_685 (O_685,N_4070,N_4686);
nand UO_686 (O_686,N_4719,N_4836);
nor UO_687 (O_687,N_4598,N_4249);
nor UO_688 (O_688,N_4599,N_4400);
or UO_689 (O_689,N_4197,N_4932);
nor UO_690 (O_690,N_4668,N_4082);
and UO_691 (O_691,N_4496,N_4302);
xor UO_692 (O_692,N_4686,N_4104);
nor UO_693 (O_693,N_4417,N_4930);
or UO_694 (O_694,N_4173,N_4616);
nand UO_695 (O_695,N_4149,N_4795);
xnor UO_696 (O_696,N_4939,N_4606);
xor UO_697 (O_697,N_4790,N_4219);
and UO_698 (O_698,N_4075,N_4450);
and UO_699 (O_699,N_4993,N_4519);
or UO_700 (O_700,N_4557,N_4755);
or UO_701 (O_701,N_4527,N_4739);
nor UO_702 (O_702,N_4951,N_4700);
or UO_703 (O_703,N_4498,N_4004);
nor UO_704 (O_704,N_4922,N_4249);
nor UO_705 (O_705,N_4743,N_4210);
nor UO_706 (O_706,N_4518,N_4949);
nor UO_707 (O_707,N_4736,N_4544);
nand UO_708 (O_708,N_4534,N_4646);
nand UO_709 (O_709,N_4118,N_4349);
xor UO_710 (O_710,N_4258,N_4646);
nand UO_711 (O_711,N_4902,N_4882);
or UO_712 (O_712,N_4592,N_4642);
or UO_713 (O_713,N_4084,N_4732);
nand UO_714 (O_714,N_4816,N_4450);
and UO_715 (O_715,N_4681,N_4144);
nor UO_716 (O_716,N_4549,N_4002);
nand UO_717 (O_717,N_4883,N_4705);
xor UO_718 (O_718,N_4058,N_4797);
xnor UO_719 (O_719,N_4137,N_4750);
nand UO_720 (O_720,N_4799,N_4653);
or UO_721 (O_721,N_4746,N_4875);
nand UO_722 (O_722,N_4068,N_4520);
nor UO_723 (O_723,N_4098,N_4423);
nand UO_724 (O_724,N_4186,N_4314);
nand UO_725 (O_725,N_4387,N_4944);
nand UO_726 (O_726,N_4415,N_4602);
or UO_727 (O_727,N_4357,N_4981);
and UO_728 (O_728,N_4559,N_4591);
nor UO_729 (O_729,N_4730,N_4025);
or UO_730 (O_730,N_4313,N_4445);
nand UO_731 (O_731,N_4036,N_4545);
xnor UO_732 (O_732,N_4338,N_4513);
or UO_733 (O_733,N_4664,N_4393);
or UO_734 (O_734,N_4086,N_4226);
nor UO_735 (O_735,N_4678,N_4557);
xnor UO_736 (O_736,N_4450,N_4722);
or UO_737 (O_737,N_4269,N_4467);
xnor UO_738 (O_738,N_4593,N_4826);
xnor UO_739 (O_739,N_4409,N_4942);
or UO_740 (O_740,N_4333,N_4997);
nor UO_741 (O_741,N_4179,N_4039);
or UO_742 (O_742,N_4299,N_4142);
nand UO_743 (O_743,N_4986,N_4961);
or UO_744 (O_744,N_4815,N_4532);
nor UO_745 (O_745,N_4723,N_4271);
and UO_746 (O_746,N_4958,N_4960);
nor UO_747 (O_747,N_4609,N_4323);
or UO_748 (O_748,N_4368,N_4790);
nor UO_749 (O_749,N_4443,N_4615);
nand UO_750 (O_750,N_4288,N_4132);
or UO_751 (O_751,N_4578,N_4829);
nand UO_752 (O_752,N_4814,N_4457);
and UO_753 (O_753,N_4318,N_4896);
and UO_754 (O_754,N_4094,N_4603);
nand UO_755 (O_755,N_4882,N_4482);
xor UO_756 (O_756,N_4170,N_4310);
nor UO_757 (O_757,N_4780,N_4737);
xnor UO_758 (O_758,N_4853,N_4361);
nor UO_759 (O_759,N_4104,N_4229);
nand UO_760 (O_760,N_4449,N_4856);
nor UO_761 (O_761,N_4283,N_4332);
nor UO_762 (O_762,N_4597,N_4301);
and UO_763 (O_763,N_4457,N_4119);
nand UO_764 (O_764,N_4627,N_4546);
nor UO_765 (O_765,N_4307,N_4849);
nor UO_766 (O_766,N_4170,N_4197);
nor UO_767 (O_767,N_4117,N_4521);
or UO_768 (O_768,N_4509,N_4188);
nor UO_769 (O_769,N_4129,N_4854);
nor UO_770 (O_770,N_4170,N_4109);
xnor UO_771 (O_771,N_4509,N_4318);
and UO_772 (O_772,N_4458,N_4163);
nor UO_773 (O_773,N_4807,N_4279);
xor UO_774 (O_774,N_4021,N_4835);
nand UO_775 (O_775,N_4983,N_4563);
nand UO_776 (O_776,N_4558,N_4902);
or UO_777 (O_777,N_4116,N_4376);
and UO_778 (O_778,N_4319,N_4057);
nor UO_779 (O_779,N_4601,N_4492);
xor UO_780 (O_780,N_4856,N_4288);
nand UO_781 (O_781,N_4883,N_4346);
nor UO_782 (O_782,N_4507,N_4725);
and UO_783 (O_783,N_4309,N_4882);
nand UO_784 (O_784,N_4741,N_4928);
or UO_785 (O_785,N_4793,N_4389);
and UO_786 (O_786,N_4004,N_4059);
xnor UO_787 (O_787,N_4868,N_4231);
or UO_788 (O_788,N_4702,N_4735);
or UO_789 (O_789,N_4871,N_4927);
or UO_790 (O_790,N_4989,N_4136);
nand UO_791 (O_791,N_4552,N_4781);
nand UO_792 (O_792,N_4617,N_4728);
and UO_793 (O_793,N_4419,N_4802);
and UO_794 (O_794,N_4910,N_4276);
nand UO_795 (O_795,N_4643,N_4136);
xor UO_796 (O_796,N_4454,N_4101);
xor UO_797 (O_797,N_4751,N_4714);
and UO_798 (O_798,N_4489,N_4701);
or UO_799 (O_799,N_4925,N_4077);
and UO_800 (O_800,N_4404,N_4788);
nor UO_801 (O_801,N_4240,N_4647);
and UO_802 (O_802,N_4418,N_4453);
and UO_803 (O_803,N_4821,N_4147);
nand UO_804 (O_804,N_4916,N_4029);
or UO_805 (O_805,N_4781,N_4709);
xnor UO_806 (O_806,N_4193,N_4442);
or UO_807 (O_807,N_4610,N_4139);
nand UO_808 (O_808,N_4525,N_4560);
nor UO_809 (O_809,N_4356,N_4709);
xor UO_810 (O_810,N_4403,N_4803);
nand UO_811 (O_811,N_4057,N_4451);
or UO_812 (O_812,N_4801,N_4735);
nand UO_813 (O_813,N_4975,N_4674);
and UO_814 (O_814,N_4214,N_4728);
xor UO_815 (O_815,N_4841,N_4903);
nor UO_816 (O_816,N_4632,N_4688);
nand UO_817 (O_817,N_4666,N_4055);
or UO_818 (O_818,N_4390,N_4664);
and UO_819 (O_819,N_4928,N_4621);
nor UO_820 (O_820,N_4258,N_4701);
or UO_821 (O_821,N_4101,N_4964);
nor UO_822 (O_822,N_4148,N_4388);
xnor UO_823 (O_823,N_4940,N_4624);
and UO_824 (O_824,N_4676,N_4986);
xor UO_825 (O_825,N_4107,N_4327);
nor UO_826 (O_826,N_4178,N_4588);
nand UO_827 (O_827,N_4119,N_4985);
and UO_828 (O_828,N_4624,N_4771);
nand UO_829 (O_829,N_4279,N_4249);
nor UO_830 (O_830,N_4853,N_4763);
nand UO_831 (O_831,N_4996,N_4852);
nand UO_832 (O_832,N_4949,N_4806);
or UO_833 (O_833,N_4578,N_4055);
nor UO_834 (O_834,N_4935,N_4134);
nor UO_835 (O_835,N_4062,N_4286);
or UO_836 (O_836,N_4235,N_4144);
or UO_837 (O_837,N_4843,N_4040);
xor UO_838 (O_838,N_4651,N_4303);
and UO_839 (O_839,N_4330,N_4027);
nor UO_840 (O_840,N_4785,N_4852);
nor UO_841 (O_841,N_4202,N_4259);
nor UO_842 (O_842,N_4167,N_4166);
or UO_843 (O_843,N_4793,N_4155);
and UO_844 (O_844,N_4132,N_4343);
nor UO_845 (O_845,N_4322,N_4009);
or UO_846 (O_846,N_4235,N_4152);
nand UO_847 (O_847,N_4909,N_4418);
nand UO_848 (O_848,N_4057,N_4188);
nor UO_849 (O_849,N_4654,N_4134);
or UO_850 (O_850,N_4569,N_4381);
xor UO_851 (O_851,N_4359,N_4978);
nand UO_852 (O_852,N_4292,N_4328);
nand UO_853 (O_853,N_4634,N_4824);
or UO_854 (O_854,N_4478,N_4957);
nand UO_855 (O_855,N_4074,N_4821);
nand UO_856 (O_856,N_4412,N_4828);
or UO_857 (O_857,N_4837,N_4730);
xnor UO_858 (O_858,N_4598,N_4668);
nor UO_859 (O_859,N_4015,N_4636);
or UO_860 (O_860,N_4964,N_4043);
and UO_861 (O_861,N_4880,N_4976);
and UO_862 (O_862,N_4048,N_4573);
nand UO_863 (O_863,N_4519,N_4754);
nor UO_864 (O_864,N_4939,N_4836);
xnor UO_865 (O_865,N_4129,N_4446);
xnor UO_866 (O_866,N_4856,N_4594);
or UO_867 (O_867,N_4260,N_4451);
nand UO_868 (O_868,N_4946,N_4596);
and UO_869 (O_869,N_4646,N_4688);
and UO_870 (O_870,N_4520,N_4149);
and UO_871 (O_871,N_4142,N_4648);
or UO_872 (O_872,N_4548,N_4728);
or UO_873 (O_873,N_4292,N_4440);
xor UO_874 (O_874,N_4399,N_4443);
nand UO_875 (O_875,N_4359,N_4786);
nand UO_876 (O_876,N_4420,N_4239);
xor UO_877 (O_877,N_4878,N_4447);
nor UO_878 (O_878,N_4389,N_4745);
nor UO_879 (O_879,N_4216,N_4687);
xnor UO_880 (O_880,N_4082,N_4198);
and UO_881 (O_881,N_4475,N_4726);
xnor UO_882 (O_882,N_4829,N_4029);
xor UO_883 (O_883,N_4786,N_4417);
xor UO_884 (O_884,N_4226,N_4905);
or UO_885 (O_885,N_4902,N_4667);
and UO_886 (O_886,N_4580,N_4808);
or UO_887 (O_887,N_4026,N_4855);
or UO_888 (O_888,N_4035,N_4604);
nor UO_889 (O_889,N_4347,N_4056);
nand UO_890 (O_890,N_4192,N_4489);
nand UO_891 (O_891,N_4638,N_4176);
nand UO_892 (O_892,N_4518,N_4517);
nand UO_893 (O_893,N_4056,N_4390);
or UO_894 (O_894,N_4645,N_4518);
nand UO_895 (O_895,N_4100,N_4908);
nor UO_896 (O_896,N_4682,N_4466);
or UO_897 (O_897,N_4813,N_4299);
nor UO_898 (O_898,N_4341,N_4419);
nor UO_899 (O_899,N_4411,N_4945);
nor UO_900 (O_900,N_4214,N_4374);
xnor UO_901 (O_901,N_4836,N_4372);
or UO_902 (O_902,N_4465,N_4680);
or UO_903 (O_903,N_4394,N_4990);
nor UO_904 (O_904,N_4852,N_4252);
nor UO_905 (O_905,N_4951,N_4237);
or UO_906 (O_906,N_4567,N_4008);
or UO_907 (O_907,N_4633,N_4610);
xnor UO_908 (O_908,N_4483,N_4354);
nor UO_909 (O_909,N_4681,N_4268);
and UO_910 (O_910,N_4277,N_4301);
nand UO_911 (O_911,N_4689,N_4799);
nand UO_912 (O_912,N_4530,N_4186);
nor UO_913 (O_913,N_4015,N_4851);
nor UO_914 (O_914,N_4635,N_4065);
and UO_915 (O_915,N_4978,N_4748);
xor UO_916 (O_916,N_4019,N_4008);
xnor UO_917 (O_917,N_4087,N_4989);
and UO_918 (O_918,N_4626,N_4234);
xor UO_919 (O_919,N_4689,N_4623);
and UO_920 (O_920,N_4647,N_4519);
nor UO_921 (O_921,N_4454,N_4524);
or UO_922 (O_922,N_4978,N_4910);
nor UO_923 (O_923,N_4693,N_4752);
nand UO_924 (O_924,N_4308,N_4682);
and UO_925 (O_925,N_4570,N_4450);
xnor UO_926 (O_926,N_4911,N_4136);
xnor UO_927 (O_927,N_4747,N_4478);
xnor UO_928 (O_928,N_4809,N_4896);
nor UO_929 (O_929,N_4944,N_4532);
nor UO_930 (O_930,N_4311,N_4360);
and UO_931 (O_931,N_4533,N_4202);
nor UO_932 (O_932,N_4900,N_4070);
and UO_933 (O_933,N_4122,N_4600);
or UO_934 (O_934,N_4812,N_4708);
and UO_935 (O_935,N_4217,N_4014);
or UO_936 (O_936,N_4449,N_4326);
nand UO_937 (O_937,N_4590,N_4402);
xnor UO_938 (O_938,N_4472,N_4032);
or UO_939 (O_939,N_4562,N_4232);
xnor UO_940 (O_940,N_4485,N_4708);
or UO_941 (O_941,N_4837,N_4049);
xor UO_942 (O_942,N_4541,N_4878);
or UO_943 (O_943,N_4718,N_4275);
nand UO_944 (O_944,N_4449,N_4351);
and UO_945 (O_945,N_4017,N_4446);
nor UO_946 (O_946,N_4614,N_4094);
nor UO_947 (O_947,N_4061,N_4583);
xnor UO_948 (O_948,N_4495,N_4611);
nor UO_949 (O_949,N_4740,N_4516);
xnor UO_950 (O_950,N_4260,N_4115);
nor UO_951 (O_951,N_4718,N_4107);
nor UO_952 (O_952,N_4985,N_4289);
xor UO_953 (O_953,N_4125,N_4201);
and UO_954 (O_954,N_4535,N_4058);
nor UO_955 (O_955,N_4785,N_4115);
nand UO_956 (O_956,N_4354,N_4417);
or UO_957 (O_957,N_4654,N_4340);
and UO_958 (O_958,N_4459,N_4189);
nor UO_959 (O_959,N_4502,N_4802);
xor UO_960 (O_960,N_4559,N_4258);
or UO_961 (O_961,N_4947,N_4942);
nand UO_962 (O_962,N_4423,N_4756);
nor UO_963 (O_963,N_4547,N_4074);
nor UO_964 (O_964,N_4345,N_4496);
nor UO_965 (O_965,N_4255,N_4891);
xor UO_966 (O_966,N_4107,N_4806);
xor UO_967 (O_967,N_4641,N_4774);
and UO_968 (O_968,N_4755,N_4251);
or UO_969 (O_969,N_4470,N_4759);
and UO_970 (O_970,N_4586,N_4596);
xnor UO_971 (O_971,N_4415,N_4330);
and UO_972 (O_972,N_4122,N_4751);
nand UO_973 (O_973,N_4584,N_4595);
xnor UO_974 (O_974,N_4269,N_4230);
xor UO_975 (O_975,N_4940,N_4368);
xnor UO_976 (O_976,N_4353,N_4650);
nor UO_977 (O_977,N_4925,N_4168);
nor UO_978 (O_978,N_4616,N_4818);
xor UO_979 (O_979,N_4082,N_4211);
nand UO_980 (O_980,N_4919,N_4842);
or UO_981 (O_981,N_4045,N_4017);
nor UO_982 (O_982,N_4743,N_4080);
and UO_983 (O_983,N_4537,N_4262);
nor UO_984 (O_984,N_4966,N_4039);
or UO_985 (O_985,N_4444,N_4641);
xor UO_986 (O_986,N_4330,N_4030);
or UO_987 (O_987,N_4581,N_4623);
or UO_988 (O_988,N_4541,N_4826);
or UO_989 (O_989,N_4679,N_4157);
or UO_990 (O_990,N_4298,N_4094);
or UO_991 (O_991,N_4593,N_4231);
and UO_992 (O_992,N_4889,N_4879);
and UO_993 (O_993,N_4786,N_4368);
xor UO_994 (O_994,N_4842,N_4908);
or UO_995 (O_995,N_4671,N_4655);
or UO_996 (O_996,N_4562,N_4938);
and UO_997 (O_997,N_4412,N_4967);
nor UO_998 (O_998,N_4495,N_4068);
or UO_999 (O_999,N_4876,N_4241);
endmodule