module basic_500_3000_500_3_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_254,In_53);
nor U1 (N_1,In_19,In_224);
xor U2 (N_2,In_100,In_433);
nand U3 (N_3,In_289,In_85);
nand U4 (N_4,In_286,In_364);
nand U5 (N_5,In_275,In_251);
nor U6 (N_6,In_367,In_299);
nor U7 (N_7,In_134,In_336);
and U8 (N_8,In_274,In_448);
xor U9 (N_9,In_123,In_140);
nor U10 (N_10,In_313,In_248);
nor U11 (N_11,In_384,In_147);
and U12 (N_12,In_344,In_440);
xor U13 (N_13,In_253,In_241);
or U14 (N_14,In_290,In_482);
nor U15 (N_15,In_304,In_175);
or U16 (N_16,In_128,In_291);
nor U17 (N_17,In_6,In_131);
nand U18 (N_18,In_185,In_239);
xor U19 (N_19,In_9,In_71);
nand U20 (N_20,In_112,In_233);
or U21 (N_21,In_425,In_473);
nor U22 (N_22,In_74,In_193);
nand U23 (N_23,In_234,In_41);
and U24 (N_24,In_62,In_387);
and U25 (N_25,In_466,In_386);
nor U26 (N_26,In_446,In_468);
xnor U27 (N_27,In_495,In_132);
nor U28 (N_28,In_212,In_334);
nor U29 (N_29,In_207,In_476);
and U30 (N_30,In_279,In_317);
or U31 (N_31,In_158,In_340);
and U32 (N_32,In_283,In_150);
nor U33 (N_33,In_481,In_219);
nand U34 (N_34,In_264,In_23);
or U35 (N_35,In_230,In_428);
nand U36 (N_36,In_121,In_327);
nor U37 (N_37,In_113,In_410);
nand U38 (N_38,In_104,In_249);
or U39 (N_39,In_339,In_357);
or U40 (N_40,In_399,In_187);
or U41 (N_41,In_491,In_371);
and U42 (N_42,In_430,In_320);
and U43 (N_43,In_353,In_389);
nand U44 (N_44,In_462,In_83);
and U45 (N_45,In_447,In_26);
or U46 (N_46,In_25,In_369);
and U47 (N_47,In_356,In_444);
nor U48 (N_48,In_394,In_77);
nor U49 (N_49,In_72,In_365);
nand U50 (N_50,In_48,In_12);
xnor U51 (N_51,In_217,In_429);
xnor U52 (N_52,In_359,In_377);
xor U53 (N_53,In_89,In_484);
or U54 (N_54,In_411,In_117);
or U55 (N_55,In_450,In_483);
nor U56 (N_56,In_162,In_125);
nor U57 (N_57,In_7,In_319);
and U58 (N_58,In_373,In_306);
nor U59 (N_59,In_28,In_152);
nor U60 (N_60,In_276,In_59);
and U61 (N_61,In_16,In_296);
nand U62 (N_62,In_54,In_285);
xor U63 (N_63,In_259,In_498);
xnor U64 (N_64,In_153,In_191);
nor U65 (N_65,In_159,In_27);
nor U66 (N_66,In_99,In_64);
or U67 (N_67,In_40,In_308);
and U68 (N_68,In_388,In_368);
xor U69 (N_69,In_106,In_343);
xor U70 (N_70,In_218,In_323);
nand U71 (N_71,In_402,In_326);
nor U72 (N_72,In_33,In_414);
and U73 (N_73,In_103,In_310);
and U74 (N_74,In_91,In_250);
nand U75 (N_75,In_237,In_181);
or U76 (N_76,In_374,In_171);
or U77 (N_77,In_269,In_427);
nor U78 (N_78,In_38,In_216);
and U79 (N_79,In_314,In_149);
nor U80 (N_80,In_20,In_166);
and U81 (N_81,In_409,In_452);
xnor U82 (N_82,In_332,In_209);
nand U83 (N_83,In_305,In_309);
nand U84 (N_84,In_78,In_438);
nor U85 (N_85,In_8,In_288);
nor U86 (N_86,In_397,In_490);
nor U87 (N_87,In_324,In_318);
nand U88 (N_88,In_203,In_380);
nor U89 (N_89,In_129,In_330);
nor U90 (N_90,In_403,In_335);
and U91 (N_91,In_110,In_111);
nand U92 (N_92,In_115,In_499);
nor U93 (N_93,In_454,In_352);
nand U94 (N_94,In_180,In_381);
nand U95 (N_95,In_328,In_126);
nand U96 (N_96,In_116,In_56);
nor U97 (N_97,In_136,In_376);
nand U98 (N_98,In_1,In_118);
nor U99 (N_99,In_92,In_451);
xor U100 (N_100,In_124,In_142);
xor U101 (N_101,In_292,In_127);
nor U102 (N_102,In_281,In_173);
or U103 (N_103,In_231,In_453);
and U104 (N_104,In_170,In_297);
and U105 (N_105,In_199,In_391);
and U106 (N_106,In_408,In_145);
nor U107 (N_107,In_60,In_457);
or U108 (N_108,In_412,In_138);
nand U109 (N_109,In_119,In_114);
nand U110 (N_110,In_229,In_354);
nor U111 (N_111,In_407,In_17);
and U112 (N_112,In_467,In_315);
nand U113 (N_113,In_24,In_489);
nor U114 (N_114,In_32,In_325);
xnor U115 (N_115,In_94,In_434);
or U116 (N_116,In_105,In_29);
xnor U117 (N_117,In_277,In_268);
or U118 (N_118,In_478,In_141);
nor U119 (N_119,In_210,In_69);
xor U120 (N_120,In_198,In_243);
nand U121 (N_121,In_68,In_192);
nor U122 (N_122,In_460,In_255);
and U123 (N_123,In_280,In_82);
xnor U124 (N_124,In_98,In_443);
and U125 (N_125,In_225,In_178);
xor U126 (N_126,In_95,In_302);
and U127 (N_127,In_362,In_420);
nor U128 (N_128,In_307,In_261);
and U129 (N_129,In_223,In_445);
nor U130 (N_130,In_190,In_439);
and U131 (N_131,In_266,In_70);
or U132 (N_132,In_139,In_151);
xor U133 (N_133,In_167,In_456);
nor U134 (N_134,In_176,In_404);
or U135 (N_135,In_256,In_197);
or U136 (N_136,In_455,In_86);
nor U137 (N_137,In_247,In_252);
nor U138 (N_138,In_44,In_66);
xor U139 (N_139,In_186,In_101);
xor U140 (N_140,In_465,In_35);
or U141 (N_141,In_265,In_246);
or U142 (N_142,In_177,In_431);
or U143 (N_143,In_272,In_188);
or U144 (N_144,In_400,In_437);
nand U145 (N_145,In_161,In_284);
xor U146 (N_146,In_39,In_497);
and U147 (N_147,In_337,In_73);
xnor U148 (N_148,In_2,In_204);
nor U149 (N_149,In_90,In_107);
and U150 (N_150,In_160,In_316);
or U151 (N_151,In_169,In_65);
xor U152 (N_152,In_10,In_485);
or U153 (N_153,In_358,In_383);
nand U154 (N_154,In_165,In_31);
xor U155 (N_155,In_287,In_293);
or U156 (N_156,In_480,In_458);
nand U157 (N_157,In_79,In_208);
xor U158 (N_158,In_257,In_267);
or U159 (N_159,In_57,In_361);
and U160 (N_160,In_424,In_154);
and U161 (N_161,In_228,In_14);
xor U162 (N_162,In_442,In_345);
xnor U163 (N_163,In_242,In_232);
nand U164 (N_164,In_236,In_338);
and U165 (N_165,In_172,In_360);
nand U166 (N_166,In_262,In_461);
nand U167 (N_167,In_182,In_312);
nand U168 (N_168,In_469,In_479);
xor U169 (N_169,In_213,In_441);
or U170 (N_170,In_379,In_395);
nor U171 (N_171,In_108,In_15);
nand U172 (N_172,In_63,In_370);
and U173 (N_173,In_390,In_195);
or U174 (N_174,In_80,In_67);
nand U175 (N_175,In_496,In_258);
and U176 (N_176,In_55,In_494);
or U177 (N_177,In_164,In_144);
or U178 (N_178,In_202,In_93);
nand U179 (N_179,In_303,In_470);
or U180 (N_180,In_435,In_426);
nor U181 (N_181,In_245,In_240);
nand U182 (N_182,In_96,In_342);
xor U183 (N_183,In_22,In_130);
nor U184 (N_184,In_235,In_156);
nor U185 (N_185,In_474,In_449);
xor U186 (N_186,In_351,In_263);
or U187 (N_187,In_346,In_419);
or U188 (N_188,In_350,In_87);
nor U189 (N_189,In_133,In_422);
or U190 (N_190,In_413,In_406);
nand U191 (N_191,In_322,In_13);
xor U192 (N_192,In_168,In_51);
and U193 (N_193,In_393,In_492);
xnor U194 (N_194,In_238,In_260);
or U195 (N_195,In_163,In_421);
and U196 (N_196,In_416,In_21);
and U197 (N_197,In_477,In_45);
or U198 (N_198,In_5,In_157);
or U199 (N_199,In_475,In_464);
nor U200 (N_200,In_401,In_11);
or U201 (N_201,In_146,In_463);
xor U202 (N_202,In_183,In_58);
and U203 (N_203,In_174,In_417);
nand U204 (N_204,In_331,In_321);
and U205 (N_205,In_301,In_135);
nor U206 (N_206,In_333,In_355);
xnor U207 (N_207,In_366,In_4);
or U208 (N_208,In_184,In_436);
or U209 (N_209,In_222,In_221);
and U210 (N_210,In_52,In_47);
nand U211 (N_211,In_423,In_372);
nand U212 (N_212,In_418,In_122);
nor U213 (N_213,In_271,In_148);
and U214 (N_214,In_196,In_205);
and U215 (N_215,In_244,In_300);
and U216 (N_216,In_363,In_194);
nand U217 (N_217,In_18,In_415);
and U218 (N_218,In_405,In_226);
nand U219 (N_219,In_102,In_214);
nor U220 (N_220,In_432,In_200);
nand U221 (N_221,In_347,In_329);
xnor U222 (N_222,In_487,In_382);
or U223 (N_223,In_76,In_0);
nand U224 (N_224,In_282,In_385);
or U225 (N_225,In_155,In_46);
xnor U226 (N_226,In_36,In_220);
and U227 (N_227,In_49,In_88);
xor U228 (N_228,In_472,In_295);
and U229 (N_229,In_298,In_398);
and U230 (N_230,In_273,In_392);
and U231 (N_231,In_179,In_459);
xor U232 (N_232,In_3,In_227);
and U233 (N_233,In_278,In_375);
nand U234 (N_234,In_488,In_109);
nor U235 (N_235,In_396,In_97);
nand U236 (N_236,In_120,In_42);
or U237 (N_237,In_81,In_486);
nor U238 (N_238,In_201,In_30);
nor U239 (N_239,In_270,In_211);
or U240 (N_240,In_143,In_75);
xor U241 (N_241,In_61,In_50);
nor U242 (N_242,In_493,In_34);
or U243 (N_243,In_84,In_43);
nor U244 (N_244,In_471,In_349);
xnor U245 (N_245,In_37,In_311);
xor U246 (N_246,In_378,In_348);
and U247 (N_247,In_189,In_206);
xnor U248 (N_248,In_215,In_294);
xnor U249 (N_249,In_341,In_137);
and U250 (N_250,In_381,In_375);
or U251 (N_251,In_67,In_225);
nor U252 (N_252,In_443,In_148);
xor U253 (N_253,In_422,In_83);
xnor U254 (N_254,In_237,In_365);
and U255 (N_255,In_150,In_125);
and U256 (N_256,In_354,In_334);
or U257 (N_257,In_282,In_121);
or U258 (N_258,In_114,In_224);
and U259 (N_259,In_423,In_69);
xor U260 (N_260,In_467,In_75);
and U261 (N_261,In_188,In_419);
nand U262 (N_262,In_216,In_386);
and U263 (N_263,In_207,In_190);
and U264 (N_264,In_158,In_218);
xor U265 (N_265,In_469,In_7);
or U266 (N_266,In_69,In_46);
nor U267 (N_267,In_137,In_438);
xnor U268 (N_268,In_78,In_106);
nand U269 (N_269,In_377,In_168);
or U270 (N_270,In_89,In_479);
and U271 (N_271,In_75,In_122);
xnor U272 (N_272,In_396,In_300);
and U273 (N_273,In_107,In_183);
nand U274 (N_274,In_181,In_367);
nor U275 (N_275,In_441,In_302);
xnor U276 (N_276,In_46,In_397);
nand U277 (N_277,In_296,In_308);
nor U278 (N_278,In_136,In_69);
and U279 (N_279,In_409,In_221);
nand U280 (N_280,In_138,In_208);
xnor U281 (N_281,In_53,In_342);
nand U282 (N_282,In_79,In_156);
and U283 (N_283,In_155,In_336);
or U284 (N_284,In_215,In_351);
xor U285 (N_285,In_195,In_426);
or U286 (N_286,In_269,In_166);
and U287 (N_287,In_132,In_488);
and U288 (N_288,In_86,In_479);
or U289 (N_289,In_487,In_50);
nand U290 (N_290,In_62,In_339);
and U291 (N_291,In_351,In_47);
and U292 (N_292,In_106,In_406);
and U293 (N_293,In_444,In_73);
nor U294 (N_294,In_31,In_8);
and U295 (N_295,In_128,In_301);
nand U296 (N_296,In_479,In_322);
xnor U297 (N_297,In_187,In_386);
or U298 (N_298,In_70,In_425);
nor U299 (N_299,In_217,In_492);
nand U300 (N_300,In_57,In_257);
nor U301 (N_301,In_231,In_155);
nor U302 (N_302,In_35,In_436);
nand U303 (N_303,In_408,In_224);
nand U304 (N_304,In_106,In_399);
and U305 (N_305,In_368,In_29);
xnor U306 (N_306,In_262,In_195);
and U307 (N_307,In_231,In_111);
xnor U308 (N_308,In_192,In_39);
or U309 (N_309,In_318,In_396);
and U310 (N_310,In_464,In_60);
nor U311 (N_311,In_2,In_70);
or U312 (N_312,In_174,In_454);
nor U313 (N_313,In_420,In_49);
nand U314 (N_314,In_274,In_213);
or U315 (N_315,In_1,In_394);
nand U316 (N_316,In_178,In_149);
nor U317 (N_317,In_288,In_236);
nor U318 (N_318,In_19,In_24);
xor U319 (N_319,In_357,In_180);
nand U320 (N_320,In_356,In_153);
or U321 (N_321,In_472,In_370);
nand U322 (N_322,In_346,In_318);
nor U323 (N_323,In_257,In_263);
xor U324 (N_324,In_203,In_158);
or U325 (N_325,In_437,In_314);
xor U326 (N_326,In_488,In_101);
nor U327 (N_327,In_259,In_437);
nor U328 (N_328,In_31,In_205);
nor U329 (N_329,In_487,In_70);
or U330 (N_330,In_177,In_335);
and U331 (N_331,In_151,In_446);
nor U332 (N_332,In_389,In_186);
nand U333 (N_333,In_446,In_430);
nand U334 (N_334,In_259,In_33);
or U335 (N_335,In_312,In_10);
nor U336 (N_336,In_438,In_378);
and U337 (N_337,In_58,In_86);
xor U338 (N_338,In_490,In_339);
nand U339 (N_339,In_350,In_376);
nor U340 (N_340,In_258,In_468);
and U341 (N_341,In_56,In_171);
or U342 (N_342,In_237,In_34);
or U343 (N_343,In_66,In_85);
xor U344 (N_344,In_2,In_160);
xor U345 (N_345,In_272,In_264);
xor U346 (N_346,In_108,In_183);
or U347 (N_347,In_377,In_51);
nor U348 (N_348,In_114,In_446);
nand U349 (N_349,In_499,In_171);
nand U350 (N_350,In_43,In_198);
and U351 (N_351,In_126,In_371);
nor U352 (N_352,In_40,In_87);
nand U353 (N_353,In_417,In_81);
nor U354 (N_354,In_24,In_291);
or U355 (N_355,In_105,In_455);
and U356 (N_356,In_439,In_287);
xor U357 (N_357,In_394,In_62);
or U358 (N_358,In_394,In_293);
nand U359 (N_359,In_377,In_391);
nor U360 (N_360,In_181,In_463);
xor U361 (N_361,In_54,In_397);
and U362 (N_362,In_219,In_215);
nand U363 (N_363,In_132,In_253);
nor U364 (N_364,In_473,In_118);
nor U365 (N_365,In_489,In_212);
nand U366 (N_366,In_220,In_343);
xor U367 (N_367,In_52,In_234);
xnor U368 (N_368,In_311,In_350);
and U369 (N_369,In_296,In_347);
xor U370 (N_370,In_318,In_196);
or U371 (N_371,In_292,In_336);
xnor U372 (N_372,In_19,In_288);
or U373 (N_373,In_2,In_377);
nand U374 (N_374,In_92,In_35);
and U375 (N_375,In_197,In_148);
nand U376 (N_376,In_415,In_373);
and U377 (N_377,In_294,In_2);
or U378 (N_378,In_90,In_185);
nor U379 (N_379,In_85,In_303);
and U380 (N_380,In_353,In_106);
nor U381 (N_381,In_362,In_285);
nand U382 (N_382,In_154,In_140);
nand U383 (N_383,In_378,In_273);
or U384 (N_384,In_75,In_100);
nor U385 (N_385,In_5,In_358);
nor U386 (N_386,In_163,In_55);
xnor U387 (N_387,In_389,In_183);
nand U388 (N_388,In_455,In_149);
nand U389 (N_389,In_159,In_342);
xnor U390 (N_390,In_182,In_390);
xnor U391 (N_391,In_150,In_287);
nand U392 (N_392,In_406,In_41);
xnor U393 (N_393,In_325,In_45);
xor U394 (N_394,In_184,In_412);
xor U395 (N_395,In_156,In_368);
xor U396 (N_396,In_18,In_483);
nor U397 (N_397,In_55,In_53);
and U398 (N_398,In_368,In_382);
or U399 (N_399,In_468,In_239);
nor U400 (N_400,In_24,In_36);
or U401 (N_401,In_449,In_313);
xnor U402 (N_402,In_4,In_352);
nand U403 (N_403,In_36,In_380);
nor U404 (N_404,In_328,In_47);
nand U405 (N_405,In_340,In_79);
nand U406 (N_406,In_106,In_209);
xor U407 (N_407,In_347,In_45);
or U408 (N_408,In_479,In_198);
or U409 (N_409,In_76,In_11);
nand U410 (N_410,In_382,In_242);
nor U411 (N_411,In_45,In_36);
and U412 (N_412,In_485,In_38);
nor U413 (N_413,In_423,In_293);
or U414 (N_414,In_279,In_41);
or U415 (N_415,In_36,In_197);
nor U416 (N_416,In_441,In_65);
and U417 (N_417,In_287,In_473);
nor U418 (N_418,In_283,In_437);
xnor U419 (N_419,In_280,In_288);
or U420 (N_420,In_341,In_381);
xnor U421 (N_421,In_297,In_331);
xnor U422 (N_422,In_101,In_11);
nor U423 (N_423,In_341,In_37);
nand U424 (N_424,In_57,In_490);
nand U425 (N_425,In_170,In_0);
or U426 (N_426,In_111,In_159);
or U427 (N_427,In_271,In_4);
or U428 (N_428,In_152,In_291);
or U429 (N_429,In_38,In_282);
nand U430 (N_430,In_127,In_154);
nand U431 (N_431,In_462,In_78);
and U432 (N_432,In_470,In_16);
xnor U433 (N_433,In_390,In_153);
xor U434 (N_434,In_61,In_274);
nand U435 (N_435,In_375,In_29);
nand U436 (N_436,In_381,In_290);
nand U437 (N_437,In_34,In_473);
or U438 (N_438,In_436,In_243);
nand U439 (N_439,In_186,In_89);
nor U440 (N_440,In_301,In_343);
or U441 (N_441,In_301,In_325);
nor U442 (N_442,In_126,In_115);
and U443 (N_443,In_454,In_134);
nand U444 (N_444,In_325,In_6);
and U445 (N_445,In_119,In_366);
or U446 (N_446,In_11,In_430);
xor U447 (N_447,In_106,In_459);
and U448 (N_448,In_411,In_8);
and U449 (N_449,In_416,In_335);
nor U450 (N_450,In_402,In_65);
xor U451 (N_451,In_47,In_383);
or U452 (N_452,In_462,In_351);
nor U453 (N_453,In_88,In_363);
or U454 (N_454,In_160,In_192);
xor U455 (N_455,In_398,In_58);
xor U456 (N_456,In_158,In_196);
nor U457 (N_457,In_433,In_365);
nor U458 (N_458,In_360,In_49);
nand U459 (N_459,In_88,In_107);
xnor U460 (N_460,In_147,In_335);
xor U461 (N_461,In_399,In_56);
nor U462 (N_462,In_449,In_32);
or U463 (N_463,In_486,In_59);
nand U464 (N_464,In_248,In_356);
nor U465 (N_465,In_22,In_115);
nor U466 (N_466,In_73,In_124);
xnor U467 (N_467,In_146,In_336);
nor U468 (N_468,In_40,In_481);
nor U469 (N_469,In_292,In_349);
or U470 (N_470,In_143,In_272);
nor U471 (N_471,In_147,In_311);
and U472 (N_472,In_384,In_135);
or U473 (N_473,In_300,In_193);
xnor U474 (N_474,In_82,In_96);
nor U475 (N_475,In_179,In_450);
nand U476 (N_476,In_107,In_314);
and U477 (N_477,In_372,In_227);
nand U478 (N_478,In_48,In_232);
nor U479 (N_479,In_475,In_220);
xor U480 (N_480,In_9,In_74);
nor U481 (N_481,In_491,In_221);
nor U482 (N_482,In_316,In_381);
nand U483 (N_483,In_321,In_484);
nand U484 (N_484,In_238,In_12);
or U485 (N_485,In_54,In_487);
nor U486 (N_486,In_430,In_292);
nor U487 (N_487,In_328,In_94);
or U488 (N_488,In_475,In_26);
nor U489 (N_489,In_418,In_117);
nand U490 (N_490,In_398,In_225);
xor U491 (N_491,In_22,In_87);
nor U492 (N_492,In_373,In_233);
and U493 (N_493,In_30,In_494);
nor U494 (N_494,In_83,In_85);
nor U495 (N_495,In_344,In_349);
nor U496 (N_496,In_381,In_159);
or U497 (N_497,In_430,In_101);
nand U498 (N_498,In_173,In_102);
or U499 (N_499,In_411,In_252);
xnor U500 (N_500,In_200,In_447);
or U501 (N_501,In_496,In_423);
or U502 (N_502,In_430,In_499);
and U503 (N_503,In_45,In_195);
nor U504 (N_504,In_70,In_290);
or U505 (N_505,In_185,In_20);
xor U506 (N_506,In_266,In_224);
nor U507 (N_507,In_364,In_98);
nor U508 (N_508,In_324,In_417);
xnor U509 (N_509,In_169,In_273);
nand U510 (N_510,In_24,In_273);
or U511 (N_511,In_94,In_352);
and U512 (N_512,In_119,In_343);
nand U513 (N_513,In_464,In_71);
nand U514 (N_514,In_283,In_239);
xnor U515 (N_515,In_362,In_396);
and U516 (N_516,In_224,In_407);
xnor U517 (N_517,In_437,In_358);
xor U518 (N_518,In_11,In_298);
nand U519 (N_519,In_405,In_312);
xnor U520 (N_520,In_497,In_121);
and U521 (N_521,In_378,In_312);
and U522 (N_522,In_262,In_385);
and U523 (N_523,In_424,In_288);
and U524 (N_524,In_421,In_398);
and U525 (N_525,In_7,In_445);
nor U526 (N_526,In_496,In_327);
or U527 (N_527,In_60,In_145);
nand U528 (N_528,In_210,In_361);
or U529 (N_529,In_463,In_445);
nor U530 (N_530,In_100,In_343);
or U531 (N_531,In_445,In_487);
xnor U532 (N_532,In_245,In_263);
nand U533 (N_533,In_118,In_54);
nand U534 (N_534,In_390,In_17);
nor U535 (N_535,In_311,In_485);
nand U536 (N_536,In_146,In_51);
xnor U537 (N_537,In_477,In_208);
xor U538 (N_538,In_497,In_286);
or U539 (N_539,In_95,In_45);
and U540 (N_540,In_228,In_177);
nor U541 (N_541,In_275,In_499);
xor U542 (N_542,In_228,In_440);
or U543 (N_543,In_497,In_155);
and U544 (N_544,In_271,In_383);
or U545 (N_545,In_192,In_105);
and U546 (N_546,In_88,In_108);
xnor U547 (N_547,In_322,In_9);
and U548 (N_548,In_132,In_448);
nand U549 (N_549,In_487,In_46);
nand U550 (N_550,In_313,In_185);
nor U551 (N_551,In_477,In_206);
nand U552 (N_552,In_222,In_270);
or U553 (N_553,In_307,In_96);
nand U554 (N_554,In_6,In_389);
xnor U555 (N_555,In_335,In_172);
or U556 (N_556,In_485,In_149);
or U557 (N_557,In_65,In_192);
xor U558 (N_558,In_425,In_14);
nand U559 (N_559,In_377,In_237);
and U560 (N_560,In_122,In_349);
or U561 (N_561,In_16,In_455);
xnor U562 (N_562,In_143,In_21);
and U563 (N_563,In_456,In_439);
nand U564 (N_564,In_162,In_334);
nor U565 (N_565,In_472,In_234);
and U566 (N_566,In_399,In_72);
or U567 (N_567,In_334,In_297);
xor U568 (N_568,In_98,In_6);
or U569 (N_569,In_86,In_239);
nand U570 (N_570,In_317,In_349);
nand U571 (N_571,In_246,In_45);
nor U572 (N_572,In_337,In_291);
or U573 (N_573,In_215,In_115);
nor U574 (N_574,In_2,In_40);
or U575 (N_575,In_151,In_448);
nand U576 (N_576,In_71,In_339);
or U577 (N_577,In_459,In_436);
xnor U578 (N_578,In_211,In_208);
xnor U579 (N_579,In_355,In_303);
xnor U580 (N_580,In_286,In_35);
and U581 (N_581,In_221,In_413);
or U582 (N_582,In_166,In_434);
or U583 (N_583,In_456,In_93);
nor U584 (N_584,In_311,In_285);
nand U585 (N_585,In_343,In_135);
nor U586 (N_586,In_157,In_199);
or U587 (N_587,In_314,In_315);
xor U588 (N_588,In_196,In_399);
and U589 (N_589,In_222,In_429);
or U590 (N_590,In_167,In_230);
and U591 (N_591,In_490,In_219);
or U592 (N_592,In_385,In_81);
and U593 (N_593,In_27,In_175);
or U594 (N_594,In_132,In_77);
xnor U595 (N_595,In_93,In_252);
xnor U596 (N_596,In_288,In_349);
xnor U597 (N_597,In_257,In_453);
or U598 (N_598,In_119,In_279);
and U599 (N_599,In_143,In_455);
and U600 (N_600,In_130,In_457);
or U601 (N_601,In_129,In_229);
nand U602 (N_602,In_368,In_399);
or U603 (N_603,In_239,In_124);
and U604 (N_604,In_64,In_141);
nand U605 (N_605,In_49,In_76);
or U606 (N_606,In_245,In_466);
nand U607 (N_607,In_494,In_231);
nand U608 (N_608,In_86,In_445);
and U609 (N_609,In_11,In_242);
or U610 (N_610,In_252,In_400);
nor U611 (N_611,In_289,In_390);
nand U612 (N_612,In_453,In_456);
and U613 (N_613,In_195,In_440);
and U614 (N_614,In_144,In_390);
xnor U615 (N_615,In_485,In_280);
or U616 (N_616,In_257,In_122);
and U617 (N_617,In_53,In_462);
xnor U618 (N_618,In_152,In_470);
and U619 (N_619,In_46,In_264);
and U620 (N_620,In_497,In_323);
and U621 (N_621,In_196,In_430);
nor U622 (N_622,In_333,In_460);
nor U623 (N_623,In_336,In_248);
or U624 (N_624,In_271,In_417);
and U625 (N_625,In_130,In_118);
or U626 (N_626,In_268,In_297);
nand U627 (N_627,In_411,In_130);
nand U628 (N_628,In_350,In_371);
nand U629 (N_629,In_403,In_118);
xnor U630 (N_630,In_223,In_312);
and U631 (N_631,In_1,In_46);
nor U632 (N_632,In_296,In_425);
and U633 (N_633,In_402,In_261);
nor U634 (N_634,In_80,In_426);
nand U635 (N_635,In_234,In_397);
xnor U636 (N_636,In_418,In_223);
and U637 (N_637,In_365,In_201);
nand U638 (N_638,In_149,In_441);
or U639 (N_639,In_101,In_319);
xnor U640 (N_640,In_80,In_107);
nor U641 (N_641,In_149,In_409);
nand U642 (N_642,In_365,In_203);
and U643 (N_643,In_51,In_227);
xnor U644 (N_644,In_211,In_331);
xnor U645 (N_645,In_390,In_113);
nand U646 (N_646,In_27,In_324);
and U647 (N_647,In_341,In_237);
and U648 (N_648,In_49,In_451);
nor U649 (N_649,In_375,In_231);
nand U650 (N_650,In_296,In_211);
and U651 (N_651,In_43,In_275);
and U652 (N_652,In_422,In_226);
nor U653 (N_653,In_88,In_352);
nor U654 (N_654,In_439,In_386);
nand U655 (N_655,In_489,In_119);
nand U656 (N_656,In_379,In_380);
or U657 (N_657,In_468,In_91);
nor U658 (N_658,In_198,In_487);
xor U659 (N_659,In_319,In_477);
nor U660 (N_660,In_431,In_410);
and U661 (N_661,In_338,In_262);
nand U662 (N_662,In_356,In_375);
nor U663 (N_663,In_61,In_157);
or U664 (N_664,In_17,In_85);
or U665 (N_665,In_213,In_312);
xnor U666 (N_666,In_250,In_391);
nand U667 (N_667,In_72,In_421);
nor U668 (N_668,In_112,In_236);
or U669 (N_669,In_259,In_47);
nand U670 (N_670,In_279,In_71);
or U671 (N_671,In_490,In_494);
xnor U672 (N_672,In_139,In_472);
nor U673 (N_673,In_313,In_447);
xnor U674 (N_674,In_170,In_33);
xnor U675 (N_675,In_398,In_206);
or U676 (N_676,In_453,In_296);
nor U677 (N_677,In_103,In_468);
or U678 (N_678,In_347,In_499);
xnor U679 (N_679,In_116,In_480);
nor U680 (N_680,In_380,In_315);
xor U681 (N_681,In_391,In_126);
xor U682 (N_682,In_493,In_275);
xnor U683 (N_683,In_286,In_134);
and U684 (N_684,In_130,In_443);
or U685 (N_685,In_109,In_300);
nand U686 (N_686,In_343,In_160);
or U687 (N_687,In_481,In_332);
and U688 (N_688,In_343,In_47);
xnor U689 (N_689,In_182,In_23);
nor U690 (N_690,In_339,In_77);
nor U691 (N_691,In_459,In_182);
nand U692 (N_692,In_215,In_295);
nand U693 (N_693,In_382,In_303);
nand U694 (N_694,In_35,In_391);
nand U695 (N_695,In_103,In_18);
nor U696 (N_696,In_107,In_150);
xor U697 (N_697,In_419,In_157);
xnor U698 (N_698,In_411,In_138);
xnor U699 (N_699,In_218,In_354);
xor U700 (N_700,In_413,In_283);
or U701 (N_701,In_431,In_141);
or U702 (N_702,In_262,In_460);
nor U703 (N_703,In_389,In_272);
or U704 (N_704,In_69,In_355);
xor U705 (N_705,In_495,In_490);
nor U706 (N_706,In_20,In_422);
nand U707 (N_707,In_302,In_47);
nand U708 (N_708,In_301,In_14);
or U709 (N_709,In_250,In_302);
xnor U710 (N_710,In_109,In_122);
and U711 (N_711,In_5,In_277);
and U712 (N_712,In_450,In_463);
nor U713 (N_713,In_0,In_212);
and U714 (N_714,In_261,In_333);
xnor U715 (N_715,In_49,In_236);
xor U716 (N_716,In_12,In_223);
and U717 (N_717,In_270,In_79);
or U718 (N_718,In_345,In_180);
nor U719 (N_719,In_207,In_211);
and U720 (N_720,In_457,In_211);
xnor U721 (N_721,In_211,In_182);
nand U722 (N_722,In_377,In_169);
nand U723 (N_723,In_296,In_168);
or U724 (N_724,In_372,In_392);
and U725 (N_725,In_41,In_462);
xor U726 (N_726,In_239,In_315);
nand U727 (N_727,In_182,In_35);
nor U728 (N_728,In_19,In_160);
nor U729 (N_729,In_68,In_347);
or U730 (N_730,In_68,In_121);
nand U731 (N_731,In_455,In_294);
nand U732 (N_732,In_346,In_72);
nor U733 (N_733,In_105,In_58);
xor U734 (N_734,In_349,In_104);
nor U735 (N_735,In_425,In_351);
xnor U736 (N_736,In_135,In_385);
nor U737 (N_737,In_460,In_6);
nand U738 (N_738,In_164,In_363);
xor U739 (N_739,In_169,In_107);
nand U740 (N_740,In_407,In_295);
and U741 (N_741,In_306,In_487);
nand U742 (N_742,In_491,In_30);
nor U743 (N_743,In_498,In_268);
and U744 (N_744,In_157,In_396);
nor U745 (N_745,In_162,In_88);
and U746 (N_746,In_175,In_169);
nand U747 (N_747,In_182,In_196);
and U748 (N_748,In_322,In_12);
or U749 (N_749,In_373,In_346);
nand U750 (N_750,In_474,In_365);
or U751 (N_751,In_449,In_83);
nor U752 (N_752,In_348,In_4);
or U753 (N_753,In_318,In_89);
and U754 (N_754,In_217,In_236);
nor U755 (N_755,In_221,In_246);
nor U756 (N_756,In_82,In_43);
nand U757 (N_757,In_420,In_20);
or U758 (N_758,In_5,In_337);
nor U759 (N_759,In_458,In_375);
xor U760 (N_760,In_125,In_12);
nand U761 (N_761,In_209,In_492);
nand U762 (N_762,In_443,In_395);
xnor U763 (N_763,In_5,In_409);
nand U764 (N_764,In_456,In_459);
or U765 (N_765,In_333,In_102);
or U766 (N_766,In_180,In_147);
or U767 (N_767,In_147,In_189);
and U768 (N_768,In_201,In_56);
nand U769 (N_769,In_188,In_250);
or U770 (N_770,In_154,In_448);
nand U771 (N_771,In_12,In_220);
xnor U772 (N_772,In_346,In_384);
xor U773 (N_773,In_153,In_357);
xor U774 (N_774,In_240,In_17);
xnor U775 (N_775,In_476,In_146);
nand U776 (N_776,In_378,In_163);
and U777 (N_777,In_218,In_281);
nor U778 (N_778,In_495,In_381);
and U779 (N_779,In_329,In_183);
nor U780 (N_780,In_364,In_276);
nand U781 (N_781,In_73,In_68);
nor U782 (N_782,In_492,In_223);
and U783 (N_783,In_466,In_436);
or U784 (N_784,In_176,In_58);
nand U785 (N_785,In_155,In_249);
xnor U786 (N_786,In_140,In_306);
xor U787 (N_787,In_241,In_19);
or U788 (N_788,In_14,In_379);
xor U789 (N_789,In_359,In_87);
and U790 (N_790,In_391,In_249);
xor U791 (N_791,In_240,In_149);
xor U792 (N_792,In_108,In_246);
nor U793 (N_793,In_115,In_30);
nor U794 (N_794,In_275,In_485);
or U795 (N_795,In_241,In_377);
and U796 (N_796,In_201,In_65);
nor U797 (N_797,In_306,In_493);
and U798 (N_798,In_474,In_292);
xor U799 (N_799,In_421,In_130);
and U800 (N_800,In_200,In_443);
nand U801 (N_801,In_200,In_153);
or U802 (N_802,In_54,In_474);
nor U803 (N_803,In_25,In_420);
xor U804 (N_804,In_169,In_105);
or U805 (N_805,In_486,In_276);
nor U806 (N_806,In_9,In_44);
or U807 (N_807,In_42,In_84);
nand U808 (N_808,In_210,In_33);
or U809 (N_809,In_255,In_96);
xnor U810 (N_810,In_372,In_356);
and U811 (N_811,In_290,In_327);
and U812 (N_812,In_282,In_367);
and U813 (N_813,In_31,In_493);
nor U814 (N_814,In_220,In_452);
xor U815 (N_815,In_425,In_417);
nor U816 (N_816,In_408,In_308);
xnor U817 (N_817,In_458,In_343);
nand U818 (N_818,In_330,In_494);
nor U819 (N_819,In_309,In_124);
xor U820 (N_820,In_134,In_126);
xor U821 (N_821,In_171,In_314);
nand U822 (N_822,In_205,In_14);
nor U823 (N_823,In_446,In_9);
and U824 (N_824,In_92,In_75);
nor U825 (N_825,In_86,In_196);
and U826 (N_826,In_54,In_370);
xor U827 (N_827,In_168,In_291);
and U828 (N_828,In_362,In_371);
and U829 (N_829,In_427,In_116);
nand U830 (N_830,In_137,In_350);
xor U831 (N_831,In_328,In_226);
nand U832 (N_832,In_492,In_160);
nor U833 (N_833,In_280,In_215);
nor U834 (N_834,In_217,In_321);
xnor U835 (N_835,In_425,In_408);
and U836 (N_836,In_372,In_77);
and U837 (N_837,In_172,In_151);
nand U838 (N_838,In_128,In_146);
nand U839 (N_839,In_176,In_310);
xnor U840 (N_840,In_473,In_353);
or U841 (N_841,In_416,In_256);
and U842 (N_842,In_258,In_195);
and U843 (N_843,In_491,In_20);
nor U844 (N_844,In_332,In_340);
or U845 (N_845,In_60,In_236);
nor U846 (N_846,In_451,In_282);
xor U847 (N_847,In_267,In_119);
nand U848 (N_848,In_220,In_54);
and U849 (N_849,In_80,In_353);
nor U850 (N_850,In_461,In_346);
or U851 (N_851,In_69,In_3);
nand U852 (N_852,In_230,In_43);
xor U853 (N_853,In_53,In_433);
nand U854 (N_854,In_442,In_234);
and U855 (N_855,In_459,In_38);
nand U856 (N_856,In_329,In_131);
xnor U857 (N_857,In_153,In_306);
nand U858 (N_858,In_16,In_70);
xor U859 (N_859,In_378,In_141);
nand U860 (N_860,In_126,In_401);
and U861 (N_861,In_388,In_484);
nand U862 (N_862,In_27,In_389);
nand U863 (N_863,In_348,In_35);
or U864 (N_864,In_363,In_470);
or U865 (N_865,In_453,In_49);
nand U866 (N_866,In_259,In_73);
xor U867 (N_867,In_382,In_43);
nand U868 (N_868,In_384,In_284);
and U869 (N_869,In_280,In_113);
nor U870 (N_870,In_270,In_57);
or U871 (N_871,In_34,In_340);
and U872 (N_872,In_469,In_6);
and U873 (N_873,In_441,In_279);
xnor U874 (N_874,In_406,In_262);
or U875 (N_875,In_315,In_175);
nand U876 (N_876,In_53,In_9);
and U877 (N_877,In_138,In_82);
xor U878 (N_878,In_170,In_383);
and U879 (N_879,In_384,In_97);
nand U880 (N_880,In_125,In_494);
nand U881 (N_881,In_308,In_466);
xor U882 (N_882,In_43,In_259);
xnor U883 (N_883,In_299,In_432);
nand U884 (N_884,In_332,In_496);
nor U885 (N_885,In_378,In_149);
nor U886 (N_886,In_74,In_428);
or U887 (N_887,In_279,In_197);
xnor U888 (N_888,In_217,In_1);
nor U889 (N_889,In_164,In_318);
and U890 (N_890,In_17,In_107);
nor U891 (N_891,In_309,In_413);
xnor U892 (N_892,In_238,In_248);
xnor U893 (N_893,In_86,In_90);
or U894 (N_894,In_360,In_461);
xor U895 (N_895,In_159,In_446);
or U896 (N_896,In_423,In_190);
xnor U897 (N_897,In_455,In_304);
or U898 (N_898,In_64,In_42);
and U899 (N_899,In_85,In_199);
or U900 (N_900,In_444,In_77);
or U901 (N_901,In_35,In_253);
and U902 (N_902,In_230,In_369);
nand U903 (N_903,In_334,In_74);
nand U904 (N_904,In_498,In_145);
nand U905 (N_905,In_443,In_211);
or U906 (N_906,In_390,In_139);
nor U907 (N_907,In_420,In_37);
or U908 (N_908,In_84,In_175);
or U909 (N_909,In_152,In_329);
xnor U910 (N_910,In_250,In_381);
xnor U911 (N_911,In_427,In_171);
or U912 (N_912,In_297,In_448);
and U913 (N_913,In_95,In_160);
and U914 (N_914,In_50,In_223);
nand U915 (N_915,In_135,In_110);
or U916 (N_916,In_55,In_0);
or U917 (N_917,In_102,In_28);
nand U918 (N_918,In_473,In_412);
nand U919 (N_919,In_126,In_103);
xor U920 (N_920,In_485,In_252);
nand U921 (N_921,In_478,In_246);
and U922 (N_922,In_190,In_292);
and U923 (N_923,In_216,In_84);
nor U924 (N_924,In_194,In_489);
nor U925 (N_925,In_429,In_177);
xor U926 (N_926,In_388,In_18);
or U927 (N_927,In_24,In_483);
xnor U928 (N_928,In_124,In_144);
and U929 (N_929,In_296,In_217);
nor U930 (N_930,In_117,In_444);
and U931 (N_931,In_430,In_362);
nor U932 (N_932,In_237,In_416);
and U933 (N_933,In_329,In_177);
or U934 (N_934,In_389,In_245);
nand U935 (N_935,In_57,In_82);
or U936 (N_936,In_293,In_181);
nor U937 (N_937,In_412,In_207);
and U938 (N_938,In_483,In_177);
nand U939 (N_939,In_109,In_85);
nor U940 (N_940,In_405,In_285);
or U941 (N_941,In_394,In_480);
nor U942 (N_942,In_219,In_164);
nor U943 (N_943,In_89,In_361);
and U944 (N_944,In_460,In_366);
nand U945 (N_945,In_77,In_272);
nor U946 (N_946,In_201,In_6);
and U947 (N_947,In_316,In_238);
and U948 (N_948,In_364,In_202);
xor U949 (N_949,In_191,In_3);
and U950 (N_950,In_92,In_453);
nor U951 (N_951,In_351,In_287);
or U952 (N_952,In_461,In_481);
nand U953 (N_953,In_360,In_447);
nor U954 (N_954,In_86,In_16);
nor U955 (N_955,In_368,In_226);
or U956 (N_956,In_339,In_165);
and U957 (N_957,In_441,In_115);
nand U958 (N_958,In_306,In_147);
nor U959 (N_959,In_293,In_10);
nand U960 (N_960,In_428,In_184);
nand U961 (N_961,In_218,In_10);
nand U962 (N_962,In_106,In_325);
and U963 (N_963,In_456,In_425);
and U964 (N_964,In_309,In_286);
nor U965 (N_965,In_26,In_405);
xnor U966 (N_966,In_451,In_146);
nor U967 (N_967,In_455,In_300);
or U968 (N_968,In_244,In_375);
nor U969 (N_969,In_282,In_440);
nor U970 (N_970,In_130,In_450);
nand U971 (N_971,In_204,In_387);
nand U972 (N_972,In_485,In_176);
nor U973 (N_973,In_310,In_363);
nand U974 (N_974,In_366,In_98);
and U975 (N_975,In_217,In_271);
or U976 (N_976,In_292,In_43);
and U977 (N_977,In_20,In_373);
xor U978 (N_978,In_252,In_250);
xor U979 (N_979,In_179,In_97);
nand U980 (N_980,In_112,In_348);
xor U981 (N_981,In_304,In_209);
nand U982 (N_982,In_341,In_117);
nand U983 (N_983,In_222,In_153);
xnor U984 (N_984,In_289,In_109);
nand U985 (N_985,In_474,In_1);
nand U986 (N_986,In_234,In_148);
or U987 (N_987,In_299,In_23);
and U988 (N_988,In_25,In_374);
or U989 (N_989,In_42,In_274);
nand U990 (N_990,In_435,In_257);
nor U991 (N_991,In_411,In_9);
nand U992 (N_992,In_275,In_174);
and U993 (N_993,In_463,In_344);
and U994 (N_994,In_175,In_468);
nor U995 (N_995,In_362,In_398);
nand U996 (N_996,In_44,In_288);
xnor U997 (N_997,In_324,In_152);
or U998 (N_998,In_449,In_315);
nor U999 (N_999,In_135,In_331);
xor U1000 (N_1000,N_897,N_999);
or U1001 (N_1001,N_112,N_149);
or U1002 (N_1002,N_506,N_631);
xnor U1003 (N_1003,N_674,N_19);
and U1004 (N_1004,N_86,N_886);
and U1005 (N_1005,N_602,N_49);
nor U1006 (N_1006,N_662,N_643);
nor U1007 (N_1007,N_837,N_590);
or U1008 (N_1008,N_422,N_25);
nand U1009 (N_1009,N_156,N_316);
nand U1010 (N_1010,N_47,N_748);
and U1011 (N_1011,N_470,N_266);
xor U1012 (N_1012,N_677,N_731);
and U1013 (N_1013,N_418,N_834);
nor U1014 (N_1014,N_391,N_651);
and U1015 (N_1015,N_629,N_796);
nor U1016 (N_1016,N_676,N_318);
xor U1017 (N_1017,N_956,N_829);
xor U1018 (N_1018,N_571,N_606);
or U1019 (N_1019,N_910,N_314);
nand U1020 (N_1020,N_803,N_146);
xnor U1021 (N_1021,N_567,N_669);
nor U1022 (N_1022,N_957,N_797);
nand U1023 (N_1023,N_284,N_300);
and U1024 (N_1024,N_831,N_574);
nand U1025 (N_1025,N_730,N_413);
nor U1026 (N_1026,N_453,N_238);
xor U1027 (N_1027,N_951,N_13);
and U1028 (N_1028,N_489,N_340);
xnor U1029 (N_1029,N_763,N_584);
nand U1030 (N_1030,N_757,N_79);
nand U1031 (N_1031,N_558,N_896);
and U1032 (N_1032,N_587,N_988);
or U1033 (N_1033,N_331,N_166);
and U1034 (N_1034,N_273,N_424);
and U1035 (N_1035,N_889,N_172);
nand U1036 (N_1036,N_689,N_546);
xnor U1037 (N_1037,N_371,N_776);
xor U1038 (N_1038,N_881,N_769);
xor U1039 (N_1039,N_802,N_147);
nand U1040 (N_1040,N_599,N_290);
xor U1041 (N_1041,N_678,N_770);
and U1042 (N_1042,N_349,N_864);
nand U1043 (N_1043,N_772,N_621);
xnor U1044 (N_1044,N_753,N_352);
or U1045 (N_1045,N_154,N_646);
or U1046 (N_1046,N_911,N_594);
xnor U1047 (N_1047,N_667,N_395);
xnor U1048 (N_1048,N_691,N_455);
xor U1049 (N_1049,N_135,N_504);
or U1050 (N_1050,N_516,N_773);
nand U1051 (N_1051,N_171,N_980);
and U1052 (N_1052,N_232,N_698);
nand U1053 (N_1053,N_465,N_823);
nor U1054 (N_1054,N_33,N_128);
xor U1055 (N_1055,N_647,N_685);
or U1056 (N_1056,N_380,N_661);
or U1057 (N_1057,N_984,N_286);
nor U1058 (N_1058,N_281,N_777);
nor U1059 (N_1059,N_627,N_27);
and U1060 (N_1060,N_360,N_197);
and U1061 (N_1061,N_800,N_603);
or U1062 (N_1062,N_810,N_109);
nor U1063 (N_1063,N_215,N_101);
xnor U1064 (N_1064,N_952,N_588);
or U1065 (N_1065,N_376,N_616);
nor U1066 (N_1066,N_502,N_712);
and U1067 (N_1067,N_299,N_804);
nand U1068 (N_1068,N_498,N_827);
xnor U1069 (N_1069,N_877,N_219);
or U1070 (N_1070,N_63,N_509);
xor U1071 (N_1071,N_807,N_293);
and U1072 (N_1072,N_520,N_611);
nand U1073 (N_1073,N_70,N_387);
nor U1074 (N_1074,N_75,N_717);
xnor U1075 (N_1075,N_695,N_347);
and U1076 (N_1076,N_907,N_471);
xor U1077 (N_1077,N_44,N_126);
nor U1078 (N_1078,N_183,N_648);
or U1079 (N_1079,N_908,N_585);
xor U1080 (N_1080,N_914,N_781);
nor U1081 (N_1081,N_467,N_73);
xor U1082 (N_1082,N_382,N_442);
xnor U1083 (N_1083,N_693,N_144);
and U1084 (N_1084,N_478,N_287);
or U1085 (N_1085,N_510,N_338);
or U1086 (N_1086,N_207,N_771);
nand U1087 (N_1087,N_67,N_652);
xnor U1088 (N_1088,N_728,N_120);
nor U1089 (N_1089,N_887,N_741);
nor U1090 (N_1090,N_158,N_397);
or U1091 (N_1091,N_870,N_95);
xor U1092 (N_1092,N_342,N_386);
or U1093 (N_1093,N_752,N_188);
nand U1094 (N_1094,N_550,N_713);
nand U1095 (N_1095,N_751,N_526);
nand U1096 (N_1096,N_885,N_176);
nand U1097 (N_1097,N_962,N_405);
xnor U1098 (N_1098,N_195,N_61);
nand U1099 (N_1099,N_968,N_452);
nor U1100 (N_1100,N_900,N_666);
and U1101 (N_1101,N_949,N_153);
nor U1102 (N_1102,N_672,N_294);
and U1103 (N_1103,N_801,N_469);
xor U1104 (N_1104,N_187,N_849);
and U1105 (N_1105,N_639,N_353);
nor U1106 (N_1106,N_879,N_103);
nand U1107 (N_1107,N_871,N_969);
or U1108 (N_1108,N_838,N_878);
nand U1109 (N_1109,N_430,N_479);
or U1110 (N_1110,N_276,N_637);
or U1111 (N_1111,N_46,N_434);
xnor U1112 (N_1112,N_130,N_665);
nor U1113 (N_1113,N_481,N_620);
nand U1114 (N_1114,N_468,N_499);
or U1115 (N_1115,N_285,N_547);
nand U1116 (N_1116,N_307,N_464);
nand U1117 (N_1117,N_105,N_533);
xor U1118 (N_1118,N_427,N_817);
and U1119 (N_1119,N_939,N_115);
and U1120 (N_1120,N_642,N_326);
and U1121 (N_1121,N_252,N_909);
nand U1122 (N_1122,N_786,N_808);
nor U1123 (N_1123,N_162,N_263);
and U1124 (N_1124,N_560,N_348);
nand U1125 (N_1125,N_230,N_0);
and U1126 (N_1126,N_448,N_883);
nand U1127 (N_1127,N_339,N_116);
and U1128 (N_1128,N_938,N_251);
and U1129 (N_1129,N_475,N_940);
xnor U1130 (N_1130,N_554,N_623);
nand U1131 (N_1131,N_607,N_174);
xor U1132 (N_1132,N_127,N_298);
nand U1133 (N_1133,N_167,N_545);
and U1134 (N_1134,N_563,N_723);
or U1135 (N_1135,N_38,N_926);
nand U1136 (N_1136,N_221,N_833);
xnor U1137 (N_1137,N_473,N_204);
nand U1138 (N_1138,N_768,N_913);
or U1139 (N_1139,N_614,N_749);
or U1140 (N_1140,N_633,N_217);
nand U1141 (N_1141,N_155,N_435);
xor U1142 (N_1142,N_564,N_544);
nand U1143 (N_1143,N_493,N_447);
nor U1144 (N_1144,N_142,N_457);
and U1145 (N_1145,N_237,N_208);
xor U1146 (N_1146,N_858,N_690);
or U1147 (N_1147,N_476,N_591);
nand U1148 (N_1148,N_505,N_734);
nor U1149 (N_1149,N_297,N_539);
or U1150 (N_1150,N_272,N_31);
nand U1151 (N_1151,N_260,N_406);
nor U1152 (N_1152,N_111,N_536);
xnor U1153 (N_1153,N_664,N_942);
xnor U1154 (N_1154,N_681,N_843);
nor U1155 (N_1155,N_223,N_983);
nor U1156 (N_1156,N_439,N_537);
and U1157 (N_1157,N_904,N_69);
nor U1158 (N_1158,N_211,N_732);
and U1159 (N_1159,N_605,N_912);
and U1160 (N_1160,N_568,N_705);
nand U1161 (N_1161,N_726,N_718);
xnor U1162 (N_1162,N_624,N_328);
and U1163 (N_1163,N_928,N_253);
or U1164 (N_1164,N_40,N_532);
nand U1165 (N_1165,N_521,N_806);
and U1166 (N_1166,N_209,N_997);
and U1167 (N_1167,N_659,N_760);
nor U1168 (N_1168,N_222,N_407);
xor U1169 (N_1169,N_675,N_444);
nor U1170 (N_1170,N_289,N_190);
and U1171 (N_1171,N_137,N_321);
nor U1172 (N_1172,N_758,N_991);
or U1173 (N_1173,N_161,N_24);
and U1174 (N_1174,N_179,N_759);
nand U1175 (N_1175,N_774,N_361);
nand U1176 (N_1176,N_366,N_851);
xor U1177 (N_1177,N_799,N_816);
or U1178 (N_1178,N_392,N_373);
nand U1179 (N_1179,N_755,N_530);
nor U1180 (N_1180,N_138,N_597);
nand U1181 (N_1181,N_372,N_388);
nor U1182 (N_1182,N_682,N_2);
or U1183 (N_1183,N_852,N_934);
nor U1184 (N_1184,N_906,N_668);
nand U1185 (N_1185,N_350,N_68);
and U1186 (N_1186,N_163,N_4);
xor U1187 (N_1187,N_565,N_52);
nand U1188 (N_1188,N_618,N_92);
nor U1189 (N_1189,N_76,N_692);
and U1190 (N_1190,N_206,N_566);
nor U1191 (N_1191,N_853,N_164);
nand U1192 (N_1192,N_820,N_993);
nor U1193 (N_1193,N_905,N_14);
or U1194 (N_1194,N_277,N_990);
and U1195 (N_1195,N_269,N_53);
nand U1196 (N_1196,N_645,N_961);
nor U1197 (N_1197,N_863,N_177);
nor U1198 (N_1198,N_854,N_242);
nand U1199 (N_1199,N_492,N_626);
nand U1200 (N_1200,N_987,N_764);
nor U1201 (N_1201,N_440,N_199);
nand U1202 (N_1202,N_185,N_106);
nand U1203 (N_1203,N_6,N_458);
or U1204 (N_1204,N_1,N_292);
or U1205 (N_1205,N_202,N_687);
nor U1206 (N_1206,N_224,N_660);
xnor U1207 (N_1207,N_866,N_191);
nand U1208 (N_1208,N_329,N_124);
nor U1209 (N_1209,N_787,N_100);
and U1210 (N_1210,N_433,N_835);
and U1211 (N_1211,N_143,N_248);
nand U1212 (N_1212,N_139,N_123);
nand U1213 (N_1213,N_245,N_960);
xor U1214 (N_1214,N_85,N_578);
xor U1215 (N_1215,N_846,N_264);
xnor U1216 (N_1216,N_131,N_37);
and U1217 (N_1217,N_579,N_746);
or U1218 (N_1218,N_743,N_529);
xor U1219 (N_1219,N_575,N_562);
nand U1220 (N_1220,N_423,N_971);
nand U1221 (N_1221,N_876,N_792);
or U1222 (N_1222,N_656,N_194);
and U1223 (N_1223,N_671,N_337);
nor U1224 (N_1224,N_994,N_548);
nor U1225 (N_1225,N_511,N_735);
and U1226 (N_1226,N_303,N_653);
or U1227 (N_1227,N_60,N_830);
xnor U1228 (N_1228,N_625,N_600);
xnor U1229 (N_1229,N_608,N_778);
or U1230 (N_1230,N_394,N_789);
xnor U1231 (N_1231,N_518,N_389);
or U1232 (N_1232,N_21,N_632);
xnor U1233 (N_1233,N_703,N_523);
and U1234 (N_1234,N_740,N_869);
nor U1235 (N_1235,N_925,N_322);
nand U1236 (N_1236,N_981,N_514);
and U1237 (N_1237,N_456,N_34);
or U1238 (N_1238,N_368,N_107);
or U1239 (N_1239,N_313,N_945);
or U1240 (N_1240,N_815,N_832);
nand U1241 (N_1241,N_11,N_496);
nor U1242 (N_1242,N_483,N_791);
or U1243 (N_1243,N_974,N_159);
xnor U1244 (N_1244,N_947,N_56);
or U1245 (N_1245,N_170,N_23);
nor U1246 (N_1246,N_254,N_121);
nor U1247 (N_1247,N_923,N_708);
or U1248 (N_1248,N_655,N_9);
nor U1249 (N_1249,N_482,N_766);
or U1250 (N_1250,N_609,N_965);
and U1251 (N_1251,N_490,N_18);
xnor U1252 (N_1252,N_739,N_459);
or U1253 (N_1253,N_216,N_573);
xnor U1254 (N_1254,N_963,N_426);
xor U1255 (N_1255,N_501,N_450);
nand U1256 (N_1256,N_762,N_844);
nor U1257 (N_1257,N_720,N_474);
nor U1258 (N_1258,N_958,N_437);
nand U1259 (N_1259,N_873,N_979);
xnor U1260 (N_1260,N_888,N_610);
and U1261 (N_1261,N_714,N_857);
nand U1262 (N_1262,N_429,N_650);
xor U1263 (N_1263,N_494,N_954);
nand U1264 (N_1264,N_491,N_924);
xor U1265 (N_1265,N_982,N_193);
nand U1266 (N_1266,N_310,N_779);
or U1267 (N_1267,N_323,N_265);
xnor U1268 (N_1268,N_343,N_267);
nand U1269 (N_1269,N_346,N_3);
nor U1270 (N_1270,N_157,N_419);
nand U1271 (N_1271,N_438,N_553);
and U1272 (N_1272,N_229,N_569);
nor U1273 (N_1273,N_72,N_635);
and U1274 (N_1274,N_362,N_83);
xor U1275 (N_1275,N_576,N_89);
and U1276 (N_1276,N_654,N_880);
or U1277 (N_1277,N_462,N_54);
nor U1278 (N_1278,N_186,N_996);
nand U1279 (N_1279,N_445,N_29);
nor U1280 (N_1280,N_102,N_96);
nand U1281 (N_1281,N_946,N_704);
nor U1282 (N_1282,N_950,N_278);
or U1283 (N_1283,N_451,N_598);
or U1284 (N_1284,N_619,N_783);
and U1285 (N_1285,N_577,N_848);
xnor U1286 (N_1286,N_203,N_821);
or U1287 (N_1287,N_354,N_10);
and U1288 (N_1288,N_358,N_955);
and U1289 (N_1289,N_320,N_998);
xnor U1290 (N_1290,N_978,N_227);
nand U1291 (N_1291,N_541,N_99);
and U1292 (N_1292,N_151,N_315);
nand U1293 (N_1293,N_859,N_108);
or U1294 (N_1294,N_570,N_812);
xor U1295 (N_1295,N_270,N_17);
xor U1296 (N_1296,N_839,N_937);
or U1297 (N_1297,N_381,N_894);
xnor U1298 (N_1298,N_91,N_80);
xor U1299 (N_1299,N_882,N_365);
nand U1300 (N_1300,N_449,N_134);
or U1301 (N_1301,N_288,N_363);
xnor U1302 (N_1302,N_291,N_148);
nand U1303 (N_1303,N_30,N_884);
or U1304 (N_1304,N_233,N_948);
nand U1305 (N_1305,N_486,N_398);
or U1306 (N_1306,N_377,N_513);
nand U1307 (N_1307,N_622,N_644);
or U1308 (N_1308,N_275,N_404);
or U1309 (N_1309,N_841,N_259);
nor U1310 (N_1310,N_65,N_255);
nand U1311 (N_1311,N_178,N_561);
or U1312 (N_1312,N_399,N_931);
nand U1313 (N_1313,N_35,N_110);
and U1314 (N_1314,N_572,N_543);
nor U1315 (N_1315,N_87,N_385);
nand U1316 (N_1316,N_722,N_122);
or U1317 (N_1317,N_711,N_141);
or U1318 (N_1318,N_615,N_916);
or U1319 (N_1319,N_43,N_82);
nand U1320 (N_1320,N_985,N_582);
nor U1321 (N_1321,N_785,N_90);
and U1322 (N_1322,N_243,N_408);
xor U1323 (N_1323,N_875,N_104);
nand U1324 (N_1324,N_244,N_706);
nand U1325 (N_1325,N_351,N_729);
xor U1326 (N_1326,N_861,N_59);
xnor U1327 (N_1327,N_736,N_274);
and U1328 (N_1328,N_788,N_865);
nor U1329 (N_1329,N_249,N_66);
nand U1330 (N_1330,N_795,N_247);
nand U1331 (N_1331,N_767,N_301);
xnor U1332 (N_1332,N_688,N_825);
nor U1333 (N_1333,N_515,N_129);
xnor U1334 (N_1334,N_94,N_972);
xnor U1335 (N_1335,N_638,N_7);
nand U1336 (N_1336,N_813,N_213);
xnor U1337 (N_1337,N_15,N_527);
xor U1338 (N_1338,N_944,N_200);
or U1339 (N_1339,N_992,N_311);
nand U1340 (N_1340,N_383,N_454);
xnor U1341 (N_1341,N_390,N_145);
nor U1342 (N_1342,N_240,N_593);
nand U1343 (N_1343,N_304,N_929);
nand U1344 (N_1344,N_556,N_847);
nand U1345 (N_1345,N_596,N_836);
nand U1346 (N_1346,N_431,N_268);
and U1347 (N_1347,N_136,N_500);
nand U1348 (N_1348,N_160,N_412);
and U1349 (N_1349,N_919,N_943);
or U1350 (N_1350,N_150,N_794);
nand U1351 (N_1351,N_503,N_50);
xor U1352 (N_1352,N_790,N_828);
nand U1353 (N_1353,N_733,N_895);
or U1354 (N_1354,N_32,N_742);
or U1355 (N_1355,N_333,N_551);
xor U1356 (N_1356,N_970,N_48);
nor U1357 (N_1357,N_201,N_256);
xor U1358 (N_1358,N_55,N_867);
nor U1359 (N_1359,N_330,N_415);
or U1360 (N_1360,N_261,N_809);
and U1361 (N_1361,N_461,N_699);
or U1362 (N_1362,N_775,N_679);
xor U1363 (N_1363,N_640,N_701);
or U1364 (N_1364,N_702,N_721);
nor U1365 (N_1365,N_903,N_959);
xnor U1366 (N_1366,N_113,N_421);
nor U1367 (N_1367,N_805,N_364);
nand U1368 (N_1368,N_552,N_966);
nand U1369 (N_1369,N_84,N_234);
xor U1370 (N_1370,N_16,N_761);
and U1371 (N_1371,N_446,N_522);
xnor U1372 (N_1372,N_495,N_953);
nand U1373 (N_1373,N_856,N_97);
and U1374 (N_1374,N_694,N_860);
xnor U1375 (N_1375,N_472,N_81);
nand U1376 (N_1376,N_402,N_332);
xor U1377 (N_1377,N_356,N_409);
xnor U1378 (N_1378,N_542,N_899);
or U1379 (N_1379,N_26,N_920);
nor U1380 (N_1380,N_868,N_862);
xnor U1381 (N_1381,N_51,N_842);
xnor U1382 (N_1382,N_355,N_344);
nand U1383 (N_1383,N_181,N_975);
and U1384 (N_1384,N_824,N_840);
or U1385 (N_1385,N_709,N_374);
or U1386 (N_1386,N_169,N_417);
xnor U1387 (N_1387,N_88,N_58);
or U1388 (N_1388,N_508,N_205);
or U1389 (N_1389,N_441,N_683);
nor U1390 (N_1390,N_258,N_874);
or U1391 (N_1391,N_410,N_700);
or U1392 (N_1392,N_765,N_228);
and U1393 (N_1393,N_917,N_538);
xor U1394 (N_1394,N_119,N_727);
or U1395 (N_1395,N_750,N_45);
or U1396 (N_1396,N_855,N_922);
xnor U1397 (N_1397,N_658,N_524);
and U1398 (N_1398,N_540,N_334);
nand U1399 (N_1399,N_396,N_613);
nor U1400 (N_1400,N_927,N_517);
xnor U1401 (N_1401,N_784,N_519);
nand U1402 (N_1402,N_680,N_71);
nand U1403 (N_1403,N_218,N_488);
nor U1404 (N_1404,N_641,N_754);
nor U1405 (N_1405,N_125,N_140);
nand U1406 (N_1406,N_152,N_357);
or U1407 (N_1407,N_403,N_308);
nor U1408 (N_1408,N_580,N_28);
nor U1409 (N_1409,N_370,N_189);
and U1410 (N_1410,N_967,N_898);
xor U1411 (N_1411,N_306,N_336);
nand U1412 (N_1412,N_636,N_175);
nor U1413 (N_1413,N_555,N_226);
nand U1414 (N_1414,N_420,N_995);
or U1415 (N_1415,N_583,N_477);
nand U1416 (N_1416,N_379,N_312);
xnor U1417 (N_1417,N_901,N_375);
or U1418 (N_1418,N_165,N_425);
nand U1419 (N_1419,N_557,N_367);
nand U1420 (N_1420,N_369,N_309);
and U1421 (N_1421,N_198,N_684);
nand U1422 (N_1422,N_466,N_210);
or U1423 (N_1423,N_257,N_601);
nand U1424 (N_1424,N_36,N_271);
nor U1425 (N_1425,N_973,N_818);
nor U1426 (N_1426,N_246,N_414);
xor U1427 (N_1427,N_64,N_559);
nor U1428 (N_1428,N_279,N_822);
nor U1429 (N_1429,N_327,N_41);
nand U1430 (N_1430,N_872,N_319);
or U1431 (N_1431,N_400,N_989);
and U1432 (N_1432,N_696,N_497);
nand U1433 (N_1433,N_214,N_617);
and U1434 (N_1434,N_586,N_819);
xnor U1435 (N_1435,N_893,N_77);
nor U1436 (N_1436,N_918,N_756);
xor U1437 (N_1437,N_416,N_485);
xnor U1438 (N_1438,N_250,N_93);
nor U1439 (N_1439,N_512,N_811);
or U1440 (N_1440,N_484,N_74);
nor U1441 (N_1441,N_411,N_239);
xnor U1442 (N_1442,N_663,N_192);
or U1443 (N_1443,N_182,N_39);
nor U1444 (N_1444,N_324,N_798);
xnor U1445 (N_1445,N_432,N_460);
nand U1446 (N_1446,N_935,N_428);
nor U1447 (N_1447,N_941,N_212);
or U1448 (N_1448,N_604,N_42);
nand U1449 (N_1449,N_738,N_168);
xor U1450 (N_1450,N_710,N_891);
or U1451 (N_1451,N_528,N_930);
or U1452 (N_1452,N_782,N_401);
or U1453 (N_1453,N_98,N_5);
nand U1454 (N_1454,N_262,N_719);
and U1455 (N_1455,N_649,N_657);
or U1456 (N_1456,N_283,N_745);
or U1457 (N_1457,N_628,N_932);
and U1458 (N_1458,N_184,N_296);
nand U1459 (N_1459,N_220,N_117);
nor U1460 (N_1460,N_133,N_463);
nor U1461 (N_1461,N_531,N_964);
nand U1462 (N_1462,N_236,N_725);
or U1463 (N_1463,N_235,N_595);
and U1464 (N_1464,N_744,N_12);
or U1465 (N_1465,N_280,N_634);
nor U1466 (N_1466,N_341,N_986);
and U1467 (N_1467,N_814,N_612);
xnor U1468 (N_1468,N_589,N_921);
or U1469 (N_1469,N_707,N_295);
nand U1470 (N_1470,N_241,N_173);
nand U1471 (N_1471,N_302,N_630);
xnor U1472 (N_1472,N_282,N_715);
nor U1473 (N_1473,N_384,N_724);
nand U1474 (N_1474,N_225,N_933);
and U1475 (N_1475,N_436,N_507);
xnor U1476 (N_1476,N_535,N_780);
nor U1477 (N_1477,N_976,N_581);
and U1478 (N_1478,N_317,N_525);
or U1479 (N_1479,N_78,N_378);
nand U1480 (N_1480,N_890,N_8);
and U1481 (N_1481,N_114,N_22);
and U1482 (N_1482,N_673,N_480);
nand U1483 (N_1483,N_686,N_62);
xor U1484 (N_1484,N_936,N_716);
nand U1485 (N_1485,N_443,N_892);
nand U1486 (N_1486,N_487,N_393);
xnor U1487 (N_1487,N_592,N_231);
nor U1488 (N_1488,N_359,N_196);
nor U1489 (N_1489,N_118,N_57);
or U1490 (N_1490,N_902,N_20);
nand U1491 (N_1491,N_180,N_335);
nor U1492 (N_1492,N_670,N_534);
nor U1493 (N_1493,N_549,N_737);
xor U1494 (N_1494,N_915,N_747);
nor U1495 (N_1495,N_305,N_793);
or U1496 (N_1496,N_845,N_850);
nor U1497 (N_1497,N_826,N_132);
xnor U1498 (N_1498,N_977,N_345);
nand U1499 (N_1499,N_325,N_697);
nor U1500 (N_1500,N_995,N_970);
xnor U1501 (N_1501,N_955,N_450);
nand U1502 (N_1502,N_87,N_803);
nor U1503 (N_1503,N_483,N_853);
or U1504 (N_1504,N_144,N_125);
or U1505 (N_1505,N_833,N_779);
nand U1506 (N_1506,N_247,N_348);
nand U1507 (N_1507,N_901,N_79);
nor U1508 (N_1508,N_357,N_842);
and U1509 (N_1509,N_704,N_37);
or U1510 (N_1510,N_341,N_568);
nor U1511 (N_1511,N_528,N_123);
nor U1512 (N_1512,N_853,N_894);
or U1513 (N_1513,N_250,N_500);
or U1514 (N_1514,N_573,N_467);
and U1515 (N_1515,N_889,N_116);
nand U1516 (N_1516,N_232,N_264);
nor U1517 (N_1517,N_38,N_170);
or U1518 (N_1518,N_397,N_913);
or U1519 (N_1519,N_80,N_301);
nand U1520 (N_1520,N_784,N_596);
or U1521 (N_1521,N_290,N_250);
or U1522 (N_1522,N_340,N_187);
or U1523 (N_1523,N_836,N_613);
and U1524 (N_1524,N_283,N_380);
nor U1525 (N_1525,N_687,N_937);
xnor U1526 (N_1526,N_638,N_585);
and U1527 (N_1527,N_807,N_982);
and U1528 (N_1528,N_384,N_646);
nor U1529 (N_1529,N_418,N_74);
or U1530 (N_1530,N_456,N_489);
nand U1531 (N_1531,N_249,N_383);
or U1532 (N_1532,N_771,N_942);
xnor U1533 (N_1533,N_137,N_234);
nand U1534 (N_1534,N_188,N_608);
xnor U1535 (N_1535,N_603,N_989);
nand U1536 (N_1536,N_935,N_117);
and U1537 (N_1537,N_927,N_987);
nand U1538 (N_1538,N_448,N_514);
nand U1539 (N_1539,N_685,N_309);
nand U1540 (N_1540,N_358,N_727);
or U1541 (N_1541,N_139,N_19);
nand U1542 (N_1542,N_79,N_401);
or U1543 (N_1543,N_267,N_214);
or U1544 (N_1544,N_848,N_892);
and U1545 (N_1545,N_355,N_374);
nand U1546 (N_1546,N_928,N_614);
and U1547 (N_1547,N_115,N_937);
xor U1548 (N_1548,N_896,N_254);
or U1549 (N_1549,N_615,N_120);
nor U1550 (N_1550,N_181,N_437);
nand U1551 (N_1551,N_803,N_344);
or U1552 (N_1552,N_194,N_143);
nand U1553 (N_1553,N_188,N_22);
xor U1554 (N_1554,N_862,N_780);
nand U1555 (N_1555,N_588,N_706);
nand U1556 (N_1556,N_919,N_671);
or U1557 (N_1557,N_64,N_951);
and U1558 (N_1558,N_749,N_99);
nand U1559 (N_1559,N_33,N_477);
nor U1560 (N_1560,N_658,N_976);
and U1561 (N_1561,N_342,N_894);
nand U1562 (N_1562,N_638,N_265);
xor U1563 (N_1563,N_548,N_388);
nand U1564 (N_1564,N_807,N_273);
xnor U1565 (N_1565,N_121,N_778);
nand U1566 (N_1566,N_44,N_866);
and U1567 (N_1567,N_461,N_194);
or U1568 (N_1568,N_521,N_832);
xnor U1569 (N_1569,N_335,N_114);
xor U1570 (N_1570,N_555,N_5);
or U1571 (N_1571,N_676,N_246);
nor U1572 (N_1572,N_921,N_209);
nand U1573 (N_1573,N_198,N_391);
nor U1574 (N_1574,N_260,N_589);
nand U1575 (N_1575,N_711,N_56);
nor U1576 (N_1576,N_174,N_9);
xnor U1577 (N_1577,N_367,N_943);
nor U1578 (N_1578,N_262,N_197);
or U1579 (N_1579,N_477,N_993);
xnor U1580 (N_1580,N_902,N_574);
nand U1581 (N_1581,N_781,N_978);
xor U1582 (N_1582,N_357,N_754);
nor U1583 (N_1583,N_986,N_220);
xor U1584 (N_1584,N_856,N_312);
and U1585 (N_1585,N_557,N_629);
nor U1586 (N_1586,N_548,N_978);
or U1587 (N_1587,N_540,N_992);
and U1588 (N_1588,N_355,N_815);
xnor U1589 (N_1589,N_718,N_132);
nand U1590 (N_1590,N_378,N_315);
xnor U1591 (N_1591,N_429,N_943);
and U1592 (N_1592,N_406,N_717);
and U1593 (N_1593,N_250,N_307);
and U1594 (N_1594,N_853,N_328);
and U1595 (N_1595,N_949,N_264);
nand U1596 (N_1596,N_198,N_649);
nand U1597 (N_1597,N_385,N_818);
and U1598 (N_1598,N_375,N_663);
nor U1599 (N_1599,N_332,N_878);
or U1600 (N_1600,N_978,N_911);
xnor U1601 (N_1601,N_699,N_837);
xor U1602 (N_1602,N_117,N_721);
nand U1603 (N_1603,N_637,N_978);
and U1604 (N_1604,N_806,N_224);
xor U1605 (N_1605,N_251,N_426);
nor U1606 (N_1606,N_508,N_96);
or U1607 (N_1607,N_79,N_436);
nand U1608 (N_1608,N_467,N_268);
or U1609 (N_1609,N_1,N_854);
nand U1610 (N_1610,N_688,N_423);
or U1611 (N_1611,N_296,N_277);
or U1612 (N_1612,N_213,N_281);
and U1613 (N_1613,N_250,N_188);
xor U1614 (N_1614,N_889,N_22);
nor U1615 (N_1615,N_639,N_187);
xor U1616 (N_1616,N_515,N_43);
xor U1617 (N_1617,N_591,N_513);
or U1618 (N_1618,N_638,N_262);
xor U1619 (N_1619,N_477,N_890);
nor U1620 (N_1620,N_884,N_678);
or U1621 (N_1621,N_972,N_691);
nor U1622 (N_1622,N_449,N_527);
nor U1623 (N_1623,N_313,N_147);
and U1624 (N_1624,N_491,N_979);
or U1625 (N_1625,N_308,N_365);
xor U1626 (N_1626,N_203,N_918);
nor U1627 (N_1627,N_868,N_419);
nor U1628 (N_1628,N_37,N_676);
or U1629 (N_1629,N_336,N_161);
xnor U1630 (N_1630,N_234,N_898);
nor U1631 (N_1631,N_746,N_168);
nand U1632 (N_1632,N_405,N_653);
and U1633 (N_1633,N_443,N_342);
and U1634 (N_1634,N_320,N_131);
xnor U1635 (N_1635,N_202,N_185);
and U1636 (N_1636,N_709,N_354);
nand U1637 (N_1637,N_871,N_767);
xnor U1638 (N_1638,N_467,N_641);
nand U1639 (N_1639,N_406,N_66);
nand U1640 (N_1640,N_138,N_754);
xor U1641 (N_1641,N_660,N_784);
nor U1642 (N_1642,N_191,N_506);
nand U1643 (N_1643,N_228,N_449);
nor U1644 (N_1644,N_479,N_253);
nand U1645 (N_1645,N_7,N_369);
or U1646 (N_1646,N_650,N_738);
and U1647 (N_1647,N_703,N_932);
xor U1648 (N_1648,N_122,N_530);
nor U1649 (N_1649,N_684,N_385);
xor U1650 (N_1650,N_798,N_113);
nand U1651 (N_1651,N_643,N_907);
xnor U1652 (N_1652,N_66,N_499);
or U1653 (N_1653,N_568,N_269);
or U1654 (N_1654,N_30,N_432);
and U1655 (N_1655,N_726,N_503);
nand U1656 (N_1656,N_435,N_125);
and U1657 (N_1657,N_655,N_894);
nand U1658 (N_1658,N_506,N_950);
xor U1659 (N_1659,N_492,N_577);
xor U1660 (N_1660,N_40,N_0);
nand U1661 (N_1661,N_369,N_172);
or U1662 (N_1662,N_689,N_71);
and U1663 (N_1663,N_952,N_649);
nor U1664 (N_1664,N_838,N_440);
or U1665 (N_1665,N_610,N_197);
and U1666 (N_1666,N_241,N_201);
and U1667 (N_1667,N_997,N_66);
and U1668 (N_1668,N_822,N_921);
nor U1669 (N_1669,N_797,N_475);
nand U1670 (N_1670,N_720,N_767);
nand U1671 (N_1671,N_838,N_365);
and U1672 (N_1672,N_316,N_417);
nand U1673 (N_1673,N_368,N_546);
nor U1674 (N_1674,N_715,N_994);
nor U1675 (N_1675,N_788,N_235);
xnor U1676 (N_1676,N_760,N_831);
xor U1677 (N_1677,N_585,N_157);
and U1678 (N_1678,N_507,N_678);
nor U1679 (N_1679,N_130,N_378);
nand U1680 (N_1680,N_134,N_229);
and U1681 (N_1681,N_439,N_333);
or U1682 (N_1682,N_565,N_963);
nand U1683 (N_1683,N_866,N_644);
or U1684 (N_1684,N_67,N_27);
and U1685 (N_1685,N_543,N_31);
xnor U1686 (N_1686,N_521,N_674);
nor U1687 (N_1687,N_738,N_259);
and U1688 (N_1688,N_692,N_717);
nand U1689 (N_1689,N_757,N_980);
xnor U1690 (N_1690,N_623,N_109);
and U1691 (N_1691,N_308,N_740);
nand U1692 (N_1692,N_83,N_113);
and U1693 (N_1693,N_342,N_844);
or U1694 (N_1694,N_822,N_810);
xnor U1695 (N_1695,N_581,N_865);
and U1696 (N_1696,N_991,N_839);
nand U1697 (N_1697,N_274,N_575);
nand U1698 (N_1698,N_17,N_890);
nor U1699 (N_1699,N_842,N_35);
xnor U1700 (N_1700,N_489,N_123);
nand U1701 (N_1701,N_83,N_892);
and U1702 (N_1702,N_588,N_897);
xnor U1703 (N_1703,N_272,N_109);
nor U1704 (N_1704,N_255,N_492);
and U1705 (N_1705,N_375,N_272);
nor U1706 (N_1706,N_916,N_469);
nand U1707 (N_1707,N_548,N_462);
and U1708 (N_1708,N_532,N_35);
nand U1709 (N_1709,N_940,N_135);
nor U1710 (N_1710,N_788,N_67);
nor U1711 (N_1711,N_621,N_493);
or U1712 (N_1712,N_674,N_428);
and U1713 (N_1713,N_879,N_451);
xnor U1714 (N_1714,N_966,N_152);
nor U1715 (N_1715,N_159,N_990);
nand U1716 (N_1716,N_665,N_475);
nand U1717 (N_1717,N_546,N_782);
or U1718 (N_1718,N_65,N_383);
nor U1719 (N_1719,N_580,N_100);
nand U1720 (N_1720,N_363,N_520);
and U1721 (N_1721,N_409,N_544);
xnor U1722 (N_1722,N_759,N_185);
nand U1723 (N_1723,N_833,N_645);
nor U1724 (N_1724,N_419,N_897);
or U1725 (N_1725,N_739,N_471);
xor U1726 (N_1726,N_465,N_503);
nor U1727 (N_1727,N_201,N_582);
and U1728 (N_1728,N_711,N_334);
and U1729 (N_1729,N_788,N_997);
nor U1730 (N_1730,N_378,N_55);
and U1731 (N_1731,N_750,N_249);
nand U1732 (N_1732,N_66,N_218);
xor U1733 (N_1733,N_442,N_461);
and U1734 (N_1734,N_282,N_776);
or U1735 (N_1735,N_634,N_844);
or U1736 (N_1736,N_126,N_68);
nand U1737 (N_1737,N_186,N_108);
xor U1738 (N_1738,N_712,N_585);
or U1739 (N_1739,N_587,N_904);
xor U1740 (N_1740,N_544,N_597);
or U1741 (N_1741,N_533,N_207);
nor U1742 (N_1742,N_966,N_100);
and U1743 (N_1743,N_180,N_534);
nand U1744 (N_1744,N_803,N_5);
and U1745 (N_1745,N_455,N_927);
or U1746 (N_1746,N_370,N_802);
or U1747 (N_1747,N_537,N_347);
xnor U1748 (N_1748,N_810,N_958);
and U1749 (N_1749,N_847,N_867);
nor U1750 (N_1750,N_481,N_243);
nor U1751 (N_1751,N_846,N_380);
xnor U1752 (N_1752,N_174,N_591);
and U1753 (N_1753,N_111,N_463);
nor U1754 (N_1754,N_106,N_854);
xor U1755 (N_1755,N_113,N_97);
and U1756 (N_1756,N_592,N_816);
nor U1757 (N_1757,N_300,N_642);
nor U1758 (N_1758,N_752,N_901);
nor U1759 (N_1759,N_928,N_952);
or U1760 (N_1760,N_677,N_350);
and U1761 (N_1761,N_960,N_669);
and U1762 (N_1762,N_958,N_693);
nand U1763 (N_1763,N_0,N_454);
xnor U1764 (N_1764,N_0,N_961);
nor U1765 (N_1765,N_911,N_939);
nand U1766 (N_1766,N_76,N_482);
and U1767 (N_1767,N_960,N_726);
xor U1768 (N_1768,N_19,N_981);
or U1769 (N_1769,N_399,N_592);
and U1770 (N_1770,N_500,N_969);
nand U1771 (N_1771,N_292,N_255);
nand U1772 (N_1772,N_85,N_70);
nor U1773 (N_1773,N_397,N_80);
and U1774 (N_1774,N_798,N_819);
xnor U1775 (N_1775,N_980,N_153);
xor U1776 (N_1776,N_16,N_57);
nand U1777 (N_1777,N_427,N_882);
nor U1778 (N_1778,N_59,N_517);
or U1779 (N_1779,N_694,N_555);
nand U1780 (N_1780,N_52,N_919);
nor U1781 (N_1781,N_888,N_22);
and U1782 (N_1782,N_914,N_509);
nand U1783 (N_1783,N_807,N_959);
xor U1784 (N_1784,N_447,N_376);
or U1785 (N_1785,N_169,N_234);
xor U1786 (N_1786,N_514,N_584);
xor U1787 (N_1787,N_412,N_645);
nor U1788 (N_1788,N_714,N_337);
xnor U1789 (N_1789,N_386,N_717);
and U1790 (N_1790,N_40,N_613);
nor U1791 (N_1791,N_615,N_858);
xor U1792 (N_1792,N_946,N_451);
xor U1793 (N_1793,N_349,N_976);
nor U1794 (N_1794,N_945,N_120);
xor U1795 (N_1795,N_130,N_543);
or U1796 (N_1796,N_230,N_881);
nand U1797 (N_1797,N_97,N_995);
nand U1798 (N_1798,N_583,N_447);
nand U1799 (N_1799,N_764,N_776);
and U1800 (N_1800,N_150,N_821);
and U1801 (N_1801,N_135,N_140);
nand U1802 (N_1802,N_168,N_204);
xnor U1803 (N_1803,N_622,N_716);
nor U1804 (N_1804,N_221,N_650);
xor U1805 (N_1805,N_864,N_28);
nor U1806 (N_1806,N_843,N_855);
or U1807 (N_1807,N_494,N_796);
and U1808 (N_1808,N_829,N_281);
and U1809 (N_1809,N_318,N_568);
nand U1810 (N_1810,N_287,N_279);
or U1811 (N_1811,N_573,N_910);
nand U1812 (N_1812,N_504,N_922);
xor U1813 (N_1813,N_532,N_626);
or U1814 (N_1814,N_985,N_293);
nand U1815 (N_1815,N_279,N_286);
nand U1816 (N_1816,N_285,N_842);
xor U1817 (N_1817,N_166,N_174);
xnor U1818 (N_1818,N_112,N_849);
nand U1819 (N_1819,N_925,N_664);
nor U1820 (N_1820,N_44,N_860);
nand U1821 (N_1821,N_955,N_908);
nor U1822 (N_1822,N_703,N_58);
xnor U1823 (N_1823,N_52,N_966);
nor U1824 (N_1824,N_743,N_755);
xnor U1825 (N_1825,N_179,N_82);
or U1826 (N_1826,N_897,N_539);
or U1827 (N_1827,N_555,N_858);
or U1828 (N_1828,N_387,N_248);
and U1829 (N_1829,N_29,N_774);
nor U1830 (N_1830,N_239,N_478);
and U1831 (N_1831,N_557,N_296);
or U1832 (N_1832,N_65,N_720);
or U1833 (N_1833,N_638,N_795);
nand U1834 (N_1834,N_302,N_547);
or U1835 (N_1835,N_237,N_856);
or U1836 (N_1836,N_677,N_262);
xor U1837 (N_1837,N_297,N_634);
xor U1838 (N_1838,N_62,N_510);
and U1839 (N_1839,N_327,N_471);
nor U1840 (N_1840,N_36,N_264);
or U1841 (N_1841,N_603,N_561);
nor U1842 (N_1842,N_493,N_676);
xor U1843 (N_1843,N_163,N_151);
or U1844 (N_1844,N_777,N_829);
xnor U1845 (N_1845,N_902,N_626);
xnor U1846 (N_1846,N_16,N_854);
or U1847 (N_1847,N_289,N_636);
or U1848 (N_1848,N_603,N_440);
xor U1849 (N_1849,N_515,N_493);
and U1850 (N_1850,N_896,N_299);
nor U1851 (N_1851,N_449,N_254);
or U1852 (N_1852,N_173,N_622);
xor U1853 (N_1853,N_811,N_165);
nor U1854 (N_1854,N_185,N_812);
and U1855 (N_1855,N_721,N_511);
or U1856 (N_1856,N_502,N_938);
xnor U1857 (N_1857,N_631,N_12);
or U1858 (N_1858,N_429,N_415);
nand U1859 (N_1859,N_157,N_275);
nand U1860 (N_1860,N_84,N_20);
nor U1861 (N_1861,N_928,N_991);
xor U1862 (N_1862,N_473,N_240);
xnor U1863 (N_1863,N_435,N_407);
nor U1864 (N_1864,N_818,N_845);
or U1865 (N_1865,N_559,N_295);
or U1866 (N_1866,N_524,N_120);
nor U1867 (N_1867,N_560,N_259);
nor U1868 (N_1868,N_526,N_200);
and U1869 (N_1869,N_467,N_28);
nand U1870 (N_1870,N_693,N_39);
nand U1871 (N_1871,N_295,N_883);
xor U1872 (N_1872,N_485,N_291);
and U1873 (N_1873,N_155,N_734);
xor U1874 (N_1874,N_528,N_263);
or U1875 (N_1875,N_604,N_806);
or U1876 (N_1876,N_532,N_977);
nand U1877 (N_1877,N_927,N_967);
nor U1878 (N_1878,N_857,N_158);
xnor U1879 (N_1879,N_810,N_827);
and U1880 (N_1880,N_79,N_808);
and U1881 (N_1881,N_424,N_912);
nor U1882 (N_1882,N_515,N_542);
nor U1883 (N_1883,N_377,N_704);
or U1884 (N_1884,N_89,N_177);
and U1885 (N_1885,N_42,N_560);
xnor U1886 (N_1886,N_539,N_446);
nor U1887 (N_1887,N_996,N_560);
or U1888 (N_1888,N_620,N_409);
or U1889 (N_1889,N_292,N_796);
and U1890 (N_1890,N_634,N_36);
nor U1891 (N_1891,N_823,N_3);
and U1892 (N_1892,N_991,N_703);
or U1893 (N_1893,N_341,N_788);
and U1894 (N_1894,N_511,N_109);
nand U1895 (N_1895,N_611,N_801);
nand U1896 (N_1896,N_825,N_452);
and U1897 (N_1897,N_587,N_939);
and U1898 (N_1898,N_92,N_601);
xor U1899 (N_1899,N_37,N_144);
and U1900 (N_1900,N_225,N_811);
nand U1901 (N_1901,N_662,N_864);
and U1902 (N_1902,N_316,N_71);
nand U1903 (N_1903,N_966,N_168);
xor U1904 (N_1904,N_614,N_501);
or U1905 (N_1905,N_196,N_60);
nand U1906 (N_1906,N_61,N_901);
or U1907 (N_1907,N_825,N_111);
and U1908 (N_1908,N_338,N_998);
and U1909 (N_1909,N_544,N_366);
or U1910 (N_1910,N_757,N_558);
or U1911 (N_1911,N_60,N_434);
nand U1912 (N_1912,N_589,N_152);
xnor U1913 (N_1913,N_521,N_309);
xor U1914 (N_1914,N_707,N_771);
nor U1915 (N_1915,N_384,N_185);
and U1916 (N_1916,N_903,N_636);
xor U1917 (N_1917,N_20,N_181);
nor U1918 (N_1918,N_725,N_962);
xor U1919 (N_1919,N_198,N_25);
and U1920 (N_1920,N_152,N_671);
nand U1921 (N_1921,N_23,N_407);
nand U1922 (N_1922,N_341,N_416);
and U1923 (N_1923,N_745,N_11);
nor U1924 (N_1924,N_424,N_51);
and U1925 (N_1925,N_486,N_47);
and U1926 (N_1926,N_837,N_395);
or U1927 (N_1927,N_542,N_125);
xnor U1928 (N_1928,N_655,N_868);
nor U1929 (N_1929,N_440,N_990);
and U1930 (N_1930,N_328,N_870);
and U1931 (N_1931,N_45,N_315);
xnor U1932 (N_1932,N_258,N_398);
xnor U1933 (N_1933,N_227,N_622);
xnor U1934 (N_1934,N_745,N_369);
nor U1935 (N_1935,N_807,N_425);
or U1936 (N_1936,N_921,N_755);
and U1937 (N_1937,N_185,N_430);
xor U1938 (N_1938,N_525,N_390);
nor U1939 (N_1939,N_188,N_194);
nand U1940 (N_1940,N_130,N_728);
and U1941 (N_1941,N_626,N_68);
xnor U1942 (N_1942,N_319,N_533);
and U1943 (N_1943,N_408,N_385);
xor U1944 (N_1944,N_711,N_123);
nor U1945 (N_1945,N_623,N_169);
nor U1946 (N_1946,N_913,N_322);
nand U1947 (N_1947,N_409,N_99);
and U1948 (N_1948,N_353,N_915);
xor U1949 (N_1949,N_428,N_404);
or U1950 (N_1950,N_160,N_732);
or U1951 (N_1951,N_264,N_766);
nand U1952 (N_1952,N_895,N_503);
and U1953 (N_1953,N_260,N_255);
nand U1954 (N_1954,N_533,N_516);
or U1955 (N_1955,N_143,N_696);
xnor U1956 (N_1956,N_409,N_515);
or U1957 (N_1957,N_415,N_672);
and U1958 (N_1958,N_544,N_639);
or U1959 (N_1959,N_375,N_371);
nand U1960 (N_1960,N_771,N_482);
nand U1961 (N_1961,N_308,N_423);
or U1962 (N_1962,N_522,N_168);
or U1963 (N_1963,N_87,N_699);
nand U1964 (N_1964,N_226,N_61);
xnor U1965 (N_1965,N_745,N_275);
and U1966 (N_1966,N_168,N_20);
nand U1967 (N_1967,N_382,N_67);
nor U1968 (N_1968,N_230,N_78);
nor U1969 (N_1969,N_913,N_565);
nand U1970 (N_1970,N_744,N_804);
nand U1971 (N_1971,N_178,N_142);
and U1972 (N_1972,N_40,N_798);
xnor U1973 (N_1973,N_873,N_649);
nand U1974 (N_1974,N_751,N_158);
or U1975 (N_1975,N_949,N_198);
and U1976 (N_1976,N_164,N_301);
nand U1977 (N_1977,N_563,N_713);
or U1978 (N_1978,N_983,N_430);
and U1979 (N_1979,N_564,N_579);
and U1980 (N_1980,N_428,N_315);
nor U1981 (N_1981,N_792,N_939);
and U1982 (N_1982,N_562,N_176);
nor U1983 (N_1983,N_765,N_120);
nor U1984 (N_1984,N_644,N_340);
nand U1985 (N_1985,N_505,N_729);
xnor U1986 (N_1986,N_631,N_508);
nor U1987 (N_1987,N_601,N_435);
nor U1988 (N_1988,N_540,N_616);
or U1989 (N_1989,N_278,N_934);
xnor U1990 (N_1990,N_995,N_5);
nor U1991 (N_1991,N_30,N_124);
and U1992 (N_1992,N_996,N_792);
and U1993 (N_1993,N_404,N_516);
or U1994 (N_1994,N_267,N_501);
and U1995 (N_1995,N_835,N_238);
nor U1996 (N_1996,N_272,N_588);
nor U1997 (N_1997,N_639,N_723);
or U1998 (N_1998,N_923,N_68);
nor U1999 (N_1999,N_777,N_369);
and U2000 (N_2000,N_1204,N_1142);
xnor U2001 (N_2001,N_1324,N_1735);
or U2002 (N_2002,N_1579,N_1250);
nor U2003 (N_2003,N_1108,N_1003);
nor U2004 (N_2004,N_1714,N_1738);
and U2005 (N_2005,N_1261,N_1590);
and U2006 (N_2006,N_1653,N_1781);
nor U2007 (N_2007,N_1356,N_1561);
and U2008 (N_2008,N_1752,N_1264);
nand U2009 (N_2009,N_1479,N_1919);
nor U2010 (N_2010,N_1015,N_1577);
nand U2011 (N_2011,N_1219,N_1258);
nand U2012 (N_2012,N_1410,N_1076);
nor U2013 (N_2013,N_1343,N_1423);
nand U2014 (N_2014,N_1935,N_1104);
nand U2015 (N_2015,N_1778,N_1418);
or U2016 (N_2016,N_1345,N_1080);
or U2017 (N_2017,N_1589,N_1618);
nor U2018 (N_2018,N_1969,N_1568);
nor U2019 (N_2019,N_1701,N_1117);
and U2020 (N_2020,N_1814,N_1668);
or U2021 (N_2021,N_1354,N_1475);
nor U2022 (N_2022,N_1510,N_1225);
nor U2023 (N_2023,N_1859,N_1257);
and U2024 (N_2024,N_1144,N_1646);
nor U2025 (N_2025,N_1013,N_1887);
or U2026 (N_2026,N_1968,N_1239);
or U2027 (N_2027,N_1404,N_1282);
nand U2028 (N_2028,N_1709,N_1830);
nor U2029 (N_2029,N_1988,N_1959);
and U2030 (N_2030,N_1295,N_1980);
nand U2031 (N_2031,N_1260,N_1524);
or U2032 (N_2032,N_1348,N_1827);
nand U2033 (N_2033,N_1218,N_1093);
and U2034 (N_2034,N_1737,N_1281);
nand U2035 (N_2035,N_1493,N_1385);
and U2036 (N_2036,N_1717,N_1136);
or U2037 (N_2037,N_1697,N_1694);
and U2038 (N_2038,N_1245,N_1269);
and U2039 (N_2039,N_1800,N_1110);
and U2040 (N_2040,N_1342,N_1162);
and U2041 (N_2041,N_1044,N_1555);
xnor U2042 (N_2042,N_1286,N_1329);
nand U2043 (N_2043,N_1776,N_1990);
and U2044 (N_2044,N_1622,N_1152);
xor U2045 (N_2045,N_1059,N_1374);
and U2046 (N_2046,N_1791,N_1321);
nand U2047 (N_2047,N_1472,N_1573);
nor U2048 (N_2048,N_1306,N_1840);
xnor U2049 (N_2049,N_1105,N_1462);
xnor U2050 (N_2050,N_1773,N_1716);
nor U2051 (N_2051,N_1165,N_1430);
nand U2052 (N_2052,N_1684,N_1001);
xnor U2053 (N_2053,N_1898,N_1743);
xnor U2054 (N_2054,N_1967,N_1976);
xor U2055 (N_2055,N_1772,N_1831);
nand U2056 (N_2056,N_1858,N_1055);
nand U2057 (N_2057,N_1871,N_1720);
and U2058 (N_2058,N_1227,N_1943);
xnor U2059 (N_2059,N_1503,N_1518);
nor U2060 (N_2060,N_1673,N_1276);
and U2061 (N_2061,N_1075,N_1259);
and U2062 (N_2062,N_1323,N_1900);
and U2063 (N_2063,N_1855,N_1757);
or U2064 (N_2064,N_1421,N_1965);
xor U2065 (N_2065,N_1049,N_1592);
and U2066 (N_2066,N_1955,N_1500);
xor U2067 (N_2067,N_1789,N_1336);
nand U2068 (N_2068,N_1106,N_1232);
and U2069 (N_2069,N_1740,N_1617);
and U2070 (N_2070,N_1920,N_1113);
nand U2071 (N_2071,N_1231,N_1991);
xnor U2072 (N_2072,N_1643,N_1907);
and U2073 (N_2073,N_1126,N_1726);
xnor U2074 (N_2074,N_1603,N_1009);
xnor U2075 (N_2075,N_1195,N_1798);
and U2076 (N_2076,N_1334,N_1069);
nor U2077 (N_2077,N_1065,N_1519);
nand U2078 (N_2078,N_1391,N_1077);
nand U2079 (N_2079,N_1580,N_1832);
xor U2080 (N_2080,N_1084,N_1924);
or U2081 (N_2081,N_1645,N_1368);
nand U2082 (N_2082,N_1143,N_1470);
or U2083 (N_2083,N_1608,N_1972);
or U2084 (N_2084,N_1996,N_1133);
xor U2085 (N_2085,N_1989,N_1613);
nor U2086 (N_2086,N_1026,N_1672);
xnor U2087 (N_2087,N_1983,N_1288);
xnor U2088 (N_2088,N_1880,N_1123);
nor U2089 (N_2089,N_1428,N_1605);
xor U2090 (N_2090,N_1340,N_1867);
nor U2091 (N_2091,N_1381,N_1298);
nand U2092 (N_2092,N_1889,N_1452);
or U2093 (N_2093,N_1767,N_1599);
and U2094 (N_2094,N_1395,N_1574);
nor U2095 (N_2095,N_1626,N_1252);
xnor U2096 (N_2096,N_1468,N_1857);
nand U2097 (N_2097,N_1455,N_1074);
or U2098 (N_2098,N_1971,N_1940);
nor U2099 (N_2099,N_1852,N_1928);
and U2100 (N_2100,N_1895,N_1494);
nand U2101 (N_2101,N_1770,N_1140);
nand U2102 (N_2102,N_1593,N_1861);
xnor U2103 (N_2103,N_1777,N_1205);
and U2104 (N_2104,N_1504,N_1525);
or U2105 (N_2105,N_1731,N_1432);
nand U2106 (N_2106,N_1660,N_1546);
nand U2107 (N_2107,N_1137,N_1497);
xnor U2108 (N_2108,N_1492,N_1841);
and U2109 (N_2109,N_1869,N_1487);
nand U2110 (N_2110,N_1834,N_1540);
or U2111 (N_2111,N_1248,N_1083);
and U2112 (N_2112,N_1621,N_1456);
xnor U2113 (N_2113,N_1669,N_1331);
and U2114 (N_2114,N_1333,N_1922);
nor U2115 (N_2115,N_1551,N_1936);
xnor U2116 (N_2116,N_1601,N_1196);
or U2117 (N_2117,N_1835,N_1696);
xnor U2118 (N_2118,N_1986,N_1828);
xnor U2119 (N_2119,N_1021,N_1255);
nand U2120 (N_2120,N_1139,N_1045);
xor U2121 (N_2121,N_1085,N_1893);
xnor U2122 (N_2122,N_1389,N_1058);
nor U2123 (N_2123,N_1016,N_1431);
and U2124 (N_2124,N_1199,N_1315);
xnor U2125 (N_2125,N_1240,N_1925);
or U2126 (N_2126,N_1805,N_1420);
nor U2127 (N_2127,N_1416,N_1483);
nor U2128 (N_2128,N_1208,N_1779);
xnor U2129 (N_2129,N_1018,N_1280);
xnor U2130 (N_2130,N_1485,N_1792);
xnor U2131 (N_2131,N_1775,N_1184);
and U2132 (N_2132,N_1806,N_1006);
xor U2133 (N_2133,N_1464,N_1386);
and U2134 (N_2134,N_1667,N_1350);
xor U2135 (N_2135,N_1631,N_1816);
nor U2136 (N_2136,N_1558,N_1293);
nor U2137 (N_2137,N_1289,N_1819);
nor U2138 (N_2138,N_1312,N_1103);
or U2139 (N_2139,N_1465,N_1896);
and U2140 (N_2140,N_1111,N_1553);
xor U2141 (N_2141,N_1193,N_1256);
nand U2142 (N_2142,N_1629,N_1849);
xnor U2143 (N_2143,N_1039,N_1918);
nor U2144 (N_2144,N_1228,N_1361);
or U2145 (N_2145,N_1619,N_1351);
nor U2146 (N_2146,N_1141,N_1482);
xor U2147 (N_2147,N_1437,N_1853);
and U2148 (N_2148,N_1217,N_1189);
nor U2149 (N_2149,N_1187,N_1010);
nand U2150 (N_2150,N_1092,N_1754);
and U2151 (N_2151,N_1745,N_1300);
or U2152 (N_2152,N_1222,N_1355);
nor U2153 (N_2153,N_1471,N_1422);
xnor U2154 (N_2154,N_1836,N_1839);
and U2155 (N_2155,N_1387,N_1644);
xor U2156 (N_2156,N_1678,N_1810);
nand U2157 (N_2157,N_1584,N_1096);
and U2158 (N_2158,N_1559,N_1606);
or U2159 (N_2159,N_1598,N_1870);
or U2160 (N_2160,N_1130,N_1099);
nor U2161 (N_2161,N_1607,N_1241);
nor U2162 (N_2162,N_1284,N_1657);
and U2163 (N_2163,N_1864,N_1457);
and U2164 (N_2164,N_1153,N_1164);
nand U2165 (N_2165,N_1956,N_1034);
and U2166 (N_2166,N_1949,N_1101);
and U2167 (N_2167,N_1636,N_1458);
nand U2168 (N_2168,N_1611,N_1878);
xnor U2169 (N_2169,N_1417,N_1048);
and U2170 (N_2170,N_1175,N_1314);
nor U2171 (N_2171,N_1929,N_1042);
and U2172 (N_2172,N_1888,N_1319);
nand U2173 (N_2173,N_1733,N_1424);
nor U2174 (N_2174,N_1901,N_1718);
nand U2175 (N_2175,N_1337,N_1583);
nand U2176 (N_2176,N_1275,N_1372);
nor U2177 (N_2177,N_1572,N_1002);
and U2178 (N_2178,N_1753,N_1449);
nand U2179 (N_2179,N_1713,N_1768);
and U2180 (N_2180,N_1397,N_1402);
or U2181 (N_2181,N_1650,N_1444);
xor U2182 (N_2182,N_1703,N_1405);
nor U2183 (N_2183,N_1185,N_1022);
nand U2184 (N_2184,N_1394,N_1446);
and U2185 (N_2185,N_1747,N_1512);
xor U2186 (N_2186,N_1548,N_1815);
and U2187 (N_2187,N_1438,N_1600);
or U2188 (N_2188,N_1729,N_1216);
and U2189 (N_2189,N_1169,N_1450);
and U2190 (N_2190,N_1095,N_1415);
or U2191 (N_2191,N_1427,N_1480);
xnor U2192 (N_2192,N_1066,N_1057);
xnor U2193 (N_2193,N_1310,N_1981);
nor U2194 (N_2194,N_1681,N_1547);
or U2195 (N_2195,N_1903,N_1506);
nor U2196 (N_2196,N_1535,N_1665);
or U2197 (N_2197,N_1119,N_1121);
or U2198 (N_2198,N_1127,N_1693);
xnor U2199 (N_2199,N_1296,N_1517);
and U2200 (N_2200,N_1398,N_1947);
or U2201 (N_2201,N_1937,N_1166);
or U2202 (N_2202,N_1656,N_1180);
nand U2203 (N_2203,N_1244,N_1522);
xor U2204 (N_2204,N_1545,N_1223);
xnor U2205 (N_2205,N_1429,N_1655);
xor U2206 (N_2206,N_1170,N_1291);
and U2207 (N_2207,N_1892,N_1763);
nor U2208 (N_2208,N_1272,N_1702);
xor U2209 (N_2209,N_1332,N_1197);
or U2210 (N_2210,N_1687,N_1530);
or U2211 (N_2211,N_1459,N_1771);
or U2212 (N_2212,N_1000,N_1910);
and U2213 (N_2213,N_1451,N_1439);
nand U2214 (N_2214,N_1008,N_1253);
nand U2215 (N_2215,N_1370,N_1214);
and U2216 (N_2216,N_1362,N_1237);
nand U2217 (N_2217,N_1683,N_1179);
and U2218 (N_2218,N_1191,N_1266);
and U2219 (N_2219,N_1094,N_1215);
nor U2220 (N_2220,N_1706,N_1651);
nor U2221 (N_2221,N_1705,N_1308);
xnor U2222 (N_2222,N_1749,N_1627);
nor U2223 (N_2223,N_1938,N_1043);
or U2224 (N_2224,N_1327,N_1883);
or U2225 (N_2225,N_1388,N_1612);
nand U2226 (N_2226,N_1652,N_1711);
nor U2227 (N_2227,N_1513,N_1884);
and U2228 (N_2228,N_1038,N_1198);
nor U2229 (N_2229,N_1496,N_1209);
nand U2230 (N_2230,N_1876,N_1285);
xor U2231 (N_2231,N_1671,N_1649);
nor U2232 (N_2232,N_1933,N_1030);
or U2233 (N_2233,N_1570,N_1974);
nor U2234 (N_2234,N_1495,N_1134);
nand U2235 (N_2235,N_1251,N_1109);
nand U2236 (N_2236,N_1610,N_1346);
nor U2237 (N_2237,N_1648,N_1046);
or U2238 (N_2238,N_1017,N_1766);
or U2239 (N_2239,N_1846,N_1363);
and U2240 (N_2240,N_1824,N_1279);
nor U2241 (N_2241,N_1014,N_1236);
xnor U2242 (N_2242,N_1700,N_1271);
and U2243 (N_2243,N_1614,N_1566);
nand U2244 (N_2244,N_1182,N_1862);
and U2245 (N_2245,N_1349,N_1413);
and U2246 (N_2246,N_1746,N_1131);
or U2247 (N_2247,N_1962,N_1945);
and U2248 (N_2248,N_1994,N_1913);
and U2249 (N_2249,N_1960,N_1278);
nor U2250 (N_2250,N_1263,N_1033);
or U2251 (N_2251,N_1838,N_1799);
nand U2252 (N_2252,N_1699,N_1004);
and U2253 (N_2253,N_1061,N_1514);
nand U2254 (N_2254,N_1999,N_1477);
and U2255 (N_2255,N_1082,N_1326);
or U2256 (N_2256,N_1760,N_1543);
or U2257 (N_2257,N_1533,N_1053);
or U2258 (N_2258,N_1707,N_1012);
and U2259 (N_2259,N_1313,N_1817);
xor U2260 (N_2260,N_1538,N_1081);
xnor U2261 (N_2261,N_1620,N_1554);
nor U2262 (N_2262,N_1796,N_1682);
nor U2263 (N_2263,N_1396,N_1642);
and U2264 (N_2264,N_1881,N_1982);
or U2265 (N_2265,N_1780,N_1463);
nor U2266 (N_2266,N_1750,N_1089);
nand U2267 (N_2267,N_1508,N_1739);
xnor U2268 (N_2268,N_1628,N_1845);
xor U2269 (N_2269,N_1246,N_1473);
xor U2270 (N_2270,N_1442,N_1802);
or U2271 (N_2271,N_1826,N_1877);
xor U2272 (N_2272,N_1647,N_1582);
xnor U2273 (N_2273,N_1369,N_1997);
nand U2274 (N_2274,N_1390,N_1330);
xnor U2275 (N_2275,N_1724,N_1571);
or U2276 (N_2276,N_1591,N_1978);
nand U2277 (N_2277,N_1813,N_1031);
or U2278 (N_2278,N_1915,N_1523);
nor U2279 (N_2279,N_1529,N_1676);
xor U2280 (N_2280,N_1963,N_1425);
and U2281 (N_2281,N_1207,N_1788);
xnor U2282 (N_2282,N_1863,N_1403);
nand U2283 (N_2283,N_1072,N_1818);
or U2284 (N_2284,N_1120,N_1382);
and U2285 (N_2285,N_1921,N_1984);
nor U2286 (N_2286,N_1804,N_1722);
xnor U2287 (N_2287,N_1238,N_1254);
nor U2288 (N_2288,N_1954,N_1062);
xnor U2289 (N_2289,N_1917,N_1734);
nor U2290 (N_2290,N_1393,N_1118);
nand U2291 (N_2291,N_1122,N_1079);
nand U2292 (N_2292,N_1489,N_1730);
nand U2293 (N_2293,N_1267,N_1054);
nor U2294 (N_2294,N_1380,N_1625);
and U2295 (N_2295,N_1467,N_1801);
and U2296 (N_2296,N_1578,N_1825);
xnor U2297 (N_2297,N_1499,N_1147);
nand U2298 (N_2298,N_1490,N_1563);
nand U2299 (N_2299,N_1379,N_1537);
nor U2300 (N_2300,N_1552,N_1376);
or U2301 (N_2301,N_1748,N_1661);
nor U2302 (N_2302,N_1035,N_1309);
nor U2303 (N_2303,N_1078,N_1056);
nand U2304 (N_2304,N_1872,N_1150);
and U2305 (N_2305,N_1299,N_1769);
nand U2306 (N_2306,N_1274,N_1371);
and U2307 (N_2307,N_1027,N_1615);
nand U2308 (N_2308,N_1148,N_1460);
nand U2309 (N_2309,N_1782,N_1102);
or U2310 (N_2310,N_1795,N_1624);
or U2311 (N_2311,N_1927,N_1304);
and U2312 (N_2312,N_1844,N_1604);
and U2313 (N_2313,N_1958,N_1821);
nand U2314 (N_2314,N_1865,N_1007);
and U2315 (N_2315,N_1951,N_1961);
and U2316 (N_2316,N_1744,N_1501);
nand U2317 (N_2317,N_1569,N_1235);
nand U2318 (N_2318,N_1623,N_1581);
nor U2319 (N_2319,N_1145,N_1339);
or U2320 (N_2320,N_1174,N_1411);
nor U2321 (N_2321,N_1596,N_1527);
xnor U2322 (N_2322,N_1822,N_1316);
xor U2323 (N_2323,N_1575,N_1194);
and U2324 (N_2324,N_1213,N_1037);
nor U2325 (N_2325,N_1311,N_1068);
xnor U2326 (N_2326,N_1692,N_1270);
nor U2327 (N_2327,N_1761,N_1833);
and U2328 (N_2328,N_1445,N_1112);
xor U2329 (N_2329,N_1401,N_1741);
and U2330 (N_2330,N_1930,N_1226);
xnor U2331 (N_2331,N_1891,N_1273);
and U2332 (N_2332,N_1028,N_1322);
and U2333 (N_2333,N_1923,N_1690);
nand U2334 (N_2334,N_1979,N_1902);
nand U2335 (N_2335,N_1294,N_1011);
or U2336 (N_2336,N_1436,N_1469);
xnor U2337 (N_2337,N_1146,N_1758);
xnor U2338 (N_2338,N_1177,N_1985);
nand U2339 (N_2339,N_1843,N_1481);
nor U2340 (N_2340,N_1186,N_1704);
xor U2341 (N_2341,N_1020,N_1658);
and U2342 (N_2342,N_1534,N_1942);
or U2343 (N_2343,N_1287,N_1856);
or U2344 (N_2344,N_1352,N_1125);
or U2345 (N_2345,N_1790,N_1894);
xor U2346 (N_2346,N_1905,N_1441);
or U2347 (N_2347,N_1176,N_1283);
nand U2348 (N_2348,N_1230,N_1203);
xor U2349 (N_2349,N_1560,N_1384);
nand U2350 (N_2350,N_1290,N_1762);
or U2351 (N_2351,N_1157,N_1220);
nand U2352 (N_2352,N_1190,N_1542);
and U2353 (N_2353,N_1719,N_1478);
nor U2354 (N_2354,N_1233,N_1850);
or U2355 (N_2355,N_1212,N_1520);
or U2356 (N_2356,N_1318,N_1414);
xnor U2357 (N_2357,N_1229,N_1454);
xor U2358 (N_2358,N_1156,N_1885);
or U2359 (N_2359,N_1674,N_1328);
nor U2360 (N_2360,N_1461,N_1484);
nor U2361 (N_2361,N_1515,N_1476);
nor U2362 (N_2362,N_1098,N_1783);
or U2363 (N_2363,N_1808,N_1755);
nor U2364 (N_2364,N_1637,N_1163);
xnor U2365 (N_2365,N_1114,N_1908);
nor U2366 (N_2366,N_1019,N_1353);
xnor U2367 (N_2367,N_1659,N_1842);
nor U2368 (N_2368,N_1685,N_1158);
xnor U2369 (N_2369,N_1115,N_1160);
or U2370 (N_2370,N_1129,N_1528);
xor U2371 (N_2371,N_1440,N_1025);
nand U2372 (N_2372,N_1466,N_1378);
xor U2373 (N_2373,N_1365,N_1998);
xnor U2374 (N_2374,N_1851,N_1070);
xor U2375 (N_2375,N_1434,N_1262);
xor U2376 (N_2376,N_1087,N_1521);
or U2377 (N_2377,N_1364,N_1097);
or U2378 (N_2378,N_1443,N_1809);
or U2379 (N_2379,N_1138,N_1183);
or U2380 (N_2380,N_1630,N_1221);
xor U2381 (N_2381,N_1124,N_1906);
nand U2382 (N_2382,N_1847,N_1820);
and U2383 (N_2383,N_1941,N_1234);
nand U2384 (N_2384,N_1686,N_1912);
or U2385 (N_2385,N_1970,N_1774);
and U2386 (N_2386,N_1695,N_1201);
and U2387 (N_2387,N_1609,N_1516);
and U2388 (N_2388,N_1360,N_1383);
or U2389 (N_2389,N_1531,N_1532);
xor U2390 (N_2390,N_1662,N_1210);
nor U2391 (N_2391,N_1728,N_1932);
xnor U2392 (N_2392,N_1567,N_1448);
and U2393 (N_2393,N_1151,N_1557);
nor U2394 (N_2394,N_1135,N_1873);
or U2395 (N_2395,N_1708,N_1407);
nor U2396 (N_2396,N_1751,N_1688);
or U2397 (N_2397,N_1914,N_1957);
or U2398 (N_2398,N_1488,N_1654);
xnor U2399 (N_2399,N_1100,N_1192);
and U2400 (N_2400,N_1377,N_1868);
or U2401 (N_2401,N_1172,N_1992);
or U2402 (N_2402,N_1344,N_1400);
xnor U2403 (N_2403,N_1677,N_1587);
xor U2404 (N_2404,N_1052,N_1890);
or U2405 (N_2405,N_1064,N_1073);
xor U2406 (N_2406,N_1875,N_1616);
and U2407 (N_2407,N_1866,N_1032);
or U2408 (N_2408,N_1338,N_1689);
or U2409 (N_2409,N_1181,N_1964);
and U2410 (N_2410,N_1585,N_1909);
or U2411 (N_2411,N_1944,N_1934);
xor U2412 (N_2412,N_1509,N_1409);
xor U2413 (N_2413,N_1277,N_1797);
xor U2414 (N_2414,N_1474,N_1161);
nor U2415 (N_2415,N_1811,N_1159);
nand U2416 (N_2416,N_1803,N_1785);
nor U2417 (N_2417,N_1886,N_1950);
and U2418 (N_2418,N_1498,N_1168);
and U2419 (N_2419,N_1200,N_1412);
and U2420 (N_2420,N_1948,N_1297);
and U2421 (N_2421,N_1664,N_1787);
nand U2422 (N_2422,N_1486,N_1698);
or U2423 (N_2423,N_1024,N_1023);
and U2424 (N_2424,N_1549,N_1358);
nor U2425 (N_2425,N_1036,N_1249);
xnor U2426 (N_2426,N_1544,N_1502);
nor U2427 (N_2427,N_1946,N_1224);
or U2428 (N_2428,N_1732,N_1848);
nand U2429 (N_2429,N_1564,N_1712);
and U2430 (N_2430,N_1202,N_1091);
nor U2431 (N_2431,N_1063,N_1691);
and U2432 (N_2432,N_1860,N_1511);
nor U2433 (N_2433,N_1829,N_1784);
nand U2434 (N_2434,N_1453,N_1307);
and U2435 (N_2435,N_1088,N_1206);
xor U2436 (N_2436,N_1874,N_1305);
or U2437 (N_2437,N_1562,N_1977);
or U2438 (N_2438,N_1406,N_1041);
xnor U2439 (N_2439,N_1050,N_1634);
and U2440 (N_2440,N_1742,N_1359);
nand U2441 (N_2441,N_1973,N_1786);
nand U2442 (N_2442,N_1837,N_1188);
or U2443 (N_2443,N_1897,N_1640);
nor U2444 (N_2444,N_1725,N_1357);
and U2445 (N_2445,N_1067,N_1341);
or U2446 (N_2446,N_1419,N_1303);
nor U2447 (N_2447,N_1392,N_1178);
nand U2448 (N_2448,N_1541,N_1586);
nor U2449 (N_2449,N_1426,N_1526);
xor U2450 (N_2450,N_1447,N_1715);
or U2451 (N_2451,N_1507,N_1247);
nand U2452 (N_2452,N_1107,N_1759);
xor U2453 (N_2453,N_1710,N_1047);
and U2454 (N_2454,N_1060,N_1987);
xnor U2455 (N_2455,N_1916,N_1764);
xnor U2456 (N_2456,N_1090,N_1670);
or U2457 (N_2457,N_1433,N_1325);
and U2458 (N_2458,N_1301,N_1854);
xor U2459 (N_2459,N_1211,N_1040);
nand U2460 (N_2460,N_1904,N_1071);
nor U2461 (N_2461,N_1793,N_1675);
nand U2462 (N_2462,N_1953,N_1723);
nor U2463 (N_2463,N_1505,N_1993);
xor U2464 (N_2464,N_1292,N_1679);
or U2465 (N_2465,N_1005,N_1594);
xnor U2466 (N_2466,N_1966,N_1051);
and U2467 (N_2467,N_1879,N_1939);
xnor U2468 (N_2468,N_1536,N_1242);
and U2469 (N_2469,N_1765,N_1931);
xnor U2470 (N_2470,N_1666,N_1347);
xor U2471 (N_2471,N_1632,N_1171);
or U2472 (N_2472,N_1756,N_1911);
xor U2473 (N_2473,N_1320,N_1995);
nand U2474 (N_2474,N_1243,N_1029);
and U2475 (N_2475,N_1408,N_1154);
xnor U2476 (N_2476,N_1155,N_1952);
xor U2477 (N_2477,N_1132,N_1975);
nor U2478 (N_2478,N_1823,N_1794);
or U2479 (N_2479,N_1149,N_1727);
nor U2480 (N_2480,N_1641,N_1576);
xnor U2481 (N_2481,N_1633,N_1597);
nand U2482 (N_2482,N_1595,N_1435);
and U2483 (N_2483,N_1635,N_1926);
or U2484 (N_2484,N_1173,N_1367);
nand U2485 (N_2485,N_1335,N_1882);
and U2486 (N_2486,N_1556,N_1373);
and U2487 (N_2487,N_1539,N_1302);
nand U2488 (N_2488,N_1680,N_1663);
or U2489 (N_2489,N_1565,N_1491);
or U2490 (N_2490,N_1899,N_1807);
or U2491 (N_2491,N_1721,N_1550);
nor U2492 (N_2492,N_1812,N_1167);
xnor U2493 (N_2493,N_1265,N_1588);
xor U2494 (N_2494,N_1375,N_1128);
xor U2495 (N_2495,N_1116,N_1736);
nor U2496 (N_2496,N_1317,N_1639);
and U2497 (N_2497,N_1086,N_1399);
nand U2498 (N_2498,N_1268,N_1602);
or U2499 (N_2499,N_1638,N_1366);
or U2500 (N_2500,N_1298,N_1519);
xnor U2501 (N_2501,N_1980,N_1864);
nor U2502 (N_2502,N_1113,N_1733);
and U2503 (N_2503,N_1147,N_1563);
xnor U2504 (N_2504,N_1931,N_1770);
or U2505 (N_2505,N_1038,N_1018);
or U2506 (N_2506,N_1676,N_1720);
xnor U2507 (N_2507,N_1036,N_1027);
or U2508 (N_2508,N_1746,N_1984);
or U2509 (N_2509,N_1202,N_1020);
and U2510 (N_2510,N_1617,N_1166);
or U2511 (N_2511,N_1242,N_1913);
or U2512 (N_2512,N_1957,N_1499);
nor U2513 (N_2513,N_1118,N_1798);
nand U2514 (N_2514,N_1984,N_1038);
nor U2515 (N_2515,N_1976,N_1087);
and U2516 (N_2516,N_1190,N_1629);
nand U2517 (N_2517,N_1346,N_1514);
xor U2518 (N_2518,N_1576,N_1731);
xnor U2519 (N_2519,N_1962,N_1379);
nor U2520 (N_2520,N_1512,N_1547);
nor U2521 (N_2521,N_1299,N_1982);
nor U2522 (N_2522,N_1932,N_1778);
and U2523 (N_2523,N_1858,N_1874);
nor U2524 (N_2524,N_1268,N_1337);
or U2525 (N_2525,N_1110,N_1073);
and U2526 (N_2526,N_1390,N_1641);
xor U2527 (N_2527,N_1700,N_1749);
nor U2528 (N_2528,N_1963,N_1443);
and U2529 (N_2529,N_1786,N_1004);
or U2530 (N_2530,N_1611,N_1237);
nand U2531 (N_2531,N_1094,N_1422);
or U2532 (N_2532,N_1626,N_1157);
nor U2533 (N_2533,N_1484,N_1513);
nor U2534 (N_2534,N_1441,N_1940);
xor U2535 (N_2535,N_1721,N_1750);
nand U2536 (N_2536,N_1519,N_1546);
and U2537 (N_2537,N_1716,N_1727);
nor U2538 (N_2538,N_1338,N_1873);
nand U2539 (N_2539,N_1344,N_1322);
or U2540 (N_2540,N_1176,N_1324);
and U2541 (N_2541,N_1061,N_1585);
nor U2542 (N_2542,N_1800,N_1667);
nor U2543 (N_2543,N_1359,N_1600);
or U2544 (N_2544,N_1652,N_1587);
xor U2545 (N_2545,N_1183,N_1967);
and U2546 (N_2546,N_1859,N_1943);
and U2547 (N_2547,N_1822,N_1928);
xor U2548 (N_2548,N_1200,N_1820);
or U2549 (N_2549,N_1902,N_1604);
xnor U2550 (N_2550,N_1617,N_1963);
or U2551 (N_2551,N_1407,N_1273);
or U2552 (N_2552,N_1977,N_1142);
nor U2553 (N_2553,N_1675,N_1177);
or U2554 (N_2554,N_1818,N_1662);
and U2555 (N_2555,N_1911,N_1952);
or U2556 (N_2556,N_1852,N_1640);
or U2557 (N_2557,N_1963,N_1779);
xnor U2558 (N_2558,N_1585,N_1074);
and U2559 (N_2559,N_1660,N_1167);
or U2560 (N_2560,N_1947,N_1196);
or U2561 (N_2561,N_1267,N_1386);
nand U2562 (N_2562,N_1658,N_1616);
or U2563 (N_2563,N_1167,N_1984);
or U2564 (N_2564,N_1880,N_1112);
xor U2565 (N_2565,N_1544,N_1646);
or U2566 (N_2566,N_1599,N_1286);
xor U2567 (N_2567,N_1964,N_1299);
and U2568 (N_2568,N_1187,N_1881);
nor U2569 (N_2569,N_1816,N_1969);
nand U2570 (N_2570,N_1863,N_1397);
and U2571 (N_2571,N_1111,N_1777);
nor U2572 (N_2572,N_1533,N_1853);
or U2573 (N_2573,N_1291,N_1667);
nand U2574 (N_2574,N_1600,N_1425);
and U2575 (N_2575,N_1577,N_1266);
xor U2576 (N_2576,N_1593,N_1931);
or U2577 (N_2577,N_1021,N_1272);
and U2578 (N_2578,N_1786,N_1438);
and U2579 (N_2579,N_1066,N_1882);
and U2580 (N_2580,N_1263,N_1489);
nor U2581 (N_2581,N_1132,N_1939);
or U2582 (N_2582,N_1165,N_1439);
nor U2583 (N_2583,N_1176,N_1064);
and U2584 (N_2584,N_1518,N_1690);
or U2585 (N_2585,N_1275,N_1350);
xnor U2586 (N_2586,N_1120,N_1805);
and U2587 (N_2587,N_1589,N_1013);
nand U2588 (N_2588,N_1236,N_1846);
and U2589 (N_2589,N_1378,N_1932);
and U2590 (N_2590,N_1752,N_1913);
or U2591 (N_2591,N_1266,N_1804);
and U2592 (N_2592,N_1254,N_1688);
and U2593 (N_2593,N_1859,N_1702);
xor U2594 (N_2594,N_1330,N_1713);
nor U2595 (N_2595,N_1059,N_1047);
and U2596 (N_2596,N_1275,N_1953);
and U2597 (N_2597,N_1079,N_1345);
nand U2598 (N_2598,N_1785,N_1714);
xnor U2599 (N_2599,N_1655,N_1966);
and U2600 (N_2600,N_1109,N_1152);
nand U2601 (N_2601,N_1787,N_1282);
and U2602 (N_2602,N_1064,N_1450);
xnor U2603 (N_2603,N_1041,N_1008);
nand U2604 (N_2604,N_1212,N_1892);
xnor U2605 (N_2605,N_1144,N_1844);
nor U2606 (N_2606,N_1301,N_1832);
xnor U2607 (N_2607,N_1675,N_1848);
nand U2608 (N_2608,N_1219,N_1901);
nor U2609 (N_2609,N_1522,N_1081);
nor U2610 (N_2610,N_1817,N_1130);
nor U2611 (N_2611,N_1450,N_1497);
and U2612 (N_2612,N_1880,N_1048);
nor U2613 (N_2613,N_1966,N_1650);
nand U2614 (N_2614,N_1384,N_1870);
or U2615 (N_2615,N_1566,N_1021);
nor U2616 (N_2616,N_1450,N_1901);
xor U2617 (N_2617,N_1039,N_1501);
nor U2618 (N_2618,N_1702,N_1988);
nand U2619 (N_2619,N_1228,N_1054);
nor U2620 (N_2620,N_1238,N_1607);
xnor U2621 (N_2621,N_1712,N_1754);
nor U2622 (N_2622,N_1475,N_1623);
or U2623 (N_2623,N_1007,N_1050);
or U2624 (N_2624,N_1755,N_1907);
and U2625 (N_2625,N_1320,N_1541);
xor U2626 (N_2626,N_1986,N_1199);
xnor U2627 (N_2627,N_1818,N_1459);
nand U2628 (N_2628,N_1742,N_1554);
and U2629 (N_2629,N_1198,N_1847);
nor U2630 (N_2630,N_1490,N_1459);
xor U2631 (N_2631,N_1563,N_1953);
and U2632 (N_2632,N_1114,N_1211);
xor U2633 (N_2633,N_1504,N_1831);
nand U2634 (N_2634,N_1725,N_1416);
xnor U2635 (N_2635,N_1900,N_1683);
or U2636 (N_2636,N_1118,N_1784);
nand U2637 (N_2637,N_1451,N_1415);
and U2638 (N_2638,N_1461,N_1530);
or U2639 (N_2639,N_1764,N_1614);
and U2640 (N_2640,N_1923,N_1360);
xnor U2641 (N_2641,N_1232,N_1850);
nor U2642 (N_2642,N_1526,N_1947);
or U2643 (N_2643,N_1001,N_1541);
or U2644 (N_2644,N_1869,N_1241);
xnor U2645 (N_2645,N_1700,N_1757);
nor U2646 (N_2646,N_1341,N_1691);
nor U2647 (N_2647,N_1764,N_1291);
and U2648 (N_2648,N_1999,N_1760);
and U2649 (N_2649,N_1791,N_1114);
xor U2650 (N_2650,N_1804,N_1275);
nor U2651 (N_2651,N_1396,N_1543);
nand U2652 (N_2652,N_1433,N_1221);
or U2653 (N_2653,N_1542,N_1078);
and U2654 (N_2654,N_1401,N_1678);
nand U2655 (N_2655,N_1511,N_1299);
or U2656 (N_2656,N_1334,N_1800);
or U2657 (N_2657,N_1997,N_1969);
xor U2658 (N_2658,N_1609,N_1535);
and U2659 (N_2659,N_1619,N_1256);
nor U2660 (N_2660,N_1285,N_1521);
nor U2661 (N_2661,N_1427,N_1352);
xnor U2662 (N_2662,N_1560,N_1271);
xor U2663 (N_2663,N_1745,N_1539);
and U2664 (N_2664,N_1648,N_1025);
nand U2665 (N_2665,N_1319,N_1197);
nor U2666 (N_2666,N_1551,N_1882);
nor U2667 (N_2667,N_1024,N_1914);
nand U2668 (N_2668,N_1293,N_1333);
nand U2669 (N_2669,N_1236,N_1542);
nor U2670 (N_2670,N_1271,N_1118);
and U2671 (N_2671,N_1673,N_1560);
or U2672 (N_2672,N_1404,N_1057);
xnor U2673 (N_2673,N_1811,N_1675);
and U2674 (N_2674,N_1475,N_1973);
nor U2675 (N_2675,N_1562,N_1319);
and U2676 (N_2676,N_1665,N_1833);
or U2677 (N_2677,N_1635,N_1226);
xor U2678 (N_2678,N_1394,N_1153);
and U2679 (N_2679,N_1581,N_1404);
or U2680 (N_2680,N_1044,N_1543);
nor U2681 (N_2681,N_1610,N_1344);
or U2682 (N_2682,N_1483,N_1667);
xor U2683 (N_2683,N_1981,N_1309);
and U2684 (N_2684,N_1521,N_1430);
or U2685 (N_2685,N_1343,N_1652);
nand U2686 (N_2686,N_1382,N_1832);
and U2687 (N_2687,N_1603,N_1451);
xnor U2688 (N_2688,N_1924,N_1326);
xor U2689 (N_2689,N_1440,N_1570);
nand U2690 (N_2690,N_1356,N_1798);
and U2691 (N_2691,N_1322,N_1250);
nand U2692 (N_2692,N_1244,N_1176);
nor U2693 (N_2693,N_1430,N_1520);
nand U2694 (N_2694,N_1380,N_1589);
and U2695 (N_2695,N_1546,N_1108);
nand U2696 (N_2696,N_1920,N_1536);
nor U2697 (N_2697,N_1217,N_1499);
nand U2698 (N_2698,N_1733,N_1418);
nor U2699 (N_2699,N_1340,N_1541);
xnor U2700 (N_2700,N_1367,N_1816);
nor U2701 (N_2701,N_1954,N_1107);
nand U2702 (N_2702,N_1660,N_1362);
nand U2703 (N_2703,N_1245,N_1924);
nor U2704 (N_2704,N_1994,N_1068);
nand U2705 (N_2705,N_1878,N_1056);
or U2706 (N_2706,N_1920,N_1567);
and U2707 (N_2707,N_1920,N_1893);
nand U2708 (N_2708,N_1201,N_1542);
xor U2709 (N_2709,N_1283,N_1462);
nand U2710 (N_2710,N_1552,N_1240);
nor U2711 (N_2711,N_1415,N_1803);
nor U2712 (N_2712,N_1592,N_1340);
or U2713 (N_2713,N_1309,N_1015);
and U2714 (N_2714,N_1562,N_1881);
and U2715 (N_2715,N_1621,N_1645);
nor U2716 (N_2716,N_1103,N_1815);
nor U2717 (N_2717,N_1797,N_1597);
nand U2718 (N_2718,N_1642,N_1488);
and U2719 (N_2719,N_1732,N_1006);
and U2720 (N_2720,N_1622,N_1689);
and U2721 (N_2721,N_1038,N_1474);
nand U2722 (N_2722,N_1603,N_1237);
or U2723 (N_2723,N_1660,N_1869);
or U2724 (N_2724,N_1608,N_1006);
or U2725 (N_2725,N_1242,N_1294);
and U2726 (N_2726,N_1714,N_1879);
nor U2727 (N_2727,N_1496,N_1545);
and U2728 (N_2728,N_1078,N_1487);
or U2729 (N_2729,N_1065,N_1737);
or U2730 (N_2730,N_1830,N_1229);
nand U2731 (N_2731,N_1547,N_1031);
and U2732 (N_2732,N_1334,N_1366);
nand U2733 (N_2733,N_1544,N_1137);
xor U2734 (N_2734,N_1762,N_1656);
xor U2735 (N_2735,N_1672,N_1095);
and U2736 (N_2736,N_1649,N_1114);
and U2737 (N_2737,N_1372,N_1202);
and U2738 (N_2738,N_1402,N_1872);
nand U2739 (N_2739,N_1772,N_1087);
nor U2740 (N_2740,N_1957,N_1836);
nor U2741 (N_2741,N_1573,N_1100);
or U2742 (N_2742,N_1039,N_1063);
or U2743 (N_2743,N_1338,N_1129);
xor U2744 (N_2744,N_1478,N_1807);
nor U2745 (N_2745,N_1077,N_1261);
nor U2746 (N_2746,N_1760,N_1012);
and U2747 (N_2747,N_1990,N_1055);
and U2748 (N_2748,N_1345,N_1236);
nand U2749 (N_2749,N_1686,N_1751);
or U2750 (N_2750,N_1833,N_1077);
xnor U2751 (N_2751,N_1446,N_1506);
xnor U2752 (N_2752,N_1082,N_1695);
nand U2753 (N_2753,N_1757,N_1350);
nor U2754 (N_2754,N_1907,N_1094);
xor U2755 (N_2755,N_1848,N_1517);
and U2756 (N_2756,N_1453,N_1718);
nor U2757 (N_2757,N_1651,N_1158);
xor U2758 (N_2758,N_1122,N_1830);
xor U2759 (N_2759,N_1263,N_1167);
or U2760 (N_2760,N_1282,N_1167);
xor U2761 (N_2761,N_1567,N_1164);
nor U2762 (N_2762,N_1849,N_1554);
nor U2763 (N_2763,N_1477,N_1023);
and U2764 (N_2764,N_1374,N_1329);
nor U2765 (N_2765,N_1288,N_1222);
nand U2766 (N_2766,N_1357,N_1096);
xor U2767 (N_2767,N_1337,N_1672);
or U2768 (N_2768,N_1809,N_1998);
nand U2769 (N_2769,N_1339,N_1611);
xor U2770 (N_2770,N_1019,N_1860);
nor U2771 (N_2771,N_1895,N_1962);
nand U2772 (N_2772,N_1903,N_1962);
nand U2773 (N_2773,N_1011,N_1550);
nor U2774 (N_2774,N_1122,N_1684);
or U2775 (N_2775,N_1014,N_1029);
xor U2776 (N_2776,N_1557,N_1808);
and U2777 (N_2777,N_1789,N_1009);
or U2778 (N_2778,N_1697,N_1844);
xnor U2779 (N_2779,N_1747,N_1777);
xnor U2780 (N_2780,N_1226,N_1934);
xor U2781 (N_2781,N_1477,N_1906);
or U2782 (N_2782,N_1211,N_1942);
xor U2783 (N_2783,N_1906,N_1625);
and U2784 (N_2784,N_1381,N_1716);
or U2785 (N_2785,N_1316,N_1333);
xor U2786 (N_2786,N_1906,N_1284);
or U2787 (N_2787,N_1132,N_1301);
xor U2788 (N_2788,N_1104,N_1079);
nor U2789 (N_2789,N_1599,N_1978);
nor U2790 (N_2790,N_1061,N_1576);
and U2791 (N_2791,N_1642,N_1557);
and U2792 (N_2792,N_1955,N_1496);
and U2793 (N_2793,N_1864,N_1065);
xnor U2794 (N_2794,N_1056,N_1238);
and U2795 (N_2795,N_1789,N_1275);
and U2796 (N_2796,N_1978,N_1915);
nor U2797 (N_2797,N_1193,N_1217);
nand U2798 (N_2798,N_1702,N_1478);
and U2799 (N_2799,N_1595,N_1454);
and U2800 (N_2800,N_1579,N_1730);
nand U2801 (N_2801,N_1373,N_1037);
nor U2802 (N_2802,N_1637,N_1731);
nor U2803 (N_2803,N_1891,N_1943);
and U2804 (N_2804,N_1340,N_1809);
nand U2805 (N_2805,N_1350,N_1302);
nand U2806 (N_2806,N_1758,N_1970);
or U2807 (N_2807,N_1168,N_1486);
or U2808 (N_2808,N_1273,N_1553);
nor U2809 (N_2809,N_1385,N_1450);
or U2810 (N_2810,N_1849,N_1993);
nor U2811 (N_2811,N_1948,N_1728);
and U2812 (N_2812,N_1165,N_1118);
xnor U2813 (N_2813,N_1702,N_1289);
nand U2814 (N_2814,N_1810,N_1034);
nand U2815 (N_2815,N_1666,N_1176);
xor U2816 (N_2816,N_1642,N_1627);
nand U2817 (N_2817,N_1766,N_1002);
nor U2818 (N_2818,N_1213,N_1971);
xor U2819 (N_2819,N_1548,N_1723);
nand U2820 (N_2820,N_1795,N_1598);
and U2821 (N_2821,N_1849,N_1205);
or U2822 (N_2822,N_1252,N_1762);
xnor U2823 (N_2823,N_1722,N_1780);
and U2824 (N_2824,N_1752,N_1038);
nor U2825 (N_2825,N_1451,N_1623);
xor U2826 (N_2826,N_1069,N_1064);
nand U2827 (N_2827,N_1538,N_1074);
nor U2828 (N_2828,N_1342,N_1518);
xor U2829 (N_2829,N_1896,N_1402);
nor U2830 (N_2830,N_1774,N_1172);
nand U2831 (N_2831,N_1310,N_1052);
and U2832 (N_2832,N_1473,N_1582);
and U2833 (N_2833,N_1027,N_1897);
xnor U2834 (N_2834,N_1043,N_1448);
nor U2835 (N_2835,N_1816,N_1120);
and U2836 (N_2836,N_1486,N_1170);
and U2837 (N_2837,N_1120,N_1493);
and U2838 (N_2838,N_1140,N_1615);
nor U2839 (N_2839,N_1552,N_1185);
or U2840 (N_2840,N_1408,N_1987);
nand U2841 (N_2841,N_1606,N_1750);
or U2842 (N_2842,N_1571,N_1984);
or U2843 (N_2843,N_1621,N_1466);
and U2844 (N_2844,N_1429,N_1040);
xnor U2845 (N_2845,N_1685,N_1854);
xnor U2846 (N_2846,N_1931,N_1189);
nor U2847 (N_2847,N_1822,N_1431);
nor U2848 (N_2848,N_1833,N_1229);
nand U2849 (N_2849,N_1995,N_1002);
or U2850 (N_2850,N_1049,N_1289);
xor U2851 (N_2851,N_1569,N_1606);
and U2852 (N_2852,N_1975,N_1536);
or U2853 (N_2853,N_1159,N_1743);
nor U2854 (N_2854,N_1497,N_1816);
and U2855 (N_2855,N_1935,N_1544);
nand U2856 (N_2856,N_1129,N_1687);
or U2857 (N_2857,N_1914,N_1740);
xnor U2858 (N_2858,N_1351,N_1854);
or U2859 (N_2859,N_1475,N_1124);
and U2860 (N_2860,N_1575,N_1736);
and U2861 (N_2861,N_1525,N_1173);
nand U2862 (N_2862,N_1884,N_1649);
or U2863 (N_2863,N_1564,N_1364);
nand U2864 (N_2864,N_1431,N_1089);
or U2865 (N_2865,N_1787,N_1124);
or U2866 (N_2866,N_1548,N_1227);
or U2867 (N_2867,N_1867,N_1719);
nand U2868 (N_2868,N_1927,N_1561);
and U2869 (N_2869,N_1405,N_1392);
or U2870 (N_2870,N_1252,N_1063);
xnor U2871 (N_2871,N_1242,N_1528);
nor U2872 (N_2872,N_1732,N_1962);
nand U2873 (N_2873,N_1391,N_1962);
nand U2874 (N_2874,N_1586,N_1201);
or U2875 (N_2875,N_1685,N_1857);
or U2876 (N_2876,N_1675,N_1406);
nand U2877 (N_2877,N_1079,N_1691);
xnor U2878 (N_2878,N_1154,N_1282);
or U2879 (N_2879,N_1053,N_1007);
nand U2880 (N_2880,N_1711,N_1294);
nand U2881 (N_2881,N_1124,N_1261);
nor U2882 (N_2882,N_1180,N_1045);
nand U2883 (N_2883,N_1200,N_1480);
or U2884 (N_2884,N_1251,N_1523);
or U2885 (N_2885,N_1230,N_1312);
and U2886 (N_2886,N_1237,N_1239);
or U2887 (N_2887,N_1265,N_1566);
and U2888 (N_2888,N_1648,N_1183);
nand U2889 (N_2889,N_1309,N_1214);
nand U2890 (N_2890,N_1752,N_1451);
xnor U2891 (N_2891,N_1525,N_1956);
or U2892 (N_2892,N_1270,N_1122);
nor U2893 (N_2893,N_1966,N_1925);
nand U2894 (N_2894,N_1895,N_1834);
nand U2895 (N_2895,N_1357,N_1945);
nor U2896 (N_2896,N_1203,N_1264);
and U2897 (N_2897,N_1890,N_1180);
nor U2898 (N_2898,N_1792,N_1698);
nand U2899 (N_2899,N_1671,N_1005);
and U2900 (N_2900,N_1574,N_1797);
or U2901 (N_2901,N_1776,N_1061);
nor U2902 (N_2902,N_1588,N_1376);
nand U2903 (N_2903,N_1007,N_1528);
nand U2904 (N_2904,N_1479,N_1834);
nand U2905 (N_2905,N_1454,N_1003);
and U2906 (N_2906,N_1105,N_1569);
or U2907 (N_2907,N_1610,N_1480);
or U2908 (N_2908,N_1228,N_1653);
nand U2909 (N_2909,N_1534,N_1039);
and U2910 (N_2910,N_1691,N_1721);
nand U2911 (N_2911,N_1446,N_1192);
nand U2912 (N_2912,N_1607,N_1083);
and U2913 (N_2913,N_1994,N_1960);
and U2914 (N_2914,N_1095,N_1803);
nor U2915 (N_2915,N_1546,N_1825);
and U2916 (N_2916,N_1445,N_1696);
nor U2917 (N_2917,N_1255,N_1351);
nand U2918 (N_2918,N_1899,N_1611);
nand U2919 (N_2919,N_1676,N_1103);
or U2920 (N_2920,N_1651,N_1690);
and U2921 (N_2921,N_1502,N_1834);
or U2922 (N_2922,N_1797,N_1364);
xnor U2923 (N_2923,N_1388,N_1599);
and U2924 (N_2924,N_1237,N_1783);
nand U2925 (N_2925,N_1346,N_1779);
xor U2926 (N_2926,N_1546,N_1090);
nand U2927 (N_2927,N_1455,N_1372);
and U2928 (N_2928,N_1002,N_1596);
xnor U2929 (N_2929,N_1348,N_1634);
nand U2930 (N_2930,N_1331,N_1802);
nand U2931 (N_2931,N_1581,N_1431);
and U2932 (N_2932,N_1121,N_1002);
nand U2933 (N_2933,N_1660,N_1818);
nor U2934 (N_2934,N_1923,N_1949);
and U2935 (N_2935,N_1411,N_1359);
and U2936 (N_2936,N_1483,N_1683);
and U2937 (N_2937,N_1013,N_1877);
nand U2938 (N_2938,N_1852,N_1190);
and U2939 (N_2939,N_1293,N_1234);
or U2940 (N_2940,N_1025,N_1138);
nor U2941 (N_2941,N_1513,N_1517);
nand U2942 (N_2942,N_1806,N_1854);
and U2943 (N_2943,N_1043,N_1255);
xor U2944 (N_2944,N_1193,N_1544);
xnor U2945 (N_2945,N_1715,N_1248);
xor U2946 (N_2946,N_1606,N_1038);
nor U2947 (N_2947,N_1820,N_1514);
nand U2948 (N_2948,N_1393,N_1593);
and U2949 (N_2949,N_1905,N_1134);
xor U2950 (N_2950,N_1291,N_1851);
nor U2951 (N_2951,N_1044,N_1855);
nand U2952 (N_2952,N_1320,N_1417);
nand U2953 (N_2953,N_1245,N_1193);
nor U2954 (N_2954,N_1649,N_1629);
and U2955 (N_2955,N_1883,N_1740);
and U2956 (N_2956,N_1337,N_1760);
nor U2957 (N_2957,N_1515,N_1167);
nor U2958 (N_2958,N_1266,N_1168);
and U2959 (N_2959,N_1010,N_1840);
or U2960 (N_2960,N_1677,N_1812);
or U2961 (N_2961,N_1453,N_1825);
or U2962 (N_2962,N_1735,N_1415);
nor U2963 (N_2963,N_1223,N_1105);
or U2964 (N_2964,N_1482,N_1517);
nor U2965 (N_2965,N_1861,N_1147);
and U2966 (N_2966,N_1603,N_1661);
or U2967 (N_2967,N_1018,N_1110);
xnor U2968 (N_2968,N_1284,N_1890);
nor U2969 (N_2969,N_1911,N_1786);
and U2970 (N_2970,N_1461,N_1565);
xor U2971 (N_2971,N_1389,N_1010);
or U2972 (N_2972,N_1097,N_1334);
nor U2973 (N_2973,N_1374,N_1105);
or U2974 (N_2974,N_1074,N_1854);
or U2975 (N_2975,N_1148,N_1259);
or U2976 (N_2976,N_1131,N_1476);
nor U2977 (N_2977,N_1761,N_1995);
nand U2978 (N_2978,N_1858,N_1939);
and U2979 (N_2979,N_1229,N_1854);
or U2980 (N_2980,N_1688,N_1847);
and U2981 (N_2981,N_1468,N_1501);
and U2982 (N_2982,N_1749,N_1384);
xor U2983 (N_2983,N_1663,N_1006);
nand U2984 (N_2984,N_1530,N_1455);
xor U2985 (N_2985,N_1533,N_1631);
xor U2986 (N_2986,N_1017,N_1775);
nand U2987 (N_2987,N_1144,N_1674);
nor U2988 (N_2988,N_1887,N_1037);
and U2989 (N_2989,N_1752,N_1227);
nand U2990 (N_2990,N_1700,N_1212);
nand U2991 (N_2991,N_1960,N_1403);
xnor U2992 (N_2992,N_1047,N_1078);
xor U2993 (N_2993,N_1726,N_1333);
nor U2994 (N_2994,N_1214,N_1195);
nor U2995 (N_2995,N_1126,N_1699);
nand U2996 (N_2996,N_1686,N_1610);
and U2997 (N_2997,N_1993,N_1075);
nor U2998 (N_2998,N_1236,N_1933);
or U2999 (N_2999,N_1725,N_1816);
nand UO_0 (O_0,N_2985,N_2941);
or UO_1 (O_1,N_2836,N_2904);
nor UO_2 (O_2,N_2827,N_2529);
or UO_3 (O_3,N_2027,N_2352);
nand UO_4 (O_4,N_2866,N_2605);
or UO_5 (O_5,N_2357,N_2007);
nor UO_6 (O_6,N_2344,N_2032);
or UO_7 (O_7,N_2256,N_2955);
and UO_8 (O_8,N_2361,N_2432);
and UO_9 (O_9,N_2918,N_2762);
nor UO_10 (O_10,N_2623,N_2916);
nor UO_11 (O_11,N_2867,N_2516);
xor UO_12 (O_12,N_2494,N_2230);
or UO_13 (O_13,N_2135,N_2094);
or UO_14 (O_14,N_2860,N_2407);
nor UO_15 (O_15,N_2459,N_2627);
nor UO_16 (O_16,N_2336,N_2987);
xor UO_17 (O_17,N_2728,N_2901);
or UO_18 (O_18,N_2808,N_2633);
or UO_19 (O_19,N_2386,N_2495);
and UO_20 (O_20,N_2306,N_2790);
nand UO_21 (O_21,N_2366,N_2883);
or UO_22 (O_22,N_2136,N_2097);
nand UO_23 (O_23,N_2881,N_2332);
and UO_24 (O_24,N_2445,N_2809);
and UO_25 (O_25,N_2310,N_2291);
and UO_26 (O_26,N_2069,N_2249);
xnor UO_27 (O_27,N_2638,N_2665);
or UO_28 (O_28,N_2744,N_2008);
xor UO_29 (O_29,N_2182,N_2927);
xnor UO_30 (O_30,N_2909,N_2364);
nand UO_31 (O_31,N_2360,N_2620);
or UO_32 (O_32,N_2565,N_2142);
or UO_33 (O_33,N_2089,N_2754);
or UO_34 (O_34,N_2018,N_2046);
nor UO_35 (O_35,N_2546,N_2823);
nand UO_36 (O_36,N_2646,N_2045);
nor UO_37 (O_37,N_2862,N_2952);
xor UO_38 (O_38,N_2537,N_2430);
and UO_39 (O_39,N_2947,N_2213);
nand UO_40 (O_40,N_2966,N_2300);
or UO_41 (O_41,N_2598,N_2267);
or UO_42 (O_42,N_2676,N_2096);
nor UO_43 (O_43,N_2457,N_2643);
or UO_44 (O_44,N_2736,N_2538);
nor UO_45 (O_45,N_2812,N_2835);
nand UO_46 (O_46,N_2257,N_2189);
and UO_47 (O_47,N_2070,N_2458);
nor UO_48 (O_48,N_2346,N_2961);
or UO_49 (O_49,N_2515,N_2659);
nand UO_50 (O_50,N_2307,N_2002);
nor UO_51 (O_51,N_2394,N_2131);
xnor UO_52 (O_52,N_2130,N_2340);
xor UO_53 (O_53,N_2421,N_2943);
nand UO_54 (O_54,N_2710,N_2844);
nand UO_55 (O_55,N_2855,N_2669);
nor UO_56 (O_56,N_2705,N_2040);
nand UO_57 (O_57,N_2724,N_2708);
and UO_58 (O_58,N_2850,N_2269);
or UO_59 (O_59,N_2365,N_2959);
or UO_60 (O_60,N_2986,N_2577);
nor UO_61 (O_61,N_2272,N_2434);
and UO_62 (O_62,N_2036,N_2422);
nand UO_63 (O_63,N_2737,N_2540);
nor UO_64 (O_64,N_2380,N_2374);
and UO_65 (O_65,N_2181,N_2799);
nand UO_66 (O_66,N_2913,N_2677);
and UO_67 (O_67,N_2103,N_2852);
or UO_68 (O_68,N_2314,N_2542);
and UO_69 (O_69,N_2834,N_2719);
xor UO_70 (O_70,N_2025,N_2639);
nor UO_71 (O_71,N_2281,N_2408);
xor UO_72 (O_72,N_2609,N_2680);
or UO_73 (O_73,N_2075,N_2304);
xor UO_74 (O_74,N_2484,N_2173);
or UO_75 (O_75,N_2576,N_2150);
xor UO_76 (O_76,N_2133,N_2183);
nor UO_77 (O_77,N_2419,N_2193);
nor UO_78 (O_78,N_2532,N_2260);
nand UO_79 (O_79,N_2675,N_2750);
nor UO_80 (O_80,N_2437,N_2104);
xnor UO_81 (O_81,N_2539,N_2388);
or UO_82 (O_82,N_2218,N_2124);
and UO_83 (O_83,N_2524,N_2425);
xor UO_84 (O_84,N_2192,N_2163);
and UO_85 (O_85,N_2868,N_2995);
or UO_86 (O_86,N_2777,N_2517);
nand UO_87 (O_87,N_2606,N_2456);
or UO_88 (O_88,N_2043,N_2297);
nor UO_89 (O_89,N_2201,N_2846);
xor UO_90 (O_90,N_2936,N_2491);
nand UO_91 (O_91,N_2452,N_2940);
xnor UO_92 (O_92,N_2333,N_2899);
nand UO_93 (O_93,N_2994,N_2423);
or UO_94 (O_94,N_2514,N_2885);
and UO_95 (O_95,N_2701,N_2420);
or UO_96 (O_96,N_2259,N_2205);
nand UO_97 (O_97,N_2871,N_2660);
xnor UO_98 (O_98,N_2015,N_2058);
or UO_99 (O_99,N_2263,N_2608);
xnor UO_100 (O_100,N_2837,N_2552);
xor UO_101 (O_101,N_2636,N_2738);
and UO_102 (O_102,N_2321,N_2923);
or UO_103 (O_103,N_2513,N_2328);
xnor UO_104 (O_104,N_2739,N_2818);
or UO_105 (O_105,N_2723,N_2689);
xnor UO_106 (O_106,N_2671,N_2649);
xnor UO_107 (O_107,N_2479,N_2893);
or UO_108 (O_108,N_2587,N_2915);
or UO_109 (O_109,N_2221,N_2604);
nand UO_110 (O_110,N_2519,N_2946);
and UO_111 (O_111,N_2702,N_2165);
nor UO_112 (O_112,N_2897,N_2861);
xnor UO_113 (O_113,N_2082,N_2718);
nor UO_114 (O_114,N_2833,N_2455);
nor UO_115 (O_115,N_2038,N_2490);
nand UO_116 (O_116,N_2924,N_2265);
nor UO_117 (O_117,N_2440,N_2787);
nand UO_118 (O_118,N_2476,N_2976);
or UO_119 (O_119,N_2481,N_2343);
nand UO_120 (O_120,N_2042,N_2877);
or UO_121 (O_121,N_2984,N_2222);
nor UO_122 (O_122,N_2957,N_2559);
xor UO_123 (O_123,N_2122,N_2982);
or UO_124 (O_124,N_2789,N_2528);
nor UO_125 (O_125,N_2435,N_2236);
or UO_126 (O_126,N_2535,N_2856);
or UO_127 (O_127,N_2246,N_2498);
nor UO_128 (O_128,N_2759,N_2840);
xnor UO_129 (O_129,N_2757,N_2406);
xnor UO_130 (O_130,N_2109,N_2726);
nand UO_131 (O_131,N_2832,N_2696);
and UO_132 (O_132,N_2411,N_2387);
nand UO_133 (O_133,N_2900,N_2733);
and UO_134 (O_134,N_2268,N_2474);
nor UO_135 (O_135,N_2238,N_2115);
nand UO_136 (O_136,N_2804,N_2743);
xor UO_137 (O_137,N_2377,N_2721);
nand UO_138 (O_138,N_2037,N_2323);
xnor UO_139 (O_139,N_2108,N_2854);
nor UO_140 (O_140,N_2751,N_2402);
nor UO_141 (O_141,N_2282,N_2666);
and UO_142 (O_142,N_2467,N_2796);
nor UO_143 (O_143,N_2353,N_2198);
nand UO_144 (O_144,N_2504,N_2595);
nor UO_145 (O_145,N_2890,N_2442);
nor UO_146 (O_146,N_2217,N_2295);
and UO_147 (O_147,N_2039,N_2258);
or UO_148 (O_148,N_2146,N_2550);
nand UO_149 (O_149,N_2313,N_2983);
or UO_150 (O_150,N_2859,N_2938);
nor UO_151 (O_151,N_2137,N_2869);
xor UO_152 (O_152,N_2932,N_2190);
xnor UO_153 (O_153,N_2057,N_2319);
nor UO_154 (O_154,N_2858,N_2488);
or UO_155 (O_155,N_2290,N_2596);
nand UO_156 (O_156,N_2906,N_2354);
or UO_157 (O_157,N_2134,N_2518);
or UO_158 (O_158,N_2814,N_2331);
or UO_159 (O_159,N_2016,N_2566);
nor UO_160 (O_160,N_2979,N_2468);
and UO_161 (O_161,N_2865,N_2254);
or UO_162 (O_162,N_2143,N_2351);
xor UO_163 (O_163,N_2229,N_2933);
nand UO_164 (O_164,N_2699,N_2911);
nor UO_165 (O_165,N_2475,N_2845);
nor UO_166 (O_166,N_2821,N_2673);
nand UO_167 (O_167,N_2303,N_2873);
nand UO_168 (O_168,N_2225,N_2647);
or UO_169 (O_169,N_2875,N_2747);
or UO_170 (O_170,N_2156,N_2228);
and UO_171 (O_171,N_2116,N_2090);
xnor UO_172 (O_172,N_2237,N_2059);
xnor UO_173 (O_173,N_2158,N_2298);
nor UO_174 (O_174,N_2155,N_2292);
xor UO_175 (O_175,N_2208,N_2065);
and UO_176 (O_176,N_2347,N_2500);
nor UO_177 (O_177,N_2655,N_2830);
nand UO_178 (O_178,N_2894,N_2782);
and UO_179 (O_179,N_2412,N_2969);
and UO_180 (O_180,N_2472,N_2775);
nand UO_181 (O_181,N_2632,N_2998);
nor UO_182 (O_182,N_2568,N_2811);
or UO_183 (O_183,N_2562,N_2641);
xnor UO_184 (O_184,N_2317,N_2921);
nand UO_185 (O_185,N_2473,N_2717);
nand UO_186 (O_186,N_2309,N_2887);
nor UO_187 (O_187,N_2417,N_2746);
nand UO_188 (O_188,N_2709,N_2574);
nor UO_189 (O_189,N_2591,N_2686);
nand UO_190 (O_190,N_2650,N_2917);
or UO_191 (O_191,N_2426,N_2978);
xor UO_192 (O_192,N_2478,N_2910);
and UO_193 (O_193,N_2822,N_2691);
nor UO_194 (O_194,N_2379,N_2575);
and UO_195 (O_195,N_2293,N_2391);
and UO_196 (O_196,N_2651,N_2993);
and UO_197 (O_197,N_2876,N_2048);
and UO_198 (O_198,N_2101,N_2684);
nor UO_199 (O_199,N_2278,N_2497);
nand UO_200 (O_200,N_2210,N_2872);
nor UO_201 (O_201,N_2960,N_2141);
and UO_202 (O_202,N_2005,N_2548);
and UO_203 (O_203,N_2630,N_2396);
xor UO_204 (O_204,N_2194,N_2054);
nor UO_205 (O_205,N_2017,N_2896);
xnor UO_206 (O_206,N_2447,N_2209);
nand UO_207 (O_207,N_2697,N_2783);
xor UO_208 (O_208,N_2224,N_2760);
or UO_209 (O_209,N_2363,N_2389);
xnor UO_210 (O_210,N_2892,N_2203);
and UO_211 (O_211,N_2195,N_2797);
xnor UO_212 (O_212,N_2919,N_2810);
nor UO_213 (O_213,N_2062,N_2202);
or UO_214 (O_214,N_2824,N_2099);
or UO_215 (O_215,N_2305,N_2398);
nand UO_216 (O_216,N_2006,N_2831);
and UO_217 (O_217,N_2414,N_2561);
and UO_218 (O_218,N_2712,N_2776);
or UO_219 (O_219,N_2191,N_2945);
and UO_220 (O_220,N_2589,N_2318);
xnor UO_221 (O_221,N_2327,N_2583);
nand UO_222 (O_222,N_2368,N_2977);
nand UO_223 (O_223,N_2345,N_2341);
nand UO_224 (O_224,N_2312,N_2645);
nor UO_225 (O_225,N_2077,N_2975);
and UO_226 (O_226,N_2286,N_2403);
and UO_227 (O_227,N_2247,N_2607);
nor UO_228 (O_228,N_2928,N_2326);
nor UO_229 (O_229,N_2756,N_2769);
or UO_230 (O_230,N_2569,N_2487);
and UO_231 (O_231,N_2968,N_2087);
nand UO_232 (O_232,N_2084,N_2092);
xor UO_233 (O_233,N_2055,N_2004);
nand UO_234 (O_234,N_2631,N_2681);
nor UO_235 (O_235,N_2180,N_2997);
nand UO_236 (O_236,N_2614,N_2079);
nor UO_237 (O_237,N_2857,N_2358);
nand UO_238 (O_238,N_2593,N_2214);
xnor UO_239 (O_239,N_2793,N_2572);
and UO_240 (O_240,N_2463,N_2428);
nand UO_241 (O_241,N_2287,N_2652);
nor UO_242 (O_242,N_2704,N_2151);
xnor UO_243 (O_243,N_2679,N_2851);
xnor UO_244 (O_244,N_2072,N_2207);
nor UO_245 (O_245,N_2599,N_2409);
nand UO_246 (O_246,N_2880,N_2695);
xor UO_247 (O_247,N_2579,N_2117);
nor UO_248 (O_248,N_2001,N_2176);
xnor UO_249 (O_249,N_2157,N_2698);
nand UO_250 (O_250,N_2742,N_2963);
xnor UO_251 (O_251,N_2688,N_2231);
or UO_252 (O_252,N_2289,N_2227);
nor UO_253 (O_253,N_2549,N_2700);
nand UO_254 (O_254,N_2640,N_2685);
xnor UO_255 (O_255,N_2621,N_2798);
and UO_256 (O_256,N_2235,N_2770);
nand UO_257 (O_257,N_2763,N_2634);
xnor UO_258 (O_258,N_2764,N_2602);
nor UO_259 (O_259,N_2240,N_2778);
xnor UO_260 (O_260,N_2073,N_2662);
nand UO_261 (O_261,N_2153,N_2536);
and UO_262 (O_262,N_2196,N_2277);
and UO_263 (O_263,N_2682,N_2590);
nor UO_264 (O_264,N_2758,N_2670);
or UO_265 (O_265,N_2772,N_2274);
and UO_266 (O_266,N_2898,N_2626);
nor UO_267 (O_267,N_2378,N_2908);
nor UO_268 (O_268,N_2107,N_2395);
xnor UO_269 (O_269,N_2616,N_2376);
and UO_270 (O_270,N_2989,N_2450);
or UO_271 (O_271,N_2544,N_2654);
or UO_272 (O_272,N_2653,N_2276);
and UO_273 (O_273,N_2088,N_2878);
and UO_274 (O_274,N_2800,N_2687);
or UO_275 (O_275,N_2988,N_2813);
and UO_276 (O_276,N_2618,N_2315);
nand UO_277 (O_277,N_2706,N_2939);
and UO_278 (O_278,N_2110,N_2356);
or UO_279 (O_279,N_2794,N_2418);
nand UO_280 (O_280,N_2248,N_2159);
and UO_281 (O_281,N_2971,N_2100);
and UO_282 (O_282,N_2505,N_2802);
or UO_283 (O_283,N_2842,N_2270);
nor UO_284 (O_284,N_2541,N_2126);
xor UO_285 (O_285,N_2774,N_2557);
xnor UO_286 (O_286,N_2725,N_2825);
xor UO_287 (O_287,N_2139,N_2339);
nand UO_288 (O_288,N_2111,N_2713);
nor UO_289 (O_289,N_2625,N_2041);
or UO_290 (O_290,N_2482,N_2922);
nand UO_291 (O_291,N_2429,N_2902);
or UO_292 (O_292,N_2161,N_2369);
or UO_293 (O_293,N_2106,N_2970);
nor UO_294 (O_294,N_2160,N_2571);
or UO_295 (O_295,N_2030,N_2464);
nand UO_296 (O_296,N_2991,N_2828);
xor UO_297 (O_297,N_2526,N_2570);
xnor UO_298 (O_298,N_2931,N_2393);
xnor UO_299 (O_299,N_2385,N_2980);
nor UO_300 (O_300,N_2220,N_2320);
xor UO_301 (O_301,N_2372,N_2252);
nand UO_302 (O_302,N_2330,N_2185);
nand UO_303 (O_303,N_2047,N_2337);
nand UO_304 (O_304,N_2817,N_2129);
and UO_305 (O_305,N_2439,N_2903);
nor UO_306 (O_306,N_2105,N_2113);
xor UO_307 (O_307,N_2567,N_2694);
or UO_308 (O_308,N_2044,N_2996);
xnor UO_309 (O_309,N_2508,N_2066);
nand UO_310 (O_310,N_2056,N_2740);
nor UO_311 (O_311,N_2410,N_2071);
or UO_312 (O_312,N_2815,N_2635);
xor UO_313 (O_313,N_2937,N_2466);
nor UO_314 (O_314,N_2471,N_2785);
nand UO_315 (O_315,N_2060,N_2453);
or UO_316 (O_316,N_2284,N_2147);
xor UO_317 (O_317,N_2973,N_2791);
or UO_318 (O_318,N_2128,N_2727);
nor UO_319 (O_319,N_2397,N_2879);
or UO_320 (O_320,N_2755,N_2948);
nand UO_321 (O_321,N_2853,N_2768);
and UO_322 (O_322,N_2035,N_2990);
xor UO_323 (O_323,N_2454,N_2807);
or UO_324 (O_324,N_2121,N_2507);
xnor UO_325 (O_325,N_2322,N_2226);
or UO_326 (O_326,N_2752,N_2912);
nand UO_327 (O_327,N_2171,N_2664);
and UO_328 (O_328,N_2801,N_2064);
xor UO_329 (O_329,N_2415,N_2648);
xor UO_330 (O_330,N_2642,N_2629);
nand UO_331 (O_331,N_2803,N_2886);
nor UO_332 (O_332,N_2371,N_2465);
or UO_333 (O_333,N_2958,N_2063);
nor UO_334 (O_334,N_2148,N_2020);
nor UO_335 (O_335,N_2543,N_2264);
xnor UO_336 (O_336,N_2527,N_2098);
xor UO_337 (O_337,N_2085,N_2753);
or UO_338 (O_338,N_2462,N_2443);
and UO_339 (O_339,N_2735,N_2847);
nand UO_340 (O_340,N_2348,N_2622);
nand UO_341 (O_341,N_2449,N_2283);
nand UO_342 (O_342,N_2436,N_2271);
xor UO_343 (O_343,N_2234,N_2863);
or UO_344 (O_344,N_2250,N_2657);
xnor UO_345 (O_345,N_2926,N_2241);
or UO_346 (O_346,N_2233,N_2152);
nand UO_347 (O_347,N_2503,N_2413);
xnor UO_348 (O_348,N_2714,N_2024);
nor UO_349 (O_349,N_2891,N_2184);
or UO_350 (O_350,N_2584,N_2496);
or UO_351 (O_351,N_2022,N_2509);
nand UO_352 (O_352,N_2033,N_2166);
xnor UO_353 (O_353,N_2469,N_2580);
nand UO_354 (O_354,N_2533,N_2175);
and UO_355 (O_355,N_2086,N_2010);
xor UO_356 (O_356,N_2311,N_2582);
xnor UO_357 (O_357,N_2232,N_2767);
or UO_358 (O_358,N_2053,N_2355);
xor UO_359 (O_359,N_2761,N_2551);
xor UO_360 (O_360,N_2784,N_2308);
or UO_361 (O_361,N_2944,N_2972);
nand UO_362 (O_362,N_2049,N_2781);
xnor UO_363 (O_363,N_2451,N_2149);
or UO_364 (O_364,N_2299,N_2296);
or UO_365 (O_365,N_2316,N_2102);
and UO_366 (O_366,N_2219,N_2050);
nor UO_367 (O_367,N_2556,N_2592);
and UO_368 (O_368,N_2967,N_2140);
nand UO_369 (O_369,N_2390,N_2942);
or UO_370 (O_370,N_2502,N_2950);
and UO_371 (O_371,N_2285,N_2427);
nand UO_372 (O_372,N_2578,N_2028);
xnor UO_373 (O_373,N_2530,N_2511);
xor UO_374 (O_374,N_2325,N_2999);
and UO_375 (O_375,N_2895,N_2253);
xor UO_376 (O_376,N_2486,N_2061);
xnor UO_377 (O_377,N_2461,N_2485);
nor UO_378 (O_378,N_2199,N_2534);
and UO_379 (O_379,N_2819,N_2838);
xnor UO_380 (O_380,N_2663,N_2362);
nor UO_381 (O_381,N_2021,N_2068);
or UO_382 (O_382,N_2349,N_2780);
nor UO_383 (O_383,N_2125,N_2658);
or UO_384 (O_384,N_2067,N_2441);
and UO_385 (O_385,N_2243,N_2935);
nand UO_386 (O_386,N_2174,N_2244);
and UO_387 (O_387,N_2693,N_2874);
and UO_388 (O_388,N_2342,N_2324);
xnor UO_389 (O_389,N_2581,N_2168);
or UO_390 (O_390,N_2741,N_2806);
nand UO_391 (O_391,N_2172,N_2288);
xnor UO_392 (O_392,N_2601,N_2448);
or UO_393 (O_393,N_2624,N_2186);
and UO_394 (O_394,N_2612,N_2619);
nor UO_395 (O_395,N_2076,N_2280);
and UO_396 (O_396,N_2907,N_2019);
xnor UO_397 (O_397,N_2732,N_2925);
nand UO_398 (O_398,N_2564,N_2525);
xor UO_399 (O_399,N_2470,N_2179);
nand UO_400 (O_400,N_2786,N_2011);
xor UO_401 (O_401,N_2674,N_2170);
and UO_402 (O_402,N_2081,N_2555);
nand UO_403 (O_403,N_2405,N_2370);
and UO_404 (O_404,N_2483,N_2154);
and UO_405 (O_405,N_2178,N_2792);
nand UO_406 (O_406,N_2212,N_2382);
nor UO_407 (O_407,N_2829,N_2929);
xnor UO_408 (O_408,N_2424,N_2223);
nor UO_409 (O_409,N_2715,N_2335);
nor UO_410 (O_410,N_2734,N_2692);
nand UO_411 (O_411,N_2748,N_2716);
nand UO_412 (O_412,N_2169,N_2431);
or UO_413 (O_413,N_2597,N_2444);
nor UO_414 (O_414,N_2920,N_2849);
and UO_415 (O_415,N_2492,N_2404);
or UO_416 (O_416,N_2392,N_2531);
nand UO_417 (O_417,N_2905,N_2480);
nor UO_418 (O_418,N_2112,N_2637);
xor UO_419 (O_419,N_2510,N_2206);
nor UO_420 (O_420,N_2438,N_2779);
nor UO_421 (O_421,N_2003,N_2611);
xor UO_422 (O_422,N_2707,N_2521);
nor UO_423 (O_423,N_2594,N_2009);
xnor UO_424 (O_424,N_2951,N_2162);
nor UO_425 (O_425,N_2603,N_2023);
xor UO_426 (O_426,N_2547,N_2954);
nor UO_427 (O_427,N_2177,N_2093);
and UO_428 (O_428,N_2816,N_2586);
and UO_429 (O_429,N_2888,N_2255);
xor UO_430 (O_430,N_2144,N_2338);
xor UO_431 (O_431,N_2884,N_2731);
or UO_432 (O_432,N_2239,N_2558);
nor UO_433 (O_433,N_2889,N_2489);
nor UO_434 (O_434,N_2416,N_2052);
nand UO_435 (O_435,N_2672,N_2964);
nor UO_436 (O_436,N_2029,N_2399);
xor UO_437 (O_437,N_2381,N_2132);
nor UO_438 (O_438,N_2839,N_2766);
xnor UO_439 (O_439,N_2350,N_2644);
xor UO_440 (O_440,N_2074,N_2012);
xor UO_441 (O_441,N_2949,N_2667);
or UO_442 (O_442,N_2610,N_2864);
nor UO_443 (O_443,N_2013,N_2843);
xor UO_444 (O_444,N_2690,N_2974);
xnor UO_445 (O_445,N_2014,N_2120);
nand UO_446 (O_446,N_2211,N_2216);
xor UO_447 (O_447,N_2934,N_2722);
or UO_448 (O_448,N_2962,N_2215);
nand UO_449 (O_449,N_2477,N_2745);
xor UO_450 (O_450,N_2613,N_2520);
nor UO_451 (O_451,N_2026,N_2729);
or UO_452 (O_452,N_2553,N_2805);
xnor UO_453 (O_453,N_2261,N_2848);
nor UO_454 (O_454,N_2501,N_2749);
and UO_455 (O_455,N_2788,N_2373);
and UO_456 (O_456,N_2765,N_2771);
nor UO_457 (O_457,N_2870,N_2953);
nor UO_458 (O_458,N_2499,N_2188);
or UO_459 (O_459,N_2615,N_2981);
and UO_460 (O_460,N_2585,N_2123);
nor UO_461 (O_461,N_2262,N_2545);
nor UO_462 (O_462,N_2078,N_2266);
nor UO_463 (O_463,N_2273,N_2200);
nand UO_464 (O_464,N_2522,N_2083);
nand UO_465 (O_465,N_2275,N_2000);
nor UO_466 (O_466,N_2523,N_2446);
nor UO_467 (O_467,N_2245,N_2051);
nand UO_468 (O_468,N_2882,N_2563);
xor UO_469 (O_469,N_2242,N_2795);
nor UO_470 (O_470,N_2095,N_2251);
and UO_471 (O_471,N_2773,N_2400);
and UO_472 (O_472,N_2114,N_2031);
or UO_473 (O_473,N_2720,N_2167);
nor UO_474 (O_474,N_2119,N_2460);
nand UO_475 (O_475,N_2118,N_2187);
xnor UO_476 (O_476,N_2433,N_2301);
nor UO_477 (O_477,N_2384,N_2683);
xnor UO_478 (O_478,N_2914,N_2678);
nand UO_479 (O_479,N_2127,N_2711);
xnor UO_480 (O_480,N_2294,N_2401);
nor UO_481 (O_481,N_2965,N_2656);
and UO_482 (O_482,N_2554,N_2279);
nand UO_483 (O_483,N_2956,N_2841);
nand UO_484 (O_484,N_2506,N_2329);
or UO_485 (O_485,N_2703,N_2091);
nor UO_486 (O_486,N_2359,N_2617);
nand UO_487 (O_487,N_2661,N_2573);
nor UO_488 (O_488,N_2628,N_2164);
xor UO_489 (O_489,N_2204,N_2600);
and UO_490 (O_490,N_2080,N_2302);
nor UO_491 (O_491,N_2367,N_2383);
nor UO_492 (O_492,N_2138,N_2930);
nand UO_493 (O_493,N_2512,N_2588);
or UO_494 (O_494,N_2375,N_2560);
xor UO_495 (O_495,N_2197,N_2826);
xnor UO_496 (O_496,N_2493,N_2034);
and UO_497 (O_497,N_2668,N_2334);
or UO_498 (O_498,N_2730,N_2145);
nor UO_499 (O_499,N_2820,N_2992);
endmodule