module basic_1500_15000_2000_30_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_1328,In_840);
nand U1 (N_1,In_784,In_1274);
xor U2 (N_2,In_523,In_879);
or U3 (N_3,In_1476,In_187);
nor U4 (N_4,In_668,In_172);
xnor U5 (N_5,In_468,In_634);
or U6 (N_6,In_803,In_522);
or U7 (N_7,In_831,In_949);
or U8 (N_8,In_46,In_916);
nor U9 (N_9,In_15,In_179);
and U10 (N_10,In_1109,In_779);
nand U11 (N_11,In_268,In_400);
or U12 (N_12,In_786,In_145);
nand U13 (N_13,In_78,In_1215);
or U14 (N_14,In_1056,In_847);
or U15 (N_15,In_1452,In_571);
or U16 (N_16,In_1140,In_550);
and U17 (N_17,In_177,In_533);
nor U18 (N_18,In_24,In_1120);
nand U19 (N_19,In_123,In_322);
or U20 (N_20,In_1379,In_1015);
nand U21 (N_21,In_469,In_1490);
and U22 (N_22,In_1323,In_333);
nor U23 (N_23,In_1045,In_501);
or U24 (N_24,In_301,In_981);
or U25 (N_25,In_1280,In_1017);
nand U26 (N_26,In_215,In_1421);
and U27 (N_27,In_247,In_1168);
and U28 (N_28,In_487,In_1129);
xnor U29 (N_29,In_845,In_1373);
nand U30 (N_30,In_167,In_355);
xor U31 (N_31,In_1308,In_676);
nor U32 (N_32,In_127,In_261);
nor U33 (N_33,In_1268,In_853);
xnor U34 (N_34,In_385,In_1239);
nor U35 (N_35,In_86,In_883);
or U36 (N_36,In_1447,In_687);
xor U37 (N_37,In_1019,In_296);
and U38 (N_38,In_628,In_1365);
and U39 (N_39,In_1428,In_673);
nor U40 (N_40,In_1333,In_1300);
nand U41 (N_41,In_595,In_1366);
and U42 (N_42,In_991,In_1223);
or U43 (N_43,In_808,In_1432);
or U44 (N_44,In_380,In_416);
or U45 (N_45,In_818,In_288);
xor U46 (N_46,In_648,In_625);
nand U47 (N_47,In_244,In_1153);
and U48 (N_48,In_781,In_14);
or U49 (N_49,In_180,In_450);
xnor U50 (N_50,In_1004,In_1309);
and U51 (N_51,In_498,In_516);
nand U52 (N_52,In_1184,In_1007);
nor U53 (N_53,In_229,In_1445);
xnor U54 (N_54,In_1479,In_914);
nor U55 (N_55,In_1195,In_844);
nor U56 (N_56,In_19,In_499);
and U57 (N_57,In_802,In_610);
nand U58 (N_58,In_1257,In_431);
and U59 (N_59,In_919,In_136);
xnor U60 (N_60,In_1123,In_1127);
nor U61 (N_61,In_164,In_699);
xnor U62 (N_62,In_969,In_940);
nand U63 (N_63,In_627,In_116);
and U64 (N_64,In_1104,In_1135);
nand U65 (N_65,In_639,In_49);
xor U66 (N_66,In_1318,In_1298);
xnor U67 (N_67,In_888,In_324);
and U68 (N_68,In_446,In_954);
and U69 (N_69,In_1466,In_335);
xor U70 (N_70,In_856,In_1495);
nand U71 (N_71,In_1464,In_758);
xnor U72 (N_72,In_681,In_151);
xor U73 (N_73,In_630,In_686);
and U74 (N_74,In_659,In_45);
and U75 (N_75,In_236,In_135);
nand U76 (N_76,In_1355,In_67);
or U77 (N_77,In_715,In_1117);
or U78 (N_78,In_478,In_1065);
or U79 (N_79,In_1097,In_1075);
xnor U80 (N_80,In_1000,In_319);
and U81 (N_81,In_430,In_1241);
or U82 (N_82,In_1414,In_1210);
and U83 (N_83,In_437,In_619);
or U84 (N_84,In_100,In_1211);
and U85 (N_85,In_1069,In_71);
nand U86 (N_86,In_16,In_740);
and U87 (N_87,In_68,In_99);
nor U88 (N_88,In_226,In_887);
or U89 (N_89,In_444,In_664);
nor U90 (N_90,In_337,In_702);
nand U91 (N_91,In_299,In_884);
nand U92 (N_92,In_944,In_1270);
xor U93 (N_93,In_436,In_350);
xnor U94 (N_94,In_776,In_1437);
nand U95 (N_95,In_742,In_959);
and U96 (N_96,In_536,In_508);
or U97 (N_97,In_1392,In_1119);
xor U98 (N_98,In_833,In_390);
xor U99 (N_99,In_730,In_413);
and U100 (N_100,In_1102,In_225);
xor U101 (N_101,In_817,In_530);
xnor U102 (N_102,In_519,In_667);
xor U103 (N_103,In_1040,In_1249);
nand U104 (N_104,In_1025,In_1058);
or U105 (N_105,In_472,In_724);
nor U106 (N_106,In_1059,In_1108);
xnor U107 (N_107,In_621,In_352);
or U108 (N_108,In_834,In_1337);
and U109 (N_109,In_913,In_370);
nand U110 (N_110,In_1219,In_609);
or U111 (N_111,In_889,In_1410);
nor U112 (N_112,In_1407,In_344);
or U113 (N_113,In_541,In_585);
nor U114 (N_114,In_706,In_555);
and U115 (N_115,In_209,In_1090);
nor U116 (N_116,In_242,In_25);
nand U117 (N_117,In_1380,In_566);
nor U118 (N_118,In_580,In_662);
xor U119 (N_119,In_1386,In_12);
nor U120 (N_120,In_457,In_1188);
or U121 (N_121,In_799,In_1431);
nor U122 (N_122,In_1424,In_691);
or U123 (N_123,In_233,In_1443);
nand U124 (N_124,In_783,In_1078);
nor U125 (N_125,In_666,In_63);
xnor U126 (N_126,In_657,In_421);
xnor U127 (N_127,In_1442,In_1107);
xor U128 (N_128,In_462,In_864);
nor U129 (N_129,In_81,In_1246);
or U130 (N_130,In_1465,In_900);
nand U131 (N_131,In_18,In_700);
nor U132 (N_132,In_1046,In_604);
nor U133 (N_133,In_956,In_763);
or U134 (N_134,In_1357,In_1294);
xor U135 (N_135,In_429,In_1041);
and U136 (N_136,In_892,In_1038);
nand U137 (N_137,In_440,In_138);
nand U138 (N_138,In_434,In_197);
nor U139 (N_139,In_745,In_235);
nor U140 (N_140,In_321,In_1167);
or U141 (N_141,In_140,In_683);
nor U142 (N_142,In_378,In_1259);
and U143 (N_143,In_17,In_106);
xor U144 (N_144,In_152,In_1279);
or U145 (N_145,In_1451,In_198);
nor U146 (N_146,In_906,In_95);
or U147 (N_147,In_1174,In_1060);
xor U148 (N_148,In_511,In_341);
nor U149 (N_149,In_547,In_616);
or U150 (N_150,In_111,In_347);
xor U151 (N_151,In_294,In_682);
and U152 (N_152,In_79,In_719);
nand U153 (N_153,In_471,In_1194);
nor U154 (N_154,In_219,In_22);
nand U155 (N_155,In_159,In_1454);
and U156 (N_156,In_35,In_32);
and U157 (N_157,In_1096,In_1179);
or U158 (N_158,In_953,In_617);
or U159 (N_159,In_1177,In_583);
and U160 (N_160,In_506,In_897);
nand U161 (N_161,In_1367,In_176);
nand U162 (N_162,In_531,In_274);
and U163 (N_163,In_114,In_539);
nand U164 (N_164,In_553,In_175);
nand U165 (N_165,In_31,In_206);
nor U166 (N_166,In_192,In_6);
nor U167 (N_167,In_1020,In_1498);
nand U168 (N_168,In_144,In_510);
xor U169 (N_169,In_388,In_286);
or U170 (N_170,In_939,In_637);
xor U171 (N_171,In_449,In_1332);
and U172 (N_172,In_185,In_690);
and U173 (N_173,In_479,In_493);
or U174 (N_174,In_1487,In_977);
xor U175 (N_175,In_356,In_992);
or U176 (N_176,In_357,In_1307);
xor U177 (N_177,In_854,In_788);
xor U178 (N_178,In_351,In_757);
nor U179 (N_179,In_955,In_354);
nor U180 (N_180,In_607,In_366);
or U181 (N_181,In_653,In_1461);
xnor U182 (N_182,In_406,In_985);
xnor U183 (N_183,In_1245,In_826);
and U184 (N_184,In_820,In_317);
nor U185 (N_185,In_1106,In_393);
and U186 (N_186,In_982,In_1310);
or U187 (N_187,In_423,In_732);
or U188 (N_188,In_570,In_142);
or U189 (N_189,In_1183,In_477);
nand U190 (N_190,In_797,In_1304);
xnor U191 (N_191,In_1349,In_386);
or U192 (N_192,In_780,In_1230);
and U193 (N_193,In_139,In_517);
nor U194 (N_194,In_401,In_558);
xnor U195 (N_195,In_832,In_133);
xor U196 (N_196,In_920,In_929);
and U197 (N_197,In_318,In_1111);
nor U198 (N_198,In_761,In_573);
and U199 (N_199,In_293,In_1295);
xnor U200 (N_200,In_183,In_1289);
xnor U201 (N_201,In_451,In_191);
nand U202 (N_202,In_254,In_1228);
xnor U203 (N_203,In_1481,In_647);
and U204 (N_204,In_372,In_942);
and U205 (N_205,In_149,In_208);
xnor U206 (N_206,In_320,In_1484);
nor U207 (N_207,In_1012,In_1399);
or U208 (N_208,In_1271,In_747);
or U209 (N_209,In_464,In_638);
and U210 (N_210,In_1095,In_103);
nor U211 (N_211,In_1101,In_769);
nand U212 (N_212,In_1287,In_407);
xor U213 (N_213,In_194,In_885);
or U214 (N_214,In_1057,In_489);
or U215 (N_215,In_435,In_199);
and U216 (N_216,In_162,In_1358);
or U217 (N_217,In_614,In_1197);
nor U218 (N_218,In_262,In_1166);
or U219 (N_219,In_1079,In_264);
nand U220 (N_220,In_1218,In_611);
or U221 (N_221,In_85,In_636);
or U222 (N_222,In_184,In_1263);
or U223 (N_223,In_37,In_886);
or U224 (N_224,In_727,In_1133);
nand U225 (N_225,In_1455,In_394);
or U226 (N_226,In_520,In_87);
or U227 (N_227,In_782,In_692);
nor U228 (N_228,In_160,In_39);
nor U229 (N_229,In_1149,In_326);
or U230 (N_230,In_824,In_1022);
nor U231 (N_231,In_1378,In_560);
xnor U232 (N_232,In_258,In_101);
and U233 (N_233,In_349,In_482);
or U234 (N_234,In_38,In_663);
and U235 (N_235,In_260,In_640);
and U236 (N_236,In_36,In_369);
xnor U237 (N_237,In_1477,In_922);
and U238 (N_238,In_30,In_214);
nor U239 (N_239,In_269,In_1496);
nand U240 (N_240,In_485,In_1336);
xnor U241 (N_241,In_1003,In_1313);
and U242 (N_242,In_1440,In_1048);
or U243 (N_243,In_1103,In_302);
nand U244 (N_244,In_1269,In_1209);
xor U245 (N_245,In_383,In_1013);
and U246 (N_246,In_1302,In_410);
nor U247 (N_247,In_716,In_1350);
and U248 (N_248,In_649,In_1084);
or U249 (N_249,In_1347,In_1311);
nor U250 (N_250,In_713,In_396);
and U251 (N_251,In_361,In_694);
xnor U252 (N_252,In_1391,In_1147);
nor U253 (N_253,In_1225,In_1284);
or U254 (N_254,In_173,In_1217);
xor U255 (N_255,In_60,In_213);
xor U256 (N_256,In_1468,In_44);
and U257 (N_257,In_597,In_1160);
xnor U258 (N_258,In_1023,In_1081);
nand U259 (N_259,In_973,In_509);
or U260 (N_260,In_976,In_749);
or U261 (N_261,In_1400,In_1460);
nor U262 (N_262,In_11,In_928);
nand U263 (N_263,In_10,In_122);
nor U264 (N_264,In_529,In_823);
xor U265 (N_265,In_454,In_1467);
and U266 (N_266,In_807,In_1352);
and U267 (N_267,In_143,In_1044);
or U268 (N_268,In_91,In_868);
and U269 (N_269,In_552,In_96);
nor U270 (N_270,In_186,In_654);
xnor U271 (N_271,In_670,In_1199);
or U272 (N_272,In_927,In_1143);
nand U273 (N_273,In_353,In_339);
nor U274 (N_274,In_532,In_384);
nand U275 (N_275,In_721,In_626);
nor U276 (N_276,In_104,In_1193);
or U277 (N_277,In_2,In_1049);
or U278 (N_278,In_909,In_739);
nand U279 (N_279,In_480,In_701);
or U280 (N_280,In_809,In_871);
or U281 (N_281,In_934,In_829);
nand U282 (N_282,In_1180,In_841);
xor U283 (N_283,In_112,In_1073);
nand U284 (N_284,In_1248,In_765);
nor U285 (N_285,In_182,In_825);
nand U286 (N_286,In_72,In_608);
xor U287 (N_287,In_925,In_723);
and U288 (N_288,In_651,In_1381);
nor U289 (N_289,In_1029,In_13);
or U290 (N_290,In_857,In_1255);
xnor U291 (N_291,In_789,In_582);
and U292 (N_292,In_1375,In_243);
nand U293 (N_293,In_1213,In_641);
nand U294 (N_294,In_455,In_750);
or U295 (N_295,In_1141,In_805);
nor U296 (N_296,In_381,In_731);
or U297 (N_297,In_1165,In_1283);
xor U298 (N_298,In_108,In_1173);
nor U299 (N_299,In_1207,In_671);
nor U300 (N_300,In_911,In_212);
and U301 (N_301,In_924,In_964);
nor U302 (N_302,In_849,In_1137);
xor U303 (N_303,In_1439,In_785);
nor U304 (N_304,In_1190,In_195);
nor U305 (N_305,In_564,In_631);
nor U306 (N_306,In_814,In_1475);
and U307 (N_307,In_432,In_166);
and U308 (N_308,In_605,In_848);
nor U309 (N_309,In_346,In_1384);
xor U310 (N_310,In_500,In_1053);
nand U311 (N_311,In_207,In_252);
xor U312 (N_312,In_722,In_827);
nand U313 (N_313,In_507,In_73);
nand U314 (N_314,In_880,In_1462);
nand U315 (N_315,In_1260,In_309);
nor U316 (N_316,In_1456,In_586);
xor U317 (N_317,In_496,In_1343);
nor U318 (N_318,In_157,In_1372);
nor U319 (N_319,In_1068,In_752);
nor U320 (N_320,In_930,In_873);
xor U321 (N_321,In_562,In_579);
or U322 (N_322,In_970,In_433);
xnor U323 (N_323,In_395,In_837);
and U324 (N_324,In_946,In_698);
nor U325 (N_325,In_375,In_592);
nor U326 (N_326,In_74,In_9);
xnor U327 (N_327,In_1390,In_1155);
or U328 (N_328,In_987,In_1159);
xnor U329 (N_329,In_1321,In_1401);
and U330 (N_330,In_994,In_1089);
nand U331 (N_331,In_494,In_755);
nand U332 (N_332,In_306,In_1009);
and U333 (N_333,In_1021,In_340);
nor U334 (N_334,In_148,In_484);
or U335 (N_335,In_502,In_1377);
xnor U336 (N_336,In_130,In_165);
xor U337 (N_337,In_310,In_1277);
nand U338 (N_338,In_876,In_734);
or U339 (N_339,In_1113,In_34);
and U340 (N_340,In_1224,In_1396);
nor U341 (N_341,In_1222,In_204);
and U342 (N_342,In_115,In_672);
xnor U343 (N_343,In_210,In_271);
and U344 (N_344,In_422,In_655);
xnor U345 (N_345,In_224,In_917);
xor U346 (N_346,In_330,In_404);
xor U347 (N_347,In_538,In_861);
and U348 (N_348,In_975,In_891);
nand U349 (N_349,In_445,In_1290);
nor U350 (N_350,In_624,In_910);
and U351 (N_351,In_1315,In_1264);
nand U352 (N_352,In_1331,In_128);
nand U353 (N_353,In_325,In_1132);
or U354 (N_354,In_1154,In_141);
nor U355 (N_355,In_870,In_417);
xor U356 (N_356,In_951,In_1419);
xor U357 (N_357,In_53,In_1244);
nand U358 (N_358,In_576,In_69);
or U359 (N_359,In_367,In_869);
or U360 (N_360,In_979,In_1116);
nand U361 (N_361,In_1463,In_1438);
nand U362 (N_362,In_1175,In_1250);
or U363 (N_363,In_1327,In_461);
nor U364 (N_364,In_1433,In_613);
nand U365 (N_365,In_312,In_1156);
and U366 (N_366,In_427,In_491);
and U367 (N_367,In_901,In_1136);
or U368 (N_368,In_315,In_908);
nor U369 (N_369,In_684,In_1319);
nor U370 (N_370,In_622,In_915);
and U371 (N_371,In_912,In_1397);
or U372 (N_372,In_232,In_736);
xor U373 (N_373,In_1145,In_392);
nor U374 (N_374,In_1157,In_158);
xor U375 (N_375,In_292,In_1043);
nor U376 (N_376,In_447,In_1243);
nand U377 (N_377,In_744,In_80);
nand U378 (N_378,In_524,In_1083);
nand U379 (N_379,In_1240,In_316);
and U380 (N_380,In_1125,In_1028);
nand U381 (N_381,In_360,In_589);
nor U382 (N_382,In_540,In_862);
xor U383 (N_383,In_600,In_549);
and U384 (N_384,In_903,In_1221);
and U385 (N_385,In_238,In_481);
nor U386 (N_386,In_515,In_796);
nand U387 (N_387,In_1130,In_720);
xnor U388 (N_388,In_1389,In_283);
and U389 (N_389,In_1296,In_448);
and U390 (N_390,In_1364,In_473);
nor U391 (N_391,In_1356,In_52);
and U392 (N_392,In_1033,In_850);
nand U393 (N_393,In_1212,In_1131);
nor U394 (N_394,In_303,In_777);
xnor U395 (N_395,In_860,In_1473);
xor U396 (N_396,In_893,In_882);
or U397 (N_397,In_277,In_932);
or U398 (N_398,In_1429,In_554);
or U399 (N_399,In_710,In_984);
nor U400 (N_400,In_1338,In_428);
nor U401 (N_401,In_1371,In_1158);
xor U402 (N_402,In_534,In_40);
and U403 (N_403,In_787,In_504);
xor U404 (N_404,In_41,In_767);
nand U405 (N_405,In_525,In_93);
nor U406 (N_406,In_962,In_822);
or U407 (N_407,In_1374,In_615);
and U408 (N_408,In_1247,In_801);
nand U409 (N_409,In_201,In_1);
xnor U410 (N_410,In_960,In_1359);
xnor U411 (N_411,In_373,In_153);
and U412 (N_412,In_1469,In_669);
nor U413 (N_413,In_1176,In_568);
or U414 (N_414,In_1093,In_697);
or U415 (N_415,In_334,In_821);
or U416 (N_416,In_1128,In_1031);
and U417 (N_417,In_181,In_311);
nor U418 (N_418,In_459,In_280);
nor U419 (N_419,In_544,In_239);
or U420 (N_420,In_1070,In_535);
nand U421 (N_421,In_526,In_1326);
nand U422 (N_422,In_1288,In_76);
and U423 (N_423,In_923,In_1071);
and U424 (N_424,In_399,In_688);
or U425 (N_425,In_50,In_1172);
xor U426 (N_426,In_1235,In_774);
xnor U427 (N_427,In_1146,In_1192);
or U428 (N_428,In_947,In_329);
or U429 (N_429,In_442,In_1353);
nand U430 (N_430,In_1420,In_1423);
or U431 (N_431,In_168,In_33);
or U432 (N_432,In_936,In_989);
nand U433 (N_433,In_1320,In_986);
and U434 (N_434,In_418,In_387);
xor U435 (N_435,In_476,In_270);
or U436 (N_436,In_1472,In_307);
xor U437 (N_437,In_878,In_368);
nor U438 (N_438,In_1351,In_933);
and U439 (N_439,In_1492,In_756);
nand U440 (N_440,In_743,In_574);
and U441 (N_441,In_1178,In_1348);
nor U442 (N_442,In_1360,In_557);
and U443 (N_443,In_545,In_497);
xnor U444 (N_444,In_1430,In_1301);
nand U445 (N_445,In_1297,In_575);
and U446 (N_446,In_193,In_1030);
nand U447 (N_447,In_147,In_810);
and U448 (N_448,In_1398,In_798);
nand U449 (N_449,In_266,In_1187);
and U450 (N_450,In_1066,In_997);
nand U451 (N_451,In_1453,In_463);
xor U452 (N_452,In_1449,In_1272);
xnor U453 (N_453,In_772,In_867);
xor U454 (N_454,In_543,In_304);
or U455 (N_455,In_741,In_1227);
nand U456 (N_456,In_1216,In_1231);
xnor U457 (N_457,In_1110,In_775);
nor U458 (N_458,In_415,In_397);
nor U459 (N_459,In_1482,In_1434);
nand U460 (N_460,In_189,In_20);
nor U461 (N_461,In_800,In_1010);
xor U462 (N_462,In_190,In_28);
xnor U463 (N_463,In_1275,In_7);
nor U464 (N_464,In_146,In_305);
or U465 (N_465,In_918,In_289);
nand U466 (N_466,In_119,In_4);
xnor U467 (N_467,In_1121,In_92);
nor U468 (N_468,In_762,In_1491);
nor U469 (N_469,In_978,In_726);
nor U470 (N_470,In_456,In_1170);
xor U471 (N_471,In_332,In_999);
nand U472 (N_472,In_1324,In_1416);
nand U473 (N_473,In_980,In_218);
xnor U474 (N_474,In_1312,In_1150);
nor U475 (N_475,In_1316,In_899);
nand U476 (N_476,In_1061,In_972);
xnor U477 (N_477,In_419,In_342);
nor U478 (N_478,In_278,In_963);
nand U479 (N_479,In_488,In_877);
and U480 (N_480,In_313,In_279);
nand U481 (N_481,In_561,In_109);
and U482 (N_482,In_1444,In_1205);
and U483 (N_483,In_656,In_1036);
nand U484 (N_484,In_113,In_735);
or U485 (N_485,In_0,In_223);
and U486 (N_486,In_1018,In_1005);
or U487 (N_487,In_569,In_169);
xnor U488 (N_488,In_843,In_374);
nor U489 (N_489,In_746,In_1064);
or U490 (N_490,In_1092,In_1417);
nor U491 (N_491,In_411,In_248);
or U492 (N_492,In_1011,In_503);
or U493 (N_493,In_88,In_54);
and U494 (N_494,In_931,In_1427);
and U495 (N_495,In_1474,In_161);
nand U496 (N_496,In_290,In_217);
and U497 (N_497,In_521,In_581);
or U498 (N_498,In_263,In_1426);
nor U499 (N_499,In_257,In_993);
or U500 (N_500,N_135,N_448);
or U501 (N_501,N_157,In_358);
nand U502 (N_502,N_359,In_1067);
nand U503 (N_503,N_147,In_567);
xor U504 (N_504,N_48,N_211);
and U505 (N_505,In_1206,N_123);
xor U506 (N_506,In_338,In_644);
nand U507 (N_507,N_215,N_119);
nand U508 (N_508,N_33,In_793);
nand U509 (N_509,N_216,N_457);
nor U510 (N_510,N_291,In_811);
and U511 (N_511,N_323,N_49);
xnor U512 (N_512,In_974,N_469);
or U513 (N_513,In_842,In_895);
nor U514 (N_514,In_1138,N_242);
or U515 (N_515,N_451,In_1139);
nor U516 (N_516,In_629,In_1220);
and U517 (N_517,In_1334,In_791);
nand U518 (N_518,In_563,N_441);
nand U519 (N_519,N_414,N_127);
xor U520 (N_520,N_459,N_42);
xnor U521 (N_521,In_1285,N_381);
and U522 (N_522,In_200,N_256);
nor U523 (N_523,In_905,N_271);
xnor U524 (N_524,In_466,N_50);
nand U525 (N_525,In_1411,N_91);
xor U526 (N_526,In_677,N_496);
xnor U527 (N_527,N_204,In_62);
nor U528 (N_528,N_185,In_265);
nor U529 (N_529,N_177,N_103);
or U530 (N_530,In_297,In_1171);
nor U531 (N_531,N_149,N_394);
xor U532 (N_532,In_1362,N_83);
xor U533 (N_533,In_1387,In_425);
nor U534 (N_534,In_707,N_345);
nor U535 (N_535,N_140,N_253);
nand U536 (N_536,N_387,N_112);
nor U537 (N_537,N_27,In_1485);
nand U538 (N_538,In_1457,In_556);
nand U539 (N_539,N_89,N_415);
or U540 (N_540,In_117,N_11);
and U541 (N_541,In_1185,In_124);
nor U542 (N_542,N_467,N_221);
xnor U543 (N_543,In_587,In_737);
or U544 (N_544,In_966,In_1370);
and U545 (N_545,In_904,N_445);
nand U546 (N_546,N_470,N_406);
and U547 (N_547,In_661,N_330);
xor U548 (N_548,N_110,In_1499);
nand U549 (N_549,N_118,N_13);
and U550 (N_550,In_1261,N_229);
nand U551 (N_551,N_363,In_1415);
or U552 (N_552,In_548,In_58);
nor U553 (N_553,In_542,N_258);
or U554 (N_554,N_172,N_455);
and U555 (N_555,N_134,In_336);
and U556 (N_556,N_380,N_499);
nand U557 (N_557,In_1346,N_405);
or U558 (N_558,N_125,In_518);
and U559 (N_559,N_4,In_241);
and U560 (N_560,N_92,N_230);
xor U561 (N_561,N_41,In_696);
or U562 (N_562,In_1342,In_1385);
nor U563 (N_563,N_106,In_29);
xnor U564 (N_564,N_14,In_118);
xor U565 (N_565,N_326,N_393);
nor U566 (N_566,N_338,N_122);
xor U567 (N_567,N_306,In_1203);
nand U568 (N_568,N_109,N_250);
or U569 (N_569,In_1403,In_1299);
nor U570 (N_570,In_1422,N_183);
and U571 (N_571,N_12,N_244);
nor U572 (N_572,N_438,N_284);
and U573 (N_573,In_458,N_153);
or U574 (N_574,In_121,In_389);
xor U575 (N_575,N_37,N_66);
nor U576 (N_576,In_483,N_174);
and U577 (N_577,In_1425,In_298);
nor U578 (N_578,In_588,In_1253);
and U579 (N_579,N_43,In_836);
nand U580 (N_580,In_1238,N_289);
xor U581 (N_581,N_161,N_146);
and U582 (N_582,N_166,In_645);
nand U583 (N_583,N_428,N_235);
or U584 (N_584,In_1281,N_464);
nand U585 (N_585,N_293,In_1470);
nor U586 (N_586,In_1483,In_1267);
xor U587 (N_587,N_320,N_360);
nand U588 (N_588,In_1008,In_211);
xor U589 (N_589,N_386,N_64);
xnor U590 (N_590,In_363,In_1329);
or U591 (N_591,In_1098,In_131);
nor U592 (N_592,N_170,N_70);
nor U593 (N_593,N_18,In_70);
and U594 (N_594,In_898,N_167);
nand U595 (N_595,In_231,In_359);
xnor U596 (N_596,In_1152,N_44);
nand U597 (N_597,In_259,N_236);
and U598 (N_598,N_26,N_28);
or U599 (N_599,N_180,N_302);
nor U600 (N_600,N_139,In_1306);
and U601 (N_601,N_126,In_1214);
nand U602 (N_602,N_19,N_347);
nand U603 (N_603,In_474,N_483);
xnor U604 (N_604,In_1042,N_87);
nor U605 (N_605,In_1002,In_968);
nor U606 (N_606,N_20,N_1);
nand U607 (N_607,In_623,N_102);
nor U608 (N_608,In_577,In_82);
xnor U609 (N_609,N_56,N_62);
or U610 (N_610,N_407,In_601);
nor U611 (N_611,In_21,N_181);
xor U612 (N_612,In_1494,N_288);
or U613 (N_613,N_389,N_382);
or U614 (N_614,N_340,In_606);
nand U615 (N_615,In_403,In_234);
nand U616 (N_616,In_228,N_362);
nor U617 (N_617,N_245,N_6);
or U618 (N_618,N_417,In_405);
or U619 (N_619,N_485,In_512);
and U620 (N_620,In_1237,In_203);
and U621 (N_621,N_247,N_154);
and U622 (N_622,N_159,N_369);
nand U623 (N_623,N_53,N_301);
nand U624 (N_624,In_1402,In_1161);
and U625 (N_625,N_398,In_1014);
and U626 (N_626,In_1072,N_397);
or U627 (N_627,N_280,N_329);
nor U628 (N_628,In_102,N_60);
and U629 (N_629,In_163,N_67);
nand U630 (N_630,In_751,In_938);
or U631 (N_631,In_343,N_333);
xor U632 (N_632,In_1181,N_379);
or U633 (N_633,In_983,N_138);
nand U634 (N_634,In_245,In_1493);
and U635 (N_635,In_1282,N_79);
nand U636 (N_636,N_189,N_55);
nor U637 (N_637,In_1361,In_1345);
or U638 (N_638,N_32,N_47);
nand U639 (N_639,In_1035,In_1016);
nand U640 (N_640,In_216,In_1144);
and U641 (N_641,In_894,In_1488);
nor U642 (N_642,In_1050,In_250);
xor U643 (N_643,N_163,N_342);
nand U644 (N_644,N_274,N_85);
and U645 (N_645,N_173,In_196);
and U646 (N_646,N_498,N_155);
or U647 (N_647,In_1047,In_345);
or U648 (N_648,N_478,N_208);
and U649 (N_649,N_410,N_156);
or U650 (N_650,N_282,N_439);
nor U651 (N_651,In_439,In_246);
nor U652 (N_652,In_134,N_465);
and U653 (N_653,N_287,N_21);
and U654 (N_654,In_1085,N_300);
and U655 (N_655,In_1292,N_132);
nand U656 (N_656,In_3,N_486);
nor U657 (N_657,N_218,In_132);
nor U658 (N_658,In_107,In_988);
and U659 (N_659,In_753,N_425);
nand U660 (N_660,N_371,N_105);
nor U661 (N_661,In_1063,In_441);
xnor U662 (N_662,In_650,In_813);
nor U663 (N_663,In_1006,N_420);
xor U664 (N_664,In_1191,In_584);
xor U665 (N_665,In_221,In_795);
xor U666 (N_666,N_482,N_81);
nor U667 (N_667,N_76,N_190);
nand U668 (N_668,N_375,N_372);
and U669 (N_669,N_401,In_729);
nor U670 (N_670,N_331,In_1458);
nor U671 (N_671,N_137,In_537);
or U672 (N_672,N_224,N_436);
nor U673 (N_673,In_907,In_748);
nand U674 (N_674,In_1489,In_790);
or U675 (N_675,N_351,In_865);
or U676 (N_676,In_945,N_99);
nor U677 (N_677,N_220,In_1162);
or U678 (N_678,In_327,N_294);
and U679 (N_679,In_1001,N_490);
xor U680 (N_680,N_194,N_238);
or U681 (N_681,In_551,N_309);
xor U682 (N_682,In_770,In_851);
xor U683 (N_683,In_890,In_866);
or U684 (N_684,N_310,N_57);
nor U685 (N_685,In_48,N_481);
nand U686 (N_686,In_1368,In_643);
nor U687 (N_687,N_249,In_61);
nor U688 (N_688,In_1262,N_261);
and U689 (N_689,In_412,N_395);
nand U690 (N_690,In_712,N_136);
nor U691 (N_691,In_314,N_113);
nor U692 (N_692,N_61,In_495);
or U693 (N_693,In_1266,N_477);
or U694 (N_694,N_148,In_1142);
or U695 (N_695,In_156,In_1305);
nor U696 (N_696,In_1406,N_327);
nor U697 (N_697,N_115,In_300);
and U698 (N_698,In_1435,In_858);
xor U699 (N_699,In_1409,N_357);
xor U700 (N_700,In_1446,In_1340);
nand U701 (N_701,In_759,In_1151);
or U702 (N_702,In_1062,N_328);
nor U703 (N_703,In_594,N_350);
nor U704 (N_704,N_101,In_733);
nor U705 (N_705,In_1204,N_52);
or U706 (N_706,In_1393,In_1105);
nor U707 (N_707,N_108,N_346);
and U708 (N_708,N_403,In_1256);
xor U709 (N_709,N_267,N_197);
or U710 (N_710,In_952,In_819);
xor U711 (N_711,N_78,N_210);
or U712 (N_712,N_332,In_1436);
nand U713 (N_713,N_39,In_703);
or U714 (N_714,N_266,In_408);
and U715 (N_715,N_268,In_1232);
and U716 (N_716,In_282,N_175);
nand U717 (N_717,N_36,In_1091);
and U718 (N_718,In_675,In_1325);
and U719 (N_719,In_680,N_217);
nand U720 (N_720,N_370,N_281);
nor U721 (N_721,N_241,N_374);
xnor U722 (N_722,In_815,In_635);
and U723 (N_723,N_297,In_859);
nor U724 (N_724,In_1341,In_1254);
nand U725 (N_725,In_838,N_143);
xor U726 (N_726,In_578,In_1229);
nor U727 (N_727,In_275,In_513);
xor U728 (N_728,N_171,N_24);
nor U729 (N_729,In_620,In_708);
and U730 (N_730,N_484,In_365);
and U731 (N_731,In_75,N_358);
and U732 (N_732,In_1265,In_1322);
nand U733 (N_733,N_295,N_120);
and U734 (N_734,N_23,In_618);
nor U735 (N_735,In_971,In_943);
xnor U736 (N_736,In_1118,In_1027);
or U737 (N_737,In_1497,In_709);
nand U738 (N_738,In_295,N_22);
nor U739 (N_739,N_226,In_658);
xnor U740 (N_740,N_116,In_26);
or U741 (N_741,N_124,In_794);
or U742 (N_742,In_59,In_65);
nand U743 (N_743,N_203,N_128);
and U744 (N_744,In_1037,In_222);
and U745 (N_745,N_45,N_196);
and U746 (N_746,In_1286,N_237);
nor U747 (N_747,N_259,N_463);
and U748 (N_748,In_828,In_990);
nand U749 (N_749,In_711,In_633);
nand U750 (N_750,N_141,N_466);
nand U751 (N_751,In_1376,In_528);
xnor U752 (N_752,In_527,N_305);
xor U753 (N_753,In_371,N_334);
nor U754 (N_754,N_65,In_764);
nor U755 (N_755,In_760,N_58);
nand U756 (N_756,In_646,In_1074);
nand U757 (N_757,N_497,In_806);
and U758 (N_758,N_77,In_240);
nand U759 (N_759,N_354,In_665);
or U760 (N_760,In_1405,N_388);
or U761 (N_761,In_1388,N_82);
or U762 (N_762,In_695,N_319);
and U763 (N_763,N_400,N_292);
and U764 (N_764,N_456,N_367);
nand U765 (N_765,N_107,In_679);
and U766 (N_766,N_431,N_355);
nor U767 (N_767,N_460,In_1382);
or U768 (N_768,In_255,N_46);
or U769 (N_769,In_1236,In_1413);
and U770 (N_770,In_1099,N_254);
and U771 (N_771,N_7,In_714);
and U772 (N_772,N_435,In_725);
nor U773 (N_773,In_704,N_225);
or U774 (N_774,In_284,N_260);
nor U775 (N_775,N_494,In_1088);
nor U776 (N_776,In_839,In_23);
and U777 (N_777,In_1076,N_493);
or U778 (N_778,N_151,N_152);
or U779 (N_779,In_438,In_178);
nand U780 (N_780,In_1189,In_1087);
xor U781 (N_781,In_771,N_145);
nor U782 (N_782,In_402,In_43);
nor U783 (N_783,In_593,In_475);
nand U784 (N_784,N_495,N_480);
and U785 (N_785,N_476,N_142);
xor U786 (N_786,In_1234,In_174);
nand U787 (N_787,N_239,N_184);
xor U788 (N_788,In_230,N_73);
or U789 (N_789,N_344,In_1242);
and U790 (N_790,N_192,In_467);
nor U791 (N_791,N_71,N_337);
xor U792 (N_792,In_120,N_449);
and U793 (N_793,In_1122,In_612);
xnor U794 (N_794,N_392,In_1052);
or U795 (N_795,N_205,In_603);
and U796 (N_796,N_276,N_100);
nand U797 (N_797,In_902,N_2);
nand U798 (N_798,In_935,In_678);
xnor U799 (N_799,In_995,In_97);
nand U800 (N_800,N_453,N_117);
nor U801 (N_801,N_385,N_90);
nand U802 (N_802,N_98,In_188);
xor U803 (N_803,N_424,N_30);
nand U804 (N_804,In_728,In_486);
and U805 (N_805,In_256,N_265);
xor U806 (N_806,In_89,In_599);
nand U807 (N_807,In_409,In_546);
nand U808 (N_808,In_693,N_270);
nand U809 (N_809,N_31,In_514);
xor U810 (N_810,N_29,In_1100);
xnor U811 (N_811,N_418,N_423);
or U812 (N_812,N_212,N_227);
or U813 (N_813,N_437,N_214);
xor U814 (N_814,N_5,In_596);
xnor U815 (N_815,In_426,N_182);
nor U816 (N_816,In_1186,In_129);
and U817 (N_817,N_315,N_487);
nor U818 (N_818,In_738,N_233);
or U819 (N_819,N_251,In_874);
or U820 (N_820,In_1480,N_468);
and U821 (N_821,In_1354,In_961);
or U822 (N_822,In_642,N_144);
xor U823 (N_823,N_352,N_409);
or U824 (N_824,N_366,N_433);
or U825 (N_825,N_207,N_391);
nor U826 (N_826,In_205,N_133);
and U827 (N_827,N_187,N_243);
nor U828 (N_828,In_285,N_75);
nor U829 (N_829,N_429,N_343);
nor U830 (N_830,In_251,N_176);
and U831 (N_831,In_377,N_307);
and U832 (N_832,N_452,N_234);
nor U833 (N_833,N_191,In_1112);
xnor U834 (N_834,N_25,N_322);
nor U835 (N_835,In_674,N_336);
nand U836 (N_836,In_926,N_0);
or U837 (N_837,In_56,N_34);
nor U838 (N_838,N_447,N_69);
nor U839 (N_839,In_1339,In_328);
nor U840 (N_840,In_1200,In_1363);
and U841 (N_841,N_262,In_364);
and U842 (N_842,In_1026,N_454);
and U843 (N_843,N_443,N_198);
nor U844 (N_844,In_1251,In_998);
nand U845 (N_845,In_652,In_872);
nand U846 (N_846,In_855,N_419);
nor U847 (N_847,In_950,N_199);
nand U848 (N_848,In_1459,N_492);
and U849 (N_849,N_72,N_427);
or U850 (N_850,N_219,In_1164);
and U851 (N_851,In_5,N_150);
nand U852 (N_852,In_1115,N_179);
nor U853 (N_853,N_240,In_1032);
xnor U854 (N_854,In_420,N_164);
xor U855 (N_855,N_416,In_424);
or U856 (N_856,In_1034,In_937);
xor U857 (N_857,N_93,N_373);
nand U858 (N_858,In_465,N_277);
nand U859 (N_859,In_1182,N_222);
nand U860 (N_860,In_1412,N_279);
or U861 (N_861,In_812,In_559);
xnor U862 (N_862,N_376,In_598);
nand U863 (N_863,In_272,In_1330);
nand U864 (N_864,In_778,In_391);
and U865 (N_865,In_754,N_38);
or U866 (N_866,N_361,N_68);
xnor U867 (N_867,N_168,In_1024);
xor U868 (N_868,In_94,In_27);
xnor U869 (N_869,In_1486,N_84);
nor U870 (N_870,N_269,In_792);
and U871 (N_871,In_110,In_170);
nand U872 (N_872,N_399,In_253);
xor U873 (N_873,In_55,In_1293);
nor U874 (N_874,N_35,N_74);
nand U875 (N_875,In_42,N_383);
or U876 (N_876,In_276,N_404);
and U877 (N_877,N_384,N_356);
nand U878 (N_878,In_460,In_863);
or U879 (N_879,N_488,N_273);
nand U880 (N_880,In_1198,N_162);
and U881 (N_881,In_846,In_202);
nand U882 (N_882,In_1169,In_267);
and U883 (N_883,N_489,In_852);
nand U884 (N_884,N_94,In_398);
nor U885 (N_885,N_188,N_434);
nand U886 (N_886,N_339,N_17);
and U887 (N_887,In_1291,In_64);
xnor U888 (N_888,In_1471,In_1314);
and U889 (N_889,In_171,N_325);
nor U890 (N_890,N_299,In_105);
or U891 (N_891,N_186,In_90);
or U892 (N_892,N_257,N_353);
and U893 (N_893,In_1276,N_290);
xnor U894 (N_894,In_452,N_426);
or U895 (N_895,In_705,In_83);
and U896 (N_896,N_95,N_201);
xnor U897 (N_897,In_875,N_213);
nor U898 (N_898,In_126,In_1258);
nand U899 (N_899,N_413,In_227);
or U900 (N_900,In_1077,In_1273);
nand U901 (N_901,N_286,In_249);
nand U902 (N_902,In_470,N_348);
and U903 (N_903,In_490,In_941);
nor U904 (N_904,In_291,N_16);
xor U905 (N_905,In_1196,In_718);
or U906 (N_906,N_232,N_349);
xor U907 (N_907,In_77,In_1055);
and U908 (N_908,In_8,In_376);
xnor U909 (N_909,In_602,N_303);
xnor U910 (N_910,N_304,N_377);
nor U911 (N_911,N_193,N_248);
and U912 (N_912,N_314,In_773);
or U913 (N_913,In_1134,In_273);
xor U914 (N_914,N_158,In_323);
xor U915 (N_915,In_1278,N_97);
and U916 (N_916,In_137,In_51);
xnor U917 (N_917,In_1317,N_202);
and U918 (N_918,N_15,In_1335);
nor U919 (N_919,In_443,N_408);
xor U920 (N_920,In_331,N_8);
or U921 (N_921,N_54,In_921);
and U922 (N_922,N_311,N_341);
nor U923 (N_923,N_275,In_1202);
nor U924 (N_924,N_228,In_1383);
and U925 (N_925,N_104,N_472);
nand U926 (N_926,N_231,N_223);
xnor U927 (N_927,In_287,In_281);
nor U928 (N_928,In_816,In_1394);
xnor U929 (N_929,In_896,N_368);
or U930 (N_930,N_252,In_362);
nor U931 (N_931,N_111,In_1148);
and U932 (N_932,N_313,N_63);
xnor U933 (N_933,N_475,N_131);
nor U934 (N_934,N_86,N_88);
nor U935 (N_935,N_206,N_442);
and U936 (N_936,N_378,N_430);
or U937 (N_937,N_165,In_948);
or U938 (N_938,N_444,N_440);
nor U939 (N_939,N_3,In_1441);
nand U940 (N_940,In_957,In_1450);
nand U941 (N_941,In_1344,In_830);
and U942 (N_942,In_965,N_263);
nand U943 (N_943,In_717,N_272);
xnor U944 (N_944,In_1126,N_209);
xor U945 (N_945,N_298,N_129);
nand U946 (N_946,N_317,N_59);
and U947 (N_947,N_396,N_178);
or U948 (N_948,In_590,N_458);
nor U949 (N_949,In_1082,N_283);
xor U950 (N_950,In_155,In_66);
xor U951 (N_951,In_1226,In_1114);
nor U952 (N_952,N_160,N_200);
and U953 (N_953,In_98,In_958);
or U954 (N_954,In_1404,N_335);
or U955 (N_955,In_1208,In_660);
xnor U956 (N_956,In_1163,In_1094);
and U957 (N_957,In_1086,N_402);
nor U958 (N_958,N_10,In_414);
or U959 (N_959,In_632,N_246);
xnor U960 (N_960,N_474,In_572);
and U961 (N_961,In_382,In_150);
and U962 (N_962,N_96,N_432);
nor U963 (N_963,N_450,N_40);
or U964 (N_964,In_1051,N_318);
or U965 (N_965,In_996,In_492);
nor U966 (N_966,In_1448,In_1124);
and U967 (N_967,In_84,N_285);
nand U968 (N_968,In_308,In_1478);
nor U969 (N_969,In_1039,In_47);
and U970 (N_970,In_1418,N_255);
xnor U971 (N_971,In_1233,In_1303);
nand U972 (N_972,N_9,In_685);
xnor U973 (N_973,N_321,In_220);
xor U974 (N_974,In_453,N_324);
xor U975 (N_975,N_390,In_1252);
and U976 (N_976,N_308,In_835);
nand U977 (N_977,In_1395,N_51);
or U978 (N_978,N_365,N_130);
nand U979 (N_979,N_461,N_312);
and U980 (N_980,In_766,N_462);
nand U981 (N_981,In_379,In_1408);
and U982 (N_982,In_1054,In_565);
and U983 (N_983,N_446,N_296);
nand U984 (N_984,In_57,N_491);
and U985 (N_985,N_121,N_471);
and U986 (N_986,N_195,In_804);
nand U987 (N_987,In_1369,In_125);
or U988 (N_988,In_967,N_479);
xnor U989 (N_989,N_411,In_689);
nand U990 (N_990,N_473,N_169);
xnor U991 (N_991,N_278,N_80);
and U992 (N_992,In_237,In_348);
nand U993 (N_993,In_591,N_114);
nand U994 (N_994,In_1080,N_422);
nand U995 (N_995,N_364,In_1201);
xnor U996 (N_996,N_264,N_316);
nor U997 (N_997,In_881,N_412);
nand U998 (N_998,In_154,N_421);
or U999 (N_999,In_505,In_768);
and U1000 (N_1000,N_964,N_940);
and U1001 (N_1001,N_519,N_677);
and U1002 (N_1002,N_745,N_701);
xor U1003 (N_1003,N_749,N_845);
nor U1004 (N_1004,N_605,N_739);
and U1005 (N_1005,N_961,N_883);
xor U1006 (N_1006,N_674,N_714);
xor U1007 (N_1007,N_537,N_588);
nor U1008 (N_1008,N_603,N_680);
xor U1009 (N_1009,N_540,N_771);
nor U1010 (N_1010,N_769,N_791);
nor U1011 (N_1011,N_687,N_644);
nor U1012 (N_1012,N_766,N_936);
nor U1013 (N_1013,N_904,N_738);
nor U1014 (N_1014,N_578,N_673);
xor U1015 (N_1015,N_855,N_682);
or U1016 (N_1016,N_841,N_531);
or U1017 (N_1017,N_805,N_610);
and U1018 (N_1018,N_720,N_843);
and U1019 (N_1019,N_669,N_663);
nor U1020 (N_1020,N_801,N_923);
or U1021 (N_1021,N_910,N_998);
or U1022 (N_1022,N_909,N_915);
or U1023 (N_1023,N_545,N_778);
xor U1024 (N_1024,N_988,N_846);
nor U1025 (N_1025,N_830,N_812);
nand U1026 (N_1026,N_725,N_630);
nor U1027 (N_1027,N_970,N_615);
nand U1028 (N_1028,N_978,N_922);
nand U1029 (N_1029,N_737,N_650);
xor U1030 (N_1030,N_799,N_562);
nor U1031 (N_1031,N_876,N_821);
nand U1032 (N_1032,N_500,N_960);
or U1033 (N_1033,N_990,N_684);
nor U1034 (N_1034,N_678,N_827);
nor U1035 (N_1035,N_554,N_625);
or U1036 (N_1036,N_937,N_885);
nor U1037 (N_1037,N_604,N_686);
xnor U1038 (N_1038,N_757,N_718);
and U1039 (N_1039,N_814,N_586);
or U1040 (N_1040,N_849,N_616);
or U1041 (N_1041,N_808,N_925);
or U1042 (N_1042,N_583,N_698);
xor U1043 (N_1043,N_787,N_994);
xnor U1044 (N_1044,N_592,N_968);
nor U1045 (N_1045,N_565,N_889);
nand U1046 (N_1046,N_785,N_842);
nand U1047 (N_1047,N_706,N_959);
or U1048 (N_1048,N_878,N_590);
and U1049 (N_1049,N_896,N_617);
nor U1050 (N_1050,N_820,N_727);
nor U1051 (N_1051,N_675,N_532);
xor U1052 (N_1052,N_666,N_600);
or U1053 (N_1053,N_819,N_831);
and U1054 (N_1054,N_579,N_764);
nor U1055 (N_1055,N_618,N_670);
nand U1056 (N_1056,N_941,N_755);
xor U1057 (N_1057,N_552,N_786);
and U1058 (N_1058,N_753,N_895);
nor U1059 (N_1059,N_869,N_679);
and U1060 (N_1060,N_694,N_699);
nand U1061 (N_1061,N_914,N_571);
or U1062 (N_1062,N_564,N_829);
nand U1063 (N_1063,N_730,N_813);
nor U1064 (N_1064,N_956,N_744);
and U1065 (N_1065,N_711,N_983);
or U1066 (N_1066,N_920,N_932);
or U1067 (N_1067,N_837,N_870);
nand U1068 (N_1068,N_511,N_832);
nand U1069 (N_1069,N_852,N_634);
xnor U1070 (N_1070,N_639,N_707);
or U1071 (N_1071,N_979,N_539);
xnor U1072 (N_1072,N_916,N_763);
xor U1073 (N_1073,N_515,N_760);
and U1074 (N_1074,N_807,N_879);
nand U1075 (N_1075,N_798,N_765);
xor U1076 (N_1076,N_563,N_697);
nand U1077 (N_1077,N_912,N_958);
xor U1078 (N_1078,N_560,N_856);
nand U1079 (N_1079,N_882,N_622);
nand U1080 (N_1080,N_952,N_629);
nand U1081 (N_1081,N_938,N_542);
or U1082 (N_1082,N_790,N_795);
nor U1083 (N_1083,N_865,N_651);
nand U1084 (N_1084,N_661,N_570);
nand U1085 (N_1085,N_803,N_822);
and U1086 (N_1086,N_736,N_894);
nor U1087 (N_1087,N_951,N_507);
nor U1088 (N_1088,N_752,N_872);
nand U1089 (N_1089,N_891,N_750);
xnor U1090 (N_1090,N_587,N_781);
or U1091 (N_1091,N_756,N_504);
nor U1092 (N_1092,N_955,N_643);
and U1093 (N_1093,N_524,N_741);
nor U1094 (N_1094,N_591,N_944);
and U1095 (N_1095,N_991,N_800);
nand U1096 (N_1096,N_620,N_754);
nand U1097 (N_1097,N_657,N_969);
nor U1098 (N_1098,N_596,N_859);
xor U1099 (N_1099,N_788,N_649);
or U1100 (N_1100,N_804,N_732);
nand U1101 (N_1101,N_659,N_641);
xnor U1102 (N_1102,N_835,N_907);
nor U1103 (N_1103,N_709,N_917);
nand U1104 (N_1104,N_762,N_726);
nand U1105 (N_1105,N_713,N_546);
xnor U1106 (N_1106,N_577,N_783);
and U1107 (N_1107,N_867,N_864);
nand U1108 (N_1108,N_866,N_628);
xnor U1109 (N_1109,N_536,N_935);
nor U1110 (N_1110,N_556,N_836);
nor U1111 (N_1111,N_580,N_768);
or U1112 (N_1112,N_899,N_522);
nor U1113 (N_1113,N_635,N_975);
nor U1114 (N_1114,N_557,N_857);
xor U1115 (N_1115,N_594,N_890);
nand U1116 (N_1116,N_535,N_868);
nor U1117 (N_1117,N_576,N_776);
nand U1118 (N_1118,N_811,N_505);
or U1119 (N_1119,N_559,N_929);
or U1120 (N_1120,N_602,N_671);
nor U1121 (N_1121,N_810,N_609);
and U1122 (N_1122,N_976,N_569);
nor U1123 (N_1123,N_547,N_921);
or U1124 (N_1124,N_695,N_534);
xnor U1125 (N_1125,N_926,N_824);
or U1126 (N_1126,N_729,N_517);
nand U1127 (N_1127,N_893,N_653);
or U1128 (N_1128,N_815,N_510);
xnor U1129 (N_1129,N_688,N_624);
or U1130 (N_1130,N_567,N_612);
or U1131 (N_1131,N_574,N_908);
or U1132 (N_1132,N_740,N_934);
nand U1133 (N_1133,N_913,N_638);
or U1134 (N_1134,N_973,N_794);
nand U1135 (N_1135,N_550,N_516);
nor U1136 (N_1136,N_862,N_502);
xnor U1137 (N_1137,N_685,N_903);
or U1138 (N_1138,N_668,N_823);
xnor U1139 (N_1139,N_627,N_746);
and U1140 (N_1140,N_691,N_851);
and U1141 (N_1141,N_967,N_667);
and U1142 (N_1142,N_514,N_621);
nand U1143 (N_1143,N_942,N_853);
nand U1144 (N_1144,N_700,N_992);
and U1145 (N_1145,N_731,N_607);
nor U1146 (N_1146,N_946,N_954);
nor U1147 (N_1147,N_723,N_900);
xnor U1148 (N_1148,N_809,N_985);
nor U1149 (N_1149,N_689,N_833);
nor U1150 (N_1150,N_555,N_608);
nand U1151 (N_1151,N_654,N_767);
xnor U1152 (N_1152,N_963,N_640);
xnor U1153 (N_1153,N_708,N_984);
nand U1154 (N_1154,N_989,N_528);
xnor U1155 (N_1155,N_533,N_693);
and U1156 (N_1156,N_541,N_652);
and U1157 (N_1157,N_598,N_646);
xnor U1158 (N_1158,N_902,N_672);
and U1159 (N_1159,N_887,N_793);
xnor U1160 (N_1160,N_690,N_508);
xnor U1161 (N_1161,N_747,N_911);
nand U1162 (N_1162,N_513,N_931);
xnor U1163 (N_1163,N_774,N_888);
and U1164 (N_1164,N_645,N_838);
nand U1165 (N_1165,N_719,N_637);
nand U1166 (N_1166,N_544,N_712);
or U1167 (N_1167,N_972,N_656);
or U1168 (N_1168,N_676,N_543);
nor U1169 (N_1169,N_681,N_683);
or U1170 (N_1170,N_779,N_806);
nand U1171 (N_1171,N_977,N_982);
nor U1172 (N_1172,N_553,N_884);
nor U1173 (N_1173,N_660,N_770);
xnor U1174 (N_1174,N_568,N_595);
nor U1175 (N_1175,N_817,N_789);
and U1176 (N_1176,N_850,N_636);
nor U1177 (N_1177,N_772,N_796);
nor U1178 (N_1178,N_816,N_530);
nand U1179 (N_1179,N_953,N_924);
and U1180 (N_1180,N_728,N_705);
and U1181 (N_1181,N_761,N_825);
xor U1182 (N_1182,N_782,N_575);
xor U1183 (N_1183,N_715,N_525);
and U1184 (N_1184,N_647,N_966);
and U1185 (N_1185,N_585,N_573);
and U1186 (N_1186,N_818,N_993);
nand U1187 (N_1187,N_927,N_945);
and U1188 (N_1188,N_633,N_987);
xor U1189 (N_1189,N_703,N_548);
xnor U1190 (N_1190,N_529,N_898);
nand U1191 (N_1191,N_844,N_780);
nand U1192 (N_1192,N_881,N_584);
nand U1193 (N_1193,N_581,N_858);
nor U1194 (N_1194,N_626,N_521);
nand U1195 (N_1195,N_611,N_854);
nor U1196 (N_1196,N_918,N_623);
or U1197 (N_1197,N_861,N_971);
and U1198 (N_1198,N_995,N_506);
xnor U1199 (N_1199,N_561,N_965);
nor U1200 (N_1200,N_566,N_751);
and U1201 (N_1201,N_549,N_518);
nand U1202 (N_1202,N_802,N_501);
or U1203 (N_1203,N_551,N_828);
or U1204 (N_1204,N_759,N_704);
nor U1205 (N_1205,N_905,N_880);
or U1206 (N_1206,N_860,N_826);
nand U1207 (N_1207,N_997,N_877);
nand U1208 (N_1208,N_797,N_980);
nand U1209 (N_1209,N_558,N_839);
or U1210 (N_1210,N_962,N_724);
and U1211 (N_1211,N_722,N_901);
xnor U1212 (N_1212,N_742,N_748);
and U1213 (N_1213,N_642,N_892);
or U1214 (N_1214,N_665,N_509);
xor U1215 (N_1215,N_601,N_658);
or U1216 (N_1216,N_758,N_734);
and U1217 (N_1217,N_784,N_919);
nor U1218 (N_1218,N_949,N_597);
xor U1219 (N_1219,N_947,N_743);
and U1220 (N_1220,N_981,N_943);
and U1221 (N_1221,N_939,N_655);
nand U1222 (N_1222,N_527,N_735);
and U1223 (N_1223,N_582,N_572);
and U1224 (N_1224,N_614,N_950);
nand U1225 (N_1225,N_523,N_777);
and U1226 (N_1226,N_717,N_792);
nor U1227 (N_1227,N_773,N_906);
nor U1228 (N_1228,N_840,N_886);
nand U1229 (N_1229,N_847,N_775);
or U1230 (N_1230,N_897,N_863);
xnor U1231 (N_1231,N_996,N_948);
xor U1232 (N_1232,N_873,N_871);
and U1233 (N_1233,N_619,N_538);
and U1234 (N_1234,N_974,N_928);
and U1235 (N_1235,N_986,N_710);
or U1236 (N_1236,N_930,N_933);
nor U1237 (N_1237,N_696,N_648);
or U1238 (N_1238,N_520,N_702);
xor U1239 (N_1239,N_613,N_662);
nand U1240 (N_1240,N_692,N_957);
nor U1241 (N_1241,N_716,N_593);
nor U1242 (N_1242,N_848,N_875);
xor U1243 (N_1243,N_664,N_526);
and U1244 (N_1244,N_874,N_512);
and U1245 (N_1245,N_606,N_733);
nor U1246 (N_1246,N_631,N_999);
nor U1247 (N_1247,N_503,N_599);
xnor U1248 (N_1248,N_834,N_632);
nand U1249 (N_1249,N_721,N_589);
xnor U1250 (N_1250,N_674,N_918);
and U1251 (N_1251,N_549,N_502);
and U1252 (N_1252,N_942,N_876);
xnor U1253 (N_1253,N_556,N_769);
or U1254 (N_1254,N_891,N_882);
nor U1255 (N_1255,N_965,N_660);
nand U1256 (N_1256,N_565,N_877);
nand U1257 (N_1257,N_942,N_950);
and U1258 (N_1258,N_921,N_561);
xor U1259 (N_1259,N_509,N_820);
or U1260 (N_1260,N_634,N_751);
xor U1261 (N_1261,N_929,N_860);
or U1262 (N_1262,N_630,N_599);
xor U1263 (N_1263,N_647,N_954);
xor U1264 (N_1264,N_634,N_980);
nand U1265 (N_1265,N_792,N_547);
and U1266 (N_1266,N_674,N_634);
nor U1267 (N_1267,N_586,N_578);
nand U1268 (N_1268,N_801,N_740);
and U1269 (N_1269,N_936,N_601);
xnor U1270 (N_1270,N_564,N_738);
xor U1271 (N_1271,N_582,N_945);
nor U1272 (N_1272,N_503,N_506);
and U1273 (N_1273,N_781,N_756);
nand U1274 (N_1274,N_785,N_754);
nand U1275 (N_1275,N_546,N_645);
and U1276 (N_1276,N_936,N_596);
nor U1277 (N_1277,N_804,N_738);
or U1278 (N_1278,N_993,N_847);
nand U1279 (N_1279,N_965,N_565);
xor U1280 (N_1280,N_969,N_933);
and U1281 (N_1281,N_572,N_958);
nor U1282 (N_1282,N_604,N_898);
xor U1283 (N_1283,N_781,N_795);
nand U1284 (N_1284,N_919,N_584);
nand U1285 (N_1285,N_929,N_849);
nand U1286 (N_1286,N_966,N_937);
xor U1287 (N_1287,N_972,N_571);
and U1288 (N_1288,N_636,N_676);
nand U1289 (N_1289,N_707,N_977);
or U1290 (N_1290,N_810,N_612);
and U1291 (N_1291,N_597,N_812);
nor U1292 (N_1292,N_549,N_680);
xnor U1293 (N_1293,N_918,N_984);
and U1294 (N_1294,N_643,N_655);
xor U1295 (N_1295,N_756,N_846);
nand U1296 (N_1296,N_776,N_867);
nand U1297 (N_1297,N_911,N_996);
nor U1298 (N_1298,N_929,N_935);
nand U1299 (N_1299,N_545,N_844);
nor U1300 (N_1300,N_815,N_946);
or U1301 (N_1301,N_662,N_748);
nand U1302 (N_1302,N_826,N_898);
or U1303 (N_1303,N_914,N_747);
nand U1304 (N_1304,N_616,N_823);
nand U1305 (N_1305,N_843,N_834);
or U1306 (N_1306,N_606,N_805);
xnor U1307 (N_1307,N_902,N_912);
xnor U1308 (N_1308,N_658,N_644);
nand U1309 (N_1309,N_991,N_838);
or U1310 (N_1310,N_579,N_769);
nor U1311 (N_1311,N_736,N_795);
xor U1312 (N_1312,N_934,N_901);
nor U1313 (N_1313,N_642,N_959);
or U1314 (N_1314,N_619,N_659);
nand U1315 (N_1315,N_917,N_901);
or U1316 (N_1316,N_823,N_719);
nor U1317 (N_1317,N_676,N_795);
nand U1318 (N_1318,N_792,N_646);
xnor U1319 (N_1319,N_682,N_671);
or U1320 (N_1320,N_743,N_815);
and U1321 (N_1321,N_893,N_701);
or U1322 (N_1322,N_512,N_986);
nand U1323 (N_1323,N_972,N_557);
nand U1324 (N_1324,N_881,N_850);
xnor U1325 (N_1325,N_912,N_740);
or U1326 (N_1326,N_824,N_540);
and U1327 (N_1327,N_945,N_840);
and U1328 (N_1328,N_735,N_760);
and U1329 (N_1329,N_556,N_653);
nand U1330 (N_1330,N_649,N_687);
or U1331 (N_1331,N_895,N_669);
xor U1332 (N_1332,N_717,N_551);
nand U1333 (N_1333,N_634,N_665);
nand U1334 (N_1334,N_984,N_568);
and U1335 (N_1335,N_765,N_683);
xor U1336 (N_1336,N_678,N_950);
nor U1337 (N_1337,N_910,N_672);
xnor U1338 (N_1338,N_635,N_519);
xnor U1339 (N_1339,N_783,N_509);
nand U1340 (N_1340,N_543,N_773);
nor U1341 (N_1341,N_648,N_908);
nor U1342 (N_1342,N_523,N_657);
nand U1343 (N_1343,N_802,N_509);
or U1344 (N_1344,N_867,N_691);
xor U1345 (N_1345,N_787,N_766);
xor U1346 (N_1346,N_628,N_980);
nor U1347 (N_1347,N_824,N_896);
xor U1348 (N_1348,N_730,N_809);
nand U1349 (N_1349,N_961,N_556);
xor U1350 (N_1350,N_680,N_779);
nand U1351 (N_1351,N_777,N_947);
nor U1352 (N_1352,N_893,N_736);
nor U1353 (N_1353,N_856,N_921);
or U1354 (N_1354,N_604,N_817);
and U1355 (N_1355,N_585,N_879);
or U1356 (N_1356,N_598,N_987);
and U1357 (N_1357,N_920,N_537);
and U1358 (N_1358,N_949,N_655);
xnor U1359 (N_1359,N_737,N_900);
nor U1360 (N_1360,N_684,N_625);
and U1361 (N_1361,N_719,N_949);
nor U1362 (N_1362,N_524,N_726);
nand U1363 (N_1363,N_814,N_726);
nor U1364 (N_1364,N_709,N_927);
and U1365 (N_1365,N_881,N_713);
nor U1366 (N_1366,N_817,N_913);
nand U1367 (N_1367,N_806,N_603);
and U1368 (N_1368,N_588,N_917);
nor U1369 (N_1369,N_640,N_574);
or U1370 (N_1370,N_804,N_583);
xor U1371 (N_1371,N_896,N_744);
nor U1372 (N_1372,N_870,N_778);
nand U1373 (N_1373,N_502,N_847);
nand U1374 (N_1374,N_523,N_939);
nor U1375 (N_1375,N_841,N_687);
nand U1376 (N_1376,N_667,N_952);
xor U1377 (N_1377,N_785,N_645);
nand U1378 (N_1378,N_823,N_990);
xnor U1379 (N_1379,N_826,N_851);
and U1380 (N_1380,N_893,N_972);
or U1381 (N_1381,N_963,N_518);
xnor U1382 (N_1382,N_656,N_673);
nand U1383 (N_1383,N_545,N_935);
nand U1384 (N_1384,N_943,N_921);
nor U1385 (N_1385,N_915,N_686);
nor U1386 (N_1386,N_732,N_893);
and U1387 (N_1387,N_656,N_805);
xor U1388 (N_1388,N_937,N_847);
xor U1389 (N_1389,N_628,N_721);
and U1390 (N_1390,N_914,N_617);
nor U1391 (N_1391,N_998,N_751);
nand U1392 (N_1392,N_994,N_946);
nand U1393 (N_1393,N_623,N_719);
nor U1394 (N_1394,N_535,N_889);
nor U1395 (N_1395,N_943,N_983);
nor U1396 (N_1396,N_542,N_820);
and U1397 (N_1397,N_599,N_973);
and U1398 (N_1398,N_770,N_682);
and U1399 (N_1399,N_672,N_836);
or U1400 (N_1400,N_628,N_630);
and U1401 (N_1401,N_857,N_865);
nand U1402 (N_1402,N_860,N_808);
or U1403 (N_1403,N_988,N_568);
xor U1404 (N_1404,N_701,N_878);
or U1405 (N_1405,N_657,N_749);
nand U1406 (N_1406,N_859,N_680);
nand U1407 (N_1407,N_826,N_843);
or U1408 (N_1408,N_927,N_649);
nand U1409 (N_1409,N_835,N_826);
xor U1410 (N_1410,N_838,N_779);
xor U1411 (N_1411,N_742,N_880);
xnor U1412 (N_1412,N_921,N_576);
and U1413 (N_1413,N_530,N_605);
or U1414 (N_1414,N_911,N_537);
nor U1415 (N_1415,N_896,N_622);
or U1416 (N_1416,N_789,N_747);
nand U1417 (N_1417,N_842,N_800);
xnor U1418 (N_1418,N_734,N_627);
nand U1419 (N_1419,N_831,N_740);
or U1420 (N_1420,N_682,N_962);
nand U1421 (N_1421,N_729,N_855);
xor U1422 (N_1422,N_970,N_868);
or U1423 (N_1423,N_535,N_503);
xnor U1424 (N_1424,N_590,N_583);
or U1425 (N_1425,N_777,N_864);
xnor U1426 (N_1426,N_692,N_681);
nand U1427 (N_1427,N_590,N_552);
nand U1428 (N_1428,N_936,N_657);
xnor U1429 (N_1429,N_631,N_704);
nand U1430 (N_1430,N_899,N_889);
xor U1431 (N_1431,N_877,N_527);
nand U1432 (N_1432,N_711,N_629);
xor U1433 (N_1433,N_594,N_566);
xnor U1434 (N_1434,N_745,N_643);
xnor U1435 (N_1435,N_920,N_686);
nor U1436 (N_1436,N_701,N_822);
nor U1437 (N_1437,N_857,N_649);
nand U1438 (N_1438,N_969,N_879);
nand U1439 (N_1439,N_938,N_720);
xnor U1440 (N_1440,N_509,N_659);
xnor U1441 (N_1441,N_612,N_680);
and U1442 (N_1442,N_897,N_762);
xor U1443 (N_1443,N_612,N_723);
nand U1444 (N_1444,N_716,N_543);
nand U1445 (N_1445,N_947,N_530);
and U1446 (N_1446,N_986,N_550);
nor U1447 (N_1447,N_671,N_700);
or U1448 (N_1448,N_821,N_670);
xor U1449 (N_1449,N_770,N_898);
nand U1450 (N_1450,N_678,N_543);
xnor U1451 (N_1451,N_747,N_860);
xor U1452 (N_1452,N_766,N_780);
and U1453 (N_1453,N_521,N_680);
or U1454 (N_1454,N_912,N_824);
nor U1455 (N_1455,N_590,N_839);
and U1456 (N_1456,N_998,N_732);
nor U1457 (N_1457,N_801,N_547);
and U1458 (N_1458,N_980,N_974);
xnor U1459 (N_1459,N_580,N_941);
xnor U1460 (N_1460,N_750,N_775);
or U1461 (N_1461,N_787,N_594);
or U1462 (N_1462,N_693,N_587);
and U1463 (N_1463,N_936,N_611);
and U1464 (N_1464,N_670,N_686);
xnor U1465 (N_1465,N_899,N_545);
nand U1466 (N_1466,N_732,N_580);
and U1467 (N_1467,N_837,N_825);
or U1468 (N_1468,N_815,N_521);
and U1469 (N_1469,N_702,N_714);
xnor U1470 (N_1470,N_986,N_508);
nor U1471 (N_1471,N_556,N_944);
xnor U1472 (N_1472,N_719,N_678);
or U1473 (N_1473,N_647,N_834);
nand U1474 (N_1474,N_678,N_769);
or U1475 (N_1475,N_513,N_905);
or U1476 (N_1476,N_504,N_772);
nor U1477 (N_1477,N_579,N_846);
or U1478 (N_1478,N_976,N_911);
and U1479 (N_1479,N_733,N_832);
nand U1480 (N_1480,N_860,N_717);
or U1481 (N_1481,N_898,N_739);
nor U1482 (N_1482,N_861,N_969);
nor U1483 (N_1483,N_945,N_532);
xnor U1484 (N_1484,N_906,N_559);
xnor U1485 (N_1485,N_947,N_857);
nor U1486 (N_1486,N_537,N_513);
or U1487 (N_1487,N_972,N_549);
or U1488 (N_1488,N_724,N_570);
nor U1489 (N_1489,N_614,N_676);
or U1490 (N_1490,N_524,N_625);
or U1491 (N_1491,N_756,N_592);
xnor U1492 (N_1492,N_528,N_818);
xor U1493 (N_1493,N_912,N_872);
nand U1494 (N_1494,N_547,N_628);
xnor U1495 (N_1495,N_711,N_936);
or U1496 (N_1496,N_680,N_652);
or U1497 (N_1497,N_654,N_622);
nor U1498 (N_1498,N_984,N_695);
nand U1499 (N_1499,N_949,N_848);
nand U1500 (N_1500,N_1040,N_1127);
and U1501 (N_1501,N_1070,N_1091);
and U1502 (N_1502,N_1097,N_1045);
or U1503 (N_1503,N_1454,N_1167);
nor U1504 (N_1504,N_1001,N_1014);
nand U1505 (N_1505,N_1220,N_1345);
nand U1506 (N_1506,N_1122,N_1241);
or U1507 (N_1507,N_1485,N_1055);
or U1508 (N_1508,N_1201,N_1495);
or U1509 (N_1509,N_1210,N_1391);
xor U1510 (N_1510,N_1400,N_1065);
or U1511 (N_1511,N_1363,N_1271);
and U1512 (N_1512,N_1099,N_1115);
or U1513 (N_1513,N_1132,N_1446);
xnor U1514 (N_1514,N_1203,N_1289);
and U1515 (N_1515,N_1135,N_1267);
nand U1516 (N_1516,N_1433,N_1116);
or U1517 (N_1517,N_1272,N_1060);
or U1518 (N_1518,N_1120,N_1405);
xnor U1519 (N_1519,N_1382,N_1402);
or U1520 (N_1520,N_1484,N_1294);
and U1521 (N_1521,N_1067,N_1321);
and U1522 (N_1522,N_1440,N_1474);
nor U1523 (N_1523,N_1119,N_1475);
nor U1524 (N_1524,N_1429,N_1244);
or U1525 (N_1525,N_1202,N_1121);
and U1526 (N_1526,N_1236,N_1385);
or U1527 (N_1527,N_1156,N_1287);
nor U1528 (N_1528,N_1048,N_1364);
xor U1529 (N_1529,N_1112,N_1101);
nand U1530 (N_1530,N_1259,N_1204);
xnor U1531 (N_1531,N_1367,N_1009);
xnor U1532 (N_1532,N_1397,N_1104);
and U1533 (N_1533,N_1021,N_1479);
nand U1534 (N_1534,N_1148,N_1169);
nand U1535 (N_1535,N_1336,N_1111);
xor U1536 (N_1536,N_1403,N_1327);
and U1537 (N_1537,N_1212,N_1129);
and U1538 (N_1538,N_1178,N_1254);
and U1539 (N_1539,N_1421,N_1420);
or U1540 (N_1540,N_1467,N_1238);
nor U1541 (N_1541,N_1373,N_1029);
or U1542 (N_1542,N_1312,N_1039);
nand U1543 (N_1543,N_1488,N_1252);
nor U1544 (N_1544,N_1198,N_1188);
and U1545 (N_1545,N_1340,N_1269);
nor U1546 (N_1546,N_1263,N_1425);
xnor U1547 (N_1547,N_1406,N_1218);
xnor U1548 (N_1548,N_1090,N_1284);
xnor U1549 (N_1549,N_1036,N_1481);
nor U1550 (N_1550,N_1080,N_1240);
xnor U1551 (N_1551,N_1118,N_1016);
nor U1552 (N_1552,N_1337,N_1493);
or U1553 (N_1553,N_1462,N_1466);
nand U1554 (N_1554,N_1207,N_1358);
nand U1555 (N_1555,N_1298,N_1186);
and U1556 (N_1556,N_1492,N_1460);
and U1557 (N_1557,N_1000,N_1133);
or U1558 (N_1558,N_1046,N_1450);
xor U1559 (N_1559,N_1352,N_1319);
nand U1560 (N_1560,N_1057,N_1458);
or U1561 (N_1561,N_1239,N_1486);
nor U1562 (N_1562,N_1066,N_1139);
and U1563 (N_1563,N_1439,N_1030);
or U1564 (N_1564,N_1184,N_1268);
or U1565 (N_1565,N_1314,N_1468);
or U1566 (N_1566,N_1437,N_1062);
and U1567 (N_1567,N_1185,N_1187);
or U1568 (N_1568,N_1226,N_1018);
xor U1569 (N_1569,N_1214,N_1227);
and U1570 (N_1570,N_1213,N_1138);
or U1571 (N_1571,N_1292,N_1211);
nor U1572 (N_1572,N_1103,N_1266);
or U1573 (N_1573,N_1426,N_1071);
or U1574 (N_1574,N_1375,N_1087);
nand U1575 (N_1575,N_1413,N_1061);
and U1576 (N_1576,N_1170,N_1346);
and U1577 (N_1577,N_1320,N_1410);
and U1578 (N_1578,N_1355,N_1461);
nand U1579 (N_1579,N_1409,N_1301);
or U1580 (N_1580,N_1037,N_1109);
nand U1581 (N_1581,N_1150,N_1360);
nor U1582 (N_1582,N_1283,N_1278);
nor U1583 (N_1583,N_1147,N_1372);
xnor U1584 (N_1584,N_1344,N_1117);
nor U1585 (N_1585,N_1072,N_1331);
nand U1586 (N_1586,N_1487,N_1280);
or U1587 (N_1587,N_1357,N_1005);
nor U1588 (N_1588,N_1158,N_1359);
nand U1589 (N_1589,N_1370,N_1463);
nand U1590 (N_1590,N_1384,N_1295);
nor U1591 (N_1591,N_1428,N_1064);
nor U1592 (N_1592,N_1224,N_1482);
and U1593 (N_1593,N_1052,N_1457);
xor U1594 (N_1594,N_1235,N_1386);
nand U1595 (N_1595,N_1137,N_1053);
and U1596 (N_1596,N_1221,N_1449);
nand U1597 (N_1597,N_1034,N_1361);
nor U1598 (N_1598,N_1206,N_1377);
nor U1599 (N_1599,N_1153,N_1033);
nor U1600 (N_1600,N_1200,N_1223);
nand U1601 (N_1601,N_1076,N_1019);
nor U1602 (N_1602,N_1190,N_1498);
nor U1603 (N_1603,N_1081,N_1423);
and U1604 (N_1604,N_1325,N_1477);
and U1605 (N_1605,N_1293,N_1307);
and U1606 (N_1606,N_1043,N_1245);
nand U1607 (N_1607,N_1165,N_1339);
nand U1608 (N_1608,N_1494,N_1166);
nor U1609 (N_1609,N_1078,N_1414);
and U1610 (N_1610,N_1007,N_1179);
nand U1611 (N_1611,N_1401,N_1251);
xnor U1612 (N_1612,N_1242,N_1197);
or U1613 (N_1613,N_1024,N_1335);
nand U1614 (N_1614,N_1092,N_1075);
nor U1615 (N_1615,N_1130,N_1246);
xnor U1616 (N_1616,N_1387,N_1038);
and U1617 (N_1617,N_1323,N_1309);
and U1618 (N_1618,N_1162,N_1277);
nand U1619 (N_1619,N_1082,N_1248);
or U1620 (N_1620,N_1054,N_1107);
nor U1621 (N_1621,N_1253,N_1383);
or U1622 (N_1622,N_1453,N_1088);
xnor U1623 (N_1623,N_1143,N_1444);
xor U1624 (N_1624,N_1390,N_1217);
nand U1625 (N_1625,N_1230,N_1448);
nor U1626 (N_1626,N_1191,N_1041);
nand U1627 (N_1627,N_1181,N_1025);
nand U1628 (N_1628,N_1459,N_1394);
nor U1629 (N_1629,N_1094,N_1183);
xor U1630 (N_1630,N_1483,N_1436);
and U1631 (N_1631,N_1144,N_1152);
nand U1632 (N_1632,N_1308,N_1013);
or U1633 (N_1633,N_1445,N_1002);
or U1634 (N_1634,N_1069,N_1250);
or U1635 (N_1635,N_1378,N_1003);
or U1636 (N_1636,N_1304,N_1419);
nand U1637 (N_1637,N_1379,N_1356);
xor U1638 (N_1638,N_1134,N_1282);
nand U1639 (N_1639,N_1126,N_1279);
or U1640 (N_1640,N_1442,N_1142);
xor U1641 (N_1641,N_1189,N_1365);
or U1642 (N_1642,N_1464,N_1196);
or U1643 (N_1643,N_1297,N_1234);
and U1644 (N_1644,N_1318,N_1044);
nor U1645 (N_1645,N_1108,N_1317);
nand U1646 (N_1646,N_1424,N_1476);
or U1647 (N_1647,N_1231,N_1085);
xor U1648 (N_1648,N_1077,N_1443);
xor U1649 (N_1649,N_1208,N_1399);
or U1650 (N_1650,N_1299,N_1222);
nor U1651 (N_1651,N_1465,N_1163);
xor U1652 (N_1652,N_1258,N_1418);
and U1653 (N_1653,N_1051,N_1435);
nand U1654 (N_1654,N_1031,N_1412);
xnor U1655 (N_1655,N_1192,N_1265);
and U1656 (N_1656,N_1438,N_1058);
nor U1657 (N_1657,N_1164,N_1128);
nor U1658 (N_1658,N_1195,N_1249);
or U1659 (N_1659,N_1324,N_1089);
and U1660 (N_1660,N_1416,N_1086);
or U1661 (N_1661,N_1286,N_1114);
nand U1662 (N_1662,N_1175,N_1489);
and U1663 (N_1663,N_1434,N_1102);
and U1664 (N_1664,N_1303,N_1146);
nand U1665 (N_1665,N_1017,N_1330);
or U1666 (N_1666,N_1491,N_1415);
xnor U1667 (N_1667,N_1371,N_1255);
nand U1668 (N_1668,N_1247,N_1262);
xor U1669 (N_1669,N_1332,N_1342);
xor U1670 (N_1670,N_1106,N_1154);
xnor U1671 (N_1671,N_1408,N_1392);
and U1672 (N_1672,N_1490,N_1140);
and U1673 (N_1673,N_1125,N_1155);
and U1674 (N_1674,N_1455,N_1059);
and U1675 (N_1675,N_1430,N_1015);
xor U1676 (N_1676,N_1470,N_1173);
and U1677 (N_1677,N_1315,N_1348);
xnor U1678 (N_1678,N_1205,N_1073);
xnor U1679 (N_1679,N_1145,N_1456);
nand U1680 (N_1680,N_1432,N_1478);
nor U1681 (N_1681,N_1441,N_1113);
nand U1682 (N_1682,N_1374,N_1098);
and U1683 (N_1683,N_1264,N_1274);
or U1684 (N_1684,N_1447,N_1056);
nor U1685 (N_1685,N_1471,N_1311);
or U1686 (N_1686,N_1349,N_1316);
and U1687 (N_1687,N_1216,N_1010);
or U1688 (N_1688,N_1313,N_1480);
and U1689 (N_1689,N_1023,N_1159);
nand U1690 (N_1690,N_1168,N_1161);
or U1691 (N_1691,N_1172,N_1276);
and U1692 (N_1692,N_1411,N_1228);
or U1693 (N_1693,N_1499,N_1219);
nand U1694 (N_1694,N_1329,N_1229);
and U1695 (N_1695,N_1095,N_1124);
xor U1696 (N_1696,N_1093,N_1020);
nor U1697 (N_1697,N_1338,N_1074);
and U1698 (N_1698,N_1027,N_1131);
xnor U1699 (N_1699,N_1368,N_1452);
or U1700 (N_1700,N_1079,N_1291);
or U1701 (N_1701,N_1398,N_1275);
nand U1702 (N_1702,N_1497,N_1004);
or U1703 (N_1703,N_1305,N_1310);
nor U1704 (N_1704,N_1347,N_1257);
or U1705 (N_1705,N_1469,N_1281);
xnor U1706 (N_1706,N_1008,N_1288);
xor U1707 (N_1707,N_1063,N_1407);
nor U1708 (N_1708,N_1160,N_1343);
or U1709 (N_1709,N_1083,N_1110);
nand U1710 (N_1710,N_1149,N_1042);
nor U1711 (N_1711,N_1322,N_1404);
and U1712 (N_1712,N_1472,N_1047);
and U1713 (N_1713,N_1353,N_1171);
nor U1714 (N_1714,N_1050,N_1496);
and U1715 (N_1715,N_1328,N_1100);
or U1716 (N_1716,N_1035,N_1209);
nand U1717 (N_1717,N_1068,N_1396);
nand U1718 (N_1718,N_1022,N_1096);
xor U1719 (N_1719,N_1306,N_1232);
or U1720 (N_1720,N_1199,N_1380);
nor U1721 (N_1721,N_1182,N_1026);
xnor U1722 (N_1722,N_1049,N_1354);
or U1723 (N_1723,N_1174,N_1151);
and U1724 (N_1724,N_1243,N_1157);
nand U1725 (N_1725,N_1334,N_1389);
and U1726 (N_1726,N_1084,N_1341);
and U1727 (N_1727,N_1256,N_1032);
xnor U1728 (N_1728,N_1123,N_1431);
xor U1729 (N_1729,N_1381,N_1141);
nand U1730 (N_1730,N_1388,N_1028);
nand U1731 (N_1731,N_1233,N_1369);
or U1732 (N_1732,N_1180,N_1237);
and U1733 (N_1733,N_1176,N_1260);
or U1734 (N_1734,N_1225,N_1011);
nor U1735 (N_1735,N_1270,N_1006);
and U1736 (N_1736,N_1194,N_1300);
or U1737 (N_1737,N_1376,N_1136);
or U1738 (N_1738,N_1105,N_1393);
nor U1739 (N_1739,N_1362,N_1366);
nand U1740 (N_1740,N_1333,N_1351);
nor U1741 (N_1741,N_1302,N_1427);
and U1742 (N_1742,N_1285,N_1193);
xnor U1743 (N_1743,N_1296,N_1273);
nand U1744 (N_1744,N_1395,N_1350);
nand U1745 (N_1745,N_1451,N_1177);
nand U1746 (N_1746,N_1422,N_1326);
nor U1747 (N_1747,N_1261,N_1417);
and U1748 (N_1748,N_1473,N_1290);
xor U1749 (N_1749,N_1215,N_1012);
nand U1750 (N_1750,N_1138,N_1478);
xor U1751 (N_1751,N_1049,N_1436);
xnor U1752 (N_1752,N_1479,N_1272);
xor U1753 (N_1753,N_1375,N_1192);
and U1754 (N_1754,N_1106,N_1392);
nand U1755 (N_1755,N_1441,N_1333);
nor U1756 (N_1756,N_1450,N_1187);
nand U1757 (N_1757,N_1360,N_1288);
and U1758 (N_1758,N_1405,N_1282);
nor U1759 (N_1759,N_1290,N_1327);
nand U1760 (N_1760,N_1427,N_1238);
nand U1761 (N_1761,N_1022,N_1293);
nor U1762 (N_1762,N_1497,N_1014);
nand U1763 (N_1763,N_1063,N_1359);
xor U1764 (N_1764,N_1323,N_1373);
or U1765 (N_1765,N_1356,N_1268);
nand U1766 (N_1766,N_1351,N_1446);
nor U1767 (N_1767,N_1267,N_1396);
nor U1768 (N_1768,N_1381,N_1130);
xor U1769 (N_1769,N_1346,N_1446);
xnor U1770 (N_1770,N_1098,N_1362);
nor U1771 (N_1771,N_1497,N_1445);
xnor U1772 (N_1772,N_1442,N_1252);
xor U1773 (N_1773,N_1015,N_1069);
xnor U1774 (N_1774,N_1313,N_1336);
and U1775 (N_1775,N_1393,N_1406);
nor U1776 (N_1776,N_1227,N_1006);
xor U1777 (N_1777,N_1106,N_1114);
nor U1778 (N_1778,N_1477,N_1233);
and U1779 (N_1779,N_1357,N_1146);
nand U1780 (N_1780,N_1365,N_1310);
and U1781 (N_1781,N_1213,N_1193);
nand U1782 (N_1782,N_1289,N_1177);
nand U1783 (N_1783,N_1479,N_1169);
nor U1784 (N_1784,N_1252,N_1332);
nor U1785 (N_1785,N_1281,N_1115);
or U1786 (N_1786,N_1335,N_1101);
xnor U1787 (N_1787,N_1251,N_1187);
or U1788 (N_1788,N_1080,N_1028);
and U1789 (N_1789,N_1088,N_1261);
nor U1790 (N_1790,N_1135,N_1114);
xor U1791 (N_1791,N_1033,N_1434);
and U1792 (N_1792,N_1410,N_1143);
nand U1793 (N_1793,N_1480,N_1390);
nand U1794 (N_1794,N_1337,N_1437);
xnor U1795 (N_1795,N_1217,N_1058);
nor U1796 (N_1796,N_1107,N_1372);
xnor U1797 (N_1797,N_1243,N_1272);
xnor U1798 (N_1798,N_1266,N_1497);
nand U1799 (N_1799,N_1067,N_1298);
xor U1800 (N_1800,N_1085,N_1097);
nor U1801 (N_1801,N_1304,N_1441);
nand U1802 (N_1802,N_1292,N_1088);
xor U1803 (N_1803,N_1189,N_1397);
and U1804 (N_1804,N_1275,N_1168);
nand U1805 (N_1805,N_1192,N_1227);
or U1806 (N_1806,N_1250,N_1039);
nand U1807 (N_1807,N_1349,N_1312);
and U1808 (N_1808,N_1027,N_1070);
xnor U1809 (N_1809,N_1244,N_1094);
nand U1810 (N_1810,N_1326,N_1072);
and U1811 (N_1811,N_1072,N_1482);
xnor U1812 (N_1812,N_1244,N_1210);
or U1813 (N_1813,N_1022,N_1181);
xnor U1814 (N_1814,N_1363,N_1070);
and U1815 (N_1815,N_1211,N_1197);
or U1816 (N_1816,N_1401,N_1221);
and U1817 (N_1817,N_1325,N_1491);
nand U1818 (N_1818,N_1331,N_1100);
nand U1819 (N_1819,N_1214,N_1340);
or U1820 (N_1820,N_1042,N_1452);
and U1821 (N_1821,N_1302,N_1314);
and U1822 (N_1822,N_1079,N_1443);
and U1823 (N_1823,N_1369,N_1267);
or U1824 (N_1824,N_1012,N_1044);
and U1825 (N_1825,N_1225,N_1356);
nand U1826 (N_1826,N_1171,N_1114);
xnor U1827 (N_1827,N_1233,N_1130);
xor U1828 (N_1828,N_1037,N_1060);
or U1829 (N_1829,N_1279,N_1376);
and U1830 (N_1830,N_1266,N_1380);
nand U1831 (N_1831,N_1035,N_1276);
nor U1832 (N_1832,N_1447,N_1136);
nand U1833 (N_1833,N_1117,N_1320);
nor U1834 (N_1834,N_1176,N_1080);
and U1835 (N_1835,N_1035,N_1283);
xnor U1836 (N_1836,N_1367,N_1101);
or U1837 (N_1837,N_1414,N_1412);
xnor U1838 (N_1838,N_1012,N_1225);
and U1839 (N_1839,N_1161,N_1001);
and U1840 (N_1840,N_1499,N_1015);
nor U1841 (N_1841,N_1111,N_1371);
or U1842 (N_1842,N_1233,N_1113);
nand U1843 (N_1843,N_1128,N_1061);
nand U1844 (N_1844,N_1281,N_1332);
and U1845 (N_1845,N_1067,N_1431);
and U1846 (N_1846,N_1315,N_1397);
nand U1847 (N_1847,N_1376,N_1318);
nor U1848 (N_1848,N_1079,N_1404);
and U1849 (N_1849,N_1472,N_1100);
or U1850 (N_1850,N_1295,N_1079);
and U1851 (N_1851,N_1197,N_1087);
xor U1852 (N_1852,N_1254,N_1281);
nor U1853 (N_1853,N_1299,N_1415);
xnor U1854 (N_1854,N_1056,N_1482);
or U1855 (N_1855,N_1158,N_1086);
nor U1856 (N_1856,N_1183,N_1252);
and U1857 (N_1857,N_1343,N_1428);
or U1858 (N_1858,N_1441,N_1187);
nand U1859 (N_1859,N_1018,N_1253);
xor U1860 (N_1860,N_1315,N_1141);
xnor U1861 (N_1861,N_1173,N_1144);
and U1862 (N_1862,N_1451,N_1010);
nor U1863 (N_1863,N_1264,N_1355);
xnor U1864 (N_1864,N_1087,N_1170);
xor U1865 (N_1865,N_1198,N_1032);
xnor U1866 (N_1866,N_1074,N_1053);
xnor U1867 (N_1867,N_1073,N_1055);
and U1868 (N_1868,N_1165,N_1498);
or U1869 (N_1869,N_1223,N_1092);
nand U1870 (N_1870,N_1284,N_1128);
and U1871 (N_1871,N_1223,N_1047);
xnor U1872 (N_1872,N_1051,N_1090);
xor U1873 (N_1873,N_1052,N_1192);
nor U1874 (N_1874,N_1280,N_1464);
nor U1875 (N_1875,N_1262,N_1328);
xnor U1876 (N_1876,N_1101,N_1274);
or U1877 (N_1877,N_1125,N_1198);
or U1878 (N_1878,N_1150,N_1228);
xnor U1879 (N_1879,N_1354,N_1291);
xor U1880 (N_1880,N_1391,N_1119);
and U1881 (N_1881,N_1377,N_1285);
nor U1882 (N_1882,N_1293,N_1289);
nor U1883 (N_1883,N_1035,N_1036);
and U1884 (N_1884,N_1224,N_1264);
and U1885 (N_1885,N_1059,N_1318);
and U1886 (N_1886,N_1406,N_1196);
xor U1887 (N_1887,N_1342,N_1383);
xor U1888 (N_1888,N_1331,N_1191);
nand U1889 (N_1889,N_1065,N_1132);
and U1890 (N_1890,N_1495,N_1082);
nor U1891 (N_1891,N_1450,N_1018);
nand U1892 (N_1892,N_1403,N_1113);
or U1893 (N_1893,N_1176,N_1249);
nor U1894 (N_1894,N_1195,N_1265);
xor U1895 (N_1895,N_1050,N_1448);
nand U1896 (N_1896,N_1342,N_1435);
nand U1897 (N_1897,N_1128,N_1250);
nor U1898 (N_1898,N_1331,N_1358);
or U1899 (N_1899,N_1224,N_1463);
nand U1900 (N_1900,N_1271,N_1064);
nor U1901 (N_1901,N_1306,N_1050);
and U1902 (N_1902,N_1020,N_1261);
and U1903 (N_1903,N_1452,N_1353);
xor U1904 (N_1904,N_1011,N_1137);
and U1905 (N_1905,N_1186,N_1245);
nor U1906 (N_1906,N_1227,N_1415);
nand U1907 (N_1907,N_1094,N_1319);
and U1908 (N_1908,N_1247,N_1304);
nand U1909 (N_1909,N_1011,N_1133);
and U1910 (N_1910,N_1273,N_1170);
or U1911 (N_1911,N_1203,N_1189);
or U1912 (N_1912,N_1150,N_1022);
or U1913 (N_1913,N_1030,N_1437);
xor U1914 (N_1914,N_1103,N_1008);
nand U1915 (N_1915,N_1274,N_1242);
nor U1916 (N_1916,N_1146,N_1306);
or U1917 (N_1917,N_1266,N_1463);
xnor U1918 (N_1918,N_1338,N_1133);
nor U1919 (N_1919,N_1012,N_1323);
xnor U1920 (N_1920,N_1451,N_1311);
nor U1921 (N_1921,N_1233,N_1434);
xor U1922 (N_1922,N_1399,N_1252);
and U1923 (N_1923,N_1092,N_1411);
xor U1924 (N_1924,N_1420,N_1221);
nor U1925 (N_1925,N_1353,N_1352);
or U1926 (N_1926,N_1414,N_1337);
nand U1927 (N_1927,N_1450,N_1026);
nand U1928 (N_1928,N_1264,N_1079);
nand U1929 (N_1929,N_1458,N_1011);
and U1930 (N_1930,N_1483,N_1445);
or U1931 (N_1931,N_1127,N_1470);
and U1932 (N_1932,N_1275,N_1087);
and U1933 (N_1933,N_1446,N_1100);
xor U1934 (N_1934,N_1237,N_1035);
nand U1935 (N_1935,N_1009,N_1071);
and U1936 (N_1936,N_1466,N_1454);
or U1937 (N_1937,N_1188,N_1307);
nand U1938 (N_1938,N_1381,N_1008);
or U1939 (N_1939,N_1224,N_1474);
nor U1940 (N_1940,N_1391,N_1420);
nor U1941 (N_1941,N_1324,N_1379);
xnor U1942 (N_1942,N_1459,N_1122);
xnor U1943 (N_1943,N_1435,N_1120);
xnor U1944 (N_1944,N_1261,N_1243);
nand U1945 (N_1945,N_1275,N_1254);
nand U1946 (N_1946,N_1051,N_1219);
and U1947 (N_1947,N_1270,N_1418);
nand U1948 (N_1948,N_1043,N_1368);
and U1949 (N_1949,N_1288,N_1258);
nand U1950 (N_1950,N_1322,N_1432);
and U1951 (N_1951,N_1403,N_1276);
or U1952 (N_1952,N_1285,N_1414);
xnor U1953 (N_1953,N_1498,N_1467);
and U1954 (N_1954,N_1456,N_1394);
or U1955 (N_1955,N_1383,N_1124);
nor U1956 (N_1956,N_1259,N_1415);
and U1957 (N_1957,N_1094,N_1399);
or U1958 (N_1958,N_1092,N_1242);
nor U1959 (N_1959,N_1352,N_1093);
nor U1960 (N_1960,N_1463,N_1319);
xnor U1961 (N_1961,N_1233,N_1129);
xnor U1962 (N_1962,N_1290,N_1016);
nor U1963 (N_1963,N_1276,N_1116);
nand U1964 (N_1964,N_1429,N_1412);
nor U1965 (N_1965,N_1300,N_1258);
or U1966 (N_1966,N_1071,N_1175);
nor U1967 (N_1967,N_1288,N_1331);
xnor U1968 (N_1968,N_1088,N_1063);
and U1969 (N_1969,N_1108,N_1158);
or U1970 (N_1970,N_1196,N_1054);
and U1971 (N_1971,N_1321,N_1186);
or U1972 (N_1972,N_1471,N_1175);
and U1973 (N_1973,N_1005,N_1265);
xnor U1974 (N_1974,N_1223,N_1211);
nor U1975 (N_1975,N_1072,N_1008);
and U1976 (N_1976,N_1296,N_1137);
xor U1977 (N_1977,N_1231,N_1298);
nor U1978 (N_1978,N_1090,N_1290);
xor U1979 (N_1979,N_1077,N_1043);
nor U1980 (N_1980,N_1391,N_1029);
nor U1981 (N_1981,N_1277,N_1180);
nor U1982 (N_1982,N_1393,N_1029);
or U1983 (N_1983,N_1287,N_1219);
nand U1984 (N_1984,N_1137,N_1124);
nand U1985 (N_1985,N_1155,N_1226);
xnor U1986 (N_1986,N_1288,N_1020);
and U1987 (N_1987,N_1087,N_1186);
xnor U1988 (N_1988,N_1303,N_1176);
nor U1989 (N_1989,N_1166,N_1010);
or U1990 (N_1990,N_1041,N_1211);
or U1991 (N_1991,N_1157,N_1232);
or U1992 (N_1992,N_1476,N_1195);
and U1993 (N_1993,N_1243,N_1317);
nor U1994 (N_1994,N_1154,N_1313);
nand U1995 (N_1995,N_1442,N_1140);
nor U1996 (N_1996,N_1178,N_1240);
or U1997 (N_1997,N_1198,N_1055);
nor U1998 (N_1998,N_1005,N_1040);
nand U1999 (N_1999,N_1161,N_1383);
and U2000 (N_2000,N_1993,N_1520);
xnor U2001 (N_2001,N_1941,N_1513);
nor U2002 (N_2002,N_1543,N_1646);
nor U2003 (N_2003,N_1874,N_1923);
and U2004 (N_2004,N_1668,N_1783);
or U2005 (N_2005,N_1722,N_1908);
xor U2006 (N_2006,N_1557,N_1804);
nor U2007 (N_2007,N_1859,N_1829);
nor U2008 (N_2008,N_1630,N_1634);
xnor U2009 (N_2009,N_1761,N_1961);
and U2010 (N_2010,N_1575,N_1744);
and U2011 (N_2011,N_1774,N_1778);
nor U2012 (N_2012,N_1702,N_1883);
nand U2013 (N_2013,N_1955,N_1951);
and U2014 (N_2014,N_1759,N_1680);
or U2015 (N_2015,N_1810,N_1544);
or U2016 (N_2016,N_1986,N_1850);
or U2017 (N_2017,N_1747,N_1773);
nor U2018 (N_2018,N_1568,N_1943);
or U2019 (N_2019,N_1755,N_1864);
nor U2020 (N_2020,N_1640,N_1801);
xor U2021 (N_2021,N_1511,N_1589);
or U2022 (N_2022,N_1972,N_1622);
nor U2023 (N_2023,N_1796,N_1518);
xor U2024 (N_2024,N_1645,N_1765);
or U2025 (N_2025,N_1992,N_1816);
nand U2026 (N_2026,N_1522,N_1756);
or U2027 (N_2027,N_1927,N_1907);
or U2028 (N_2028,N_1667,N_1949);
xor U2029 (N_2029,N_1635,N_1736);
nand U2030 (N_2030,N_1670,N_1619);
nand U2031 (N_2031,N_1509,N_1721);
and U2032 (N_2032,N_1987,N_1866);
nand U2033 (N_2033,N_1613,N_1904);
nor U2034 (N_2034,N_1659,N_1561);
nand U2035 (N_2035,N_1838,N_1662);
nand U2036 (N_2036,N_1612,N_1983);
xnor U2037 (N_2037,N_1694,N_1922);
xor U2038 (N_2038,N_1775,N_1894);
or U2039 (N_2039,N_1593,N_1728);
and U2040 (N_2040,N_1914,N_1909);
xor U2041 (N_2041,N_1639,N_1696);
or U2042 (N_2042,N_1934,N_1512);
and U2043 (N_2043,N_1614,N_1517);
nand U2044 (N_2044,N_1760,N_1689);
xor U2045 (N_2045,N_1935,N_1800);
or U2046 (N_2046,N_1821,N_1879);
xor U2047 (N_2047,N_1998,N_1686);
or U2048 (N_2048,N_1808,N_1881);
nor U2049 (N_2049,N_1631,N_1552);
nor U2050 (N_2050,N_1558,N_1835);
nor U2051 (N_2051,N_1900,N_1878);
xor U2052 (N_2052,N_1989,N_1959);
nor U2053 (N_2053,N_1936,N_1601);
nand U2054 (N_2054,N_1726,N_1527);
nand U2055 (N_2055,N_1582,N_1805);
xor U2056 (N_2056,N_1764,N_1576);
nor U2057 (N_2057,N_1691,N_1658);
or U2058 (N_2058,N_1807,N_1929);
nor U2059 (N_2059,N_1855,N_1621);
xor U2060 (N_2060,N_1750,N_1771);
xor U2061 (N_2061,N_1820,N_1629);
or U2062 (N_2062,N_1610,N_1617);
and U2063 (N_2063,N_1873,N_1566);
nor U2064 (N_2064,N_1585,N_1792);
nand U2065 (N_2065,N_1982,N_1584);
and U2066 (N_2066,N_1845,N_1533);
nor U2067 (N_2067,N_1597,N_1657);
nand U2068 (N_2068,N_1681,N_1768);
and U2069 (N_2069,N_1731,N_1594);
xor U2070 (N_2070,N_1931,N_1570);
nor U2071 (N_2071,N_1892,N_1997);
or U2072 (N_2072,N_1548,N_1916);
or U2073 (N_2073,N_1673,N_1841);
nand U2074 (N_2074,N_1574,N_1860);
xnor U2075 (N_2075,N_1797,N_1872);
and U2076 (N_2076,N_1648,N_1770);
xnor U2077 (N_2077,N_1595,N_1508);
and U2078 (N_2078,N_1779,N_1615);
or U2079 (N_2079,N_1620,N_1708);
and U2080 (N_2080,N_1896,N_1812);
nand U2081 (N_2081,N_1870,N_1814);
nor U2082 (N_2082,N_1551,N_1823);
xnor U2083 (N_2083,N_1793,N_1709);
xnor U2084 (N_2084,N_1910,N_1724);
xnor U2085 (N_2085,N_1868,N_1514);
xnor U2086 (N_2086,N_1633,N_1573);
or U2087 (N_2087,N_1787,N_1735);
nand U2088 (N_2088,N_1880,N_1976);
and U2089 (N_2089,N_1828,N_1505);
nor U2090 (N_2090,N_1857,N_1791);
nor U2091 (N_2091,N_1966,N_1684);
or U2092 (N_2092,N_1833,N_1827);
and U2093 (N_2093,N_1685,N_1580);
xnor U2094 (N_2094,N_1628,N_1919);
nand U2095 (N_2095,N_1515,N_1598);
nor U2096 (N_2096,N_1882,N_1831);
or U2097 (N_2097,N_1697,N_1886);
and U2098 (N_2098,N_1893,N_1785);
nand U2099 (N_2099,N_1939,N_1741);
or U2100 (N_2100,N_1984,N_1901);
and U2101 (N_2101,N_1587,N_1999);
nand U2102 (N_2102,N_1913,N_1803);
xnor U2103 (N_2103,N_1863,N_1743);
xnor U2104 (N_2104,N_1780,N_1665);
nor U2105 (N_2105,N_1707,N_1825);
xnor U2106 (N_2106,N_1649,N_1849);
and U2107 (N_2107,N_1592,N_1839);
xnor U2108 (N_2108,N_1539,N_1826);
nand U2109 (N_2109,N_1607,N_1677);
or U2110 (N_2110,N_1946,N_1819);
nor U2111 (N_2111,N_1562,N_1799);
or U2112 (N_2112,N_1525,N_1813);
xor U2113 (N_2113,N_1565,N_1895);
nor U2114 (N_2114,N_1956,N_1748);
or U2115 (N_2115,N_1944,N_1704);
nor U2116 (N_2116,N_1618,N_1578);
nand U2117 (N_2117,N_1830,N_1650);
nor U2118 (N_2118,N_1542,N_1516);
nand U2119 (N_2119,N_1546,N_1683);
xor U2120 (N_2120,N_1671,N_1504);
xor U2121 (N_2121,N_1917,N_1811);
nand U2122 (N_2122,N_1798,N_1746);
and U2123 (N_2123,N_1611,N_1887);
xor U2124 (N_2124,N_1660,N_1865);
nor U2125 (N_2125,N_1847,N_1824);
nand U2126 (N_2126,N_1753,N_1651);
or U2127 (N_2127,N_1716,N_1563);
or U2128 (N_2128,N_1979,N_1794);
xnor U2129 (N_2129,N_1626,N_1769);
and U2130 (N_2130,N_1818,N_1790);
xnor U2131 (N_2131,N_1925,N_1950);
and U2132 (N_2132,N_1862,N_1763);
xnor U2133 (N_2133,N_1609,N_1625);
or U2134 (N_2134,N_1559,N_1523);
and U2135 (N_2135,N_1682,N_1711);
or U2136 (N_2136,N_1877,N_1837);
or U2137 (N_2137,N_1653,N_1906);
xnor U2138 (N_2138,N_1898,N_1688);
nand U2139 (N_2139,N_1588,N_1861);
nor U2140 (N_2140,N_1752,N_1905);
and U2141 (N_2141,N_1699,N_1899);
or U2142 (N_2142,N_1530,N_1500);
and U2143 (N_2143,N_1842,N_1643);
nor U2144 (N_2144,N_1749,N_1714);
xnor U2145 (N_2145,N_1738,N_1742);
and U2146 (N_2146,N_1532,N_1933);
or U2147 (N_2147,N_1911,N_1836);
or U2148 (N_2148,N_1990,N_1586);
xor U2149 (N_2149,N_1676,N_1591);
xnor U2150 (N_2150,N_1767,N_1975);
nand U2151 (N_2151,N_1817,N_1854);
xor U2152 (N_2152,N_1981,N_1772);
xor U2153 (N_2153,N_1550,N_1687);
nand U2154 (N_2154,N_1510,N_1926);
nand U2155 (N_2155,N_1977,N_1579);
xnor U2156 (N_2156,N_1739,N_1554);
and U2157 (N_2157,N_1915,N_1656);
and U2158 (N_2158,N_1788,N_1953);
or U2159 (N_2159,N_1603,N_1534);
xor U2160 (N_2160,N_1705,N_1781);
xnor U2161 (N_2161,N_1506,N_1891);
or U2162 (N_2162,N_1718,N_1560);
and U2163 (N_2163,N_1885,N_1641);
and U2164 (N_2164,N_1784,N_1786);
nand U2165 (N_2165,N_1531,N_1663);
and U2166 (N_2166,N_1745,N_1669);
or U2167 (N_2167,N_1583,N_1572);
xor U2168 (N_2168,N_1642,N_1867);
nand U2169 (N_2169,N_1832,N_1690);
xor U2170 (N_2170,N_1535,N_1802);
or U2171 (N_2171,N_1871,N_1567);
xor U2172 (N_2172,N_1678,N_1930);
nand U2173 (N_2173,N_1942,N_1856);
nor U2174 (N_2174,N_1876,N_1632);
or U2175 (N_2175,N_1590,N_1757);
nand U2176 (N_2176,N_1693,N_1529);
nand U2177 (N_2177,N_1608,N_1853);
xor U2178 (N_2178,N_1957,N_1924);
nand U2179 (N_2179,N_1890,N_1692);
and U2180 (N_2180,N_1541,N_1666);
or U2181 (N_2181,N_1652,N_1852);
xor U2182 (N_2182,N_1606,N_1902);
nor U2183 (N_2183,N_1991,N_1577);
and U2184 (N_2184,N_1889,N_1655);
nor U2185 (N_2185,N_1888,N_1549);
nand U2186 (N_2186,N_1701,N_1884);
nor U2187 (N_2187,N_1675,N_1994);
nand U2188 (N_2188,N_1912,N_1754);
or U2189 (N_2189,N_1985,N_1644);
nand U2190 (N_2190,N_1964,N_1932);
xor U2191 (N_2191,N_1623,N_1553);
and U2192 (N_2192,N_1875,N_1903);
nand U2193 (N_2193,N_1920,N_1737);
nand U2194 (N_2194,N_1851,N_1848);
nand U2195 (N_2195,N_1637,N_1978);
or U2196 (N_2196,N_1730,N_1602);
or U2197 (N_2197,N_1782,N_1717);
nor U2198 (N_2198,N_1967,N_1937);
nand U2199 (N_2199,N_1526,N_1815);
or U2200 (N_2200,N_1713,N_1661);
nor U2201 (N_2201,N_1538,N_1564);
or U2202 (N_2202,N_1858,N_1970);
or U2203 (N_2203,N_1928,N_1703);
nand U2204 (N_2204,N_1501,N_1725);
or U2205 (N_2205,N_1869,N_1948);
or U2206 (N_2206,N_1507,N_1806);
or U2207 (N_2207,N_1674,N_1624);
nor U2208 (N_2208,N_1740,N_1581);
nand U2209 (N_2209,N_1995,N_1664);
or U2210 (N_2210,N_1844,N_1596);
nand U2211 (N_2211,N_1766,N_1555);
and U2212 (N_2212,N_1973,N_1758);
and U2213 (N_2213,N_1695,N_1988);
and U2214 (N_2214,N_1996,N_1654);
or U2215 (N_2215,N_1751,N_1502);
and U2216 (N_2216,N_1547,N_1762);
or U2217 (N_2217,N_1834,N_1599);
and U2218 (N_2218,N_1536,N_1647);
nand U2219 (N_2219,N_1729,N_1777);
nor U2220 (N_2220,N_1947,N_1727);
nand U2221 (N_2221,N_1960,N_1720);
nor U2222 (N_2222,N_1706,N_1734);
and U2223 (N_2223,N_1846,N_1776);
xnor U2224 (N_2224,N_1969,N_1897);
xnor U2225 (N_2225,N_1954,N_1712);
nand U2226 (N_2226,N_1503,N_1945);
or U2227 (N_2227,N_1822,N_1719);
nor U2228 (N_2228,N_1809,N_1918);
nor U2229 (N_2229,N_1958,N_1605);
or U2230 (N_2230,N_1638,N_1840);
nand U2231 (N_2231,N_1938,N_1698);
nand U2232 (N_2232,N_1962,N_1528);
nor U2233 (N_2233,N_1974,N_1545);
and U2234 (N_2234,N_1980,N_1965);
xor U2235 (N_2235,N_1733,N_1569);
xor U2236 (N_2236,N_1710,N_1571);
and U2237 (N_2237,N_1940,N_1968);
xor U2238 (N_2238,N_1732,N_1789);
xnor U2239 (N_2239,N_1921,N_1971);
nand U2240 (N_2240,N_1636,N_1723);
nor U2241 (N_2241,N_1672,N_1700);
nand U2242 (N_2242,N_1519,N_1600);
nand U2243 (N_2243,N_1556,N_1679);
xor U2244 (N_2244,N_1537,N_1604);
xnor U2245 (N_2245,N_1540,N_1521);
xor U2246 (N_2246,N_1524,N_1843);
nor U2247 (N_2247,N_1963,N_1715);
nor U2248 (N_2248,N_1627,N_1616);
xor U2249 (N_2249,N_1952,N_1795);
nand U2250 (N_2250,N_1787,N_1936);
xor U2251 (N_2251,N_1792,N_1885);
nor U2252 (N_2252,N_1851,N_1963);
nor U2253 (N_2253,N_1517,N_1978);
or U2254 (N_2254,N_1682,N_1964);
xor U2255 (N_2255,N_1898,N_1643);
nor U2256 (N_2256,N_1571,N_1517);
and U2257 (N_2257,N_1756,N_1578);
nor U2258 (N_2258,N_1613,N_1746);
and U2259 (N_2259,N_1721,N_1832);
nand U2260 (N_2260,N_1865,N_1621);
nor U2261 (N_2261,N_1850,N_1774);
nor U2262 (N_2262,N_1800,N_1584);
or U2263 (N_2263,N_1966,N_1885);
xnor U2264 (N_2264,N_1603,N_1521);
xor U2265 (N_2265,N_1813,N_1880);
and U2266 (N_2266,N_1755,N_1742);
xor U2267 (N_2267,N_1836,N_1738);
and U2268 (N_2268,N_1710,N_1583);
or U2269 (N_2269,N_1690,N_1737);
or U2270 (N_2270,N_1592,N_1618);
xnor U2271 (N_2271,N_1836,N_1725);
nor U2272 (N_2272,N_1781,N_1872);
nor U2273 (N_2273,N_1959,N_1853);
or U2274 (N_2274,N_1777,N_1588);
nor U2275 (N_2275,N_1501,N_1830);
xnor U2276 (N_2276,N_1634,N_1505);
xnor U2277 (N_2277,N_1500,N_1872);
xnor U2278 (N_2278,N_1958,N_1761);
nor U2279 (N_2279,N_1706,N_1503);
nor U2280 (N_2280,N_1571,N_1663);
nor U2281 (N_2281,N_1882,N_1926);
nand U2282 (N_2282,N_1728,N_1813);
or U2283 (N_2283,N_1574,N_1927);
or U2284 (N_2284,N_1565,N_1648);
nand U2285 (N_2285,N_1749,N_1621);
or U2286 (N_2286,N_1783,N_1931);
nand U2287 (N_2287,N_1510,N_1761);
nand U2288 (N_2288,N_1978,N_1653);
or U2289 (N_2289,N_1825,N_1889);
or U2290 (N_2290,N_1957,N_1642);
nand U2291 (N_2291,N_1960,N_1980);
and U2292 (N_2292,N_1621,N_1996);
or U2293 (N_2293,N_1814,N_1950);
and U2294 (N_2294,N_1595,N_1900);
or U2295 (N_2295,N_1859,N_1816);
xor U2296 (N_2296,N_1516,N_1782);
or U2297 (N_2297,N_1579,N_1578);
and U2298 (N_2298,N_1682,N_1809);
nor U2299 (N_2299,N_1766,N_1687);
or U2300 (N_2300,N_1838,N_1642);
nand U2301 (N_2301,N_1640,N_1963);
and U2302 (N_2302,N_1914,N_1704);
nor U2303 (N_2303,N_1569,N_1910);
xnor U2304 (N_2304,N_1721,N_1564);
or U2305 (N_2305,N_1729,N_1670);
nor U2306 (N_2306,N_1587,N_1589);
nand U2307 (N_2307,N_1947,N_1746);
and U2308 (N_2308,N_1923,N_1706);
or U2309 (N_2309,N_1715,N_1748);
and U2310 (N_2310,N_1572,N_1940);
nand U2311 (N_2311,N_1961,N_1709);
nand U2312 (N_2312,N_1723,N_1820);
and U2313 (N_2313,N_1864,N_1554);
xor U2314 (N_2314,N_1754,N_1702);
or U2315 (N_2315,N_1752,N_1567);
or U2316 (N_2316,N_1539,N_1814);
nand U2317 (N_2317,N_1696,N_1982);
nand U2318 (N_2318,N_1733,N_1909);
nand U2319 (N_2319,N_1563,N_1782);
or U2320 (N_2320,N_1690,N_1512);
or U2321 (N_2321,N_1761,N_1789);
nor U2322 (N_2322,N_1697,N_1565);
nand U2323 (N_2323,N_1726,N_1625);
and U2324 (N_2324,N_1592,N_1997);
or U2325 (N_2325,N_1643,N_1559);
nor U2326 (N_2326,N_1773,N_1739);
and U2327 (N_2327,N_1661,N_1863);
xnor U2328 (N_2328,N_1874,N_1639);
xnor U2329 (N_2329,N_1507,N_1727);
or U2330 (N_2330,N_1800,N_1741);
or U2331 (N_2331,N_1940,N_1552);
or U2332 (N_2332,N_1853,N_1657);
and U2333 (N_2333,N_1535,N_1646);
nor U2334 (N_2334,N_1619,N_1998);
nand U2335 (N_2335,N_1509,N_1668);
xnor U2336 (N_2336,N_1514,N_1539);
nor U2337 (N_2337,N_1632,N_1554);
nor U2338 (N_2338,N_1850,N_1625);
nand U2339 (N_2339,N_1855,N_1682);
nor U2340 (N_2340,N_1624,N_1637);
and U2341 (N_2341,N_1997,N_1553);
and U2342 (N_2342,N_1743,N_1972);
or U2343 (N_2343,N_1888,N_1692);
nor U2344 (N_2344,N_1652,N_1700);
xor U2345 (N_2345,N_1999,N_1808);
or U2346 (N_2346,N_1890,N_1985);
or U2347 (N_2347,N_1871,N_1606);
or U2348 (N_2348,N_1551,N_1526);
and U2349 (N_2349,N_1945,N_1950);
xnor U2350 (N_2350,N_1877,N_1676);
xnor U2351 (N_2351,N_1701,N_1704);
nand U2352 (N_2352,N_1996,N_1898);
xor U2353 (N_2353,N_1582,N_1937);
nand U2354 (N_2354,N_1574,N_1924);
and U2355 (N_2355,N_1885,N_1802);
xor U2356 (N_2356,N_1873,N_1516);
nand U2357 (N_2357,N_1536,N_1788);
xor U2358 (N_2358,N_1752,N_1808);
or U2359 (N_2359,N_1987,N_1705);
and U2360 (N_2360,N_1849,N_1964);
nor U2361 (N_2361,N_1511,N_1887);
nor U2362 (N_2362,N_1869,N_1627);
nand U2363 (N_2363,N_1607,N_1525);
nor U2364 (N_2364,N_1829,N_1512);
xor U2365 (N_2365,N_1586,N_1885);
nor U2366 (N_2366,N_1841,N_1552);
or U2367 (N_2367,N_1825,N_1631);
nor U2368 (N_2368,N_1993,N_1913);
xnor U2369 (N_2369,N_1729,N_1697);
xnor U2370 (N_2370,N_1999,N_1726);
xnor U2371 (N_2371,N_1998,N_1669);
nand U2372 (N_2372,N_1771,N_1939);
nor U2373 (N_2373,N_1988,N_1722);
nand U2374 (N_2374,N_1920,N_1536);
and U2375 (N_2375,N_1756,N_1773);
nor U2376 (N_2376,N_1956,N_1857);
xnor U2377 (N_2377,N_1968,N_1552);
and U2378 (N_2378,N_1929,N_1587);
xor U2379 (N_2379,N_1979,N_1709);
nor U2380 (N_2380,N_1651,N_1884);
or U2381 (N_2381,N_1564,N_1935);
nor U2382 (N_2382,N_1884,N_1915);
and U2383 (N_2383,N_1591,N_1516);
or U2384 (N_2384,N_1785,N_1872);
nor U2385 (N_2385,N_1565,N_1877);
xor U2386 (N_2386,N_1615,N_1912);
nand U2387 (N_2387,N_1679,N_1993);
nand U2388 (N_2388,N_1709,N_1513);
and U2389 (N_2389,N_1705,N_1999);
or U2390 (N_2390,N_1645,N_1921);
xor U2391 (N_2391,N_1708,N_1823);
or U2392 (N_2392,N_1753,N_1734);
and U2393 (N_2393,N_1992,N_1546);
nor U2394 (N_2394,N_1519,N_1937);
xnor U2395 (N_2395,N_1543,N_1766);
nand U2396 (N_2396,N_1866,N_1533);
nand U2397 (N_2397,N_1643,N_1522);
and U2398 (N_2398,N_1679,N_1673);
nor U2399 (N_2399,N_1709,N_1757);
or U2400 (N_2400,N_1582,N_1680);
xor U2401 (N_2401,N_1742,N_1588);
or U2402 (N_2402,N_1995,N_1804);
and U2403 (N_2403,N_1782,N_1890);
xor U2404 (N_2404,N_1725,N_1977);
nor U2405 (N_2405,N_1587,N_1734);
and U2406 (N_2406,N_1968,N_1854);
nor U2407 (N_2407,N_1682,N_1975);
xor U2408 (N_2408,N_1513,N_1925);
nand U2409 (N_2409,N_1865,N_1616);
nor U2410 (N_2410,N_1540,N_1626);
xor U2411 (N_2411,N_1731,N_1622);
and U2412 (N_2412,N_1950,N_1702);
xor U2413 (N_2413,N_1958,N_1520);
xor U2414 (N_2414,N_1745,N_1541);
xor U2415 (N_2415,N_1984,N_1966);
and U2416 (N_2416,N_1710,N_1825);
nand U2417 (N_2417,N_1767,N_1698);
xnor U2418 (N_2418,N_1558,N_1524);
nand U2419 (N_2419,N_1577,N_1937);
and U2420 (N_2420,N_1735,N_1758);
nor U2421 (N_2421,N_1967,N_1582);
or U2422 (N_2422,N_1791,N_1511);
or U2423 (N_2423,N_1904,N_1822);
nand U2424 (N_2424,N_1701,N_1802);
or U2425 (N_2425,N_1895,N_1795);
and U2426 (N_2426,N_1952,N_1976);
nand U2427 (N_2427,N_1901,N_1593);
nand U2428 (N_2428,N_1781,N_1544);
xnor U2429 (N_2429,N_1803,N_1795);
or U2430 (N_2430,N_1808,N_1592);
xnor U2431 (N_2431,N_1770,N_1941);
xor U2432 (N_2432,N_1915,N_1741);
xnor U2433 (N_2433,N_1624,N_1867);
or U2434 (N_2434,N_1838,N_1994);
xor U2435 (N_2435,N_1695,N_1888);
nand U2436 (N_2436,N_1986,N_1655);
nand U2437 (N_2437,N_1857,N_1606);
and U2438 (N_2438,N_1513,N_1963);
or U2439 (N_2439,N_1977,N_1777);
xnor U2440 (N_2440,N_1658,N_1576);
or U2441 (N_2441,N_1925,N_1983);
xnor U2442 (N_2442,N_1693,N_1766);
nand U2443 (N_2443,N_1757,N_1644);
and U2444 (N_2444,N_1580,N_1613);
and U2445 (N_2445,N_1621,N_1746);
and U2446 (N_2446,N_1837,N_1566);
nor U2447 (N_2447,N_1537,N_1617);
or U2448 (N_2448,N_1546,N_1595);
xnor U2449 (N_2449,N_1916,N_1906);
and U2450 (N_2450,N_1739,N_1987);
nor U2451 (N_2451,N_1762,N_1795);
or U2452 (N_2452,N_1633,N_1896);
xnor U2453 (N_2453,N_1518,N_1500);
and U2454 (N_2454,N_1727,N_1723);
or U2455 (N_2455,N_1815,N_1823);
nor U2456 (N_2456,N_1672,N_1729);
nand U2457 (N_2457,N_1668,N_1955);
nor U2458 (N_2458,N_1902,N_1880);
or U2459 (N_2459,N_1911,N_1689);
xor U2460 (N_2460,N_1824,N_1760);
or U2461 (N_2461,N_1911,N_1824);
and U2462 (N_2462,N_1923,N_1607);
and U2463 (N_2463,N_1561,N_1860);
and U2464 (N_2464,N_1651,N_1994);
or U2465 (N_2465,N_1993,N_1557);
or U2466 (N_2466,N_1658,N_1624);
nand U2467 (N_2467,N_1995,N_1795);
or U2468 (N_2468,N_1597,N_1861);
or U2469 (N_2469,N_1839,N_1923);
nor U2470 (N_2470,N_1646,N_1717);
nand U2471 (N_2471,N_1861,N_1878);
nand U2472 (N_2472,N_1502,N_1947);
nand U2473 (N_2473,N_1836,N_1932);
or U2474 (N_2474,N_1959,N_1600);
nor U2475 (N_2475,N_1577,N_1570);
and U2476 (N_2476,N_1715,N_1949);
or U2477 (N_2477,N_1724,N_1803);
xnor U2478 (N_2478,N_1986,N_1849);
xnor U2479 (N_2479,N_1541,N_1995);
xor U2480 (N_2480,N_1822,N_1981);
xnor U2481 (N_2481,N_1716,N_1779);
nand U2482 (N_2482,N_1592,N_1718);
nor U2483 (N_2483,N_1810,N_1761);
nor U2484 (N_2484,N_1635,N_1992);
xnor U2485 (N_2485,N_1798,N_1800);
xor U2486 (N_2486,N_1740,N_1619);
xor U2487 (N_2487,N_1696,N_1677);
xor U2488 (N_2488,N_1626,N_1793);
nor U2489 (N_2489,N_1815,N_1938);
xnor U2490 (N_2490,N_1652,N_1955);
nor U2491 (N_2491,N_1689,N_1756);
nand U2492 (N_2492,N_1961,N_1546);
and U2493 (N_2493,N_1875,N_1581);
nand U2494 (N_2494,N_1728,N_1674);
nor U2495 (N_2495,N_1873,N_1661);
and U2496 (N_2496,N_1935,N_1895);
nand U2497 (N_2497,N_1989,N_1701);
and U2498 (N_2498,N_1500,N_1803);
and U2499 (N_2499,N_1509,N_1860);
or U2500 (N_2500,N_2464,N_2346);
and U2501 (N_2501,N_2202,N_2310);
or U2502 (N_2502,N_2008,N_2475);
nor U2503 (N_2503,N_2342,N_2438);
and U2504 (N_2504,N_2183,N_2326);
or U2505 (N_2505,N_2457,N_2292);
and U2506 (N_2506,N_2124,N_2200);
and U2507 (N_2507,N_2481,N_2482);
xnor U2508 (N_2508,N_2397,N_2434);
and U2509 (N_2509,N_2013,N_2067);
nor U2510 (N_2510,N_2432,N_2233);
xnor U2511 (N_2511,N_2250,N_2360);
nor U2512 (N_2512,N_2171,N_2366);
or U2513 (N_2513,N_2450,N_2204);
and U2514 (N_2514,N_2092,N_2393);
nand U2515 (N_2515,N_2042,N_2452);
and U2516 (N_2516,N_2084,N_2428);
xnor U2517 (N_2517,N_2251,N_2206);
xnor U2518 (N_2518,N_2178,N_2441);
or U2519 (N_2519,N_2037,N_2080);
nor U2520 (N_2520,N_2291,N_2036);
or U2521 (N_2521,N_2299,N_2297);
or U2522 (N_2522,N_2137,N_2352);
xnor U2523 (N_2523,N_2105,N_2261);
xor U2524 (N_2524,N_2378,N_2485);
nand U2525 (N_2525,N_2316,N_2284);
or U2526 (N_2526,N_2295,N_2093);
xnor U2527 (N_2527,N_2417,N_2309);
or U2528 (N_2528,N_2319,N_2440);
xor U2529 (N_2529,N_2391,N_2235);
nand U2530 (N_2530,N_2061,N_2083);
or U2531 (N_2531,N_2079,N_2329);
xnor U2532 (N_2532,N_2275,N_2418);
nand U2533 (N_2533,N_2426,N_2019);
or U2534 (N_2534,N_2198,N_2483);
nand U2535 (N_2535,N_2263,N_2270);
and U2536 (N_2536,N_2007,N_2009);
and U2537 (N_2537,N_2060,N_2447);
nor U2538 (N_2538,N_2069,N_2020);
and U2539 (N_2539,N_2276,N_2185);
nand U2540 (N_2540,N_2119,N_2145);
nor U2541 (N_2541,N_2281,N_2015);
nand U2542 (N_2542,N_2433,N_2173);
xnor U2543 (N_2543,N_2166,N_2287);
nand U2544 (N_2544,N_2039,N_2386);
nor U2545 (N_2545,N_2102,N_2109);
or U2546 (N_2546,N_2211,N_2098);
xnor U2547 (N_2547,N_2062,N_2429);
nor U2548 (N_2548,N_2257,N_2362);
or U2549 (N_2549,N_2014,N_2018);
and U2550 (N_2550,N_2216,N_2279);
and U2551 (N_2551,N_2025,N_2304);
nand U2552 (N_2552,N_2205,N_2187);
and U2553 (N_2553,N_2394,N_2456);
or U2554 (N_2554,N_2095,N_2144);
and U2555 (N_2555,N_2298,N_2315);
and U2556 (N_2556,N_2163,N_2268);
and U2557 (N_2557,N_2252,N_2143);
or U2558 (N_2558,N_2115,N_2051);
nand U2559 (N_2559,N_2357,N_2053);
nand U2560 (N_2560,N_2127,N_2280);
or U2561 (N_2561,N_2135,N_2488);
nor U2562 (N_2562,N_2234,N_2099);
and U2563 (N_2563,N_2484,N_2003);
nor U2564 (N_2564,N_2006,N_2254);
xor U2565 (N_2565,N_2023,N_2385);
nand U2566 (N_2566,N_2113,N_2289);
nor U2567 (N_2567,N_2203,N_2367);
xor U2568 (N_2568,N_2118,N_2082);
xnor U2569 (N_2569,N_2435,N_2207);
xor U2570 (N_2570,N_2277,N_2474);
nand U2571 (N_2571,N_2492,N_2238);
or U2572 (N_2572,N_2017,N_2253);
nand U2573 (N_2573,N_2142,N_2050);
or U2574 (N_2574,N_2273,N_2181);
nand U2575 (N_2575,N_2220,N_2395);
nand U2576 (N_2576,N_2455,N_2125);
or U2577 (N_2577,N_2191,N_2403);
nand U2578 (N_2578,N_2215,N_2467);
nor U2579 (N_2579,N_2258,N_2381);
or U2580 (N_2580,N_2179,N_2073);
nand U2581 (N_2581,N_2213,N_2415);
or U2582 (N_2582,N_2209,N_2333);
or U2583 (N_2583,N_2089,N_2461);
or U2584 (N_2584,N_2172,N_2317);
or U2585 (N_2585,N_2493,N_2134);
nor U2586 (N_2586,N_2180,N_2244);
or U2587 (N_2587,N_2407,N_2075);
or U2588 (N_2588,N_2214,N_2221);
nand U2589 (N_2589,N_2419,N_2128);
or U2590 (N_2590,N_2152,N_2405);
nor U2591 (N_2591,N_2323,N_2340);
nand U2592 (N_2592,N_2208,N_2459);
xor U2593 (N_2593,N_2248,N_2265);
or U2594 (N_2594,N_2071,N_2054);
nand U2595 (N_2595,N_2196,N_2138);
nand U2596 (N_2596,N_2491,N_2372);
and U2597 (N_2597,N_2383,N_2189);
nor U2598 (N_2598,N_2322,N_2370);
xor U2599 (N_2599,N_2174,N_2024);
and U2600 (N_2600,N_2212,N_2305);
nand U2601 (N_2601,N_2168,N_2463);
nand U2602 (N_2602,N_2005,N_2081);
or U2603 (N_2603,N_2267,N_2348);
xnor U2604 (N_2604,N_2249,N_2401);
or U2605 (N_2605,N_2409,N_2197);
and U2606 (N_2606,N_2165,N_2162);
and U2607 (N_2607,N_2091,N_2392);
xnor U2608 (N_2608,N_2160,N_2184);
xnor U2609 (N_2609,N_2496,N_2049);
nor U2610 (N_2610,N_2176,N_2497);
xnor U2611 (N_2611,N_2294,N_2041);
xor U2612 (N_2612,N_2318,N_2247);
or U2613 (N_2613,N_2044,N_2094);
nor U2614 (N_2614,N_2195,N_2122);
or U2615 (N_2615,N_2465,N_2454);
nand U2616 (N_2616,N_2453,N_2058);
nor U2617 (N_2617,N_2255,N_2349);
nand U2618 (N_2618,N_2130,N_2421);
or U2619 (N_2619,N_2424,N_2078);
xor U2620 (N_2620,N_2031,N_2106);
xnor U2621 (N_2621,N_2107,N_2087);
and U2622 (N_2622,N_2296,N_2034);
and U2623 (N_2623,N_2451,N_2111);
or U2624 (N_2624,N_2164,N_2241);
nor U2625 (N_2625,N_2004,N_2324);
xnor U2626 (N_2626,N_2412,N_2226);
or U2627 (N_2627,N_2356,N_2011);
nand U2628 (N_2628,N_2337,N_2411);
nand U2629 (N_2629,N_2408,N_2057);
nor U2630 (N_2630,N_2449,N_2271);
nor U2631 (N_2631,N_2103,N_2473);
and U2632 (N_2632,N_2359,N_2001);
and U2633 (N_2633,N_2422,N_2070);
xnor U2634 (N_2634,N_2159,N_2101);
xor U2635 (N_2635,N_2476,N_2350);
nor U2636 (N_2636,N_2033,N_2300);
nor U2637 (N_2637,N_2311,N_2085);
nor U2638 (N_2638,N_2443,N_2021);
or U2639 (N_2639,N_2132,N_2027);
xor U2640 (N_2640,N_2190,N_2028);
and U2641 (N_2641,N_2288,N_2201);
or U2642 (N_2642,N_2157,N_2260);
xnor U2643 (N_2643,N_2448,N_2387);
nand U2644 (N_2644,N_2074,N_2345);
nor U2645 (N_2645,N_2139,N_2470);
xnor U2646 (N_2646,N_2240,N_2256);
nor U2647 (N_2647,N_2266,N_2338);
nor U2648 (N_2648,N_2462,N_2148);
xor U2649 (N_2649,N_2396,N_2436);
or U2650 (N_2650,N_2010,N_2232);
nor U2651 (N_2651,N_2375,N_2056);
nand U2652 (N_2652,N_2479,N_2038);
and U2653 (N_2653,N_2245,N_2108);
nor U2654 (N_2654,N_2498,N_2339);
or U2655 (N_2655,N_2242,N_2175);
or U2656 (N_2656,N_2413,N_2035);
xnor U2657 (N_2657,N_2458,N_2321);
and U2658 (N_2658,N_2499,N_2332);
nor U2659 (N_2659,N_2437,N_2380);
nor U2660 (N_2660,N_2307,N_2026);
nand U2661 (N_2661,N_2334,N_2140);
nand U2662 (N_2662,N_2314,N_2194);
nor U2663 (N_2663,N_2328,N_2365);
xor U2664 (N_2664,N_2114,N_2066);
nand U2665 (N_2665,N_2188,N_2354);
or U2666 (N_2666,N_2022,N_2278);
xnor U2667 (N_2667,N_2371,N_2222);
xnor U2668 (N_2668,N_2495,N_2126);
xnor U2669 (N_2669,N_2210,N_2431);
or U2670 (N_2670,N_2442,N_2430);
and U2671 (N_2671,N_2086,N_2351);
and U2672 (N_2672,N_2331,N_2480);
nor U2673 (N_2673,N_2303,N_2097);
or U2674 (N_2674,N_2065,N_2192);
xnor U2675 (N_2675,N_2090,N_2344);
or U2676 (N_2676,N_2477,N_2150);
nand U2677 (N_2677,N_2327,N_2306);
nor U2678 (N_2678,N_2110,N_2170);
nand U2679 (N_2679,N_2445,N_2224);
nor U2680 (N_2680,N_2379,N_2384);
nand U2681 (N_2681,N_2264,N_2167);
or U2682 (N_2682,N_2117,N_2048);
xnor U2683 (N_2683,N_2466,N_2046);
or U2684 (N_2684,N_2377,N_2487);
and U2685 (N_2685,N_2153,N_2225);
nand U2686 (N_2686,N_2472,N_2376);
and U2687 (N_2687,N_2121,N_2229);
nand U2688 (N_2688,N_2223,N_2283);
and U2689 (N_2689,N_2423,N_2228);
xnor U2690 (N_2690,N_2068,N_2388);
or U2691 (N_2691,N_2030,N_2055);
nor U2692 (N_2692,N_2088,N_2012);
nor U2693 (N_2693,N_2149,N_2293);
and U2694 (N_2694,N_2131,N_2335);
xor U2695 (N_2695,N_2427,N_2490);
nor U2696 (N_2696,N_2404,N_2274);
xnor U2697 (N_2697,N_2374,N_2400);
or U2698 (N_2698,N_2460,N_2416);
xnor U2699 (N_2699,N_2308,N_2382);
nand U2700 (N_2700,N_2151,N_2446);
xor U2701 (N_2701,N_2471,N_2439);
xnor U2702 (N_2702,N_2341,N_2169);
nor U2703 (N_2703,N_2231,N_2052);
nand U2704 (N_2704,N_2199,N_2353);
or U2705 (N_2705,N_2147,N_2029);
or U2706 (N_2706,N_2373,N_2269);
xor U2707 (N_2707,N_2177,N_2156);
nand U2708 (N_2708,N_2398,N_2469);
nor U2709 (N_2709,N_2186,N_2227);
or U2710 (N_2710,N_2355,N_2363);
and U2711 (N_2711,N_2161,N_2389);
nor U2712 (N_2712,N_2282,N_2243);
or U2713 (N_2713,N_2285,N_2313);
nand U2714 (N_2714,N_2123,N_2112);
nand U2715 (N_2715,N_2406,N_2478);
nor U2716 (N_2716,N_2059,N_2302);
or U2717 (N_2717,N_2043,N_2218);
xnor U2718 (N_2718,N_2414,N_2141);
or U2719 (N_2719,N_2358,N_2158);
xor U2720 (N_2720,N_2246,N_2155);
and U2721 (N_2721,N_2325,N_2077);
xor U2722 (N_2722,N_2364,N_2237);
nand U2723 (N_2723,N_2486,N_2045);
and U2724 (N_2724,N_2104,N_2182);
and U2725 (N_2725,N_2272,N_2286);
and U2726 (N_2726,N_2154,N_2390);
and U2727 (N_2727,N_2369,N_2076);
or U2728 (N_2728,N_2100,N_2347);
and U2729 (N_2729,N_2236,N_2330);
xnor U2730 (N_2730,N_2032,N_2320);
or U2731 (N_2731,N_2336,N_2425);
or U2732 (N_2732,N_2420,N_2489);
xor U2733 (N_2733,N_2064,N_2136);
xnor U2734 (N_2734,N_2262,N_2129);
xnor U2735 (N_2735,N_2002,N_2399);
and U2736 (N_2736,N_2343,N_2016);
xor U2737 (N_2737,N_2361,N_2219);
nand U2738 (N_2738,N_2402,N_2239);
nor U2739 (N_2739,N_2301,N_2468);
and U2740 (N_2740,N_2444,N_2072);
xnor U2741 (N_2741,N_2133,N_2000);
nand U2742 (N_2742,N_2290,N_2494);
nor U2743 (N_2743,N_2096,N_2368);
and U2744 (N_2744,N_2040,N_2193);
xor U2745 (N_2745,N_2410,N_2312);
or U2746 (N_2746,N_2063,N_2047);
nand U2747 (N_2747,N_2259,N_2230);
and U2748 (N_2748,N_2116,N_2120);
nand U2749 (N_2749,N_2146,N_2217);
xnor U2750 (N_2750,N_2099,N_2251);
xor U2751 (N_2751,N_2480,N_2192);
or U2752 (N_2752,N_2457,N_2167);
nor U2753 (N_2753,N_2464,N_2036);
and U2754 (N_2754,N_2028,N_2295);
or U2755 (N_2755,N_2093,N_2234);
nand U2756 (N_2756,N_2355,N_2001);
and U2757 (N_2757,N_2264,N_2078);
or U2758 (N_2758,N_2223,N_2113);
xnor U2759 (N_2759,N_2481,N_2271);
and U2760 (N_2760,N_2281,N_2419);
and U2761 (N_2761,N_2315,N_2167);
or U2762 (N_2762,N_2023,N_2465);
nor U2763 (N_2763,N_2208,N_2079);
nor U2764 (N_2764,N_2488,N_2038);
nor U2765 (N_2765,N_2220,N_2346);
xor U2766 (N_2766,N_2018,N_2336);
nand U2767 (N_2767,N_2034,N_2316);
xnor U2768 (N_2768,N_2307,N_2244);
or U2769 (N_2769,N_2136,N_2334);
or U2770 (N_2770,N_2278,N_2074);
nand U2771 (N_2771,N_2131,N_2353);
and U2772 (N_2772,N_2446,N_2118);
nor U2773 (N_2773,N_2286,N_2355);
nor U2774 (N_2774,N_2446,N_2341);
and U2775 (N_2775,N_2410,N_2229);
or U2776 (N_2776,N_2393,N_2010);
or U2777 (N_2777,N_2474,N_2275);
nand U2778 (N_2778,N_2007,N_2494);
and U2779 (N_2779,N_2110,N_2260);
and U2780 (N_2780,N_2188,N_2357);
and U2781 (N_2781,N_2472,N_2120);
or U2782 (N_2782,N_2398,N_2053);
xnor U2783 (N_2783,N_2461,N_2442);
xnor U2784 (N_2784,N_2350,N_2263);
xor U2785 (N_2785,N_2005,N_2375);
nand U2786 (N_2786,N_2402,N_2015);
xor U2787 (N_2787,N_2298,N_2409);
nand U2788 (N_2788,N_2105,N_2217);
or U2789 (N_2789,N_2308,N_2469);
nand U2790 (N_2790,N_2275,N_2073);
and U2791 (N_2791,N_2207,N_2163);
nor U2792 (N_2792,N_2002,N_2203);
nand U2793 (N_2793,N_2438,N_2302);
nor U2794 (N_2794,N_2162,N_2292);
or U2795 (N_2795,N_2362,N_2119);
nand U2796 (N_2796,N_2256,N_2058);
nor U2797 (N_2797,N_2410,N_2428);
and U2798 (N_2798,N_2090,N_2302);
or U2799 (N_2799,N_2374,N_2240);
xnor U2800 (N_2800,N_2055,N_2299);
or U2801 (N_2801,N_2114,N_2005);
and U2802 (N_2802,N_2379,N_2274);
and U2803 (N_2803,N_2058,N_2098);
xor U2804 (N_2804,N_2344,N_2485);
or U2805 (N_2805,N_2345,N_2292);
nand U2806 (N_2806,N_2065,N_2311);
and U2807 (N_2807,N_2137,N_2139);
or U2808 (N_2808,N_2358,N_2230);
nand U2809 (N_2809,N_2487,N_2457);
nor U2810 (N_2810,N_2470,N_2280);
and U2811 (N_2811,N_2102,N_2266);
or U2812 (N_2812,N_2326,N_2136);
or U2813 (N_2813,N_2147,N_2416);
nor U2814 (N_2814,N_2284,N_2352);
or U2815 (N_2815,N_2090,N_2176);
and U2816 (N_2816,N_2022,N_2029);
xnor U2817 (N_2817,N_2443,N_2154);
or U2818 (N_2818,N_2228,N_2246);
nand U2819 (N_2819,N_2264,N_2258);
or U2820 (N_2820,N_2411,N_2210);
and U2821 (N_2821,N_2227,N_2018);
xor U2822 (N_2822,N_2224,N_2319);
nor U2823 (N_2823,N_2062,N_2186);
nor U2824 (N_2824,N_2267,N_2357);
nand U2825 (N_2825,N_2398,N_2158);
nand U2826 (N_2826,N_2169,N_2011);
xnor U2827 (N_2827,N_2060,N_2145);
nor U2828 (N_2828,N_2063,N_2241);
or U2829 (N_2829,N_2333,N_2027);
xnor U2830 (N_2830,N_2213,N_2461);
xor U2831 (N_2831,N_2112,N_2339);
nor U2832 (N_2832,N_2001,N_2168);
nand U2833 (N_2833,N_2034,N_2491);
or U2834 (N_2834,N_2041,N_2028);
or U2835 (N_2835,N_2005,N_2463);
and U2836 (N_2836,N_2336,N_2335);
or U2837 (N_2837,N_2029,N_2491);
xor U2838 (N_2838,N_2098,N_2441);
nand U2839 (N_2839,N_2143,N_2052);
nand U2840 (N_2840,N_2499,N_2139);
and U2841 (N_2841,N_2474,N_2443);
nor U2842 (N_2842,N_2366,N_2274);
nand U2843 (N_2843,N_2140,N_2455);
xor U2844 (N_2844,N_2045,N_2099);
or U2845 (N_2845,N_2182,N_2417);
nand U2846 (N_2846,N_2063,N_2078);
nand U2847 (N_2847,N_2091,N_2288);
nor U2848 (N_2848,N_2458,N_2243);
and U2849 (N_2849,N_2114,N_2486);
nor U2850 (N_2850,N_2267,N_2497);
or U2851 (N_2851,N_2130,N_2242);
xnor U2852 (N_2852,N_2425,N_2254);
nor U2853 (N_2853,N_2033,N_2403);
xnor U2854 (N_2854,N_2319,N_2041);
nand U2855 (N_2855,N_2079,N_2490);
nand U2856 (N_2856,N_2410,N_2329);
nor U2857 (N_2857,N_2262,N_2423);
nand U2858 (N_2858,N_2355,N_2013);
xor U2859 (N_2859,N_2141,N_2241);
nor U2860 (N_2860,N_2181,N_2199);
nand U2861 (N_2861,N_2396,N_2431);
and U2862 (N_2862,N_2232,N_2326);
or U2863 (N_2863,N_2185,N_2493);
nand U2864 (N_2864,N_2127,N_2423);
and U2865 (N_2865,N_2460,N_2024);
and U2866 (N_2866,N_2479,N_2432);
xnor U2867 (N_2867,N_2348,N_2172);
nand U2868 (N_2868,N_2317,N_2055);
nor U2869 (N_2869,N_2418,N_2421);
and U2870 (N_2870,N_2308,N_2440);
and U2871 (N_2871,N_2145,N_2257);
nand U2872 (N_2872,N_2250,N_2024);
or U2873 (N_2873,N_2433,N_2343);
nand U2874 (N_2874,N_2439,N_2138);
nand U2875 (N_2875,N_2166,N_2080);
nor U2876 (N_2876,N_2361,N_2316);
nand U2877 (N_2877,N_2246,N_2166);
xnor U2878 (N_2878,N_2204,N_2390);
or U2879 (N_2879,N_2093,N_2022);
or U2880 (N_2880,N_2251,N_2178);
nor U2881 (N_2881,N_2011,N_2413);
and U2882 (N_2882,N_2475,N_2040);
or U2883 (N_2883,N_2047,N_2012);
and U2884 (N_2884,N_2426,N_2468);
xor U2885 (N_2885,N_2356,N_2103);
nor U2886 (N_2886,N_2443,N_2481);
nor U2887 (N_2887,N_2194,N_2262);
and U2888 (N_2888,N_2406,N_2018);
nor U2889 (N_2889,N_2324,N_2215);
and U2890 (N_2890,N_2079,N_2341);
or U2891 (N_2891,N_2474,N_2463);
and U2892 (N_2892,N_2039,N_2014);
and U2893 (N_2893,N_2306,N_2278);
xnor U2894 (N_2894,N_2094,N_2127);
or U2895 (N_2895,N_2038,N_2105);
and U2896 (N_2896,N_2051,N_2314);
or U2897 (N_2897,N_2110,N_2348);
nor U2898 (N_2898,N_2145,N_2307);
nand U2899 (N_2899,N_2383,N_2430);
nand U2900 (N_2900,N_2456,N_2345);
or U2901 (N_2901,N_2238,N_2097);
nor U2902 (N_2902,N_2173,N_2440);
or U2903 (N_2903,N_2174,N_2198);
xnor U2904 (N_2904,N_2324,N_2182);
nor U2905 (N_2905,N_2218,N_2051);
or U2906 (N_2906,N_2025,N_2493);
xor U2907 (N_2907,N_2121,N_2055);
xor U2908 (N_2908,N_2406,N_2186);
nor U2909 (N_2909,N_2102,N_2422);
nand U2910 (N_2910,N_2239,N_2000);
nor U2911 (N_2911,N_2435,N_2464);
or U2912 (N_2912,N_2300,N_2215);
xnor U2913 (N_2913,N_2263,N_2174);
nor U2914 (N_2914,N_2301,N_2064);
and U2915 (N_2915,N_2299,N_2084);
and U2916 (N_2916,N_2383,N_2186);
nand U2917 (N_2917,N_2169,N_2474);
xor U2918 (N_2918,N_2052,N_2191);
nor U2919 (N_2919,N_2150,N_2487);
nor U2920 (N_2920,N_2219,N_2067);
or U2921 (N_2921,N_2044,N_2059);
nor U2922 (N_2922,N_2212,N_2136);
or U2923 (N_2923,N_2049,N_2075);
and U2924 (N_2924,N_2357,N_2324);
or U2925 (N_2925,N_2033,N_2484);
or U2926 (N_2926,N_2193,N_2152);
and U2927 (N_2927,N_2220,N_2443);
xor U2928 (N_2928,N_2373,N_2265);
and U2929 (N_2929,N_2001,N_2271);
or U2930 (N_2930,N_2336,N_2465);
and U2931 (N_2931,N_2451,N_2262);
xor U2932 (N_2932,N_2071,N_2277);
nor U2933 (N_2933,N_2092,N_2224);
nand U2934 (N_2934,N_2305,N_2125);
or U2935 (N_2935,N_2114,N_2350);
and U2936 (N_2936,N_2159,N_2071);
and U2937 (N_2937,N_2076,N_2444);
xor U2938 (N_2938,N_2386,N_2123);
xnor U2939 (N_2939,N_2248,N_2409);
nor U2940 (N_2940,N_2119,N_2441);
nand U2941 (N_2941,N_2254,N_2226);
and U2942 (N_2942,N_2323,N_2143);
or U2943 (N_2943,N_2387,N_2201);
nand U2944 (N_2944,N_2288,N_2435);
or U2945 (N_2945,N_2395,N_2267);
nor U2946 (N_2946,N_2137,N_2322);
nor U2947 (N_2947,N_2353,N_2476);
xnor U2948 (N_2948,N_2290,N_2435);
or U2949 (N_2949,N_2399,N_2232);
nor U2950 (N_2950,N_2290,N_2233);
or U2951 (N_2951,N_2026,N_2066);
nand U2952 (N_2952,N_2259,N_2059);
and U2953 (N_2953,N_2202,N_2499);
xnor U2954 (N_2954,N_2352,N_2019);
xnor U2955 (N_2955,N_2480,N_2362);
and U2956 (N_2956,N_2193,N_2229);
nand U2957 (N_2957,N_2189,N_2059);
nor U2958 (N_2958,N_2344,N_2169);
or U2959 (N_2959,N_2099,N_2479);
and U2960 (N_2960,N_2329,N_2203);
nor U2961 (N_2961,N_2010,N_2008);
or U2962 (N_2962,N_2318,N_2453);
or U2963 (N_2963,N_2425,N_2123);
nor U2964 (N_2964,N_2370,N_2085);
and U2965 (N_2965,N_2131,N_2068);
nor U2966 (N_2966,N_2327,N_2359);
nor U2967 (N_2967,N_2208,N_2222);
nor U2968 (N_2968,N_2331,N_2256);
nand U2969 (N_2969,N_2485,N_2315);
or U2970 (N_2970,N_2363,N_2144);
xor U2971 (N_2971,N_2130,N_2399);
xnor U2972 (N_2972,N_2046,N_2442);
nor U2973 (N_2973,N_2243,N_2264);
xor U2974 (N_2974,N_2192,N_2254);
or U2975 (N_2975,N_2236,N_2032);
nor U2976 (N_2976,N_2038,N_2433);
nor U2977 (N_2977,N_2351,N_2325);
nor U2978 (N_2978,N_2408,N_2264);
and U2979 (N_2979,N_2165,N_2004);
nor U2980 (N_2980,N_2361,N_2265);
nand U2981 (N_2981,N_2390,N_2355);
and U2982 (N_2982,N_2096,N_2151);
and U2983 (N_2983,N_2112,N_2488);
nand U2984 (N_2984,N_2005,N_2285);
and U2985 (N_2985,N_2274,N_2192);
nand U2986 (N_2986,N_2023,N_2321);
nand U2987 (N_2987,N_2173,N_2225);
and U2988 (N_2988,N_2158,N_2021);
nand U2989 (N_2989,N_2072,N_2044);
nand U2990 (N_2990,N_2407,N_2328);
nand U2991 (N_2991,N_2013,N_2196);
and U2992 (N_2992,N_2223,N_2426);
and U2993 (N_2993,N_2282,N_2087);
and U2994 (N_2994,N_2253,N_2144);
nand U2995 (N_2995,N_2263,N_2427);
and U2996 (N_2996,N_2019,N_2134);
nand U2997 (N_2997,N_2391,N_2334);
nand U2998 (N_2998,N_2017,N_2099);
or U2999 (N_2999,N_2202,N_2335);
xnor U3000 (N_3000,N_2724,N_2823);
xor U3001 (N_3001,N_2749,N_2584);
nor U3002 (N_3002,N_2733,N_2643);
and U3003 (N_3003,N_2654,N_2664);
or U3004 (N_3004,N_2856,N_2544);
and U3005 (N_3005,N_2891,N_2660);
or U3006 (N_3006,N_2800,N_2904);
xor U3007 (N_3007,N_2626,N_2814);
xnor U3008 (N_3008,N_2854,N_2922);
and U3009 (N_3009,N_2882,N_2524);
nand U3010 (N_3010,N_2534,N_2825);
or U3011 (N_3011,N_2914,N_2907);
nor U3012 (N_3012,N_2738,N_2833);
nor U3013 (N_3013,N_2564,N_2616);
or U3014 (N_3014,N_2992,N_2821);
or U3015 (N_3015,N_2936,N_2890);
nor U3016 (N_3016,N_2717,N_2950);
nor U3017 (N_3017,N_2745,N_2578);
nand U3018 (N_3018,N_2901,N_2592);
xnor U3019 (N_3019,N_2542,N_2507);
nor U3020 (N_3020,N_2655,N_2576);
xor U3021 (N_3021,N_2743,N_2892);
and U3022 (N_3022,N_2978,N_2646);
or U3023 (N_3023,N_2969,N_2644);
nand U3024 (N_3024,N_2678,N_2887);
nand U3025 (N_3025,N_2596,N_2767);
or U3026 (N_3026,N_2740,N_2828);
nand U3027 (N_3027,N_2668,N_2897);
and U3028 (N_3028,N_2750,N_2820);
or U3029 (N_3029,N_2605,N_2555);
and U3030 (N_3030,N_2774,N_2709);
nand U3031 (N_3031,N_2903,N_2554);
xor U3032 (N_3032,N_2710,N_2567);
and U3033 (N_3033,N_2725,N_2672);
xor U3034 (N_3034,N_2667,N_2770);
xnor U3035 (N_3035,N_2959,N_2504);
xor U3036 (N_3036,N_2998,N_2874);
or U3037 (N_3037,N_2719,N_2894);
nand U3038 (N_3038,N_2631,N_2527);
nand U3039 (N_3039,N_2520,N_2515);
nor U3040 (N_3040,N_2824,N_2840);
and U3041 (N_3041,N_2819,N_2784);
or U3042 (N_3042,N_2863,N_2620);
nor U3043 (N_3043,N_2853,N_2679);
and U3044 (N_3044,N_2871,N_2707);
nand U3045 (N_3045,N_2810,N_2662);
and U3046 (N_3046,N_2666,N_2744);
and U3047 (N_3047,N_2610,N_2532);
nand U3048 (N_3048,N_2635,N_2798);
nor U3049 (N_3049,N_2921,N_2625);
nand U3050 (N_3050,N_2940,N_2975);
and U3051 (N_3051,N_2613,N_2817);
xnor U3052 (N_3052,N_2811,N_2851);
and U3053 (N_3053,N_2797,N_2756);
xor U3054 (N_3054,N_2609,N_2618);
or U3055 (N_3055,N_2972,N_2946);
nor U3056 (N_3056,N_2640,N_2989);
xor U3057 (N_3057,N_2802,N_2873);
or U3058 (N_3058,N_2875,N_2686);
nor U3059 (N_3059,N_2933,N_2697);
nor U3060 (N_3060,N_2553,N_2729);
or U3061 (N_3061,N_2706,N_2572);
xor U3062 (N_3062,N_2685,N_2731);
nand U3063 (N_3063,N_2547,N_2715);
nand U3064 (N_3064,N_2557,N_2966);
and U3065 (N_3065,N_2805,N_2781);
nand U3066 (N_3066,N_2562,N_2792);
or U3067 (N_3067,N_2769,N_2732);
xor U3068 (N_3068,N_2742,N_2790);
nor U3069 (N_3069,N_2812,N_2513);
nor U3070 (N_3070,N_2793,N_2832);
nand U3071 (N_3071,N_2846,N_2638);
and U3072 (N_3072,N_2628,N_2949);
nor U3073 (N_3073,N_2560,N_2876);
or U3074 (N_3074,N_2748,N_2773);
nor U3075 (N_3075,N_2964,N_2671);
and U3076 (N_3076,N_2632,N_2735);
and U3077 (N_3077,N_2939,N_2923);
or U3078 (N_3078,N_2859,N_2841);
nor U3079 (N_3079,N_2830,N_2885);
and U3080 (N_3080,N_2981,N_2508);
xnor U3081 (N_3081,N_2565,N_2925);
nand U3082 (N_3082,N_2838,N_2545);
or U3083 (N_3083,N_2988,N_2886);
or U3084 (N_3084,N_2764,N_2794);
and U3085 (N_3085,N_2834,N_2653);
and U3086 (N_3086,N_2768,N_2866);
xor U3087 (N_3087,N_2888,N_2583);
nor U3088 (N_3088,N_2980,N_2751);
xnor U3089 (N_3089,N_2573,N_2642);
and U3090 (N_3090,N_2860,N_2996);
nand U3091 (N_3091,N_2566,N_2525);
xor U3092 (N_3092,N_2763,N_2928);
and U3093 (N_3093,N_2899,N_2523);
or U3094 (N_3094,N_2561,N_2574);
and U3095 (N_3095,N_2734,N_2870);
nor U3096 (N_3096,N_2747,N_2912);
and U3097 (N_3097,N_2995,N_2737);
nand U3098 (N_3098,N_2765,N_2977);
and U3099 (N_3099,N_2600,N_2550);
or U3100 (N_3100,N_2500,N_2771);
and U3101 (N_3101,N_2815,N_2836);
nand U3102 (N_3102,N_2597,N_2906);
xor U3103 (N_3103,N_2880,N_2657);
or U3104 (N_3104,N_2934,N_2868);
xor U3105 (N_3105,N_2736,N_2700);
and U3106 (N_3106,N_2987,N_2589);
and U3107 (N_3107,N_2968,N_2982);
xor U3108 (N_3108,N_2505,N_2692);
nand U3109 (N_3109,N_2570,N_2693);
and U3110 (N_3110,N_2760,N_2663);
and U3111 (N_3111,N_2918,N_2986);
xor U3112 (N_3112,N_2630,N_2952);
nor U3113 (N_3113,N_2639,N_2852);
or U3114 (N_3114,N_2571,N_2758);
xnor U3115 (N_3115,N_2687,N_2675);
xnor U3116 (N_3116,N_2967,N_2543);
and U3117 (N_3117,N_2935,N_2761);
nand U3118 (N_3118,N_2510,N_2955);
nor U3119 (N_3119,N_2577,N_2911);
or U3120 (N_3120,N_2984,N_2612);
xor U3121 (N_3121,N_2953,N_2783);
xnor U3122 (N_3122,N_2712,N_2549);
and U3123 (N_3123,N_2593,N_2924);
or U3124 (N_3124,N_2927,N_2929);
nor U3125 (N_3125,N_2985,N_2705);
nor U3126 (N_3126,N_2855,N_2938);
or U3127 (N_3127,N_2777,N_2575);
nor U3128 (N_3128,N_2536,N_2806);
xnor U3129 (N_3129,N_2976,N_2591);
or U3130 (N_3130,N_2603,N_2858);
or U3131 (N_3131,N_2594,N_2512);
nor U3132 (N_3132,N_2658,N_2961);
nand U3133 (N_3133,N_2633,N_2822);
and U3134 (N_3134,N_2842,N_2845);
and U3135 (N_3135,N_2599,N_2530);
or U3136 (N_3136,N_2910,N_2533);
or U3137 (N_3137,N_2881,N_2909);
or U3138 (N_3138,N_2844,N_2869);
and U3139 (N_3139,N_2619,N_2990);
nand U3140 (N_3140,N_2791,N_2682);
xnor U3141 (N_3141,N_2943,N_2716);
and U3142 (N_3142,N_2711,N_2651);
nor U3143 (N_3143,N_2701,N_2908);
nor U3144 (N_3144,N_2623,N_2615);
and U3145 (N_3145,N_2579,N_2741);
xnor U3146 (N_3146,N_2611,N_2691);
nor U3147 (N_3147,N_2641,N_2535);
nor U3148 (N_3148,N_2690,N_2727);
and U3149 (N_3149,N_2538,N_2546);
nand U3150 (N_3150,N_2649,N_2837);
or U3151 (N_3151,N_2721,N_2926);
and U3152 (N_3152,N_2608,N_2867);
xnor U3153 (N_3153,N_2816,N_2884);
nor U3154 (N_3154,N_2826,N_2702);
xnor U3155 (N_3155,N_2720,N_2598);
nand U3156 (N_3156,N_2522,N_2636);
and U3157 (N_3157,N_2829,N_2541);
or U3158 (N_3158,N_2941,N_2669);
nor U3159 (N_3159,N_2606,N_2796);
xnor U3160 (N_3160,N_2993,N_2896);
xor U3161 (N_3161,N_2835,N_2958);
nand U3162 (N_3162,N_2857,N_2942);
nand U3163 (N_3163,N_2537,N_2580);
nor U3164 (N_3164,N_2723,N_2762);
nor U3165 (N_3165,N_2779,N_2915);
nor U3166 (N_3166,N_2970,N_2746);
and U3167 (N_3167,N_2947,N_2694);
and U3168 (N_3168,N_2991,N_2695);
nand U3169 (N_3169,N_2799,N_2994);
or U3170 (N_3170,N_2703,N_2813);
nand U3171 (N_3171,N_2889,N_2514);
and U3172 (N_3172,N_2607,N_2772);
xor U3173 (N_3173,N_2698,N_2604);
xor U3174 (N_3174,N_2752,N_2917);
nor U3175 (N_3175,N_2913,N_2704);
nand U3176 (N_3176,N_2503,N_2808);
or U3177 (N_3177,N_2883,N_2877);
and U3178 (N_3178,N_2521,N_2932);
nor U3179 (N_3179,N_2900,N_2518);
nand U3180 (N_3180,N_2965,N_2588);
and U3181 (N_3181,N_2937,N_2590);
nor U3182 (N_3182,N_2722,N_2581);
nand U3183 (N_3183,N_2905,N_2502);
nand U3184 (N_3184,N_2595,N_2809);
and U3185 (N_3185,N_2587,N_2782);
and U3186 (N_3186,N_2531,N_2753);
nor U3187 (N_3187,N_2755,N_2728);
nand U3188 (N_3188,N_2879,N_2872);
nor U3189 (N_3189,N_2552,N_2568);
xor U3190 (N_3190,N_2960,N_2979);
and U3191 (N_3191,N_2634,N_2569);
and U3192 (N_3192,N_2637,N_2775);
xnor U3193 (N_3193,N_2848,N_2999);
nor U3194 (N_3194,N_2766,N_2676);
or U3195 (N_3195,N_2674,N_2511);
xor U3196 (N_3196,N_2659,N_2818);
nor U3197 (N_3197,N_2843,N_2787);
nor U3198 (N_3198,N_2621,N_2516);
nor U3199 (N_3199,N_2931,N_2739);
or U3200 (N_3200,N_2661,N_2624);
xnor U3201 (N_3201,N_2714,N_2801);
xor U3202 (N_3202,N_2713,N_2974);
or U3203 (N_3203,N_2696,N_2789);
nand U3204 (N_3204,N_2627,N_2684);
nor U3205 (N_3205,N_2526,N_2517);
and U3206 (N_3206,N_2650,N_2726);
and U3207 (N_3207,N_2916,N_2898);
and U3208 (N_3208,N_2963,N_2670);
and U3209 (N_3209,N_2559,N_2944);
nand U3210 (N_3210,N_2602,N_2689);
and U3211 (N_3211,N_2582,N_2648);
xor U3212 (N_3212,N_2528,N_2788);
nor U3213 (N_3213,N_2708,N_2656);
or U3214 (N_3214,N_2930,N_2865);
nand U3215 (N_3215,N_2778,N_2501);
or U3216 (N_3216,N_2647,N_2850);
nor U3217 (N_3217,N_2807,N_2971);
nand U3218 (N_3218,N_2847,N_2548);
xor U3219 (N_3219,N_2839,N_2539);
and U3220 (N_3220,N_2601,N_2803);
and U3221 (N_3221,N_2919,N_2957);
xor U3222 (N_3222,N_2730,N_2786);
nor U3223 (N_3223,N_2540,N_2506);
xor U3224 (N_3224,N_2878,N_2785);
or U3225 (N_3225,N_2831,N_2893);
nor U3226 (N_3226,N_2680,N_2556);
and U3227 (N_3227,N_2757,N_2954);
xnor U3228 (N_3228,N_2629,N_2586);
and U3229 (N_3229,N_2519,N_2849);
nand U3230 (N_3230,N_2509,N_2945);
xor U3231 (N_3231,N_2983,N_2948);
nor U3232 (N_3232,N_2622,N_2614);
nand U3233 (N_3233,N_2645,N_2962);
and U3234 (N_3234,N_2804,N_2699);
and U3235 (N_3235,N_2997,N_2529);
xnor U3236 (N_3236,N_2652,N_2551);
nand U3237 (N_3237,N_2585,N_2718);
xnor U3238 (N_3238,N_2951,N_2754);
or U3239 (N_3239,N_2776,N_2617);
and U3240 (N_3240,N_2902,N_2795);
and U3241 (N_3241,N_2688,N_2827);
and U3242 (N_3242,N_2563,N_2683);
nand U3243 (N_3243,N_2956,N_2681);
xnor U3244 (N_3244,N_2673,N_2861);
xnor U3245 (N_3245,N_2862,N_2895);
nor U3246 (N_3246,N_2665,N_2973);
nor U3247 (N_3247,N_2864,N_2759);
xnor U3248 (N_3248,N_2920,N_2780);
or U3249 (N_3249,N_2677,N_2558);
nand U3250 (N_3250,N_2925,N_2926);
xor U3251 (N_3251,N_2888,N_2649);
xnor U3252 (N_3252,N_2579,N_2526);
xnor U3253 (N_3253,N_2853,N_2522);
or U3254 (N_3254,N_2747,N_2607);
xor U3255 (N_3255,N_2559,N_2685);
xnor U3256 (N_3256,N_2689,N_2956);
xor U3257 (N_3257,N_2746,N_2729);
or U3258 (N_3258,N_2670,N_2620);
or U3259 (N_3259,N_2993,N_2822);
or U3260 (N_3260,N_2897,N_2982);
nand U3261 (N_3261,N_2705,N_2557);
xor U3262 (N_3262,N_2597,N_2535);
nand U3263 (N_3263,N_2685,N_2666);
and U3264 (N_3264,N_2764,N_2663);
nor U3265 (N_3265,N_2837,N_2736);
nor U3266 (N_3266,N_2784,N_2660);
nor U3267 (N_3267,N_2541,N_2795);
or U3268 (N_3268,N_2772,N_2535);
nor U3269 (N_3269,N_2647,N_2771);
and U3270 (N_3270,N_2691,N_2612);
xnor U3271 (N_3271,N_2648,N_2821);
xor U3272 (N_3272,N_2513,N_2685);
and U3273 (N_3273,N_2793,N_2696);
or U3274 (N_3274,N_2813,N_2944);
nor U3275 (N_3275,N_2654,N_2665);
nand U3276 (N_3276,N_2529,N_2580);
and U3277 (N_3277,N_2949,N_2872);
nor U3278 (N_3278,N_2665,N_2965);
and U3279 (N_3279,N_2841,N_2777);
xnor U3280 (N_3280,N_2797,N_2953);
and U3281 (N_3281,N_2774,N_2561);
xnor U3282 (N_3282,N_2572,N_2700);
xor U3283 (N_3283,N_2912,N_2648);
xnor U3284 (N_3284,N_2742,N_2977);
or U3285 (N_3285,N_2512,N_2725);
or U3286 (N_3286,N_2569,N_2581);
and U3287 (N_3287,N_2942,N_2904);
or U3288 (N_3288,N_2879,N_2635);
nand U3289 (N_3289,N_2750,N_2579);
and U3290 (N_3290,N_2529,N_2900);
xor U3291 (N_3291,N_2566,N_2744);
and U3292 (N_3292,N_2778,N_2745);
or U3293 (N_3293,N_2577,N_2841);
xor U3294 (N_3294,N_2836,N_2930);
and U3295 (N_3295,N_2877,N_2577);
nand U3296 (N_3296,N_2692,N_2895);
nand U3297 (N_3297,N_2922,N_2600);
nor U3298 (N_3298,N_2831,N_2773);
or U3299 (N_3299,N_2861,N_2662);
and U3300 (N_3300,N_2951,N_2899);
nor U3301 (N_3301,N_2749,N_2941);
xnor U3302 (N_3302,N_2528,N_2607);
xnor U3303 (N_3303,N_2680,N_2725);
or U3304 (N_3304,N_2918,N_2868);
and U3305 (N_3305,N_2712,N_2938);
and U3306 (N_3306,N_2534,N_2956);
and U3307 (N_3307,N_2717,N_2886);
nand U3308 (N_3308,N_2957,N_2990);
nand U3309 (N_3309,N_2714,N_2834);
and U3310 (N_3310,N_2792,N_2754);
xnor U3311 (N_3311,N_2846,N_2865);
nand U3312 (N_3312,N_2770,N_2602);
nor U3313 (N_3313,N_2691,N_2542);
nand U3314 (N_3314,N_2551,N_2782);
nor U3315 (N_3315,N_2910,N_2833);
and U3316 (N_3316,N_2644,N_2961);
nand U3317 (N_3317,N_2807,N_2588);
or U3318 (N_3318,N_2627,N_2778);
nand U3319 (N_3319,N_2602,N_2523);
nand U3320 (N_3320,N_2973,N_2559);
nand U3321 (N_3321,N_2762,N_2593);
and U3322 (N_3322,N_2900,N_2506);
xnor U3323 (N_3323,N_2773,N_2971);
nand U3324 (N_3324,N_2641,N_2775);
nand U3325 (N_3325,N_2794,N_2950);
nor U3326 (N_3326,N_2994,N_2544);
or U3327 (N_3327,N_2986,N_2973);
or U3328 (N_3328,N_2667,N_2906);
nand U3329 (N_3329,N_2596,N_2735);
and U3330 (N_3330,N_2888,N_2678);
and U3331 (N_3331,N_2960,N_2746);
and U3332 (N_3332,N_2998,N_2706);
nand U3333 (N_3333,N_2767,N_2738);
xor U3334 (N_3334,N_2992,N_2823);
and U3335 (N_3335,N_2504,N_2675);
and U3336 (N_3336,N_2736,N_2719);
xnor U3337 (N_3337,N_2694,N_2965);
and U3338 (N_3338,N_2639,N_2666);
nor U3339 (N_3339,N_2812,N_2834);
or U3340 (N_3340,N_2617,N_2659);
xor U3341 (N_3341,N_2838,N_2548);
nand U3342 (N_3342,N_2625,N_2579);
nor U3343 (N_3343,N_2743,N_2548);
nand U3344 (N_3344,N_2785,N_2514);
or U3345 (N_3345,N_2921,N_2669);
nand U3346 (N_3346,N_2853,N_2953);
nand U3347 (N_3347,N_2980,N_2965);
or U3348 (N_3348,N_2684,N_2979);
nor U3349 (N_3349,N_2654,N_2803);
nand U3350 (N_3350,N_2849,N_2562);
xnor U3351 (N_3351,N_2909,N_2572);
nor U3352 (N_3352,N_2591,N_2894);
xor U3353 (N_3353,N_2782,N_2870);
or U3354 (N_3354,N_2791,N_2636);
and U3355 (N_3355,N_2609,N_2606);
or U3356 (N_3356,N_2650,N_2873);
and U3357 (N_3357,N_2688,N_2649);
nor U3358 (N_3358,N_2702,N_2547);
and U3359 (N_3359,N_2729,N_2533);
or U3360 (N_3360,N_2851,N_2688);
and U3361 (N_3361,N_2639,N_2956);
nand U3362 (N_3362,N_2700,N_2958);
nand U3363 (N_3363,N_2784,N_2697);
nand U3364 (N_3364,N_2959,N_2969);
nor U3365 (N_3365,N_2618,N_2837);
and U3366 (N_3366,N_2591,N_2983);
or U3367 (N_3367,N_2731,N_2859);
nand U3368 (N_3368,N_2764,N_2894);
or U3369 (N_3369,N_2709,N_2521);
xnor U3370 (N_3370,N_2772,N_2811);
and U3371 (N_3371,N_2552,N_2741);
or U3372 (N_3372,N_2577,N_2790);
nor U3373 (N_3373,N_2742,N_2796);
or U3374 (N_3374,N_2854,N_2825);
nor U3375 (N_3375,N_2677,N_2807);
and U3376 (N_3376,N_2602,N_2817);
nand U3377 (N_3377,N_2876,N_2984);
or U3378 (N_3378,N_2711,N_2959);
nor U3379 (N_3379,N_2689,N_2601);
or U3380 (N_3380,N_2582,N_2993);
or U3381 (N_3381,N_2540,N_2962);
nor U3382 (N_3382,N_2921,N_2676);
or U3383 (N_3383,N_2748,N_2844);
and U3384 (N_3384,N_2521,N_2792);
or U3385 (N_3385,N_2980,N_2526);
or U3386 (N_3386,N_2925,N_2500);
and U3387 (N_3387,N_2950,N_2914);
xor U3388 (N_3388,N_2742,N_2621);
xnor U3389 (N_3389,N_2871,N_2533);
xnor U3390 (N_3390,N_2582,N_2654);
nand U3391 (N_3391,N_2603,N_2882);
or U3392 (N_3392,N_2860,N_2596);
and U3393 (N_3393,N_2534,N_2529);
nor U3394 (N_3394,N_2825,N_2801);
nand U3395 (N_3395,N_2673,N_2999);
nand U3396 (N_3396,N_2973,N_2736);
nand U3397 (N_3397,N_2728,N_2782);
nand U3398 (N_3398,N_2946,N_2752);
nor U3399 (N_3399,N_2570,N_2975);
nor U3400 (N_3400,N_2940,N_2547);
and U3401 (N_3401,N_2871,N_2932);
xor U3402 (N_3402,N_2936,N_2546);
xnor U3403 (N_3403,N_2661,N_2513);
xnor U3404 (N_3404,N_2933,N_2675);
and U3405 (N_3405,N_2604,N_2753);
or U3406 (N_3406,N_2938,N_2768);
xor U3407 (N_3407,N_2627,N_2729);
or U3408 (N_3408,N_2556,N_2922);
or U3409 (N_3409,N_2536,N_2726);
xor U3410 (N_3410,N_2727,N_2598);
nor U3411 (N_3411,N_2624,N_2675);
nor U3412 (N_3412,N_2658,N_2786);
nand U3413 (N_3413,N_2896,N_2568);
nor U3414 (N_3414,N_2906,N_2729);
nand U3415 (N_3415,N_2969,N_2550);
or U3416 (N_3416,N_2904,N_2797);
and U3417 (N_3417,N_2601,N_2580);
nor U3418 (N_3418,N_2889,N_2966);
nor U3419 (N_3419,N_2565,N_2795);
nand U3420 (N_3420,N_2825,N_2996);
nor U3421 (N_3421,N_2505,N_2722);
and U3422 (N_3422,N_2853,N_2708);
and U3423 (N_3423,N_2573,N_2846);
nand U3424 (N_3424,N_2671,N_2854);
and U3425 (N_3425,N_2831,N_2723);
or U3426 (N_3426,N_2904,N_2994);
nor U3427 (N_3427,N_2734,N_2895);
or U3428 (N_3428,N_2737,N_2908);
and U3429 (N_3429,N_2734,N_2721);
nand U3430 (N_3430,N_2776,N_2771);
nand U3431 (N_3431,N_2771,N_2814);
nand U3432 (N_3432,N_2805,N_2760);
or U3433 (N_3433,N_2716,N_2737);
nand U3434 (N_3434,N_2680,N_2718);
and U3435 (N_3435,N_2600,N_2941);
nor U3436 (N_3436,N_2681,N_2701);
nor U3437 (N_3437,N_2711,N_2544);
or U3438 (N_3438,N_2971,N_2949);
and U3439 (N_3439,N_2681,N_2691);
or U3440 (N_3440,N_2832,N_2663);
xnor U3441 (N_3441,N_2849,N_2750);
xor U3442 (N_3442,N_2694,N_2831);
xor U3443 (N_3443,N_2608,N_2995);
and U3444 (N_3444,N_2765,N_2875);
nor U3445 (N_3445,N_2720,N_2561);
nand U3446 (N_3446,N_2626,N_2931);
nor U3447 (N_3447,N_2681,N_2844);
xnor U3448 (N_3448,N_2584,N_2585);
nor U3449 (N_3449,N_2639,N_2572);
nor U3450 (N_3450,N_2502,N_2763);
nor U3451 (N_3451,N_2862,N_2813);
nand U3452 (N_3452,N_2887,N_2884);
nor U3453 (N_3453,N_2854,N_2574);
or U3454 (N_3454,N_2627,N_2647);
xnor U3455 (N_3455,N_2901,N_2810);
or U3456 (N_3456,N_2720,N_2664);
nor U3457 (N_3457,N_2952,N_2828);
or U3458 (N_3458,N_2526,N_2859);
xnor U3459 (N_3459,N_2734,N_2600);
xnor U3460 (N_3460,N_2689,N_2943);
or U3461 (N_3461,N_2910,N_2844);
xnor U3462 (N_3462,N_2587,N_2803);
and U3463 (N_3463,N_2556,N_2585);
or U3464 (N_3464,N_2665,N_2938);
xnor U3465 (N_3465,N_2840,N_2855);
or U3466 (N_3466,N_2529,N_2688);
and U3467 (N_3467,N_2693,N_2917);
and U3468 (N_3468,N_2731,N_2608);
xnor U3469 (N_3469,N_2582,N_2959);
or U3470 (N_3470,N_2835,N_2918);
and U3471 (N_3471,N_2664,N_2618);
nor U3472 (N_3472,N_2745,N_2893);
nor U3473 (N_3473,N_2845,N_2926);
and U3474 (N_3474,N_2832,N_2869);
nand U3475 (N_3475,N_2806,N_2803);
nor U3476 (N_3476,N_2793,N_2508);
and U3477 (N_3477,N_2888,N_2558);
and U3478 (N_3478,N_2829,N_2938);
or U3479 (N_3479,N_2550,N_2735);
or U3480 (N_3480,N_2528,N_2727);
nand U3481 (N_3481,N_2602,N_2679);
or U3482 (N_3482,N_2550,N_2561);
or U3483 (N_3483,N_2520,N_2639);
nor U3484 (N_3484,N_2672,N_2674);
or U3485 (N_3485,N_2750,N_2965);
nand U3486 (N_3486,N_2975,N_2700);
nor U3487 (N_3487,N_2760,N_2550);
or U3488 (N_3488,N_2513,N_2956);
xnor U3489 (N_3489,N_2578,N_2972);
nand U3490 (N_3490,N_2541,N_2587);
nor U3491 (N_3491,N_2552,N_2577);
nand U3492 (N_3492,N_2900,N_2816);
xnor U3493 (N_3493,N_2838,N_2759);
and U3494 (N_3494,N_2772,N_2911);
xor U3495 (N_3495,N_2644,N_2918);
nand U3496 (N_3496,N_2806,N_2708);
and U3497 (N_3497,N_2673,N_2973);
xnor U3498 (N_3498,N_2788,N_2752);
xnor U3499 (N_3499,N_2664,N_2674);
or U3500 (N_3500,N_3438,N_3047);
nand U3501 (N_3501,N_3113,N_3285);
xor U3502 (N_3502,N_3280,N_3069);
nor U3503 (N_3503,N_3131,N_3450);
nor U3504 (N_3504,N_3020,N_3475);
or U3505 (N_3505,N_3390,N_3011);
nor U3506 (N_3506,N_3061,N_3425);
nor U3507 (N_3507,N_3054,N_3368);
xor U3508 (N_3508,N_3022,N_3350);
nor U3509 (N_3509,N_3072,N_3402);
nand U3510 (N_3510,N_3272,N_3299);
xnor U3511 (N_3511,N_3310,N_3330);
nor U3512 (N_3512,N_3370,N_3034);
and U3513 (N_3513,N_3363,N_3043);
nor U3514 (N_3514,N_3371,N_3440);
or U3515 (N_3515,N_3358,N_3093);
nor U3516 (N_3516,N_3426,N_3111);
nor U3517 (N_3517,N_3073,N_3052);
xor U3518 (N_3518,N_3441,N_3182);
or U3519 (N_3519,N_3319,N_3120);
xor U3520 (N_3520,N_3337,N_3463);
nand U3521 (N_3521,N_3449,N_3030);
and U3522 (N_3522,N_3278,N_3257);
or U3523 (N_3523,N_3179,N_3303);
and U3524 (N_3524,N_3322,N_3036);
xor U3525 (N_3525,N_3456,N_3457);
nor U3526 (N_3526,N_3238,N_3128);
or U3527 (N_3527,N_3185,N_3211);
or U3528 (N_3528,N_3486,N_3246);
nor U3529 (N_3529,N_3243,N_3263);
nor U3530 (N_3530,N_3461,N_3352);
and U3531 (N_3531,N_3119,N_3366);
nor U3532 (N_3532,N_3234,N_3469);
and U3533 (N_3533,N_3409,N_3194);
nor U3534 (N_3534,N_3088,N_3124);
and U3535 (N_3535,N_3178,N_3465);
or U3536 (N_3536,N_3288,N_3123);
nor U3537 (N_3537,N_3284,N_3283);
and U3538 (N_3538,N_3296,N_3496);
and U3539 (N_3539,N_3397,N_3217);
xnor U3540 (N_3540,N_3172,N_3304);
and U3541 (N_3541,N_3403,N_3129);
and U3542 (N_3542,N_3386,N_3139);
and U3543 (N_3543,N_3410,N_3023);
nand U3544 (N_3544,N_3376,N_3484);
nand U3545 (N_3545,N_3147,N_3029);
xor U3546 (N_3546,N_3408,N_3490);
and U3547 (N_3547,N_3464,N_3081);
xor U3548 (N_3548,N_3375,N_3167);
xnor U3549 (N_3549,N_3333,N_3364);
and U3550 (N_3550,N_3082,N_3313);
and U3551 (N_3551,N_3277,N_3068);
xor U3552 (N_3552,N_3476,N_3204);
or U3553 (N_3553,N_3325,N_3151);
xor U3554 (N_3554,N_3080,N_3374);
and U3555 (N_3555,N_3261,N_3404);
and U3556 (N_3556,N_3242,N_3156);
nor U3557 (N_3557,N_3339,N_3146);
and U3558 (N_3558,N_3003,N_3389);
nand U3559 (N_3559,N_3033,N_3354);
and U3560 (N_3560,N_3434,N_3423);
xor U3561 (N_3561,N_3005,N_3250);
nand U3562 (N_3562,N_3323,N_3481);
nand U3563 (N_3563,N_3420,N_3032);
nand U3564 (N_3564,N_3431,N_3021);
and U3565 (N_3565,N_3104,N_3437);
and U3566 (N_3566,N_3031,N_3230);
and U3567 (N_3567,N_3012,N_3110);
nand U3568 (N_3568,N_3215,N_3164);
nor U3569 (N_3569,N_3380,N_3237);
and U3570 (N_3570,N_3485,N_3017);
nand U3571 (N_3571,N_3208,N_3293);
xor U3572 (N_3572,N_3187,N_3415);
nor U3573 (N_3573,N_3133,N_3361);
and U3574 (N_3574,N_3331,N_3258);
nand U3575 (N_3575,N_3265,N_3377);
or U3576 (N_3576,N_3216,N_3384);
and U3577 (N_3577,N_3489,N_3221);
or U3578 (N_3578,N_3143,N_3060);
xnor U3579 (N_3579,N_3168,N_3024);
and U3580 (N_3580,N_3355,N_3196);
xnor U3581 (N_3581,N_3276,N_3161);
or U3582 (N_3582,N_3422,N_3351);
nand U3583 (N_3583,N_3395,N_3341);
or U3584 (N_3584,N_3347,N_3270);
or U3585 (N_3585,N_3180,N_3412);
nor U3586 (N_3586,N_3136,N_3436);
xnor U3587 (N_3587,N_3455,N_3000);
or U3588 (N_3588,N_3378,N_3447);
nor U3589 (N_3589,N_3326,N_3349);
xor U3590 (N_3590,N_3162,N_3317);
or U3591 (N_3591,N_3228,N_3114);
or U3592 (N_3592,N_3454,N_3078);
and U3593 (N_3593,N_3112,N_3346);
xnor U3594 (N_3594,N_3106,N_3253);
nor U3595 (N_3595,N_3096,N_3065);
xnor U3596 (N_3596,N_3055,N_3398);
or U3597 (N_3597,N_3035,N_3399);
or U3598 (N_3598,N_3247,N_3057);
or U3599 (N_3599,N_3248,N_3342);
nand U3600 (N_3600,N_3497,N_3019);
xnor U3601 (N_3601,N_3307,N_3004);
and U3602 (N_3602,N_3117,N_3206);
and U3603 (N_3603,N_3101,N_3477);
or U3604 (N_3604,N_3443,N_3446);
nor U3605 (N_3605,N_3026,N_3079);
nor U3606 (N_3606,N_3311,N_3362);
nor U3607 (N_3607,N_3344,N_3214);
nand U3608 (N_3608,N_3294,N_3467);
nand U3609 (N_3609,N_3109,N_3199);
and U3610 (N_3610,N_3292,N_3235);
xor U3611 (N_3611,N_3046,N_3498);
and U3612 (N_3612,N_3255,N_3121);
or U3613 (N_3613,N_3207,N_3066);
nor U3614 (N_3614,N_3462,N_3049);
and U3615 (N_3615,N_3122,N_3040);
xnor U3616 (N_3616,N_3316,N_3212);
nand U3617 (N_3617,N_3062,N_3432);
nor U3618 (N_3618,N_3166,N_3295);
nor U3619 (N_3619,N_3324,N_3421);
xnor U3620 (N_3620,N_3345,N_3186);
or U3621 (N_3621,N_3063,N_3279);
xor U3622 (N_3622,N_3083,N_3138);
nand U3623 (N_3623,N_3448,N_3134);
nor U3624 (N_3624,N_3209,N_3287);
nor U3625 (N_3625,N_3100,N_3002);
nand U3626 (N_3626,N_3274,N_3419);
nor U3627 (N_3627,N_3148,N_3458);
xnor U3628 (N_3628,N_3271,N_3176);
xnor U3629 (N_3629,N_3126,N_3190);
xnor U3630 (N_3630,N_3058,N_3302);
nor U3631 (N_3631,N_3094,N_3130);
nand U3632 (N_3632,N_3150,N_3039);
and U3633 (N_3633,N_3343,N_3144);
nand U3634 (N_3634,N_3396,N_3306);
or U3635 (N_3635,N_3244,N_3142);
or U3636 (N_3636,N_3241,N_3321);
and U3637 (N_3637,N_3290,N_3291);
nand U3638 (N_3638,N_3091,N_3008);
and U3639 (N_3639,N_3125,N_3379);
or U3640 (N_3640,N_3018,N_3487);
xor U3641 (N_3641,N_3259,N_3226);
or U3642 (N_3642,N_3200,N_3460);
xor U3643 (N_3643,N_3256,N_3075);
or U3644 (N_3644,N_3045,N_3471);
nand U3645 (N_3645,N_3348,N_3195);
nand U3646 (N_3646,N_3001,N_3297);
xnor U3647 (N_3647,N_3098,N_3251);
and U3648 (N_3648,N_3245,N_3382);
and U3649 (N_3649,N_3359,N_3466);
nor U3650 (N_3650,N_3225,N_3479);
nor U3651 (N_3651,N_3159,N_3087);
nand U3652 (N_3652,N_3494,N_3273);
or U3653 (N_3653,N_3239,N_3407);
xnor U3654 (N_3654,N_3340,N_3427);
xnor U3655 (N_3655,N_3218,N_3452);
nor U3656 (N_3656,N_3413,N_3160);
xor U3657 (N_3657,N_3157,N_3070);
nand U3658 (N_3658,N_3492,N_3202);
nor U3659 (N_3659,N_3388,N_3428);
xor U3660 (N_3660,N_3472,N_3095);
nand U3661 (N_3661,N_3071,N_3373);
nor U3662 (N_3662,N_3480,N_3177);
nor U3663 (N_3663,N_3411,N_3116);
xor U3664 (N_3664,N_3468,N_3491);
or U3665 (N_3665,N_3338,N_3483);
xnor U3666 (N_3666,N_3028,N_3356);
nand U3667 (N_3667,N_3184,N_3353);
or U3668 (N_3668,N_3372,N_3149);
and U3669 (N_3669,N_3459,N_3015);
and U3670 (N_3670,N_3406,N_3328);
nand U3671 (N_3671,N_3418,N_3429);
or U3672 (N_3672,N_3268,N_3289);
and U3673 (N_3673,N_3391,N_3169);
or U3674 (N_3674,N_3170,N_3016);
nand U3675 (N_3675,N_3442,N_3050);
nor U3676 (N_3676,N_3329,N_3308);
nor U3677 (N_3677,N_3077,N_3414);
or U3678 (N_3678,N_3056,N_3335);
and U3679 (N_3679,N_3264,N_3232);
xor U3680 (N_3680,N_3181,N_3025);
nand U3681 (N_3681,N_3163,N_3267);
and U3682 (N_3682,N_3145,N_3013);
or U3683 (N_3683,N_3127,N_3198);
nand U3684 (N_3684,N_3010,N_3041);
nand U3685 (N_3685,N_3493,N_3229);
nand U3686 (N_3686,N_3155,N_3387);
nand U3687 (N_3687,N_3192,N_3064);
nand U3688 (N_3688,N_3191,N_3223);
and U3689 (N_3689,N_3286,N_3269);
nand U3690 (N_3690,N_3260,N_3435);
nor U3691 (N_3691,N_3115,N_3249);
xnor U3692 (N_3692,N_3108,N_3165);
and U3693 (N_3693,N_3220,N_3135);
nand U3694 (N_3694,N_3006,N_3014);
nand U3695 (N_3695,N_3365,N_3171);
nand U3696 (N_3696,N_3394,N_3282);
xor U3697 (N_3697,N_3141,N_3400);
or U3698 (N_3698,N_3281,N_3044);
and U3699 (N_3699,N_3474,N_3417);
or U3700 (N_3700,N_3059,N_3275);
xor U3701 (N_3701,N_3038,N_3367);
and U3702 (N_3702,N_3478,N_3314);
nand U3703 (N_3703,N_3318,N_3007);
and U3704 (N_3704,N_3357,N_3084);
nor U3705 (N_3705,N_3174,N_3027);
and U3706 (N_3706,N_3381,N_3140);
xnor U3707 (N_3707,N_3392,N_3227);
and U3708 (N_3708,N_3193,N_3315);
or U3709 (N_3709,N_3327,N_3444);
and U3710 (N_3710,N_3219,N_3300);
or U3711 (N_3711,N_3042,N_3188);
nand U3712 (N_3712,N_3336,N_3086);
and U3713 (N_3713,N_3103,N_3118);
and U3714 (N_3714,N_3213,N_3222);
nand U3715 (N_3715,N_3301,N_3102);
or U3716 (N_3716,N_3231,N_3153);
nor U3717 (N_3717,N_3090,N_3252);
or U3718 (N_3718,N_3298,N_3439);
xor U3719 (N_3719,N_3053,N_3254);
nand U3720 (N_3720,N_3424,N_3453);
or U3721 (N_3721,N_3152,N_3233);
and U3722 (N_3722,N_3089,N_3360);
and U3723 (N_3723,N_3158,N_3393);
and U3724 (N_3724,N_3305,N_3137);
or U3725 (N_3725,N_3488,N_3416);
xor U3726 (N_3726,N_3499,N_3197);
nor U3727 (N_3727,N_3037,N_3210);
and U3728 (N_3728,N_3074,N_3203);
or U3729 (N_3729,N_3433,N_3430);
or U3730 (N_3730,N_3009,N_3092);
and U3731 (N_3731,N_3470,N_3189);
or U3732 (N_3732,N_3320,N_3051);
xor U3733 (N_3733,N_3201,N_3262);
xnor U3734 (N_3734,N_3097,N_3205);
xor U3735 (N_3735,N_3334,N_3369);
or U3736 (N_3736,N_3132,N_3224);
nor U3737 (N_3737,N_3105,N_3085);
xor U3738 (N_3738,N_3482,N_3154);
and U3739 (N_3739,N_3332,N_3107);
nand U3740 (N_3740,N_3309,N_3076);
nor U3741 (N_3741,N_3383,N_3405);
xor U3742 (N_3742,N_3240,N_3385);
and U3743 (N_3743,N_3236,N_3175);
nor U3744 (N_3744,N_3495,N_3401);
nor U3745 (N_3745,N_3266,N_3173);
and U3746 (N_3746,N_3048,N_3445);
xnor U3747 (N_3747,N_3312,N_3067);
xor U3748 (N_3748,N_3451,N_3183);
nand U3749 (N_3749,N_3099,N_3473);
or U3750 (N_3750,N_3237,N_3356);
nor U3751 (N_3751,N_3152,N_3151);
nand U3752 (N_3752,N_3473,N_3141);
or U3753 (N_3753,N_3333,N_3289);
xor U3754 (N_3754,N_3369,N_3364);
nor U3755 (N_3755,N_3161,N_3094);
nand U3756 (N_3756,N_3467,N_3122);
and U3757 (N_3757,N_3310,N_3118);
nand U3758 (N_3758,N_3273,N_3176);
and U3759 (N_3759,N_3491,N_3227);
and U3760 (N_3760,N_3439,N_3314);
or U3761 (N_3761,N_3099,N_3374);
or U3762 (N_3762,N_3102,N_3214);
nand U3763 (N_3763,N_3264,N_3038);
and U3764 (N_3764,N_3173,N_3030);
nand U3765 (N_3765,N_3272,N_3257);
and U3766 (N_3766,N_3483,N_3397);
and U3767 (N_3767,N_3267,N_3330);
nand U3768 (N_3768,N_3063,N_3487);
or U3769 (N_3769,N_3121,N_3382);
nand U3770 (N_3770,N_3255,N_3357);
nand U3771 (N_3771,N_3057,N_3364);
xnor U3772 (N_3772,N_3432,N_3228);
nand U3773 (N_3773,N_3494,N_3029);
nor U3774 (N_3774,N_3251,N_3410);
nor U3775 (N_3775,N_3118,N_3314);
or U3776 (N_3776,N_3251,N_3185);
nor U3777 (N_3777,N_3376,N_3310);
nor U3778 (N_3778,N_3058,N_3101);
nand U3779 (N_3779,N_3472,N_3133);
nand U3780 (N_3780,N_3205,N_3256);
xnor U3781 (N_3781,N_3354,N_3169);
nor U3782 (N_3782,N_3460,N_3189);
and U3783 (N_3783,N_3377,N_3450);
xor U3784 (N_3784,N_3406,N_3154);
and U3785 (N_3785,N_3097,N_3384);
and U3786 (N_3786,N_3402,N_3212);
nor U3787 (N_3787,N_3279,N_3233);
xor U3788 (N_3788,N_3333,N_3200);
nor U3789 (N_3789,N_3198,N_3338);
nor U3790 (N_3790,N_3309,N_3331);
nand U3791 (N_3791,N_3117,N_3275);
and U3792 (N_3792,N_3415,N_3458);
and U3793 (N_3793,N_3343,N_3116);
and U3794 (N_3794,N_3290,N_3429);
nand U3795 (N_3795,N_3224,N_3372);
or U3796 (N_3796,N_3445,N_3202);
or U3797 (N_3797,N_3498,N_3008);
nand U3798 (N_3798,N_3013,N_3390);
or U3799 (N_3799,N_3159,N_3010);
nand U3800 (N_3800,N_3084,N_3393);
or U3801 (N_3801,N_3472,N_3055);
xnor U3802 (N_3802,N_3232,N_3202);
or U3803 (N_3803,N_3250,N_3197);
nand U3804 (N_3804,N_3063,N_3272);
and U3805 (N_3805,N_3149,N_3004);
and U3806 (N_3806,N_3127,N_3342);
and U3807 (N_3807,N_3333,N_3220);
nor U3808 (N_3808,N_3020,N_3181);
xor U3809 (N_3809,N_3331,N_3181);
nor U3810 (N_3810,N_3177,N_3441);
nor U3811 (N_3811,N_3139,N_3051);
nor U3812 (N_3812,N_3099,N_3264);
xnor U3813 (N_3813,N_3259,N_3171);
and U3814 (N_3814,N_3466,N_3115);
nor U3815 (N_3815,N_3261,N_3018);
or U3816 (N_3816,N_3259,N_3101);
nand U3817 (N_3817,N_3430,N_3234);
or U3818 (N_3818,N_3455,N_3294);
and U3819 (N_3819,N_3017,N_3063);
xor U3820 (N_3820,N_3117,N_3349);
nor U3821 (N_3821,N_3085,N_3145);
or U3822 (N_3822,N_3401,N_3020);
and U3823 (N_3823,N_3382,N_3193);
nand U3824 (N_3824,N_3439,N_3104);
nand U3825 (N_3825,N_3351,N_3063);
and U3826 (N_3826,N_3269,N_3084);
or U3827 (N_3827,N_3465,N_3497);
xor U3828 (N_3828,N_3432,N_3195);
and U3829 (N_3829,N_3490,N_3230);
nor U3830 (N_3830,N_3239,N_3019);
xnor U3831 (N_3831,N_3481,N_3495);
and U3832 (N_3832,N_3297,N_3482);
or U3833 (N_3833,N_3020,N_3371);
nor U3834 (N_3834,N_3021,N_3026);
or U3835 (N_3835,N_3306,N_3204);
xor U3836 (N_3836,N_3299,N_3349);
and U3837 (N_3837,N_3407,N_3430);
and U3838 (N_3838,N_3328,N_3161);
or U3839 (N_3839,N_3306,N_3478);
nand U3840 (N_3840,N_3003,N_3146);
nand U3841 (N_3841,N_3418,N_3054);
nor U3842 (N_3842,N_3258,N_3454);
nand U3843 (N_3843,N_3268,N_3481);
nand U3844 (N_3844,N_3321,N_3144);
or U3845 (N_3845,N_3174,N_3410);
or U3846 (N_3846,N_3460,N_3181);
nand U3847 (N_3847,N_3247,N_3429);
nor U3848 (N_3848,N_3073,N_3320);
and U3849 (N_3849,N_3301,N_3173);
xnor U3850 (N_3850,N_3173,N_3357);
nand U3851 (N_3851,N_3118,N_3301);
nand U3852 (N_3852,N_3180,N_3199);
nor U3853 (N_3853,N_3281,N_3473);
or U3854 (N_3854,N_3420,N_3399);
nand U3855 (N_3855,N_3027,N_3232);
nor U3856 (N_3856,N_3353,N_3189);
nand U3857 (N_3857,N_3035,N_3279);
xnor U3858 (N_3858,N_3367,N_3380);
and U3859 (N_3859,N_3461,N_3086);
and U3860 (N_3860,N_3158,N_3255);
or U3861 (N_3861,N_3373,N_3374);
xnor U3862 (N_3862,N_3355,N_3125);
or U3863 (N_3863,N_3349,N_3493);
nor U3864 (N_3864,N_3442,N_3098);
and U3865 (N_3865,N_3258,N_3456);
nor U3866 (N_3866,N_3360,N_3328);
nor U3867 (N_3867,N_3038,N_3438);
nor U3868 (N_3868,N_3173,N_3259);
and U3869 (N_3869,N_3287,N_3050);
or U3870 (N_3870,N_3444,N_3329);
and U3871 (N_3871,N_3314,N_3161);
nand U3872 (N_3872,N_3353,N_3451);
nor U3873 (N_3873,N_3051,N_3377);
xor U3874 (N_3874,N_3442,N_3408);
nor U3875 (N_3875,N_3447,N_3290);
nand U3876 (N_3876,N_3465,N_3267);
and U3877 (N_3877,N_3335,N_3491);
or U3878 (N_3878,N_3197,N_3326);
nand U3879 (N_3879,N_3177,N_3244);
and U3880 (N_3880,N_3346,N_3199);
nor U3881 (N_3881,N_3044,N_3410);
or U3882 (N_3882,N_3081,N_3322);
xnor U3883 (N_3883,N_3414,N_3386);
xor U3884 (N_3884,N_3037,N_3057);
or U3885 (N_3885,N_3169,N_3241);
xor U3886 (N_3886,N_3121,N_3175);
xor U3887 (N_3887,N_3012,N_3246);
xnor U3888 (N_3888,N_3342,N_3445);
nor U3889 (N_3889,N_3271,N_3247);
and U3890 (N_3890,N_3470,N_3221);
nand U3891 (N_3891,N_3462,N_3075);
xor U3892 (N_3892,N_3369,N_3264);
and U3893 (N_3893,N_3004,N_3464);
and U3894 (N_3894,N_3436,N_3025);
nor U3895 (N_3895,N_3439,N_3170);
xnor U3896 (N_3896,N_3255,N_3312);
nor U3897 (N_3897,N_3116,N_3496);
nor U3898 (N_3898,N_3151,N_3352);
nand U3899 (N_3899,N_3153,N_3264);
nor U3900 (N_3900,N_3220,N_3180);
nor U3901 (N_3901,N_3378,N_3424);
xor U3902 (N_3902,N_3470,N_3387);
nand U3903 (N_3903,N_3013,N_3071);
xor U3904 (N_3904,N_3244,N_3249);
and U3905 (N_3905,N_3275,N_3374);
nor U3906 (N_3906,N_3364,N_3300);
and U3907 (N_3907,N_3011,N_3180);
and U3908 (N_3908,N_3388,N_3153);
nor U3909 (N_3909,N_3397,N_3046);
xor U3910 (N_3910,N_3189,N_3075);
nor U3911 (N_3911,N_3242,N_3053);
nor U3912 (N_3912,N_3114,N_3354);
or U3913 (N_3913,N_3417,N_3072);
xnor U3914 (N_3914,N_3145,N_3422);
nor U3915 (N_3915,N_3113,N_3216);
or U3916 (N_3916,N_3385,N_3468);
xnor U3917 (N_3917,N_3118,N_3179);
nor U3918 (N_3918,N_3410,N_3453);
nor U3919 (N_3919,N_3416,N_3281);
and U3920 (N_3920,N_3147,N_3311);
nor U3921 (N_3921,N_3408,N_3223);
and U3922 (N_3922,N_3309,N_3317);
nor U3923 (N_3923,N_3370,N_3091);
nor U3924 (N_3924,N_3074,N_3161);
nor U3925 (N_3925,N_3257,N_3235);
or U3926 (N_3926,N_3003,N_3190);
nor U3927 (N_3927,N_3253,N_3404);
nor U3928 (N_3928,N_3152,N_3276);
or U3929 (N_3929,N_3207,N_3249);
nor U3930 (N_3930,N_3071,N_3434);
nor U3931 (N_3931,N_3327,N_3397);
nor U3932 (N_3932,N_3018,N_3310);
or U3933 (N_3933,N_3297,N_3385);
or U3934 (N_3934,N_3025,N_3010);
xnor U3935 (N_3935,N_3444,N_3357);
and U3936 (N_3936,N_3497,N_3193);
nand U3937 (N_3937,N_3110,N_3428);
nor U3938 (N_3938,N_3470,N_3175);
xor U3939 (N_3939,N_3443,N_3306);
and U3940 (N_3940,N_3334,N_3432);
and U3941 (N_3941,N_3358,N_3440);
xor U3942 (N_3942,N_3246,N_3383);
xnor U3943 (N_3943,N_3259,N_3004);
and U3944 (N_3944,N_3256,N_3105);
xnor U3945 (N_3945,N_3447,N_3028);
and U3946 (N_3946,N_3185,N_3451);
or U3947 (N_3947,N_3201,N_3354);
nor U3948 (N_3948,N_3147,N_3009);
nand U3949 (N_3949,N_3371,N_3379);
xor U3950 (N_3950,N_3473,N_3146);
nor U3951 (N_3951,N_3451,N_3472);
and U3952 (N_3952,N_3225,N_3191);
nand U3953 (N_3953,N_3333,N_3415);
nand U3954 (N_3954,N_3220,N_3011);
nand U3955 (N_3955,N_3230,N_3205);
and U3956 (N_3956,N_3340,N_3144);
xnor U3957 (N_3957,N_3355,N_3264);
or U3958 (N_3958,N_3047,N_3187);
and U3959 (N_3959,N_3302,N_3159);
or U3960 (N_3960,N_3165,N_3037);
and U3961 (N_3961,N_3365,N_3405);
and U3962 (N_3962,N_3295,N_3117);
nand U3963 (N_3963,N_3269,N_3146);
xnor U3964 (N_3964,N_3298,N_3009);
or U3965 (N_3965,N_3419,N_3230);
nand U3966 (N_3966,N_3188,N_3278);
nand U3967 (N_3967,N_3250,N_3143);
and U3968 (N_3968,N_3268,N_3100);
or U3969 (N_3969,N_3230,N_3496);
or U3970 (N_3970,N_3280,N_3476);
or U3971 (N_3971,N_3091,N_3420);
and U3972 (N_3972,N_3130,N_3098);
or U3973 (N_3973,N_3161,N_3337);
xnor U3974 (N_3974,N_3155,N_3048);
xnor U3975 (N_3975,N_3248,N_3382);
xor U3976 (N_3976,N_3239,N_3112);
nor U3977 (N_3977,N_3004,N_3024);
or U3978 (N_3978,N_3419,N_3118);
xnor U3979 (N_3979,N_3311,N_3131);
xnor U3980 (N_3980,N_3149,N_3293);
nor U3981 (N_3981,N_3183,N_3390);
nor U3982 (N_3982,N_3143,N_3474);
nor U3983 (N_3983,N_3290,N_3377);
nand U3984 (N_3984,N_3237,N_3418);
or U3985 (N_3985,N_3233,N_3310);
nor U3986 (N_3986,N_3167,N_3304);
nor U3987 (N_3987,N_3208,N_3076);
nor U3988 (N_3988,N_3341,N_3399);
or U3989 (N_3989,N_3344,N_3306);
or U3990 (N_3990,N_3388,N_3205);
and U3991 (N_3991,N_3069,N_3350);
nand U3992 (N_3992,N_3292,N_3209);
and U3993 (N_3993,N_3280,N_3150);
and U3994 (N_3994,N_3141,N_3230);
or U3995 (N_3995,N_3180,N_3267);
nor U3996 (N_3996,N_3264,N_3391);
or U3997 (N_3997,N_3193,N_3096);
or U3998 (N_3998,N_3065,N_3342);
and U3999 (N_3999,N_3085,N_3057);
nand U4000 (N_4000,N_3833,N_3817);
nand U4001 (N_4001,N_3647,N_3678);
xor U4002 (N_4002,N_3625,N_3930);
or U4003 (N_4003,N_3715,N_3606);
or U4004 (N_4004,N_3649,N_3552);
or U4005 (N_4005,N_3858,N_3758);
and U4006 (N_4006,N_3811,N_3568);
or U4007 (N_4007,N_3791,N_3921);
nand U4008 (N_4008,N_3897,N_3653);
nand U4009 (N_4009,N_3726,N_3820);
nor U4010 (N_4010,N_3727,N_3940);
or U4011 (N_4011,N_3819,N_3525);
nand U4012 (N_4012,N_3970,N_3751);
and U4013 (N_4013,N_3759,N_3809);
or U4014 (N_4014,N_3907,N_3619);
nor U4015 (N_4015,N_3692,N_3533);
nand U4016 (N_4016,N_3771,N_3676);
or U4017 (N_4017,N_3866,N_3696);
nand U4018 (N_4018,N_3735,N_3863);
nand U4019 (N_4019,N_3754,N_3616);
nand U4020 (N_4020,N_3629,N_3974);
nor U4021 (N_4021,N_3873,N_3986);
and U4022 (N_4022,N_3802,N_3946);
nand U4023 (N_4023,N_3982,N_3859);
nand U4024 (N_4024,N_3740,N_3519);
nand U4025 (N_4025,N_3908,N_3768);
xor U4026 (N_4026,N_3773,N_3520);
and U4027 (N_4027,N_3892,N_3646);
or U4028 (N_4028,N_3731,N_3951);
and U4029 (N_4029,N_3687,N_3502);
nor U4030 (N_4030,N_3681,N_3673);
or U4031 (N_4031,N_3975,N_3633);
and U4032 (N_4032,N_3793,N_3529);
nor U4033 (N_4033,N_3746,N_3536);
xnor U4034 (N_4034,N_3508,N_3770);
or U4035 (N_4035,N_3621,N_3654);
and U4036 (N_4036,N_3860,N_3530);
or U4037 (N_4037,N_3882,N_3643);
nand U4038 (N_4038,N_3713,N_3729);
nor U4039 (N_4039,N_3602,N_3899);
and U4040 (N_4040,N_3842,N_3900);
xnor U4041 (N_4041,N_3853,N_3592);
and U4042 (N_4042,N_3814,N_3821);
and U4043 (N_4043,N_3560,N_3664);
nor U4044 (N_4044,N_3737,N_3719);
nand U4045 (N_4045,N_3682,N_3541);
nor U4046 (N_4046,N_3569,N_3763);
xnor U4047 (N_4047,N_3652,N_3547);
and U4048 (N_4048,N_3948,N_3810);
or U4049 (N_4049,N_3925,N_3512);
xor U4050 (N_4050,N_3697,N_3571);
or U4051 (N_4051,N_3599,N_3874);
nor U4052 (N_4052,N_3867,N_3794);
xor U4053 (N_4053,N_3688,N_3706);
and U4054 (N_4054,N_3638,N_3884);
and U4055 (N_4055,N_3941,N_3999);
nor U4056 (N_4056,N_3808,N_3608);
nor U4057 (N_4057,N_3852,N_3699);
or U4058 (N_4058,N_3683,N_3955);
or U4059 (N_4059,N_3934,N_3909);
nand U4060 (N_4060,N_3632,N_3644);
nand U4061 (N_4061,N_3558,N_3889);
nor U4062 (N_4062,N_3958,N_3650);
xor U4063 (N_4063,N_3661,N_3985);
nor U4064 (N_4064,N_3756,N_3677);
and U4065 (N_4065,N_3983,N_3642);
nor U4066 (N_4066,N_3967,N_3916);
nand U4067 (N_4067,N_3767,N_3589);
xor U4068 (N_4068,N_3733,N_3834);
and U4069 (N_4069,N_3708,N_3546);
or U4070 (N_4070,N_3670,N_3857);
nor U4071 (N_4071,N_3947,N_3666);
and U4072 (N_4072,N_3564,N_3898);
nor U4073 (N_4073,N_3700,N_3949);
xor U4074 (N_4074,N_3917,N_3543);
nor U4075 (N_4075,N_3601,N_3903);
or U4076 (N_4076,N_3618,N_3789);
nor U4077 (N_4077,N_3877,N_3838);
xnor U4078 (N_4078,N_3504,N_3827);
or U4079 (N_4079,N_3918,N_3843);
or U4080 (N_4080,N_3575,N_3559);
xor U4081 (N_4081,N_3660,N_3831);
or U4082 (N_4082,N_3718,N_3829);
and U4083 (N_4083,N_3736,N_3938);
nor U4084 (N_4084,N_3963,N_3624);
xnor U4085 (N_4085,N_3610,N_3871);
or U4086 (N_4086,N_3855,N_3787);
or U4087 (N_4087,N_3805,N_3956);
nand U4088 (N_4088,N_3570,N_3876);
xor U4089 (N_4089,N_3905,N_3895);
xor U4090 (N_4090,N_3836,N_3851);
or U4091 (N_4091,N_3840,N_3937);
nand U4092 (N_4092,N_3962,N_3521);
nor U4093 (N_4093,N_3728,N_3943);
nor U4094 (N_4094,N_3583,N_3639);
or U4095 (N_4095,N_3505,N_3741);
or U4096 (N_4096,N_3659,N_3698);
xnor U4097 (N_4097,N_3865,N_3611);
nor U4098 (N_4098,N_3813,N_3792);
and U4099 (N_4099,N_3801,N_3932);
xnor U4100 (N_4100,N_3747,N_3785);
nor U4101 (N_4101,N_3693,N_3997);
or U4102 (N_4102,N_3607,N_3662);
nand U4103 (N_4103,N_3712,N_3984);
nor U4104 (N_4104,N_3849,N_3604);
or U4105 (N_4105,N_3954,N_3637);
nor U4106 (N_4106,N_3671,N_3825);
nand U4107 (N_4107,N_3596,N_3515);
xnor U4108 (N_4108,N_3879,N_3665);
xor U4109 (N_4109,N_3630,N_3636);
and U4110 (N_4110,N_3945,N_3517);
nor U4111 (N_4111,N_3622,N_3545);
nor U4112 (N_4112,N_3830,N_3769);
nand U4113 (N_4113,N_3510,N_3847);
or U4114 (N_4114,N_3658,N_3710);
or U4115 (N_4115,N_3548,N_3887);
nor U4116 (N_4116,N_3919,N_3878);
nor U4117 (N_4117,N_3837,N_3532);
and U4118 (N_4118,N_3904,N_3509);
xor U4119 (N_4119,N_3861,N_3960);
and U4120 (N_4120,N_3565,N_3913);
nor U4121 (N_4121,N_3544,N_3640);
nor U4122 (N_4122,N_3701,N_3511);
and U4123 (N_4123,N_3760,N_3645);
nand U4124 (N_4124,N_3657,N_3527);
xor U4125 (N_4125,N_3503,N_3780);
or U4126 (N_4126,N_3804,N_3862);
and U4127 (N_4127,N_3922,N_3524);
nor U4128 (N_4128,N_3690,N_3709);
or U4129 (N_4129,N_3500,N_3846);
nor U4130 (N_4130,N_3839,N_3989);
nand U4131 (N_4131,N_3703,N_3806);
nand U4132 (N_4132,N_3753,N_3824);
nand U4133 (N_4133,N_3781,N_3912);
nand U4134 (N_4134,N_3542,N_3694);
nand U4135 (N_4135,N_3844,N_3572);
nor U4136 (N_4136,N_3902,N_3550);
and U4137 (N_4137,N_3957,N_3961);
nor U4138 (N_4138,N_3920,N_3686);
and U4139 (N_4139,N_3523,N_3577);
nand U4140 (N_4140,N_3518,N_3581);
nand U4141 (N_4141,N_3929,N_3812);
and U4142 (N_4142,N_3883,N_3695);
or U4143 (N_4143,N_3628,N_3988);
or U4144 (N_4144,N_3927,N_3723);
or U4145 (N_4145,N_3672,N_3864);
and U4146 (N_4146,N_3627,N_3972);
or U4147 (N_4147,N_3528,N_3755);
nand U4148 (N_4148,N_3689,N_3551);
nand U4149 (N_4149,N_3924,N_3563);
and U4150 (N_4150,N_3935,N_3561);
and U4151 (N_4151,N_3894,N_3777);
nor U4152 (N_4152,N_3772,N_3993);
xnor U4153 (N_4153,N_3591,N_3612);
nor U4154 (N_4154,N_3582,N_3557);
and U4155 (N_4155,N_3868,N_3501);
or U4156 (N_4156,N_3964,N_3750);
xnor U4157 (N_4157,N_3680,N_3722);
and U4158 (N_4158,N_3641,N_3888);
or U4159 (N_4159,N_3605,N_3573);
nor U4160 (N_4160,N_3953,N_3835);
xnor U4161 (N_4161,N_3526,N_3562);
xor U4162 (N_4162,N_3744,N_3617);
xnor U4163 (N_4163,N_3936,N_3885);
or U4164 (N_4164,N_3782,N_3790);
and U4165 (N_4165,N_3631,N_3702);
and U4166 (N_4166,N_3634,N_3595);
xor U4167 (N_4167,N_3973,N_3707);
nand U4168 (N_4168,N_3590,N_3669);
xnor U4169 (N_4169,N_3798,N_3614);
nand U4170 (N_4170,N_3748,N_3648);
nor U4171 (N_4171,N_3620,N_3663);
nor U4172 (N_4172,N_3797,N_3845);
nor U4173 (N_4173,N_3765,N_3593);
and U4174 (N_4174,N_3950,N_3734);
nand U4175 (N_4175,N_3626,N_3784);
xnor U4176 (N_4176,N_3600,N_3911);
nand U4177 (N_4177,N_3776,N_3995);
nor U4178 (N_4178,N_3779,N_3942);
or U4179 (N_4179,N_3971,N_3796);
xnor U4180 (N_4180,N_3991,N_3788);
xnor U4181 (N_4181,N_3506,N_3538);
and U4182 (N_4182,N_3705,N_3588);
nor U4183 (N_4183,N_3549,N_3783);
and U4184 (N_4184,N_3535,N_3981);
nand U4185 (N_4185,N_3980,N_3739);
nand U4186 (N_4186,N_3881,N_3513);
or U4187 (N_4187,N_3968,N_3800);
and U4188 (N_4188,N_3603,N_3507);
or U4189 (N_4189,N_3933,N_3959);
or U4190 (N_4190,N_3965,N_3704);
nor U4191 (N_4191,N_3786,N_3615);
nand U4192 (N_4192,N_3743,N_3635);
and U4193 (N_4193,N_3761,N_3574);
or U4194 (N_4194,N_3807,N_3766);
or U4195 (N_4195,N_3685,N_3613);
nand U4196 (N_4196,N_3870,N_3742);
and U4197 (N_4197,N_3969,N_3799);
or U4198 (N_4198,N_3752,N_3774);
or U4199 (N_4199,N_3816,N_3976);
and U4200 (N_4200,N_3540,N_3872);
nand U4201 (N_4201,N_3762,N_3966);
or U4202 (N_4202,N_3890,N_3778);
nor U4203 (N_4203,N_3841,N_3578);
nor U4204 (N_4204,N_3725,N_3994);
nand U4205 (N_4205,N_3609,N_3914);
nor U4206 (N_4206,N_3679,N_3724);
and U4207 (N_4207,N_3585,N_3893);
xor U4208 (N_4208,N_3514,N_3556);
xnor U4209 (N_4209,N_3716,N_3952);
nor U4210 (N_4210,N_3553,N_3566);
nand U4211 (N_4211,N_3832,N_3714);
xor U4212 (N_4212,N_3823,N_3854);
xor U4213 (N_4213,N_3539,N_3730);
nor U4214 (N_4214,N_3534,N_3655);
or U4215 (N_4215,N_3717,N_3555);
xor U4216 (N_4216,N_3554,N_3667);
nor U4217 (N_4217,N_3977,N_3998);
xor U4218 (N_4218,N_3576,N_3928);
nor U4219 (N_4219,N_3869,N_3522);
nor U4220 (N_4220,N_3749,N_3979);
xnor U4221 (N_4221,N_3886,N_3651);
or U4222 (N_4222,N_3992,N_3775);
nor U4223 (N_4223,N_3516,N_3926);
xnor U4224 (N_4224,N_3880,N_3915);
or U4225 (N_4225,N_3910,N_3691);
xor U4226 (N_4226,N_3896,N_3848);
nand U4227 (N_4227,N_3537,N_3675);
nor U4228 (N_4228,N_3587,N_3567);
or U4229 (N_4229,N_3901,N_3931);
or U4230 (N_4230,N_3711,N_3584);
nor U4231 (N_4231,N_3822,N_3732);
xnor U4232 (N_4232,N_3990,N_3803);
nor U4233 (N_4233,N_3586,N_3738);
nand U4234 (N_4234,N_3987,N_3668);
nor U4235 (N_4235,N_3764,N_3656);
nand U4236 (N_4236,N_3795,N_3996);
or U4237 (N_4237,N_3674,N_3906);
xor U4238 (N_4238,N_3818,N_3580);
or U4239 (N_4239,N_3684,N_3856);
nor U4240 (N_4240,N_3923,N_3875);
nand U4241 (N_4241,N_3531,N_3594);
and U4242 (N_4242,N_3891,N_3757);
nor U4243 (N_4243,N_3944,N_3579);
xnor U4244 (N_4244,N_3745,N_3597);
or U4245 (N_4245,N_3939,N_3815);
and U4246 (N_4246,N_3720,N_3850);
or U4247 (N_4247,N_3826,N_3598);
xnor U4248 (N_4248,N_3828,N_3623);
and U4249 (N_4249,N_3978,N_3721);
or U4250 (N_4250,N_3534,N_3739);
and U4251 (N_4251,N_3572,N_3840);
nor U4252 (N_4252,N_3942,N_3720);
nand U4253 (N_4253,N_3825,N_3980);
and U4254 (N_4254,N_3772,N_3681);
xnor U4255 (N_4255,N_3630,N_3565);
xor U4256 (N_4256,N_3898,N_3753);
or U4257 (N_4257,N_3532,N_3895);
or U4258 (N_4258,N_3742,N_3927);
and U4259 (N_4259,N_3746,N_3548);
nor U4260 (N_4260,N_3969,N_3734);
or U4261 (N_4261,N_3945,N_3946);
nand U4262 (N_4262,N_3810,N_3754);
nand U4263 (N_4263,N_3609,N_3958);
or U4264 (N_4264,N_3750,N_3780);
and U4265 (N_4265,N_3884,N_3921);
and U4266 (N_4266,N_3803,N_3983);
or U4267 (N_4267,N_3908,N_3905);
nor U4268 (N_4268,N_3654,N_3709);
nor U4269 (N_4269,N_3924,N_3674);
nor U4270 (N_4270,N_3690,N_3505);
nor U4271 (N_4271,N_3818,N_3695);
or U4272 (N_4272,N_3512,N_3668);
xor U4273 (N_4273,N_3624,N_3965);
nor U4274 (N_4274,N_3541,N_3973);
xnor U4275 (N_4275,N_3694,N_3510);
xnor U4276 (N_4276,N_3546,N_3521);
nand U4277 (N_4277,N_3563,N_3555);
or U4278 (N_4278,N_3693,N_3962);
and U4279 (N_4279,N_3598,N_3522);
xor U4280 (N_4280,N_3632,N_3576);
or U4281 (N_4281,N_3587,N_3990);
or U4282 (N_4282,N_3627,N_3537);
and U4283 (N_4283,N_3773,N_3673);
nor U4284 (N_4284,N_3654,N_3972);
xnor U4285 (N_4285,N_3654,N_3705);
and U4286 (N_4286,N_3959,N_3982);
or U4287 (N_4287,N_3522,N_3567);
xnor U4288 (N_4288,N_3754,N_3582);
nor U4289 (N_4289,N_3957,N_3675);
or U4290 (N_4290,N_3596,N_3746);
nor U4291 (N_4291,N_3900,N_3759);
and U4292 (N_4292,N_3559,N_3647);
nand U4293 (N_4293,N_3692,N_3721);
nor U4294 (N_4294,N_3983,N_3940);
and U4295 (N_4295,N_3962,N_3746);
nand U4296 (N_4296,N_3977,N_3503);
or U4297 (N_4297,N_3667,N_3539);
nand U4298 (N_4298,N_3631,N_3890);
nand U4299 (N_4299,N_3994,N_3515);
nand U4300 (N_4300,N_3910,N_3817);
nand U4301 (N_4301,N_3668,N_3692);
or U4302 (N_4302,N_3600,N_3647);
nand U4303 (N_4303,N_3801,N_3959);
nand U4304 (N_4304,N_3556,N_3913);
and U4305 (N_4305,N_3765,N_3840);
or U4306 (N_4306,N_3643,N_3522);
xnor U4307 (N_4307,N_3513,N_3722);
nor U4308 (N_4308,N_3603,N_3595);
xnor U4309 (N_4309,N_3922,N_3679);
nand U4310 (N_4310,N_3540,N_3876);
xnor U4311 (N_4311,N_3531,N_3687);
xnor U4312 (N_4312,N_3994,N_3885);
xnor U4313 (N_4313,N_3805,N_3651);
xor U4314 (N_4314,N_3734,N_3717);
and U4315 (N_4315,N_3624,N_3544);
xnor U4316 (N_4316,N_3880,N_3567);
xnor U4317 (N_4317,N_3543,N_3738);
and U4318 (N_4318,N_3785,N_3543);
and U4319 (N_4319,N_3632,N_3758);
or U4320 (N_4320,N_3672,N_3756);
nor U4321 (N_4321,N_3560,N_3824);
xnor U4322 (N_4322,N_3540,N_3646);
nor U4323 (N_4323,N_3844,N_3573);
or U4324 (N_4324,N_3828,N_3624);
xnor U4325 (N_4325,N_3878,N_3801);
nor U4326 (N_4326,N_3577,N_3809);
xor U4327 (N_4327,N_3583,N_3530);
or U4328 (N_4328,N_3848,N_3654);
and U4329 (N_4329,N_3807,N_3991);
nor U4330 (N_4330,N_3869,N_3611);
or U4331 (N_4331,N_3646,N_3954);
and U4332 (N_4332,N_3871,N_3919);
nand U4333 (N_4333,N_3841,N_3747);
and U4334 (N_4334,N_3587,N_3693);
nor U4335 (N_4335,N_3526,N_3803);
nand U4336 (N_4336,N_3900,N_3819);
nor U4337 (N_4337,N_3780,N_3806);
and U4338 (N_4338,N_3777,N_3852);
and U4339 (N_4339,N_3841,N_3847);
nand U4340 (N_4340,N_3927,N_3652);
nand U4341 (N_4341,N_3670,N_3604);
nor U4342 (N_4342,N_3566,N_3530);
nor U4343 (N_4343,N_3932,N_3723);
and U4344 (N_4344,N_3834,N_3687);
and U4345 (N_4345,N_3947,N_3591);
nand U4346 (N_4346,N_3717,N_3812);
nand U4347 (N_4347,N_3864,N_3625);
or U4348 (N_4348,N_3599,N_3706);
nand U4349 (N_4349,N_3968,N_3888);
nor U4350 (N_4350,N_3886,N_3707);
and U4351 (N_4351,N_3579,N_3623);
nor U4352 (N_4352,N_3750,N_3617);
nor U4353 (N_4353,N_3688,N_3627);
or U4354 (N_4354,N_3666,N_3566);
xor U4355 (N_4355,N_3565,N_3530);
nand U4356 (N_4356,N_3698,N_3986);
or U4357 (N_4357,N_3652,N_3770);
or U4358 (N_4358,N_3532,N_3923);
nand U4359 (N_4359,N_3865,N_3884);
nand U4360 (N_4360,N_3659,N_3718);
xor U4361 (N_4361,N_3580,N_3959);
or U4362 (N_4362,N_3553,N_3510);
xnor U4363 (N_4363,N_3766,N_3728);
nor U4364 (N_4364,N_3950,N_3762);
xor U4365 (N_4365,N_3706,N_3586);
xor U4366 (N_4366,N_3879,N_3518);
and U4367 (N_4367,N_3989,N_3563);
nor U4368 (N_4368,N_3579,N_3735);
nor U4369 (N_4369,N_3840,N_3668);
nand U4370 (N_4370,N_3913,N_3539);
nor U4371 (N_4371,N_3695,N_3536);
nor U4372 (N_4372,N_3716,N_3525);
and U4373 (N_4373,N_3895,N_3947);
nand U4374 (N_4374,N_3981,N_3909);
nand U4375 (N_4375,N_3537,N_3551);
or U4376 (N_4376,N_3825,N_3783);
nand U4377 (N_4377,N_3650,N_3844);
nand U4378 (N_4378,N_3719,N_3640);
xnor U4379 (N_4379,N_3978,N_3824);
and U4380 (N_4380,N_3884,N_3976);
and U4381 (N_4381,N_3685,N_3640);
and U4382 (N_4382,N_3853,N_3641);
nand U4383 (N_4383,N_3915,N_3796);
or U4384 (N_4384,N_3768,N_3569);
xor U4385 (N_4385,N_3608,N_3700);
xnor U4386 (N_4386,N_3530,N_3883);
nor U4387 (N_4387,N_3528,N_3823);
xnor U4388 (N_4388,N_3857,N_3568);
and U4389 (N_4389,N_3708,N_3976);
or U4390 (N_4390,N_3829,N_3523);
nand U4391 (N_4391,N_3778,N_3518);
nand U4392 (N_4392,N_3911,N_3943);
nor U4393 (N_4393,N_3507,N_3967);
or U4394 (N_4394,N_3632,N_3891);
xor U4395 (N_4395,N_3637,N_3641);
or U4396 (N_4396,N_3744,N_3927);
xor U4397 (N_4397,N_3964,N_3692);
nor U4398 (N_4398,N_3902,N_3604);
nor U4399 (N_4399,N_3967,N_3852);
nor U4400 (N_4400,N_3903,N_3600);
xor U4401 (N_4401,N_3902,N_3850);
nand U4402 (N_4402,N_3811,N_3972);
and U4403 (N_4403,N_3662,N_3836);
nor U4404 (N_4404,N_3548,N_3917);
and U4405 (N_4405,N_3868,N_3692);
xor U4406 (N_4406,N_3609,N_3550);
nand U4407 (N_4407,N_3947,N_3788);
nor U4408 (N_4408,N_3923,N_3982);
nand U4409 (N_4409,N_3658,N_3927);
nand U4410 (N_4410,N_3665,N_3585);
nor U4411 (N_4411,N_3777,N_3590);
or U4412 (N_4412,N_3735,N_3890);
or U4413 (N_4413,N_3937,N_3951);
nand U4414 (N_4414,N_3914,N_3849);
or U4415 (N_4415,N_3550,N_3954);
nor U4416 (N_4416,N_3704,N_3655);
nand U4417 (N_4417,N_3612,N_3927);
and U4418 (N_4418,N_3839,N_3788);
or U4419 (N_4419,N_3652,N_3904);
and U4420 (N_4420,N_3797,N_3636);
xor U4421 (N_4421,N_3823,N_3550);
or U4422 (N_4422,N_3817,N_3842);
nand U4423 (N_4423,N_3926,N_3680);
xor U4424 (N_4424,N_3681,N_3830);
nand U4425 (N_4425,N_3830,N_3608);
and U4426 (N_4426,N_3758,N_3685);
or U4427 (N_4427,N_3821,N_3718);
or U4428 (N_4428,N_3981,N_3570);
or U4429 (N_4429,N_3505,N_3969);
and U4430 (N_4430,N_3660,N_3848);
nand U4431 (N_4431,N_3666,N_3860);
nor U4432 (N_4432,N_3805,N_3616);
nor U4433 (N_4433,N_3996,N_3807);
xnor U4434 (N_4434,N_3896,N_3690);
xor U4435 (N_4435,N_3659,N_3723);
xnor U4436 (N_4436,N_3608,N_3857);
nand U4437 (N_4437,N_3550,N_3788);
and U4438 (N_4438,N_3845,N_3637);
nor U4439 (N_4439,N_3577,N_3945);
and U4440 (N_4440,N_3780,N_3640);
and U4441 (N_4441,N_3621,N_3605);
and U4442 (N_4442,N_3936,N_3741);
and U4443 (N_4443,N_3745,N_3605);
or U4444 (N_4444,N_3801,N_3955);
and U4445 (N_4445,N_3584,N_3985);
and U4446 (N_4446,N_3894,N_3560);
nor U4447 (N_4447,N_3838,N_3628);
nor U4448 (N_4448,N_3966,N_3520);
nor U4449 (N_4449,N_3916,N_3726);
and U4450 (N_4450,N_3638,N_3906);
or U4451 (N_4451,N_3572,N_3836);
or U4452 (N_4452,N_3549,N_3868);
and U4453 (N_4453,N_3876,N_3776);
xor U4454 (N_4454,N_3584,N_3748);
xor U4455 (N_4455,N_3994,N_3523);
nand U4456 (N_4456,N_3838,N_3553);
nand U4457 (N_4457,N_3528,N_3879);
or U4458 (N_4458,N_3996,N_3916);
xor U4459 (N_4459,N_3614,N_3881);
xor U4460 (N_4460,N_3969,N_3943);
xnor U4461 (N_4461,N_3792,N_3790);
or U4462 (N_4462,N_3533,N_3516);
xnor U4463 (N_4463,N_3668,N_3927);
or U4464 (N_4464,N_3747,N_3938);
nor U4465 (N_4465,N_3981,N_3859);
nand U4466 (N_4466,N_3887,N_3981);
or U4467 (N_4467,N_3584,N_3954);
and U4468 (N_4468,N_3965,N_3581);
xnor U4469 (N_4469,N_3708,N_3726);
xnor U4470 (N_4470,N_3501,N_3689);
and U4471 (N_4471,N_3535,N_3770);
xnor U4472 (N_4472,N_3758,N_3907);
and U4473 (N_4473,N_3776,N_3903);
nor U4474 (N_4474,N_3857,N_3814);
nor U4475 (N_4475,N_3746,N_3792);
nor U4476 (N_4476,N_3783,N_3633);
or U4477 (N_4477,N_3663,N_3683);
or U4478 (N_4478,N_3972,N_3640);
or U4479 (N_4479,N_3847,N_3901);
and U4480 (N_4480,N_3628,N_3570);
nand U4481 (N_4481,N_3991,N_3871);
nor U4482 (N_4482,N_3541,N_3854);
and U4483 (N_4483,N_3855,N_3779);
or U4484 (N_4484,N_3769,N_3834);
nand U4485 (N_4485,N_3918,N_3534);
or U4486 (N_4486,N_3635,N_3590);
nor U4487 (N_4487,N_3696,N_3851);
nand U4488 (N_4488,N_3924,N_3734);
nand U4489 (N_4489,N_3537,N_3658);
xnor U4490 (N_4490,N_3742,N_3884);
and U4491 (N_4491,N_3638,N_3787);
nor U4492 (N_4492,N_3601,N_3646);
xor U4493 (N_4493,N_3854,N_3814);
nand U4494 (N_4494,N_3995,N_3565);
or U4495 (N_4495,N_3594,N_3789);
nor U4496 (N_4496,N_3904,N_3917);
nand U4497 (N_4497,N_3982,N_3619);
nand U4498 (N_4498,N_3825,N_3934);
nand U4499 (N_4499,N_3763,N_3811);
nand U4500 (N_4500,N_4206,N_4311);
xor U4501 (N_4501,N_4025,N_4297);
xor U4502 (N_4502,N_4201,N_4034);
xor U4503 (N_4503,N_4290,N_4392);
and U4504 (N_4504,N_4427,N_4074);
xor U4505 (N_4505,N_4177,N_4055);
or U4506 (N_4506,N_4469,N_4394);
nor U4507 (N_4507,N_4040,N_4416);
nand U4508 (N_4508,N_4438,N_4411);
nor U4509 (N_4509,N_4205,N_4355);
or U4510 (N_4510,N_4393,N_4423);
or U4511 (N_4511,N_4227,N_4428);
xor U4512 (N_4512,N_4185,N_4245);
nor U4513 (N_4513,N_4009,N_4093);
xor U4514 (N_4514,N_4207,N_4140);
nor U4515 (N_4515,N_4117,N_4197);
or U4516 (N_4516,N_4084,N_4404);
or U4517 (N_4517,N_4159,N_4129);
nand U4518 (N_4518,N_4370,N_4286);
nor U4519 (N_4519,N_4489,N_4044);
nand U4520 (N_4520,N_4014,N_4249);
nand U4521 (N_4521,N_4080,N_4193);
xor U4522 (N_4522,N_4000,N_4007);
nor U4523 (N_4523,N_4301,N_4315);
and U4524 (N_4524,N_4320,N_4062);
nand U4525 (N_4525,N_4110,N_4484);
nor U4526 (N_4526,N_4285,N_4189);
or U4527 (N_4527,N_4351,N_4352);
xor U4528 (N_4528,N_4406,N_4401);
xnor U4529 (N_4529,N_4194,N_4109);
nand U4530 (N_4530,N_4032,N_4130);
xor U4531 (N_4531,N_4065,N_4420);
nand U4532 (N_4532,N_4190,N_4115);
nand U4533 (N_4533,N_4001,N_4457);
and U4534 (N_4534,N_4440,N_4322);
or U4535 (N_4535,N_4144,N_4386);
and U4536 (N_4536,N_4168,N_4476);
or U4537 (N_4537,N_4186,N_4292);
xnor U4538 (N_4538,N_4271,N_4273);
xnor U4539 (N_4539,N_4403,N_4373);
nor U4540 (N_4540,N_4031,N_4090);
or U4541 (N_4541,N_4374,N_4380);
xnor U4542 (N_4542,N_4119,N_4121);
nor U4543 (N_4543,N_4410,N_4118);
nand U4544 (N_4544,N_4365,N_4470);
or U4545 (N_4545,N_4296,N_4236);
nor U4546 (N_4546,N_4181,N_4396);
and U4547 (N_4547,N_4255,N_4033);
nor U4548 (N_4548,N_4157,N_4221);
and U4549 (N_4549,N_4172,N_4147);
nand U4550 (N_4550,N_4037,N_4268);
nand U4551 (N_4551,N_4053,N_4468);
nand U4552 (N_4552,N_4314,N_4218);
nand U4553 (N_4553,N_4072,N_4424);
or U4554 (N_4554,N_4112,N_4123);
xor U4555 (N_4555,N_4283,N_4008);
nor U4556 (N_4556,N_4316,N_4223);
or U4557 (N_4557,N_4158,N_4455);
and U4558 (N_4558,N_4305,N_4284);
and U4559 (N_4559,N_4332,N_4407);
nand U4560 (N_4560,N_4170,N_4444);
xor U4561 (N_4561,N_4054,N_4421);
and U4562 (N_4562,N_4230,N_4310);
and U4563 (N_4563,N_4319,N_4293);
nor U4564 (N_4564,N_4472,N_4242);
nor U4565 (N_4565,N_4134,N_4291);
or U4566 (N_4566,N_4264,N_4002);
nand U4567 (N_4567,N_4244,N_4340);
or U4568 (N_4568,N_4057,N_4487);
or U4569 (N_4569,N_4272,N_4141);
nand U4570 (N_4570,N_4097,N_4228);
nor U4571 (N_4571,N_4388,N_4349);
or U4572 (N_4572,N_4362,N_4318);
or U4573 (N_4573,N_4453,N_4067);
nor U4574 (N_4574,N_4267,N_4356);
xnor U4575 (N_4575,N_4371,N_4131);
or U4576 (N_4576,N_4111,N_4073);
or U4577 (N_4577,N_4212,N_4474);
or U4578 (N_4578,N_4486,N_4382);
xnor U4579 (N_4579,N_4248,N_4341);
xnor U4580 (N_4580,N_4338,N_4217);
nor U4581 (N_4581,N_4116,N_4413);
and U4582 (N_4582,N_4385,N_4437);
nor U4583 (N_4583,N_4400,N_4451);
or U4584 (N_4584,N_4304,N_4497);
nor U4585 (N_4585,N_4298,N_4443);
or U4586 (N_4586,N_4475,N_4160);
nand U4587 (N_4587,N_4069,N_4075);
nor U4588 (N_4588,N_4050,N_4191);
xnor U4589 (N_4589,N_4381,N_4259);
nand U4590 (N_4590,N_4082,N_4279);
nand U4591 (N_4591,N_4155,N_4094);
or U4592 (N_4592,N_4435,N_4375);
xnor U4593 (N_4593,N_4330,N_4017);
xor U4594 (N_4594,N_4089,N_4496);
and U4595 (N_4595,N_4402,N_4132);
and U4596 (N_4596,N_4239,N_4376);
nor U4597 (N_4597,N_4466,N_4418);
xnor U4598 (N_4598,N_4195,N_4460);
nand U4599 (N_4599,N_4026,N_4036);
and U4600 (N_4600,N_4083,N_4148);
nand U4601 (N_4601,N_4462,N_4389);
and U4602 (N_4602,N_4164,N_4397);
xor U4603 (N_4603,N_4240,N_4463);
xnor U4604 (N_4604,N_4204,N_4103);
and U4605 (N_4605,N_4346,N_4041);
or U4606 (N_4606,N_4019,N_4419);
or U4607 (N_4607,N_4137,N_4081);
nand U4608 (N_4608,N_4149,N_4350);
xnor U4609 (N_4609,N_4233,N_4495);
xnor U4610 (N_4610,N_4479,N_4237);
or U4611 (N_4611,N_4088,N_4347);
xor U4612 (N_4612,N_4313,N_4027);
xor U4613 (N_4613,N_4369,N_4180);
or U4614 (N_4614,N_4384,N_4282);
xnor U4615 (N_4615,N_4358,N_4323);
nor U4616 (N_4616,N_4395,N_4260);
or U4617 (N_4617,N_4243,N_4254);
and U4618 (N_4618,N_4183,N_4077);
xor U4619 (N_4619,N_4096,N_4224);
and U4620 (N_4620,N_4056,N_4359);
and U4621 (N_4621,N_4169,N_4482);
nor U4622 (N_4622,N_4167,N_4448);
and U4623 (N_4623,N_4429,N_4481);
and U4624 (N_4624,N_4126,N_4478);
xor U4625 (N_4625,N_4042,N_4222);
or U4626 (N_4626,N_4079,N_4361);
xor U4627 (N_4627,N_4415,N_4030);
and U4628 (N_4628,N_4447,N_4176);
nand U4629 (N_4629,N_4277,N_4235);
or U4630 (N_4630,N_4215,N_4187);
nor U4631 (N_4631,N_4171,N_4348);
and U4632 (N_4632,N_4208,N_4266);
and U4633 (N_4633,N_4039,N_4265);
or U4634 (N_4634,N_4490,N_4152);
or U4635 (N_4635,N_4049,N_4087);
nor U4636 (N_4636,N_4269,N_4299);
nand U4637 (N_4637,N_4471,N_4275);
and U4638 (N_4638,N_4258,N_4029);
nand U4639 (N_4639,N_4433,N_4199);
nor U4640 (N_4640,N_4353,N_4021);
nor U4641 (N_4641,N_4485,N_4477);
xnor U4642 (N_4642,N_4335,N_4366);
or U4643 (N_4643,N_4331,N_4108);
nand U4644 (N_4644,N_4231,N_4494);
nand U4645 (N_4645,N_4306,N_4071);
xnor U4646 (N_4646,N_4390,N_4328);
and U4647 (N_4647,N_4178,N_4015);
or U4648 (N_4648,N_4483,N_4309);
and U4649 (N_4649,N_4043,N_4379);
and U4650 (N_4650,N_4124,N_4122);
and U4651 (N_4651,N_4302,N_4220);
or U4652 (N_4652,N_4128,N_4325);
and U4653 (N_4653,N_4434,N_4442);
nor U4654 (N_4654,N_4498,N_4016);
xor U4655 (N_4655,N_4229,N_4143);
nor U4656 (N_4656,N_4010,N_4289);
or U4657 (N_4657,N_4326,N_4038);
nor U4658 (N_4658,N_4102,N_4464);
or U4659 (N_4659,N_4196,N_4127);
and U4660 (N_4660,N_4426,N_4114);
or U4661 (N_4661,N_4458,N_4307);
nor U4662 (N_4662,N_4336,N_4216);
or U4663 (N_4663,N_4162,N_4414);
nand U4664 (N_4664,N_4099,N_4364);
or U4665 (N_4665,N_4070,N_4321);
nand U4666 (N_4666,N_4329,N_4105);
or U4667 (N_4667,N_4076,N_4261);
nand U4668 (N_4668,N_4408,N_4461);
xor U4669 (N_4669,N_4104,N_4120);
and U4670 (N_4670,N_4163,N_4154);
xnor U4671 (N_4671,N_4003,N_4086);
nor U4672 (N_4672,N_4023,N_4250);
or U4673 (N_4673,N_4312,N_4013);
nand U4674 (N_4674,N_4368,N_4439);
nor U4675 (N_4675,N_4022,N_4387);
nand U4676 (N_4676,N_4430,N_4198);
and U4677 (N_4677,N_4150,N_4247);
nor U4678 (N_4678,N_4095,N_4467);
and U4679 (N_4679,N_4136,N_4064);
and U4680 (N_4680,N_4334,N_4241);
and U4681 (N_4681,N_4146,N_4139);
and U4682 (N_4682,N_4287,N_4135);
and U4683 (N_4683,N_4012,N_4151);
nand U4684 (N_4684,N_4454,N_4270);
and U4685 (N_4685,N_4342,N_4179);
nor U4686 (N_4686,N_4142,N_4226);
and U4687 (N_4687,N_4417,N_4354);
xor U4688 (N_4688,N_4333,N_4047);
nand U4689 (N_4689,N_4278,N_4133);
nor U4690 (N_4690,N_4232,N_4465);
xor U4691 (N_4691,N_4492,N_4399);
and U4692 (N_4692,N_4246,N_4068);
nand U4693 (N_4693,N_4078,N_4166);
nand U4694 (N_4694,N_4035,N_4446);
and U4695 (N_4695,N_4138,N_4225);
xnor U4696 (N_4696,N_4422,N_4409);
or U4697 (N_4697,N_4209,N_4098);
or U4698 (N_4698,N_4028,N_4175);
or U4699 (N_4699,N_4101,N_4405);
or U4700 (N_4700,N_4445,N_4165);
nor U4701 (N_4701,N_4257,N_4006);
nand U4702 (N_4702,N_4276,N_4288);
and U4703 (N_4703,N_4372,N_4436);
or U4704 (N_4704,N_4377,N_4048);
and U4705 (N_4705,N_4046,N_4024);
or U4706 (N_4706,N_4383,N_4262);
xor U4707 (N_4707,N_4052,N_4161);
or U4708 (N_4708,N_4219,N_4234);
or U4709 (N_4709,N_4188,N_4210);
nor U4710 (N_4710,N_4339,N_4263);
or U4711 (N_4711,N_4345,N_4203);
or U4712 (N_4712,N_4303,N_4274);
nand U4713 (N_4713,N_4480,N_4238);
and U4714 (N_4714,N_4107,N_4153);
xnor U4715 (N_4715,N_4450,N_4060);
xnor U4716 (N_4716,N_4398,N_4174);
nor U4717 (N_4717,N_4327,N_4294);
nand U4718 (N_4718,N_4211,N_4378);
or U4719 (N_4719,N_4360,N_4051);
xor U4720 (N_4720,N_4091,N_4192);
or U4721 (N_4721,N_4058,N_4251);
or U4722 (N_4722,N_4425,N_4308);
xor U4723 (N_4723,N_4182,N_4066);
nand U4724 (N_4724,N_4200,N_4317);
or U4725 (N_4725,N_4367,N_4061);
and U4726 (N_4726,N_4045,N_4125);
and U4727 (N_4727,N_4473,N_4202);
and U4728 (N_4728,N_4281,N_4391);
and U4729 (N_4729,N_4412,N_4213);
nand U4730 (N_4730,N_4113,N_4488);
nor U4731 (N_4731,N_4092,N_4337);
or U4732 (N_4732,N_4432,N_4085);
nand U4733 (N_4733,N_4173,N_4491);
nand U4734 (N_4734,N_4295,N_4106);
nor U4735 (N_4735,N_4018,N_4005);
nor U4736 (N_4736,N_4253,N_4459);
xnor U4737 (N_4737,N_4004,N_4456);
nand U4738 (N_4738,N_4063,N_4252);
nand U4739 (N_4739,N_4441,N_4363);
nor U4740 (N_4740,N_4452,N_4256);
and U4741 (N_4741,N_4156,N_4214);
nor U4742 (N_4742,N_4184,N_4449);
xor U4743 (N_4743,N_4493,N_4011);
or U4744 (N_4744,N_4145,N_4020);
and U4745 (N_4745,N_4280,N_4324);
nor U4746 (N_4746,N_4344,N_4499);
nor U4747 (N_4747,N_4431,N_4343);
or U4748 (N_4748,N_4357,N_4100);
and U4749 (N_4749,N_4300,N_4059);
nor U4750 (N_4750,N_4414,N_4376);
and U4751 (N_4751,N_4377,N_4067);
or U4752 (N_4752,N_4305,N_4270);
xor U4753 (N_4753,N_4105,N_4183);
and U4754 (N_4754,N_4244,N_4481);
xor U4755 (N_4755,N_4396,N_4262);
nand U4756 (N_4756,N_4352,N_4251);
nand U4757 (N_4757,N_4000,N_4034);
and U4758 (N_4758,N_4069,N_4256);
xor U4759 (N_4759,N_4209,N_4438);
nor U4760 (N_4760,N_4042,N_4285);
or U4761 (N_4761,N_4112,N_4295);
or U4762 (N_4762,N_4093,N_4151);
nand U4763 (N_4763,N_4025,N_4362);
xor U4764 (N_4764,N_4180,N_4186);
nor U4765 (N_4765,N_4410,N_4290);
nor U4766 (N_4766,N_4148,N_4486);
nand U4767 (N_4767,N_4387,N_4098);
nor U4768 (N_4768,N_4178,N_4249);
or U4769 (N_4769,N_4445,N_4248);
or U4770 (N_4770,N_4079,N_4411);
and U4771 (N_4771,N_4497,N_4265);
xnor U4772 (N_4772,N_4189,N_4086);
nor U4773 (N_4773,N_4072,N_4162);
or U4774 (N_4774,N_4089,N_4362);
xor U4775 (N_4775,N_4291,N_4314);
and U4776 (N_4776,N_4271,N_4399);
and U4777 (N_4777,N_4299,N_4458);
nor U4778 (N_4778,N_4200,N_4316);
nor U4779 (N_4779,N_4251,N_4407);
xor U4780 (N_4780,N_4128,N_4184);
nor U4781 (N_4781,N_4436,N_4049);
xnor U4782 (N_4782,N_4234,N_4175);
nand U4783 (N_4783,N_4376,N_4407);
or U4784 (N_4784,N_4206,N_4293);
nor U4785 (N_4785,N_4349,N_4283);
nor U4786 (N_4786,N_4461,N_4401);
and U4787 (N_4787,N_4260,N_4495);
nand U4788 (N_4788,N_4097,N_4431);
nand U4789 (N_4789,N_4336,N_4023);
or U4790 (N_4790,N_4294,N_4012);
nor U4791 (N_4791,N_4450,N_4071);
or U4792 (N_4792,N_4180,N_4049);
and U4793 (N_4793,N_4081,N_4286);
nand U4794 (N_4794,N_4054,N_4303);
or U4795 (N_4795,N_4432,N_4252);
or U4796 (N_4796,N_4223,N_4329);
nand U4797 (N_4797,N_4055,N_4381);
nor U4798 (N_4798,N_4329,N_4046);
and U4799 (N_4799,N_4144,N_4165);
or U4800 (N_4800,N_4392,N_4210);
and U4801 (N_4801,N_4453,N_4492);
or U4802 (N_4802,N_4114,N_4063);
nor U4803 (N_4803,N_4375,N_4095);
nor U4804 (N_4804,N_4316,N_4314);
xor U4805 (N_4805,N_4144,N_4471);
and U4806 (N_4806,N_4096,N_4044);
nor U4807 (N_4807,N_4304,N_4465);
and U4808 (N_4808,N_4282,N_4375);
or U4809 (N_4809,N_4179,N_4287);
xnor U4810 (N_4810,N_4464,N_4404);
nor U4811 (N_4811,N_4067,N_4491);
and U4812 (N_4812,N_4483,N_4256);
nand U4813 (N_4813,N_4049,N_4332);
and U4814 (N_4814,N_4242,N_4473);
and U4815 (N_4815,N_4419,N_4259);
nand U4816 (N_4816,N_4210,N_4218);
nand U4817 (N_4817,N_4405,N_4099);
nand U4818 (N_4818,N_4358,N_4217);
xor U4819 (N_4819,N_4238,N_4112);
or U4820 (N_4820,N_4357,N_4279);
or U4821 (N_4821,N_4479,N_4151);
and U4822 (N_4822,N_4380,N_4289);
nor U4823 (N_4823,N_4005,N_4305);
or U4824 (N_4824,N_4322,N_4459);
or U4825 (N_4825,N_4262,N_4264);
nand U4826 (N_4826,N_4236,N_4095);
nor U4827 (N_4827,N_4117,N_4121);
nand U4828 (N_4828,N_4482,N_4272);
and U4829 (N_4829,N_4098,N_4240);
nor U4830 (N_4830,N_4292,N_4473);
nor U4831 (N_4831,N_4097,N_4497);
xor U4832 (N_4832,N_4473,N_4305);
xnor U4833 (N_4833,N_4019,N_4068);
nand U4834 (N_4834,N_4262,N_4041);
and U4835 (N_4835,N_4042,N_4129);
and U4836 (N_4836,N_4174,N_4486);
nand U4837 (N_4837,N_4207,N_4136);
xnor U4838 (N_4838,N_4297,N_4329);
nand U4839 (N_4839,N_4387,N_4149);
xor U4840 (N_4840,N_4492,N_4056);
and U4841 (N_4841,N_4160,N_4422);
xor U4842 (N_4842,N_4076,N_4332);
nor U4843 (N_4843,N_4149,N_4245);
or U4844 (N_4844,N_4123,N_4404);
and U4845 (N_4845,N_4112,N_4376);
xor U4846 (N_4846,N_4148,N_4299);
nor U4847 (N_4847,N_4457,N_4422);
and U4848 (N_4848,N_4275,N_4031);
nand U4849 (N_4849,N_4413,N_4149);
nand U4850 (N_4850,N_4467,N_4193);
xnor U4851 (N_4851,N_4174,N_4149);
nand U4852 (N_4852,N_4146,N_4149);
or U4853 (N_4853,N_4213,N_4095);
and U4854 (N_4854,N_4456,N_4231);
or U4855 (N_4855,N_4076,N_4172);
and U4856 (N_4856,N_4149,N_4071);
nand U4857 (N_4857,N_4388,N_4371);
nor U4858 (N_4858,N_4395,N_4134);
xor U4859 (N_4859,N_4399,N_4182);
xor U4860 (N_4860,N_4094,N_4153);
or U4861 (N_4861,N_4157,N_4047);
nor U4862 (N_4862,N_4290,N_4243);
or U4863 (N_4863,N_4383,N_4210);
or U4864 (N_4864,N_4091,N_4198);
nand U4865 (N_4865,N_4147,N_4491);
nor U4866 (N_4866,N_4316,N_4252);
nor U4867 (N_4867,N_4285,N_4171);
and U4868 (N_4868,N_4128,N_4236);
xor U4869 (N_4869,N_4123,N_4129);
or U4870 (N_4870,N_4163,N_4221);
xnor U4871 (N_4871,N_4307,N_4424);
and U4872 (N_4872,N_4231,N_4018);
and U4873 (N_4873,N_4354,N_4094);
nand U4874 (N_4874,N_4260,N_4194);
nand U4875 (N_4875,N_4230,N_4218);
xor U4876 (N_4876,N_4421,N_4401);
or U4877 (N_4877,N_4305,N_4237);
nand U4878 (N_4878,N_4055,N_4002);
nor U4879 (N_4879,N_4088,N_4099);
and U4880 (N_4880,N_4245,N_4000);
nand U4881 (N_4881,N_4196,N_4274);
or U4882 (N_4882,N_4321,N_4088);
xnor U4883 (N_4883,N_4411,N_4366);
nand U4884 (N_4884,N_4176,N_4170);
and U4885 (N_4885,N_4137,N_4285);
and U4886 (N_4886,N_4490,N_4397);
nand U4887 (N_4887,N_4490,N_4479);
and U4888 (N_4888,N_4246,N_4242);
nor U4889 (N_4889,N_4397,N_4387);
nor U4890 (N_4890,N_4336,N_4159);
nor U4891 (N_4891,N_4128,N_4147);
xor U4892 (N_4892,N_4012,N_4382);
xor U4893 (N_4893,N_4476,N_4384);
and U4894 (N_4894,N_4019,N_4290);
nor U4895 (N_4895,N_4222,N_4301);
or U4896 (N_4896,N_4448,N_4278);
nand U4897 (N_4897,N_4420,N_4032);
nand U4898 (N_4898,N_4026,N_4310);
nor U4899 (N_4899,N_4028,N_4254);
nor U4900 (N_4900,N_4276,N_4024);
and U4901 (N_4901,N_4252,N_4352);
nor U4902 (N_4902,N_4245,N_4206);
and U4903 (N_4903,N_4120,N_4360);
nand U4904 (N_4904,N_4483,N_4394);
or U4905 (N_4905,N_4301,N_4297);
nand U4906 (N_4906,N_4421,N_4470);
or U4907 (N_4907,N_4166,N_4377);
nand U4908 (N_4908,N_4213,N_4200);
or U4909 (N_4909,N_4046,N_4461);
nor U4910 (N_4910,N_4140,N_4467);
and U4911 (N_4911,N_4087,N_4419);
xnor U4912 (N_4912,N_4266,N_4016);
or U4913 (N_4913,N_4118,N_4027);
nor U4914 (N_4914,N_4212,N_4052);
or U4915 (N_4915,N_4249,N_4162);
or U4916 (N_4916,N_4252,N_4187);
xnor U4917 (N_4917,N_4272,N_4475);
and U4918 (N_4918,N_4377,N_4007);
nand U4919 (N_4919,N_4354,N_4038);
and U4920 (N_4920,N_4348,N_4141);
xor U4921 (N_4921,N_4280,N_4495);
and U4922 (N_4922,N_4446,N_4484);
and U4923 (N_4923,N_4202,N_4199);
nand U4924 (N_4924,N_4171,N_4318);
nand U4925 (N_4925,N_4097,N_4381);
and U4926 (N_4926,N_4329,N_4109);
and U4927 (N_4927,N_4063,N_4486);
or U4928 (N_4928,N_4421,N_4392);
nand U4929 (N_4929,N_4355,N_4351);
nand U4930 (N_4930,N_4450,N_4030);
and U4931 (N_4931,N_4103,N_4047);
nor U4932 (N_4932,N_4469,N_4497);
nand U4933 (N_4933,N_4076,N_4377);
nand U4934 (N_4934,N_4421,N_4053);
nand U4935 (N_4935,N_4488,N_4331);
nand U4936 (N_4936,N_4368,N_4396);
or U4937 (N_4937,N_4411,N_4254);
nand U4938 (N_4938,N_4384,N_4071);
and U4939 (N_4939,N_4311,N_4167);
and U4940 (N_4940,N_4449,N_4432);
nor U4941 (N_4941,N_4490,N_4327);
nand U4942 (N_4942,N_4491,N_4361);
or U4943 (N_4943,N_4425,N_4104);
and U4944 (N_4944,N_4119,N_4083);
xor U4945 (N_4945,N_4145,N_4392);
nor U4946 (N_4946,N_4286,N_4496);
nor U4947 (N_4947,N_4118,N_4222);
or U4948 (N_4948,N_4259,N_4149);
nand U4949 (N_4949,N_4413,N_4201);
or U4950 (N_4950,N_4063,N_4324);
and U4951 (N_4951,N_4425,N_4435);
nor U4952 (N_4952,N_4495,N_4196);
nand U4953 (N_4953,N_4080,N_4417);
or U4954 (N_4954,N_4153,N_4264);
nand U4955 (N_4955,N_4466,N_4320);
nand U4956 (N_4956,N_4330,N_4295);
or U4957 (N_4957,N_4211,N_4109);
nand U4958 (N_4958,N_4352,N_4460);
or U4959 (N_4959,N_4399,N_4125);
xor U4960 (N_4960,N_4022,N_4165);
or U4961 (N_4961,N_4169,N_4019);
nand U4962 (N_4962,N_4035,N_4023);
nand U4963 (N_4963,N_4023,N_4332);
or U4964 (N_4964,N_4264,N_4232);
nand U4965 (N_4965,N_4440,N_4244);
or U4966 (N_4966,N_4079,N_4106);
or U4967 (N_4967,N_4207,N_4355);
and U4968 (N_4968,N_4070,N_4271);
nor U4969 (N_4969,N_4323,N_4256);
xor U4970 (N_4970,N_4433,N_4136);
or U4971 (N_4971,N_4485,N_4062);
nor U4972 (N_4972,N_4024,N_4446);
or U4973 (N_4973,N_4451,N_4463);
or U4974 (N_4974,N_4089,N_4069);
or U4975 (N_4975,N_4177,N_4371);
nand U4976 (N_4976,N_4246,N_4338);
nand U4977 (N_4977,N_4028,N_4067);
nor U4978 (N_4978,N_4285,N_4227);
nand U4979 (N_4979,N_4255,N_4053);
xor U4980 (N_4980,N_4221,N_4490);
and U4981 (N_4981,N_4097,N_4180);
nand U4982 (N_4982,N_4122,N_4440);
and U4983 (N_4983,N_4007,N_4117);
nor U4984 (N_4984,N_4263,N_4304);
and U4985 (N_4985,N_4243,N_4375);
or U4986 (N_4986,N_4287,N_4447);
and U4987 (N_4987,N_4033,N_4312);
or U4988 (N_4988,N_4489,N_4046);
or U4989 (N_4989,N_4090,N_4378);
nand U4990 (N_4990,N_4259,N_4216);
nand U4991 (N_4991,N_4471,N_4065);
or U4992 (N_4992,N_4493,N_4415);
xor U4993 (N_4993,N_4033,N_4390);
and U4994 (N_4994,N_4333,N_4304);
and U4995 (N_4995,N_4395,N_4184);
nor U4996 (N_4996,N_4222,N_4048);
nand U4997 (N_4997,N_4004,N_4020);
and U4998 (N_4998,N_4222,N_4408);
nor U4999 (N_4999,N_4302,N_4154);
or U5000 (N_5000,N_4611,N_4753);
xnor U5001 (N_5001,N_4746,N_4555);
nand U5002 (N_5002,N_4520,N_4735);
nand U5003 (N_5003,N_4872,N_4624);
xor U5004 (N_5004,N_4894,N_4732);
xnor U5005 (N_5005,N_4629,N_4862);
and U5006 (N_5006,N_4821,N_4642);
or U5007 (N_5007,N_4846,N_4960);
xnor U5008 (N_5008,N_4524,N_4516);
nor U5009 (N_5009,N_4562,N_4793);
xor U5010 (N_5010,N_4582,N_4911);
or U5011 (N_5011,N_4980,N_4822);
or U5012 (N_5012,N_4815,N_4655);
or U5013 (N_5013,N_4670,N_4640);
nand U5014 (N_5014,N_4630,N_4552);
and U5015 (N_5015,N_4754,N_4908);
nand U5016 (N_5016,N_4579,N_4829);
nand U5017 (N_5017,N_4853,N_4868);
nor U5018 (N_5018,N_4887,N_4828);
and U5019 (N_5019,N_4729,N_4540);
nand U5020 (N_5020,N_4507,N_4599);
or U5021 (N_5021,N_4519,N_4880);
nand U5022 (N_5022,N_4944,N_4914);
xor U5023 (N_5023,N_4530,N_4699);
and U5024 (N_5024,N_4509,N_4781);
and U5025 (N_5025,N_4733,N_4533);
xnor U5026 (N_5026,N_4590,N_4865);
and U5027 (N_5027,N_4875,N_4920);
and U5028 (N_5028,N_4989,N_4964);
xor U5029 (N_5029,N_4788,N_4730);
xor U5030 (N_5030,N_4956,N_4628);
or U5031 (N_5031,N_4852,N_4531);
nand U5032 (N_5032,N_4907,N_4610);
and U5033 (N_5033,N_4656,N_4679);
and U5034 (N_5034,N_4843,N_4882);
xnor U5035 (N_5035,N_4817,N_4915);
or U5036 (N_5036,N_4896,N_4928);
or U5037 (N_5037,N_4921,N_4502);
and U5038 (N_5038,N_4615,N_4917);
xnor U5039 (N_5039,N_4778,N_4687);
and U5040 (N_5040,N_4986,N_4612);
or U5041 (N_5041,N_4803,N_4764);
or U5042 (N_5042,N_4892,N_4663);
and U5043 (N_5043,N_4751,N_4525);
nor U5044 (N_5044,N_4654,N_4870);
and U5045 (N_5045,N_4691,N_4818);
nand U5046 (N_5046,N_4607,N_4571);
xnor U5047 (N_5047,N_4762,N_4769);
nor U5048 (N_5048,N_4805,N_4845);
nor U5049 (N_5049,N_4643,N_4800);
or U5050 (N_5050,N_4697,N_4926);
xor U5051 (N_5051,N_4913,N_4665);
xnor U5052 (N_5052,N_4613,N_4835);
and U5053 (N_5053,N_4877,N_4849);
nand U5054 (N_5054,N_4939,N_4726);
nand U5055 (N_5055,N_4690,N_4526);
nor U5056 (N_5056,N_4522,N_4711);
nor U5057 (N_5057,N_4988,N_4709);
nand U5058 (N_5058,N_4949,N_4997);
nand U5059 (N_5059,N_4736,N_4708);
xnor U5060 (N_5060,N_4837,N_4604);
and U5061 (N_5061,N_4694,N_4824);
and U5062 (N_5062,N_4632,N_4873);
and U5063 (N_5063,N_4572,N_4798);
nor U5064 (N_5064,N_4922,N_4995);
and U5065 (N_5065,N_4750,N_4504);
nor U5066 (N_5066,N_4692,N_4741);
or U5067 (N_5067,N_4623,N_4614);
or U5068 (N_5068,N_4527,N_4796);
or U5069 (N_5069,N_4731,N_4958);
xor U5070 (N_5070,N_4678,N_4659);
xnor U5071 (N_5071,N_4569,N_4681);
and U5072 (N_5072,N_4923,N_4660);
xor U5073 (N_5073,N_4787,N_4722);
and U5074 (N_5074,N_4963,N_4547);
xnor U5075 (N_5075,N_4541,N_4752);
or U5076 (N_5076,N_4653,N_4685);
xor U5077 (N_5077,N_4667,N_4780);
or U5078 (N_5078,N_4639,N_4727);
nand U5079 (N_5079,N_4885,N_4534);
nor U5080 (N_5080,N_4968,N_4724);
nand U5081 (N_5081,N_4957,N_4702);
nor U5082 (N_5082,N_4951,N_4761);
nor U5083 (N_5083,N_4638,N_4646);
nand U5084 (N_5084,N_4884,N_4991);
nor U5085 (N_5085,N_4973,N_4714);
nor U5086 (N_5086,N_4940,N_4734);
nor U5087 (N_5087,N_4603,N_4595);
nor U5088 (N_5088,N_4901,N_4856);
xnor U5089 (N_5089,N_4587,N_4617);
nand U5090 (N_5090,N_4712,N_4927);
and U5091 (N_5091,N_4889,N_4556);
or U5092 (N_5092,N_4943,N_4860);
xnor U5093 (N_5093,N_4893,N_4797);
and U5094 (N_5094,N_4857,N_4992);
and U5095 (N_5095,N_4826,N_4647);
xnor U5096 (N_5096,N_4506,N_4693);
or U5097 (N_5097,N_4704,N_4905);
xnor U5098 (N_5098,N_4810,N_4602);
or U5099 (N_5099,N_4718,N_4777);
nand U5100 (N_5100,N_4563,N_4941);
nand U5101 (N_5101,N_4725,N_4848);
nor U5102 (N_5102,N_4545,N_4710);
or U5103 (N_5103,N_4559,N_4536);
nand U5104 (N_5104,N_4954,N_4783);
xnor U5105 (N_5105,N_4671,N_4517);
xor U5106 (N_5106,N_4969,N_4938);
and U5107 (N_5107,N_4649,N_4974);
and U5108 (N_5108,N_4955,N_4543);
xor U5109 (N_5109,N_4635,N_4950);
xnor U5110 (N_5110,N_4756,N_4591);
nand U5111 (N_5111,N_4698,N_4542);
or U5112 (N_5112,N_4505,N_4792);
and U5113 (N_5113,N_4947,N_4539);
xor U5114 (N_5114,N_4916,N_4574);
nand U5115 (N_5115,N_4672,N_4513);
or U5116 (N_5116,N_4749,N_4503);
nand U5117 (N_5117,N_4909,N_4855);
or U5118 (N_5118,N_4619,N_4929);
nor U5119 (N_5119,N_4739,N_4508);
xor U5120 (N_5120,N_4760,N_4666);
nand U5121 (N_5121,N_4971,N_4636);
and U5122 (N_5122,N_4959,N_4510);
xnor U5123 (N_5123,N_4535,N_4844);
nor U5124 (N_5124,N_4935,N_4738);
and U5125 (N_5125,N_4983,N_4809);
nor U5126 (N_5126,N_4621,N_4807);
or U5127 (N_5127,N_4906,N_4812);
and U5128 (N_5128,N_4600,N_4626);
xnor U5129 (N_5129,N_4668,N_4594);
and U5130 (N_5130,N_4825,N_4834);
xor U5131 (N_5131,N_4554,N_4833);
nand U5132 (N_5132,N_4850,N_4816);
xor U5133 (N_5133,N_4755,N_4802);
nor U5134 (N_5134,N_4703,N_4883);
and U5135 (N_5135,N_4721,N_4806);
nand U5136 (N_5136,N_4650,N_4933);
nand U5137 (N_5137,N_4881,N_4934);
nand U5138 (N_5138,N_4585,N_4537);
and U5139 (N_5139,N_4673,N_4838);
nor U5140 (N_5140,N_4808,N_4979);
xor U5141 (N_5141,N_4515,N_4771);
and U5142 (N_5142,N_4549,N_4766);
and U5143 (N_5143,N_4529,N_4674);
or U5144 (N_5144,N_4745,N_4948);
nor U5145 (N_5145,N_4637,N_4990);
nand U5146 (N_5146,N_4620,N_4879);
nand U5147 (N_5147,N_4723,N_4593);
nor U5148 (N_5148,N_4581,N_4532);
nor U5149 (N_5149,N_4669,N_4832);
nand U5150 (N_5150,N_4830,N_4616);
xnor U5151 (N_5151,N_4930,N_4631);
or U5152 (N_5152,N_4876,N_4627);
nor U5153 (N_5153,N_4558,N_4707);
nor U5154 (N_5154,N_4789,N_4977);
and U5155 (N_5155,N_4869,N_4978);
xnor U5156 (N_5156,N_4686,N_4689);
or U5157 (N_5157,N_4866,N_4976);
xor U5158 (N_5158,N_4565,N_4918);
or U5159 (N_5159,N_4765,N_4767);
nor U5160 (N_5160,N_4946,N_4705);
nor U5161 (N_5161,N_4779,N_4580);
nor U5162 (N_5162,N_4898,N_4575);
nor U5163 (N_5163,N_4782,N_4936);
and U5164 (N_5164,N_4596,N_4759);
and U5165 (N_5165,N_4567,N_4863);
and U5166 (N_5166,N_4847,N_4592);
or U5167 (N_5167,N_4890,N_4937);
xnor U5168 (N_5168,N_4823,N_4684);
and U5169 (N_5169,N_4841,N_4608);
xor U5170 (N_5170,N_4799,N_4757);
or U5171 (N_5171,N_4910,N_4773);
nor U5172 (N_5172,N_4589,N_4688);
nor U5173 (N_5173,N_4523,N_4897);
and U5174 (N_5174,N_4706,N_4900);
nor U5175 (N_5175,N_4831,N_4664);
and U5176 (N_5176,N_4743,N_4942);
nor U5177 (N_5177,N_4747,N_4982);
or U5178 (N_5178,N_4891,N_4598);
nor U5179 (N_5179,N_4544,N_4791);
xor U5180 (N_5180,N_4652,N_4605);
xnor U5181 (N_5181,N_4763,N_4961);
xnor U5182 (N_5182,N_4912,N_4864);
or U5183 (N_5183,N_4696,N_4966);
or U5184 (N_5184,N_4972,N_4984);
xnor U5185 (N_5185,N_4701,N_4561);
nand U5186 (N_5186,N_4998,N_4557);
and U5187 (N_5187,N_4583,N_4700);
nor U5188 (N_5188,N_4695,N_4742);
or U5189 (N_5189,N_4601,N_4993);
nand U5190 (N_5190,N_4584,N_4801);
nor U5191 (N_5191,N_4895,N_4658);
or U5192 (N_5192,N_4501,N_4661);
xor U5193 (N_5193,N_4744,N_4925);
nand U5194 (N_5194,N_4962,N_4719);
nand U5195 (N_5195,N_4740,N_4874);
nor U5196 (N_5196,N_4790,N_4967);
and U5197 (N_5197,N_4794,N_4511);
nand U5198 (N_5198,N_4776,N_4715);
or U5199 (N_5199,N_4840,N_4871);
xnor U5200 (N_5200,N_4804,N_4859);
and U5201 (N_5201,N_4622,N_4644);
nor U5202 (N_5202,N_4625,N_4774);
nor U5203 (N_5203,N_4945,N_4919);
nor U5204 (N_5204,N_4888,N_4932);
nand U5205 (N_5205,N_4953,N_4795);
nand U5206 (N_5206,N_4651,N_4903);
or U5207 (N_5207,N_4586,N_4548);
and U5208 (N_5208,N_4720,N_4772);
xnor U5209 (N_5209,N_4854,N_4758);
xnor U5210 (N_5210,N_4551,N_4713);
and U5211 (N_5211,N_4662,N_4588);
nand U5212 (N_5212,N_4578,N_4878);
or U5213 (N_5213,N_4560,N_4851);
xnor U5214 (N_5214,N_4996,N_4737);
or U5215 (N_5215,N_4568,N_4577);
or U5216 (N_5216,N_4839,N_4634);
and U5217 (N_5217,N_4618,N_4819);
or U5218 (N_5218,N_4609,N_4827);
or U5219 (N_5219,N_4518,N_4728);
xnor U5220 (N_5220,N_4981,N_4861);
or U5221 (N_5221,N_4597,N_4814);
xor U5222 (N_5222,N_4899,N_4546);
and U5223 (N_5223,N_4820,N_4902);
and U5224 (N_5224,N_4645,N_4680);
or U5225 (N_5225,N_4994,N_4641);
nor U5226 (N_5226,N_4931,N_4606);
nand U5227 (N_5227,N_4924,N_4811);
nand U5228 (N_5228,N_4784,N_4716);
and U5229 (N_5229,N_4676,N_4657);
nor U5230 (N_5230,N_4770,N_4999);
xor U5231 (N_5231,N_4717,N_4813);
nor U5232 (N_5232,N_4683,N_4576);
and U5233 (N_5233,N_4521,N_4682);
nand U5234 (N_5234,N_4677,N_4836);
and U5235 (N_5235,N_4987,N_4500);
or U5236 (N_5236,N_4858,N_4570);
xnor U5237 (N_5237,N_4904,N_4768);
and U5238 (N_5238,N_4573,N_4528);
xor U5239 (N_5239,N_4553,N_4748);
and U5240 (N_5240,N_4675,N_4952);
nor U5241 (N_5241,N_4538,N_4648);
nand U5242 (N_5242,N_4512,N_4970);
or U5243 (N_5243,N_4842,N_4886);
or U5244 (N_5244,N_4965,N_4566);
nor U5245 (N_5245,N_4867,N_4514);
nand U5246 (N_5246,N_4985,N_4975);
or U5247 (N_5247,N_4550,N_4564);
xor U5248 (N_5248,N_4785,N_4786);
xnor U5249 (N_5249,N_4633,N_4775);
and U5250 (N_5250,N_4600,N_4702);
nor U5251 (N_5251,N_4951,N_4838);
and U5252 (N_5252,N_4941,N_4629);
nor U5253 (N_5253,N_4996,N_4526);
or U5254 (N_5254,N_4602,N_4998);
nand U5255 (N_5255,N_4693,N_4614);
nand U5256 (N_5256,N_4679,N_4971);
and U5257 (N_5257,N_4830,N_4851);
or U5258 (N_5258,N_4864,N_4981);
nor U5259 (N_5259,N_4543,N_4515);
or U5260 (N_5260,N_4888,N_4737);
nor U5261 (N_5261,N_4702,N_4648);
or U5262 (N_5262,N_4861,N_4661);
nor U5263 (N_5263,N_4833,N_4717);
xor U5264 (N_5264,N_4806,N_4534);
xnor U5265 (N_5265,N_4815,N_4916);
or U5266 (N_5266,N_4847,N_4636);
nor U5267 (N_5267,N_4987,N_4835);
nand U5268 (N_5268,N_4506,N_4715);
nor U5269 (N_5269,N_4517,N_4624);
nand U5270 (N_5270,N_4902,N_4578);
nand U5271 (N_5271,N_4711,N_4860);
nor U5272 (N_5272,N_4526,N_4789);
or U5273 (N_5273,N_4609,N_4671);
nand U5274 (N_5274,N_4857,N_4982);
nor U5275 (N_5275,N_4592,N_4642);
nand U5276 (N_5276,N_4898,N_4639);
and U5277 (N_5277,N_4848,N_4600);
nand U5278 (N_5278,N_4528,N_4554);
or U5279 (N_5279,N_4865,N_4982);
and U5280 (N_5280,N_4666,N_4942);
or U5281 (N_5281,N_4891,N_4551);
xnor U5282 (N_5282,N_4950,N_4660);
nor U5283 (N_5283,N_4690,N_4595);
and U5284 (N_5284,N_4835,N_4658);
or U5285 (N_5285,N_4560,N_4929);
or U5286 (N_5286,N_4706,N_4942);
and U5287 (N_5287,N_4624,N_4911);
and U5288 (N_5288,N_4523,N_4671);
xnor U5289 (N_5289,N_4925,N_4950);
or U5290 (N_5290,N_4783,N_4769);
xor U5291 (N_5291,N_4853,N_4960);
or U5292 (N_5292,N_4745,N_4971);
nor U5293 (N_5293,N_4847,N_4724);
or U5294 (N_5294,N_4758,N_4960);
and U5295 (N_5295,N_4835,N_4971);
xor U5296 (N_5296,N_4912,N_4679);
and U5297 (N_5297,N_4836,N_4721);
xor U5298 (N_5298,N_4674,N_4798);
nor U5299 (N_5299,N_4610,N_4829);
nand U5300 (N_5300,N_4583,N_4798);
xor U5301 (N_5301,N_4939,N_4598);
nor U5302 (N_5302,N_4887,N_4911);
nand U5303 (N_5303,N_4978,N_4688);
xnor U5304 (N_5304,N_4652,N_4788);
or U5305 (N_5305,N_4643,N_4878);
or U5306 (N_5306,N_4670,N_4655);
and U5307 (N_5307,N_4850,N_4508);
xnor U5308 (N_5308,N_4602,N_4587);
or U5309 (N_5309,N_4934,N_4789);
or U5310 (N_5310,N_4558,N_4866);
or U5311 (N_5311,N_4579,N_4906);
xor U5312 (N_5312,N_4982,N_4606);
or U5313 (N_5313,N_4920,N_4549);
xor U5314 (N_5314,N_4998,N_4649);
or U5315 (N_5315,N_4548,N_4820);
nor U5316 (N_5316,N_4673,N_4597);
nor U5317 (N_5317,N_4528,N_4628);
xor U5318 (N_5318,N_4871,N_4797);
nand U5319 (N_5319,N_4666,N_4889);
and U5320 (N_5320,N_4718,N_4567);
or U5321 (N_5321,N_4996,N_4512);
and U5322 (N_5322,N_4994,N_4776);
nand U5323 (N_5323,N_4866,N_4753);
and U5324 (N_5324,N_4920,N_4605);
nand U5325 (N_5325,N_4546,N_4980);
nand U5326 (N_5326,N_4867,N_4640);
xor U5327 (N_5327,N_4646,N_4958);
and U5328 (N_5328,N_4918,N_4950);
or U5329 (N_5329,N_4895,N_4779);
nor U5330 (N_5330,N_4719,N_4637);
and U5331 (N_5331,N_4951,N_4528);
and U5332 (N_5332,N_4878,N_4774);
nor U5333 (N_5333,N_4888,N_4947);
and U5334 (N_5334,N_4550,N_4501);
and U5335 (N_5335,N_4749,N_4863);
or U5336 (N_5336,N_4673,N_4861);
nand U5337 (N_5337,N_4993,N_4666);
and U5338 (N_5338,N_4541,N_4831);
nor U5339 (N_5339,N_4637,N_4608);
and U5340 (N_5340,N_4890,N_4664);
and U5341 (N_5341,N_4617,N_4836);
nand U5342 (N_5342,N_4631,N_4646);
nand U5343 (N_5343,N_4963,N_4658);
nand U5344 (N_5344,N_4971,N_4721);
nand U5345 (N_5345,N_4763,N_4603);
and U5346 (N_5346,N_4765,N_4801);
or U5347 (N_5347,N_4810,N_4626);
nand U5348 (N_5348,N_4572,N_4918);
nor U5349 (N_5349,N_4964,N_4753);
xor U5350 (N_5350,N_4642,N_4910);
xor U5351 (N_5351,N_4931,N_4924);
nand U5352 (N_5352,N_4548,N_4617);
nor U5353 (N_5353,N_4823,N_4564);
nand U5354 (N_5354,N_4672,N_4785);
or U5355 (N_5355,N_4757,N_4687);
xor U5356 (N_5356,N_4970,N_4842);
and U5357 (N_5357,N_4978,N_4592);
nand U5358 (N_5358,N_4559,N_4548);
xor U5359 (N_5359,N_4841,N_4745);
nor U5360 (N_5360,N_4928,N_4629);
nor U5361 (N_5361,N_4641,N_4551);
xor U5362 (N_5362,N_4947,N_4667);
xnor U5363 (N_5363,N_4653,N_4648);
and U5364 (N_5364,N_4832,N_4575);
xnor U5365 (N_5365,N_4906,N_4511);
nor U5366 (N_5366,N_4842,N_4690);
or U5367 (N_5367,N_4902,N_4700);
or U5368 (N_5368,N_4578,N_4688);
and U5369 (N_5369,N_4705,N_4537);
or U5370 (N_5370,N_4760,N_4864);
and U5371 (N_5371,N_4911,N_4637);
nor U5372 (N_5372,N_4663,N_4799);
or U5373 (N_5373,N_4632,N_4653);
and U5374 (N_5374,N_4749,N_4901);
and U5375 (N_5375,N_4715,N_4652);
or U5376 (N_5376,N_4732,N_4627);
or U5377 (N_5377,N_4741,N_4666);
nand U5378 (N_5378,N_4773,N_4790);
and U5379 (N_5379,N_4859,N_4744);
nand U5380 (N_5380,N_4813,N_4600);
nand U5381 (N_5381,N_4566,N_4946);
and U5382 (N_5382,N_4637,N_4899);
and U5383 (N_5383,N_4781,N_4685);
nand U5384 (N_5384,N_4690,N_4958);
and U5385 (N_5385,N_4673,N_4890);
or U5386 (N_5386,N_4684,N_4897);
nor U5387 (N_5387,N_4876,N_4831);
and U5388 (N_5388,N_4956,N_4729);
or U5389 (N_5389,N_4600,N_4747);
nand U5390 (N_5390,N_4683,N_4910);
nand U5391 (N_5391,N_4892,N_4963);
xor U5392 (N_5392,N_4689,N_4582);
xnor U5393 (N_5393,N_4898,N_4649);
or U5394 (N_5394,N_4893,N_4629);
xor U5395 (N_5395,N_4632,N_4660);
or U5396 (N_5396,N_4913,N_4634);
nor U5397 (N_5397,N_4666,N_4695);
nor U5398 (N_5398,N_4830,N_4996);
nand U5399 (N_5399,N_4745,N_4665);
nand U5400 (N_5400,N_4827,N_4943);
nor U5401 (N_5401,N_4557,N_4573);
xnor U5402 (N_5402,N_4742,N_4758);
and U5403 (N_5403,N_4833,N_4684);
nand U5404 (N_5404,N_4891,N_4756);
and U5405 (N_5405,N_4779,N_4854);
xnor U5406 (N_5406,N_4835,N_4644);
or U5407 (N_5407,N_4982,N_4824);
and U5408 (N_5408,N_4755,N_4705);
and U5409 (N_5409,N_4599,N_4625);
xnor U5410 (N_5410,N_4798,N_4940);
nor U5411 (N_5411,N_4782,N_4716);
or U5412 (N_5412,N_4666,N_4646);
and U5413 (N_5413,N_4745,N_4668);
nor U5414 (N_5414,N_4798,N_4531);
nor U5415 (N_5415,N_4703,N_4639);
and U5416 (N_5416,N_4952,N_4946);
xor U5417 (N_5417,N_4509,N_4647);
and U5418 (N_5418,N_4929,N_4666);
nand U5419 (N_5419,N_4690,N_4619);
nor U5420 (N_5420,N_4953,N_4584);
or U5421 (N_5421,N_4590,N_4596);
and U5422 (N_5422,N_4797,N_4530);
and U5423 (N_5423,N_4550,N_4726);
nor U5424 (N_5424,N_4687,N_4633);
nor U5425 (N_5425,N_4975,N_4736);
nand U5426 (N_5426,N_4917,N_4598);
xnor U5427 (N_5427,N_4847,N_4879);
or U5428 (N_5428,N_4728,N_4617);
and U5429 (N_5429,N_4635,N_4938);
or U5430 (N_5430,N_4966,N_4693);
or U5431 (N_5431,N_4501,N_4794);
nor U5432 (N_5432,N_4880,N_4777);
nand U5433 (N_5433,N_4962,N_4743);
xnor U5434 (N_5434,N_4654,N_4718);
xor U5435 (N_5435,N_4956,N_4607);
and U5436 (N_5436,N_4549,N_4752);
nand U5437 (N_5437,N_4641,N_4571);
or U5438 (N_5438,N_4710,N_4875);
nand U5439 (N_5439,N_4713,N_4812);
and U5440 (N_5440,N_4968,N_4804);
or U5441 (N_5441,N_4951,N_4760);
nand U5442 (N_5442,N_4733,N_4925);
nor U5443 (N_5443,N_4551,N_4518);
nor U5444 (N_5444,N_4925,N_4718);
nand U5445 (N_5445,N_4743,N_4693);
and U5446 (N_5446,N_4966,N_4769);
nor U5447 (N_5447,N_4649,N_4624);
nor U5448 (N_5448,N_4979,N_4788);
nor U5449 (N_5449,N_4758,N_4588);
nor U5450 (N_5450,N_4996,N_4603);
and U5451 (N_5451,N_4746,N_4729);
or U5452 (N_5452,N_4702,N_4859);
xor U5453 (N_5453,N_4855,N_4810);
and U5454 (N_5454,N_4590,N_4612);
and U5455 (N_5455,N_4925,N_4822);
nor U5456 (N_5456,N_4869,N_4670);
or U5457 (N_5457,N_4557,N_4796);
nand U5458 (N_5458,N_4610,N_4881);
xnor U5459 (N_5459,N_4609,N_4957);
or U5460 (N_5460,N_4703,N_4754);
or U5461 (N_5461,N_4653,N_4604);
or U5462 (N_5462,N_4912,N_4850);
and U5463 (N_5463,N_4843,N_4923);
or U5464 (N_5464,N_4933,N_4726);
xnor U5465 (N_5465,N_4704,N_4735);
nand U5466 (N_5466,N_4950,N_4983);
nor U5467 (N_5467,N_4633,N_4683);
xor U5468 (N_5468,N_4999,N_4658);
xnor U5469 (N_5469,N_4879,N_4865);
nand U5470 (N_5470,N_4700,N_4763);
and U5471 (N_5471,N_4782,N_4563);
nor U5472 (N_5472,N_4883,N_4548);
and U5473 (N_5473,N_4880,N_4950);
nor U5474 (N_5474,N_4864,N_4781);
or U5475 (N_5475,N_4589,N_4777);
nand U5476 (N_5476,N_4925,N_4876);
and U5477 (N_5477,N_4992,N_4751);
nor U5478 (N_5478,N_4713,N_4613);
nand U5479 (N_5479,N_4638,N_4987);
nor U5480 (N_5480,N_4910,N_4803);
xnor U5481 (N_5481,N_4595,N_4609);
nor U5482 (N_5482,N_4531,N_4892);
nor U5483 (N_5483,N_4748,N_4783);
xnor U5484 (N_5484,N_4633,N_4576);
or U5485 (N_5485,N_4620,N_4728);
and U5486 (N_5486,N_4552,N_4632);
xnor U5487 (N_5487,N_4571,N_4700);
and U5488 (N_5488,N_4930,N_4694);
nand U5489 (N_5489,N_4667,N_4717);
xnor U5490 (N_5490,N_4741,N_4609);
or U5491 (N_5491,N_4665,N_4661);
nor U5492 (N_5492,N_4549,N_4710);
nor U5493 (N_5493,N_4619,N_4893);
or U5494 (N_5494,N_4823,N_4960);
or U5495 (N_5495,N_4637,N_4888);
nor U5496 (N_5496,N_4755,N_4841);
nand U5497 (N_5497,N_4672,N_4587);
or U5498 (N_5498,N_4518,N_4967);
nand U5499 (N_5499,N_4713,N_4864);
nor U5500 (N_5500,N_5221,N_5097);
and U5501 (N_5501,N_5313,N_5272);
and U5502 (N_5502,N_5464,N_5040);
or U5503 (N_5503,N_5268,N_5100);
nor U5504 (N_5504,N_5075,N_5046);
xor U5505 (N_5505,N_5480,N_5085);
and U5506 (N_5506,N_5438,N_5310);
xnor U5507 (N_5507,N_5465,N_5099);
or U5508 (N_5508,N_5278,N_5121);
xor U5509 (N_5509,N_5139,N_5147);
or U5510 (N_5510,N_5366,N_5160);
xor U5511 (N_5511,N_5295,N_5031);
nand U5512 (N_5512,N_5190,N_5440);
or U5513 (N_5513,N_5195,N_5140);
or U5514 (N_5514,N_5332,N_5286);
and U5515 (N_5515,N_5362,N_5111);
xnor U5516 (N_5516,N_5309,N_5342);
nand U5517 (N_5517,N_5359,N_5244);
nand U5518 (N_5518,N_5167,N_5312);
xnor U5519 (N_5519,N_5070,N_5360);
and U5520 (N_5520,N_5386,N_5300);
nand U5521 (N_5521,N_5290,N_5035);
or U5522 (N_5522,N_5135,N_5347);
or U5523 (N_5523,N_5297,N_5096);
nor U5524 (N_5524,N_5240,N_5494);
or U5525 (N_5525,N_5263,N_5447);
nand U5526 (N_5526,N_5477,N_5307);
or U5527 (N_5527,N_5433,N_5022);
xnor U5528 (N_5528,N_5110,N_5231);
nand U5529 (N_5529,N_5407,N_5496);
and U5530 (N_5530,N_5189,N_5059);
nand U5531 (N_5531,N_5044,N_5490);
xnor U5532 (N_5532,N_5245,N_5230);
or U5533 (N_5533,N_5113,N_5261);
or U5534 (N_5534,N_5020,N_5061);
or U5535 (N_5535,N_5011,N_5390);
nand U5536 (N_5536,N_5374,N_5055);
nor U5537 (N_5537,N_5393,N_5383);
nor U5538 (N_5538,N_5473,N_5306);
or U5539 (N_5539,N_5152,N_5101);
nand U5540 (N_5540,N_5304,N_5485);
nor U5541 (N_5541,N_5235,N_5158);
or U5542 (N_5542,N_5116,N_5010);
and U5543 (N_5543,N_5172,N_5267);
nor U5544 (N_5544,N_5131,N_5027);
nand U5545 (N_5545,N_5087,N_5375);
nand U5546 (N_5546,N_5081,N_5034);
xor U5547 (N_5547,N_5186,N_5319);
nor U5548 (N_5548,N_5180,N_5037);
nand U5549 (N_5549,N_5004,N_5282);
and U5550 (N_5550,N_5321,N_5466);
nand U5551 (N_5551,N_5327,N_5353);
xnor U5552 (N_5552,N_5184,N_5463);
nand U5553 (N_5553,N_5276,N_5367);
or U5554 (N_5554,N_5256,N_5076);
nand U5555 (N_5555,N_5226,N_5060);
xor U5556 (N_5556,N_5420,N_5227);
and U5557 (N_5557,N_5092,N_5161);
xor U5558 (N_5558,N_5204,N_5325);
nor U5559 (N_5559,N_5157,N_5098);
or U5560 (N_5560,N_5106,N_5082);
nor U5561 (N_5561,N_5484,N_5398);
nor U5562 (N_5562,N_5248,N_5133);
nor U5563 (N_5563,N_5224,N_5219);
nor U5564 (N_5564,N_5232,N_5188);
xor U5565 (N_5565,N_5394,N_5053);
and U5566 (N_5566,N_5437,N_5138);
xnor U5567 (N_5567,N_5399,N_5179);
nand U5568 (N_5568,N_5424,N_5411);
and U5569 (N_5569,N_5436,N_5007);
nand U5570 (N_5570,N_5124,N_5066);
nor U5571 (N_5571,N_5493,N_5350);
or U5572 (N_5572,N_5456,N_5127);
xor U5573 (N_5573,N_5457,N_5271);
nand U5574 (N_5574,N_5410,N_5459);
nand U5575 (N_5575,N_5370,N_5469);
nor U5576 (N_5576,N_5215,N_5062);
nor U5577 (N_5577,N_5210,N_5151);
xnor U5578 (N_5578,N_5299,N_5354);
xor U5579 (N_5579,N_5365,N_5146);
xor U5580 (N_5580,N_5183,N_5339);
xnor U5581 (N_5581,N_5095,N_5049);
xor U5582 (N_5582,N_5495,N_5107);
and U5583 (N_5583,N_5051,N_5264);
nand U5584 (N_5584,N_5030,N_5478);
and U5585 (N_5585,N_5218,N_5277);
or U5586 (N_5586,N_5132,N_5435);
and U5587 (N_5587,N_5439,N_5467);
or U5588 (N_5588,N_5086,N_5320);
and U5589 (N_5589,N_5200,N_5404);
nand U5590 (N_5590,N_5322,N_5036);
nor U5591 (N_5591,N_5474,N_5442);
and U5592 (N_5592,N_5067,N_5239);
nor U5593 (N_5593,N_5164,N_5250);
and U5594 (N_5594,N_5378,N_5129);
and U5595 (N_5595,N_5423,N_5364);
or U5596 (N_5596,N_5173,N_5242);
nand U5597 (N_5597,N_5185,N_5125);
nand U5598 (N_5598,N_5134,N_5130);
xor U5599 (N_5599,N_5228,N_5197);
xnor U5600 (N_5600,N_5168,N_5074);
or U5601 (N_5601,N_5213,N_5279);
or U5602 (N_5602,N_5175,N_5069);
nand U5603 (N_5603,N_5117,N_5199);
nor U5604 (N_5604,N_5249,N_5203);
nor U5605 (N_5605,N_5434,N_5006);
or U5606 (N_5606,N_5426,N_5418);
xnor U5607 (N_5607,N_5090,N_5388);
nand U5608 (N_5608,N_5225,N_5241);
nor U5609 (N_5609,N_5413,N_5104);
or U5610 (N_5610,N_5174,N_5057);
nor U5611 (N_5611,N_5311,N_5144);
and U5612 (N_5612,N_5014,N_5170);
and U5613 (N_5613,N_5289,N_5479);
nor U5614 (N_5614,N_5444,N_5032);
nand U5615 (N_5615,N_5206,N_5214);
nand U5616 (N_5616,N_5475,N_5408);
and U5617 (N_5617,N_5275,N_5016);
and U5618 (N_5618,N_5077,N_5149);
nand U5619 (N_5619,N_5455,N_5252);
nand U5620 (N_5620,N_5026,N_5191);
nor U5621 (N_5621,N_5187,N_5202);
and U5622 (N_5622,N_5155,N_5233);
xor U5623 (N_5623,N_5201,N_5222);
nor U5624 (N_5624,N_5108,N_5009);
and U5625 (N_5625,N_5453,N_5047);
nor U5626 (N_5626,N_5483,N_5247);
or U5627 (N_5627,N_5251,N_5217);
nand U5628 (N_5628,N_5294,N_5461);
and U5629 (N_5629,N_5391,N_5352);
nor U5630 (N_5630,N_5336,N_5039);
or U5631 (N_5631,N_5358,N_5220);
and U5632 (N_5632,N_5379,N_5033);
or U5633 (N_5633,N_5141,N_5102);
nand U5634 (N_5634,N_5429,N_5491);
and U5635 (N_5635,N_5093,N_5381);
or U5636 (N_5636,N_5481,N_5385);
nor U5637 (N_5637,N_5331,N_5112);
or U5638 (N_5638,N_5337,N_5340);
xnor U5639 (N_5639,N_5162,N_5323);
and U5640 (N_5640,N_5266,N_5422);
and U5641 (N_5641,N_5291,N_5476);
or U5642 (N_5642,N_5194,N_5148);
nand U5643 (N_5643,N_5403,N_5126);
nand U5644 (N_5644,N_5425,N_5431);
or U5645 (N_5645,N_5064,N_5177);
and U5646 (N_5646,N_5417,N_5389);
nand U5647 (N_5647,N_5303,N_5223);
nor U5648 (N_5648,N_5018,N_5397);
xor U5649 (N_5649,N_5171,N_5094);
nor U5650 (N_5650,N_5258,N_5013);
xor U5651 (N_5651,N_5254,N_5216);
nor U5652 (N_5652,N_5371,N_5029);
nand U5653 (N_5653,N_5209,N_5396);
nand U5654 (N_5654,N_5314,N_5302);
nand U5655 (N_5655,N_5153,N_5166);
xnor U5656 (N_5656,N_5460,N_5317);
or U5657 (N_5657,N_5377,N_5471);
nand U5658 (N_5658,N_5328,N_5255);
and U5659 (N_5659,N_5165,N_5150);
xnor U5660 (N_5660,N_5038,N_5376);
and U5661 (N_5661,N_5028,N_5283);
and U5662 (N_5662,N_5445,N_5402);
and U5663 (N_5663,N_5274,N_5163);
or U5664 (N_5664,N_5118,N_5181);
nor U5665 (N_5665,N_5497,N_5043);
xor U5666 (N_5666,N_5169,N_5285);
nor U5667 (N_5667,N_5315,N_5343);
xnor U5668 (N_5668,N_5382,N_5071);
nor U5669 (N_5669,N_5414,N_5428);
and U5670 (N_5670,N_5421,N_5293);
nor U5671 (N_5671,N_5281,N_5123);
nand U5672 (N_5672,N_5023,N_5487);
or U5673 (N_5673,N_5355,N_5156);
nor U5674 (N_5674,N_5079,N_5498);
or U5675 (N_5675,N_5265,N_5259);
nand U5676 (N_5676,N_5432,N_5091);
or U5677 (N_5677,N_5142,N_5305);
or U5678 (N_5678,N_5405,N_5119);
or U5679 (N_5679,N_5260,N_5143);
or U5680 (N_5680,N_5050,N_5229);
or U5681 (N_5681,N_5387,N_5073);
nor U5682 (N_5682,N_5330,N_5489);
and U5683 (N_5683,N_5056,N_5419);
or U5684 (N_5684,N_5395,N_5080);
nor U5685 (N_5685,N_5005,N_5198);
nor U5686 (N_5686,N_5368,N_5178);
and U5687 (N_5687,N_5045,N_5237);
and U5688 (N_5688,N_5063,N_5412);
xor U5689 (N_5689,N_5246,N_5114);
nor U5690 (N_5690,N_5012,N_5373);
nor U5691 (N_5691,N_5488,N_5262);
or U5692 (N_5692,N_5344,N_5492);
nor U5693 (N_5693,N_5472,N_5441);
nor U5694 (N_5694,N_5468,N_5019);
or U5695 (N_5695,N_5345,N_5316);
nand U5696 (N_5696,N_5334,N_5416);
and U5697 (N_5697,N_5392,N_5326);
xnor U5698 (N_5698,N_5065,N_5400);
nor U5699 (N_5699,N_5470,N_5000);
nand U5700 (N_5700,N_5351,N_5002);
and U5701 (N_5701,N_5269,N_5482);
nor U5702 (N_5702,N_5448,N_5298);
and U5703 (N_5703,N_5243,N_5292);
or U5704 (N_5704,N_5458,N_5136);
nor U5705 (N_5705,N_5041,N_5287);
nand U5706 (N_5706,N_5211,N_5212);
or U5707 (N_5707,N_5446,N_5329);
and U5708 (N_5708,N_5450,N_5443);
nor U5709 (N_5709,N_5021,N_5115);
nand U5710 (N_5710,N_5357,N_5284);
and U5711 (N_5711,N_5003,N_5145);
nor U5712 (N_5712,N_5486,N_5154);
or U5713 (N_5713,N_5338,N_5301);
xnor U5714 (N_5714,N_5058,N_5451);
or U5715 (N_5715,N_5048,N_5088);
xor U5716 (N_5716,N_5318,N_5308);
and U5717 (N_5717,N_5273,N_5369);
nand U5718 (N_5718,N_5207,N_5462);
xor U5719 (N_5719,N_5137,N_5234);
nor U5720 (N_5720,N_5356,N_5083);
and U5721 (N_5721,N_5324,N_5205);
or U5722 (N_5722,N_5361,N_5257);
nor U5723 (N_5723,N_5089,N_5333);
or U5724 (N_5724,N_5072,N_5499);
nor U5725 (N_5725,N_5159,N_5008);
or U5726 (N_5726,N_5341,N_5288);
and U5727 (N_5727,N_5024,N_5208);
nor U5728 (N_5728,N_5182,N_5363);
and U5729 (N_5729,N_5454,N_5054);
or U5730 (N_5730,N_5415,N_5015);
and U5731 (N_5731,N_5176,N_5193);
nand U5732 (N_5732,N_5346,N_5078);
or U5733 (N_5733,N_5348,N_5192);
nand U5734 (N_5734,N_5430,N_5372);
or U5735 (N_5735,N_5349,N_5238);
nand U5736 (N_5736,N_5296,N_5384);
or U5737 (N_5737,N_5409,N_5042);
xor U5738 (N_5738,N_5236,N_5196);
xor U5739 (N_5739,N_5380,N_5253);
or U5740 (N_5740,N_5401,N_5105);
nor U5741 (N_5741,N_5122,N_5084);
xnor U5742 (N_5742,N_5068,N_5120);
and U5743 (N_5743,N_5406,N_5449);
or U5744 (N_5744,N_5103,N_5427);
and U5745 (N_5745,N_5052,N_5025);
and U5746 (N_5746,N_5452,N_5335);
and U5747 (N_5747,N_5001,N_5270);
and U5748 (N_5748,N_5280,N_5109);
or U5749 (N_5749,N_5017,N_5128);
nor U5750 (N_5750,N_5203,N_5429);
xnor U5751 (N_5751,N_5009,N_5104);
nand U5752 (N_5752,N_5366,N_5222);
xor U5753 (N_5753,N_5173,N_5159);
nand U5754 (N_5754,N_5095,N_5459);
xor U5755 (N_5755,N_5307,N_5106);
nand U5756 (N_5756,N_5458,N_5198);
nand U5757 (N_5757,N_5376,N_5281);
and U5758 (N_5758,N_5158,N_5332);
or U5759 (N_5759,N_5448,N_5082);
nor U5760 (N_5760,N_5019,N_5053);
nand U5761 (N_5761,N_5209,N_5217);
and U5762 (N_5762,N_5411,N_5488);
xor U5763 (N_5763,N_5012,N_5109);
nor U5764 (N_5764,N_5141,N_5226);
xnor U5765 (N_5765,N_5414,N_5424);
or U5766 (N_5766,N_5432,N_5054);
nand U5767 (N_5767,N_5104,N_5172);
nand U5768 (N_5768,N_5064,N_5027);
nor U5769 (N_5769,N_5363,N_5030);
xor U5770 (N_5770,N_5463,N_5222);
nand U5771 (N_5771,N_5283,N_5464);
xnor U5772 (N_5772,N_5282,N_5397);
nor U5773 (N_5773,N_5289,N_5218);
or U5774 (N_5774,N_5111,N_5449);
or U5775 (N_5775,N_5239,N_5122);
xnor U5776 (N_5776,N_5132,N_5491);
nand U5777 (N_5777,N_5268,N_5372);
nand U5778 (N_5778,N_5406,N_5337);
nor U5779 (N_5779,N_5126,N_5173);
xor U5780 (N_5780,N_5113,N_5358);
and U5781 (N_5781,N_5274,N_5061);
and U5782 (N_5782,N_5221,N_5363);
or U5783 (N_5783,N_5366,N_5387);
and U5784 (N_5784,N_5219,N_5022);
xor U5785 (N_5785,N_5324,N_5201);
xnor U5786 (N_5786,N_5280,N_5140);
and U5787 (N_5787,N_5204,N_5066);
nand U5788 (N_5788,N_5209,N_5017);
nor U5789 (N_5789,N_5173,N_5384);
or U5790 (N_5790,N_5032,N_5335);
xnor U5791 (N_5791,N_5487,N_5447);
and U5792 (N_5792,N_5035,N_5451);
nand U5793 (N_5793,N_5019,N_5279);
nor U5794 (N_5794,N_5347,N_5292);
nand U5795 (N_5795,N_5061,N_5329);
nor U5796 (N_5796,N_5393,N_5364);
nand U5797 (N_5797,N_5042,N_5019);
and U5798 (N_5798,N_5062,N_5260);
xor U5799 (N_5799,N_5175,N_5014);
nor U5800 (N_5800,N_5229,N_5011);
or U5801 (N_5801,N_5064,N_5407);
nand U5802 (N_5802,N_5498,N_5213);
and U5803 (N_5803,N_5335,N_5451);
or U5804 (N_5804,N_5275,N_5450);
and U5805 (N_5805,N_5029,N_5094);
nand U5806 (N_5806,N_5459,N_5426);
and U5807 (N_5807,N_5049,N_5408);
or U5808 (N_5808,N_5478,N_5389);
xnor U5809 (N_5809,N_5441,N_5260);
xor U5810 (N_5810,N_5042,N_5420);
nand U5811 (N_5811,N_5428,N_5433);
and U5812 (N_5812,N_5173,N_5200);
or U5813 (N_5813,N_5140,N_5145);
nand U5814 (N_5814,N_5005,N_5120);
nand U5815 (N_5815,N_5008,N_5320);
or U5816 (N_5816,N_5067,N_5423);
xnor U5817 (N_5817,N_5384,N_5410);
xor U5818 (N_5818,N_5470,N_5489);
nand U5819 (N_5819,N_5034,N_5304);
nor U5820 (N_5820,N_5123,N_5435);
nor U5821 (N_5821,N_5083,N_5243);
nand U5822 (N_5822,N_5279,N_5363);
or U5823 (N_5823,N_5166,N_5322);
nor U5824 (N_5824,N_5108,N_5240);
nor U5825 (N_5825,N_5275,N_5147);
and U5826 (N_5826,N_5305,N_5139);
and U5827 (N_5827,N_5166,N_5037);
nand U5828 (N_5828,N_5023,N_5245);
nand U5829 (N_5829,N_5320,N_5088);
nor U5830 (N_5830,N_5258,N_5315);
and U5831 (N_5831,N_5218,N_5484);
or U5832 (N_5832,N_5304,N_5298);
or U5833 (N_5833,N_5016,N_5360);
nand U5834 (N_5834,N_5455,N_5150);
and U5835 (N_5835,N_5499,N_5478);
nand U5836 (N_5836,N_5394,N_5433);
xnor U5837 (N_5837,N_5268,N_5106);
xnor U5838 (N_5838,N_5474,N_5148);
and U5839 (N_5839,N_5240,N_5233);
nor U5840 (N_5840,N_5117,N_5382);
or U5841 (N_5841,N_5443,N_5454);
nand U5842 (N_5842,N_5061,N_5194);
xor U5843 (N_5843,N_5492,N_5098);
or U5844 (N_5844,N_5328,N_5238);
nand U5845 (N_5845,N_5026,N_5245);
xor U5846 (N_5846,N_5038,N_5319);
xnor U5847 (N_5847,N_5214,N_5108);
xor U5848 (N_5848,N_5002,N_5232);
xor U5849 (N_5849,N_5219,N_5018);
nor U5850 (N_5850,N_5003,N_5377);
or U5851 (N_5851,N_5155,N_5497);
and U5852 (N_5852,N_5293,N_5254);
or U5853 (N_5853,N_5024,N_5198);
xor U5854 (N_5854,N_5322,N_5160);
or U5855 (N_5855,N_5213,N_5070);
or U5856 (N_5856,N_5045,N_5136);
nor U5857 (N_5857,N_5330,N_5083);
and U5858 (N_5858,N_5046,N_5020);
xnor U5859 (N_5859,N_5470,N_5018);
xnor U5860 (N_5860,N_5029,N_5071);
and U5861 (N_5861,N_5280,N_5163);
nand U5862 (N_5862,N_5112,N_5018);
nand U5863 (N_5863,N_5339,N_5040);
or U5864 (N_5864,N_5137,N_5307);
nor U5865 (N_5865,N_5327,N_5275);
xnor U5866 (N_5866,N_5020,N_5332);
xor U5867 (N_5867,N_5021,N_5279);
and U5868 (N_5868,N_5311,N_5120);
nor U5869 (N_5869,N_5011,N_5030);
nand U5870 (N_5870,N_5190,N_5018);
xor U5871 (N_5871,N_5258,N_5314);
nor U5872 (N_5872,N_5424,N_5149);
nor U5873 (N_5873,N_5125,N_5131);
nand U5874 (N_5874,N_5390,N_5468);
nand U5875 (N_5875,N_5335,N_5435);
nor U5876 (N_5876,N_5492,N_5425);
and U5877 (N_5877,N_5299,N_5308);
and U5878 (N_5878,N_5350,N_5369);
and U5879 (N_5879,N_5000,N_5036);
nor U5880 (N_5880,N_5046,N_5188);
nor U5881 (N_5881,N_5014,N_5411);
or U5882 (N_5882,N_5330,N_5265);
xor U5883 (N_5883,N_5068,N_5091);
xnor U5884 (N_5884,N_5007,N_5483);
or U5885 (N_5885,N_5420,N_5404);
or U5886 (N_5886,N_5398,N_5435);
nor U5887 (N_5887,N_5224,N_5424);
or U5888 (N_5888,N_5493,N_5196);
or U5889 (N_5889,N_5398,N_5382);
xor U5890 (N_5890,N_5458,N_5014);
xnor U5891 (N_5891,N_5239,N_5432);
or U5892 (N_5892,N_5451,N_5389);
or U5893 (N_5893,N_5381,N_5068);
nand U5894 (N_5894,N_5120,N_5416);
nor U5895 (N_5895,N_5169,N_5071);
xnor U5896 (N_5896,N_5193,N_5369);
and U5897 (N_5897,N_5077,N_5380);
xor U5898 (N_5898,N_5094,N_5086);
nand U5899 (N_5899,N_5208,N_5319);
and U5900 (N_5900,N_5247,N_5429);
nor U5901 (N_5901,N_5269,N_5432);
nand U5902 (N_5902,N_5213,N_5365);
xor U5903 (N_5903,N_5371,N_5317);
or U5904 (N_5904,N_5181,N_5495);
nor U5905 (N_5905,N_5010,N_5387);
nand U5906 (N_5906,N_5039,N_5286);
or U5907 (N_5907,N_5093,N_5472);
or U5908 (N_5908,N_5010,N_5108);
and U5909 (N_5909,N_5300,N_5001);
nand U5910 (N_5910,N_5328,N_5130);
nor U5911 (N_5911,N_5429,N_5391);
xor U5912 (N_5912,N_5025,N_5446);
xor U5913 (N_5913,N_5463,N_5170);
xnor U5914 (N_5914,N_5408,N_5266);
nand U5915 (N_5915,N_5314,N_5217);
nor U5916 (N_5916,N_5079,N_5165);
nand U5917 (N_5917,N_5104,N_5252);
or U5918 (N_5918,N_5456,N_5060);
nor U5919 (N_5919,N_5317,N_5248);
or U5920 (N_5920,N_5385,N_5324);
nand U5921 (N_5921,N_5382,N_5303);
or U5922 (N_5922,N_5153,N_5177);
or U5923 (N_5923,N_5471,N_5393);
or U5924 (N_5924,N_5175,N_5410);
nand U5925 (N_5925,N_5228,N_5103);
nor U5926 (N_5926,N_5239,N_5309);
or U5927 (N_5927,N_5274,N_5349);
and U5928 (N_5928,N_5094,N_5432);
nand U5929 (N_5929,N_5041,N_5340);
and U5930 (N_5930,N_5207,N_5495);
or U5931 (N_5931,N_5017,N_5169);
nor U5932 (N_5932,N_5477,N_5329);
and U5933 (N_5933,N_5304,N_5224);
nand U5934 (N_5934,N_5274,N_5177);
nor U5935 (N_5935,N_5376,N_5481);
nor U5936 (N_5936,N_5001,N_5487);
nor U5937 (N_5937,N_5326,N_5429);
xnor U5938 (N_5938,N_5238,N_5060);
and U5939 (N_5939,N_5499,N_5054);
nand U5940 (N_5940,N_5481,N_5105);
and U5941 (N_5941,N_5453,N_5433);
nand U5942 (N_5942,N_5337,N_5080);
and U5943 (N_5943,N_5424,N_5273);
and U5944 (N_5944,N_5123,N_5035);
or U5945 (N_5945,N_5284,N_5067);
xor U5946 (N_5946,N_5439,N_5284);
xor U5947 (N_5947,N_5419,N_5069);
and U5948 (N_5948,N_5071,N_5493);
xor U5949 (N_5949,N_5495,N_5498);
nor U5950 (N_5950,N_5286,N_5030);
nand U5951 (N_5951,N_5263,N_5129);
nand U5952 (N_5952,N_5096,N_5017);
or U5953 (N_5953,N_5451,N_5160);
nor U5954 (N_5954,N_5142,N_5249);
nand U5955 (N_5955,N_5283,N_5077);
or U5956 (N_5956,N_5140,N_5448);
nor U5957 (N_5957,N_5489,N_5085);
nand U5958 (N_5958,N_5346,N_5428);
or U5959 (N_5959,N_5189,N_5450);
nor U5960 (N_5960,N_5169,N_5255);
xor U5961 (N_5961,N_5227,N_5104);
xnor U5962 (N_5962,N_5112,N_5151);
nand U5963 (N_5963,N_5344,N_5270);
and U5964 (N_5964,N_5239,N_5411);
or U5965 (N_5965,N_5188,N_5274);
and U5966 (N_5966,N_5134,N_5411);
nand U5967 (N_5967,N_5486,N_5066);
nand U5968 (N_5968,N_5234,N_5140);
xor U5969 (N_5969,N_5390,N_5172);
xor U5970 (N_5970,N_5403,N_5301);
xnor U5971 (N_5971,N_5249,N_5492);
nor U5972 (N_5972,N_5288,N_5089);
xnor U5973 (N_5973,N_5236,N_5323);
and U5974 (N_5974,N_5378,N_5198);
nor U5975 (N_5975,N_5277,N_5150);
nand U5976 (N_5976,N_5179,N_5489);
or U5977 (N_5977,N_5173,N_5045);
nand U5978 (N_5978,N_5255,N_5058);
or U5979 (N_5979,N_5170,N_5064);
or U5980 (N_5980,N_5020,N_5300);
xor U5981 (N_5981,N_5434,N_5460);
xnor U5982 (N_5982,N_5367,N_5116);
and U5983 (N_5983,N_5296,N_5052);
and U5984 (N_5984,N_5432,N_5123);
and U5985 (N_5985,N_5192,N_5163);
or U5986 (N_5986,N_5156,N_5335);
xnor U5987 (N_5987,N_5110,N_5144);
xnor U5988 (N_5988,N_5339,N_5151);
xnor U5989 (N_5989,N_5342,N_5238);
nor U5990 (N_5990,N_5242,N_5409);
nand U5991 (N_5991,N_5248,N_5301);
xnor U5992 (N_5992,N_5120,N_5459);
xor U5993 (N_5993,N_5310,N_5088);
nor U5994 (N_5994,N_5436,N_5165);
or U5995 (N_5995,N_5184,N_5306);
or U5996 (N_5996,N_5221,N_5246);
xnor U5997 (N_5997,N_5251,N_5011);
and U5998 (N_5998,N_5395,N_5117);
xnor U5999 (N_5999,N_5241,N_5194);
nand U6000 (N_6000,N_5916,N_5768);
xnor U6001 (N_6001,N_5668,N_5999);
or U6002 (N_6002,N_5855,N_5681);
or U6003 (N_6003,N_5536,N_5640);
xnor U6004 (N_6004,N_5782,N_5862);
or U6005 (N_6005,N_5949,N_5998);
xor U6006 (N_6006,N_5910,N_5856);
and U6007 (N_6007,N_5930,N_5599);
nand U6008 (N_6008,N_5873,N_5893);
or U6009 (N_6009,N_5528,N_5787);
xor U6010 (N_6010,N_5967,N_5617);
and U6011 (N_6011,N_5915,N_5690);
nor U6012 (N_6012,N_5650,N_5937);
nand U6013 (N_6013,N_5946,N_5996);
or U6014 (N_6014,N_5541,N_5621);
nand U6015 (N_6015,N_5649,N_5978);
and U6016 (N_6016,N_5812,N_5721);
xnor U6017 (N_6017,N_5711,N_5685);
xnor U6018 (N_6018,N_5836,N_5509);
nand U6019 (N_6019,N_5706,N_5713);
and U6020 (N_6020,N_5882,N_5725);
xor U6021 (N_6021,N_5973,N_5620);
nor U6022 (N_6022,N_5615,N_5515);
or U6023 (N_6023,N_5993,N_5982);
or U6024 (N_6024,N_5689,N_5866);
nor U6025 (N_6025,N_5687,N_5994);
nor U6026 (N_6026,N_5688,N_5924);
nand U6027 (N_6027,N_5677,N_5719);
or U6028 (N_6028,N_5563,N_5814);
and U6029 (N_6029,N_5817,N_5618);
and U6030 (N_6030,N_5844,N_5979);
xnor U6031 (N_6031,N_5686,N_5842);
and U6032 (N_6032,N_5631,N_5543);
and U6033 (N_6033,N_5943,N_5869);
nand U6034 (N_6034,N_5673,N_5786);
xor U6035 (N_6035,N_5763,N_5665);
or U6036 (N_6036,N_5709,N_5744);
nand U6037 (N_6037,N_5789,N_5902);
nor U6038 (N_6038,N_5761,N_5586);
nor U6039 (N_6039,N_5974,N_5992);
nor U6040 (N_6040,N_5818,N_5566);
and U6041 (N_6041,N_5820,N_5561);
or U6042 (N_6042,N_5634,N_5735);
nor U6043 (N_6043,N_5590,N_5717);
or U6044 (N_6044,N_5513,N_5624);
nand U6045 (N_6045,N_5506,N_5642);
or U6046 (N_6046,N_5582,N_5762);
and U6047 (N_6047,N_5554,N_5635);
xor U6048 (N_6048,N_5504,N_5813);
or U6049 (N_6049,N_5770,N_5553);
nand U6050 (N_6050,N_5895,N_5790);
and U6051 (N_6051,N_5560,N_5914);
nand U6052 (N_6052,N_5801,N_5609);
nand U6053 (N_6053,N_5746,N_5722);
and U6054 (N_6054,N_5905,N_5675);
or U6055 (N_6055,N_5824,N_5971);
nand U6056 (N_6056,N_5573,N_5904);
xnor U6057 (N_6057,N_5773,N_5714);
nor U6058 (N_6058,N_5991,N_5832);
nor U6059 (N_6059,N_5661,N_5843);
and U6060 (N_6060,N_5784,N_5696);
or U6061 (N_6061,N_5908,N_5750);
and U6062 (N_6062,N_5779,N_5984);
xor U6063 (N_6063,N_5648,N_5575);
xnor U6064 (N_6064,N_5864,N_5512);
nand U6065 (N_6065,N_5546,N_5516);
xnor U6066 (N_6066,N_5596,N_5990);
xnor U6067 (N_6067,N_5652,N_5568);
xor U6068 (N_6068,N_5743,N_5619);
or U6069 (N_6069,N_5637,N_5802);
xor U6070 (N_6070,N_5753,N_5727);
and U6071 (N_6071,N_5752,N_5986);
xor U6072 (N_6072,N_5574,N_5759);
xor U6073 (N_6073,N_5863,N_5851);
nand U6074 (N_6074,N_5948,N_5874);
or U6075 (N_6075,N_5583,N_5955);
or U6076 (N_6076,N_5976,N_5788);
nand U6077 (N_6077,N_5822,N_5780);
xnor U6078 (N_6078,N_5913,N_5796);
nand U6079 (N_6079,N_5923,N_5731);
or U6080 (N_6080,N_5886,N_5636);
xnor U6081 (N_6081,N_5699,N_5704);
or U6082 (N_6082,N_5738,N_5691);
nand U6083 (N_6083,N_5607,N_5867);
and U6084 (N_6084,N_5981,N_5745);
nand U6085 (N_6085,N_5580,N_5524);
xnor U6086 (N_6086,N_5645,N_5859);
xnor U6087 (N_6087,N_5933,N_5584);
or U6088 (N_6088,N_5678,N_5868);
or U6089 (N_6089,N_5540,N_5847);
or U6090 (N_6090,N_5920,N_5997);
and U6091 (N_6091,N_5680,N_5833);
xor U6092 (N_6092,N_5800,N_5811);
and U6093 (N_6093,N_5537,N_5903);
xor U6094 (N_6094,N_5877,N_5906);
and U6095 (N_6095,N_5989,N_5751);
nor U6096 (N_6096,N_5896,N_5581);
nor U6097 (N_6097,N_5959,N_5939);
nand U6098 (N_6098,N_5671,N_5659);
nand U6099 (N_6099,N_5942,N_5600);
xnor U6100 (N_6100,N_5527,N_5769);
nand U6101 (N_6101,N_5733,N_5736);
nor U6102 (N_6102,N_5625,N_5849);
or U6103 (N_6103,N_5576,N_5593);
or U6104 (N_6104,N_5819,N_5841);
xor U6105 (N_6105,N_5785,N_5657);
or U6106 (N_6106,N_5660,N_5826);
xor U6107 (N_6107,N_5845,N_5823);
and U6108 (N_6108,N_5771,N_5589);
and U6109 (N_6109,N_5718,N_5775);
xnor U6110 (N_6110,N_5792,N_5684);
nand U6111 (N_6111,N_5928,N_5623);
nor U6112 (N_6112,N_5508,N_5632);
and U6113 (N_6113,N_5518,N_5754);
nor U6114 (N_6114,N_5676,N_5557);
xnor U6115 (N_6115,N_5591,N_5918);
nand U6116 (N_6116,N_5952,N_5551);
and U6117 (N_6117,N_5555,N_5737);
nor U6118 (N_6118,N_5900,N_5726);
and U6119 (N_6119,N_5764,N_5977);
nand U6120 (N_6120,N_5988,N_5598);
nand U6121 (N_6121,N_5556,N_5892);
and U6122 (N_6122,N_5940,N_5562);
nand U6123 (N_6123,N_5532,N_5683);
nand U6124 (N_6124,N_5647,N_5610);
and U6125 (N_6125,N_5783,N_5629);
nor U6126 (N_6126,N_5578,N_5672);
and U6127 (N_6127,N_5502,N_5837);
or U6128 (N_6128,N_5963,N_5549);
nand U6129 (N_6129,N_5700,N_5564);
and U6130 (N_6130,N_5626,N_5565);
nor U6131 (N_6131,N_5611,N_5797);
and U6132 (N_6132,N_5740,N_5897);
or U6133 (N_6133,N_5523,N_5756);
nand U6134 (N_6134,N_5798,N_5748);
and U6135 (N_6135,N_5881,N_5664);
nand U6136 (N_6136,N_5934,N_5970);
xor U6137 (N_6137,N_5550,N_5693);
nor U6138 (N_6138,N_5932,N_5935);
or U6139 (N_6139,N_5875,N_5912);
nand U6140 (N_6140,N_5529,N_5876);
nand U6141 (N_6141,N_5511,N_5601);
nor U6142 (N_6142,N_5968,N_5644);
and U6143 (N_6143,N_5834,N_5547);
nor U6144 (N_6144,N_5747,N_5503);
nor U6145 (N_6145,N_5641,N_5791);
nand U6146 (N_6146,N_5957,N_5653);
nor U6147 (N_6147,N_5911,N_5606);
or U6148 (N_6148,N_5692,N_5669);
or U6149 (N_6149,N_5519,N_5850);
xnor U6150 (N_6150,N_5778,N_5835);
nand U6151 (N_6151,N_5838,N_5694);
or U6152 (N_6152,N_5674,N_5720);
nor U6153 (N_6153,N_5938,N_5885);
nor U6154 (N_6154,N_5517,N_5616);
and U6155 (N_6155,N_5953,N_5701);
and U6156 (N_6156,N_5670,N_5894);
and U6157 (N_6157,N_5871,N_5739);
nand U6158 (N_6158,N_5898,N_5947);
xnor U6159 (N_6159,N_5630,N_5567);
nand U6160 (N_6160,N_5585,N_5816);
and U6161 (N_6161,N_5776,N_5579);
nor U6162 (N_6162,N_5899,N_5954);
nor U6163 (N_6163,N_5917,N_5526);
xor U6164 (N_6164,N_5907,N_5588);
or U6165 (N_6165,N_5919,N_5945);
nor U6166 (N_6166,N_5821,N_5883);
and U6167 (N_6167,N_5995,N_5602);
and U6168 (N_6168,N_5538,N_5890);
nor U6169 (N_6169,N_5975,N_5950);
nand U6170 (N_6170,N_5655,N_5522);
nor U6171 (N_6171,N_5742,N_5951);
nor U6172 (N_6172,N_5865,N_5805);
nand U6173 (N_6173,N_5697,N_5741);
nand U6174 (N_6174,N_5716,N_5570);
or U6175 (N_6175,N_5707,N_5732);
nor U6176 (N_6176,N_5531,N_5682);
nor U6177 (N_6177,N_5533,N_5558);
or U6178 (N_6178,N_5807,N_5983);
and U6179 (N_6179,N_5825,N_5854);
nand U6180 (N_6180,N_5929,N_5887);
xnor U6181 (N_6181,N_5622,N_5852);
or U6182 (N_6182,N_5901,N_5605);
nor U6183 (N_6183,N_5931,N_5829);
and U6184 (N_6184,N_5848,N_5839);
nor U6185 (N_6185,N_5639,N_5521);
and U6186 (N_6186,N_5651,N_5514);
xor U6187 (N_6187,N_5643,N_5815);
or U6188 (N_6188,N_5808,N_5860);
or U6189 (N_6189,N_5666,N_5760);
or U6190 (N_6190,N_5972,N_5827);
and U6191 (N_6191,N_5872,N_5799);
nor U6192 (N_6192,N_5962,N_5758);
nand U6193 (N_6193,N_5628,N_5708);
xnor U6194 (N_6194,N_5729,N_5638);
or U6195 (N_6195,N_5510,N_5724);
and U6196 (N_6196,N_5548,N_5597);
and U6197 (N_6197,N_5958,N_5781);
or U6198 (N_6198,N_5656,N_5831);
and U6199 (N_6199,N_5987,N_5695);
xnor U6200 (N_6200,N_5803,N_5774);
nand U6201 (N_6201,N_5840,N_5927);
or U6202 (N_6202,N_5880,N_5956);
and U6203 (N_6203,N_5667,N_5534);
nand U6204 (N_6204,N_5730,N_5594);
xor U6205 (N_6205,N_5941,N_5544);
nand U6206 (N_6206,N_5870,N_5961);
nor U6207 (N_6207,N_5545,N_5734);
xnor U6208 (N_6208,N_5595,N_5587);
or U6209 (N_6209,N_5794,N_5633);
and U6210 (N_6210,N_5944,N_5654);
or U6211 (N_6211,N_5765,N_5853);
and U6212 (N_6212,N_5804,N_5936);
nor U6213 (N_6213,N_5712,N_5525);
xnor U6214 (N_6214,N_5969,N_5608);
and U6215 (N_6215,N_5530,N_5889);
and U6216 (N_6216,N_5809,N_5612);
xor U6217 (N_6217,N_5658,N_5909);
nand U6218 (N_6218,N_5960,N_5662);
nor U6219 (N_6219,N_5926,N_5922);
xnor U6220 (N_6220,N_5679,N_5964);
nor U6221 (N_6221,N_5879,N_5806);
nand U6222 (N_6222,N_5793,N_5577);
xor U6223 (N_6223,N_5592,N_5663);
xnor U6224 (N_6224,N_5705,N_5878);
xnor U6225 (N_6225,N_5569,N_5846);
xor U6226 (N_6226,N_5728,N_5749);
nand U6227 (N_6227,N_5966,N_5572);
nand U6228 (N_6228,N_5795,N_5965);
and U6229 (N_6229,N_5921,N_5571);
xor U6230 (N_6230,N_5884,N_5604);
and U6231 (N_6231,N_5603,N_5858);
or U6232 (N_6232,N_5505,N_5613);
or U6233 (N_6233,N_5698,N_5535);
or U6234 (N_6234,N_5542,N_5715);
xnor U6235 (N_6235,N_5857,N_5539);
xor U6236 (N_6236,N_5925,N_5702);
xnor U6237 (N_6237,N_5710,N_5766);
nand U6238 (N_6238,N_5985,N_5552);
or U6239 (N_6239,N_5501,N_5767);
or U6240 (N_6240,N_5810,N_5559);
xor U6241 (N_6241,N_5772,N_5723);
nor U6242 (N_6242,N_5830,N_5828);
and U6243 (N_6243,N_5703,N_5755);
or U6244 (N_6244,N_5520,N_5500);
xor U6245 (N_6245,N_5646,N_5757);
or U6246 (N_6246,N_5627,N_5861);
and U6247 (N_6247,N_5614,N_5888);
or U6248 (N_6248,N_5980,N_5777);
nand U6249 (N_6249,N_5891,N_5507);
nor U6250 (N_6250,N_5798,N_5550);
xnor U6251 (N_6251,N_5863,N_5709);
and U6252 (N_6252,N_5714,N_5686);
nor U6253 (N_6253,N_5822,N_5833);
xnor U6254 (N_6254,N_5661,N_5616);
nor U6255 (N_6255,N_5764,N_5986);
xor U6256 (N_6256,N_5597,N_5799);
xor U6257 (N_6257,N_5586,N_5914);
nor U6258 (N_6258,N_5951,N_5973);
nand U6259 (N_6259,N_5942,N_5701);
nor U6260 (N_6260,N_5983,N_5772);
nor U6261 (N_6261,N_5902,N_5878);
nand U6262 (N_6262,N_5969,N_5628);
nand U6263 (N_6263,N_5763,N_5833);
or U6264 (N_6264,N_5770,N_5522);
nand U6265 (N_6265,N_5588,N_5523);
xor U6266 (N_6266,N_5636,N_5908);
xnor U6267 (N_6267,N_5997,N_5757);
or U6268 (N_6268,N_5721,N_5926);
nor U6269 (N_6269,N_5995,N_5510);
xnor U6270 (N_6270,N_5969,N_5816);
nand U6271 (N_6271,N_5552,N_5860);
or U6272 (N_6272,N_5811,N_5815);
xnor U6273 (N_6273,N_5950,N_5991);
nor U6274 (N_6274,N_5643,N_5626);
xor U6275 (N_6275,N_5934,N_5684);
xnor U6276 (N_6276,N_5970,N_5609);
or U6277 (N_6277,N_5985,N_5533);
or U6278 (N_6278,N_5935,N_5693);
or U6279 (N_6279,N_5874,N_5951);
or U6280 (N_6280,N_5650,N_5550);
or U6281 (N_6281,N_5979,N_5967);
and U6282 (N_6282,N_5943,N_5650);
or U6283 (N_6283,N_5959,N_5544);
or U6284 (N_6284,N_5912,N_5662);
nor U6285 (N_6285,N_5553,N_5779);
or U6286 (N_6286,N_5738,N_5954);
and U6287 (N_6287,N_5617,N_5896);
and U6288 (N_6288,N_5697,N_5867);
or U6289 (N_6289,N_5768,N_5754);
nor U6290 (N_6290,N_5988,N_5912);
and U6291 (N_6291,N_5564,N_5821);
or U6292 (N_6292,N_5922,N_5662);
nand U6293 (N_6293,N_5608,N_5797);
nor U6294 (N_6294,N_5941,N_5727);
or U6295 (N_6295,N_5553,N_5953);
and U6296 (N_6296,N_5717,N_5685);
nor U6297 (N_6297,N_5942,N_5906);
and U6298 (N_6298,N_5916,N_5855);
xnor U6299 (N_6299,N_5841,N_5683);
and U6300 (N_6300,N_5667,N_5850);
nand U6301 (N_6301,N_5947,N_5540);
and U6302 (N_6302,N_5623,N_5960);
nor U6303 (N_6303,N_5780,N_5673);
and U6304 (N_6304,N_5511,N_5915);
nor U6305 (N_6305,N_5755,N_5730);
nor U6306 (N_6306,N_5766,N_5667);
nor U6307 (N_6307,N_5961,N_5660);
nor U6308 (N_6308,N_5971,N_5671);
or U6309 (N_6309,N_5810,N_5589);
nand U6310 (N_6310,N_5936,N_5939);
nand U6311 (N_6311,N_5688,N_5808);
nand U6312 (N_6312,N_5734,N_5711);
and U6313 (N_6313,N_5624,N_5994);
nand U6314 (N_6314,N_5982,N_5996);
nor U6315 (N_6315,N_5909,N_5530);
or U6316 (N_6316,N_5863,N_5797);
and U6317 (N_6317,N_5654,N_5842);
and U6318 (N_6318,N_5868,N_5743);
nor U6319 (N_6319,N_5881,N_5794);
xnor U6320 (N_6320,N_5734,N_5830);
nor U6321 (N_6321,N_5542,N_5983);
and U6322 (N_6322,N_5890,N_5516);
nand U6323 (N_6323,N_5741,N_5995);
and U6324 (N_6324,N_5995,N_5922);
nor U6325 (N_6325,N_5915,N_5503);
nand U6326 (N_6326,N_5737,N_5663);
nor U6327 (N_6327,N_5981,N_5518);
or U6328 (N_6328,N_5983,N_5852);
nor U6329 (N_6329,N_5874,N_5554);
xor U6330 (N_6330,N_5661,N_5701);
nand U6331 (N_6331,N_5806,N_5994);
nand U6332 (N_6332,N_5921,N_5718);
nand U6333 (N_6333,N_5922,N_5632);
xor U6334 (N_6334,N_5852,N_5576);
nand U6335 (N_6335,N_5896,N_5747);
nand U6336 (N_6336,N_5935,N_5941);
nor U6337 (N_6337,N_5869,N_5872);
xnor U6338 (N_6338,N_5796,N_5989);
nor U6339 (N_6339,N_5507,N_5837);
and U6340 (N_6340,N_5604,N_5506);
xor U6341 (N_6341,N_5721,N_5513);
nand U6342 (N_6342,N_5533,N_5563);
xnor U6343 (N_6343,N_5728,N_5907);
xor U6344 (N_6344,N_5978,N_5838);
xor U6345 (N_6345,N_5685,N_5862);
nor U6346 (N_6346,N_5826,N_5510);
or U6347 (N_6347,N_5651,N_5826);
nand U6348 (N_6348,N_5603,N_5511);
and U6349 (N_6349,N_5521,N_5507);
xor U6350 (N_6350,N_5603,N_5664);
nor U6351 (N_6351,N_5528,N_5521);
or U6352 (N_6352,N_5750,N_5751);
or U6353 (N_6353,N_5626,N_5839);
or U6354 (N_6354,N_5910,N_5621);
nand U6355 (N_6355,N_5650,N_5947);
and U6356 (N_6356,N_5555,N_5721);
nand U6357 (N_6357,N_5593,N_5597);
and U6358 (N_6358,N_5521,N_5728);
nor U6359 (N_6359,N_5952,N_5888);
nor U6360 (N_6360,N_5646,N_5924);
nand U6361 (N_6361,N_5742,N_5981);
xor U6362 (N_6362,N_5818,N_5803);
xnor U6363 (N_6363,N_5833,N_5797);
nor U6364 (N_6364,N_5514,N_5899);
and U6365 (N_6365,N_5521,N_5756);
or U6366 (N_6366,N_5644,N_5557);
nand U6367 (N_6367,N_5518,N_5554);
nand U6368 (N_6368,N_5639,N_5788);
xor U6369 (N_6369,N_5691,N_5546);
or U6370 (N_6370,N_5906,N_5588);
and U6371 (N_6371,N_5717,N_5828);
or U6372 (N_6372,N_5626,N_5734);
and U6373 (N_6373,N_5807,N_5843);
nand U6374 (N_6374,N_5706,N_5524);
or U6375 (N_6375,N_5675,N_5536);
and U6376 (N_6376,N_5977,N_5752);
nor U6377 (N_6377,N_5984,N_5708);
nand U6378 (N_6378,N_5798,N_5929);
and U6379 (N_6379,N_5791,N_5568);
and U6380 (N_6380,N_5573,N_5702);
or U6381 (N_6381,N_5737,N_5539);
and U6382 (N_6382,N_5783,N_5628);
xor U6383 (N_6383,N_5570,N_5584);
xnor U6384 (N_6384,N_5561,N_5619);
and U6385 (N_6385,N_5626,N_5557);
and U6386 (N_6386,N_5898,N_5670);
nor U6387 (N_6387,N_5604,N_5729);
nand U6388 (N_6388,N_5647,N_5930);
nand U6389 (N_6389,N_5675,N_5515);
or U6390 (N_6390,N_5931,N_5751);
or U6391 (N_6391,N_5632,N_5896);
nand U6392 (N_6392,N_5501,N_5895);
nand U6393 (N_6393,N_5991,N_5985);
or U6394 (N_6394,N_5906,N_5570);
or U6395 (N_6395,N_5754,N_5838);
and U6396 (N_6396,N_5815,N_5697);
nor U6397 (N_6397,N_5933,N_5831);
xnor U6398 (N_6398,N_5522,N_5684);
nor U6399 (N_6399,N_5680,N_5908);
xor U6400 (N_6400,N_5809,N_5512);
and U6401 (N_6401,N_5868,N_5844);
xnor U6402 (N_6402,N_5649,N_5835);
and U6403 (N_6403,N_5777,N_5662);
nor U6404 (N_6404,N_5550,N_5598);
xor U6405 (N_6405,N_5639,N_5590);
and U6406 (N_6406,N_5600,N_5844);
and U6407 (N_6407,N_5585,N_5625);
and U6408 (N_6408,N_5930,N_5848);
and U6409 (N_6409,N_5735,N_5693);
nand U6410 (N_6410,N_5847,N_5542);
or U6411 (N_6411,N_5535,N_5500);
nand U6412 (N_6412,N_5821,N_5956);
xor U6413 (N_6413,N_5757,N_5829);
and U6414 (N_6414,N_5675,N_5589);
nor U6415 (N_6415,N_5728,N_5631);
xnor U6416 (N_6416,N_5853,N_5655);
or U6417 (N_6417,N_5875,N_5660);
or U6418 (N_6418,N_5596,N_5693);
xor U6419 (N_6419,N_5968,N_5982);
or U6420 (N_6420,N_5992,N_5784);
or U6421 (N_6421,N_5954,N_5923);
nor U6422 (N_6422,N_5870,N_5640);
xnor U6423 (N_6423,N_5682,N_5972);
nor U6424 (N_6424,N_5965,N_5628);
and U6425 (N_6425,N_5636,N_5634);
nand U6426 (N_6426,N_5910,N_5618);
and U6427 (N_6427,N_5864,N_5804);
or U6428 (N_6428,N_5964,N_5622);
or U6429 (N_6429,N_5862,N_5518);
nand U6430 (N_6430,N_5800,N_5877);
or U6431 (N_6431,N_5529,N_5560);
xnor U6432 (N_6432,N_5794,N_5951);
nand U6433 (N_6433,N_5570,N_5975);
nand U6434 (N_6434,N_5642,N_5804);
nand U6435 (N_6435,N_5951,N_5629);
nor U6436 (N_6436,N_5529,N_5788);
xor U6437 (N_6437,N_5865,N_5588);
or U6438 (N_6438,N_5987,N_5924);
nand U6439 (N_6439,N_5805,N_5646);
nand U6440 (N_6440,N_5819,N_5776);
and U6441 (N_6441,N_5927,N_5901);
xnor U6442 (N_6442,N_5653,N_5510);
and U6443 (N_6443,N_5888,N_5625);
nand U6444 (N_6444,N_5961,N_5904);
nor U6445 (N_6445,N_5985,N_5555);
or U6446 (N_6446,N_5650,N_5849);
or U6447 (N_6447,N_5551,N_5939);
and U6448 (N_6448,N_5694,N_5991);
xor U6449 (N_6449,N_5836,N_5880);
nand U6450 (N_6450,N_5778,N_5877);
nand U6451 (N_6451,N_5639,N_5556);
and U6452 (N_6452,N_5645,N_5831);
and U6453 (N_6453,N_5544,N_5893);
or U6454 (N_6454,N_5885,N_5744);
nand U6455 (N_6455,N_5883,N_5785);
and U6456 (N_6456,N_5797,N_5746);
xnor U6457 (N_6457,N_5564,N_5587);
nor U6458 (N_6458,N_5660,N_5692);
xor U6459 (N_6459,N_5589,N_5959);
xor U6460 (N_6460,N_5790,N_5847);
nor U6461 (N_6461,N_5758,N_5915);
nor U6462 (N_6462,N_5824,N_5834);
xor U6463 (N_6463,N_5509,N_5884);
nor U6464 (N_6464,N_5968,N_5748);
xor U6465 (N_6465,N_5881,N_5821);
or U6466 (N_6466,N_5514,N_5854);
or U6467 (N_6467,N_5532,N_5571);
xnor U6468 (N_6468,N_5676,N_5529);
or U6469 (N_6469,N_5789,N_5767);
and U6470 (N_6470,N_5567,N_5855);
and U6471 (N_6471,N_5665,N_5801);
or U6472 (N_6472,N_5985,N_5825);
or U6473 (N_6473,N_5867,N_5794);
or U6474 (N_6474,N_5652,N_5759);
and U6475 (N_6475,N_5690,N_5941);
nor U6476 (N_6476,N_5805,N_5809);
nor U6477 (N_6477,N_5798,N_5597);
nor U6478 (N_6478,N_5503,N_5653);
and U6479 (N_6479,N_5577,N_5633);
and U6480 (N_6480,N_5967,N_5798);
nand U6481 (N_6481,N_5692,N_5984);
or U6482 (N_6482,N_5995,N_5603);
or U6483 (N_6483,N_5726,N_5819);
nor U6484 (N_6484,N_5917,N_5627);
xor U6485 (N_6485,N_5666,N_5538);
or U6486 (N_6486,N_5910,N_5569);
nand U6487 (N_6487,N_5615,N_5890);
or U6488 (N_6488,N_5501,N_5722);
nor U6489 (N_6489,N_5628,N_5533);
nor U6490 (N_6490,N_5712,N_5617);
xnor U6491 (N_6491,N_5558,N_5670);
xnor U6492 (N_6492,N_5815,N_5725);
or U6493 (N_6493,N_5849,N_5600);
nand U6494 (N_6494,N_5549,N_5874);
and U6495 (N_6495,N_5846,N_5836);
and U6496 (N_6496,N_5676,N_5594);
xor U6497 (N_6497,N_5696,N_5572);
nand U6498 (N_6498,N_5900,N_5787);
xnor U6499 (N_6499,N_5815,N_5601);
nand U6500 (N_6500,N_6155,N_6174);
or U6501 (N_6501,N_6491,N_6151);
or U6502 (N_6502,N_6392,N_6398);
xnor U6503 (N_6503,N_6200,N_6268);
and U6504 (N_6504,N_6424,N_6329);
or U6505 (N_6505,N_6131,N_6421);
nor U6506 (N_6506,N_6263,N_6201);
nor U6507 (N_6507,N_6395,N_6211);
nand U6508 (N_6508,N_6347,N_6095);
or U6509 (N_6509,N_6344,N_6055);
nand U6510 (N_6510,N_6429,N_6085);
nand U6511 (N_6511,N_6247,N_6291);
and U6512 (N_6512,N_6396,N_6147);
xor U6513 (N_6513,N_6399,N_6167);
xor U6514 (N_6514,N_6324,N_6454);
and U6515 (N_6515,N_6352,N_6229);
nor U6516 (N_6516,N_6099,N_6029);
nor U6517 (N_6517,N_6463,N_6388);
nand U6518 (N_6518,N_6191,N_6238);
or U6519 (N_6519,N_6407,N_6473);
nand U6520 (N_6520,N_6216,N_6348);
or U6521 (N_6521,N_6297,N_6362);
nor U6522 (N_6522,N_6036,N_6097);
nor U6523 (N_6523,N_6129,N_6124);
xnor U6524 (N_6524,N_6257,N_6168);
nor U6525 (N_6525,N_6082,N_6180);
or U6526 (N_6526,N_6276,N_6018);
and U6527 (N_6527,N_6374,N_6123);
and U6528 (N_6528,N_6377,N_6030);
nand U6529 (N_6529,N_6003,N_6172);
and U6530 (N_6530,N_6243,N_6420);
or U6531 (N_6531,N_6450,N_6156);
or U6532 (N_6532,N_6146,N_6499);
nand U6533 (N_6533,N_6204,N_6176);
nand U6534 (N_6534,N_6092,N_6119);
nor U6535 (N_6535,N_6014,N_6267);
xor U6536 (N_6536,N_6278,N_6230);
or U6537 (N_6537,N_6311,N_6495);
nand U6538 (N_6538,N_6397,N_6441);
xnor U6539 (N_6539,N_6056,N_6051);
nand U6540 (N_6540,N_6031,N_6426);
and U6541 (N_6541,N_6294,N_6222);
or U6542 (N_6542,N_6440,N_6116);
nand U6543 (N_6543,N_6135,N_6067);
nand U6544 (N_6544,N_6442,N_6197);
and U6545 (N_6545,N_6303,N_6449);
and U6546 (N_6546,N_6315,N_6468);
or U6547 (N_6547,N_6162,N_6017);
or U6548 (N_6548,N_6049,N_6233);
or U6549 (N_6549,N_6078,N_6312);
and U6550 (N_6550,N_6109,N_6387);
nor U6551 (N_6551,N_6260,N_6178);
and U6552 (N_6552,N_6448,N_6453);
nand U6553 (N_6553,N_6476,N_6187);
nor U6554 (N_6554,N_6313,N_6475);
nand U6555 (N_6555,N_6064,N_6089);
xor U6556 (N_6556,N_6052,N_6075);
nor U6557 (N_6557,N_6478,N_6380);
nand U6558 (N_6558,N_6159,N_6436);
nor U6559 (N_6559,N_6357,N_6431);
xnor U6560 (N_6560,N_6220,N_6009);
nor U6561 (N_6561,N_6386,N_6363);
or U6562 (N_6562,N_6337,N_6183);
or U6563 (N_6563,N_6402,N_6121);
or U6564 (N_6564,N_6193,N_6050);
xor U6565 (N_6565,N_6406,N_6203);
or U6566 (N_6566,N_6005,N_6271);
nor U6567 (N_6567,N_6213,N_6057);
and U6568 (N_6568,N_6393,N_6164);
nor U6569 (N_6569,N_6384,N_6325);
xnor U6570 (N_6570,N_6317,N_6032);
xnor U6571 (N_6571,N_6048,N_6289);
and U6572 (N_6572,N_6079,N_6210);
nand U6573 (N_6573,N_6411,N_6100);
and U6574 (N_6574,N_6319,N_6409);
or U6575 (N_6575,N_6094,N_6170);
xor U6576 (N_6576,N_6364,N_6405);
xnor U6577 (N_6577,N_6464,N_6137);
and U6578 (N_6578,N_6296,N_6343);
nor U6579 (N_6579,N_6195,N_6404);
xor U6580 (N_6580,N_6118,N_6428);
nor U6581 (N_6581,N_6308,N_6087);
or U6582 (N_6582,N_6285,N_6300);
nand U6583 (N_6583,N_6130,N_6232);
nor U6584 (N_6584,N_6321,N_6372);
or U6585 (N_6585,N_6088,N_6016);
and U6586 (N_6586,N_6173,N_6443);
and U6587 (N_6587,N_6346,N_6488);
nor U6588 (N_6588,N_6080,N_6445);
xnor U6589 (N_6589,N_6419,N_6090);
and U6590 (N_6590,N_6145,N_6305);
nand U6591 (N_6591,N_6074,N_6353);
nand U6592 (N_6592,N_6227,N_6394);
or U6593 (N_6593,N_6345,N_6113);
nor U6594 (N_6594,N_6333,N_6190);
nand U6595 (N_6595,N_6108,N_6225);
nor U6596 (N_6596,N_6073,N_6043);
nand U6597 (N_6597,N_6234,N_6390);
or U6598 (N_6598,N_6258,N_6309);
or U6599 (N_6599,N_6292,N_6077);
and U6600 (N_6600,N_6433,N_6245);
nor U6601 (N_6601,N_6483,N_6028);
or U6602 (N_6602,N_6338,N_6306);
nand U6603 (N_6603,N_6006,N_6114);
or U6604 (N_6604,N_6418,N_6007);
nor U6605 (N_6605,N_6091,N_6040);
or U6606 (N_6606,N_6215,N_6194);
nor U6607 (N_6607,N_6160,N_6142);
xnor U6608 (N_6608,N_6477,N_6015);
or U6609 (N_6609,N_6033,N_6327);
or U6610 (N_6610,N_6046,N_6360);
and U6611 (N_6611,N_6060,N_6132);
and U6612 (N_6612,N_6186,N_6320);
nor U6613 (N_6613,N_6408,N_6457);
or U6614 (N_6614,N_6027,N_6259);
xnor U6615 (N_6615,N_6410,N_6318);
and U6616 (N_6616,N_6277,N_6104);
nor U6617 (N_6617,N_6284,N_6202);
and U6618 (N_6618,N_6244,N_6106);
and U6619 (N_6619,N_6199,N_6072);
nand U6620 (N_6620,N_6492,N_6322);
nand U6621 (N_6621,N_6066,N_6103);
and U6622 (N_6622,N_6179,N_6196);
xor U6623 (N_6623,N_6169,N_6218);
or U6624 (N_6624,N_6331,N_6316);
or U6625 (N_6625,N_6228,N_6379);
nor U6626 (N_6626,N_6062,N_6008);
nor U6627 (N_6627,N_6112,N_6479);
xnor U6628 (N_6628,N_6452,N_6039);
or U6629 (N_6629,N_6021,N_6472);
or U6630 (N_6630,N_6188,N_6466);
nand U6631 (N_6631,N_6239,N_6063);
xor U6632 (N_6632,N_6148,N_6375);
and U6633 (N_6633,N_6487,N_6083);
and U6634 (N_6634,N_6430,N_6266);
xnor U6635 (N_6635,N_6274,N_6301);
xor U6636 (N_6636,N_6355,N_6280);
nand U6637 (N_6637,N_6382,N_6446);
nand U6638 (N_6638,N_6093,N_6208);
nor U6639 (N_6639,N_6154,N_6269);
xor U6640 (N_6640,N_6000,N_6181);
or U6641 (N_6641,N_6166,N_6041);
or U6642 (N_6642,N_6470,N_6059);
and U6643 (N_6643,N_6417,N_6061);
and U6644 (N_6644,N_6323,N_6149);
nand U6645 (N_6645,N_6253,N_6070);
xnor U6646 (N_6646,N_6020,N_6432);
and U6647 (N_6647,N_6310,N_6185);
xnor U6648 (N_6648,N_6367,N_6340);
nand U6649 (N_6649,N_6144,N_6351);
nor U6650 (N_6650,N_6011,N_6403);
xor U6651 (N_6651,N_6342,N_6102);
nor U6652 (N_6652,N_6358,N_6023);
xnor U6653 (N_6653,N_6486,N_6143);
nand U6654 (N_6654,N_6381,N_6383);
or U6655 (N_6655,N_6022,N_6171);
and U6656 (N_6656,N_6068,N_6349);
or U6657 (N_6657,N_6339,N_6054);
nand U6658 (N_6658,N_6425,N_6435);
or U6659 (N_6659,N_6111,N_6400);
nor U6660 (N_6660,N_6035,N_6086);
nand U6661 (N_6661,N_6444,N_6494);
nor U6662 (N_6662,N_6298,N_6336);
and U6663 (N_6663,N_6161,N_6434);
nor U6664 (N_6664,N_6013,N_6125);
and U6665 (N_6665,N_6461,N_6189);
nor U6666 (N_6666,N_6053,N_6198);
nand U6667 (N_6667,N_6423,N_6262);
xnor U6668 (N_6668,N_6350,N_6219);
nor U6669 (N_6669,N_6136,N_6065);
nor U6670 (N_6670,N_6456,N_6235);
or U6671 (N_6671,N_6150,N_6026);
xnor U6672 (N_6672,N_6415,N_6019);
and U6673 (N_6673,N_6290,N_6141);
or U6674 (N_6674,N_6412,N_6126);
or U6675 (N_6675,N_6480,N_6366);
nor U6676 (N_6676,N_6369,N_6256);
and U6677 (N_6677,N_6128,N_6458);
or U6678 (N_6678,N_6012,N_6140);
or U6679 (N_6679,N_6224,N_6101);
nand U6680 (N_6680,N_6307,N_6302);
xor U6681 (N_6681,N_6042,N_6226);
and U6682 (N_6682,N_6299,N_6044);
and U6683 (N_6683,N_6373,N_6157);
and U6684 (N_6684,N_6001,N_6165);
and U6685 (N_6685,N_6272,N_6370);
nor U6686 (N_6686,N_6138,N_6482);
or U6687 (N_6687,N_6288,N_6241);
nor U6688 (N_6688,N_6038,N_6025);
nand U6689 (N_6689,N_6221,N_6175);
or U6690 (N_6690,N_6214,N_6153);
xor U6691 (N_6691,N_6455,N_6209);
and U6692 (N_6692,N_6096,N_6184);
or U6693 (N_6693,N_6361,N_6117);
nand U6694 (N_6694,N_6481,N_6459);
and U6695 (N_6695,N_6002,N_6127);
nand U6696 (N_6696,N_6485,N_6081);
nand U6697 (N_6697,N_6439,N_6283);
nor U6698 (N_6698,N_6497,N_6401);
or U6699 (N_6699,N_6270,N_6024);
and U6700 (N_6700,N_6279,N_6314);
nor U6701 (N_6701,N_6231,N_6217);
nand U6702 (N_6702,N_6484,N_6293);
or U6703 (N_6703,N_6451,N_6490);
xnor U6704 (N_6704,N_6287,N_6192);
nor U6705 (N_6705,N_6295,N_6139);
xor U6706 (N_6706,N_6076,N_6177);
nor U6707 (N_6707,N_6326,N_6205);
xor U6708 (N_6708,N_6105,N_6493);
nor U6709 (N_6709,N_6376,N_6120);
or U6710 (N_6710,N_6416,N_6265);
nand U6711 (N_6711,N_6158,N_6447);
xnor U6712 (N_6712,N_6261,N_6223);
nand U6713 (N_6713,N_6246,N_6359);
nand U6714 (N_6714,N_6489,N_6037);
or U6715 (N_6715,N_6133,N_6236);
xor U6716 (N_6716,N_6414,N_6107);
xnor U6717 (N_6717,N_6422,N_6462);
xnor U6718 (N_6718,N_6438,N_6004);
or U6719 (N_6719,N_6356,N_6328);
and U6720 (N_6720,N_6047,N_6252);
xnor U6721 (N_6721,N_6334,N_6413);
xor U6722 (N_6722,N_6115,N_6122);
nor U6723 (N_6723,N_6354,N_6249);
and U6724 (N_6724,N_6471,N_6304);
and U6725 (N_6725,N_6378,N_6385);
or U6726 (N_6726,N_6069,N_6391);
or U6727 (N_6727,N_6389,N_6255);
or U6728 (N_6728,N_6465,N_6152);
nor U6729 (N_6729,N_6273,N_6251);
nand U6730 (N_6730,N_6332,N_6250);
xor U6731 (N_6731,N_6469,N_6281);
nor U6732 (N_6732,N_6242,N_6282);
and U6733 (N_6733,N_6240,N_6206);
nor U6734 (N_6734,N_6467,N_6371);
or U6735 (N_6735,N_6034,N_6496);
or U6736 (N_6736,N_6474,N_6098);
and U6737 (N_6737,N_6275,N_6071);
xnor U6738 (N_6738,N_6286,N_6330);
nor U6739 (N_6739,N_6045,N_6341);
or U6740 (N_6740,N_6058,N_6110);
xnor U6741 (N_6741,N_6248,N_6460);
or U6742 (N_6742,N_6084,N_6207);
or U6743 (N_6743,N_6365,N_6254);
nand U6744 (N_6744,N_6010,N_6237);
nor U6745 (N_6745,N_6427,N_6264);
nand U6746 (N_6746,N_6368,N_6163);
xor U6747 (N_6747,N_6498,N_6134);
or U6748 (N_6748,N_6182,N_6212);
xnor U6749 (N_6749,N_6335,N_6437);
and U6750 (N_6750,N_6412,N_6264);
nand U6751 (N_6751,N_6161,N_6003);
or U6752 (N_6752,N_6007,N_6291);
nand U6753 (N_6753,N_6227,N_6299);
or U6754 (N_6754,N_6083,N_6353);
nor U6755 (N_6755,N_6216,N_6226);
nand U6756 (N_6756,N_6268,N_6405);
and U6757 (N_6757,N_6335,N_6075);
xor U6758 (N_6758,N_6222,N_6081);
nand U6759 (N_6759,N_6301,N_6442);
and U6760 (N_6760,N_6458,N_6167);
and U6761 (N_6761,N_6460,N_6456);
xnor U6762 (N_6762,N_6284,N_6058);
nor U6763 (N_6763,N_6365,N_6075);
xor U6764 (N_6764,N_6122,N_6259);
nand U6765 (N_6765,N_6292,N_6263);
or U6766 (N_6766,N_6286,N_6432);
nand U6767 (N_6767,N_6278,N_6025);
nand U6768 (N_6768,N_6094,N_6027);
nor U6769 (N_6769,N_6056,N_6463);
and U6770 (N_6770,N_6262,N_6271);
or U6771 (N_6771,N_6301,N_6183);
nor U6772 (N_6772,N_6103,N_6286);
nand U6773 (N_6773,N_6218,N_6487);
and U6774 (N_6774,N_6229,N_6360);
or U6775 (N_6775,N_6463,N_6454);
nor U6776 (N_6776,N_6224,N_6202);
xor U6777 (N_6777,N_6369,N_6078);
xor U6778 (N_6778,N_6077,N_6263);
nor U6779 (N_6779,N_6291,N_6166);
xnor U6780 (N_6780,N_6298,N_6431);
nand U6781 (N_6781,N_6280,N_6408);
or U6782 (N_6782,N_6346,N_6127);
xor U6783 (N_6783,N_6020,N_6313);
nor U6784 (N_6784,N_6181,N_6356);
nand U6785 (N_6785,N_6167,N_6065);
or U6786 (N_6786,N_6281,N_6040);
nor U6787 (N_6787,N_6415,N_6270);
and U6788 (N_6788,N_6222,N_6098);
nor U6789 (N_6789,N_6137,N_6143);
or U6790 (N_6790,N_6112,N_6368);
or U6791 (N_6791,N_6294,N_6295);
xnor U6792 (N_6792,N_6418,N_6049);
or U6793 (N_6793,N_6093,N_6021);
or U6794 (N_6794,N_6021,N_6135);
nand U6795 (N_6795,N_6314,N_6344);
nor U6796 (N_6796,N_6229,N_6236);
nor U6797 (N_6797,N_6303,N_6312);
or U6798 (N_6798,N_6319,N_6426);
or U6799 (N_6799,N_6374,N_6114);
nand U6800 (N_6800,N_6336,N_6013);
and U6801 (N_6801,N_6264,N_6393);
nand U6802 (N_6802,N_6262,N_6317);
and U6803 (N_6803,N_6430,N_6177);
xor U6804 (N_6804,N_6369,N_6023);
and U6805 (N_6805,N_6410,N_6056);
xnor U6806 (N_6806,N_6439,N_6196);
xor U6807 (N_6807,N_6436,N_6480);
nor U6808 (N_6808,N_6197,N_6361);
or U6809 (N_6809,N_6450,N_6187);
xor U6810 (N_6810,N_6303,N_6243);
xor U6811 (N_6811,N_6061,N_6054);
nand U6812 (N_6812,N_6432,N_6493);
and U6813 (N_6813,N_6238,N_6470);
nor U6814 (N_6814,N_6097,N_6055);
or U6815 (N_6815,N_6211,N_6354);
or U6816 (N_6816,N_6151,N_6161);
nand U6817 (N_6817,N_6040,N_6480);
nand U6818 (N_6818,N_6147,N_6391);
nor U6819 (N_6819,N_6475,N_6389);
and U6820 (N_6820,N_6365,N_6233);
and U6821 (N_6821,N_6072,N_6037);
nand U6822 (N_6822,N_6001,N_6030);
nand U6823 (N_6823,N_6133,N_6383);
or U6824 (N_6824,N_6459,N_6421);
xor U6825 (N_6825,N_6471,N_6380);
and U6826 (N_6826,N_6404,N_6071);
or U6827 (N_6827,N_6387,N_6203);
xor U6828 (N_6828,N_6331,N_6358);
or U6829 (N_6829,N_6226,N_6045);
nand U6830 (N_6830,N_6126,N_6168);
and U6831 (N_6831,N_6112,N_6085);
or U6832 (N_6832,N_6066,N_6171);
xnor U6833 (N_6833,N_6325,N_6477);
nor U6834 (N_6834,N_6388,N_6063);
and U6835 (N_6835,N_6046,N_6204);
xnor U6836 (N_6836,N_6019,N_6324);
nand U6837 (N_6837,N_6331,N_6495);
xor U6838 (N_6838,N_6379,N_6226);
nor U6839 (N_6839,N_6393,N_6126);
or U6840 (N_6840,N_6327,N_6185);
nor U6841 (N_6841,N_6345,N_6284);
nor U6842 (N_6842,N_6283,N_6185);
nand U6843 (N_6843,N_6475,N_6022);
nand U6844 (N_6844,N_6024,N_6396);
and U6845 (N_6845,N_6482,N_6036);
and U6846 (N_6846,N_6071,N_6184);
or U6847 (N_6847,N_6320,N_6258);
and U6848 (N_6848,N_6192,N_6394);
and U6849 (N_6849,N_6028,N_6294);
nor U6850 (N_6850,N_6423,N_6443);
xor U6851 (N_6851,N_6250,N_6029);
and U6852 (N_6852,N_6399,N_6285);
nor U6853 (N_6853,N_6428,N_6362);
or U6854 (N_6854,N_6407,N_6108);
or U6855 (N_6855,N_6153,N_6317);
or U6856 (N_6856,N_6465,N_6191);
xor U6857 (N_6857,N_6408,N_6397);
nand U6858 (N_6858,N_6300,N_6194);
or U6859 (N_6859,N_6468,N_6420);
or U6860 (N_6860,N_6013,N_6054);
nand U6861 (N_6861,N_6278,N_6316);
xor U6862 (N_6862,N_6480,N_6301);
or U6863 (N_6863,N_6374,N_6336);
nand U6864 (N_6864,N_6476,N_6482);
nand U6865 (N_6865,N_6225,N_6039);
or U6866 (N_6866,N_6104,N_6343);
nand U6867 (N_6867,N_6142,N_6490);
nand U6868 (N_6868,N_6351,N_6105);
or U6869 (N_6869,N_6492,N_6223);
xor U6870 (N_6870,N_6005,N_6213);
xor U6871 (N_6871,N_6202,N_6142);
and U6872 (N_6872,N_6209,N_6016);
or U6873 (N_6873,N_6435,N_6388);
xnor U6874 (N_6874,N_6397,N_6486);
xor U6875 (N_6875,N_6040,N_6291);
and U6876 (N_6876,N_6251,N_6310);
xor U6877 (N_6877,N_6320,N_6001);
and U6878 (N_6878,N_6348,N_6440);
and U6879 (N_6879,N_6445,N_6180);
xnor U6880 (N_6880,N_6498,N_6175);
xor U6881 (N_6881,N_6051,N_6267);
nand U6882 (N_6882,N_6197,N_6423);
nor U6883 (N_6883,N_6041,N_6465);
nand U6884 (N_6884,N_6481,N_6334);
xnor U6885 (N_6885,N_6068,N_6364);
nor U6886 (N_6886,N_6158,N_6127);
xor U6887 (N_6887,N_6134,N_6116);
nor U6888 (N_6888,N_6331,N_6225);
or U6889 (N_6889,N_6350,N_6189);
and U6890 (N_6890,N_6166,N_6319);
and U6891 (N_6891,N_6042,N_6180);
and U6892 (N_6892,N_6065,N_6029);
nor U6893 (N_6893,N_6133,N_6250);
or U6894 (N_6894,N_6254,N_6127);
or U6895 (N_6895,N_6047,N_6178);
nand U6896 (N_6896,N_6072,N_6401);
nor U6897 (N_6897,N_6077,N_6221);
nand U6898 (N_6898,N_6426,N_6252);
or U6899 (N_6899,N_6258,N_6060);
nand U6900 (N_6900,N_6463,N_6377);
nand U6901 (N_6901,N_6476,N_6352);
xnor U6902 (N_6902,N_6470,N_6329);
nor U6903 (N_6903,N_6396,N_6318);
xnor U6904 (N_6904,N_6441,N_6047);
xnor U6905 (N_6905,N_6471,N_6463);
xnor U6906 (N_6906,N_6103,N_6327);
xnor U6907 (N_6907,N_6410,N_6037);
nor U6908 (N_6908,N_6301,N_6445);
or U6909 (N_6909,N_6423,N_6487);
nor U6910 (N_6910,N_6119,N_6208);
nor U6911 (N_6911,N_6173,N_6068);
nor U6912 (N_6912,N_6448,N_6476);
xor U6913 (N_6913,N_6362,N_6407);
or U6914 (N_6914,N_6062,N_6000);
nor U6915 (N_6915,N_6298,N_6410);
or U6916 (N_6916,N_6101,N_6429);
nor U6917 (N_6917,N_6092,N_6228);
and U6918 (N_6918,N_6369,N_6035);
and U6919 (N_6919,N_6401,N_6206);
nor U6920 (N_6920,N_6304,N_6069);
xnor U6921 (N_6921,N_6203,N_6105);
nor U6922 (N_6922,N_6194,N_6465);
nor U6923 (N_6923,N_6308,N_6252);
nor U6924 (N_6924,N_6081,N_6332);
nor U6925 (N_6925,N_6058,N_6450);
and U6926 (N_6926,N_6332,N_6209);
or U6927 (N_6927,N_6344,N_6150);
nand U6928 (N_6928,N_6490,N_6385);
nor U6929 (N_6929,N_6204,N_6408);
nand U6930 (N_6930,N_6300,N_6270);
nor U6931 (N_6931,N_6002,N_6482);
xor U6932 (N_6932,N_6077,N_6010);
nor U6933 (N_6933,N_6368,N_6191);
nor U6934 (N_6934,N_6162,N_6031);
nand U6935 (N_6935,N_6316,N_6291);
and U6936 (N_6936,N_6079,N_6312);
nor U6937 (N_6937,N_6058,N_6190);
and U6938 (N_6938,N_6185,N_6379);
xor U6939 (N_6939,N_6297,N_6383);
xor U6940 (N_6940,N_6065,N_6445);
xnor U6941 (N_6941,N_6408,N_6226);
or U6942 (N_6942,N_6476,N_6003);
and U6943 (N_6943,N_6097,N_6308);
or U6944 (N_6944,N_6098,N_6314);
xnor U6945 (N_6945,N_6491,N_6438);
or U6946 (N_6946,N_6024,N_6003);
nor U6947 (N_6947,N_6030,N_6195);
and U6948 (N_6948,N_6032,N_6155);
nand U6949 (N_6949,N_6156,N_6415);
nor U6950 (N_6950,N_6221,N_6277);
or U6951 (N_6951,N_6335,N_6276);
and U6952 (N_6952,N_6118,N_6092);
nand U6953 (N_6953,N_6314,N_6297);
and U6954 (N_6954,N_6428,N_6402);
nor U6955 (N_6955,N_6195,N_6335);
nor U6956 (N_6956,N_6237,N_6320);
nand U6957 (N_6957,N_6097,N_6029);
or U6958 (N_6958,N_6091,N_6432);
nor U6959 (N_6959,N_6286,N_6238);
xnor U6960 (N_6960,N_6024,N_6021);
or U6961 (N_6961,N_6377,N_6357);
and U6962 (N_6962,N_6189,N_6078);
nor U6963 (N_6963,N_6367,N_6095);
nor U6964 (N_6964,N_6098,N_6297);
xnor U6965 (N_6965,N_6221,N_6449);
and U6966 (N_6966,N_6161,N_6495);
nand U6967 (N_6967,N_6382,N_6335);
nand U6968 (N_6968,N_6273,N_6148);
nor U6969 (N_6969,N_6307,N_6284);
xnor U6970 (N_6970,N_6231,N_6007);
or U6971 (N_6971,N_6462,N_6465);
nor U6972 (N_6972,N_6384,N_6336);
nor U6973 (N_6973,N_6478,N_6055);
nand U6974 (N_6974,N_6106,N_6482);
nand U6975 (N_6975,N_6360,N_6084);
nand U6976 (N_6976,N_6063,N_6346);
and U6977 (N_6977,N_6360,N_6456);
or U6978 (N_6978,N_6248,N_6216);
and U6979 (N_6979,N_6396,N_6161);
xnor U6980 (N_6980,N_6348,N_6444);
or U6981 (N_6981,N_6127,N_6264);
xor U6982 (N_6982,N_6352,N_6011);
nor U6983 (N_6983,N_6351,N_6202);
or U6984 (N_6984,N_6314,N_6110);
nand U6985 (N_6985,N_6368,N_6091);
and U6986 (N_6986,N_6124,N_6249);
or U6987 (N_6987,N_6188,N_6013);
and U6988 (N_6988,N_6344,N_6441);
nor U6989 (N_6989,N_6182,N_6081);
nand U6990 (N_6990,N_6320,N_6112);
nand U6991 (N_6991,N_6050,N_6216);
nor U6992 (N_6992,N_6382,N_6033);
nor U6993 (N_6993,N_6132,N_6189);
xor U6994 (N_6994,N_6178,N_6393);
nand U6995 (N_6995,N_6232,N_6472);
xor U6996 (N_6996,N_6123,N_6181);
nand U6997 (N_6997,N_6237,N_6140);
and U6998 (N_6998,N_6232,N_6324);
or U6999 (N_6999,N_6319,N_6468);
and U7000 (N_7000,N_6987,N_6959);
and U7001 (N_7001,N_6800,N_6966);
nand U7002 (N_7002,N_6858,N_6843);
and U7003 (N_7003,N_6938,N_6955);
nor U7004 (N_7004,N_6517,N_6830);
nor U7005 (N_7005,N_6808,N_6538);
nand U7006 (N_7006,N_6905,N_6962);
nor U7007 (N_7007,N_6502,N_6529);
xnor U7008 (N_7008,N_6672,N_6571);
and U7009 (N_7009,N_6570,N_6591);
or U7010 (N_7010,N_6534,N_6573);
nor U7011 (N_7011,N_6688,N_6994);
xor U7012 (N_7012,N_6705,N_6741);
or U7013 (N_7013,N_6694,N_6971);
and U7014 (N_7014,N_6706,N_6684);
nor U7015 (N_7015,N_6539,N_6930);
xnor U7016 (N_7016,N_6977,N_6543);
nand U7017 (N_7017,N_6632,N_6578);
nand U7018 (N_7018,N_6968,N_6921);
and U7019 (N_7019,N_6649,N_6639);
nor U7020 (N_7020,N_6513,N_6895);
or U7021 (N_7021,N_6863,N_6546);
nor U7022 (N_7022,N_6730,N_6663);
xor U7023 (N_7023,N_6609,N_6923);
nand U7024 (N_7024,N_6714,N_6756);
and U7025 (N_7025,N_6960,N_6953);
nor U7026 (N_7026,N_6935,N_6658);
and U7027 (N_7027,N_6845,N_6715);
and U7028 (N_7028,N_6880,N_6695);
or U7029 (N_7029,N_6797,N_6877);
nand U7030 (N_7030,N_6666,N_6648);
or U7031 (N_7031,N_6854,N_6778);
or U7032 (N_7032,N_6656,N_6884);
nand U7033 (N_7033,N_6798,N_6941);
xor U7034 (N_7034,N_6561,N_6846);
or U7035 (N_7035,N_6844,N_6505);
nand U7036 (N_7036,N_6826,N_6541);
nor U7037 (N_7037,N_6693,N_6754);
or U7038 (N_7038,N_6547,N_6650);
and U7039 (N_7039,N_6725,N_6707);
or U7040 (N_7040,N_6833,N_6525);
and U7041 (N_7041,N_6631,N_6786);
nor U7042 (N_7042,N_6795,N_6755);
nand U7043 (N_7043,N_6532,N_6703);
and U7044 (N_7044,N_6601,N_6785);
nand U7045 (N_7045,N_6726,N_6992);
and U7046 (N_7046,N_6879,N_6788);
nor U7047 (N_7047,N_6524,N_6586);
nor U7048 (N_7048,N_6899,N_6767);
xnor U7049 (N_7049,N_6682,N_6668);
and U7050 (N_7050,N_6732,N_6629);
and U7051 (N_7051,N_6727,N_6881);
and U7052 (N_7052,N_6946,N_6906);
nor U7053 (N_7053,N_6516,N_6842);
nand U7054 (N_7054,N_6655,N_6796);
or U7055 (N_7055,N_6810,N_6821);
xnor U7056 (N_7056,N_6871,N_6780);
and U7057 (N_7057,N_6589,N_6885);
and U7058 (N_7058,N_6768,N_6604);
nor U7059 (N_7059,N_6592,N_6803);
nand U7060 (N_7060,N_6995,N_6948);
and U7061 (N_7061,N_6876,N_6851);
or U7062 (N_7062,N_6728,N_6990);
or U7063 (N_7063,N_6752,N_6642);
and U7064 (N_7064,N_6766,N_6550);
or U7065 (N_7065,N_6764,N_6908);
and U7066 (N_7066,N_6940,N_6646);
xor U7067 (N_7067,N_6974,N_6862);
nor U7068 (N_7068,N_6925,N_6951);
nor U7069 (N_7069,N_6818,N_6659);
xnor U7070 (N_7070,N_6594,N_6544);
xor U7071 (N_7071,N_6583,N_6961);
nand U7072 (N_7072,N_6520,N_6984);
nor U7073 (N_7073,N_6734,N_6912);
xor U7074 (N_7074,N_6619,N_6779);
or U7075 (N_7075,N_6782,N_6878);
xor U7076 (N_7076,N_6564,N_6548);
nand U7077 (N_7077,N_6852,N_6837);
xnor U7078 (N_7078,N_6620,N_6911);
and U7079 (N_7079,N_6893,N_6613);
xor U7080 (N_7080,N_6836,N_6986);
xor U7081 (N_7081,N_6552,N_6819);
xnor U7082 (N_7082,N_6676,N_6933);
nand U7083 (N_7083,N_6507,N_6860);
nand U7084 (N_7084,N_6892,N_6637);
xnor U7085 (N_7085,N_6612,N_6869);
xor U7086 (N_7086,N_6630,N_6643);
nand U7087 (N_7087,N_6874,N_6614);
nor U7088 (N_7088,N_6934,N_6508);
xnor U7089 (N_7089,N_6587,N_6518);
nand U7090 (N_7090,N_6735,N_6815);
nor U7091 (N_7091,N_6970,N_6944);
nor U7092 (N_7092,N_6920,N_6634);
nor U7093 (N_7093,N_6599,N_6989);
xor U7094 (N_7094,N_6673,N_6981);
and U7095 (N_7095,N_6719,N_6736);
or U7096 (N_7096,N_6793,N_6611);
nor U7097 (N_7097,N_6882,N_6608);
or U7098 (N_7098,N_6991,N_6825);
nand U7099 (N_7099,N_6914,N_6514);
nor U7100 (N_7100,N_6746,N_6685);
xor U7101 (N_7101,N_6555,N_6838);
and U7102 (N_7102,N_6551,N_6657);
nand U7103 (N_7103,N_6913,N_6849);
nand U7104 (N_7104,N_6771,N_6744);
and U7105 (N_7105,N_6985,N_6597);
xor U7106 (N_7106,N_6873,N_6813);
and U7107 (N_7107,N_6807,N_6679);
xnor U7108 (N_7108,N_6943,N_6500);
xor U7109 (N_7109,N_6824,N_6922);
nand U7110 (N_7110,N_6816,N_6698);
or U7111 (N_7111,N_6557,N_6531);
or U7112 (N_7112,N_6956,N_6641);
xnor U7113 (N_7113,N_6820,N_6605);
nor U7114 (N_7114,N_6806,N_6888);
nor U7115 (N_7115,N_6702,N_6841);
nor U7116 (N_7116,N_6776,N_6965);
and U7117 (N_7117,N_6640,N_6958);
and U7118 (N_7118,N_6758,N_6616);
nor U7119 (N_7119,N_6717,N_6804);
and U7120 (N_7120,N_6654,N_6638);
and U7121 (N_7121,N_6709,N_6848);
xnor U7122 (N_7122,N_6503,N_6568);
xnor U7123 (N_7123,N_6945,N_6652);
nand U7124 (N_7124,N_6540,N_6829);
xor U7125 (N_7125,N_6775,N_6929);
xor U7126 (N_7126,N_6670,N_6581);
xnor U7127 (N_7127,N_6853,N_6509);
or U7128 (N_7128,N_6542,N_6737);
nor U7129 (N_7129,N_6855,N_6661);
xnor U7130 (N_7130,N_6708,N_6566);
nand U7131 (N_7131,N_6753,N_6618);
nor U7132 (N_7132,N_6588,N_6926);
or U7133 (N_7133,N_6972,N_6950);
nor U7134 (N_7134,N_6867,N_6784);
and U7135 (N_7135,N_6856,N_6724);
nor U7136 (N_7136,N_6774,N_6748);
xor U7137 (N_7137,N_6954,N_6590);
and U7138 (N_7138,N_6939,N_6789);
nor U7139 (N_7139,N_6701,N_6665);
or U7140 (N_7140,N_6947,N_6901);
nand U7141 (N_7141,N_6680,N_6687);
xor U7142 (N_7142,N_6558,N_6691);
nand U7143 (N_7143,N_6577,N_6615);
nand U7144 (N_7144,N_6919,N_6569);
nand U7145 (N_7145,N_6560,N_6917);
nand U7146 (N_7146,N_6811,N_6553);
nand U7147 (N_7147,N_6580,N_6690);
nor U7148 (N_7148,N_6519,N_6689);
or U7149 (N_7149,N_6633,N_6750);
and U7150 (N_7150,N_6675,N_6743);
and U7151 (N_7151,N_6515,N_6562);
xnor U7152 (N_7152,N_6607,N_6565);
and U7153 (N_7153,N_6674,N_6868);
or U7154 (N_7154,N_6822,N_6533);
and U7155 (N_7155,N_6781,N_6624);
and U7156 (N_7156,N_6772,N_6567);
and U7157 (N_7157,N_6595,N_6898);
nor U7158 (N_7158,N_6904,N_6576);
nand U7159 (N_7159,N_6777,N_6678);
and U7160 (N_7160,N_6671,N_6857);
nor U7161 (N_7161,N_6769,N_6973);
or U7162 (N_7162,N_6890,N_6861);
xor U7163 (N_7163,N_6697,N_6739);
xor U7164 (N_7164,N_6909,N_6967);
xnor U7165 (N_7165,N_6745,N_6980);
xnor U7166 (N_7166,N_6765,N_6537);
nor U7167 (N_7167,N_6978,N_6713);
and U7168 (N_7168,N_6903,N_6790);
or U7169 (N_7169,N_6662,N_6626);
xnor U7170 (N_7170,N_6644,N_6692);
or U7171 (N_7171,N_6504,N_6621);
and U7172 (N_7172,N_6761,N_6681);
or U7173 (N_7173,N_6828,N_6850);
xor U7174 (N_7174,N_6827,N_6722);
nor U7175 (N_7175,N_6942,N_6832);
or U7176 (N_7176,N_6506,N_6927);
nand U7177 (N_7177,N_6596,N_6536);
xor U7178 (N_7178,N_6603,N_6924);
nor U7179 (N_7179,N_6501,N_6751);
nor U7180 (N_7180,N_6969,N_6907);
nand U7181 (N_7181,N_6928,N_6699);
and U7182 (N_7182,N_6902,N_6993);
or U7183 (N_7183,N_6647,N_6864);
and U7184 (N_7184,N_6653,N_6814);
xnor U7185 (N_7185,N_6636,N_6802);
and U7186 (N_7186,N_6559,N_6792);
or U7187 (N_7187,N_6606,N_6545);
and U7188 (N_7188,N_6686,N_6835);
xor U7189 (N_7189,N_6963,N_6817);
and U7190 (N_7190,N_6535,N_6711);
xnor U7191 (N_7191,N_6579,N_6982);
nand U7192 (N_7192,N_6875,N_6512);
nand U7193 (N_7193,N_6574,N_6593);
nand U7194 (N_7194,N_6932,N_6847);
or U7195 (N_7195,N_6530,N_6823);
xor U7196 (N_7196,N_6598,N_6770);
nand U7197 (N_7197,N_6975,N_6883);
or U7198 (N_7198,N_6582,N_6812);
or U7199 (N_7199,N_6872,N_6683);
and U7200 (N_7200,N_6976,N_6556);
nand U7201 (N_7201,N_6918,N_6840);
xnor U7202 (N_7202,N_6900,N_6602);
nand U7203 (N_7203,N_6738,N_6897);
xnor U7204 (N_7204,N_6910,N_6623);
nor U7205 (N_7205,N_6635,N_6996);
and U7206 (N_7206,N_6747,N_6763);
or U7207 (N_7207,N_6700,N_6510);
or U7208 (N_7208,N_6521,N_6891);
nor U7209 (N_7209,N_6526,N_6664);
nor U7210 (N_7210,N_6787,N_6740);
xor U7211 (N_7211,N_6600,N_6931);
nor U7212 (N_7212,N_6522,N_6894);
nand U7213 (N_7213,N_6669,N_6575);
nor U7214 (N_7214,N_6799,N_6896);
and U7215 (N_7215,N_6870,N_6622);
and U7216 (N_7216,N_6660,N_6957);
or U7217 (N_7217,N_6718,N_6723);
nand U7218 (N_7218,N_6617,N_6791);
nand U7219 (N_7219,N_6834,N_6527);
xor U7220 (N_7220,N_6645,N_6865);
nor U7221 (N_7221,N_6949,N_6887);
nor U7222 (N_7222,N_6937,N_6999);
nor U7223 (N_7223,N_6628,N_6859);
nand U7224 (N_7224,N_6528,N_6710);
and U7225 (N_7225,N_6983,N_6889);
nand U7226 (N_7226,N_6721,N_6762);
xnor U7227 (N_7227,N_6733,N_6801);
nand U7228 (N_7228,N_6677,N_6839);
xor U7229 (N_7229,N_6563,N_6805);
xnor U7230 (N_7230,N_6979,N_6964);
nor U7231 (N_7231,N_6759,N_6627);
xor U7232 (N_7232,N_6742,N_6783);
xor U7233 (N_7233,N_6831,N_6952);
or U7234 (N_7234,N_6794,N_6585);
nor U7235 (N_7235,N_6720,N_6809);
nor U7236 (N_7236,N_6625,N_6729);
and U7237 (N_7237,N_6731,N_6549);
nand U7238 (N_7238,N_6712,N_6584);
nand U7239 (N_7239,N_6523,N_6511);
nand U7240 (N_7240,N_6667,N_6716);
xnor U7241 (N_7241,N_6915,N_6773);
xor U7242 (N_7242,N_6610,N_6936);
or U7243 (N_7243,N_6749,N_6998);
xnor U7244 (N_7244,N_6572,N_6886);
nor U7245 (N_7245,N_6696,N_6757);
or U7246 (N_7246,N_6997,N_6866);
xnor U7247 (N_7247,N_6554,N_6651);
or U7248 (N_7248,N_6916,N_6760);
and U7249 (N_7249,N_6988,N_6704);
nand U7250 (N_7250,N_6735,N_6575);
and U7251 (N_7251,N_6699,N_6612);
xnor U7252 (N_7252,N_6930,N_6548);
or U7253 (N_7253,N_6519,N_6735);
or U7254 (N_7254,N_6592,N_6907);
xor U7255 (N_7255,N_6626,N_6535);
or U7256 (N_7256,N_6926,N_6962);
and U7257 (N_7257,N_6920,N_6530);
nand U7258 (N_7258,N_6751,N_6913);
xnor U7259 (N_7259,N_6594,N_6654);
xor U7260 (N_7260,N_6922,N_6623);
nor U7261 (N_7261,N_6717,N_6593);
and U7262 (N_7262,N_6866,N_6830);
or U7263 (N_7263,N_6830,N_6760);
nor U7264 (N_7264,N_6714,N_6557);
nand U7265 (N_7265,N_6575,N_6675);
nor U7266 (N_7266,N_6533,N_6560);
xnor U7267 (N_7267,N_6655,N_6500);
or U7268 (N_7268,N_6946,N_6950);
nor U7269 (N_7269,N_6868,N_6681);
xnor U7270 (N_7270,N_6524,N_6704);
nand U7271 (N_7271,N_6544,N_6699);
nand U7272 (N_7272,N_6830,N_6812);
nor U7273 (N_7273,N_6621,N_6998);
nand U7274 (N_7274,N_6689,N_6837);
xnor U7275 (N_7275,N_6858,N_6521);
xnor U7276 (N_7276,N_6930,N_6769);
or U7277 (N_7277,N_6870,N_6510);
nand U7278 (N_7278,N_6525,N_6845);
xnor U7279 (N_7279,N_6851,N_6956);
and U7280 (N_7280,N_6677,N_6734);
and U7281 (N_7281,N_6552,N_6662);
nor U7282 (N_7282,N_6511,N_6956);
xor U7283 (N_7283,N_6759,N_6673);
xor U7284 (N_7284,N_6729,N_6972);
or U7285 (N_7285,N_6970,N_6790);
xor U7286 (N_7286,N_6913,N_6556);
xnor U7287 (N_7287,N_6622,N_6520);
xor U7288 (N_7288,N_6536,N_6686);
and U7289 (N_7289,N_6833,N_6719);
nor U7290 (N_7290,N_6809,N_6791);
nand U7291 (N_7291,N_6922,N_6833);
nor U7292 (N_7292,N_6984,N_6794);
nor U7293 (N_7293,N_6874,N_6686);
or U7294 (N_7294,N_6772,N_6807);
nor U7295 (N_7295,N_6663,N_6521);
nand U7296 (N_7296,N_6952,N_6697);
and U7297 (N_7297,N_6955,N_6577);
nand U7298 (N_7298,N_6829,N_6634);
nor U7299 (N_7299,N_6562,N_6661);
nor U7300 (N_7300,N_6541,N_6520);
or U7301 (N_7301,N_6643,N_6985);
or U7302 (N_7302,N_6715,N_6919);
and U7303 (N_7303,N_6932,N_6641);
nand U7304 (N_7304,N_6904,N_6570);
or U7305 (N_7305,N_6599,N_6881);
and U7306 (N_7306,N_6707,N_6755);
and U7307 (N_7307,N_6998,N_6567);
nand U7308 (N_7308,N_6845,N_6520);
and U7309 (N_7309,N_6736,N_6779);
or U7310 (N_7310,N_6670,N_6551);
or U7311 (N_7311,N_6772,N_6948);
nand U7312 (N_7312,N_6703,N_6632);
nand U7313 (N_7313,N_6920,N_6915);
or U7314 (N_7314,N_6852,N_6611);
nor U7315 (N_7315,N_6832,N_6712);
nand U7316 (N_7316,N_6837,N_6817);
or U7317 (N_7317,N_6988,N_6857);
nor U7318 (N_7318,N_6880,N_6625);
nor U7319 (N_7319,N_6517,N_6684);
or U7320 (N_7320,N_6722,N_6552);
nand U7321 (N_7321,N_6986,N_6822);
xor U7322 (N_7322,N_6575,N_6931);
xor U7323 (N_7323,N_6779,N_6808);
and U7324 (N_7324,N_6769,N_6898);
nor U7325 (N_7325,N_6766,N_6993);
nand U7326 (N_7326,N_6678,N_6680);
and U7327 (N_7327,N_6637,N_6993);
or U7328 (N_7328,N_6853,N_6501);
nand U7329 (N_7329,N_6912,N_6568);
or U7330 (N_7330,N_6780,N_6730);
or U7331 (N_7331,N_6959,N_6729);
or U7332 (N_7332,N_6656,N_6559);
nor U7333 (N_7333,N_6755,N_6814);
nand U7334 (N_7334,N_6868,N_6700);
xnor U7335 (N_7335,N_6863,N_6763);
nor U7336 (N_7336,N_6780,N_6824);
nor U7337 (N_7337,N_6618,N_6925);
or U7338 (N_7338,N_6735,N_6800);
nand U7339 (N_7339,N_6639,N_6630);
nand U7340 (N_7340,N_6621,N_6594);
xor U7341 (N_7341,N_6990,N_6783);
xor U7342 (N_7342,N_6902,N_6782);
or U7343 (N_7343,N_6959,N_6518);
or U7344 (N_7344,N_6640,N_6523);
nor U7345 (N_7345,N_6668,N_6858);
and U7346 (N_7346,N_6709,N_6505);
nand U7347 (N_7347,N_6622,N_6683);
nand U7348 (N_7348,N_6651,N_6790);
nand U7349 (N_7349,N_6892,N_6760);
nand U7350 (N_7350,N_6962,N_6811);
xor U7351 (N_7351,N_6522,N_6879);
and U7352 (N_7352,N_6610,N_6691);
or U7353 (N_7353,N_6826,N_6611);
and U7354 (N_7354,N_6810,N_6613);
nor U7355 (N_7355,N_6537,N_6596);
and U7356 (N_7356,N_6909,N_6549);
nand U7357 (N_7357,N_6978,N_6648);
nor U7358 (N_7358,N_6970,N_6583);
xnor U7359 (N_7359,N_6606,N_6719);
or U7360 (N_7360,N_6509,N_6866);
nor U7361 (N_7361,N_6942,N_6512);
and U7362 (N_7362,N_6700,N_6716);
nand U7363 (N_7363,N_6854,N_6521);
nor U7364 (N_7364,N_6680,N_6918);
xor U7365 (N_7365,N_6722,N_6677);
and U7366 (N_7366,N_6514,N_6736);
or U7367 (N_7367,N_6922,N_6782);
nor U7368 (N_7368,N_6665,N_6730);
xnor U7369 (N_7369,N_6673,N_6855);
or U7370 (N_7370,N_6997,N_6816);
nand U7371 (N_7371,N_6993,N_6729);
xnor U7372 (N_7372,N_6965,N_6915);
and U7373 (N_7373,N_6635,N_6832);
and U7374 (N_7374,N_6842,N_6569);
xor U7375 (N_7375,N_6528,N_6818);
and U7376 (N_7376,N_6561,N_6524);
and U7377 (N_7377,N_6916,N_6742);
and U7378 (N_7378,N_6533,N_6938);
nor U7379 (N_7379,N_6924,N_6728);
nor U7380 (N_7380,N_6866,N_6843);
or U7381 (N_7381,N_6839,N_6877);
nand U7382 (N_7382,N_6594,N_6951);
or U7383 (N_7383,N_6561,N_6602);
nor U7384 (N_7384,N_6646,N_6731);
and U7385 (N_7385,N_6939,N_6784);
xor U7386 (N_7386,N_6658,N_6676);
or U7387 (N_7387,N_6869,N_6591);
nor U7388 (N_7388,N_6601,N_6907);
and U7389 (N_7389,N_6759,N_6769);
xor U7390 (N_7390,N_6556,N_6920);
nor U7391 (N_7391,N_6806,N_6773);
and U7392 (N_7392,N_6645,N_6939);
or U7393 (N_7393,N_6742,N_6609);
nand U7394 (N_7394,N_6799,N_6529);
nor U7395 (N_7395,N_6671,N_6710);
or U7396 (N_7396,N_6954,N_6716);
xnor U7397 (N_7397,N_6829,N_6933);
xnor U7398 (N_7398,N_6542,N_6668);
or U7399 (N_7399,N_6704,N_6580);
or U7400 (N_7400,N_6727,N_6775);
or U7401 (N_7401,N_6647,N_6829);
xnor U7402 (N_7402,N_6713,N_6968);
or U7403 (N_7403,N_6877,N_6981);
and U7404 (N_7404,N_6654,N_6549);
nor U7405 (N_7405,N_6580,N_6755);
xnor U7406 (N_7406,N_6721,N_6975);
xor U7407 (N_7407,N_6822,N_6545);
nor U7408 (N_7408,N_6559,N_6721);
nor U7409 (N_7409,N_6613,N_6945);
xor U7410 (N_7410,N_6630,N_6948);
or U7411 (N_7411,N_6942,N_6810);
nor U7412 (N_7412,N_6657,N_6618);
nand U7413 (N_7413,N_6585,N_6506);
xnor U7414 (N_7414,N_6659,N_6927);
nand U7415 (N_7415,N_6778,N_6527);
nor U7416 (N_7416,N_6944,N_6982);
xor U7417 (N_7417,N_6731,N_6619);
or U7418 (N_7418,N_6719,N_6901);
nor U7419 (N_7419,N_6618,N_6892);
nand U7420 (N_7420,N_6788,N_6725);
nor U7421 (N_7421,N_6979,N_6809);
nand U7422 (N_7422,N_6935,N_6535);
nor U7423 (N_7423,N_6534,N_6952);
nand U7424 (N_7424,N_6647,N_6581);
or U7425 (N_7425,N_6683,N_6893);
nor U7426 (N_7426,N_6908,N_6721);
or U7427 (N_7427,N_6796,N_6556);
nor U7428 (N_7428,N_6802,N_6788);
xor U7429 (N_7429,N_6517,N_6580);
xor U7430 (N_7430,N_6873,N_6608);
and U7431 (N_7431,N_6584,N_6542);
nand U7432 (N_7432,N_6984,N_6920);
nand U7433 (N_7433,N_6836,N_6904);
nor U7434 (N_7434,N_6780,N_6992);
or U7435 (N_7435,N_6865,N_6766);
xnor U7436 (N_7436,N_6563,N_6973);
or U7437 (N_7437,N_6996,N_6573);
and U7438 (N_7438,N_6847,N_6742);
xnor U7439 (N_7439,N_6960,N_6781);
nand U7440 (N_7440,N_6585,N_6904);
and U7441 (N_7441,N_6867,N_6592);
xnor U7442 (N_7442,N_6957,N_6972);
or U7443 (N_7443,N_6717,N_6641);
or U7444 (N_7444,N_6587,N_6796);
xor U7445 (N_7445,N_6669,N_6971);
or U7446 (N_7446,N_6773,N_6942);
xor U7447 (N_7447,N_6717,N_6600);
and U7448 (N_7448,N_6552,N_6542);
xor U7449 (N_7449,N_6736,N_6834);
nor U7450 (N_7450,N_6925,N_6916);
nor U7451 (N_7451,N_6846,N_6571);
and U7452 (N_7452,N_6798,N_6822);
nor U7453 (N_7453,N_6973,N_6765);
and U7454 (N_7454,N_6622,N_6958);
or U7455 (N_7455,N_6708,N_6951);
nand U7456 (N_7456,N_6631,N_6612);
or U7457 (N_7457,N_6605,N_6537);
or U7458 (N_7458,N_6544,N_6585);
nor U7459 (N_7459,N_6770,N_6540);
and U7460 (N_7460,N_6639,N_6631);
or U7461 (N_7461,N_6607,N_6680);
nand U7462 (N_7462,N_6795,N_6689);
xnor U7463 (N_7463,N_6644,N_6927);
nand U7464 (N_7464,N_6876,N_6501);
xnor U7465 (N_7465,N_6546,N_6989);
or U7466 (N_7466,N_6514,N_6797);
and U7467 (N_7467,N_6942,N_6524);
xnor U7468 (N_7468,N_6720,N_6568);
and U7469 (N_7469,N_6994,N_6596);
or U7470 (N_7470,N_6910,N_6554);
and U7471 (N_7471,N_6518,N_6972);
and U7472 (N_7472,N_6828,N_6674);
or U7473 (N_7473,N_6653,N_6562);
xnor U7474 (N_7474,N_6874,N_6591);
nor U7475 (N_7475,N_6502,N_6752);
or U7476 (N_7476,N_6643,N_6967);
or U7477 (N_7477,N_6878,N_6580);
or U7478 (N_7478,N_6602,N_6667);
and U7479 (N_7479,N_6977,N_6507);
nand U7480 (N_7480,N_6518,N_6680);
xor U7481 (N_7481,N_6665,N_6663);
xnor U7482 (N_7482,N_6977,N_6546);
nand U7483 (N_7483,N_6633,N_6962);
or U7484 (N_7484,N_6907,N_6643);
nand U7485 (N_7485,N_6700,N_6808);
nand U7486 (N_7486,N_6988,N_6896);
nand U7487 (N_7487,N_6576,N_6796);
nor U7488 (N_7488,N_6637,N_6879);
nand U7489 (N_7489,N_6717,N_6892);
and U7490 (N_7490,N_6956,N_6758);
and U7491 (N_7491,N_6789,N_6924);
xor U7492 (N_7492,N_6773,N_6686);
nor U7493 (N_7493,N_6751,N_6861);
nand U7494 (N_7494,N_6527,N_6571);
or U7495 (N_7495,N_6940,N_6565);
nand U7496 (N_7496,N_6757,N_6657);
and U7497 (N_7497,N_6878,N_6531);
nor U7498 (N_7498,N_6510,N_6629);
xor U7499 (N_7499,N_6583,N_6700);
and U7500 (N_7500,N_7153,N_7448);
or U7501 (N_7501,N_7087,N_7417);
and U7502 (N_7502,N_7062,N_7030);
nor U7503 (N_7503,N_7262,N_7124);
nor U7504 (N_7504,N_7101,N_7036);
nand U7505 (N_7505,N_7435,N_7080);
nor U7506 (N_7506,N_7477,N_7068);
nand U7507 (N_7507,N_7076,N_7228);
and U7508 (N_7508,N_7260,N_7014);
nand U7509 (N_7509,N_7466,N_7467);
or U7510 (N_7510,N_7147,N_7471);
or U7511 (N_7511,N_7067,N_7016);
xor U7512 (N_7512,N_7055,N_7148);
nand U7513 (N_7513,N_7495,N_7059);
or U7514 (N_7514,N_7395,N_7180);
or U7515 (N_7515,N_7399,N_7490);
or U7516 (N_7516,N_7378,N_7116);
nand U7517 (N_7517,N_7052,N_7363);
nor U7518 (N_7518,N_7374,N_7447);
and U7519 (N_7519,N_7420,N_7294);
nand U7520 (N_7520,N_7176,N_7119);
or U7521 (N_7521,N_7008,N_7201);
nor U7522 (N_7522,N_7379,N_7137);
xor U7523 (N_7523,N_7430,N_7078);
nand U7524 (N_7524,N_7145,N_7332);
nor U7525 (N_7525,N_7449,N_7309);
or U7526 (N_7526,N_7488,N_7348);
xor U7527 (N_7527,N_7326,N_7292);
and U7528 (N_7528,N_7286,N_7405);
xnor U7529 (N_7529,N_7172,N_7084);
and U7530 (N_7530,N_7088,N_7383);
and U7531 (N_7531,N_7433,N_7413);
nand U7532 (N_7532,N_7476,N_7419);
nor U7533 (N_7533,N_7327,N_7194);
and U7534 (N_7534,N_7250,N_7375);
and U7535 (N_7535,N_7110,N_7209);
nor U7536 (N_7536,N_7173,N_7469);
nand U7537 (N_7537,N_7491,N_7229);
nor U7538 (N_7538,N_7425,N_7158);
or U7539 (N_7539,N_7489,N_7044);
xor U7540 (N_7540,N_7114,N_7482);
or U7541 (N_7541,N_7261,N_7445);
or U7542 (N_7542,N_7112,N_7093);
nor U7543 (N_7543,N_7269,N_7351);
and U7544 (N_7544,N_7031,N_7219);
or U7545 (N_7545,N_7174,N_7095);
nor U7546 (N_7546,N_7142,N_7025);
nor U7547 (N_7547,N_7352,N_7057);
or U7548 (N_7548,N_7451,N_7224);
xnor U7549 (N_7549,N_7480,N_7325);
and U7550 (N_7550,N_7240,N_7434);
and U7551 (N_7551,N_7129,N_7072);
nand U7552 (N_7552,N_7429,N_7086);
or U7553 (N_7553,N_7313,N_7151);
or U7554 (N_7554,N_7299,N_7296);
nand U7555 (N_7555,N_7013,N_7077);
nor U7556 (N_7556,N_7233,N_7499);
or U7557 (N_7557,N_7321,N_7456);
or U7558 (N_7558,N_7431,N_7333);
or U7559 (N_7559,N_7081,N_7226);
and U7560 (N_7560,N_7054,N_7318);
xor U7561 (N_7561,N_7028,N_7270);
nand U7562 (N_7562,N_7190,N_7006);
xnor U7563 (N_7563,N_7130,N_7439);
or U7564 (N_7564,N_7497,N_7272);
or U7565 (N_7565,N_7322,N_7310);
and U7566 (N_7566,N_7422,N_7002);
xnor U7567 (N_7567,N_7376,N_7097);
xor U7568 (N_7568,N_7104,N_7335);
nor U7569 (N_7569,N_7302,N_7493);
and U7570 (N_7570,N_7303,N_7381);
or U7571 (N_7571,N_7218,N_7312);
nor U7572 (N_7572,N_7152,N_7045);
nand U7573 (N_7573,N_7017,N_7196);
and U7574 (N_7574,N_7336,N_7274);
nand U7575 (N_7575,N_7266,N_7401);
and U7576 (N_7576,N_7195,N_7191);
xor U7577 (N_7577,N_7392,N_7126);
nor U7578 (N_7578,N_7049,N_7367);
nor U7579 (N_7579,N_7166,N_7100);
xnor U7580 (N_7580,N_7212,N_7406);
or U7581 (N_7581,N_7438,N_7139);
xnor U7582 (N_7582,N_7217,N_7001);
xnor U7583 (N_7583,N_7092,N_7107);
xnor U7584 (N_7584,N_7026,N_7307);
nor U7585 (N_7585,N_7103,N_7213);
nor U7586 (N_7586,N_7056,N_7342);
nand U7587 (N_7587,N_7027,N_7064);
nand U7588 (N_7588,N_7205,N_7181);
nor U7589 (N_7589,N_7208,N_7221);
xor U7590 (N_7590,N_7178,N_7366);
and U7591 (N_7591,N_7436,N_7105);
xnor U7592 (N_7592,N_7353,N_7115);
nor U7593 (N_7593,N_7437,N_7127);
nor U7594 (N_7594,N_7284,N_7047);
or U7595 (N_7595,N_7005,N_7177);
nor U7596 (N_7596,N_7404,N_7323);
and U7597 (N_7597,N_7365,N_7023);
or U7598 (N_7598,N_7029,N_7470);
nor U7599 (N_7599,N_7271,N_7192);
nand U7600 (N_7600,N_7423,N_7082);
or U7601 (N_7601,N_7046,N_7458);
or U7602 (N_7602,N_7400,N_7133);
and U7603 (N_7603,N_7403,N_7004);
nand U7604 (N_7604,N_7215,N_7360);
and U7605 (N_7605,N_7037,N_7349);
nor U7606 (N_7606,N_7305,N_7009);
or U7607 (N_7607,N_7328,N_7258);
and U7608 (N_7608,N_7492,N_7278);
and U7609 (N_7609,N_7454,N_7069);
nor U7610 (N_7610,N_7242,N_7199);
nand U7611 (N_7611,N_7356,N_7239);
xor U7612 (N_7612,N_7032,N_7441);
nand U7613 (N_7613,N_7314,N_7169);
nand U7614 (N_7614,N_7019,N_7264);
and U7615 (N_7615,N_7234,N_7143);
nand U7616 (N_7616,N_7020,N_7065);
or U7617 (N_7617,N_7163,N_7243);
or U7618 (N_7618,N_7184,N_7478);
nand U7619 (N_7619,N_7164,N_7308);
nand U7620 (N_7620,N_7334,N_7474);
and U7621 (N_7621,N_7397,N_7039);
xnor U7622 (N_7622,N_7263,N_7295);
nand U7623 (N_7623,N_7079,N_7085);
or U7624 (N_7624,N_7007,N_7157);
xor U7625 (N_7625,N_7227,N_7074);
or U7626 (N_7626,N_7200,N_7198);
xnor U7627 (N_7627,N_7123,N_7135);
xor U7628 (N_7628,N_7455,N_7304);
and U7629 (N_7629,N_7280,N_7207);
or U7630 (N_7630,N_7254,N_7149);
nand U7631 (N_7631,N_7255,N_7186);
nor U7632 (N_7632,N_7113,N_7387);
nor U7633 (N_7633,N_7090,N_7109);
xor U7634 (N_7634,N_7483,N_7222);
nor U7635 (N_7635,N_7211,N_7315);
nor U7636 (N_7636,N_7393,N_7160);
nand U7637 (N_7637,N_7398,N_7033);
and U7638 (N_7638,N_7364,N_7232);
nor U7639 (N_7639,N_7389,N_7414);
nand U7640 (N_7640,N_7377,N_7183);
nand U7641 (N_7641,N_7236,N_7358);
or U7642 (N_7642,N_7410,N_7144);
or U7643 (N_7643,N_7098,N_7121);
nand U7644 (N_7644,N_7380,N_7385);
or U7645 (N_7645,N_7111,N_7141);
nor U7646 (N_7646,N_7346,N_7457);
nor U7647 (N_7647,N_7247,N_7345);
nand U7648 (N_7648,N_7179,N_7070);
nand U7649 (N_7649,N_7287,N_7073);
and U7650 (N_7650,N_7132,N_7216);
xnor U7651 (N_7651,N_7409,N_7317);
or U7652 (N_7652,N_7096,N_7462);
xor U7653 (N_7653,N_7369,N_7257);
or U7654 (N_7654,N_7288,N_7165);
xnor U7655 (N_7655,N_7300,N_7391);
and U7656 (N_7656,N_7094,N_7162);
nand U7657 (N_7657,N_7464,N_7161);
nor U7658 (N_7658,N_7155,N_7343);
and U7659 (N_7659,N_7331,N_7248);
xor U7660 (N_7660,N_7443,N_7220);
nor U7661 (N_7661,N_7000,N_7265);
nand U7662 (N_7662,N_7102,N_7170);
nor U7663 (N_7663,N_7244,N_7426);
or U7664 (N_7664,N_7235,N_7089);
or U7665 (N_7665,N_7256,N_7370);
nor U7666 (N_7666,N_7418,N_7018);
and U7667 (N_7667,N_7320,N_7485);
nand U7668 (N_7668,N_7463,N_7408);
and U7669 (N_7669,N_7117,N_7498);
xnor U7670 (N_7670,N_7128,N_7075);
nor U7671 (N_7671,N_7486,N_7035);
nor U7672 (N_7672,N_7246,N_7416);
and U7673 (N_7673,N_7187,N_7060);
nor U7674 (N_7674,N_7440,N_7231);
xor U7675 (N_7675,N_7118,N_7051);
and U7676 (N_7676,N_7204,N_7230);
or U7677 (N_7677,N_7021,N_7249);
or U7678 (N_7678,N_7341,N_7290);
xor U7679 (N_7679,N_7040,N_7010);
nor U7680 (N_7680,N_7193,N_7459);
xor U7681 (N_7681,N_7197,N_7063);
or U7682 (N_7682,N_7347,N_7238);
and U7683 (N_7683,N_7159,N_7394);
nor U7684 (N_7684,N_7042,N_7282);
and U7685 (N_7685,N_7267,N_7338);
nand U7686 (N_7686,N_7131,N_7481);
nand U7687 (N_7687,N_7468,N_7146);
nor U7688 (N_7688,N_7122,N_7460);
and U7689 (N_7689,N_7245,N_7202);
xnor U7690 (N_7690,N_7275,N_7253);
nand U7691 (N_7691,N_7273,N_7182);
and U7692 (N_7692,N_7106,N_7214);
and U7693 (N_7693,N_7427,N_7337);
or U7694 (N_7694,N_7024,N_7472);
nand U7695 (N_7695,N_7283,N_7461);
nand U7696 (N_7696,N_7138,N_7411);
xor U7697 (N_7697,N_7407,N_7034);
xor U7698 (N_7698,N_7357,N_7362);
or U7699 (N_7699,N_7251,N_7268);
xor U7700 (N_7700,N_7339,N_7277);
or U7701 (N_7701,N_7237,N_7354);
or U7702 (N_7702,N_7125,N_7175);
xor U7703 (N_7703,N_7048,N_7297);
or U7704 (N_7704,N_7371,N_7446);
nand U7705 (N_7705,N_7140,N_7453);
or U7706 (N_7706,N_7091,N_7487);
or U7707 (N_7707,N_7324,N_7421);
nand U7708 (N_7708,N_7120,N_7099);
nor U7709 (N_7709,N_7071,N_7412);
xor U7710 (N_7710,N_7452,N_7390);
or U7711 (N_7711,N_7344,N_7289);
nand U7712 (N_7712,N_7465,N_7210);
or U7713 (N_7713,N_7373,N_7276);
nand U7714 (N_7714,N_7311,N_7150);
or U7715 (N_7715,N_7285,N_7306);
nor U7716 (N_7716,N_7134,N_7038);
and U7717 (N_7717,N_7361,N_7444);
xnor U7718 (N_7718,N_7223,N_7279);
nand U7719 (N_7719,N_7428,N_7043);
nand U7720 (N_7720,N_7494,N_7372);
nand U7721 (N_7721,N_7396,N_7022);
nand U7722 (N_7722,N_7066,N_7156);
or U7723 (N_7723,N_7203,N_7359);
and U7724 (N_7724,N_7473,N_7241);
xnor U7725 (N_7725,N_7189,N_7058);
nor U7726 (N_7726,N_7496,N_7432);
or U7727 (N_7727,N_7050,N_7061);
nand U7728 (N_7728,N_7136,N_7329);
nand U7729 (N_7729,N_7167,N_7154);
and U7730 (N_7730,N_7368,N_7185);
and U7731 (N_7731,N_7291,N_7188);
nor U7732 (N_7732,N_7424,N_7384);
nand U7733 (N_7733,N_7316,N_7252);
and U7734 (N_7734,N_7003,N_7298);
nand U7735 (N_7735,N_7402,N_7293);
and U7736 (N_7736,N_7484,N_7168);
nor U7737 (N_7737,N_7442,N_7281);
nor U7738 (N_7738,N_7475,N_7330);
xnor U7739 (N_7739,N_7108,N_7171);
or U7740 (N_7740,N_7301,N_7083);
or U7741 (N_7741,N_7350,N_7415);
nor U7742 (N_7742,N_7011,N_7206);
nor U7743 (N_7743,N_7386,N_7479);
xnor U7744 (N_7744,N_7319,N_7259);
and U7745 (N_7745,N_7053,N_7041);
and U7746 (N_7746,N_7355,N_7382);
nor U7747 (N_7747,N_7012,N_7015);
xor U7748 (N_7748,N_7340,N_7225);
nor U7749 (N_7749,N_7388,N_7450);
nand U7750 (N_7750,N_7276,N_7321);
nand U7751 (N_7751,N_7291,N_7059);
nand U7752 (N_7752,N_7308,N_7455);
nand U7753 (N_7753,N_7164,N_7176);
xor U7754 (N_7754,N_7102,N_7026);
or U7755 (N_7755,N_7205,N_7167);
or U7756 (N_7756,N_7162,N_7178);
xnor U7757 (N_7757,N_7072,N_7179);
xor U7758 (N_7758,N_7460,N_7289);
nand U7759 (N_7759,N_7243,N_7140);
nand U7760 (N_7760,N_7414,N_7271);
and U7761 (N_7761,N_7235,N_7184);
or U7762 (N_7762,N_7038,N_7196);
or U7763 (N_7763,N_7057,N_7330);
and U7764 (N_7764,N_7036,N_7053);
and U7765 (N_7765,N_7326,N_7033);
nor U7766 (N_7766,N_7126,N_7377);
or U7767 (N_7767,N_7209,N_7406);
nand U7768 (N_7768,N_7329,N_7301);
nand U7769 (N_7769,N_7037,N_7271);
and U7770 (N_7770,N_7078,N_7114);
nand U7771 (N_7771,N_7273,N_7486);
nand U7772 (N_7772,N_7207,N_7215);
or U7773 (N_7773,N_7154,N_7454);
or U7774 (N_7774,N_7425,N_7311);
and U7775 (N_7775,N_7431,N_7149);
nor U7776 (N_7776,N_7401,N_7279);
and U7777 (N_7777,N_7446,N_7208);
xnor U7778 (N_7778,N_7105,N_7135);
or U7779 (N_7779,N_7498,N_7143);
nor U7780 (N_7780,N_7322,N_7235);
nor U7781 (N_7781,N_7395,N_7177);
or U7782 (N_7782,N_7124,N_7186);
nand U7783 (N_7783,N_7057,N_7276);
nand U7784 (N_7784,N_7154,N_7413);
or U7785 (N_7785,N_7282,N_7495);
and U7786 (N_7786,N_7220,N_7354);
or U7787 (N_7787,N_7179,N_7400);
nand U7788 (N_7788,N_7111,N_7494);
nand U7789 (N_7789,N_7493,N_7070);
or U7790 (N_7790,N_7274,N_7217);
and U7791 (N_7791,N_7475,N_7013);
or U7792 (N_7792,N_7238,N_7072);
or U7793 (N_7793,N_7232,N_7489);
nand U7794 (N_7794,N_7345,N_7297);
nor U7795 (N_7795,N_7219,N_7026);
or U7796 (N_7796,N_7031,N_7181);
xnor U7797 (N_7797,N_7488,N_7478);
or U7798 (N_7798,N_7009,N_7395);
xnor U7799 (N_7799,N_7129,N_7346);
xor U7800 (N_7800,N_7430,N_7321);
xnor U7801 (N_7801,N_7042,N_7465);
nor U7802 (N_7802,N_7221,N_7035);
and U7803 (N_7803,N_7068,N_7221);
nand U7804 (N_7804,N_7035,N_7151);
nor U7805 (N_7805,N_7293,N_7449);
nand U7806 (N_7806,N_7024,N_7091);
nand U7807 (N_7807,N_7372,N_7275);
and U7808 (N_7808,N_7034,N_7350);
nand U7809 (N_7809,N_7205,N_7042);
nor U7810 (N_7810,N_7174,N_7198);
nand U7811 (N_7811,N_7423,N_7020);
or U7812 (N_7812,N_7467,N_7181);
or U7813 (N_7813,N_7383,N_7337);
xnor U7814 (N_7814,N_7196,N_7413);
and U7815 (N_7815,N_7424,N_7188);
or U7816 (N_7816,N_7251,N_7099);
nor U7817 (N_7817,N_7364,N_7185);
xnor U7818 (N_7818,N_7158,N_7393);
nor U7819 (N_7819,N_7071,N_7097);
xor U7820 (N_7820,N_7467,N_7311);
nor U7821 (N_7821,N_7250,N_7464);
and U7822 (N_7822,N_7049,N_7446);
nor U7823 (N_7823,N_7261,N_7437);
nor U7824 (N_7824,N_7212,N_7281);
nor U7825 (N_7825,N_7319,N_7152);
xnor U7826 (N_7826,N_7452,N_7388);
xor U7827 (N_7827,N_7473,N_7209);
nand U7828 (N_7828,N_7114,N_7359);
nand U7829 (N_7829,N_7075,N_7385);
nor U7830 (N_7830,N_7363,N_7482);
or U7831 (N_7831,N_7227,N_7478);
nor U7832 (N_7832,N_7455,N_7433);
nand U7833 (N_7833,N_7117,N_7404);
nor U7834 (N_7834,N_7189,N_7209);
xor U7835 (N_7835,N_7224,N_7124);
nor U7836 (N_7836,N_7038,N_7107);
and U7837 (N_7837,N_7229,N_7273);
xnor U7838 (N_7838,N_7363,N_7094);
xnor U7839 (N_7839,N_7195,N_7076);
xor U7840 (N_7840,N_7480,N_7395);
xnor U7841 (N_7841,N_7481,N_7017);
xnor U7842 (N_7842,N_7181,N_7476);
nor U7843 (N_7843,N_7307,N_7126);
xnor U7844 (N_7844,N_7341,N_7214);
nor U7845 (N_7845,N_7238,N_7102);
nor U7846 (N_7846,N_7019,N_7208);
nand U7847 (N_7847,N_7323,N_7225);
nor U7848 (N_7848,N_7229,N_7282);
and U7849 (N_7849,N_7492,N_7350);
or U7850 (N_7850,N_7311,N_7219);
nand U7851 (N_7851,N_7059,N_7394);
and U7852 (N_7852,N_7170,N_7464);
xor U7853 (N_7853,N_7142,N_7108);
xor U7854 (N_7854,N_7248,N_7137);
xor U7855 (N_7855,N_7328,N_7262);
xor U7856 (N_7856,N_7122,N_7456);
xor U7857 (N_7857,N_7466,N_7453);
nand U7858 (N_7858,N_7222,N_7043);
or U7859 (N_7859,N_7242,N_7043);
xor U7860 (N_7860,N_7234,N_7401);
nand U7861 (N_7861,N_7230,N_7127);
and U7862 (N_7862,N_7377,N_7089);
nor U7863 (N_7863,N_7096,N_7129);
or U7864 (N_7864,N_7365,N_7469);
and U7865 (N_7865,N_7397,N_7192);
xnor U7866 (N_7866,N_7250,N_7472);
xor U7867 (N_7867,N_7073,N_7305);
nand U7868 (N_7868,N_7382,N_7096);
nand U7869 (N_7869,N_7495,N_7358);
nor U7870 (N_7870,N_7315,N_7069);
and U7871 (N_7871,N_7480,N_7361);
or U7872 (N_7872,N_7161,N_7013);
and U7873 (N_7873,N_7365,N_7186);
and U7874 (N_7874,N_7001,N_7011);
nand U7875 (N_7875,N_7305,N_7191);
nor U7876 (N_7876,N_7092,N_7313);
nand U7877 (N_7877,N_7315,N_7182);
or U7878 (N_7878,N_7045,N_7019);
nor U7879 (N_7879,N_7499,N_7478);
xnor U7880 (N_7880,N_7430,N_7437);
nor U7881 (N_7881,N_7100,N_7002);
nor U7882 (N_7882,N_7037,N_7259);
and U7883 (N_7883,N_7129,N_7447);
nor U7884 (N_7884,N_7208,N_7487);
nand U7885 (N_7885,N_7121,N_7329);
or U7886 (N_7886,N_7202,N_7007);
nand U7887 (N_7887,N_7138,N_7134);
xnor U7888 (N_7888,N_7495,N_7353);
and U7889 (N_7889,N_7244,N_7102);
nor U7890 (N_7890,N_7168,N_7086);
or U7891 (N_7891,N_7046,N_7101);
xnor U7892 (N_7892,N_7165,N_7325);
nand U7893 (N_7893,N_7174,N_7053);
xnor U7894 (N_7894,N_7123,N_7082);
and U7895 (N_7895,N_7199,N_7009);
nor U7896 (N_7896,N_7209,N_7239);
nand U7897 (N_7897,N_7029,N_7283);
and U7898 (N_7898,N_7309,N_7194);
xor U7899 (N_7899,N_7207,N_7413);
and U7900 (N_7900,N_7238,N_7234);
xnor U7901 (N_7901,N_7471,N_7460);
nor U7902 (N_7902,N_7293,N_7008);
nand U7903 (N_7903,N_7238,N_7248);
xnor U7904 (N_7904,N_7280,N_7130);
nor U7905 (N_7905,N_7020,N_7188);
nor U7906 (N_7906,N_7449,N_7415);
nand U7907 (N_7907,N_7403,N_7119);
xnor U7908 (N_7908,N_7145,N_7264);
nor U7909 (N_7909,N_7198,N_7105);
nand U7910 (N_7910,N_7489,N_7462);
or U7911 (N_7911,N_7007,N_7054);
nand U7912 (N_7912,N_7181,N_7210);
and U7913 (N_7913,N_7430,N_7375);
and U7914 (N_7914,N_7401,N_7047);
nor U7915 (N_7915,N_7458,N_7179);
nand U7916 (N_7916,N_7284,N_7499);
xnor U7917 (N_7917,N_7003,N_7246);
xnor U7918 (N_7918,N_7047,N_7182);
nor U7919 (N_7919,N_7473,N_7089);
xor U7920 (N_7920,N_7323,N_7215);
xor U7921 (N_7921,N_7461,N_7280);
nor U7922 (N_7922,N_7047,N_7449);
and U7923 (N_7923,N_7158,N_7325);
and U7924 (N_7924,N_7359,N_7174);
or U7925 (N_7925,N_7358,N_7117);
xor U7926 (N_7926,N_7194,N_7381);
xnor U7927 (N_7927,N_7176,N_7253);
xnor U7928 (N_7928,N_7409,N_7255);
or U7929 (N_7929,N_7426,N_7071);
and U7930 (N_7930,N_7451,N_7218);
and U7931 (N_7931,N_7362,N_7240);
nor U7932 (N_7932,N_7294,N_7433);
or U7933 (N_7933,N_7450,N_7285);
nand U7934 (N_7934,N_7401,N_7235);
nand U7935 (N_7935,N_7125,N_7177);
and U7936 (N_7936,N_7293,N_7371);
and U7937 (N_7937,N_7124,N_7094);
nand U7938 (N_7938,N_7312,N_7403);
nand U7939 (N_7939,N_7374,N_7445);
nand U7940 (N_7940,N_7052,N_7291);
and U7941 (N_7941,N_7119,N_7301);
nor U7942 (N_7942,N_7249,N_7020);
or U7943 (N_7943,N_7346,N_7226);
nand U7944 (N_7944,N_7129,N_7154);
nand U7945 (N_7945,N_7300,N_7382);
nand U7946 (N_7946,N_7462,N_7479);
nand U7947 (N_7947,N_7258,N_7297);
nand U7948 (N_7948,N_7413,N_7361);
or U7949 (N_7949,N_7094,N_7159);
nand U7950 (N_7950,N_7028,N_7426);
xnor U7951 (N_7951,N_7235,N_7051);
xnor U7952 (N_7952,N_7432,N_7214);
nor U7953 (N_7953,N_7297,N_7152);
nand U7954 (N_7954,N_7394,N_7389);
or U7955 (N_7955,N_7062,N_7389);
xnor U7956 (N_7956,N_7219,N_7426);
nand U7957 (N_7957,N_7266,N_7303);
and U7958 (N_7958,N_7362,N_7349);
nand U7959 (N_7959,N_7152,N_7149);
or U7960 (N_7960,N_7003,N_7056);
and U7961 (N_7961,N_7190,N_7479);
and U7962 (N_7962,N_7452,N_7406);
and U7963 (N_7963,N_7228,N_7391);
or U7964 (N_7964,N_7196,N_7498);
or U7965 (N_7965,N_7107,N_7216);
or U7966 (N_7966,N_7418,N_7173);
and U7967 (N_7967,N_7216,N_7361);
xnor U7968 (N_7968,N_7057,N_7265);
nor U7969 (N_7969,N_7086,N_7443);
and U7970 (N_7970,N_7414,N_7285);
nand U7971 (N_7971,N_7145,N_7330);
and U7972 (N_7972,N_7209,N_7131);
or U7973 (N_7973,N_7406,N_7203);
or U7974 (N_7974,N_7190,N_7312);
or U7975 (N_7975,N_7456,N_7342);
nor U7976 (N_7976,N_7092,N_7036);
or U7977 (N_7977,N_7183,N_7389);
nor U7978 (N_7978,N_7454,N_7291);
nor U7979 (N_7979,N_7277,N_7409);
nor U7980 (N_7980,N_7438,N_7454);
and U7981 (N_7981,N_7176,N_7429);
nor U7982 (N_7982,N_7345,N_7045);
nor U7983 (N_7983,N_7085,N_7393);
or U7984 (N_7984,N_7069,N_7133);
nand U7985 (N_7985,N_7316,N_7157);
and U7986 (N_7986,N_7208,N_7379);
nand U7987 (N_7987,N_7472,N_7431);
or U7988 (N_7988,N_7066,N_7485);
or U7989 (N_7989,N_7407,N_7241);
and U7990 (N_7990,N_7219,N_7383);
xor U7991 (N_7991,N_7330,N_7412);
or U7992 (N_7992,N_7250,N_7211);
xnor U7993 (N_7993,N_7114,N_7348);
and U7994 (N_7994,N_7359,N_7329);
nand U7995 (N_7995,N_7461,N_7063);
nand U7996 (N_7996,N_7117,N_7245);
and U7997 (N_7997,N_7215,N_7102);
nor U7998 (N_7998,N_7064,N_7473);
and U7999 (N_7999,N_7207,N_7063);
and U8000 (N_8000,N_7652,N_7980);
or U8001 (N_8001,N_7592,N_7645);
nand U8002 (N_8002,N_7955,N_7503);
nor U8003 (N_8003,N_7522,N_7854);
or U8004 (N_8004,N_7941,N_7504);
nand U8005 (N_8005,N_7568,N_7765);
nand U8006 (N_8006,N_7763,N_7525);
and U8007 (N_8007,N_7575,N_7659);
nand U8008 (N_8008,N_7580,N_7508);
and U8009 (N_8009,N_7721,N_7831);
or U8010 (N_8010,N_7649,N_7914);
or U8011 (N_8011,N_7550,N_7714);
xor U8012 (N_8012,N_7982,N_7595);
nand U8013 (N_8013,N_7728,N_7954);
nor U8014 (N_8014,N_7998,N_7791);
nor U8015 (N_8015,N_7705,N_7576);
or U8016 (N_8016,N_7978,N_7551);
nor U8017 (N_8017,N_7545,N_7846);
nand U8018 (N_8018,N_7739,N_7822);
nand U8019 (N_8019,N_7779,N_7662);
and U8020 (N_8020,N_7611,N_7905);
nand U8021 (N_8021,N_7530,N_7594);
and U8022 (N_8022,N_7623,N_7894);
xor U8023 (N_8023,N_7687,N_7896);
or U8024 (N_8024,N_7931,N_7947);
or U8025 (N_8025,N_7547,N_7729);
or U8026 (N_8026,N_7816,N_7851);
or U8027 (N_8027,N_7628,N_7790);
and U8028 (N_8028,N_7569,N_7967);
or U8029 (N_8029,N_7926,N_7873);
or U8030 (N_8030,N_7584,N_7839);
nor U8031 (N_8031,N_7707,N_7958);
nor U8032 (N_8032,N_7803,N_7886);
xnor U8033 (N_8033,N_7637,N_7746);
nor U8034 (N_8034,N_7853,N_7682);
or U8035 (N_8035,N_7593,N_7891);
nand U8036 (N_8036,N_7715,N_7829);
xor U8037 (N_8037,N_7857,N_7573);
xnor U8038 (N_8038,N_7909,N_7708);
nor U8039 (N_8039,N_7961,N_7513);
xnor U8040 (N_8040,N_7975,N_7579);
or U8041 (N_8041,N_7697,N_7505);
nand U8042 (N_8042,N_7651,N_7953);
xor U8043 (N_8043,N_7556,N_7937);
xor U8044 (N_8044,N_7834,N_7608);
nor U8045 (N_8045,N_7745,N_7950);
and U8046 (N_8046,N_7563,N_7850);
nand U8047 (N_8047,N_7868,N_7643);
and U8048 (N_8048,N_7985,N_7781);
xnor U8049 (N_8049,N_7747,N_7567);
and U8050 (N_8050,N_7602,N_7861);
xor U8051 (N_8051,N_7944,N_7828);
nand U8052 (N_8052,N_7972,N_7713);
xor U8053 (N_8053,N_7717,N_7883);
nor U8054 (N_8054,N_7722,N_7849);
nor U8055 (N_8055,N_7843,N_7684);
nor U8056 (N_8056,N_7830,N_7744);
xor U8057 (N_8057,N_7749,N_7660);
xor U8058 (N_8058,N_7689,N_7964);
and U8059 (N_8059,N_7981,N_7820);
nand U8060 (N_8060,N_7590,N_7604);
nand U8061 (N_8061,N_7933,N_7806);
and U8062 (N_8062,N_7596,N_7917);
nor U8063 (N_8063,N_7774,N_7994);
and U8064 (N_8064,N_7963,N_7510);
nand U8065 (N_8065,N_7733,N_7701);
or U8066 (N_8066,N_7629,N_7702);
nand U8067 (N_8067,N_7724,N_7974);
nor U8068 (N_8068,N_7795,N_7535);
nor U8069 (N_8069,N_7882,N_7805);
nand U8070 (N_8070,N_7929,N_7726);
xnor U8071 (N_8071,N_7895,N_7844);
or U8072 (N_8072,N_7549,N_7542);
xor U8073 (N_8073,N_7907,N_7712);
or U8074 (N_8074,N_7793,N_7678);
or U8075 (N_8075,N_7991,N_7809);
xor U8076 (N_8076,N_7766,N_7586);
nand U8077 (N_8077,N_7661,N_7757);
nand U8078 (N_8078,N_7585,N_7945);
or U8079 (N_8079,N_7544,N_7928);
and U8080 (N_8080,N_7581,N_7635);
nor U8081 (N_8081,N_7906,N_7564);
xnor U8082 (N_8082,N_7825,N_7633);
and U8083 (N_8083,N_7915,N_7812);
and U8084 (N_8084,N_7673,N_7741);
nand U8085 (N_8085,N_7656,N_7537);
nor U8086 (N_8086,N_7737,N_7540);
or U8087 (N_8087,N_7560,N_7858);
nand U8088 (N_8088,N_7863,N_7969);
nor U8089 (N_8089,N_7776,N_7855);
and U8090 (N_8090,N_7626,N_7815);
nor U8091 (N_8091,N_7876,N_7620);
and U8092 (N_8092,N_7865,N_7532);
or U8093 (N_8093,N_7848,N_7959);
and U8094 (N_8094,N_7898,N_7986);
xnor U8095 (N_8095,N_7818,N_7897);
nand U8096 (N_8096,N_7787,N_7845);
xnor U8097 (N_8097,N_7589,N_7615);
nand U8098 (N_8098,N_7695,N_7856);
nand U8099 (N_8099,N_7574,N_7646);
nand U8100 (N_8100,N_7672,N_7566);
or U8101 (N_8101,N_7731,N_7792);
nor U8102 (N_8102,N_7872,N_7529);
xor U8103 (N_8103,N_7804,N_7599);
nor U8104 (N_8104,N_7908,N_7640);
or U8105 (N_8105,N_7506,N_7988);
and U8106 (N_8106,N_7921,N_7810);
nand U8107 (N_8107,N_7922,N_7877);
nand U8108 (N_8108,N_7817,N_7904);
nand U8109 (N_8109,N_7704,N_7720);
nand U8110 (N_8110,N_7860,N_7807);
nand U8111 (N_8111,N_7840,N_7918);
nor U8112 (N_8112,N_7924,N_7916);
or U8113 (N_8113,N_7606,N_7962);
xnor U8114 (N_8114,N_7632,N_7966);
or U8115 (N_8115,N_7993,N_7992);
or U8116 (N_8116,N_7952,N_7501);
or U8117 (N_8117,N_7881,N_7847);
or U8118 (N_8118,N_7515,N_7605);
xnor U8119 (N_8119,N_7871,N_7583);
nand U8120 (N_8120,N_7610,N_7677);
nand U8121 (N_8121,N_7977,N_7674);
and U8122 (N_8122,N_7533,N_7698);
nor U8123 (N_8123,N_7813,N_7794);
nor U8124 (N_8124,N_7764,N_7920);
xnor U8125 (N_8125,N_7625,N_7543);
nand U8126 (N_8126,N_7838,N_7968);
nor U8127 (N_8127,N_7788,N_7837);
nor U8128 (N_8128,N_7949,N_7885);
or U8129 (N_8129,N_7923,N_7603);
and U8130 (N_8130,N_7956,N_7957);
nor U8131 (N_8131,N_7852,N_7823);
xor U8132 (N_8132,N_7658,N_7655);
or U8133 (N_8133,N_7771,N_7740);
nor U8134 (N_8134,N_7836,N_7889);
and U8135 (N_8135,N_7786,N_7627);
or U8136 (N_8136,N_7725,N_7866);
nor U8137 (N_8137,N_7801,N_7700);
and U8138 (N_8138,N_7892,N_7940);
and U8139 (N_8139,N_7631,N_7783);
and U8140 (N_8140,N_7965,N_7727);
nand U8141 (N_8141,N_7553,N_7613);
or U8142 (N_8142,N_7808,N_7557);
xor U8143 (N_8143,N_7539,N_7832);
nor U8144 (N_8144,N_7979,N_7531);
nor U8145 (N_8145,N_7752,N_7692);
nand U8146 (N_8146,N_7693,N_7711);
nand U8147 (N_8147,N_7859,N_7597);
nand U8148 (N_8148,N_7970,N_7778);
or U8149 (N_8149,N_7767,N_7591);
and U8150 (N_8150,N_7676,N_7903);
nand U8151 (N_8151,N_7696,N_7636);
nor U8152 (N_8152,N_7690,N_7887);
xor U8153 (N_8153,N_7518,N_7642);
nor U8154 (N_8154,N_7664,N_7878);
nor U8155 (N_8155,N_7507,N_7756);
nor U8156 (N_8156,N_7598,N_7694);
xnor U8157 (N_8157,N_7548,N_7538);
or U8158 (N_8158,N_7621,N_7723);
and U8159 (N_8159,N_7619,N_7572);
xor U8160 (N_8160,N_7617,N_7691);
and U8161 (N_8161,N_7912,N_7748);
nor U8162 (N_8162,N_7984,N_7934);
nor U8163 (N_8163,N_7699,N_7742);
xnor U8164 (N_8164,N_7890,N_7997);
or U8165 (N_8165,N_7624,N_7942);
xnor U8166 (N_8166,N_7743,N_7519);
or U8167 (N_8167,N_7555,N_7750);
or U8168 (N_8168,N_7870,N_7900);
and U8169 (N_8169,N_7570,N_7775);
and U8170 (N_8170,N_7768,N_7888);
xor U8171 (N_8171,N_7614,N_7800);
xnor U8172 (N_8172,N_7559,N_7841);
or U8173 (N_8173,N_7546,N_7869);
xor U8174 (N_8174,N_7925,N_7935);
or U8175 (N_8175,N_7502,N_7719);
and U8176 (N_8176,N_7996,N_7973);
nand U8177 (N_8177,N_7666,N_7639);
nor U8178 (N_8178,N_7681,N_7650);
and U8179 (N_8179,N_7670,N_7913);
nand U8180 (N_8180,N_7911,N_7893);
nand U8181 (N_8181,N_7577,N_7622);
xnor U8182 (N_8182,N_7634,N_7943);
nor U8183 (N_8183,N_7777,N_7755);
nor U8184 (N_8184,N_7554,N_7665);
nand U8185 (N_8185,N_7983,N_7987);
and U8186 (N_8186,N_7517,N_7688);
nor U8187 (N_8187,N_7738,N_7867);
and U8188 (N_8188,N_7582,N_7679);
and U8189 (N_8189,N_7938,N_7821);
nand U8190 (N_8190,N_7999,N_7683);
and U8191 (N_8191,N_7971,N_7571);
and U8192 (N_8192,N_7811,N_7862);
nor U8193 (N_8193,N_7995,N_7762);
and U8194 (N_8194,N_7798,N_7880);
nand U8195 (N_8195,N_7827,N_7565);
nand U8196 (N_8196,N_7799,N_7647);
xor U8197 (N_8197,N_7899,N_7772);
or U8198 (N_8198,N_7511,N_7716);
and U8199 (N_8199,N_7509,N_7932);
nand U8200 (N_8200,N_7703,N_7990);
xor U8201 (N_8201,N_7675,N_7946);
xnor U8202 (N_8202,N_7930,N_7706);
or U8203 (N_8203,N_7520,N_7874);
or U8204 (N_8204,N_7512,N_7562);
or U8205 (N_8205,N_7734,N_7780);
and U8206 (N_8206,N_7789,N_7819);
or U8207 (N_8207,N_7770,N_7864);
nand U8208 (N_8208,N_7751,N_7607);
nor U8209 (N_8209,N_7630,N_7951);
and U8210 (N_8210,N_7609,N_7814);
nor U8211 (N_8211,N_7797,N_7578);
and U8212 (N_8212,N_7600,N_7561);
nand U8213 (N_8213,N_7758,N_7833);
xor U8214 (N_8214,N_7835,N_7718);
nand U8215 (N_8215,N_7773,N_7796);
and U8216 (N_8216,N_7910,N_7618);
xor U8217 (N_8217,N_7976,N_7686);
and U8218 (N_8218,N_7824,N_7782);
or U8219 (N_8219,N_7759,N_7653);
nor U8220 (N_8220,N_7526,N_7552);
xnor U8221 (N_8221,N_7588,N_7784);
or U8222 (N_8222,N_7902,N_7534);
nor U8223 (N_8223,N_7736,N_7601);
and U8224 (N_8224,N_7641,N_7657);
xor U8225 (N_8225,N_7669,N_7654);
xor U8226 (N_8226,N_7558,N_7521);
nor U8227 (N_8227,N_7802,N_7667);
nand U8228 (N_8228,N_7901,N_7732);
nor U8229 (N_8229,N_7638,N_7753);
nand U8230 (N_8230,N_7710,N_7612);
nand U8231 (N_8231,N_7527,N_7927);
nor U8232 (N_8232,N_7685,N_7528);
and U8233 (N_8233,N_7644,N_7769);
nand U8234 (N_8234,N_7648,N_7541);
xnor U8235 (N_8235,N_7785,N_7939);
and U8236 (N_8236,N_7730,N_7536);
nor U8237 (N_8237,N_7826,N_7989);
or U8238 (N_8238,N_7616,N_7500);
nand U8239 (N_8239,N_7587,N_7523);
xor U8240 (N_8240,N_7875,N_7671);
or U8241 (N_8241,N_7524,N_7948);
xor U8242 (N_8242,N_7514,N_7516);
nand U8243 (N_8243,N_7754,N_7879);
and U8244 (N_8244,N_7680,N_7960);
nor U8245 (N_8245,N_7735,N_7919);
nor U8246 (N_8246,N_7761,N_7760);
nand U8247 (N_8247,N_7709,N_7936);
or U8248 (N_8248,N_7663,N_7668);
and U8249 (N_8249,N_7884,N_7842);
xor U8250 (N_8250,N_7912,N_7787);
or U8251 (N_8251,N_7886,N_7910);
and U8252 (N_8252,N_7554,N_7750);
and U8253 (N_8253,N_7821,N_7530);
nand U8254 (N_8254,N_7901,N_7678);
nand U8255 (N_8255,N_7534,N_7658);
nand U8256 (N_8256,N_7842,N_7506);
nand U8257 (N_8257,N_7767,N_7679);
nand U8258 (N_8258,N_7805,N_7843);
nor U8259 (N_8259,N_7559,N_7946);
or U8260 (N_8260,N_7784,N_7738);
and U8261 (N_8261,N_7629,N_7818);
nand U8262 (N_8262,N_7836,N_7921);
or U8263 (N_8263,N_7923,N_7540);
nand U8264 (N_8264,N_7724,N_7653);
or U8265 (N_8265,N_7607,N_7841);
xor U8266 (N_8266,N_7666,N_7806);
nand U8267 (N_8267,N_7524,N_7908);
and U8268 (N_8268,N_7963,N_7556);
nor U8269 (N_8269,N_7939,N_7578);
xnor U8270 (N_8270,N_7567,N_7931);
and U8271 (N_8271,N_7757,N_7615);
and U8272 (N_8272,N_7826,N_7864);
nand U8273 (N_8273,N_7783,N_7540);
or U8274 (N_8274,N_7543,N_7870);
and U8275 (N_8275,N_7652,N_7894);
and U8276 (N_8276,N_7636,N_7634);
or U8277 (N_8277,N_7785,N_7983);
and U8278 (N_8278,N_7528,N_7579);
xor U8279 (N_8279,N_7813,N_7760);
and U8280 (N_8280,N_7665,N_7567);
xor U8281 (N_8281,N_7827,N_7561);
nor U8282 (N_8282,N_7521,N_7767);
nand U8283 (N_8283,N_7574,N_7641);
nand U8284 (N_8284,N_7725,N_7904);
nand U8285 (N_8285,N_7758,N_7695);
nand U8286 (N_8286,N_7565,N_7806);
or U8287 (N_8287,N_7849,N_7583);
and U8288 (N_8288,N_7579,N_7620);
and U8289 (N_8289,N_7528,N_7519);
or U8290 (N_8290,N_7582,N_7746);
or U8291 (N_8291,N_7825,N_7618);
or U8292 (N_8292,N_7558,N_7852);
or U8293 (N_8293,N_7533,N_7607);
or U8294 (N_8294,N_7568,N_7861);
nand U8295 (N_8295,N_7513,N_7704);
or U8296 (N_8296,N_7747,N_7788);
and U8297 (N_8297,N_7754,N_7784);
nand U8298 (N_8298,N_7537,N_7900);
nor U8299 (N_8299,N_7708,N_7527);
nand U8300 (N_8300,N_7580,N_7659);
xnor U8301 (N_8301,N_7939,N_7940);
xor U8302 (N_8302,N_7894,N_7881);
and U8303 (N_8303,N_7535,N_7857);
or U8304 (N_8304,N_7882,N_7841);
or U8305 (N_8305,N_7901,N_7500);
or U8306 (N_8306,N_7516,N_7818);
nand U8307 (N_8307,N_7867,N_7950);
and U8308 (N_8308,N_7546,N_7793);
and U8309 (N_8309,N_7734,N_7579);
xnor U8310 (N_8310,N_7851,N_7727);
and U8311 (N_8311,N_7543,N_7980);
xnor U8312 (N_8312,N_7729,N_7571);
and U8313 (N_8313,N_7906,N_7942);
nor U8314 (N_8314,N_7855,N_7911);
nand U8315 (N_8315,N_7977,N_7732);
and U8316 (N_8316,N_7983,N_7746);
nand U8317 (N_8317,N_7569,N_7778);
and U8318 (N_8318,N_7893,N_7989);
nand U8319 (N_8319,N_7675,N_7797);
or U8320 (N_8320,N_7516,N_7692);
nor U8321 (N_8321,N_7915,N_7862);
nor U8322 (N_8322,N_7764,N_7631);
xnor U8323 (N_8323,N_7823,N_7869);
nand U8324 (N_8324,N_7634,N_7641);
nor U8325 (N_8325,N_7839,N_7850);
xnor U8326 (N_8326,N_7936,N_7746);
nor U8327 (N_8327,N_7917,N_7985);
nand U8328 (N_8328,N_7972,N_7780);
nand U8329 (N_8329,N_7568,N_7784);
xor U8330 (N_8330,N_7802,N_7795);
or U8331 (N_8331,N_7753,N_7642);
and U8332 (N_8332,N_7659,N_7615);
xor U8333 (N_8333,N_7764,N_7608);
and U8334 (N_8334,N_7659,N_7651);
and U8335 (N_8335,N_7669,N_7666);
xnor U8336 (N_8336,N_7645,N_7906);
and U8337 (N_8337,N_7548,N_7625);
nand U8338 (N_8338,N_7558,N_7561);
and U8339 (N_8339,N_7903,N_7981);
nand U8340 (N_8340,N_7789,N_7534);
nor U8341 (N_8341,N_7686,N_7746);
nand U8342 (N_8342,N_7778,N_7595);
and U8343 (N_8343,N_7681,N_7716);
nor U8344 (N_8344,N_7719,N_7504);
or U8345 (N_8345,N_7718,N_7812);
nand U8346 (N_8346,N_7717,N_7622);
or U8347 (N_8347,N_7523,N_7571);
nand U8348 (N_8348,N_7733,N_7850);
xnor U8349 (N_8349,N_7811,N_7679);
nor U8350 (N_8350,N_7512,N_7710);
and U8351 (N_8351,N_7618,N_7578);
xnor U8352 (N_8352,N_7711,N_7550);
nand U8353 (N_8353,N_7708,N_7549);
xnor U8354 (N_8354,N_7606,N_7660);
and U8355 (N_8355,N_7759,N_7633);
nor U8356 (N_8356,N_7771,N_7897);
or U8357 (N_8357,N_7863,N_7883);
nand U8358 (N_8358,N_7838,N_7594);
or U8359 (N_8359,N_7953,N_7618);
nor U8360 (N_8360,N_7952,N_7899);
nor U8361 (N_8361,N_7519,N_7816);
nor U8362 (N_8362,N_7981,N_7544);
nand U8363 (N_8363,N_7838,N_7585);
and U8364 (N_8364,N_7542,N_7513);
xnor U8365 (N_8365,N_7590,N_7654);
xnor U8366 (N_8366,N_7962,N_7802);
and U8367 (N_8367,N_7795,N_7667);
xor U8368 (N_8368,N_7669,N_7579);
xnor U8369 (N_8369,N_7843,N_7643);
nand U8370 (N_8370,N_7688,N_7607);
xnor U8371 (N_8371,N_7857,N_7983);
nand U8372 (N_8372,N_7673,N_7722);
or U8373 (N_8373,N_7807,N_7901);
nor U8374 (N_8374,N_7572,N_7902);
xnor U8375 (N_8375,N_7578,N_7679);
nor U8376 (N_8376,N_7611,N_7630);
nand U8377 (N_8377,N_7502,N_7750);
nand U8378 (N_8378,N_7875,N_7883);
xor U8379 (N_8379,N_7652,N_7517);
nor U8380 (N_8380,N_7745,N_7953);
nor U8381 (N_8381,N_7985,N_7939);
xor U8382 (N_8382,N_7912,N_7999);
or U8383 (N_8383,N_7846,N_7571);
nand U8384 (N_8384,N_7921,N_7984);
or U8385 (N_8385,N_7763,N_7858);
nor U8386 (N_8386,N_7603,N_7629);
or U8387 (N_8387,N_7846,N_7917);
xnor U8388 (N_8388,N_7545,N_7653);
or U8389 (N_8389,N_7715,N_7628);
xor U8390 (N_8390,N_7914,N_7502);
nand U8391 (N_8391,N_7828,N_7962);
and U8392 (N_8392,N_7996,N_7685);
nor U8393 (N_8393,N_7875,N_7799);
xor U8394 (N_8394,N_7543,N_7944);
or U8395 (N_8395,N_7543,N_7969);
nor U8396 (N_8396,N_7819,N_7767);
xor U8397 (N_8397,N_7536,N_7646);
or U8398 (N_8398,N_7994,N_7665);
xor U8399 (N_8399,N_7959,N_7721);
and U8400 (N_8400,N_7817,N_7638);
or U8401 (N_8401,N_7720,N_7988);
nand U8402 (N_8402,N_7578,N_7858);
xor U8403 (N_8403,N_7933,N_7808);
nand U8404 (N_8404,N_7965,N_7810);
or U8405 (N_8405,N_7867,N_7811);
nor U8406 (N_8406,N_7806,N_7739);
xor U8407 (N_8407,N_7511,N_7929);
nor U8408 (N_8408,N_7711,N_7506);
nor U8409 (N_8409,N_7776,N_7730);
xnor U8410 (N_8410,N_7505,N_7592);
nor U8411 (N_8411,N_7764,N_7712);
or U8412 (N_8412,N_7646,N_7655);
or U8413 (N_8413,N_7715,N_7980);
nand U8414 (N_8414,N_7750,N_7905);
or U8415 (N_8415,N_7811,N_7830);
nor U8416 (N_8416,N_7698,N_7973);
and U8417 (N_8417,N_7788,N_7854);
xnor U8418 (N_8418,N_7908,N_7586);
or U8419 (N_8419,N_7977,N_7833);
or U8420 (N_8420,N_7966,N_7541);
and U8421 (N_8421,N_7971,N_7649);
or U8422 (N_8422,N_7782,N_7675);
or U8423 (N_8423,N_7621,N_7514);
nor U8424 (N_8424,N_7902,N_7634);
and U8425 (N_8425,N_7865,N_7741);
nor U8426 (N_8426,N_7854,N_7727);
nor U8427 (N_8427,N_7752,N_7552);
xnor U8428 (N_8428,N_7550,N_7643);
and U8429 (N_8429,N_7821,N_7569);
or U8430 (N_8430,N_7997,N_7692);
nand U8431 (N_8431,N_7908,N_7835);
nand U8432 (N_8432,N_7936,N_7699);
or U8433 (N_8433,N_7719,N_7815);
or U8434 (N_8434,N_7791,N_7830);
xnor U8435 (N_8435,N_7521,N_7556);
nand U8436 (N_8436,N_7536,N_7970);
or U8437 (N_8437,N_7720,N_7507);
or U8438 (N_8438,N_7690,N_7638);
nor U8439 (N_8439,N_7723,N_7900);
and U8440 (N_8440,N_7889,N_7727);
or U8441 (N_8441,N_7951,N_7721);
nand U8442 (N_8442,N_7854,N_7790);
xnor U8443 (N_8443,N_7830,N_7573);
or U8444 (N_8444,N_7894,N_7931);
and U8445 (N_8445,N_7753,N_7801);
nor U8446 (N_8446,N_7731,N_7570);
nand U8447 (N_8447,N_7938,N_7829);
xnor U8448 (N_8448,N_7674,N_7818);
xor U8449 (N_8449,N_7660,N_7580);
nand U8450 (N_8450,N_7623,N_7529);
or U8451 (N_8451,N_7755,N_7649);
xor U8452 (N_8452,N_7552,N_7898);
xor U8453 (N_8453,N_7830,N_7659);
xnor U8454 (N_8454,N_7649,N_7581);
xor U8455 (N_8455,N_7832,N_7733);
xnor U8456 (N_8456,N_7685,N_7600);
and U8457 (N_8457,N_7555,N_7836);
or U8458 (N_8458,N_7729,N_7940);
and U8459 (N_8459,N_7955,N_7864);
nor U8460 (N_8460,N_7851,N_7842);
and U8461 (N_8461,N_7790,N_7791);
or U8462 (N_8462,N_7954,N_7980);
and U8463 (N_8463,N_7789,N_7640);
xnor U8464 (N_8464,N_7953,N_7529);
xnor U8465 (N_8465,N_7637,N_7668);
nand U8466 (N_8466,N_7641,N_7975);
and U8467 (N_8467,N_7649,N_7709);
or U8468 (N_8468,N_7546,N_7534);
or U8469 (N_8469,N_7819,N_7979);
nor U8470 (N_8470,N_7523,N_7835);
or U8471 (N_8471,N_7697,N_7580);
nor U8472 (N_8472,N_7561,N_7998);
and U8473 (N_8473,N_7550,N_7654);
nand U8474 (N_8474,N_7895,N_7629);
nor U8475 (N_8475,N_7938,N_7678);
and U8476 (N_8476,N_7863,N_7653);
or U8477 (N_8477,N_7740,N_7898);
or U8478 (N_8478,N_7762,N_7541);
or U8479 (N_8479,N_7566,N_7830);
xor U8480 (N_8480,N_7591,N_7784);
xor U8481 (N_8481,N_7890,N_7747);
nand U8482 (N_8482,N_7792,N_7555);
or U8483 (N_8483,N_7880,N_7870);
nand U8484 (N_8484,N_7918,N_7976);
and U8485 (N_8485,N_7787,N_7520);
nand U8486 (N_8486,N_7957,N_7980);
or U8487 (N_8487,N_7791,N_7758);
nor U8488 (N_8488,N_7872,N_7860);
nor U8489 (N_8489,N_7723,N_7852);
nand U8490 (N_8490,N_7707,N_7851);
nor U8491 (N_8491,N_7599,N_7985);
xor U8492 (N_8492,N_7542,N_7563);
nor U8493 (N_8493,N_7892,N_7655);
xnor U8494 (N_8494,N_7543,N_7616);
xnor U8495 (N_8495,N_7604,N_7682);
nor U8496 (N_8496,N_7725,N_7506);
nand U8497 (N_8497,N_7632,N_7896);
nand U8498 (N_8498,N_7519,N_7726);
nor U8499 (N_8499,N_7529,N_7934);
nand U8500 (N_8500,N_8333,N_8007);
nand U8501 (N_8501,N_8237,N_8309);
nor U8502 (N_8502,N_8389,N_8489);
and U8503 (N_8503,N_8108,N_8026);
and U8504 (N_8504,N_8071,N_8063);
xor U8505 (N_8505,N_8348,N_8069);
or U8506 (N_8506,N_8251,N_8138);
or U8507 (N_8507,N_8132,N_8086);
nor U8508 (N_8508,N_8137,N_8141);
and U8509 (N_8509,N_8264,N_8328);
or U8510 (N_8510,N_8293,N_8435);
nand U8511 (N_8511,N_8487,N_8325);
and U8512 (N_8512,N_8257,N_8017);
nand U8513 (N_8513,N_8386,N_8404);
nor U8514 (N_8514,N_8024,N_8049);
or U8515 (N_8515,N_8127,N_8203);
and U8516 (N_8516,N_8482,N_8093);
nor U8517 (N_8517,N_8199,N_8245);
xnor U8518 (N_8518,N_8406,N_8265);
nand U8519 (N_8519,N_8219,N_8168);
and U8520 (N_8520,N_8167,N_8080);
nor U8521 (N_8521,N_8010,N_8258);
nor U8522 (N_8522,N_8448,N_8058);
nor U8523 (N_8523,N_8117,N_8261);
or U8524 (N_8524,N_8327,N_8409);
nand U8525 (N_8525,N_8274,N_8408);
nand U8526 (N_8526,N_8003,N_8458);
xnor U8527 (N_8527,N_8355,N_8156);
nand U8528 (N_8528,N_8198,N_8470);
nor U8529 (N_8529,N_8280,N_8322);
nor U8530 (N_8530,N_8457,N_8414);
nor U8531 (N_8531,N_8392,N_8417);
or U8532 (N_8532,N_8142,N_8332);
nor U8533 (N_8533,N_8048,N_8191);
or U8534 (N_8534,N_8352,N_8145);
or U8535 (N_8535,N_8401,N_8144);
nor U8536 (N_8536,N_8043,N_8460);
or U8537 (N_8537,N_8186,N_8312);
nand U8538 (N_8538,N_8234,N_8350);
or U8539 (N_8539,N_8396,N_8089);
nor U8540 (N_8540,N_8372,N_8387);
xor U8541 (N_8541,N_8120,N_8078);
and U8542 (N_8542,N_8464,N_8463);
or U8543 (N_8543,N_8176,N_8231);
xnor U8544 (N_8544,N_8220,N_8323);
nor U8545 (N_8545,N_8055,N_8039);
xor U8546 (N_8546,N_8107,N_8180);
xnor U8547 (N_8547,N_8393,N_8259);
nand U8548 (N_8548,N_8455,N_8228);
nand U8549 (N_8549,N_8091,N_8019);
or U8550 (N_8550,N_8371,N_8445);
or U8551 (N_8551,N_8495,N_8469);
nand U8552 (N_8552,N_8242,N_8196);
or U8553 (N_8553,N_8002,N_8032);
nand U8554 (N_8554,N_8179,N_8152);
and U8555 (N_8555,N_8082,N_8216);
xnor U8556 (N_8556,N_8166,N_8287);
xor U8557 (N_8557,N_8429,N_8115);
nor U8558 (N_8558,N_8415,N_8494);
nor U8559 (N_8559,N_8267,N_8300);
xnor U8560 (N_8560,N_8320,N_8011);
nor U8561 (N_8561,N_8496,N_8096);
nand U8562 (N_8562,N_8499,N_8381);
or U8563 (N_8563,N_8075,N_8221);
or U8564 (N_8564,N_8131,N_8051);
nand U8565 (N_8565,N_8398,N_8321);
and U8566 (N_8566,N_8420,N_8072);
and U8567 (N_8567,N_8126,N_8253);
or U8568 (N_8568,N_8119,N_8373);
or U8569 (N_8569,N_8297,N_8143);
xnor U8570 (N_8570,N_8097,N_8447);
or U8571 (N_8571,N_8356,N_8057);
nand U8572 (N_8572,N_8379,N_8122);
or U8573 (N_8573,N_8181,N_8319);
nor U8574 (N_8574,N_8247,N_8336);
and U8575 (N_8575,N_8149,N_8326);
nand U8576 (N_8576,N_8187,N_8374);
and U8577 (N_8577,N_8238,N_8292);
nor U8578 (N_8578,N_8169,N_8233);
and U8579 (N_8579,N_8354,N_8315);
and U8580 (N_8580,N_8441,N_8471);
nor U8581 (N_8581,N_8092,N_8050);
or U8582 (N_8582,N_8212,N_8250);
nor U8583 (N_8583,N_8202,N_8347);
or U8584 (N_8584,N_8283,N_8481);
xor U8585 (N_8585,N_8474,N_8079);
and U8586 (N_8586,N_8095,N_8140);
xnor U8587 (N_8587,N_8045,N_8485);
and U8588 (N_8588,N_8164,N_8206);
and U8589 (N_8589,N_8088,N_8109);
and U8590 (N_8590,N_8044,N_8439);
nand U8591 (N_8591,N_8477,N_8436);
xor U8592 (N_8592,N_8405,N_8222);
nand U8593 (N_8593,N_8298,N_8151);
nor U8594 (N_8594,N_8139,N_8468);
or U8595 (N_8595,N_8317,N_8262);
nand U8596 (N_8596,N_8330,N_8302);
and U8597 (N_8597,N_8299,N_8183);
or U8598 (N_8598,N_8130,N_8382);
xor U8599 (N_8599,N_8204,N_8214);
and U8600 (N_8600,N_8225,N_8337);
nand U8601 (N_8601,N_8025,N_8367);
and U8602 (N_8602,N_8345,N_8036);
nor U8603 (N_8603,N_8479,N_8205);
xnor U8604 (N_8604,N_8476,N_8286);
xnor U8605 (N_8605,N_8028,N_8217);
or U8606 (N_8606,N_8358,N_8483);
nand U8607 (N_8607,N_8165,N_8197);
or U8608 (N_8608,N_8146,N_8466);
or U8609 (N_8609,N_8106,N_8054);
nand U8610 (N_8610,N_8065,N_8031);
nand U8611 (N_8611,N_8004,N_8094);
nand U8612 (N_8612,N_8419,N_8136);
nor U8613 (N_8613,N_8153,N_8430);
nor U8614 (N_8614,N_8207,N_8246);
or U8615 (N_8615,N_8314,N_8121);
nand U8616 (N_8616,N_8304,N_8178);
and U8617 (N_8617,N_8005,N_8370);
and U8618 (N_8618,N_8035,N_8313);
xnor U8619 (N_8619,N_8467,N_8163);
nand U8620 (N_8620,N_8488,N_8363);
nor U8621 (N_8621,N_8318,N_8232);
xor U8622 (N_8622,N_8177,N_8229);
nand U8623 (N_8623,N_8009,N_8444);
nor U8624 (N_8624,N_8074,N_8289);
or U8625 (N_8625,N_8224,N_8239);
nor U8626 (N_8626,N_8201,N_8353);
nor U8627 (N_8627,N_8223,N_8162);
nand U8628 (N_8628,N_8281,N_8349);
xnor U8629 (N_8629,N_8475,N_8266);
xnor U8630 (N_8630,N_8013,N_8189);
nand U8631 (N_8631,N_8400,N_8147);
and U8632 (N_8632,N_8084,N_8016);
or U8633 (N_8633,N_8380,N_8486);
nand U8634 (N_8634,N_8346,N_8331);
nand U8635 (N_8635,N_8062,N_8184);
or U8636 (N_8636,N_8306,N_8324);
or U8637 (N_8637,N_8443,N_8413);
nor U8638 (N_8638,N_8307,N_8465);
nor U8639 (N_8639,N_8034,N_8378);
xnor U8640 (N_8640,N_8193,N_8135);
or U8641 (N_8641,N_8422,N_8244);
or U8642 (N_8642,N_8215,N_8394);
and U8643 (N_8643,N_8484,N_8454);
nor U8644 (N_8644,N_8182,N_8085);
xor U8645 (N_8645,N_8158,N_8113);
nand U8646 (N_8646,N_8296,N_8450);
and U8647 (N_8647,N_8282,N_8269);
xnor U8648 (N_8648,N_8123,N_8171);
or U8649 (N_8649,N_8277,N_8357);
or U8650 (N_8650,N_8273,N_8027);
and U8651 (N_8651,N_8070,N_8060);
xor U8652 (N_8652,N_8437,N_8159);
nand U8653 (N_8653,N_8284,N_8428);
nor U8654 (N_8654,N_8341,N_8343);
and U8655 (N_8655,N_8365,N_8490);
xor U8656 (N_8656,N_8335,N_8059);
nand U8657 (N_8657,N_8295,N_8377);
nor U8658 (N_8658,N_8360,N_8001);
or U8659 (N_8659,N_8061,N_8000);
nor U8660 (N_8660,N_8211,N_8278);
xnor U8661 (N_8661,N_8390,N_8150);
nor U8662 (N_8662,N_8105,N_8200);
xor U8663 (N_8663,N_8342,N_8192);
nand U8664 (N_8664,N_8218,N_8068);
and U8665 (N_8665,N_8427,N_8449);
or U8666 (N_8666,N_8263,N_8399);
or U8667 (N_8667,N_8442,N_8255);
nand U8668 (N_8668,N_8424,N_8423);
nor U8669 (N_8669,N_8038,N_8103);
nand U8670 (N_8670,N_8112,N_8473);
and U8671 (N_8671,N_8497,N_8491);
nor U8672 (N_8672,N_8279,N_8056);
nand U8673 (N_8673,N_8275,N_8340);
nor U8674 (N_8674,N_8172,N_8361);
nand U8675 (N_8675,N_8190,N_8362);
xor U8676 (N_8676,N_8310,N_8480);
nand U8677 (N_8677,N_8285,N_8101);
nor U8678 (N_8678,N_8432,N_8174);
and U8679 (N_8679,N_8128,N_8431);
nor U8680 (N_8680,N_8294,N_8154);
or U8681 (N_8681,N_8376,N_8226);
and U8682 (N_8682,N_8388,N_8129);
xor U8683 (N_8683,N_8241,N_8368);
or U8684 (N_8684,N_8334,N_8029);
nor U8685 (N_8685,N_8230,N_8451);
nand U8686 (N_8686,N_8160,N_8478);
xnor U8687 (N_8687,N_8369,N_8030);
nor U8688 (N_8688,N_8456,N_8366);
or U8689 (N_8689,N_8271,N_8194);
or U8690 (N_8690,N_8402,N_8046);
xor U8691 (N_8691,N_8008,N_8073);
nand U8692 (N_8692,N_8033,N_8066);
and U8693 (N_8693,N_8014,N_8087);
and U8694 (N_8694,N_8134,N_8155);
or U8695 (N_8695,N_8157,N_8339);
nor U8696 (N_8696,N_8037,N_8351);
and U8697 (N_8697,N_8208,N_8411);
and U8698 (N_8698,N_8012,N_8124);
nor U8699 (N_8699,N_8083,N_8498);
nand U8700 (N_8700,N_8359,N_8006);
nor U8701 (N_8701,N_8116,N_8344);
nor U8702 (N_8702,N_8170,N_8493);
or U8703 (N_8703,N_8173,N_8375);
nor U8704 (N_8704,N_8453,N_8022);
nand U8705 (N_8705,N_8260,N_8301);
nor U8706 (N_8706,N_8053,N_8042);
and U8707 (N_8707,N_8303,N_8110);
xor U8708 (N_8708,N_8185,N_8047);
nand U8709 (N_8709,N_8385,N_8213);
nand U8710 (N_8710,N_8111,N_8148);
xnor U8711 (N_8711,N_8288,N_8438);
nand U8712 (N_8712,N_8099,N_8240);
nand U8713 (N_8713,N_8041,N_8254);
or U8714 (N_8714,N_8418,N_8195);
or U8715 (N_8715,N_8472,N_8291);
nor U8716 (N_8716,N_8383,N_8077);
nor U8717 (N_8717,N_8446,N_8227);
or U8718 (N_8718,N_8272,N_8403);
nor U8719 (N_8719,N_8076,N_8209);
or U8720 (N_8720,N_8236,N_8114);
or U8721 (N_8721,N_8018,N_8270);
and U8722 (N_8722,N_8276,N_8248);
and U8723 (N_8723,N_8015,N_8452);
and U8724 (N_8724,N_8243,N_8052);
and U8725 (N_8725,N_8098,N_8407);
nor U8726 (N_8726,N_8102,N_8249);
xor U8727 (N_8727,N_8311,N_8021);
xor U8728 (N_8728,N_8397,N_8412);
xor U8729 (N_8729,N_8235,N_8256);
nand U8730 (N_8730,N_8384,N_8133);
nand U8731 (N_8731,N_8459,N_8064);
nand U8732 (N_8732,N_8305,N_8023);
nor U8733 (N_8733,N_8100,N_8416);
xnor U8734 (N_8734,N_8391,N_8440);
nor U8735 (N_8735,N_8308,N_8434);
nand U8736 (N_8736,N_8364,N_8395);
or U8737 (N_8737,N_8268,N_8188);
nor U8738 (N_8738,N_8492,N_8125);
or U8739 (N_8739,N_8425,N_8252);
and U8740 (N_8740,N_8433,N_8461);
nand U8741 (N_8741,N_8338,N_8290);
and U8742 (N_8742,N_8040,N_8329);
and U8743 (N_8743,N_8104,N_8410);
nand U8744 (N_8744,N_8316,N_8421);
xnor U8745 (N_8745,N_8090,N_8175);
or U8746 (N_8746,N_8081,N_8067);
nand U8747 (N_8747,N_8210,N_8426);
and U8748 (N_8748,N_8462,N_8161);
and U8749 (N_8749,N_8020,N_8118);
or U8750 (N_8750,N_8042,N_8051);
or U8751 (N_8751,N_8408,N_8471);
nand U8752 (N_8752,N_8200,N_8059);
nor U8753 (N_8753,N_8013,N_8442);
and U8754 (N_8754,N_8356,N_8436);
or U8755 (N_8755,N_8415,N_8287);
and U8756 (N_8756,N_8271,N_8073);
nor U8757 (N_8757,N_8129,N_8409);
or U8758 (N_8758,N_8309,N_8111);
nor U8759 (N_8759,N_8444,N_8012);
nand U8760 (N_8760,N_8498,N_8064);
nand U8761 (N_8761,N_8308,N_8423);
and U8762 (N_8762,N_8340,N_8341);
nor U8763 (N_8763,N_8469,N_8347);
and U8764 (N_8764,N_8396,N_8190);
or U8765 (N_8765,N_8010,N_8422);
and U8766 (N_8766,N_8441,N_8186);
xor U8767 (N_8767,N_8394,N_8013);
and U8768 (N_8768,N_8457,N_8415);
nor U8769 (N_8769,N_8386,N_8419);
or U8770 (N_8770,N_8165,N_8185);
xnor U8771 (N_8771,N_8250,N_8023);
nor U8772 (N_8772,N_8151,N_8450);
and U8773 (N_8773,N_8498,N_8028);
xor U8774 (N_8774,N_8196,N_8402);
nor U8775 (N_8775,N_8173,N_8492);
nand U8776 (N_8776,N_8422,N_8182);
nand U8777 (N_8777,N_8319,N_8178);
and U8778 (N_8778,N_8338,N_8366);
or U8779 (N_8779,N_8288,N_8077);
nand U8780 (N_8780,N_8064,N_8240);
nor U8781 (N_8781,N_8192,N_8104);
nor U8782 (N_8782,N_8428,N_8252);
nand U8783 (N_8783,N_8497,N_8037);
and U8784 (N_8784,N_8416,N_8113);
and U8785 (N_8785,N_8214,N_8423);
xor U8786 (N_8786,N_8326,N_8333);
or U8787 (N_8787,N_8098,N_8498);
and U8788 (N_8788,N_8458,N_8253);
nor U8789 (N_8789,N_8297,N_8420);
and U8790 (N_8790,N_8002,N_8115);
and U8791 (N_8791,N_8470,N_8042);
nand U8792 (N_8792,N_8280,N_8233);
xor U8793 (N_8793,N_8085,N_8328);
and U8794 (N_8794,N_8009,N_8295);
xnor U8795 (N_8795,N_8107,N_8165);
or U8796 (N_8796,N_8078,N_8353);
and U8797 (N_8797,N_8313,N_8030);
nand U8798 (N_8798,N_8123,N_8490);
and U8799 (N_8799,N_8426,N_8279);
and U8800 (N_8800,N_8032,N_8470);
nand U8801 (N_8801,N_8250,N_8186);
or U8802 (N_8802,N_8282,N_8072);
nand U8803 (N_8803,N_8348,N_8455);
or U8804 (N_8804,N_8297,N_8278);
or U8805 (N_8805,N_8461,N_8490);
and U8806 (N_8806,N_8085,N_8022);
xnor U8807 (N_8807,N_8424,N_8356);
and U8808 (N_8808,N_8411,N_8441);
nand U8809 (N_8809,N_8482,N_8049);
and U8810 (N_8810,N_8317,N_8345);
and U8811 (N_8811,N_8404,N_8479);
xor U8812 (N_8812,N_8187,N_8343);
nand U8813 (N_8813,N_8015,N_8042);
nor U8814 (N_8814,N_8467,N_8452);
or U8815 (N_8815,N_8108,N_8443);
and U8816 (N_8816,N_8270,N_8327);
and U8817 (N_8817,N_8408,N_8141);
xor U8818 (N_8818,N_8263,N_8114);
and U8819 (N_8819,N_8269,N_8200);
and U8820 (N_8820,N_8177,N_8258);
or U8821 (N_8821,N_8264,N_8063);
or U8822 (N_8822,N_8125,N_8257);
or U8823 (N_8823,N_8226,N_8448);
nand U8824 (N_8824,N_8140,N_8021);
nand U8825 (N_8825,N_8191,N_8376);
xnor U8826 (N_8826,N_8236,N_8433);
nor U8827 (N_8827,N_8253,N_8273);
nand U8828 (N_8828,N_8274,N_8226);
and U8829 (N_8829,N_8370,N_8464);
and U8830 (N_8830,N_8239,N_8091);
nor U8831 (N_8831,N_8310,N_8234);
nor U8832 (N_8832,N_8145,N_8351);
or U8833 (N_8833,N_8459,N_8312);
or U8834 (N_8834,N_8109,N_8226);
nand U8835 (N_8835,N_8272,N_8095);
nand U8836 (N_8836,N_8043,N_8434);
nand U8837 (N_8837,N_8281,N_8290);
nand U8838 (N_8838,N_8448,N_8192);
xor U8839 (N_8839,N_8424,N_8447);
xnor U8840 (N_8840,N_8028,N_8146);
xor U8841 (N_8841,N_8307,N_8374);
or U8842 (N_8842,N_8176,N_8105);
xor U8843 (N_8843,N_8193,N_8236);
nor U8844 (N_8844,N_8070,N_8175);
nand U8845 (N_8845,N_8157,N_8435);
xnor U8846 (N_8846,N_8228,N_8494);
or U8847 (N_8847,N_8365,N_8346);
and U8848 (N_8848,N_8377,N_8169);
xor U8849 (N_8849,N_8131,N_8091);
and U8850 (N_8850,N_8330,N_8249);
nor U8851 (N_8851,N_8141,N_8339);
or U8852 (N_8852,N_8373,N_8274);
or U8853 (N_8853,N_8341,N_8148);
xnor U8854 (N_8854,N_8175,N_8235);
and U8855 (N_8855,N_8140,N_8386);
nand U8856 (N_8856,N_8403,N_8273);
or U8857 (N_8857,N_8384,N_8171);
xnor U8858 (N_8858,N_8104,N_8446);
nor U8859 (N_8859,N_8447,N_8116);
nand U8860 (N_8860,N_8462,N_8046);
and U8861 (N_8861,N_8485,N_8438);
nor U8862 (N_8862,N_8048,N_8098);
nor U8863 (N_8863,N_8355,N_8384);
and U8864 (N_8864,N_8365,N_8489);
or U8865 (N_8865,N_8241,N_8153);
nand U8866 (N_8866,N_8036,N_8183);
and U8867 (N_8867,N_8384,N_8104);
nand U8868 (N_8868,N_8357,N_8313);
nor U8869 (N_8869,N_8194,N_8302);
nand U8870 (N_8870,N_8180,N_8260);
xor U8871 (N_8871,N_8340,N_8013);
nor U8872 (N_8872,N_8421,N_8147);
nor U8873 (N_8873,N_8189,N_8266);
nor U8874 (N_8874,N_8289,N_8375);
and U8875 (N_8875,N_8061,N_8155);
nand U8876 (N_8876,N_8369,N_8103);
or U8877 (N_8877,N_8389,N_8197);
or U8878 (N_8878,N_8226,N_8370);
nor U8879 (N_8879,N_8416,N_8382);
and U8880 (N_8880,N_8484,N_8036);
or U8881 (N_8881,N_8468,N_8207);
or U8882 (N_8882,N_8291,N_8459);
nor U8883 (N_8883,N_8247,N_8285);
and U8884 (N_8884,N_8059,N_8229);
and U8885 (N_8885,N_8015,N_8462);
nand U8886 (N_8886,N_8435,N_8498);
or U8887 (N_8887,N_8288,N_8406);
or U8888 (N_8888,N_8163,N_8402);
nor U8889 (N_8889,N_8445,N_8158);
or U8890 (N_8890,N_8092,N_8278);
nor U8891 (N_8891,N_8413,N_8476);
nand U8892 (N_8892,N_8255,N_8151);
nor U8893 (N_8893,N_8338,N_8425);
nand U8894 (N_8894,N_8105,N_8480);
nand U8895 (N_8895,N_8126,N_8325);
xor U8896 (N_8896,N_8089,N_8466);
nor U8897 (N_8897,N_8455,N_8023);
or U8898 (N_8898,N_8288,N_8072);
xnor U8899 (N_8899,N_8011,N_8102);
and U8900 (N_8900,N_8089,N_8347);
or U8901 (N_8901,N_8412,N_8143);
nor U8902 (N_8902,N_8125,N_8185);
nand U8903 (N_8903,N_8366,N_8303);
and U8904 (N_8904,N_8495,N_8022);
or U8905 (N_8905,N_8115,N_8006);
and U8906 (N_8906,N_8372,N_8342);
and U8907 (N_8907,N_8174,N_8305);
nor U8908 (N_8908,N_8374,N_8316);
or U8909 (N_8909,N_8004,N_8170);
nor U8910 (N_8910,N_8491,N_8073);
nor U8911 (N_8911,N_8006,N_8377);
nor U8912 (N_8912,N_8311,N_8364);
xnor U8913 (N_8913,N_8460,N_8324);
nand U8914 (N_8914,N_8158,N_8068);
nand U8915 (N_8915,N_8197,N_8003);
or U8916 (N_8916,N_8382,N_8192);
nor U8917 (N_8917,N_8227,N_8027);
xor U8918 (N_8918,N_8203,N_8134);
nor U8919 (N_8919,N_8477,N_8372);
xnor U8920 (N_8920,N_8429,N_8004);
nand U8921 (N_8921,N_8050,N_8408);
or U8922 (N_8922,N_8375,N_8390);
nor U8923 (N_8923,N_8142,N_8026);
xnor U8924 (N_8924,N_8348,N_8240);
nor U8925 (N_8925,N_8003,N_8020);
xnor U8926 (N_8926,N_8200,N_8292);
xnor U8927 (N_8927,N_8219,N_8314);
and U8928 (N_8928,N_8477,N_8345);
nand U8929 (N_8929,N_8442,N_8292);
or U8930 (N_8930,N_8259,N_8312);
nand U8931 (N_8931,N_8198,N_8284);
or U8932 (N_8932,N_8485,N_8245);
nand U8933 (N_8933,N_8197,N_8083);
xor U8934 (N_8934,N_8123,N_8175);
xor U8935 (N_8935,N_8283,N_8369);
xnor U8936 (N_8936,N_8255,N_8209);
nor U8937 (N_8937,N_8324,N_8284);
or U8938 (N_8938,N_8290,N_8341);
and U8939 (N_8939,N_8266,N_8115);
and U8940 (N_8940,N_8019,N_8191);
and U8941 (N_8941,N_8128,N_8178);
nor U8942 (N_8942,N_8208,N_8306);
xnor U8943 (N_8943,N_8121,N_8333);
and U8944 (N_8944,N_8226,N_8335);
nor U8945 (N_8945,N_8477,N_8263);
and U8946 (N_8946,N_8470,N_8365);
nand U8947 (N_8947,N_8354,N_8196);
nand U8948 (N_8948,N_8490,N_8372);
or U8949 (N_8949,N_8247,N_8363);
or U8950 (N_8950,N_8297,N_8194);
or U8951 (N_8951,N_8163,N_8490);
xor U8952 (N_8952,N_8000,N_8187);
nand U8953 (N_8953,N_8281,N_8135);
or U8954 (N_8954,N_8137,N_8014);
nand U8955 (N_8955,N_8184,N_8448);
nor U8956 (N_8956,N_8205,N_8290);
xnor U8957 (N_8957,N_8006,N_8138);
or U8958 (N_8958,N_8235,N_8088);
and U8959 (N_8959,N_8238,N_8073);
nand U8960 (N_8960,N_8470,N_8446);
and U8961 (N_8961,N_8071,N_8481);
nand U8962 (N_8962,N_8329,N_8378);
and U8963 (N_8963,N_8165,N_8084);
nor U8964 (N_8964,N_8497,N_8134);
nand U8965 (N_8965,N_8104,N_8368);
or U8966 (N_8966,N_8373,N_8055);
nor U8967 (N_8967,N_8481,N_8234);
or U8968 (N_8968,N_8062,N_8494);
or U8969 (N_8969,N_8359,N_8287);
nor U8970 (N_8970,N_8262,N_8011);
nor U8971 (N_8971,N_8074,N_8237);
nand U8972 (N_8972,N_8100,N_8095);
or U8973 (N_8973,N_8118,N_8052);
nor U8974 (N_8974,N_8070,N_8000);
nor U8975 (N_8975,N_8059,N_8091);
nor U8976 (N_8976,N_8269,N_8160);
xnor U8977 (N_8977,N_8335,N_8198);
and U8978 (N_8978,N_8140,N_8056);
nand U8979 (N_8979,N_8372,N_8001);
nand U8980 (N_8980,N_8445,N_8295);
nand U8981 (N_8981,N_8228,N_8090);
or U8982 (N_8982,N_8022,N_8033);
or U8983 (N_8983,N_8286,N_8446);
xnor U8984 (N_8984,N_8064,N_8472);
or U8985 (N_8985,N_8002,N_8183);
or U8986 (N_8986,N_8087,N_8423);
nor U8987 (N_8987,N_8411,N_8271);
xor U8988 (N_8988,N_8409,N_8335);
and U8989 (N_8989,N_8430,N_8186);
xor U8990 (N_8990,N_8296,N_8236);
and U8991 (N_8991,N_8123,N_8477);
nor U8992 (N_8992,N_8202,N_8488);
or U8993 (N_8993,N_8127,N_8376);
nand U8994 (N_8994,N_8023,N_8169);
or U8995 (N_8995,N_8275,N_8320);
nor U8996 (N_8996,N_8420,N_8328);
or U8997 (N_8997,N_8122,N_8161);
and U8998 (N_8998,N_8099,N_8370);
xnor U8999 (N_8999,N_8263,N_8435);
nor U9000 (N_9000,N_8832,N_8761);
nand U9001 (N_9001,N_8542,N_8641);
nand U9002 (N_9002,N_8666,N_8640);
xor U9003 (N_9003,N_8680,N_8509);
or U9004 (N_9004,N_8563,N_8629);
and U9005 (N_9005,N_8622,N_8784);
nand U9006 (N_9006,N_8725,N_8528);
and U9007 (N_9007,N_8543,N_8778);
xor U9008 (N_9008,N_8994,N_8651);
nand U9009 (N_9009,N_8535,N_8963);
nor U9010 (N_9010,N_8697,N_8532);
nor U9011 (N_9011,N_8781,N_8598);
nand U9012 (N_9012,N_8817,N_8688);
nor U9013 (N_9013,N_8689,N_8610);
nand U9014 (N_9014,N_8770,N_8816);
nor U9015 (N_9015,N_8732,N_8615);
xnor U9016 (N_9016,N_8857,N_8804);
and U9017 (N_9017,N_8913,N_8556);
nor U9018 (N_9018,N_8845,N_8964);
nor U9019 (N_9019,N_8707,N_8966);
and U9020 (N_9020,N_8704,N_8934);
or U9021 (N_9021,N_8821,N_8534);
nand U9022 (N_9022,N_8541,N_8976);
nand U9023 (N_9023,N_8861,N_8691);
xnor U9024 (N_9024,N_8518,N_8973);
nand U9025 (N_9025,N_8918,N_8800);
and U9026 (N_9026,N_8671,N_8917);
and U9027 (N_9027,N_8802,N_8843);
and U9028 (N_9028,N_8649,N_8925);
or U9029 (N_9029,N_8951,N_8654);
xnor U9030 (N_9030,N_8812,N_8893);
nor U9031 (N_9031,N_8739,N_8795);
and U9032 (N_9032,N_8677,N_8808);
nor U9033 (N_9033,N_8959,N_8969);
nor U9034 (N_9034,N_8814,N_8529);
and U9035 (N_9035,N_8879,N_8679);
nor U9036 (N_9036,N_8895,N_8836);
or U9037 (N_9037,N_8743,N_8864);
xor U9038 (N_9038,N_8884,N_8702);
nor U9039 (N_9039,N_8866,N_8599);
or U9040 (N_9040,N_8575,N_8674);
and U9041 (N_9041,N_8765,N_8608);
or U9042 (N_9042,N_8506,N_8862);
xor U9043 (N_9043,N_8742,N_8692);
and U9044 (N_9044,N_8844,N_8948);
nor U9045 (N_9045,N_8955,N_8990);
or U9046 (N_9046,N_8714,N_8724);
xnor U9047 (N_9047,N_8617,N_8570);
and U9048 (N_9048,N_8786,N_8605);
or U9049 (N_9049,N_8909,N_8665);
and U9050 (N_9050,N_8762,N_8758);
and U9051 (N_9051,N_8578,N_8823);
or U9052 (N_9052,N_8829,N_8635);
or U9053 (N_9053,N_8612,N_8504);
xor U9054 (N_9054,N_8639,N_8926);
nand U9055 (N_9055,N_8752,N_8712);
nor U9056 (N_9056,N_8953,N_8811);
nand U9057 (N_9057,N_8924,N_8946);
or U9058 (N_9058,N_8858,N_8636);
or U9059 (N_9059,N_8863,N_8956);
nand U9060 (N_9060,N_8503,N_8820);
nor U9061 (N_9061,N_8719,N_8915);
and U9062 (N_9062,N_8731,N_8664);
and U9063 (N_9063,N_8967,N_8849);
xnor U9064 (N_9064,N_8941,N_8944);
or U9065 (N_9065,N_8632,N_8744);
xor U9066 (N_9066,N_8908,N_8746);
and U9067 (N_9067,N_8899,N_8898);
or U9068 (N_9068,N_8872,N_8876);
xor U9069 (N_9069,N_8868,N_8565);
and U9070 (N_9070,N_8995,N_8873);
and U9071 (N_9071,N_8633,N_8831);
nand U9072 (N_9072,N_8979,N_8985);
nand U9073 (N_9073,N_8984,N_8538);
nor U9074 (N_9074,N_8930,N_8776);
or U9075 (N_9075,N_8569,N_8830);
and U9076 (N_9076,N_8757,N_8896);
nor U9077 (N_9077,N_8813,N_8774);
or U9078 (N_9078,N_8668,N_8625);
or U9079 (N_9079,N_8584,N_8737);
and U9080 (N_9080,N_8711,N_8760);
and U9081 (N_9081,N_8833,N_8968);
nor U9082 (N_9082,N_8897,N_8870);
and U9083 (N_9083,N_8787,N_8526);
xnor U9084 (N_9084,N_8591,N_8658);
or U9085 (N_9085,N_8996,N_8588);
nand U9086 (N_9086,N_8928,N_8581);
and U9087 (N_9087,N_8949,N_8838);
nor U9088 (N_9088,N_8708,N_8601);
or U9089 (N_9089,N_8763,N_8684);
nand U9090 (N_9090,N_8989,N_8929);
nand U9091 (N_9091,N_8693,N_8960);
nand U9092 (N_9092,N_8906,N_8524);
or U9093 (N_9093,N_8593,N_8840);
nand U9094 (N_9094,N_8950,N_8508);
or U9095 (N_9095,N_8777,N_8611);
nand U9096 (N_9096,N_8669,N_8613);
or U9097 (N_9097,N_8931,N_8860);
xnor U9098 (N_9098,N_8754,N_8888);
nor U9099 (N_9099,N_8631,N_8887);
or U9100 (N_9100,N_8740,N_8537);
nor U9101 (N_9101,N_8846,N_8722);
and U9102 (N_9102,N_8997,N_8877);
xnor U9103 (N_9103,N_8954,N_8907);
xor U9104 (N_9104,N_8616,N_8785);
and U9105 (N_9105,N_8571,N_8585);
xnor U9106 (N_9106,N_8828,N_8583);
xor U9107 (N_9107,N_8520,N_8919);
nor U9108 (N_9108,N_8695,N_8505);
or U9109 (N_9109,N_8618,N_8975);
xor U9110 (N_9110,N_8661,N_8573);
nand U9111 (N_9111,N_8839,N_8983);
or U9112 (N_9112,N_8775,N_8513);
and U9113 (N_9113,N_8728,N_8676);
and U9114 (N_9114,N_8962,N_8594);
nand U9115 (N_9115,N_8590,N_8619);
or U9116 (N_9116,N_8738,N_8815);
or U9117 (N_9117,N_8834,N_8747);
and U9118 (N_9118,N_8652,N_8683);
and U9119 (N_9119,N_8942,N_8721);
and U9120 (N_9120,N_8567,N_8965);
or U9121 (N_9121,N_8952,N_8792);
xor U9122 (N_9122,N_8938,N_8947);
or U9123 (N_9123,N_8933,N_8624);
or U9124 (N_9124,N_8937,N_8726);
or U9125 (N_9125,N_8670,N_8793);
xnor U9126 (N_9126,N_8595,N_8700);
xnor U9127 (N_9127,N_8771,N_8678);
or U9128 (N_9128,N_8998,N_8699);
nand U9129 (N_9129,N_8606,N_8703);
nand U9130 (N_9130,N_8856,N_8980);
nand U9131 (N_9131,N_8993,N_8987);
and U9132 (N_9132,N_8852,N_8882);
nand U9133 (N_9133,N_8579,N_8554);
or U9134 (N_9134,N_8523,N_8748);
and U9135 (N_9135,N_8592,N_8791);
xnor U9136 (N_9136,N_8662,N_8727);
and U9137 (N_9137,N_8730,N_8540);
xnor U9138 (N_9138,N_8560,N_8603);
xor U9139 (N_9139,N_8656,N_8660);
nor U9140 (N_9140,N_8902,N_8709);
nand U9141 (N_9141,N_8847,N_8970);
nor U9142 (N_9142,N_8568,N_8885);
and U9143 (N_9143,N_8886,N_8685);
nor U9144 (N_9144,N_8600,N_8911);
or U9145 (N_9145,N_8690,N_8779);
nor U9146 (N_9146,N_8500,N_8647);
nand U9147 (N_9147,N_8871,N_8536);
xor U9148 (N_9148,N_8723,N_8552);
nand U9149 (N_9149,N_8741,N_8945);
or U9150 (N_9150,N_8672,N_8927);
nand U9151 (N_9151,N_8566,N_8530);
or U9152 (N_9152,N_8853,N_8533);
xnor U9153 (N_9153,N_8932,N_8644);
and U9154 (N_9154,N_8630,N_8551);
and U9155 (N_9155,N_8623,N_8715);
or U9156 (N_9156,N_8614,N_8735);
xor U9157 (N_9157,N_8974,N_8891);
and U9158 (N_9158,N_8904,N_8865);
or U9159 (N_9159,N_8798,N_8681);
nor U9160 (N_9160,N_8710,N_8650);
nand U9161 (N_9161,N_8790,N_8646);
nand U9162 (N_9162,N_8991,N_8957);
nor U9163 (N_9163,N_8653,N_8559);
xnor U9164 (N_9164,N_8733,N_8905);
and U9165 (N_9165,N_8971,N_8626);
and U9166 (N_9166,N_8522,N_8782);
nor U9167 (N_9167,N_8992,N_8604);
and U9168 (N_9168,N_8648,N_8696);
nand U9169 (N_9169,N_8841,N_8659);
or U9170 (N_9170,N_8548,N_8705);
nand U9171 (N_9171,N_8637,N_8634);
xor U9172 (N_9172,N_8914,N_8824);
or U9173 (N_9173,N_8806,N_8686);
and U9174 (N_9174,N_8645,N_8597);
and U9175 (N_9175,N_8557,N_8912);
nand U9176 (N_9176,N_8892,N_8881);
or U9177 (N_9177,N_8713,N_8794);
or U9178 (N_9178,N_8920,N_8745);
or U9179 (N_9179,N_8922,N_8521);
and U9180 (N_9180,N_8848,N_8586);
xnor U9181 (N_9181,N_8826,N_8687);
or U9182 (N_9182,N_8517,N_8511);
nand U9183 (N_9183,N_8675,N_8799);
or U9184 (N_9184,N_8514,N_8803);
nand U9185 (N_9185,N_8550,N_8910);
and U9186 (N_9186,N_8716,N_8545);
nand U9187 (N_9187,N_8589,N_8516);
nand U9188 (N_9188,N_8796,N_8572);
nand U9189 (N_9189,N_8935,N_8507);
nor U9190 (N_9190,N_8621,N_8602);
xnor U9191 (N_9191,N_8961,N_8519);
nand U9192 (N_9192,N_8576,N_8851);
nand U9193 (N_9193,N_8878,N_8574);
and U9194 (N_9194,N_8673,N_8978);
nor U9195 (N_9195,N_8580,N_8883);
or U9196 (N_9196,N_8810,N_8547);
nor U9197 (N_9197,N_8515,N_8807);
and U9198 (N_9198,N_8982,N_8694);
or U9199 (N_9199,N_8531,N_8682);
nand U9200 (N_9200,N_8720,N_8903);
xor U9201 (N_9201,N_8880,N_8874);
and U9202 (N_9202,N_8766,N_8736);
and U9203 (N_9203,N_8502,N_8958);
xor U9204 (N_9204,N_8875,N_8577);
or U9205 (N_9205,N_8759,N_8642);
nand U9206 (N_9206,N_8729,N_8825);
nor U9207 (N_9207,N_8890,N_8609);
nor U9208 (N_9208,N_8663,N_8544);
and U9209 (N_9209,N_8837,N_8628);
nand U9210 (N_9210,N_8867,N_8859);
or U9211 (N_9211,N_8797,N_8587);
nand U9212 (N_9212,N_8850,N_8582);
or U9213 (N_9213,N_8527,N_8769);
nand U9214 (N_9214,N_8555,N_8939);
xnor U9215 (N_9215,N_8717,N_8698);
xor U9216 (N_9216,N_8749,N_8667);
and U9217 (N_9217,N_8943,N_8510);
and U9218 (N_9218,N_8553,N_8539);
nor U9219 (N_9219,N_8734,N_8921);
and U9220 (N_9220,N_8805,N_8854);
nor U9221 (N_9221,N_8988,N_8855);
or U9222 (N_9222,N_8607,N_8706);
nor U9223 (N_9223,N_8638,N_8755);
xnor U9224 (N_9224,N_8501,N_8549);
and U9225 (N_9225,N_8780,N_8756);
nor U9226 (N_9226,N_8981,N_8783);
or U9227 (N_9227,N_8900,N_8869);
and U9228 (N_9228,N_8561,N_8809);
xor U9229 (N_9229,N_8767,N_8558);
and U9230 (N_9230,N_8972,N_8819);
xor U9231 (N_9231,N_8564,N_8620);
nand U9232 (N_9232,N_8788,N_8822);
and U9233 (N_9233,N_8842,N_8701);
nand U9234 (N_9234,N_8999,N_8750);
nand U9235 (N_9235,N_8773,N_8718);
nand U9236 (N_9236,N_8657,N_8764);
nor U9237 (N_9237,N_8894,N_8923);
nor U9238 (N_9238,N_8512,N_8827);
nand U9239 (N_9239,N_8801,N_8772);
and U9240 (N_9240,N_8525,N_8562);
and U9241 (N_9241,N_8751,N_8768);
or U9242 (N_9242,N_8916,N_8835);
nand U9243 (N_9243,N_8901,N_8655);
nand U9244 (N_9244,N_8643,N_8936);
xor U9245 (N_9245,N_8546,N_8977);
xnor U9246 (N_9246,N_8889,N_8596);
nand U9247 (N_9247,N_8940,N_8818);
nor U9248 (N_9248,N_8753,N_8789);
nor U9249 (N_9249,N_8986,N_8627);
xnor U9250 (N_9250,N_8532,N_8720);
nand U9251 (N_9251,N_8691,N_8805);
nor U9252 (N_9252,N_8840,N_8929);
and U9253 (N_9253,N_8796,N_8560);
or U9254 (N_9254,N_8723,N_8850);
and U9255 (N_9255,N_8576,N_8790);
and U9256 (N_9256,N_8749,N_8598);
or U9257 (N_9257,N_8778,N_8723);
nor U9258 (N_9258,N_8808,N_8554);
nor U9259 (N_9259,N_8984,N_8632);
nand U9260 (N_9260,N_8805,N_8567);
and U9261 (N_9261,N_8668,N_8921);
or U9262 (N_9262,N_8864,N_8531);
nor U9263 (N_9263,N_8901,N_8894);
or U9264 (N_9264,N_8682,N_8833);
nor U9265 (N_9265,N_8597,N_8803);
nor U9266 (N_9266,N_8908,N_8829);
nor U9267 (N_9267,N_8683,N_8743);
or U9268 (N_9268,N_8899,N_8571);
xnor U9269 (N_9269,N_8611,N_8990);
nor U9270 (N_9270,N_8750,N_8645);
nor U9271 (N_9271,N_8504,N_8626);
and U9272 (N_9272,N_8517,N_8850);
nor U9273 (N_9273,N_8505,N_8845);
or U9274 (N_9274,N_8751,N_8744);
nor U9275 (N_9275,N_8561,N_8669);
xnor U9276 (N_9276,N_8642,N_8788);
xnor U9277 (N_9277,N_8745,N_8589);
nand U9278 (N_9278,N_8574,N_8675);
or U9279 (N_9279,N_8573,N_8865);
or U9280 (N_9280,N_8522,N_8648);
xor U9281 (N_9281,N_8644,N_8603);
or U9282 (N_9282,N_8844,N_8639);
or U9283 (N_9283,N_8936,N_8621);
xor U9284 (N_9284,N_8556,N_8595);
xnor U9285 (N_9285,N_8752,N_8905);
or U9286 (N_9286,N_8730,N_8514);
nor U9287 (N_9287,N_8511,N_8593);
xor U9288 (N_9288,N_8699,N_8562);
or U9289 (N_9289,N_8516,N_8680);
and U9290 (N_9290,N_8570,N_8819);
nand U9291 (N_9291,N_8940,N_8547);
or U9292 (N_9292,N_8880,N_8642);
nor U9293 (N_9293,N_8654,N_8878);
nand U9294 (N_9294,N_8691,N_8972);
or U9295 (N_9295,N_8634,N_8582);
and U9296 (N_9296,N_8790,N_8922);
xnor U9297 (N_9297,N_8782,N_8817);
nor U9298 (N_9298,N_8539,N_8823);
nor U9299 (N_9299,N_8605,N_8642);
and U9300 (N_9300,N_8552,N_8534);
nand U9301 (N_9301,N_8529,N_8873);
nor U9302 (N_9302,N_8768,N_8987);
nand U9303 (N_9303,N_8573,N_8851);
nor U9304 (N_9304,N_8814,N_8795);
or U9305 (N_9305,N_8616,N_8743);
nor U9306 (N_9306,N_8606,N_8936);
nand U9307 (N_9307,N_8687,N_8720);
and U9308 (N_9308,N_8984,N_8863);
xnor U9309 (N_9309,N_8769,N_8788);
nor U9310 (N_9310,N_8914,N_8871);
or U9311 (N_9311,N_8719,N_8720);
nand U9312 (N_9312,N_8927,N_8951);
nand U9313 (N_9313,N_8840,N_8951);
xor U9314 (N_9314,N_8670,N_8972);
nand U9315 (N_9315,N_8621,N_8915);
xor U9316 (N_9316,N_8777,N_8770);
and U9317 (N_9317,N_8739,N_8566);
or U9318 (N_9318,N_8869,N_8942);
nand U9319 (N_9319,N_8954,N_8782);
nor U9320 (N_9320,N_8903,N_8622);
nor U9321 (N_9321,N_8510,N_8969);
and U9322 (N_9322,N_8996,N_8952);
nor U9323 (N_9323,N_8541,N_8792);
or U9324 (N_9324,N_8694,N_8899);
xnor U9325 (N_9325,N_8914,N_8664);
nand U9326 (N_9326,N_8751,N_8828);
and U9327 (N_9327,N_8594,N_8969);
nor U9328 (N_9328,N_8953,N_8955);
or U9329 (N_9329,N_8803,N_8958);
nand U9330 (N_9330,N_8556,N_8555);
nand U9331 (N_9331,N_8954,N_8983);
or U9332 (N_9332,N_8578,N_8613);
nor U9333 (N_9333,N_8983,N_8973);
or U9334 (N_9334,N_8989,N_8811);
or U9335 (N_9335,N_8747,N_8599);
and U9336 (N_9336,N_8741,N_8507);
nand U9337 (N_9337,N_8565,N_8511);
or U9338 (N_9338,N_8714,N_8641);
and U9339 (N_9339,N_8538,N_8565);
or U9340 (N_9340,N_8564,N_8926);
xor U9341 (N_9341,N_8666,N_8664);
or U9342 (N_9342,N_8839,N_8832);
nand U9343 (N_9343,N_8944,N_8575);
or U9344 (N_9344,N_8768,N_8934);
and U9345 (N_9345,N_8929,N_8693);
nand U9346 (N_9346,N_8553,N_8649);
and U9347 (N_9347,N_8877,N_8762);
nand U9348 (N_9348,N_8732,N_8789);
nor U9349 (N_9349,N_8981,N_8674);
nand U9350 (N_9350,N_8662,N_8915);
and U9351 (N_9351,N_8505,N_8917);
nor U9352 (N_9352,N_8952,N_8778);
and U9353 (N_9353,N_8966,N_8562);
and U9354 (N_9354,N_8655,N_8563);
nor U9355 (N_9355,N_8873,N_8607);
nor U9356 (N_9356,N_8848,N_8669);
nor U9357 (N_9357,N_8973,N_8766);
xnor U9358 (N_9358,N_8504,N_8605);
or U9359 (N_9359,N_8917,N_8902);
and U9360 (N_9360,N_8575,N_8731);
nor U9361 (N_9361,N_8928,N_8965);
nand U9362 (N_9362,N_8813,N_8710);
or U9363 (N_9363,N_8620,N_8815);
or U9364 (N_9364,N_8974,N_8645);
xor U9365 (N_9365,N_8822,N_8687);
nand U9366 (N_9366,N_8976,N_8628);
or U9367 (N_9367,N_8659,N_8942);
nor U9368 (N_9368,N_8968,N_8971);
and U9369 (N_9369,N_8705,N_8915);
xor U9370 (N_9370,N_8532,N_8841);
nor U9371 (N_9371,N_8949,N_8686);
and U9372 (N_9372,N_8617,N_8862);
xnor U9373 (N_9373,N_8975,N_8513);
nor U9374 (N_9374,N_8923,N_8847);
nand U9375 (N_9375,N_8526,N_8903);
and U9376 (N_9376,N_8985,N_8514);
nand U9377 (N_9377,N_8942,N_8770);
or U9378 (N_9378,N_8625,N_8820);
and U9379 (N_9379,N_8562,N_8572);
or U9380 (N_9380,N_8604,N_8969);
and U9381 (N_9381,N_8810,N_8928);
and U9382 (N_9382,N_8650,N_8662);
xor U9383 (N_9383,N_8909,N_8734);
or U9384 (N_9384,N_8900,N_8785);
nand U9385 (N_9385,N_8980,N_8951);
nand U9386 (N_9386,N_8503,N_8656);
nand U9387 (N_9387,N_8641,N_8509);
or U9388 (N_9388,N_8967,N_8741);
xor U9389 (N_9389,N_8746,N_8782);
xor U9390 (N_9390,N_8911,N_8579);
nand U9391 (N_9391,N_8874,N_8659);
nand U9392 (N_9392,N_8814,N_8883);
nor U9393 (N_9393,N_8991,N_8716);
or U9394 (N_9394,N_8726,N_8769);
nand U9395 (N_9395,N_8918,N_8583);
nand U9396 (N_9396,N_8836,N_8947);
nor U9397 (N_9397,N_8994,N_8805);
xnor U9398 (N_9398,N_8960,N_8833);
and U9399 (N_9399,N_8544,N_8874);
or U9400 (N_9400,N_8505,N_8718);
xor U9401 (N_9401,N_8783,N_8677);
xor U9402 (N_9402,N_8978,N_8588);
xnor U9403 (N_9403,N_8578,N_8709);
nand U9404 (N_9404,N_8896,N_8754);
and U9405 (N_9405,N_8526,N_8893);
and U9406 (N_9406,N_8517,N_8737);
and U9407 (N_9407,N_8555,N_8706);
nand U9408 (N_9408,N_8787,N_8542);
or U9409 (N_9409,N_8948,N_8747);
nand U9410 (N_9410,N_8587,N_8873);
xnor U9411 (N_9411,N_8553,N_8758);
and U9412 (N_9412,N_8829,N_8944);
nor U9413 (N_9413,N_8631,N_8634);
nor U9414 (N_9414,N_8667,N_8842);
or U9415 (N_9415,N_8541,N_8889);
nand U9416 (N_9416,N_8884,N_8666);
nor U9417 (N_9417,N_8566,N_8824);
nand U9418 (N_9418,N_8619,N_8645);
nand U9419 (N_9419,N_8969,N_8847);
xor U9420 (N_9420,N_8911,N_8659);
or U9421 (N_9421,N_8989,N_8603);
nor U9422 (N_9422,N_8892,N_8845);
nand U9423 (N_9423,N_8902,N_8939);
nand U9424 (N_9424,N_8938,N_8762);
nand U9425 (N_9425,N_8560,N_8639);
nor U9426 (N_9426,N_8599,N_8722);
nor U9427 (N_9427,N_8974,N_8789);
xnor U9428 (N_9428,N_8991,N_8681);
and U9429 (N_9429,N_8921,N_8653);
nand U9430 (N_9430,N_8907,N_8942);
or U9431 (N_9431,N_8526,N_8505);
or U9432 (N_9432,N_8931,N_8588);
xnor U9433 (N_9433,N_8736,N_8553);
or U9434 (N_9434,N_8532,N_8770);
nor U9435 (N_9435,N_8902,N_8611);
nor U9436 (N_9436,N_8646,N_8664);
or U9437 (N_9437,N_8627,N_8832);
xnor U9438 (N_9438,N_8592,N_8558);
nor U9439 (N_9439,N_8795,N_8619);
or U9440 (N_9440,N_8611,N_8568);
and U9441 (N_9441,N_8953,N_8796);
and U9442 (N_9442,N_8561,N_8794);
or U9443 (N_9443,N_8840,N_8558);
and U9444 (N_9444,N_8516,N_8958);
nand U9445 (N_9445,N_8683,N_8581);
or U9446 (N_9446,N_8551,N_8939);
nor U9447 (N_9447,N_8735,N_8998);
or U9448 (N_9448,N_8547,N_8742);
or U9449 (N_9449,N_8556,N_8793);
or U9450 (N_9450,N_8508,N_8631);
and U9451 (N_9451,N_8969,N_8511);
and U9452 (N_9452,N_8916,N_8584);
nor U9453 (N_9453,N_8923,N_8751);
or U9454 (N_9454,N_8878,N_8669);
nand U9455 (N_9455,N_8620,N_8759);
or U9456 (N_9456,N_8778,N_8775);
nor U9457 (N_9457,N_8502,N_8541);
nor U9458 (N_9458,N_8539,N_8669);
nand U9459 (N_9459,N_8747,N_8950);
and U9460 (N_9460,N_8641,N_8546);
or U9461 (N_9461,N_8811,N_8855);
xnor U9462 (N_9462,N_8642,N_8649);
nor U9463 (N_9463,N_8905,N_8793);
and U9464 (N_9464,N_8605,N_8846);
nor U9465 (N_9465,N_8930,N_8631);
and U9466 (N_9466,N_8984,N_8524);
or U9467 (N_9467,N_8551,N_8642);
nor U9468 (N_9468,N_8667,N_8563);
or U9469 (N_9469,N_8780,N_8798);
or U9470 (N_9470,N_8565,N_8826);
and U9471 (N_9471,N_8796,N_8903);
nand U9472 (N_9472,N_8892,N_8978);
and U9473 (N_9473,N_8580,N_8735);
and U9474 (N_9474,N_8808,N_8600);
xor U9475 (N_9475,N_8521,N_8512);
nor U9476 (N_9476,N_8839,N_8918);
or U9477 (N_9477,N_8938,N_8716);
nand U9478 (N_9478,N_8563,N_8650);
xnor U9479 (N_9479,N_8775,N_8913);
nor U9480 (N_9480,N_8695,N_8547);
nand U9481 (N_9481,N_8925,N_8965);
nand U9482 (N_9482,N_8662,N_8810);
and U9483 (N_9483,N_8650,N_8978);
nand U9484 (N_9484,N_8981,N_8602);
and U9485 (N_9485,N_8916,N_8569);
nor U9486 (N_9486,N_8915,N_8846);
and U9487 (N_9487,N_8627,N_8618);
or U9488 (N_9488,N_8833,N_8591);
nand U9489 (N_9489,N_8752,N_8515);
xor U9490 (N_9490,N_8953,N_8614);
and U9491 (N_9491,N_8662,N_8781);
or U9492 (N_9492,N_8839,N_8536);
and U9493 (N_9493,N_8698,N_8750);
and U9494 (N_9494,N_8522,N_8951);
and U9495 (N_9495,N_8900,N_8964);
nand U9496 (N_9496,N_8855,N_8605);
or U9497 (N_9497,N_8725,N_8662);
nor U9498 (N_9498,N_8822,N_8985);
xor U9499 (N_9499,N_8601,N_8740);
nand U9500 (N_9500,N_9175,N_9022);
or U9501 (N_9501,N_9165,N_9043);
or U9502 (N_9502,N_9248,N_9087);
nor U9503 (N_9503,N_9005,N_9388);
or U9504 (N_9504,N_9468,N_9184);
nor U9505 (N_9505,N_9091,N_9077);
nor U9506 (N_9506,N_9339,N_9482);
and U9507 (N_9507,N_9372,N_9306);
xor U9508 (N_9508,N_9334,N_9282);
xor U9509 (N_9509,N_9057,N_9030);
nand U9510 (N_9510,N_9144,N_9418);
or U9511 (N_9511,N_9347,N_9283);
nor U9512 (N_9512,N_9391,N_9220);
nor U9513 (N_9513,N_9108,N_9237);
nor U9514 (N_9514,N_9470,N_9092);
nand U9515 (N_9515,N_9225,N_9122);
nand U9516 (N_9516,N_9099,N_9369);
or U9517 (N_9517,N_9274,N_9477);
or U9518 (N_9518,N_9221,N_9459);
or U9519 (N_9519,N_9136,N_9176);
and U9520 (N_9520,N_9309,N_9150);
nor U9521 (N_9521,N_9152,N_9238);
xor U9522 (N_9522,N_9276,N_9169);
xnor U9523 (N_9523,N_9444,N_9246);
nand U9524 (N_9524,N_9054,N_9449);
and U9525 (N_9525,N_9455,N_9322);
or U9526 (N_9526,N_9013,N_9191);
or U9527 (N_9527,N_9198,N_9362);
nor U9528 (N_9528,N_9179,N_9126);
xor U9529 (N_9529,N_9416,N_9249);
or U9530 (N_9530,N_9121,N_9399);
or U9531 (N_9531,N_9042,N_9446);
xor U9532 (N_9532,N_9348,N_9166);
or U9533 (N_9533,N_9371,N_9051);
nand U9534 (N_9534,N_9330,N_9208);
xor U9535 (N_9535,N_9116,N_9385);
nand U9536 (N_9536,N_9392,N_9113);
or U9537 (N_9537,N_9496,N_9298);
nor U9538 (N_9538,N_9110,N_9268);
xnor U9539 (N_9539,N_9431,N_9442);
xnor U9540 (N_9540,N_9223,N_9017);
nor U9541 (N_9541,N_9243,N_9066);
or U9542 (N_9542,N_9183,N_9286);
nor U9543 (N_9543,N_9417,N_9211);
nand U9544 (N_9544,N_9281,N_9458);
xnor U9545 (N_9545,N_9404,N_9199);
xor U9546 (N_9546,N_9015,N_9341);
nor U9547 (N_9547,N_9472,N_9316);
and U9548 (N_9548,N_9457,N_9397);
or U9549 (N_9549,N_9354,N_9186);
nand U9550 (N_9550,N_9337,N_9378);
and U9551 (N_9551,N_9124,N_9086);
nor U9552 (N_9552,N_9395,N_9190);
xnor U9553 (N_9553,N_9296,N_9173);
and U9554 (N_9554,N_9139,N_9252);
or U9555 (N_9555,N_9021,N_9090);
xor U9556 (N_9556,N_9490,N_9102);
or U9557 (N_9557,N_9025,N_9480);
and U9558 (N_9558,N_9055,N_9426);
nor U9559 (N_9559,N_9300,N_9471);
nand U9560 (N_9560,N_9026,N_9429);
and U9561 (N_9561,N_9188,N_9445);
nand U9562 (N_9562,N_9224,N_9142);
or U9563 (N_9563,N_9212,N_9251);
nand U9564 (N_9564,N_9332,N_9326);
and U9565 (N_9565,N_9273,N_9235);
xor U9566 (N_9566,N_9178,N_9396);
nand U9567 (N_9567,N_9301,N_9400);
nor U9568 (N_9568,N_9203,N_9314);
nand U9569 (N_9569,N_9185,N_9156);
nand U9570 (N_9570,N_9196,N_9058);
nand U9571 (N_9571,N_9089,N_9230);
and U9572 (N_9572,N_9375,N_9264);
and U9573 (N_9573,N_9101,N_9127);
nor U9574 (N_9574,N_9344,N_9453);
and U9575 (N_9575,N_9202,N_9390);
xor U9576 (N_9576,N_9061,N_9419);
nand U9577 (N_9577,N_9037,N_9168);
nor U9578 (N_9578,N_9327,N_9159);
or U9579 (N_9579,N_9174,N_9063);
nor U9580 (N_9580,N_9259,N_9240);
nand U9581 (N_9581,N_9236,N_9125);
nor U9582 (N_9582,N_9140,N_9161);
or U9583 (N_9583,N_9187,N_9189);
and U9584 (N_9584,N_9201,N_9265);
nor U9585 (N_9585,N_9483,N_9335);
nand U9586 (N_9586,N_9070,N_9381);
or U9587 (N_9587,N_9052,N_9473);
nand U9588 (N_9588,N_9180,N_9411);
xnor U9589 (N_9589,N_9412,N_9351);
xor U9590 (N_9590,N_9352,N_9096);
and U9591 (N_9591,N_9085,N_9250);
and U9592 (N_9592,N_9115,N_9487);
and U9593 (N_9593,N_9493,N_9149);
and U9594 (N_9594,N_9106,N_9428);
nand U9595 (N_9595,N_9181,N_9171);
or U9596 (N_9596,N_9491,N_9423);
nand U9597 (N_9597,N_9374,N_9147);
or U9598 (N_9598,N_9083,N_9297);
xor U9599 (N_9599,N_9361,N_9498);
nand U9600 (N_9600,N_9364,N_9422);
nand U9601 (N_9601,N_9394,N_9387);
and U9602 (N_9602,N_9258,N_9462);
or U9603 (N_9603,N_9353,N_9117);
nand U9604 (N_9604,N_9340,N_9228);
or U9605 (N_9605,N_9155,N_9001);
nand U9606 (N_9606,N_9207,N_9217);
nand U9607 (N_9607,N_9050,N_9131);
xor U9608 (N_9608,N_9024,N_9130);
xnor U9609 (N_9609,N_9094,N_9226);
or U9610 (N_9610,N_9318,N_9244);
xnor U9611 (N_9611,N_9204,N_9329);
and U9612 (N_9612,N_9038,N_9256);
xor U9613 (N_9613,N_9290,N_9216);
nand U9614 (N_9614,N_9359,N_9135);
nand U9615 (N_9615,N_9414,N_9098);
nand U9616 (N_9616,N_9153,N_9078);
nand U9617 (N_9617,N_9193,N_9409);
nor U9618 (N_9618,N_9103,N_9325);
xnor U9619 (N_9619,N_9401,N_9014);
or U9620 (N_9620,N_9007,N_9137);
and U9621 (N_9621,N_9345,N_9475);
or U9622 (N_9622,N_9338,N_9012);
xnor U9623 (N_9623,N_9272,N_9255);
and U9624 (N_9624,N_9313,N_9295);
xnor U9625 (N_9625,N_9486,N_9355);
or U9626 (N_9626,N_9435,N_9280);
nor U9627 (N_9627,N_9049,N_9287);
nor U9628 (N_9628,N_9160,N_9143);
or U9629 (N_9629,N_9182,N_9023);
nand U9630 (N_9630,N_9020,N_9109);
or U9631 (N_9631,N_9386,N_9242);
nor U9632 (N_9632,N_9154,N_9499);
and U9633 (N_9633,N_9425,N_9321);
and U9634 (N_9634,N_9018,N_9408);
nand U9635 (N_9635,N_9358,N_9467);
nand U9636 (N_9636,N_9003,N_9073);
nor U9637 (N_9637,N_9076,N_9254);
xor U9638 (N_9638,N_9114,N_9485);
nand U9639 (N_9639,N_9346,N_9492);
or U9640 (N_9640,N_9209,N_9461);
nand U9641 (N_9641,N_9393,N_9036);
or U9642 (N_9642,N_9261,N_9481);
nand U9643 (N_9643,N_9439,N_9464);
or U9644 (N_9644,N_9488,N_9262);
or U9645 (N_9645,N_9271,N_9430);
and U9646 (N_9646,N_9291,N_9138);
nor U9647 (N_9647,N_9440,N_9257);
xnor U9648 (N_9648,N_9082,N_9420);
xor U9649 (N_9649,N_9097,N_9031);
xnor U9650 (N_9650,N_9357,N_9305);
nor U9651 (N_9651,N_9000,N_9370);
nand U9652 (N_9652,N_9029,N_9456);
xor U9653 (N_9653,N_9320,N_9466);
nand U9654 (N_9654,N_9075,N_9004);
xor U9655 (N_9655,N_9474,N_9343);
nand U9656 (N_9656,N_9373,N_9402);
nand U9657 (N_9657,N_9035,N_9383);
xnor U9658 (N_9658,N_9071,N_9148);
nand U9659 (N_9659,N_9095,N_9247);
and U9660 (N_9660,N_9319,N_9484);
or U9661 (N_9661,N_9403,N_9336);
nor U9662 (N_9662,N_9494,N_9288);
and U9663 (N_9663,N_9436,N_9134);
or U9664 (N_9664,N_9376,N_9123);
and U9665 (N_9665,N_9200,N_9307);
nor U9666 (N_9666,N_9294,N_9410);
nand U9667 (N_9667,N_9333,N_9206);
xor U9668 (N_9668,N_9415,N_9479);
or U9669 (N_9669,N_9463,N_9064);
or U9670 (N_9670,N_9232,N_9311);
nor U9671 (N_9671,N_9145,N_9424);
and U9672 (N_9672,N_9047,N_9151);
or U9673 (N_9673,N_9368,N_9405);
and U9674 (N_9674,N_9460,N_9310);
nor U9675 (N_9675,N_9040,N_9019);
xor U9676 (N_9676,N_9105,N_9380);
xnor U9677 (N_9677,N_9195,N_9497);
and U9678 (N_9678,N_9065,N_9079);
or U9679 (N_9679,N_9111,N_9413);
or U9680 (N_9680,N_9495,N_9053);
nor U9681 (N_9681,N_9120,N_9011);
nand U9682 (N_9682,N_9008,N_9215);
or U9683 (N_9683,N_9447,N_9219);
nor U9684 (N_9684,N_9443,N_9239);
xnor U9685 (N_9685,N_9027,N_9093);
xnor U9686 (N_9686,N_9041,N_9284);
nand U9687 (N_9687,N_9100,N_9366);
xor U9688 (N_9688,N_9299,N_9363);
nand U9689 (N_9689,N_9253,N_9056);
and U9690 (N_9690,N_9270,N_9129);
or U9691 (N_9691,N_9278,N_9277);
nand U9692 (N_9692,N_9118,N_9241);
and U9693 (N_9693,N_9192,N_9448);
xnor U9694 (N_9694,N_9197,N_9450);
nor U9695 (N_9695,N_9062,N_9222);
nand U9696 (N_9696,N_9275,N_9324);
nor U9697 (N_9697,N_9231,N_9107);
xor U9698 (N_9698,N_9128,N_9379);
nor U9699 (N_9699,N_9177,N_9048);
xnor U9700 (N_9700,N_9146,N_9302);
or U9701 (N_9701,N_9432,N_9263);
nand U9702 (N_9702,N_9437,N_9072);
and U9703 (N_9703,N_9006,N_9465);
and U9704 (N_9704,N_9328,N_9194);
nand U9705 (N_9705,N_9469,N_9342);
or U9706 (N_9706,N_9304,N_9260);
or U9707 (N_9707,N_9356,N_9266);
and U9708 (N_9708,N_9205,N_9112);
xnor U9709 (N_9709,N_9088,N_9451);
xor U9710 (N_9710,N_9028,N_9245);
xor U9711 (N_9711,N_9269,N_9210);
nor U9712 (N_9712,N_9104,N_9009);
and U9713 (N_9713,N_9454,N_9367);
nand U9714 (N_9714,N_9389,N_9421);
nand U9715 (N_9715,N_9045,N_9331);
nand U9716 (N_9716,N_9308,N_9084);
and U9717 (N_9717,N_9032,N_9312);
and U9718 (N_9718,N_9489,N_9227);
xor U9719 (N_9719,N_9452,N_9349);
or U9720 (N_9720,N_9292,N_9060);
nand U9721 (N_9721,N_9163,N_9214);
or U9722 (N_9722,N_9289,N_9044);
xor U9723 (N_9723,N_9059,N_9267);
xor U9724 (N_9724,N_9046,N_9382);
xnor U9725 (N_9725,N_9317,N_9384);
or U9726 (N_9726,N_9433,N_9074);
or U9727 (N_9727,N_9164,N_9010);
and U9728 (N_9728,N_9303,N_9167);
xnor U9729 (N_9729,N_9119,N_9081);
and U9730 (N_9730,N_9157,N_9377);
nor U9731 (N_9731,N_9441,N_9350);
and U9732 (N_9732,N_9039,N_9323);
nand U9733 (N_9733,N_9438,N_9233);
or U9734 (N_9734,N_9285,N_9434);
nor U9735 (N_9735,N_9002,N_9080);
nand U9736 (N_9736,N_9293,N_9068);
or U9737 (N_9737,N_9478,N_9218);
nand U9738 (N_9738,N_9406,N_9172);
nor U9739 (N_9739,N_9069,N_9315);
nor U9740 (N_9740,N_9213,N_9360);
or U9741 (N_9741,N_9407,N_9170);
nor U9742 (N_9742,N_9067,N_9398);
xor U9743 (N_9743,N_9162,N_9033);
nand U9744 (N_9744,N_9234,N_9133);
nand U9745 (N_9745,N_9158,N_9427);
nand U9746 (N_9746,N_9132,N_9279);
xor U9747 (N_9747,N_9016,N_9229);
nor U9748 (N_9748,N_9365,N_9141);
xor U9749 (N_9749,N_9476,N_9034);
xnor U9750 (N_9750,N_9047,N_9248);
or U9751 (N_9751,N_9350,N_9392);
nand U9752 (N_9752,N_9491,N_9010);
or U9753 (N_9753,N_9457,N_9429);
or U9754 (N_9754,N_9182,N_9436);
and U9755 (N_9755,N_9188,N_9396);
xnor U9756 (N_9756,N_9492,N_9476);
and U9757 (N_9757,N_9394,N_9045);
nor U9758 (N_9758,N_9073,N_9484);
or U9759 (N_9759,N_9436,N_9132);
nand U9760 (N_9760,N_9111,N_9452);
or U9761 (N_9761,N_9431,N_9008);
nor U9762 (N_9762,N_9334,N_9308);
nor U9763 (N_9763,N_9393,N_9273);
and U9764 (N_9764,N_9210,N_9044);
or U9765 (N_9765,N_9034,N_9200);
or U9766 (N_9766,N_9464,N_9245);
nand U9767 (N_9767,N_9399,N_9462);
xnor U9768 (N_9768,N_9489,N_9042);
nor U9769 (N_9769,N_9475,N_9070);
and U9770 (N_9770,N_9355,N_9129);
nand U9771 (N_9771,N_9377,N_9474);
or U9772 (N_9772,N_9058,N_9038);
and U9773 (N_9773,N_9052,N_9159);
or U9774 (N_9774,N_9284,N_9113);
and U9775 (N_9775,N_9014,N_9146);
nor U9776 (N_9776,N_9410,N_9017);
nand U9777 (N_9777,N_9098,N_9042);
and U9778 (N_9778,N_9168,N_9008);
nand U9779 (N_9779,N_9303,N_9009);
nor U9780 (N_9780,N_9069,N_9049);
or U9781 (N_9781,N_9182,N_9357);
and U9782 (N_9782,N_9425,N_9052);
or U9783 (N_9783,N_9379,N_9178);
or U9784 (N_9784,N_9180,N_9392);
and U9785 (N_9785,N_9274,N_9231);
and U9786 (N_9786,N_9424,N_9461);
xor U9787 (N_9787,N_9202,N_9376);
and U9788 (N_9788,N_9444,N_9114);
or U9789 (N_9789,N_9278,N_9231);
xnor U9790 (N_9790,N_9358,N_9395);
or U9791 (N_9791,N_9128,N_9374);
nor U9792 (N_9792,N_9004,N_9431);
xor U9793 (N_9793,N_9014,N_9192);
xor U9794 (N_9794,N_9254,N_9255);
xnor U9795 (N_9795,N_9116,N_9062);
or U9796 (N_9796,N_9296,N_9136);
nor U9797 (N_9797,N_9402,N_9054);
and U9798 (N_9798,N_9424,N_9221);
nand U9799 (N_9799,N_9354,N_9457);
and U9800 (N_9800,N_9402,N_9189);
or U9801 (N_9801,N_9071,N_9005);
xor U9802 (N_9802,N_9219,N_9044);
xor U9803 (N_9803,N_9340,N_9057);
and U9804 (N_9804,N_9019,N_9293);
and U9805 (N_9805,N_9286,N_9101);
and U9806 (N_9806,N_9222,N_9211);
and U9807 (N_9807,N_9149,N_9026);
xor U9808 (N_9808,N_9393,N_9220);
nand U9809 (N_9809,N_9382,N_9465);
xnor U9810 (N_9810,N_9309,N_9182);
xnor U9811 (N_9811,N_9014,N_9304);
and U9812 (N_9812,N_9308,N_9371);
or U9813 (N_9813,N_9350,N_9050);
or U9814 (N_9814,N_9421,N_9104);
nor U9815 (N_9815,N_9194,N_9250);
nand U9816 (N_9816,N_9131,N_9434);
or U9817 (N_9817,N_9159,N_9173);
nor U9818 (N_9818,N_9425,N_9352);
nand U9819 (N_9819,N_9459,N_9498);
nor U9820 (N_9820,N_9295,N_9075);
xor U9821 (N_9821,N_9436,N_9454);
nand U9822 (N_9822,N_9383,N_9241);
xor U9823 (N_9823,N_9307,N_9171);
and U9824 (N_9824,N_9087,N_9195);
and U9825 (N_9825,N_9138,N_9497);
xor U9826 (N_9826,N_9181,N_9107);
nor U9827 (N_9827,N_9203,N_9395);
and U9828 (N_9828,N_9224,N_9058);
nor U9829 (N_9829,N_9273,N_9244);
or U9830 (N_9830,N_9376,N_9413);
xnor U9831 (N_9831,N_9455,N_9126);
and U9832 (N_9832,N_9041,N_9134);
and U9833 (N_9833,N_9432,N_9053);
and U9834 (N_9834,N_9288,N_9396);
xnor U9835 (N_9835,N_9064,N_9184);
and U9836 (N_9836,N_9030,N_9229);
or U9837 (N_9837,N_9437,N_9049);
or U9838 (N_9838,N_9297,N_9183);
or U9839 (N_9839,N_9098,N_9321);
xnor U9840 (N_9840,N_9127,N_9280);
nor U9841 (N_9841,N_9332,N_9394);
nand U9842 (N_9842,N_9229,N_9061);
xor U9843 (N_9843,N_9494,N_9358);
and U9844 (N_9844,N_9171,N_9436);
nor U9845 (N_9845,N_9299,N_9001);
nand U9846 (N_9846,N_9284,N_9353);
and U9847 (N_9847,N_9117,N_9194);
nand U9848 (N_9848,N_9478,N_9144);
xor U9849 (N_9849,N_9026,N_9220);
and U9850 (N_9850,N_9269,N_9425);
and U9851 (N_9851,N_9314,N_9445);
nor U9852 (N_9852,N_9397,N_9065);
and U9853 (N_9853,N_9318,N_9278);
and U9854 (N_9854,N_9473,N_9344);
or U9855 (N_9855,N_9489,N_9251);
nor U9856 (N_9856,N_9209,N_9274);
xor U9857 (N_9857,N_9406,N_9448);
nand U9858 (N_9858,N_9166,N_9286);
or U9859 (N_9859,N_9237,N_9432);
nor U9860 (N_9860,N_9008,N_9268);
and U9861 (N_9861,N_9432,N_9013);
and U9862 (N_9862,N_9306,N_9126);
nand U9863 (N_9863,N_9241,N_9363);
or U9864 (N_9864,N_9181,N_9263);
and U9865 (N_9865,N_9119,N_9352);
nor U9866 (N_9866,N_9019,N_9088);
xor U9867 (N_9867,N_9192,N_9443);
xnor U9868 (N_9868,N_9146,N_9293);
nor U9869 (N_9869,N_9205,N_9065);
nor U9870 (N_9870,N_9428,N_9190);
and U9871 (N_9871,N_9274,N_9398);
nand U9872 (N_9872,N_9425,N_9327);
nand U9873 (N_9873,N_9235,N_9301);
and U9874 (N_9874,N_9256,N_9107);
nor U9875 (N_9875,N_9163,N_9140);
and U9876 (N_9876,N_9426,N_9157);
nor U9877 (N_9877,N_9400,N_9470);
or U9878 (N_9878,N_9018,N_9442);
nand U9879 (N_9879,N_9086,N_9282);
and U9880 (N_9880,N_9163,N_9454);
xor U9881 (N_9881,N_9173,N_9433);
or U9882 (N_9882,N_9088,N_9035);
nand U9883 (N_9883,N_9243,N_9146);
and U9884 (N_9884,N_9151,N_9303);
or U9885 (N_9885,N_9376,N_9495);
xor U9886 (N_9886,N_9005,N_9301);
or U9887 (N_9887,N_9358,N_9191);
nor U9888 (N_9888,N_9370,N_9335);
nor U9889 (N_9889,N_9054,N_9164);
and U9890 (N_9890,N_9469,N_9000);
nor U9891 (N_9891,N_9219,N_9062);
nor U9892 (N_9892,N_9085,N_9110);
or U9893 (N_9893,N_9037,N_9204);
nor U9894 (N_9894,N_9023,N_9392);
and U9895 (N_9895,N_9432,N_9465);
and U9896 (N_9896,N_9190,N_9326);
and U9897 (N_9897,N_9140,N_9101);
nand U9898 (N_9898,N_9284,N_9419);
xor U9899 (N_9899,N_9171,N_9167);
nand U9900 (N_9900,N_9078,N_9280);
nand U9901 (N_9901,N_9087,N_9241);
nor U9902 (N_9902,N_9064,N_9349);
nor U9903 (N_9903,N_9264,N_9177);
nor U9904 (N_9904,N_9445,N_9057);
nor U9905 (N_9905,N_9358,N_9272);
and U9906 (N_9906,N_9161,N_9073);
nand U9907 (N_9907,N_9423,N_9424);
and U9908 (N_9908,N_9270,N_9085);
or U9909 (N_9909,N_9198,N_9429);
and U9910 (N_9910,N_9395,N_9300);
xnor U9911 (N_9911,N_9215,N_9229);
nor U9912 (N_9912,N_9105,N_9050);
or U9913 (N_9913,N_9089,N_9401);
or U9914 (N_9914,N_9466,N_9389);
nand U9915 (N_9915,N_9089,N_9448);
and U9916 (N_9916,N_9445,N_9128);
nor U9917 (N_9917,N_9356,N_9384);
nand U9918 (N_9918,N_9356,N_9380);
nor U9919 (N_9919,N_9279,N_9438);
nand U9920 (N_9920,N_9484,N_9280);
and U9921 (N_9921,N_9414,N_9077);
nor U9922 (N_9922,N_9217,N_9297);
or U9923 (N_9923,N_9459,N_9271);
nor U9924 (N_9924,N_9067,N_9125);
nor U9925 (N_9925,N_9000,N_9247);
or U9926 (N_9926,N_9237,N_9110);
nand U9927 (N_9927,N_9038,N_9255);
xor U9928 (N_9928,N_9490,N_9133);
and U9929 (N_9929,N_9441,N_9130);
and U9930 (N_9930,N_9130,N_9168);
xor U9931 (N_9931,N_9201,N_9234);
and U9932 (N_9932,N_9019,N_9060);
nor U9933 (N_9933,N_9469,N_9222);
nor U9934 (N_9934,N_9177,N_9010);
xor U9935 (N_9935,N_9085,N_9258);
and U9936 (N_9936,N_9052,N_9310);
and U9937 (N_9937,N_9184,N_9365);
nand U9938 (N_9938,N_9418,N_9006);
or U9939 (N_9939,N_9262,N_9357);
or U9940 (N_9940,N_9391,N_9079);
xnor U9941 (N_9941,N_9468,N_9107);
nand U9942 (N_9942,N_9008,N_9496);
xor U9943 (N_9943,N_9459,N_9136);
and U9944 (N_9944,N_9225,N_9249);
and U9945 (N_9945,N_9378,N_9020);
and U9946 (N_9946,N_9238,N_9456);
and U9947 (N_9947,N_9371,N_9348);
nor U9948 (N_9948,N_9307,N_9334);
nand U9949 (N_9949,N_9456,N_9005);
nor U9950 (N_9950,N_9210,N_9259);
xnor U9951 (N_9951,N_9049,N_9206);
nor U9952 (N_9952,N_9189,N_9143);
and U9953 (N_9953,N_9447,N_9300);
or U9954 (N_9954,N_9159,N_9400);
nor U9955 (N_9955,N_9052,N_9118);
and U9956 (N_9956,N_9006,N_9009);
or U9957 (N_9957,N_9478,N_9472);
xnor U9958 (N_9958,N_9230,N_9259);
nor U9959 (N_9959,N_9126,N_9121);
nor U9960 (N_9960,N_9162,N_9046);
nor U9961 (N_9961,N_9467,N_9014);
nor U9962 (N_9962,N_9459,N_9415);
and U9963 (N_9963,N_9451,N_9115);
or U9964 (N_9964,N_9040,N_9099);
or U9965 (N_9965,N_9098,N_9358);
and U9966 (N_9966,N_9290,N_9425);
xor U9967 (N_9967,N_9114,N_9106);
and U9968 (N_9968,N_9275,N_9463);
nand U9969 (N_9969,N_9413,N_9095);
nand U9970 (N_9970,N_9476,N_9163);
xnor U9971 (N_9971,N_9144,N_9403);
xnor U9972 (N_9972,N_9292,N_9283);
nor U9973 (N_9973,N_9024,N_9047);
xor U9974 (N_9974,N_9178,N_9224);
xor U9975 (N_9975,N_9446,N_9023);
and U9976 (N_9976,N_9010,N_9049);
and U9977 (N_9977,N_9382,N_9481);
nor U9978 (N_9978,N_9282,N_9291);
and U9979 (N_9979,N_9034,N_9011);
nor U9980 (N_9980,N_9464,N_9060);
and U9981 (N_9981,N_9482,N_9353);
nand U9982 (N_9982,N_9238,N_9054);
and U9983 (N_9983,N_9458,N_9487);
xor U9984 (N_9984,N_9244,N_9499);
and U9985 (N_9985,N_9338,N_9474);
xnor U9986 (N_9986,N_9116,N_9396);
nand U9987 (N_9987,N_9347,N_9247);
nor U9988 (N_9988,N_9257,N_9457);
nor U9989 (N_9989,N_9347,N_9210);
or U9990 (N_9990,N_9088,N_9189);
xnor U9991 (N_9991,N_9297,N_9031);
or U9992 (N_9992,N_9092,N_9279);
nand U9993 (N_9993,N_9247,N_9037);
and U9994 (N_9994,N_9046,N_9399);
nand U9995 (N_9995,N_9096,N_9085);
and U9996 (N_9996,N_9043,N_9175);
xor U9997 (N_9997,N_9213,N_9263);
and U9998 (N_9998,N_9220,N_9013);
nand U9999 (N_9999,N_9182,N_9010);
xnor U10000 (N_10000,N_9551,N_9723);
xor U10001 (N_10001,N_9908,N_9837);
xnor U10002 (N_10002,N_9813,N_9883);
xnor U10003 (N_10003,N_9943,N_9787);
nand U10004 (N_10004,N_9713,N_9934);
and U10005 (N_10005,N_9754,N_9718);
nor U10006 (N_10006,N_9566,N_9931);
nor U10007 (N_10007,N_9673,N_9796);
and U10008 (N_10008,N_9812,N_9563);
nand U10009 (N_10009,N_9638,N_9579);
or U10010 (N_10010,N_9657,N_9568);
xor U10011 (N_10011,N_9573,N_9732);
and U10012 (N_10012,N_9710,N_9532);
and U10013 (N_10013,N_9535,N_9800);
xnor U10014 (N_10014,N_9917,N_9916);
or U10015 (N_10015,N_9819,N_9741);
xnor U10016 (N_10016,N_9761,N_9988);
nand U10017 (N_10017,N_9697,N_9544);
xnor U10018 (N_10018,N_9504,N_9767);
and U10019 (N_10019,N_9817,N_9788);
nand U10020 (N_10020,N_9963,N_9832);
and U10021 (N_10021,N_9882,N_9696);
xor U10022 (N_10022,N_9654,N_9869);
and U10023 (N_10023,N_9996,N_9990);
nand U10024 (N_10024,N_9584,N_9958);
or U10025 (N_10025,N_9550,N_9711);
nand U10026 (N_10026,N_9685,N_9726);
and U10027 (N_10027,N_9811,N_9627);
or U10028 (N_10028,N_9605,N_9871);
or U10029 (N_10029,N_9738,N_9892);
nand U10030 (N_10030,N_9938,N_9665);
and U10031 (N_10031,N_9851,N_9625);
or U10032 (N_10032,N_9778,N_9602);
or U10033 (N_10033,N_9828,N_9528);
or U10034 (N_10034,N_9588,N_9846);
and U10035 (N_10035,N_9976,N_9631);
nor U10036 (N_10036,N_9652,N_9595);
xor U10037 (N_10037,N_9860,N_9699);
nand U10038 (N_10038,N_9742,N_9896);
and U10039 (N_10039,N_9825,N_9609);
xor U10040 (N_10040,N_9799,N_9607);
or U10041 (N_10041,N_9666,N_9816);
and U10042 (N_10042,N_9914,N_9777);
and U10043 (N_10043,N_9518,N_9868);
xnor U10044 (N_10044,N_9630,N_9601);
or U10045 (N_10045,N_9972,N_9591);
nor U10046 (N_10046,N_9590,N_9983);
or U10047 (N_10047,N_9542,N_9692);
and U10048 (N_10048,N_9875,N_9626);
xor U10049 (N_10049,N_9939,N_9569);
or U10050 (N_10050,N_9597,N_9715);
or U10051 (N_10051,N_9929,N_9617);
and U10052 (N_10052,N_9753,N_9893);
or U10053 (N_10053,N_9651,N_9596);
and U10054 (N_10054,N_9768,N_9744);
nor U10055 (N_10055,N_9992,N_9621);
nor U10056 (N_10056,N_9920,N_9945);
nand U10057 (N_10057,N_9689,N_9783);
and U10058 (N_10058,N_9520,N_9580);
or U10059 (N_10059,N_9526,N_9684);
xor U10060 (N_10060,N_9884,N_9806);
xnor U10061 (N_10061,N_9881,N_9556);
xnor U10062 (N_10062,N_9946,N_9629);
xnor U10063 (N_10063,N_9575,N_9640);
xnor U10064 (N_10064,N_9781,N_9865);
xnor U10065 (N_10065,N_9856,N_9949);
nand U10066 (N_10066,N_9915,N_9815);
xnor U10067 (N_10067,N_9564,N_9690);
or U10068 (N_10068,N_9858,N_9735);
or U10069 (N_10069,N_9606,N_9801);
nor U10070 (N_10070,N_9863,N_9903);
and U10071 (N_10071,N_9681,N_9775);
or U10072 (N_10072,N_9834,N_9969);
nand U10073 (N_10073,N_9608,N_9758);
and U10074 (N_10074,N_9864,N_9786);
xor U10075 (N_10075,N_9951,N_9529);
xnor U10076 (N_10076,N_9862,N_9933);
nor U10077 (N_10077,N_9513,N_9734);
nand U10078 (N_10078,N_9913,N_9663);
or U10079 (N_10079,N_9502,N_9537);
nor U10080 (N_10080,N_9760,N_9516);
or U10081 (N_10081,N_9857,N_9805);
xnor U10082 (N_10082,N_9780,N_9633);
xor U10083 (N_10083,N_9910,N_9872);
or U10084 (N_10084,N_9867,N_9534);
xor U10085 (N_10085,N_9680,N_9838);
and U10086 (N_10086,N_9912,N_9978);
nand U10087 (N_10087,N_9600,N_9772);
nand U10088 (N_10088,N_9733,N_9888);
nor U10089 (N_10089,N_9662,N_9512);
nand U10090 (N_10090,N_9674,N_9682);
xnor U10091 (N_10091,N_9672,N_9507);
nand U10092 (N_10092,N_9902,N_9506);
xor U10093 (N_10093,N_9759,N_9552);
xor U10094 (N_10094,N_9950,N_9519);
xnor U10095 (N_10095,N_9647,N_9764);
nand U10096 (N_10096,N_9527,N_9802);
xor U10097 (N_10097,N_9536,N_9740);
and U10098 (N_10098,N_9611,N_9848);
xnor U10099 (N_10099,N_9830,N_9918);
xor U10100 (N_10100,N_9706,N_9982);
xnor U10101 (N_10101,N_9968,N_9948);
xnor U10102 (N_10102,N_9879,N_9712);
or U10103 (N_10103,N_9642,N_9986);
nor U10104 (N_10104,N_9501,N_9720);
nand U10105 (N_10105,N_9545,N_9930);
xnor U10106 (N_10106,N_9668,N_9622);
xnor U10107 (N_10107,N_9687,N_9667);
nand U10108 (N_10108,N_9708,N_9826);
xor U10109 (N_10109,N_9547,N_9905);
or U10110 (N_10110,N_9581,N_9671);
xnor U10111 (N_10111,N_9843,N_9889);
nor U10112 (N_10112,N_9750,N_9618);
xor U10113 (N_10113,N_9653,N_9936);
nor U10114 (N_10114,N_9897,N_9840);
or U10115 (N_10115,N_9559,N_9603);
nand U10116 (N_10116,N_9558,N_9731);
nor U10117 (N_10117,N_9586,N_9702);
and U10118 (N_10118,N_9739,N_9904);
and U10119 (N_10119,N_9818,N_9831);
or U10120 (N_10120,N_9533,N_9984);
or U10121 (N_10121,N_9679,N_9909);
nor U10122 (N_10122,N_9967,N_9779);
xor U10123 (N_10123,N_9895,N_9954);
and U10124 (N_10124,N_9798,N_9604);
nand U10125 (N_10125,N_9511,N_9704);
or U10126 (N_10126,N_9574,N_9981);
and U10127 (N_10127,N_9925,N_9947);
and U10128 (N_10128,N_9922,N_9694);
and U10129 (N_10129,N_9634,N_9661);
nand U10130 (N_10130,N_9521,N_9751);
xnor U10131 (N_10131,N_9845,N_9729);
nand U10132 (N_10132,N_9850,N_9941);
xnor U10133 (N_10133,N_9530,N_9782);
or U10134 (N_10134,N_9635,N_9899);
or U10135 (N_10135,N_9911,N_9900);
and U10136 (N_10136,N_9898,N_9999);
or U10137 (N_10137,N_9553,N_9649);
and U10138 (N_10138,N_9847,N_9944);
xor U10139 (N_10139,N_9686,N_9646);
and U10140 (N_10140,N_9560,N_9567);
nand U10141 (N_10141,N_9614,N_9565);
or U10142 (N_10142,N_9525,N_9612);
nand U10143 (N_10143,N_9763,N_9940);
xnor U10144 (N_10144,N_9628,N_9876);
and U10145 (N_10145,N_9790,N_9926);
nor U10146 (N_10146,N_9698,N_9906);
nor U10147 (N_10147,N_9613,N_9776);
nor U10148 (N_10148,N_9745,N_9980);
nand U10149 (N_10149,N_9594,N_9773);
nand U10150 (N_10150,N_9757,N_9921);
nor U10151 (N_10151,N_9998,N_9578);
or U10152 (N_10152,N_9991,N_9548);
or U10153 (N_10153,N_9874,N_9890);
nand U10154 (N_10154,N_9887,N_9994);
nand U10155 (N_10155,N_9861,N_9656);
xnor U10156 (N_10156,N_9693,N_9844);
and U10157 (N_10157,N_9873,N_9823);
and U10158 (N_10158,N_9774,N_9932);
nand U10159 (N_10159,N_9645,N_9599);
or U10160 (N_10160,N_9620,N_9624);
nor U10161 (N_10161,N_9765,N_9695);
and U10162 (N_10162,N_9769,N_9770);
nor U10163 (N_10163,N_9880,N_9549);
nor U10164 (N_10164,N_9971,N_9508);
or U10165 (N_10165,N_9877,N_9531);
or U10166 (N_10166,N_9808,N_9570);
or U10167 (N_10167,N_9705,N_9966);
xnor U10168 (N_10168,N_9919,N_9655);
nor U10169 (N_10169,N_9928,N_9736);
or U10170 (N_10170,N_9700,N_9854);
nor U10171 (N_10171,N_9722,N_9514);
xnor U10172 (N_10172,N_9814,N_9554);
or U10173 (N_10173,N_9730,N_9648);
and U10174 (N_10174,N_9853,N_9956);
and U10175 (N_10175,N_9987,N_9632);
and U10176 (N_10176,N_9503,N_9855);
and U10177 (N_10177,N_9678,N_9737);
or U10178 (N_10178,N_9809,N_9576);
and U10179 (N_10179,N_9952,N_9541);
and U10180 (N_10180,N_9641,N_9789);
and U10181 (N_10181,N_9747,N_9650);
nand U10182 (N_10182,N_9619,N_9561);
xor U10183 (N_10183,N_9820,N_9794);
or U10184 (N_10184,N_9571,N_9785);
nand U10185 (N_10185,N_9791,N_9979);
nand U10186 (N_10186,N_9658,N_9637);
xor U10187 (N_10187,N_9993,N_9539);
nor U10188 (N_10188,N_9803,N_9821);
nand U10189 (N_10189,N_9623,N_9746);
or U10190 (N_10190,N_9749,N_9517);
xor U10191 (N_10191,N_9995,N_9510);
and U10192 (N_10192,N_9886,N_9885);
nand U10193 (N_10193,N_9644,N_9725);
nand U10194 (N_10194,N_9859,N_9582);
xor U10195 (N_10195,N_9962,N_9555);
xnor U10196 (N_10196,N_9839,N_9701);
nand U10197 (N_10197,N_9959,N_9810);
or U10198 (N_10198,N_9974,N_9676);
xor U10199 (N_10199,N_9543,N_9636);
xor U10200 (N_10200,N_9538,N_9822);
and U10201 (N_10201,N_9792,N_9827);
nor U10202 (N_10202,N_9975,N_9804);
or U10203 (N_10203,N_9714,N_9748);
and U10204 (N_10204,N_9577,N_9557);
and U10205 (N_10205,N_9670,N_9522);
nor U10206 (N_10206,N_9664,N_9841);
nor U10207 (N_10207,N_9942,N_9500);
and U10208 (N_10208,N_9572,N_9585);
or U10209 (N_10209,N_9953,N_9610);
or U10210 (N_10210,N_9546,N_9593);
xnor U10211 (N_10211,N_9756,N_9515);
and U10212 (N_10212,N_9707,N_9784);
xor U10213 (N_10213,N_9955,N_9795);
nand U10214 (N_10214,N_9894,N_9957);
nor U10215 (N_10215,N_9961,N_9719);
nor U10216 (N_10216,N_9709,N_9524);
or U10217 (N_10217,N_9562,N_9977);
and U10218 (N_10218,N_9509,N_9836);
or U10219 (N_10219,N_9639,N_9935);
and U10220 (N_10220,N_9824,N_9937);
or U10221 (N_10221,N_9835,N_9970);
nor U10222 (N_10222,N_9523,N_9771);
and U10223 (N_10223,N_9583,N_9829);
nor U10224 (N_10224,N_9587,N_9589);
or U10225 (N_10225,N_9660,N_9870);
and U10226 (N_10226,N_9592,N_9766);
and U10227 (N_10227,N_9960,N_9807);
nor U10228 (N_10228,N_9762,N_9965);
nand U10229 (N_10229,N_9683,N_9677);
nand U10230 (N_10230,N_9616,N_9891);
or U10231 (N_10231,N_9727,N_9743);
nand U10232 (N_10232,N_9721,N_9669);
and U10233 (N_10233,N_9907,N_9755);
or U10234 (N_10234,N_9643,N_9615);
nand U10235 (N_10235,N_9973,N_9964);
and U10236 (N_10236,N_9716,N_9985);
and U10237 (N_10237,N_9923,N_9717);
or U10238 (N_10238,N_9833,N_9724);
or U10239 (N_10239,N_9659,N_9797);
or U10240 (N_10240,N_9752,N_9989);
nor U10241 (N_10241,N_9540,N_9849);
or U10242 (N_10242,N_9852,N_9793);
nand U10243 (N_10243,N_9997,N_9598);
nor U10244 (N_10244,N_9691,N_9901);
nor U10245 (N_10245,N_9675,N_9728);
and U10246 (N_10246,N_9703,N_9866);
nand U10247 (N_10247,N_9505,N_9688);
nor U10248 (N_10248,N_9878,N_9924);
nor U10249 (N_10249,N_9927,N_9842);
nor U10250 (N_10250,N_9606,N_9817);
nor U10251 (N_10251,N_9972,N_9973);
and U10252 (N_10252,N_9652,N_9506);
nand U10253 (N_10253,N_9529,N_9969);
or U10254 (N_10254,N_9515,N_9722);
nand U10255 (N_10255,N_9796,N_9617);
or U10256 (N_10256,N_9892,N_9712);
and U10257 (N_10257,N_9818,N_9539);
nor U10258 (N_10258,N_9848,N_9514);
or U10259 (N_10259,N_9552,N_9571);
nor U10260 (N_10260,N_9515,N_9819);
nor U10261 (N_10261,N_9703,N_9647);
xnor U10262 (N_10262,N_9669,N_9608);
nand U10263 (N_10263,N_9862,N_9726);
nor U10264 (N_10264,N_9529,N_9721);
xor U10265 (N_10265,N_9508,N_9512);
nand U10266 (N_10266,N_9790,N_9879);
or U10267 (N_10267,N_9760,N_9706);
and U10268 (N_10268,N_9934,N_9896);
or U10269 (N_10269,N_9945,N_9997);
nand U10270 (N_10270,N_9587,N_9702);
xor U10271 (N_10271,N_9524,N_9708);
and U10272 (N_10272,N_9556,N_9883);
or U10273 (N_10273,N_9650,N_9971);
or U10274 (N_10274,N_9694,N_9894);
or U10275 (N_10275,N_9639,N_9507);
or U10276 (N_10276,N_9509,N_9540);
or U10277 (N_10277,N_9643,N_9572);
nor U10278 (N_10278,N_9887,N_9638);
nor U10279 (N_10279,N_9714,N_9552);
and U10280 (N_10280,N_9908,N_9745);
nor U10281 (N_10281,N_9686,N_9987);
nand U10282 (N_10282,N_9539,N_9948);
or U10283 (N_10283,N_9890,N_9961);
nand U10284 (N_10284,N_9855,N_9532);
nand U10285 (N_10285,N_9649,N_9516);
xnor U10286 (N_10286,N_9640,N_9790);
xor U10287 (N_10287,N_9847,N_9689);
nand U10288 (N_10288,N_9956,N_9575);
xnor U10289 (N_10289,N_9984,N_9835);
and U10290 (N_10290,N_9885,N_9994);
or U10291 (N_10291,N_9806,N_9849);
and U10292 (N_10292,N_9575,N_9564);
xor U10293 (N_10293,N_9524,N_9536);
nor U10294 (N_10294,N_9678,N_9643);
nor U10295 (N_10295,N_9667,N_9750);
nor U10296 (N_10296,N_9983,N_9540);
nor U10297 (N_10297,N_9931,N_9542);
nor U10298 (N_10298,N_9731,N_9604);
nand U10299 (N_10299,N_9994,N_9637);
or U10300 (N_10300,N_9870,N_9908);
and U10301 (N_10301,N_9628,N_9749);
nor U10302 (N_10302,N_9823,N_9512);
nand U10303 (N_10303,N_9548,N_9860);
xnor U10304 (N_10304,N_9607,N_9834);
and U10305 (N_10305,N_9747,N_9576);
or U10306 (N_10306,N_9596,N_9575);
nor U10307 (N_10307,N_9957,N_9908);
xnor U10308 (N_10308,N_9923,N_9527);
and U10309 (N_10309,N_9630,N_9658);
xor U10310 (N_10310,N_9726,N_9534);
xor U10311 (N_10311,N_9772,N_9751);
nor U10312 (N_10312,N_9646,N_9517);
and U10313 (N_10313,N_9702,N_9840);
or U10314 (N_10314,N_9946,N_9892);
xnor U10315 (N_10315,N_9856,N_9616);
or U10316 (N_10316,N_9537,N_9529);
nor U10317 (N_10317,N_9716,N_9910);
nor U10318 (N_10318,N_9749,N_9980);
nor U10319 (N_10319,N_9527,N_9821);
nor U10320 (N_10320,N_9757,N_9675);
xor U10321 (N_10321,N_9671,N_9867);
xor U10322 (N_10322,N_9959,N_9585);
nand U10323 (N_10323,N_9637,N_9696);
nand U10324 (N_10324,N_9604,N_9903);
nor U10325 (N_10325,N_9788,N_9985);
or U10326 (N_10326,N_9820,N_9904);
or U10327 (N_10327,N_9905,N_9676);
xor U10328 (N_10328,N_9521,N_9579);
and U10329 (N_10329,N_9571,N_9761);
nor U10330 (N_10330,N_9575,N_9699);
or U10331 (N_10331,N_9937,N_9841);
nand U10332 (N_10332,N_9823,N_9520);
xnor U10333 (N_10333,N_9977,N_9546);
and U10334 (N_10334,N_9728,N_9775);
and U10335 (N_10335,N_9947,N_9780);
xnor U10336 (N_10336,N_9975,N_9926);
nand U10337 (N_10337,N_9537,N_9934);
nand U10338 (N_10338,N_9877,N_9980);
xor U10339 (N_10339,N_9563,N_9713);
or U10340 (N_10340,N_9829,N_9657);
nor U10341 (N_10341,N_9660,N_9525);
and U10342 (N_10342,N_9657,N_9612);
and U10343 (N_10343,N_9959,N_9884);
nor U10344 (N_10344,N_9698,N_9814);
nand U10345 (N_10345,N_9890,N_9981);
nor U10346 (N_10346,N_9739,N_9515);
nor U10347 (N_10347,N_9790,N_9615);
and U10348 (N_10348,N_9618,N_9754);
nor U10349 (N_10349,N_9870,N_9532);
or U10350 (N_10350,N_9866,N_9801);
xnor U10351 (N_10351,N_9990,N_9536);
nand U10352 (N_10352,N_9839,N_9761);
or U10353 (N_10353,N_9521,N_9736);
nand U10354 (N_10354,N_9777,N_9561);
nand U10355 (N_10355,N_9764,N_9890);
nand U10356 (N_10356,N_9817,N_9665);
nand U10357 (N_10357,N_9502,N_9571);
nand U10358 (N_10358,N_9872,N_9783);
nor U10359 (N_10359,N_9998,N_9660);
xnor U10360 (N_10360,N_9836,N_9911);
nand U10361 (N_10361,N_9537,N_9808);
or U10362 (N_10362,N_9567,N_9842);
nand U10363 (N_10363,N_9624,N_9543);
and U10364 (N_10364,N_9557,N_9991);
and U10365 (N_10365,N_9901,N_9553);
xnor U10366 (N_10366,N_9697,N_9866);
nor U10367 (N_10367,N_9921,N_9846);
or U10368 (N_10368,N_9571,N_9555);
and U10369 (N_10369,N_9933,N_9829);
xnor U10370 (N_10370,N_9531,N_9842);
or U10371 (N_10371,N_9561,N_9598);
nand U10372 (N_10372,N_9794,N_9847);
nor U10373 (N_10373,N_9954,N_9572);
nand U10374 (N_10374,N_9513,N_9814);
and U10375 (N_10375,N_9558,N_9674);
nand U10376 (N_10376,N_9895,N_9731);
or U10377 (N_10377,N_9793,N_9927);
or U10378 (N_10378,N_9858,N_9524);
or U10379 (N_10379,N_9760,N_9751);
nand U10380 (N_10380,N_9697,N_9869);
or U10381 (N_10381,N_9855,N_9971);
xor U10382 (N_10382,N_9965,N_9626);
nor U10383 (N_10383,N_9855,N_9912);
xor U10384 (N_10384,N_9520,N_9840);
nand U10385 (N_10385,N_9553,N_9640);
nand U10386 (N_10386,N_9636,N_9533);
or U10387 (N_10387,N_9568,N_9643);
and U10388 (N_10388,N_9759,N_9609);
xor U10389 (N_10389,N_9823,N_9554);
nor U10390 (N_10390,N_9961,N_9665);
nor U10391 (N_10391,N_9744,N_9685);
and U10392 (N_10392,N_9719,N_9545);
and U10393 (N_10393,N_9874,N_9589);
xor U10394 (N_10394,N_9947,N_9512);
xor U10395 (N_10395,N_9647,N_9847);
xnor U10396 (N_10396,N_9872,N_9584);
xnor U10397 (N_10397,N_9993,N_9514);
nand U10398 (N_10398,N_9955,N_9555);
xnor U10399 (N_10399,N_9566,N_9746);
nand U10400 (N_10400,N_9797,N_9898);
or U10401 (N_10401,N_9992,N_9763);
xnor U10402 (N_10402,N_9611,N_9623);
nor U10403 (N_10403,N_9545,N_9879);
nand U10404 (N_10404,N_9910,N_9607);
and U10405 (N_10405,N_9599,N_9624);
nor U10406 (N_10406,N_9502,N_9909);
or U10407 (N_10407,N_9597,N_9828);
and U10408 (N_10408,N_9583,N_9730);
and U10409 (N_10409,N_9585,N_9971);
xnor U10410 (N_10410,N_9754,N_9904);
xnor U10411 (N_10411,N_9875,N_9963);
and U10412 (N_10412,N_9711,N_9660);
xnor U10413 (N_10413,N_9996,N_9875);
or U10414 (N_10414,N_9544,N_9730);
or U10415 (N_10415,N_9662,N_9766);
xor U10416 (N_10416,N_9773,N_9758);
or U10417 (N_10417,N_9973,N_9851);
and U10418 (N_10418,N_9721,N_9646);
xnor U10419 (N_10419,N_9849,N_9867);
or U10420 (N_10420,N_9671,N_9760);
nand U10421 (N_10421,N_9624,N_9589);
nor U10422 (N_10422,N_9835,N_9826);
and U10423 (N_10423,N_9600,N_9922);
nand U10424 (N_10424,N_9655,N_9694);
nor U10425 (N_10425,N_9505,N_9576);
xor U10426 (N_10426,N_9930,N_9537);
and U10427 (N_10427,N_9774,N_9730);
or U10428 (N_10428,N_9925,N_9575);
or U10429 (N_10429,N_9727,N_9853);
and U10430 (N_10430,N_9896,N_9624);
nor U10431 (N_10431,N_9701,N_9793);
nand U10432 (N_10432,N_9969,N_9972);
and U10433 (N_10433,N_9513,N_9588);
nor U10434 (N_10434,N_9647,N_9983);
or U10435 (N_10435,N_9688,N_9681);
xor U10436 (N_10436,N_9845,N_9632);
and U10437 (N_10437,N_9787,N_9608);
nor U10438 (N_10438,N_9927,N_9574);
or U10439 (N_10439,N_9782,N_9524);
nor U10440 (N_10440,N_9860,N_9901);
or U10441 (N_10441,N_9962,N_9744);
nand U10442 (N_10442,N_9829,N_9728);
and U10443 (N_10443,N_9910,N_9900);
nand U10444 (N_10444,N_9625,N_9885);
or U10445 (N_10445,N_9725,N_9534);
xor U10446 (N_10446,N_9520,N_9624);
or U10447 (N_10447,N_9535,N_9778);
or U10448 (N_10448,N_9575,N_9620);
and U10449 (N_10449,N_9550,N_9964);
or U10450 (N_10450,N_9719,N_9534);
nand U10451 (N_10451,N_9521,N_9792);
and U10452 (N_10452,N_9712,N_9949);
and U10453 (N_10453,N_9969,N_9787);
and U10454 (N_10454,N_9534,N_9754);
xor U10455 (N_10455,N_9527,N_9716);
and U10456 (N_10456,N_9948,N_9915);
xor U10457 (N_10457,N_9714,N_9730);
nor U10458 (N_10458,N_9811,N_9594);
and U10459 (N_10459,N_9717,N_9649);
nand U10460 (N_10460,N_9929,N_9582);
and U10461 (N_10461,N_9585,N_9693);
xnor U10462 (N_10462,N_9973,N_9657);
xnor U10463 (N_10463,N_9745,N_9656);
and U10464 (N_10464,N_9954,N_9930);
nand U10465 (N_10465,N_9857,N_9530);
nor U10466 (N_10466,N_9673,N_9953);
nand U10467 (N_10467,N_9764,N_9536);
nand U10468 (N_10468,N_9674,N_9735);
nand U10469 (N_10469,N_9991,N_9730);
or U10470 (N_10470,N_9860,N_9642);
or U10471 (N_10471,N_9726,N_9750);
or U10472 (N_10472,N_9932,N_9720);
nand U10473 (N_10473,N_9819,N_9604);
or U10474 (N_10474,N_9519,N_9687);
or U10475 (N_10475,N_9814,N_9961);
xnor U10476 (N_10476,N_9870,N_9620);
nor U10477 (N_10477,N_9979,N_9749);
or U10478 (N_10478,N_9962,N_9748);
nor U10479 (N_10479,N_9824,N_9972);
xnor U10480 (N_10480,N_9667,N_9643);
or U10481 (N_10481,N_9735,N_9763);
xor U10482 (N_10482,N_9991,N_9618);
and U10483 (N_10483,N_9992,N_9613);
xnor U10484 (N_10484,N_9967,N_9995);
nand U10485 (N_10485,N_9521,N_9682);
or U10486 (N_10486,N_9532,N_9567);
or U10487 (N_10487,N_9740,N_9734);
nand U10488 (N_10488,N_9578,N_9987);
and U10489 (N_10489,N_9694,N_9906);
or U10490 (N_10490,N_9681,N_9662);
nor U10491 (N_10491,N_9886,N_9952);
or U10492 (N_10492,N_9624,N_9584);
or U10493 (N_10493,N_9698,N_9987);
nand U10494 (N_10494,N_9836,N_9706);
nor U10495 (N_10495,N_9896,N_9958);
and U10496 (N_10496,N_9918,N_9930);
nand U10497 (N_10497,N_9543,N_9844);
and U10498 (N_10498,N_9803,N_9864);
nor U10499 (N_10499,N_9949,N_9703);
nor U10500 (N_10500,N_10072,N_10482);
and U10501 (N_10501,N_10127,N_10208);
xnor U10502 (N_10502,N_10119,N_10252);
xnor U10503 (N_10503,N_10367,N_10013);
xnor U10504 (N_10504,N_10408,N_10118);
or U10505 (N_10505,N_10128,N_10368);
and U10506 (N_10506,N_10170,N_10328);
nor U10507 (N_10507,N_10182,N_10176);
xor U10508 (N_10508,N_10438,N_10432);
or U10509 (N_10509,N_10452,N_10455);
nor U10510 (N_10510,N_10010,N_10281);
nand U10511 (N_10511,N_10371,N_10166);
and U10512 (N_10512,N_10487,N_10456);
or U10513 (N_10513,N_10384,N_10388);
nor U10514 (N_10514,N_10261,N_10011);
and U10515 (N_10515,N_10038,N_10308);
nand U10516 (N_10516,N_10226,N_10116);
xnor U10517 (N_10517,N_10242,N_10447);
or U10518 (N_10518,N_10258,N_10167);
or U10519 (N_10519,N_10077,N_10472);
xor U10520 (N_10520,N_10414,N_10496);
xnor U10521 (N_10521,N_10099,N_10131);
and U10522 (N_10522,N_10022,N_10295);
nand U10523 (N_10523,N_10468,N_10085);
and U10524 (N_10524,N_10331,N_10179);
xor U10525 (N_10525,N_10039,N_10255);
xnor U10526 (N_10526,N_10104,N_10177);
xnor U10527 (N_10527,N_10494,N_10370);
xnor U10528 (N_10528,N_10398,N_10112);
xnor U10529 (N_10529,N_10274,N_10441);
or U10530 (N_10530,N_10093,N_10443);
or U10531 (N_10531,N_10339,N_10479);
xor U10532 (N_10532,N_10428,N_10307);
nand U10533 (N_10533,N_10098,N_10490);
xor U10534 (N_10534,N_10366,N_10068);
xnor U10535 (N_10535,N_10312,N_10136);
nor U10536 (N_10536,N_10042,N_10195);
nor U10537 (N_10537,N_10287,N_10376);
or U10538 (N_10538,N_10288,N_10125);
nand U10539 (N_10539,N_10427,N_10188);
and U10540 (N_10540,N_10257,N_10431);
xnor U10541 (N_10541,N_10092,N_10411);
nor U10542 (N_10542,N_10240,N_10083);
nor U10543 (N_10543,N_10107,N_10016);
and U10544 (N_10544,N_10251,N_10269);
and U10545 (N_10545,N_10346,N_10007);
nor U10546 (N_10546,N_10140,N_10478);
nor U10547 (N_10547,N_10306,N_10142);
nand U10548 (N_10548,N_10230,N_10027);
nor U10549 (N_10549,N_10043,N_10461);
and U10550 (N_10550,N_10459,N_10154);
xor U10551 (N_10551,N_10259,N_10201);
xnor U10552 (N_10552,N_10066,N_10397);
and U10553 (N_10553,N_10160,N_10265);
and U10554 (N_10554,N_10117,N_10101);
nor U10555 (N_10555,N_10173,N_10451);
and U10556 (N_10556,N_10164,N_10489);
nor U10557 (N_10557,N_10148,N_10363);
nand U10558 (N_10558,N_10227,N_10151);
or U10559 (N_10559,N_10033,N_10350);
nand U10560 (N_10560,N_10285,N_10467);
nor U10561 (N_10561,N_10190,N_10152);
xor U10562 (N_10562,N_10061,N_10364);
or U10563 (N_10563,N_10053,N_10215);
xnor U10564 (N_10564,N_10374,N_10480);
xnor U10565 (N_10565,N_10224,N_10492);
xor U10566 (N_10566,N_10020,N_10426);
nor U10567 (N_10567,N_10395,N_10229);
and U10568 (N_10568,N_10041,N_10294);
nor U10569 (N_10569,N_10143,N_10423);
and U10570 (N_10570,N_10214,N_10425);
xor U10571 (N_10571,N_10354,N_10194);
and U10572 (N_10572,N_10162,N_10028);
nand U10573 (N_10573,N_10005,N_10361);
nand U10574 (N_10574,N_10442,N_10341);
or U10575 (N_10575,N_10440,N_10336);
xnor U10576 (N_10576,N_10416,N_10037);
xor U10577 (N_10577,N_10199,N_10197);
and U10578 (N_10578,N_10279,N_10181);
nor U10579 (N_10579,N_10134,N_10175);
or U10580 (N_10580,N_10052,N_10246);
nor U10581 (N_10581,N_10163,N_10169);
and U10582 (N_10582,N_10453,N_10244);
nor U10583 (N_10583,N_10067,N_10129);
and U10584 (N_10584,N_10087,N_10120);
xor U10585 (N_10585,N_10450,N_10130);
xnor U10586 (N_10586,N_10198,N_10015);
xor U10587 (N_10587,N_10114,N_10298);
or U10588 (N_10588,N_10156,N_10111);
nor U10589 (N_10589,N_10218,N_10260);
xnor U10590 (N_10590,N_10399,N_10051);
or U10591 (N_10591,N_10171,N_10436);
nor U10592 (N_10592,N_10221,N_10219);
and U10593 (N_10593,N_10365,N_10109);
nor U10594 (N_10594,N_10059,N_10222);
and U10595 (N_10595,N_10437,N_10132);
nand U10596 (N_10596,N_10406,N_10139);
nor U10597 (N_10597,N_10330,N_10446);
xnor U10598 (N_10598,N_10311,N_10345);
nor U10599 (N_10599,N_10250,N_10233);
or U10600 (N_10600,N_10385,N_10123);
or U10601 (N_10601,N_10122,N_10338);
or U10602 (N_10602,N_10393,N_10046);
or U10603 (N_10603,N_10031,N_10073);
or U10604 (N_10604,N_10324,N_10486);
nand U10605 (N_10605,N_10323,N_10084);
xor U10606 (N_10606,N_10014,N_10469);
nand U10607 (N_10607,N_10373,N_10238);
or U10608 (N_10608,N_10090,N_10054);
xnor U10609 (N_10609,N_10212,N_10445);
nor U10610 (N_10610,N_10124,N_10493);
nor U10611 (N_10611,N_10006,N_10065);
xnor U10612 (N_10612,N_10348,N_10483);
and U10613 (N_10613,N_10351,N_10200);
and U10614 (N_10614,N_10047,N_10000);
and U10615 (N_10615,N_10412,N_10050);
or U10616 (N_10616,N_10225,N_10001);
xnor U10617 (N_10617,N_10021,N_10055);
nand U10618 (N_10618,N_10405,N_10189);
and U10619 (N_10619,N_10457,N_10322);
nor U10620 (N_10620,N_10435,N_10210);
and U10621 (N_10621,N_10473,N_10138);
or U10622 (N_10622,N_10403,N_10213);
and U10623 (N_10623,N_10157,N_10301);
and U10624 (N_10624,N_10475,N_10237);
and U10625 (N_10625,N_10392,N_10187);
and U10626 (N_10626,N_10024,N_10235);
xnor U10627 (N_10627,N_10286,N_10144);
and U10628 (N_10628,N_10071,N_10193);
nand U10629 (N_10629,N_10299,N_10186);
and U10630 (N_10630,N_10044,N_10430);
and U10631 (N_10631,N_10029,N_10495);
xor U10632 (N_10632,N_10108,N_10078);
and U10633 (N_10633,N_10206,N_10004);
nand U10634 (N_10634,N_10267,N_10003);
nor U10635 (N_10635,N_10088,N_10049);
and U10636 (N_10636,N_10254,N_10058);
and U10637 (N_10637,N_10422,N_10035);
xnor U10638 (N_10638,N_10334,N_10463);
or U10639 (N_10639,N_10379,N_10153);
and U10640 (N_10640,N_10161,N_10342);
xor U10641 (N_10641,N_10081,N_10121);
nand U10642 (N_10642,N_10429,N_10106);
or U10643 (N_10643,N_10434,N_10333);
nand U10644 (N_10644,N_10360,N_10290);
nor U10645 (N_10645,N_10268,N_10386);
nor U10646 (N_10646,N_10327,N_10375);
and U10647 (N_10647,N_10137,N_10340);
xnor U10648 (N_10648,N_10466,N_10381);
and U10649 (N_10649,N_10262,N_10241);
or U10650 (N_10650,N_10184,N_10086);
xor U10651 (N_10651,N_10174,N_10018);
nor U10652 (N_10652,N_10211,N_10079);
and U10653 (N_10653,N_10220,N_10471);
or U10654 (N_10654,N_10355,N_10320);
and U10655 (N_10655,N_10217,N_10277);
nand U10656 (N_10656,N_10329,N_10196);
nor U10657 (N_10657,N_10383,N_10291);
nand U10658 (N_10658,N_10264,N_10275);
nand U10659 (N_10659,N_10387,N_10091);
and U10660 (N_10660,N_10069,N_10315);
and U10661 (N_10661,N_10113,N_10382);
and U10662 (N_10662,N_10062,N_10343);
or U10663 (N_10663,N_10249,N_10168);
nor U10664 (N_10664,N_10499,N_10353);
nand U10665 (N_10665,N_10056,N_10335);
and U10666 (N_10666,N_10402,N_10100);
xnor U10667 (N_10667,N_10278,N_10293);
xor U10668 (N_10668,N_10110,N_10272);
nand U10669 (N_10669,N_10075,N_10158);
nor U10670 (N_10670,N_10488,N_10063);
nand U10671 (N_10671,N_10094,N_10165);
xnor U10672 (N_10672,N_10178,N_10413);
nand U10673 (N_10673,N_10234,N_10314);
or U10674 (N_10674,N_10297,N_10415);
or U10675 (N_10675,N_10284,N_10470);
xnor U10676 (N_10676,N_10458,N_10032);
nor U10677 (N_10677,N_10439,N_10096);
nor U10678 (N_10678,N_10498,N_10159);
xnor U10679 (N_10679,N_10045,N_10060);
nor U10680 (N_10680,N_10019,N_10358);
xor U10681 (N_10681,N_10417,N_10147);
and U10682 (N_10682,N_10239,N_10080);
xor U10683 (N_10683,N_10316,N_10337);
nand U10684 (N_10684,N_10232,N_10409);
nor U10685 (N_10685,N_10476,N_10025);
or U10686 (N_10686,N_10076,N_10266);
xor U10687 (N_10687,N_10185,N_10145);
nor U10688 (N_10688,N_10380,N_10300);
nand U10689 (N_10689,N_10172,N_10243);
xor U10690 (N_10690,N_10256,N_10026);
xnor U10691 (N_10691,N_10228,N_10325);
nand U10692 (N_10692,N_10008,N_10253);
nor U10693 (N_10693,N_10344,N_10231);
nand U10694 (N_10694,N_10497,N_10133);
and U10695 (N_10695,N_10481,N_10207);
and U10696 (N_10696,N_10270,N_10150);
xor U10697 (N_10697,N_10326,N_10465);
xor U10698 (N_10698,N_10180,N_10389);
or U10699 (N_10699,N_10263,N_10477);
or U10700 (N_10700,N_10280,N_10433);
and U10701 (N_10701,N_10313,N_10404);
nor U10702 (N_10702,N_10484,N_10126);
nand U10703 (N_10703,N_10183,N_10377);
and U10704 (N_10704,N_10248,N_10095);
xor U10705 (N_10705,N_10357,N_10105);
xor U10706 (N_10706,N_10321,N_10203);
xnor U10707 (N_10707,N_10485,N_10289);
and U10708 (N_10708,N_10245,N_10369);
or U10709 (N_10709,N_10283,N_10310);
xnor U10710 (N_10710,N_10271,N_10216);
xnor U10711 (N_10711,N_10491,N_10449);
xnor U10712 (N_10712,N_10191,N_10419);
xor U10713 (N_10713,N_10030,N_10002);
or U10714 (N_10714,N_10292,N_10204);
xnor U10715 (N_10715,N_10296,N_10394);
and U10716 (N_10716,N_10012,N_10420);
nand U10717 (N_10717,N_10400,N_10352);
nor U10718 (N_10718,N_10202,N_10303);
and U10719 (N_10719,N_10192,N_10205);
nand U10720 (N_10720,N_10141,N_10082);
nor U10721 (N_10721,N_10155,N_10057);
and U10722 (N_10722,N_10378,N_10462);
or U10723 (N_10723,N_10149,N_10089);
nor U10724 (N_10724,N_10347,N_10474);
or U10725 (N_10725,N_10410,N_10318);
nor U10726 (N_10726,N_10036,N_10236);
or U10727 (N_10727,N_10223,N_10356);
xor U10728 (N_10728,N_10372,N_10040);
or U10729 (N_10729,N_10097,N_10309);
nor U10730 (N_10730,N_10444,N_10070);
or U10731 (N_10731,N_10421,N_10332);
and U10732 (N_10732,N_10304,N_10407);
xnor U10733 (N_10733,N_10302,N_10401);
nor U10734 (N_10734,N_10418,N_10209);
nand U10735 (N_10735,N_10146,N_10247);
or U10736 (N_10736,N_10282,N_10464);
nand U10737 (N_10737,N_10448,N_10103);
nor U10738 (N_10738,N_10424,N_10102);
xor U10739 (N_10739,N_10454,N_10115);
xor U10740 (N_10740,N_10317,N_10390);
nand U10741 (N_10741,N_10359,N_10349);
nor U10742 (N_10742,N_10017,N_10460);
or U10743 (N_10743,N_10064,N_10305);
nor U10744 (N_10744,N_10034,N_10135);
nand U10745 (N_10745,N_10396,N_10391);
or U10746 (N_10746,N_10074,N_10319);
nand U10747 (N_10747,N_10023,N_10273);
xnor U10748 (N_10748,N_10276,N_10048);
or U10749 (N_10749,N_10009,N_10362);
xor U10750 (N_10750,N_10471,N_10273);
and U10751 (N_10751,N_10438,N_10060);
xnor U10752 (N_10752,N_10475,N_10096);
and U10753 (N_10753,N_10461,N_10091);
nand U10754 (N_10754,N_10128,N_10152);
or U10755 (N_10755,N_10000,N_10185);
nand U10756 (N_10756,N_10272,N_10273);
nor U10757 (N_10757,N_10049,N_10283);
and U10758 (N_10758,N_10013,N_10069);
nand U10759 (N_10759,N_10012,N_10110);
or U10760 (N_10760,N_10159,N_10018);
nand U10761 (N_10761,N_10315,N_10235);
and U10762 (N_10762,N_10230,N_10221);
and U10763 (N_10763,N_10367,N_10480);
nor U10764 (N_10764,N_10278,N_10273);
xor U10765 (N_10765,N_10102,N_10459);
xor U10766 (N_10766,N_10323,N_10213);
and U10767 (N_10767,N_10105,N_10139);
and U10768 (N_10768,N_10107,N_10482);
or U10769 (N_10769,N_10297,N_10420);
nand U10770 (N_10770,N_10047,N_10174);
and U10771 (N_10771,N_10206,N_10005);
and U10772 (N_10772,N_10042,N_10280);
xor U10773 (N_10773,N_10226,N_10157);
or U10774 (N_10774,N_10385,N_10391);
xnor U10775 (N_10775,N_10242,N_10113);
or U10776 (N_10776,N_10373,N_10458);
nor U10777 (N_10777,N_10225,N_10407);
and U10778 (N_10778,N_10013,N_10094);
or U10779 (N_10779,N_10354,N_10445);
nand U10780 (N_10780,N_10138,N_10164);
nor U10781 (N_10781,N_10116,N_10409);
xnor U10782 (N_10782,N_10460,N_10281);
nor U10783 (N_10783,N_10290,N_10226);
or U10784 (N_10784,N_10195,N_10211);
nand U10785 (N_10785,N_10462,N_10042);
xor U10786 (N_10786,N_10476,N_10320);
or U10787 (N_10787,N_10106,N_10186);
nand U10788 (N_10788,N_10287,N_10446);
or U10789 (N_10789,N_10024,N_10082);
nor U10790 (N_10790,N_10025,N_10405);
xnor U10791 (N_10791,N_10233,N_10059);
nor U10792 (N_10792,N_10140,N_10489);
xnor U10793 (N_10793,N_10065,N_10067);
nand U10794 (N_10794,N_10497,N_10424);
xnor U10795 (N_10795,N_10377,N_10018);
nor U10796 (N_10796,N_10437,N_10148);
nor U10797 (N_10797,N_10078,N_10289);
nor U10798 (N_10798,N_10163,N_10335);
or U10799 (N_10799,N_10083,N_10388);
nand U10800 (N_10800,N_10432,N_10282);
and U10801 (N_10801,N_10052,N_10187);
nor U10802 (N_10802,N_10069,N_10264);
nor U10803 (N_10803,N_10359,N_10301);
nand U10804 (N_10804,N_10391,N_10191);
nand U10805 (N_10805,N_10418,N_10222);
xor U10806 (N_10806,N_10198,N_10338);
xor U10807 (N_10807,N_10244,N_10195);
nor U10808 (N_10808,N_10329,N_10477);
xor U10809 (N_10809,N_10223,N_10040);
or U10810 (N_10810,N_10174,N_10499);
xnor U10811 (N_10811,N_10012,N_10089);
nand U10812 (N_10812,N_10037,N_10090);
and U10813 (N_10813,N_10089,N_10248);
nand U10814 (N_10814,N_10215,N_10487);
and U10815 (N_10815,N_10203,N_10140);
or U10816 (N_10816,N_10484,N_10458);
nor U10817 (N_10817,N_10264,N_10405);
xor U10818 (N_10818,N_10015,N_10362);
and U10819 (N_10819,N_10382,N_10460);
or U10820 (N_10820,N_10271,N_10066);
xnor U10821 (N_10821,N_10344,N_10020);
nand U10822 (N_10822,N_10128,N_10298);
nor U10823 (N_10823,N_10213,N_10015);
nor U10824 (N_10824,N_10442,N_10407);
nand U10825 (N_10825,N_10320,N_10077);
nand U10826 (N_10826,N_10051,N_10075);
and U10827 (N_10827,N_10227,N_10164);
and U10828 (N_10828,N_10401,N_10433);
nor U10829 (N_10829,N_10456,N_10173);
or U10830 (N_10830,N_10399,N_10367);
and U10831 (N_10831,N_10109,N_10356);
xnor U10832 (N_10832,N_10044,N_10489);
and U10833 (N_10833,N_10348,N_10391);
or U10834 (N_10834,N_10448,N_10276);
nand U10835 (N_10835,N_10455,N_10431);
nor U10836 (N_10836,N_10282,N_10039);
and U10837 (N_10837,N_10383,N_10423);
or U10838 (N_10838,N_10103,N_10353);
nor U10839 (N_10839,N_10068,N_10343);
and U10840 (N_10840,N_10016,N_10064);
xnor U10841 (N_10841,N_10123,N_10117);
nand U10842 (N_10842,N_10363,N_10319);
xor U10843 (N_10843,N_10162,N_10284);
nand U10844 (N_10844,N_10329,N_10354);
and U10845 (N_10845,N_10416,N_10345);
xnor U10846 (N_10846,N_10095,N_10098);
nor U10847 (N_10847,N_10475,N_10343);
or U10848 (N_10848,N_10270,N_10282);
or U10849 (N_10849,N_10161,N_10236);
nand U10850 (N_10850,N_10241,N_10212);
nor U10851 (N_10851,N_10265,N_10060);
xnor U10852 (N_10852,N_10444,N_10315);
and U10853 (N_10853,N_10056,N_10352);
nor U10854 (N_10854,N_10119,N_10037);
nand U10855 (N_10855,N_10248,N_10029);
or U10856 (N_10856,N_10246,N_10377);
or U10857 (N_10857,N_10470,N_10304);
nand U10858 (N_10858,N_10182,N_10311);
xor U10859 (N_10859,N_10410,N_10131);
nor U10860 (N_10860,N_10333,N_10058);
or U10861 (N_10861,N_10069,N_10021);
nor U10862 (N_10862,N_10271,N_10059);
nand U10863 (N_10863,N_10232,N_10279);
nor U10864 (N_10864,N_10461,N_10025);
nor U10865 (N_10865,N_10265,N_10236);
xnor U10866 (N_10866,N_10103,N_10376);
nor U10867 (N_10867,N_10491,N_10002);
or U10868 (N_10868,N_10192,N_10267);
and U10869 (N_10869,N_10281,N_10362);
nand U10870 (N_10870,N_10100,N_10012);
and U10871 (N_10871,N_10217,N_10220);
xor U10872 (N_10872,N_10498,N_10028);
and U10873 (N_10873,N_10412,N_10044);
xor U10874 (N_10874,N_10158,N_10168);
xnor U10875 (N_10875,N_10369,N_10155);
nor U10876 (N_10876,N_10312,N_10333);
or U10877 (N_10877,N_10432,N_10049);
or U10878 (N_10878,N_10499,N_10450);
nor U10879 (N_10879,N_10182,N_10468);
nor U10880 (N_10880,N_10473,N_10257);
xnor U10881 (N_10881,N_10491,N_10028);
and U10882 (N_10882,N_10146,N_10166);
nand U10883 (N_10883,N_10054,N_10409);
and U10884 (N_10884,N_10356,N_10473);
and U10885 (N_10885,N_10333,N_10401);
xnor U10886 (N_10886,N_10332,N_10261);
xor U10887 (N_10887,N_10425,N_10131);
nand U10888 (N_10888,N_10239,N_10232);
or U10889 (N_10889,N_10320,N_10303);
or U10890 (N_10890,N_10092,N_10159);
nand U10891 (N_10891,N_10287,N_10347);
nor U10892 (N_10892,N_10427,N_10006);
xnor U10893 (N_10893,N_10241,N_10143);
or U10894 (N_10894,N_10287,N_10005);
nor U10895 (N_10895,N_10069,N_10397);
nor U10896 (N_10896,N_10317,N_10418);
nand U10897 (N_10897,N_10138,N_10008);
nand U10898 (N_10898,N_10398,N_10219);
or U10899 (N_10899,N_10348,N_10120);
nand U10900 (N_10900,N_10368,N_10142);
and U10901 (N_10901,N_10000,N_10305);
or U10902 (N_10902,N_10044,N_10212);
nor U10903 (N_10903,N_10054,N_10225);
or U10904 (N_10904,N_10447,N_10201);
and U10905 (N_10905,N_10063,N_10198);
xnor U10906 (N_10906,N_10442,N_10355);
and U10907 (N_10907,N_10040,N_10455);
and U10908 (N_10908,N_10372,N_10272);
xnor U10909 (N_10909,N_10088,N_10445);
and U10910 (N_10910,N_10330,N_10382);
nor U10911 (N_10911,N_10223,N_10259);
nor U10912 (N_10912,N_10462,N_10344);
or U10913 (N_10913,N_10455,N_10427);
nor U10914 (N_10914,N_10121,N_10045);
nor U10915 (N_10915,N_10310,N_10499);
or U10916 (N_10916,N_10081,N_10405);
nor U10917 (N_10917,N_10412,N_10140);
nor U10918 (N_10918,N_10123,N_10091);
and U10919 (N_10919,N_10162,N_10270);
xnor U10920 (N_10920,N_10478,N_10471);
and U10921 (N_10921,N_10449,N_10217);
and U10922 (N_10922,N_10207,N_10272);
and U10923 (N_10923,N_10082,N_10035);
xnor U10924 (N_10924,N_10111,N_10037);
nor U10925 (N_10925,N_10458,N_10264);
nand U10926 (N_10926,N_10314,N_10030);
xor U10927 (N_10927,N_10047,N_10013);
and U10928 (N_10928,N_10319,N_10357);
and U10929 (N_10929,N_10469,N_10266);
nor U10930 (N_10930,N_10018,N_10375);
or U10931 (N_10931,N_10431,N_10340);
nand U10932 (N_10932,N_10401,N_10321);
xor U10933 (N_10933,N_10222,N_10496);
or U10934 (N_10934,N_10070,N_10476);
nor U10935 (N_10935,N_10449,N_10444);
nor U10936 (N_10936,N_10321,N_10482);
nand U10937 (N_10937,N_10203,N_10256);
nor U10938 (N_10938,N_10341,N_10466);
and U10939 (N_10939,N_10095,N_10394);
nor U10940 (N_10940,N_10164,N_10342);
nand U10941 (N_10941,N_10258,N_10383);
xnor U10942 (N_10942,N_10337,N_10023);
and U10943 (N_10943,N_10424,N_10189);
nand U10944 (N_10944,N_10420,N_10344);
nand U10945 (N_10945,N_10032,N_10347);
nand U10946 (N_10946,N_10107,N_10086);
nor U10947 (N_10947,N_10234,N_10036);
xnor U10948 (N_10948,N_10467,N_10056);
or U10949 (N_10949,N_10174,N_10028);
nand U10950 (N_10950,N_10316,N_10490);
and U10951 (N_10951,N_10268,N_10365);
or U10952 (N_10952,N_10487,N_10074);
and U10953 (N_10953,N_10048,N_10245);
and U10954 (N_10954,N_10351,N_10418);
xor U10955 (N_10955,N_10445,N_10052);
and U10956 (N_10956,N_10100,N_10010);
nand U10957 (N_10957,N_10172,N_10222);
or U10958 (N_10958,N_10182,N_10433);
nor U10959 (N_10959,N_10054,N_10126);
nand U10960 (N_10960,N_10187,N_10298);
or U10961 (N_10961,N_10382,N_10010);
nor U10962 (N_10962,N_10168,N_10233);
nor U10963 (N_10963,N_10248,N_10497);
nor U10964 (N_10964,N_10430,N_10328);
and U10965 (N_10965,N_10401,N_10199);
nand U10966 (N_10966,N_10163,N_10275);
nor U10967 (N_10967,N_10316,N_10231);
nor U10968 (N_10968,N_10050,N_10465);
nand U10969 (N_10969,N_10179,N_10310);
and U10970 (N_10970,N_10497,N_10219);
xnor U10971 (N_10971,N_10371,N_10268);
or U10972 (N_10972,N_10435,N_10407);
nand U10973 (N_10973,N_10084,N_10400);
nor U10974 (N_10974,N_10203,N_10124);
and U10975 (N_10975,N_10070,N_10088);
and U10976 (N_10976,N_10281,N_10114);
and U10977 (N_10977,N_10171,N_10441);
nor U10978 (N_10978,N_10470,N_10412);
xor U10979 (N_10979,N_10378,N_10143);
xnor U10980 (N_10980,N_10417,N_10351);
and U10981 (N_10981,N_10048,N_10024);
xor U10982 (N_10982,N_10229,N_10311);
or U10983 (N_10983,N_10283,N_10469);
xnor U10984 (N_10984,N_10075,N_10282);
and U10985 (N_10985,N_10495,N_10030);
xnor U10986 (N_10986,N_10002,N_10379);
xor U10987 (N_10987,N_10295,N_10207);
nor U10988 (N_10988,N_10425,N_10112);
xor U10989 (N_10989,N_10159,N_10360);
or U10990 (N_10990,N_10405,N_10486);
or U10991 (N_10991,N_10301,N_10138);
or U10992 (N_10992,N_10382,N_10349);
nor U10993 (N_10993,N_10312,N_10400);
xnor U10994 (N_10994,N_10066,N_10281);
or U10995 (N_10995,N_10271,N_10085);
nor U10996 (N_10996,N_10418,N_10402);
nand U10997 (N_10997,N_10010,N_10245);
nor U10998 (N_10998,N_10426,N_10429);
and U10999 (N_10999,N_10374,N_10221);
and U11000 (N_11000,N_10850,N_10604);
nor U11001 (N_11001,N_10605,N_10825);
xor U11002 (N_11002,N_10637,N_10808);
or U11003 (N_11003,N_10983,N_10698);
nor U11004 (N_11004,N_10908,N_10663);
xnor U11005 (N_11005,N_10690,N_10627);
or U11006 (N_11006,N_10615,N_10590);
nor U11007 (N_11007,N_10578,N_10549);
or U11008 (N_11008,N_10992,N_10841);
nor U11009 (N_11009,N_10952,N_10626);
nand U11010 (N_11010,N_10839,N_10993);
or U11011 (N_11011,N_10638,N_10702);
and U11012 (N_11012,N_10595,N_10719);
or U11013 (N_11013,N_10946,N_10576);
or U11014 (N_11014,N_10716,N_10508);
xnor U11015 (N_11015,N_10704,N_10887);
or U11016 (N_11016,N_10697,N_10869);
nand U11017 (N_11017,N_10512,N_10914);
and U11018 (N_11018,N_10905,N_10658);
or U11019 (N_11019,N_10571,N_10525);
xnor U11020 (N_11020,N_10938,N_10912);
or U11021 (N_11021,N_10827,N_10821);
nand U11022 (N_11022,N_10685,N_10501);
nor U11023 (N_11023,N_10655,N_10788);
nand U11024 (N_11024,N_10923,N_10594);
nor U11025 (N_11025,N_10832,N_10990);
xnor U11026 (N_11026,N_10812,N_10647);
xor U11027 (N_11027,N_10889,N_10561);
and U11028 (N_11028,N_10509,N_10886);
and U11029 (N_11029,N_10642,N_10566);
and U11030 (N_11030,N_10855,N_10673);
and U11031 (N_11031,N_10533,N_10511);
or U11032 (N_11032,N_10980,N_10510);
xnor U11033 (N_11033,N_10819,N_10744);
xnor U11034 (N_11034,N_10795,N_10932);
nor U11035 (N_11035,N_10653,N_10896);
nand U11036 (N_11036,N_10739,N_10756);
nand U11037 (N_11037,N_10589,N_10957);
xor U11038 (N_11038,N_10676,N_10570);
and U11039 (N_11039,N_10974,N_10966);
xor U11040 (N_11040,N_10767,N_10822);
or U11041 (N_11041,N_10635,N_10999);
and U11042 (N_11042,N_10505,N_10797);
or U11043 (N_11043,N_10534,N_10579);
or U11044 (N_11044,N_10623,N_10991);
nor U11045 (N_11045,N_10577,N_10970);
nor U11046 (N_11046,N_10568,N_10921);
and U11047 (N_11047,N_10679,N_10728);
and U11048 (N_11048,N_10644,N_10718);
nand U11049 (N_11049,N_10554,N_10592);
or U11050 (N_11050,N_10665,N_10749);
or U11051 (N_11051,N_10763,N_10979);
or U11052 (N_11052,N_10768,N_10774);
and U11053 (N_11053,N_10560,N_10972);
nor U11054 (N_11054,N_10870,N_10654);
and U11055 (N_11055,N_10927,N_10516);
nand U11056 (N_11056,N_10751,N_10610);
and U11057 (N_11057,N_10607,N_10503);
nand U11058 (N_11058,N_10624,N_10546);
or U11059 (N_11059,N_10646,N_10695);
xnor U11060 (N_11060,N_10700,N_10956);
xor U11061 (N_11061,N_10694,N_10670);
or U11062 (N_11062,N_10681,N_10733);
or U11063 (N_11063,N_10890,N_10666);
and U11064 (N_11064,N_10944,N_10917);
xor U11065 (N_11065,N_10844,N_10929);
nor U11066 (N_11066,N_10961,N_10996);
xor U11067 (N_11067,N_10981,N_10523);
nand U11068 (N_11068,N_10831,N_10772);
nand U11069 (N_11069,N_10630,N_10893);
nor U11070 (N_11070,N_10785,N_10888);
and U11071 (N_11071,N_10514,N_10902);
nand U11072 (N_11072,N_10965,N_10969);
and U11073 (N_11073,N_10786,N_10810);
nand U11074 (N_11074,N_10779,N_10684);
nand U11075 (N_11075,N_10667,N_10959);
xnor U11076 (N_11076,N_10731,N_10924);
or U11077 (N_11077,N_10910,N_10793);
and U11078 (N_11078,N_10746,N_10918);
nor U11079 (N_11079,N_10747,N_10677);
nand U11080 (N_11080,N_10936,N_10757);
nor U11081 (N_11081,N_10836,N_10903);
nand U11082 (N_11082,N_10608,N_10633);
nor U11083 (N_11083,N_10943,N_10773);
and U11084 (N_11084,N_10552,N_10602);
or U11085 (N_11085,N_10729,N_10529);
nand U11086 (N_11086,N_10569,N_10527);
nand U11087 (N_11087,N_10748,N_10564);
or U11088 (N_11088,N_10581,N_10616);
and U11089 (N_11089,N_10851,N_10906);
xor U11090 (N_11090,N_10815,N_10706);
xnor U11091 (N_11091,N_10937,N_10875);
and U11092 (N_11092,N_10975,N_10674);
or U11093 (N_11093,N_10898,N_10593);
xor U11094 (N_11094,N_10899,N_10531);
xnor U11095 (N_11095,N_10804,N_10600);
xor U11096 (N_11096,N_10897,N_10761);
nand U11097 (N_11097,N_10829,N_10881);
nand U11098 (N_11098,N_10708,N_10539);
and U11099 (N_11099,N_10545,N_10843);
nor U11100 (N_11100,N_10864,N_10606);
xnor U11101 (N_11101,N_10920,N_10659);
xnor U11102 (N_11102,N_10771,N_10978);
nor U11103 (N_11103,N_10973,N_10504);
xor U11104 (N_11104,N_10775,N_10584);
nor U11105 (N_11105,N_10692,N_10620);
or U11106 (N_11106,N_10682,N_10721);
or U11107 (N_11107,N_10892,N_10651);
nand U11108 (N_11108,N_10555,N_10652);
xor U11109 (N_11109,N_10805,N_10934);
and U11110 (N_11110,N_10942,N_10876);
xor U11111 (N_11111,N_10878,N_10553);
or U11112 (N_11112,N_10699,N_10567);
and U11113 (N_11113,N_10913,N_10930);
xor U11114 (N_11114,N_10813,N_10950);
nor U11115 (N_11115,N_10524,N_10781);
nor U11116 (N_11116,N_10826,N_10925);
xnor U11117 (N_11117,N_10986,N_10955);
nor U11118 (N_11118,N_10587,N_10544);
nor U11119 (N_11119,N_10960,N_10834);
nand U11120 (N_11120,N_10634,N_10645);
nand U11121 (N_11121,N_10532,N_10740);
or U11122 (N_11122,N_10828,N_10854);
and U11123 (N_11123,N_10783,N_10872);
nor U11124 (N_11124,N_10933,N_10530);
xnor U11125 (N_11125,N_10853,N_10540);
nand U11126 (N_11126,N_10643,N_10588);
or U11127 (N_11127,N_10947,N_10777);
xor U11128 (N_11128,N_10657,N_10660);
nand U11129 (N_11129,N_10689,N_10664);
nor U11130 (N_11130,N_10625,N_10585);
nand U11131 (N_11131,N_10752,N_10948);
or U11132 (N_11132,N_10565,N_10711);
and U11133 (N_11133,N_10572,N_10526);
nand U11134 (N_11134,N_10997,N_10737);
xnor U11135 (N_11135,N_10556,N_10537);
or U11136 (N_11136,N_10732,N_10949);
or U11137 (N_11137,N_10557,N_10707);
xnor U11138 (N_11138,N_10867,N_10693);
nand U11139 (N_11139,N_10856,N_10631);
nor U11140 (N_11140,N_10596,N_10866);
nand U11141 (N_11141,N_10720,N_10662);
nand U11142 (N_11142,N_10860,N_10803);
xnor U11143 (N_11143,N_10703,N_10521);
and U11144 (N_11144,N_10686,N_10519);
and U11145 (N_11145,N_10784,N_10649);
nor U11146 (N_11146,N_10926,N_10935);
nor U11147 (N_11147,N_10842,N_10678);
nand U11148 (N_11148,N_10621,N_10586);
or U11149 (N_11149,N_10789,N_10538);
and U11150 (N_11150,N_10722,N_10614);
xnor U11151 (N_11151,N_10675,N_10687);
and U11152 (N_11152,N_10904,N_10745);
nand U11153 (N_11153,N_10940,N_10998);
nor U11154 (N_11154,N_10573,N_10563);
and U11155 (N_11155,N_10518,N_10591);
and U11156 (N_11156,N_10814,N_10724);
and U11157 (N_11157,N_10922,N_10536);
and U11158 (N_11158,N_10984,N_10951);
or U11159 (N_11159,N_10770,N_10816);
or U11160 (N_11160,N_10612,N_10717);
and U11161 (N_11161,N_10862,N_10507);
xnor U11162 (N_11162,N_10726,N_10683);
nand U11163 (N_11163,N_10730,N_10953);
xnor U11164 (N_11164,N_10599,N_10696);
or U11165 (N_11165,N_10502,N_10758);
nand U11166 (N_11166,N_10900,N_10597);
nor U11167 (N_11167,N_10710,N_10513);
nand U11168 (N_11168,N_10865,N_10840);
or U11169 (N_11169,N_10661,N_10846);
and U11170 (N_11170,N_10598,N_10916);
and U11171 (N_11171,N_10559,N_10963);
nor U11172 (N_11172,N_10764,N_10945);
nand U11173 (N_11173,N_10601,N_10871);
nand U11174 (N_11174,N_10941,N_10542);
nand U11175 (N_11175,N_10891,N_10712);
or U11176 (N_11176,N_10837,N_10835);
nand U11177 (N_11177,N_10909,N_10823);
or U11178 (N_11178,N_10550,N_10801);
nand U11179 (N_11179,N_10641,N_10769);
or U11180 (N_11180,N_10792,N_10873);
nor U11181 (N_11181,N_10582,N_10632);
nor U11182 (N_11182,N_10976,N_10848);
xnor U11183 (N_11183,N_10939,N_10882);
nor U11184 (N_11184,N_10762,N_10743);
nor U11185 (N_11185,N_10820,N_10800);
xor U11186 (N_11186,N_10811,N_10520);
nand U11187 (N_11187,N_10613,N_10715);
nor U11188 (N_11188,N_10964,N_10562);
or U11189 (N_11189,N_10734,N_10691);
xnor U11190 (N_11190,N_10622,N_10575);
nor U11191 (N_11191,N_10830,N_10884);
xor U11192 (N_11192,N_10852,N_10628);
and U11193 (N_11193,N_10859,N_10522);
nand U11194 (N_11194,N_10995,N_10736);
nand U11195 (N_11195,N_10790,N_10799);
and U11196 (N_11196,N_10766,N_10506);
or U11197 (N_11197,N_10688,N_10988);
and U11198 (N_11198,N_10583,N_10535);
nor U11199 (N_11199,N_10931,N_10547);
nand U11200 (N_11200,N_10639,N_10609);
and U11201 (N_11201,N_10750,N_10709);
nand U11202 (N_11202,N_10911,N_10760);
nand U11203 (N_11203,N_10879,N_10741);
or U11204 (N_11204,N_10919,N_10725);
nor U11205 (N_11205,N_10794,N_10928);
and U11206 (N_11206,N_10517,N_10705);
nand U11207 (N_11207,N_10874,N_10500);
nand U11208 (N_11208,N_10742,N_10754);
and U11209 (N_11209,N_10958,N_10668);
nor U11210 (N_11210,N_10967,N_10541);
xor U11211 (N_11211,N_10603,N_10735);
nand U11212 (N_11212,N_10987,N_10543);
nand U11213 (N_11213,N_10672,N_10907);
and U11214 (N_11214,N_10738,N_10640);
or U11215 (N_11215,N_10656,N_10791);
xnor U11216 (N_11216,N_10807,N_10894);
or U11217 (N_11217,N_10787,N_10713);
and U11218 (N_11218,N_10982,N_10977);
xnor U11219 (N_11219,N_10776,N_10617);
xnor U11220 (N_11220,N_10985,N_10817);
nand U11221 (N_11221,N_10818,N_10574);
nand U11222 (N_11222,N_10782,N_10824);
nor U11223 (N_11223,N_10753,N_10551);
nor U11224 (N_11224,N_10618,N_10755);
xnor U11225 (N_11225,N_10838,N_10648);
and U11226 (N_11226,N_10968,N_10802);
or U11227 (N_11227,N_10806,N_10994);
nand U11228 (N_11228,N_10847,N_10680);
xor U11229 (N_11229,N_10971,N_10558);
and U11230 (N_11230,N_10989,N_10798);
xor U11231 (N_11231,N_10650,N_10528);
nor U11232 (N_11232,N_10877,N_10669);
nand U11233 (N_11233,N_10962,N_10895);
nor U11234 (N_11234,N_10759,N_10883);
and U11235 (N_11235,N_10901,N_10796);
and U11236 (N_11236,N_10857,N_10849);
and U11237 (N_11237,N_10861,N_10845);
nor U11238 (N_11238,N_10780,N_10714);
xor U11239 (N_11239,N_10858,N_10629);
and U11240 (N_11240,N_10611,N_10701);
nor U11241 (N_11241,N_10671,N_10619);
and U11242 (N_11242,N_10863,N_10636);
xnor U11243 (N_11243,N_10727,N_10809);
or U11244 (N_11244,N_10833,N_10880);
and U11245 (N_11245,N_10868,N_10548);
xor U11246 (N_11246,N_10885,N_10723);
and U11247 (N_11247,N_10765,N_10778);
xor U11248 (N_11248,N_10915,N_10954);
or U11249 (N_11249,N_10580,N_10515);
nor U11250 (N_11250,N_10794,N_10779);
nor U11251 (N_11251,N_10667,N_10714);
and U11252 (N_11252,N_10875,N_10736);
nor U11253 (N_11253,N_10826,N_10702);
and U11254 (N_11254,N_10581,N_10637);
nand U11255 (N_11255,N_10623,N_10767);
nor U11256 (N_11256,N_10872,N_10883);
nor U11257 (N_11257,N_10975,N_10689);
and U11258 (N_11258,N_10516,N_10887);
and U11259 (N_11259,N_10707,N_10641);
nand U11260 (N_11260,N_10648,N_10583);
nand U11261 (N_11261,N_10543,N_10643);
nor U11262 (N_11262,N_10730,N_10709);
and U11263 (N_11263,N_10891,N_10571);
nor U11264 (N_11264,N_10938,N_10804);
or U11265 (N_11265,N_10643,N_10841);
or U11266 (N_11266,N_10983,N_10680);
xnor U11267 (N_11267,N_10595,N_10682);
and U11268 (N_11268,N_10679,N_10741);
xor U11269 (N_11269,N_10823,N_10581);
nor U11270 (N_11270,N_10698,N_10965);
xnor U11271 (N_11271,N_10992,N_10505);
nor U11272 (N_11272,N_10750,N_10697);
and U11273 (N_11273,N_10805,N_10964);
xnor U11274 (N_11274,N_10900,N_10544);
nor U11275 (N_11275,N_10694,N_10709);
nand U11276 (N_11276,N_10577,N_10706);
nor U11277 (N_11277,N_10809,N_10682);
nand U11278 (N_11278,N_10513,N_10676);
nor U11279 (N_11279,N_10947,N_10774);
or U11280 (N_11280,N_10857,N_10647);
nand U11281 (N_11281,N_10658,N_10985);
nand U11282 (N_11282,N_10782,N_10559);
nand U11283 (N_11283,N_10565,N_10834);
xor U11284 (N_11284,N_10997,N_10532);
nor U11285 (N_11285,N_10743,N_10649);
xnor U11286 (N_11286,N_10881,N_10574);
nor U11287 (N_11287,N_10642,N_10926);
xor U11288 (N_11288,N_10756,N_10880);
nand U11289 (N_11289,N_10537,N_10592);
nor U11290 (N_11290,N_10783,N_10596);
nand U11291 (N_11291,N_10598,N_10641);
or U11292 (N_11292,N_10841,N_10858);
or U11293 (N_11293,N_10964,N_10857);
xnor U11294 (N_11294,N_10968,N_10931);
xnor U11295 (N_11295,N_10690,N_10997);
and U11296 (N_11296,N_10713,N_10782);
xnor U11297 (N_11297,N_10762,N_10732);
and U11298 (N_11298,N_10890,N_10788);
or U11299 (N_11299,N_10578,N_10707);
or U11300 (N_11300,N_10914,N_10969);
xor U11301 (N_11301,N_10653,N_10711);
xnor U11302 (N_11302,N_10658,N_10556);
nand U11303 (N_11303,N_10704,N_10813);
nand U11304 (N_11304,N_10627,N_10941);
or U11305 (N_11305,N_10954,N_10722);
and U11306 (N_11306,N_10790,N_10764);
nand U11307 (N_11307,N_10683,N_10634);
nand U11308 (N_11308,N_10942,N_10651);
nand U11309 (N_11309,N_10567,N_10513);
and U11310 (N_11310,N_10748,N_10509);
nand U11311 (N_11311,N_10651,N_10716);
nor U11312 (N_11312,N_10781,N_10665);
or U11313 (N_11313,N_10684,N_10801);
nor U11314 (N_11314,N_10939,N_10658);
xor U11315 (N_11315,N_10986,N_10609);
nand U11316 (N_11316,N_10649,N_10514);
and U11317 (N_11317,N_10710,N_10886);
or U11318 (N_11318,N_10557,N_10981);
nand U11319 (N_11319,N_10638,N_10544);
xnor U11320 (N_11320,N_10833,N_10750);
or U11321 (N_11321,N_10597,N_10729);
and U11322 (N_11322,N_10840,N_10838);
xnor U11323 (N_11323,N_10993,N_10511);
nand U11324 (N_11324,N_10669,N_10522);
or U11325 (N_11325,N_10725,N_10748);
or U11326 (N_11326,N_10803,N_10555);
xnor U11327 (N_11327,N_10717,N_10943);
and U11328 (N_11328,N_10504,N_10594);
and U11329 (N_11329,N_10764,N_10872);
and U11330 (N_11330,N_10938,N_10931);
nor U11331 (N_11331,N_10617,N_10562);
nor U11332 (N_11332,N_10745,N_10942);
and U11333 (N_11333,N_10529,N_10525);
or U11334 (N_11334,N_10638,N_10901);
xnor U11335 (N_11335,N_10958,N_10517);
nor U11336 (N_11336,N_10652,N_10847);
and U11337 (N_11337,N_10658,N_10765);
xor U11338 (N_11338,N_10553,N_10532);
or U11339 (N_11339,N_10519,N_10720);
nor U11340 (N_11340,N_10524,N_10589);
xnor U11341 (N_11341,N_10853,N_10717);
nand U11342 (N_11342,N_10835,N_10897);
xnor U11343 (N_11343,N_10984,N_10638);
and U11344 (N_11344,N_10640,N_10687);
and U11345 (N_11345,N_10947,N_10948);
and U11346 (N_11346,N_10853,N_10930);
xnor U11347 (N_11347,N_10966,N_10550);
nor U11348 (N_11348,N_10731,N_10501);
or U11349 (N_11349,N_10506,N_10518);
or U11350 (N_11350,N_10866,N_10787);
nand U11351 (N_11351,N_10626,N_10581);
and U11352 (N_11352,N_10889,N_10873);
and U11353 (N_11353,N_10654,N_10701);
and U11354 (N_11354,N_10927,N_10693);
and U11355 (N_11355,N_10578,N_10630);
xor U11356 (N_11356,N_10692,N_10933);
or U11357 (N_11357,N_10761,N_10781);
nand U11358 (N_11358,N_10945,N_10802);
nand U11359 (N_11359,N_10650,N_10943);
and U11360 (N_11360,N_10627,N_10925);
nor U11361 (N_11361,N_10708,N_10610);
or U11362 (N_11362,N_10868,N_10521);
or U11363 (N_11363,N_10546,N_10686);
or U11364 (N_11364,N_10707,N_10735);
and U11365 (N_11365,N_10813,N_10954);
xnor U11366 (N_11366,N_10956,N_10585);
nor U11367 (N_11367,N_10930,N_10980);
and U11368 (N_11368,N_10835,N_10684);
and U11369 (N_11369,N_10864,N_10717);
and U11370 (N_11370,N_10521,N_10976);
nand U11371 (N_11371,N_10550,N_10746);
nor U11372 (N_11372,N_10839,N_10651);
and U11373 (N_11373,N_10575,N_10651);
or U11374 (N_11374,N_10789,N_10507);
nand U11375 (N_11375,N_10960,N_10852);
or U11376 (N_11376,N_10780,N_10914);
or U11377 (N_11377,N_10971,N_10722);
xor U11378 (N_11378,N_10697,N_10532);
xnor U11379 (N_11379,N_10562,N_10655);
or U11380 (N_11380,N_10598,N_10610);
nor U11381 (N_11381,N_10945,N_10670);
and U11382 (N_11382,N_10643,N_10521);
nand U11383 (N_11383,N_10630,N_10761);
and U11384 (N_11384,N_10914,N_10857);
nand U11385 (N_11385,N_10990,N_10833);
and U11386 (N_11386,N_10542,N_10855);
xnor U11387 (N_11387,N_10977,N_10657);
or U11388 (N_11388,N_10520,N_10825);
nand U11389 (N_11389,N_10583,N_10871);
and U11390 (N_11390,N_10943,N_10706);
or U11391 (N_11391,N_10841,N_10993);
nand U11392 (N_11392,N_10520,N_10961);
or U11393 (N_11393,N_10618,N_10963);
nor U11394 (N_11394,N_10553,N_10992);
xor U11395 (N_11395,N_10708,N_10822);
nand U11396 (N_11396,N_10906,N_10664);
nor U11397 (N_11397,N_10631,N_10848);
xor U11398 (N_11398,N_10742,N_10723);
xor U11399 (N_11399,N_10921,N_10543);
nor U11400 (N_11400,N_10647,N_10786);
and U11401 (N_11401,N_10512,N_10804);
nor U11402 (N_11402,N_10675,N_10868);
nand U11403 (N_11403,N_10968,N_10512);
xnor U11404 (N_11404,N_10698,N_10542);
xnor U11405 (N_11405,N_10791,N_10919);
xnor U11406 (N_11406,N_10895,N_10890);
xor U11407 (N_11407,N_10598,N_10608);
xnor U11408 (N_11408,N_10675,N_10964);
or U11409 (N_11409,N_10562,N_10620);
nand U11410 (N_11410,N_10613,N_10983);
xnor U11411 (N_11411,N_10552,N_10995);
or U11412 (N_11412,N_10970,N_10857);
xnor U11413 (N_11413,N_10919,N_10589);
nand U11414 (N_11414,N_10727,N_10747);
nor U11415 (N_11415,N_10998,N_10576);
xnor U11416 (N_11416,N_10893,N_10813);
and U11417 (N_11417,N_10506,N_10700);
nor U11418 (N_11418,N_10768,N_10798);
nor U11419 (N_11419,N_10573,N_10544);
xnor U11420 (N_11420,N_10908,N_10938);
nor U11421 (N_11421,N_10906,N_10879);
and U11422 (N_11422,N_10992,N_10701);
or U11423 (N_11423,N_10730,N_10597);
or U11424 (N_11424,N_10595,N_10696);
xnor U11425 (N_11425,N_10985,N_10808);
nor U11426 (N_11426,N_10560,N_10976);
nand U11427 (N_11427,N_10891,N_10711);
and U11428 (N_11428,N_10517,N_10942);
nor U11429 (N_11429,N_10545,N_10683);
and U11430 (N_11430,N_10685,N_10858);
nor U11431 (N_11431,N_10841,N_10718);
or U11432 (N_11432,N_10939,N_10714);
nand U11433 (N_11433,N_10570,N_10621);
or U11434 (N_11434,N_10768,N_10845);
or U11435 (N_11435,N_10884,N_10694);
and U11436 (N_11436,N_10873,N_10546);
nor U11437 (N_11437,N_10693,N_10795);
or U11438 (N_11438,N_10647,N_10973);
nor U11439 (N_11439,N_10824,N_10520);
or U11440 (N_11440,N_10614,N_10984);
or U11441 (N_11441,N_10593,N_10613);
nor U11442 (N_11442,N_10952,N_10745);
nand U11443 (N_11443,N_10506,N_10658);
or U11444 (N_11444,N_10618,N_10841);
xnor U11445 (N_11445,N_10952,N_10713);
xnor U11446 (N_11446,N_10553,N_10621);
nand U11447 (N_11447,N_10776,N_10592);
or U11448 (N_11448,N_10818,N_10901);
and U11449 (N_11449,N_10660,N_10993);
or U11450 (N_11450,N_10824,N_10565);
nand U11451 (N_11451,N_10825,N_10777);
xor U11452 (N_11452,N_10584,N_10985);
nand U11453 (N_11453,N_10778,N_10962);
or U11454 (N_11454,N_10857,N_10641);
nand U11455 (N_11455,N_10618,N_10661);
nor U11456 (N_11456,N_10575,N_10523);
nand U11457 (N_11457,N_10750,N_10721);
or U11458 (N_11458,N_10854,N_10787);
and U11459 (N_11459,N_10530,N_10911);
and U11460 (N_11460,N_10671,N_10854);
nand U11461 (N_11461,N_10985,N_10698);
nand U11462 (N_11462,N_10915,N_10732);
nand U11463 (N_11463,N_10886,N_10938);
and U11464 (N_11464,N_10603,N_10891);
and U11465 (N_11465,N_10997,N_10723);
nand U11466 (N_11466,N_10852,N_10501);
xnor U11467 (N_11467,N_10661,N_10989);
nor U11468 (N_11468,N_10692,N_10834);
and U11469 (N_11469,N_10714,N_10663);
or U11470 (N_11470,N_10856,N_10811);
nand U11471 (N_11471,N_10877,N_10739);
nand U11472 (N_11472,N_10913,N_10866);
xor U11473 (N_11473,N_10895,N_10946);
and U11474 (N_11474,N_10614,N_10783);
and U11475 (N_11475,N_10984,N_10589);
xnor U11476 (N_11476,N_10852,N_10834);
or U11477 (N_11477,N_10616,N_10672);
and U11478 (N_11478,N_10597,N_10616);
or U11479 (N_11479,N_10506,N_10939);
nor U11480 (N_11480,N_10526,N_10583);
nand U11481 (N_11481,N_10882,N_10832);
or U11482 (N_11482,N_10585,N_10829);
nor U11483 (N_11483,N_10932,N_10540);
or U11484 (N_11484,N_10578,N_10834);
nor U11485 (N_11485,N_10750,N_10635);
nand U11486 (N_11486,N_10519,N_10883);
xnor U11487 (N_11487,N_10578,N_10552);
and U11488 (N_11488,N_10529,N_10840);
and U11489 (N_11489,N_10912,N_10796);
xor U11490 (N_11490,N_10916,N_10764);
nor U11491 (N_11491,N_10735,N_10685);
nor U11492 (N_11492,N_10748,N_10795);
xnor U11493 (N_11493,N_10866,N_10529);
or U11494 (N_11494,N_10965,N_10962);
xnor U11495 (N_11495,N_10669,N_10700);
and U11496 (N_11496,N_10976,N_10924);
and U11497 (N_11497,N_10838,N_10678);
and U11498 (N_11498,N_10790,N_10618);
nand U11499 (N_11499,N_10698,N_10789);
nor U11500 (N_11500,N_11072,N_11416);
and U11501 (N_11501,N_11440,N_11215);
and U11502 (N_11502,N_11335,N_11441);
xor U11503 (N_11503,N_11467,N_11397);
nor U11504 (N_11504,N_11245,N_11007);
nand U11505 (N_11505,N_11450,N_11209);
nand U11506 (N_11506,N_11204,N_11049);
and U11507 (N_11507,N_11449,N_11357);
and U11508 (N_11508,N_11261,N_11286);
nor U11509 (N_11509,N_11491,N_11418);
or U11510 (N_11510,N_11227,N_11190);
and U11511 (N_11511,N_11135,N_11443);
nor U11512 (N_11512,N_11137,N_11050);
nor U11513 (N_11513,N_11062,N_11297);
nand U11514 (N_11514,N_11311,N_11205);
nand U11515 (N_11515,N_11216,N_11411);
or U11516 (N_11516,N_11146,N_11424);
and U11517 (N_11517,N_11325,N_11320);
and U11518 (N_11518,N_11363,N_11296);
xor U11519 (N_11519,N_11422,N_11428);
nand U11520 (N_11520,N_11122,N_11052);
nand U11521 (N_11521,N_11039,N_11488);
nand U11522 (N_11522,N_11337,N_11029);
nor U11523 (N_11523,N_11106,N_11021);
nor U11524 (N_11524,N_11228,N_11408);
and U11525 (N_11525,N_11444,N_11338);
nand U11526 (N_11526,N_11085,N_11233);
nor U11527 (N_11527,N_11268,N_11486);
nor U11528 (N_11528,N_11390,N_11217);
xnor U11529 (N_11529,N_11082,N_11153);
and U11530 (N_11530,N_11154,N_11377);
nand U11531 (N_11531,N_11068,N_11383);
or U11532 (N_11532,N_11437,N_11386);
and U11533 (N_11533,N_11108,N_11412);
xnor U11534 (N_11534,N_11170,N_11407);
and U11535 (N_11535,N_11025,N_11127);
or U11536 (N_11536,N_11103,N_11121);
xor U11537 (N_11537,N_11092,N_11178);
or U11538 (N_11538,N_11023,N_11352);
or U11539 (N_11539,N_11376,N_11175);
xor U11540 (N_11540,N_11264,N_11414);
and U11541 (N_11541,N_11493,N_11000);
or U11542 (N_11542,N_11123,N_11241);
nor U11543 (N_11543,N_11287,N_11421);
or U11544 (N_11544,N_11447,N_11285);
nand U11545 (N_11545,N_11333,N_11150);
xnor U11546 (N_11546,N_11315,N_11339);
and U11547 (N_11547,N_11476,N_11477);
xor U11548 (N_11548,N_11078,N_11400);
nand U11549 (N_11549,N_11079,N_11037);
or U11550 (N_11550,N_11246,N_11047);
xnor U11551 (N_11551,N_11382,N_11022);
nand U11552 (N_11552,N_11157,N_11188);
nand U11553 (N_11553,N_11095,N_11176);
xor U11554 (N_11554,N_11323,N_11265);
and U11555 (N_11555,N_11358,N_11445);
and U11556 (N_11556,N_11226,N_11334);
and U11557 (N_11557,N_11064,N_11163);
nor U11558 (N_11558,N_11448,N_11456);
nor U11559 (N_11559,N_11249,N_11292);
nand U11560 (N_11560,N_11279,N_11080);
and U11561 (N_11561,N_11101,N_11484);
nand U11562 (N_11562,N_11319,N_11259);
xor U11563 (N_11563,N_11015,N_11168);
nand U11564 (N_11564,N_11393,N_11403);
nand U11565 (N_11565,N_11237,N_11253);
and U11566 (N_11566,N_11071,N_11370);
nand U11567 (N_11567,N_11158,N_11183);
nand U11568 (N_11568,N_11099,N_11385);
and U11569 (N_11569,N_11165,N_11281);
nor U11570 (N_11570,N_11307,N_11374);
xor U11571 (N_11571,N_11090,N_11371);
or U11572 (N_11572,N_11434,N_11081);
xnor U11573 (N_11573,N_11141,N_11271);
nand U11574 (N_11574,N_11191,N_11343);
nor U11575 (N_11575,N_11482,N_11111);
and U11576 (N_11576,N_11304,N_11425);
nor U11577 (N_11577,N_11203,N_11086);
nand U11578 (N_11578,N_11347,N_11219);
or U11579 (N_11579,N_11032,N_11475);
or U11580 (N_11580,N_11273,N_11151);
and U11581 (N_11581,N_11497,N_11238);
and U11582 (N_11582,N_11288,N_11387);
xnor U11583 (N_11583,N_11470,N_11034);
xnor U11584 (N_11584,N_11199,N_11088);
or U11585 (N_11585,N_11011,N_11066);
nand U11586 (N_11586,N_11131,N_11433);
and U11587 (N_11587,N_11289,N_11465);
and U11588 (N_11588,N_11458,N_11362);
nand U11589 (N_11589,N_11294,N_11251);
nand U11590 (N_11590,N_11196,N_11295);
or U11591 (N_11591,N_11327,N_11051);
xor U11592 (N_11592,N_11193,N_11169);
nand U11593 (N_11593,N_11100,N_11044);
nand U11594 (N_11594,N_11405,N_11223);
and U11595 (N_11595,N_11473,N_11471);
and U11596 (N_11596,N_11208,N_11236);
nand U11597 (N_11597,N_11161,N_11275);
nand U11598 (N_11598,N_11423,N_11116);
and U11599 (N_11599,N_11128,N_11496);
nand U11600 (N_11600,N_11160,N_11406);
nor U11601 (N_11601,N_11427,N_11087);
or U11602 (N_11602,N_11211,N_11316);
nand U11603 (N_11603,N_11464,N_11457);
nor U11604 (N_11604,N_11002,N_11167);
and U11605 (N_11605,N_11305,N_11075);
xnor U11606 (N_11606,N_11389,N_11177);
nand U11607 (N_11607,N_11004,N_11166);
nor U11608 (N_11608,N_11495,N_11171);
nand U11609 (N_11609,N_11026,N_11104);
and U11610 (N_11610,N_11340,N_11189);
or U11611 (N_11611,N_11056,N_11126);
and U11612 (N_11612,N_11195,N_11481);
xnor U11613 (N_11613,N_11453,N_11270);
or U11614 (N_11614,N_11276,N_11173);
nor U11615 (N_11615,N_11256,N_11391);
nand U11616 (N_11616,N_11243,N_11113);
and U11617 (N_11617,N_11360,N_11240);
xnor U11618 (N_11618,N_11359,N_11048);
and U11619 (N_11619,N_11058,N_11059);
xnor U11620 (N_11620,N_11398,N_11489);
and U11621 (N_11621,N_11186,N_11054);
xnor U11622 (N_11622,N_11089,N_11415);
nor U11623 (N_11623,N_11419,N_11028);
nand U11624 (N_11624,N_11446,N_11006);
or U11625 (N_11625,N_11280,N_11024);
nand U11626 (N_11626,N_11417,N_11399);
nor U11627 (N_11627,N_11290,N_11365);
nand U11628 (N_11628,N_11384,N_11120);
or U11629 (N_11629,N_11388,N_11198);
and U11630 (N_11630,N_11460,N_11063);
nor U11631 (N_11631,N_11224,N_11105);
nor U11632 (N_11632,N_11067,N_11159);
nor U11633 (N_11633,N_11485,N_11083);
and U11634 (N_11634,N_11461,N_11269);
nand U11635 (N_11635,N_11060,N_11013);
or U11636 (N_11636,N_11221,N_11220);
xor U11637 (N_11637,N_11016,N_11348);
and U11638 (N_11638,N_11124,N_11452);
xnor U11639 (N_11639,N_11324,N_11330);
or U11640 (N_11640,N_11074,N_11353);
and U11641 (N_11641,N_11252,N_11213);
nand U11642 (N_11642,N_11244,N_11134);
or U11643 (N_11643,N_11107,N_11472);
xor U11644 (N_11644,N_11114,N_11490);
or U11645 (N_11645,N_11200,N_11156);
xor U11646 (N_11646,N_11118,N_11431);
xor U11647 (N_11647,N_11364,N_11369);
or U11648 (N_11648,N_11117,N_11351);
and U11649 (N_11649,N_11225,N_11030);
nand U11650 (N_11650,N_11487,N_11084);
xor U11651 (N_11651,N_11235,N_11184);
or U11652 (N_11652,N_11368,N_11152);
and U11653 (N_11653,N_11136,N_11202);
nor U11654 (N_11654,N_11313,N_11318);
nand U11655 (N_11655,N_11291,N_11144);
or U11656 (N_11656,N_11222,N_11008);
xnor U11657 (N_11657,N_11057,N_11125);
or U11658 (N_11658,N_11420,N_11040);
or U11659 (N_11659,N_11462,N_11185);
nor U11660 (N_11660,N_11454,N_11302);
nand U11661 (N_11661,N_11043,N_11306);
xor U11662 (N_11662,N_11140,N_11426);
xnor U11663 (N_11663,N_11155,N_11375);
or U11664 (N_11664,N_11206,N_11344);
and U11665 (N_11665,N_11053,N_11031);
nor U11666 (N_11666,N_11479,N_11017);
or U11667 (N_11667,N_11182,N_11257);
nor U11668 (N_11668,N_11027,N_11277);
nor U11669 (N_11669,N_11317,N_11005);
nand U11670 (N_11670,N_11001,N_11110);
xor U11671 (N_11671,N_11009,N_11480);
xor U11672 (N_11672,N_11263,N_11463);
and U11673 (N_11673,N_11468,N_11413);
or U11674 (N_11674,N_11336,N_11258);
nor U11675 (N_11675,N_11218,N_11260);
xnor U11676 (N_11676,N_11361,N_11180);
and U11677 (N_11677,N_11042,N_11442);
and U11678 (N_11678,N_11018,N_11282);
xor U11679 (N_11679,N_11139,N_11115);
nor U11680 (N_11680,N_11250,N_11142);
nor U11681 (N_11681,N_11036,N_11308);
nor U11682 (N_11682,N_11367,N_11010);
and U11683 (N_11683,N_11298,N_11109);
nor U11684 (N_11684,N_11234,N_11394);
and U11685 (N_11685,N_11300,N_11395);
nor U11686 (N_11686,N_11455,N_11093);
nor U11687 (N_11687,N_11346,N_11239);
and U11688 (N_11688,N_11194,N_11469);
xor U11689 (N_11689,N_11201,N_11247);
nor U11690 (N_11690,N_11232,N_11212);
xor U11691 (N_11691,N_11402,N_11341);
and U11692 (N_11692,N_11164,N_11309);
xor U11693 (N_11693,N_11197,N_11435);
xnor U11694 (N_11694,N_11439,N_11354);
nand U11695 (N_11695,N_11035,N_11070);
nand U11696 (N_11696,N_11148,N_11102);
and U11697 (N_11697,N_11094,N_11172);
xnor U11698 (N_11698,N_11248,N_11429);
and U11699 (N_11699,N_11392,N_11430);
nor U11700 (N_11700,N_11065,N_11349);
or U11701 (N_11701,N_11179,N_11162);
and U11702 (N_11702,N_11274,N_11077);
and U11703 (N_11703,N_11020,N_11378);
xor U11704 (N_11704,N_11474,N_11373);
and U11705 (N_11705,N_11061,N_11372);
or U11706 (N_11706,N_11192,N_11138);
xor U11707 (N_11707,N_11350,N_11483);
and U11708 (N_11708,N_11207,N_11329);
nand U11709 (N_11709,N_11041,N_11019);
xor U11710 (N_11710,N_11229,N_11242);
nand U11711 (N_11711,N_11409,N_11410);
xor U11712 (N_11712,N_11466,N_11321);
or U11713 (N_11713,N_11436,N_11098);
or U11714 (N_11714,N_11073,N_11331);
or U11715 (N_11715,N_11181,N_11303);
nand U11716 (N_11716,N_11254,N_11328);
xor U11717 (N_11717,N_11097,N_11396);
xnor U11718 (N_11718,N_11096,N_11055);
xnor U11719 (N_11719,N_11069,N_11498);
nand U11720 (N_11720,N_11293,N_11283);
nand U11721 (N_11721,N_11230,N_11322);
and U11722 (N_11722,N_11014,N_11301);
or U11723 (N_11723,N_11003,N_11380);
nor U11724 (N_11724,N_11379,N_11174);
nand U11725 (N_11725,N_11312,N_11314);
nand U11726 (N_11726,N_11012,N_11401);
and U11727 (N_11727,N_11499,N_11345);
nand U11728 (N_11728,N_11187,N_11046);
nand U11729 (N_11729,N_11310,N_11145);
nor U11730 (N_11730,N_11214,N_11332);
nor U11731 (N_11731,N_11326,N_11132);
or U11732 (N_11732,N_11129,N_11494);
nand U11733 (N_11733,N_11130,N_11147);
nor U11734 (N_11734,N_11366,N_11076);
nand U11735 (N_11735,N_11045,N_11033);
xnor U11736 (N_11736,N_11143,N_11267);
and U11737 (N_11737,N_11266,N_11355);
nor U11738 (N_11738,N_11272,N_11451);
nor U11739 (N_11739,N_11459,N_11091);
and U11740 (N_11740,N_11112,N_11381);
nor U11741 (N_11741,N_11231,N_11342);
and U11742 (N_11742,N_11438,N_11038);
xor U11743 (N_11743,N_11284,N_11119);
and U11744 (N_11744,N_11299,N_11278);
xor U11745 (N_11745,N_11492,N_11356);
xor U11746 (N_11746,N_11149,N_11210);
nor U11747 (N_11747,N_11133,N_11255);
nor U11748 (N_11748,N_11262,N_11478);
xnor U11749 (N_11749,N_11432,N_11404);
nor U11750 (N_11750,N_11171,N_11417);
xnor U11751 (N_11751,N_11424,N_11173);
nand U11752 (N_11752,N_11085,N_11206);
and U11753 (N_11753,N_11473,N_11141);
nand U11754 (N_11754,N_11324,N_11389);
nand U11755 (N_11755,N_11171,N_11315);
xor U11756 (N_11756,N_11467,N_11465);
xnor U11757 (N_11757,N_11180,N_11055);
or U11758 (N_11758,N_11123,N_11101);
xnor U11759 (N_11759,N_11431,N_11365);
and U11760 (N_11760,N_11382,N_11435);
and U11761 (N_11761,N_11495,N_11065);
and U11762 (N_11762,N_11486,N_11234);
xnor U11763 (N_11763,N_11015,N_11296);
and U11764 (N_11764,N_11137,N_11224);
and U11765 (N_11765,N_11279,N_11230);
nand U11766 (N_11766,N_11129,N_11431);
and U11767 (N_11767,N_11321,N_11469);
and U11768 (N_11768,N_11297,N_11147);
xor U11769 (N_11769,N_11173,N_11305);
nor U11770 (N_11770,N_11329,N_11369);
nand U11771 (N_11771,N_11081,N_11198);
or U11772 (N_11772,N_11160,N_11323);
xor U11773 (N_11773,N_11137,N_11092);
nand U11774 (N_11774,N_11180,N_11275);
nand U11775 (N_11775,N_11269,N_11033);
nand U11776 (N_11776,N_11442,N_11016);
nand U11777 (N_11777,N_11075,N_11103);
nor U11778 (N_11778,N_11276,N_11047);
or U11779 (N_11779,N_11477,N_11459);
xor U11780 (N_11780,N_11224,N_11159);
and U11781 (N_11781,N_11486,N_11340);
or U11782 (N_11782,N_11133,N_11215);
or U11783 (N_11783,N_11151,N_11388);
or U11784 (N_11784,N_11116,N_11496);
xor U11785 (N_11785,N_11451,N_11281);
xnor U11786 (N_11786,N_11279,N_11428);
xor U11787 (N_11787,N_11286,N_11260);
nor U11788 (N_11788,N_11464,N_11123);
or U11789 (N_11789,N_11444,N_11402);
nor U11790 (N_11790,N_11440,N_11462);
nor U11791 (N_11791,N_11464,N_11046);
or U11792 (N_11792,N_11083,N_11047);
nand U11793 (N_11793,N_11015,N_11470);
nor U11794 (N_11794,N_11222,N_11171);
or U11795 (N_11795,N_11023,N_11282);
nand U11796 (N_11796,N_11341,N_11241);
or U11797 (N_11797,N_11316,N_11076);
xnor U11798 (N_11798,N_11285,N_11036);
xnor U11799 (N_11799,N_11147,N_11432);
and U11800 (N_11800,N_11274,N_11004);
nand U11801 (N_11801,N_11419,N_11298);
and U11802 (N_11802,N_11352,N_11167);
nand U11803 (N_11803,N_11476,N_11150);
nand U11804 (N_11804,N_11349,N_11214);
and U11805 (N_11805,N_11138,N_11403);
nand U11806 (N_11806,N_11104,N_11356);
or U11807 (N_11807,N_11461,N_11491);
or U11808 (N_11808,N_11388,N_11041);
nor U11809 (N_11809,N_11277,N_11382);
and U11810 (N_11810,N_11217,N_11330);
or U11811 (N_11811,N_11330,N_11111);
nand U11812 (N_11812,N_11141,N_11152);
and U11813 (N_11813,N_11209,N_11213);
or U11814 (N_11814,N_11279,N_11409);
nand U11815 (N_11815,N_11045,N_11253);
nand U11816 (N_11816,N_11463,N_11113);
nor U11817 (N_11817,N_11241,N_11215);
nor U11818 (N_11818,N_11407,N_11127);
xor U11819 (N_11819,N_11188,N_11061);
nor U11820 (N_11820,N_11299,N_11339);
nand U11821 (N_11821,N_11311,N_11435);
nand U11822 (N_11822,N_11163,N_11188);
nand U11823 (N_11823,N_11244,N_11005);
or U11824 (N_11824,N_11146,N_11427);
xor U11825 (N_11825,N_11447,N_11005);
xor U11826 (N_11826,N_11423,N_11082);
xnor U11827 (N_11827,N_11000,N_11040);
or U11828 (N_11828,N_11293,N_11104);
nor U11829 (N_11829,N_11160,N_11215);
nor U11830 (N_11830,N_11288,N_11180);
nand U11831 (N_11831,N_11013,N_11339);
and U11832 (N_11832,N_11138,N_11179);
xnor U11833 (N_11833,N_11434,N_11246);
xor U11834 (N_11834,N_11064,N_11133);
or U11835 (N_11835,N_11369,N_11056);
or U11836 (N_11836,N_11410,N_11379);
or U11837 (N_11837,N_11295,N_11113);
and U11838 (N_11838,N_11152,N_11065);
nor U11839 (N_11839,N_11123,N_11213);
nand U11840 (N_11840,N_11227,N_11349);
nor U11841 (N_11841,N_11367,N_11227);
nor U11842 (N_11842,N_11399,N_11102);
and U11843 (N_11843,N_11318,N_11381);
and U11844 (N_11844,N_11421,N_11281);
or U11845 (N_11845,N_11323,N_11422);
and U11846 (N_11846,N_11297,N_11213);
nand U11847 (N_11847,N_11166,N_11467);
or U11848 (N_11848,N_11264,N_11337);
or U11849 (N_11849,N_11366,N_11441);
or U11850 (N_11850,N_11132,N_11437);
or U11851 (N_11851,N_11490,N_11299);
and U11852 (N_11852,N_11359,N_11298);
nor U11853 (N_11853,N_11245,N_11376);
or U11854 (N_11854,N_11063,N_11239);
nand U11855 (N_11855,N_11053,N_11050);
nor U11856 (N_11856,N_11072,N_11333);
nand U11857 (N_11857,N_11454,N_11300);
nor U11858 (N_11858,N_11165,N_11007);
nor U11859 (N_11859,N_11151,N_11164);
or U11860 (N_11860,N_11255,N_11006);
nor U11861 (N_11861,N_11288,N_11169);
nor U11862 (N_11862,N_11447,N_11101);
nor U11863 (N_11863,N_11379,N_11363);
or U11864 (N_11864,N_11123,N_11282);
nor U11865 (N_11865,N_11091,N_11025);
or U11866 (N_11866,N_11318,N_11405);
nor U11867 (N_11867,N_11492,N_11357);
and U11868 (N_11868,N_11450,N_11116);
or U11869 (N_11869,N_11095,N_11002);
or U11870 (N_11870,N_11065,N_11260);
nor U11871 (N_11871,N_11339,N_11014);
or U11872 (N_11872,N_11072,N_11364);
nor U11873 (N_11873,N_11290,N_11401);
or U11874 (N_11874,N_11262,N_11358);
nand U11875 (N_11875,N_11159,N_11177);
nand U11876 (N_11876,N_11090,N_11357);
nand U11877 (N_11877,N_11209,N_11100);
or U11878 (N_11878,N_11107,N_11089);
or U11879 (N_11879,N_11212,N_11462);
nor U11880 (N_11880,N_11239,N_11160);
nor U11881 (N_11881,N_11212,N_11308);
or U11882 (N_11882,N_11087,N_11436);
nand U11883 (N_11883,N_11422,N_11066);
xnor U11884 (N_11884,N_11166,N_11362);
xnor U11885 (N_11885,N_11381,N_11473);
nor U11886 (N_11886,N_11390,N_11252);
nand U11887 (N_11887,N_11039,N_11422);
or U11888 (N_11888,N_11326,N_11101);
and U11889 (N_11889,N_11158,N_11129);
or U11890 (N_11890,N_11374,N_11042);
and U11891 (N_11891,N_11144,N_11470);
nand U11892 (N_11892,N_11073,N_11053);
and U11893 (N_11893,N_11158,N_11359);
and U11894 (N_11894,N_11428,N_11424);
or U11895 (N_11895,N_11195,N_11120);
nand U11896 (N_11896,N_11312,N_11465);
nor U11897 (N_11897,N_11207,N_11281);
xnor U11898 (N_11898,N_11484,N_11476);
xnor U11899 (N_11899,N_11499,N_11224);
nor U11900 (N_11900,N_11114,N_11232);
nand U11901 (N_11901,N_11136,N_11263);
xor U11902 (N_11902,N_11214,N_11023);
and U11903 (N_11903,N_11061,N_11458);
or U11904 (N_11904,N_11324,N_11420);
xor U11905 (N_11905,N_11069,N_11375);
xor U11906 (N_11906,N_11074,N_11419);
xnor U11907 (N_11907,N_11455,N_11486);
nand U11908 (N_11908,N_11227,N_11062);
and U11909 (N_11909,N_11305,N_11085);
and U11910 (N_11910,N_11432,N_11084);
xor U11911 (N_11911,N_11256,N_11225);
nor U11912 (N_11912,N_11428,N_11169);
and U11913 (N_11913,N_11327,N_11356);
xnor U11914 (N_11914,N_11267,N_11207);
or U11915 (N_11915,N_11281,N_11378);
nor U11916 (N_11916,N_11423,N_11410);
nand U11917 (N_11917,N_11001,N_11420);
xnor U11918 (N_11918,N_11357,N_11270);
nor U11919 (N_11919,N_11138,N_11273);
nor U11920 (N_11920,N_11000,N_11371);
xor U11921 (N_11921,N_11261,N_11175);
nor U11922 (N_11922,N_11355,N_11459);
or U11923 (N_11923,N_11411,N_11410);
or U11924 (N_11924,N_11023,N_11274);
xor U11925 (N_11925,N_11487,N_11353);
and U11926 (N_11926,N_11143,N_11250);
and U11927 (N_11927,N_11351,N_11387);
nor U11928 (N_11928,N_11163,N_11078);
xnor U11929 (N_11929,N_11171,N_11123);
and U11930 (N_11930,N_11248,N_11344);
nand U11931 (N_11931,N_11206,N_11191);
xnor U11932 (N_11932,N_11433,N_11110);
or U11933 (N_11933,N_11142,N_11456);
nor U11934 (N_11934,N_11370,N_11286);
xor U11935 (N_11935,N_11444,N_11214);
nand U11936 (N_11936,N_11401,N_11154);
or U11937 (N_11937,N_11214,N_11263);
or U11938 (N_11938,N_11264,N_11358);
or U11939 (N_11939,N_11459,N_11165);
or U11940 (N_11940,N_11189,N_11096);
or U11941 (N_11941,N_11147,N_11428);
xor U11942 (N_11942,N_11401,N_11359);
nand U11943 (N_11943,N_11458,N_11420);
xor U11944 (N_11944,N_11368,N_11131);
or U11945 (N_11945,N_11059,N_11224);
xnor U11946 (N_11946,N_11111,N_11367);
and U11947 (N_11947,N_11480,N_11097);
nand U11948 (N_11948,N_11155,N_11009);
nor U11949 (N_11949,N_11175,N_11332);
nor U11950 (N_11950,N_11202,N_11292);
xnor U11951 (N_11951,N_11202,N_11479);
or U11952 (N_11952,N_11195,N_11027);
nand U11953 (N_11953,N_11457,N_11399);
and U11954 (N_11954,N_11410,N_11433);
or U11955 (N_11955,N_11205,N_11148);
xor U11956 (N_11956,N_11353,N_11305);
nor U11957 (N_11957,N_11062,N_11426);
and U11958 (N_11958,N_11271,N_11401);
nand U11959 (N_11959,N_11367,N_11100);
xor U11960 (N_11960,N_11282,N_11294);
nor U11961 (N_11961,N_11307,N_11249);
nand U11962 (N_11962,N_11407,N_11399);
nand U11963 (N_11963,N_11062,N_11269);
and U11964 (N_11964,N_11014,N_11134);
or U11965 (N_11965,N_11391,N_11287);
nand U11966 (N_11966,N_11208,N_11358);
xnor U11967 (N_11967,N_11311,N_11120);
xor U11968 (N_11968,N_11235,N_11133);
nor U11969 (N_11969,N_11134,N_11066);
nor U11970 (N_11970,N_11380,N_11452);
nor U11971 (N_11971,N_11482,N_11068);
xor U11972 (N_11972,N_11492,N_11197);
nand U11973 (N_11973,N_11493,N_11221);
or U11974 (N_11974,N_11137,N_11176);
nand U11975 (N_11975,N_11414,N_11438);
nor U11976 (N_11976,N_11342,N_11499);
or U11977 (N_11977,N_11352,N_11155);
xnor U11978 (N_11978,N_11314,N_11151);
xor U11979 (N_11979,N_11406,N_11223);
or U11980 (N_11980,N_11418,N_11432);
or U11981 (N_11981,N_11263,N_11284);
nand U11982 (N_11982,N_11102,N_11376);
nand U11983 (N_11983,N_11498,N_11261);
xor U11984 (N_11984,N_11215,N_11092);
or U11985 (N_11985,N_11053,N_11479);
nand U11986 (N_11986,N_11366,N_11307);
or U11987 (N_11987,N_11429,N_11068);
or U11988 (N_11988,N_11288,N_11473);
nand U11989 (N_11989,N_11050,N_11088);
nand U11990 (N_11990,N_11260,N_11244);
or U11991 (N_11991,N_11021,N_11365);
xnor U11992 (N_11992,N_11452,N_11125);
nand U11993 (N_11993,N_11089,N_11150);
or U11994 (N_11994,N_11412,N_11304);
nor U11995 (N_11995,N_11412,N_11424);
xor U11996 (N_11996,N_11125,N_11092);
nand U11997 (N_11997,N_11221,N_11115);
xor U11998 (N_11998,N_11349,N_11177);
xnor U11999 (N_11999,N_11125,N_11374);
xnor U12000 (N_12000,N_11799,N_11621);
nor U12001 (N_12001,N_11603,N_11806);
xor U12002 (N_12002,N_11989,N_11994);
nand U12003 (N_12003,N_11644,N_11765);
nor U12004 (N_12004,N_11899,N_11953);
nor U12005 (N_12005,N_11803,N_11564);
xnor U12006 (N_12006,N_11585,N_11533);
and U12007 (N_12007,N_11753,N_11982);
nand U12008 (N_12008,N_11938,N_11738);
nor U12009 (N_12009,N_11784,N_11816);
and U12010 (N_12010,N_11931,N_11873);
xor U12011 (N_12011,N_11665,N_11697);
nor U12012 (N_12012,N_11715,N_11721);
or U12013 (N_12013,N_11567,N_11976);
nor U12014 (N_12014,N_11595,N_11579);
and U12015 (N_12015,N_11594,N_11601);
xor U12016 (N_12016,N_11861,N_11553);
and U12017 (N_12017,N_11981,N_11760);
or U12018 (N_12018,N_11919,N_11825);
and U12019 (N_12019,N_11957,N_11705);
nand U12020 (N_12020,N_11714,N_11868);
and U12021 (N_12021,N_11850,N_11584);
or U12022 (N_12022,N_11900,N_11993);
nand U12023 (N_12023,N_11796,N_11947);
or U12024 (N_12024,N_11995,N_11649);
nor U12025 (N_12025,N_11561,N_11888);
and U12026 (N_12026,N_11679,N_11801);
or U12027 (N_12027,N_11696,N_11925);
nand U12028 (N_12028,N_11565,N_11959);
nand U12029 (N_12029,N_11548,N_11719);
nand U12030 (N_12030,N_11515,N_11988);
or U12031 (N_12031,N_11537,N_11997);
and U12032 (N_12032,N_11912,N_11883);
nor U12033 (N_12033,N_11630,N_11648);
nand U12034 (N_12034,N_11836,N_11787);
nor U12035 (N_12035,N_11757,N_11897);
and U12036 (N_12036,N_11749,N_11756);
and U12037 (N_12037,N_11597,N_11783);
or U12038 (N_12038,N_11538,N_11531);
nor U12039 (N_12039,N_11704,N_11785);
nand U12040 (N_12040,N_11881,N_11586);
and U12041 (N_12041,N_11820,N_11686);
or U12042 (N_12042,N_11987,N_11673);
xor U12043 (N_12043,N_11605,N_11827);
xor U12044 (N_12044,N_11840,N_11920);
and U12045 (N_12045,N_11914,N_11556);
or U12046 (N_12046,N_11632,N_11558);
or U12047 (N_12047,N_11598,N_11932);
nor U12048 (N_12048,N_11694,N_11950);
nor U12049 (N_12049,N_11518,N_11964);
nor U12050 (N_12050,N_11623,N_11990);
nor U12051 (N_12051,N_11517,N_11917);
and U12052 (N_12052,N_11849,N_11535);
xnor U12053 (N_12053,N_11971,N_11725);
nor U12054 (N_12054,N_11542,N_11574);
nor U12055 (N_12055,N_11748,N_11745);
xnor U12056 (N_12056,N_11527,N_11832);
nor U12057 (N_12057,N_11659,N_11855);
or U12058 (N_12058,N_11674,N_11828);
nand U12059 (N_12059,N_11812,N_11894);
nand U12060 (N_12060,N_11511,N_11602);
and U12061 (N_12061,N_11516,N_11846);
xor U12062 (N_12062,N_11751,N_11963);
nand U12063 (N_12063,N_11734,N_11670);
xor U12064 (N_12064,N_11766,N_11545);
nor U12065 (N_12065,N_11747,N_11637);
or U12066 (N_12066,N_11933,N_11552);
nor U12067 (N_12067,N_11606,N_11616);
nand U12068 (N_12068,N_11560,N_11834);
and U12069 (N_12069,N_11788,N_11918);
nor U12070 (N_12070,N_11666,N_11654);
nand U12071 (N_12071,N_11587,N_11677);
or U12072 (N_12072,N_11767,N_11774);
nor U12073 (N_12073,N_11859,N_11559);
or U12074 (N_12074,N_11829,N_11948);
or U12075 (N_12075,N_11688,N_11916);
or U12076 (N_12076,N_11737,N_11510);
nor U12077 (N_12077,N_11682,N_11877);
and U12078 (N_12078,N_11884,N_11978);
xnor U12079 (N_12079,N_11966,N_11706);
xnor U12080 (N_12080,N_11607,N_11506);
xor U12081 (N_12081,N_11724,N_11683);
or U12082 (N_12082,N_11713,N_11599);
and U12083 (N_12083,N_11856,N_11685);
xnor U12084 (N_12084,N_11944,N_11793);
xnor U12085 (N_12085,N_11811,N_11923);
xor U12086 (N_12086,N_11662,N_11936);
or U12087 (N_12087,N_11887,N_11992);
and U12088 (N_12088,N_11693,N_11610);
or U12089 (N_12089,N_11805,N_11731);
nand U12090 (N_12090,N_11795,N_11671);
or U12091 (N_12091,N_11909,N_11851);
or U12092 (N_12092,N_11740,N_11777);
nor U12093 (N_12093,N_11942,N_11698);
nor U12094 (N_12094,N_11582,N_11720);
nand U12095 (N_12095,N_11652,N_11819);
nor U12096 (N_12096,N_11779,N_11660);
nand U12097 (N_12097,N_11906,N_11875);
nor U12098 (N_12098,N_11908,N_11818);
nand U12099 (N_12099,N_11742,N_11588);
nand U12100 (N_12100,N_11858,N_11695);
xor U12101 (N_12101,N_11969,N_11879);
xnor U12102 (N_12102,N_11631,N_11580);
xnor U12103 (N_12103,N_11924,N_11629);
and U12104 (N_12104,N_11667,N_11960);
and U12105 (N_12105,N_11583,N_11501);
or U12106 (N_12106,N_11744,N_11521);
xnor U12107 (N_12107,N_11804,N_11622);
nor U12108 (N_12108,N_11904,N_11566);
nand U12109 (N_12109,N_11581,N_11741);
and U12110 (N_12110,N_11736,N_11646);
nand U12111 (N_12111,N_11718,N_11973);
nor U12112 (N_12112,N_11821,N_11650);
nor U12113 (N_12113,N_11614,N_11672);
nor U12114 (N_12114,N_11842,N_11739);
or U12115 (N_12115,N_11624,N_11937);
nor U12116 (N_12116,N_11999,N_11690);
xor U12117 (N_12117,N_11571,N_11658);
nor U12118 (N_12118,N_11536,N_11841);
or U12119 (N_12119,N_11754,N_11764);
nand U12120 (N_12120,N_11592,N_11986);
xor U12121 (N_12121,N_11589,N_11503);
xnor U12122 (N_12122,N_11655,N_11864);
nor U12123 (N_12123,N_11703,N_11551);
xnor U12124 (N_12124,N_11642,N_11845);
nand U12125 (N_12125,N_11857,N_11958);
nand U12126 (N_12126,N_11885,N_11907);
nor U12127 (N_12127,N_11604,N_11889);
and U12128 (N_12128,N_11943,N_11926);
nor U12129 (N_12129,N_11636,N_11802);
and U12130 (N_12130,N_11880,N_11955);
nand U12131 (N_12131,N_11949,N_11972);
and U12132 (N_12132,N_11500,N_11544);
xnor U12133 (N_12133,N_11522,N_11733);
nand U12134 (N_12134,N_11554,N_11869);
or U12135 (N_12135,N_11870,N_11645);
nor U12136 (N_12136,N_11555,N_11893);
and U12137 (N_12137,N_11680,N_11984);
xnor U12138 (N_12138,N_11882,N_11617);
xnor U12139 (N_12139,N_11707,N_11709);
and U12140 (N_12140,N_11525,N_11613);
xor U12141 (N_12141,N_11771,N_11915);
xor U12142 (N_12142,N_11643,N_11941);
or U12143 (N_12143,N_11626,N_11891);
nor U12144 (N_12144,N_11902,N_11886);
or U12145 (N_12145,N_11627,N_11550);
nand U12146 (N_12146,N_11901,N_11844);
and U12147 (N_12147,N_11927,N_11635);
nor U12148 (N_12148,N_11769,N_11577);
xnor U12149 (N_12149,N_11691,N_11547);
nand U12150 (N_12150,N_11833,N_11996);
and U12151 (N_12151,N_11809,N_11755);
or U12152 (N_12152,N_11968,N_11562);
nor U12153 (N_12153,N_11676,N_11529);
xor U12154 (N_12154,N_11611,N_11549);
nor U12155 (N_12155,N_11848,N_11678);
and U12156 (N_12156,N_11930,N_11839);
or U12157 (N_12157,N_11791,N_11640);
xor U12158 (N_12158,N_11615,N_11681);
xnor U12159 (N_12159,N_11639,N_11810);
and U12160 (N_12160,N_11822,N_11838);
or U12161 (N_12161,N_11952,N_11609);
nand U12162 (N_12162,N_11797,N_11961);
nand U12163 (N_12163,N_11743,N_11815);
and U12164 (N_12164,N_11540,N_11922);
nor U12165 (N_12165,N_11723,N_11770);
and U12166 (N_12166,N_11687,N_11998);
and U12167 (N_12167,N_11509,N_11702);
nor U12168 (N_12168,N_11726,N_11722);
nor U12169 (N_12169,N_11730,N_11965);
nand U12170 (N_12170,N_11700,N_11523);
and U12171 (N_12171,N_11563,N_11591);
nor U12172 (N_12172,N_11854,N_11946);
nor U12173 (N_12173,N_11534,N_11710);
xor U12174 (N_12174,N_11628,N_11573);
nand U12175 (N_12175,N_11977,N_11929);
xor U12176 (N_12176,N_11612,N_11638);
nand U12177 (N_12177,N_11541,N_11847);
and U12178 (N_12178,N_11641,N_11716);
xor U12179 (N_12179,N_11814,N_11905);
xnor U12180 (N_12180,N_11520,N_11956);
nor U12181 (N_12181,N_11800,N_11528);
nor U12182 (N_12182,N_11620,N_11962);
nor U12183 (N_12183,N_11903,N_11778);
xor U12184 (N_12184,N_11934,N_11790);
xnor U12185 (N_12185,N_11600,N_11758);
nand U12186 (N_12186,N_11664,N_11618);
and U12187 (N_12187,N_11773,N_11568);
nand U12188 (N_12188,N_11860,N_11504);
and U12189 (N_12189,N_11890,N_11576);
and U12190 (N_12190,N_11669,N_11699);
or U12191 (N_12191,N_11728,N_11507);
or U12192 (N_12192,N_11625,N_11578);
or U12193 (N_12193,N_11935,N_11975);
nand U12194 (N_12194,N_11898,N_11794);
or U12195 (N_12195,N_11813,N_11974);
nor U12196 (N_12196,N_11735,N_11911);
and U12197 (N_12197,N_11775,N_11826);
and U12198 (N_12198,N_11983,N_11852);
xor U12199 (N_12199,N_11862,N_11807);
or U12200 (N_12200,N_11980,N_11782);
nand U12201 (N_12201,N_11780,N_11653);
or U12202 (N_12202,N_11657,N_11692);
and U12203 (N_12203,N_11513,N_11608);
xnor U12204 (N_12204,N_11872,N_11940);
and U12205 (N_12205,N_11878,N_11546);
and U12206 (N_12206,N_11781,N_11786);
and U12207 (N_12207,N_11892,N_11951);
nand U12208 (N_12208,N_11557,N_11684);
nor U12209 (N_12209,N_11596,N_11619);
nand U12210 (N_12210,N_11876,N_11711);
nand U12211 (N_12211,N_11824,N_11746);
and U12212 (N_12212,N_11656,N_11837);
xor U12213 (N_12213,N_11570,N_11729);
xor U12214 (N_12214,N_11633,N_11835);
nand U12215 (N_12215,N_11865,N_11543);
or U12216 (N_12216,N_11896,N_11817);
nand U12217 (N_12217,N_11830,N_11689);
or U12218 (N_12218,N_11789,N_11939);
xnor U12219 (N_12219,N_11539,N_11514);
or U12220 (N_12220,N_11593,N_11651);
or U12221 (N_12221,N_11921,N_11863);
xor U12222 (N_12222,N_11843,N_11967);
xnor U12223 (N_12223,N_11575,N_11675);
nor U12224 (N_12224,N_11895,N_11505);
nand U12225 (N_12225,N_11763,N_11732);
nand U12226 (N_12226,N_11910,N_11727);
nand U12227 (N_12227,N_11762,N_11717);
and U12228 (N_12228,N_11768,N_11772);
and U12229 (N_12229,N_11831,N_11970);
xnor U12230 (N_12230,N_11712,N_11752);
nand U12231 (N_12231,N_11945,N_11798);
nor U12232 (N_12232,N_11572,N_11663);
nor U12233 (N_12233,N_11502,N_11808);
nor U12234 (N_12234,N_11524,N_11867);
or U12235 (N_12235,N_11532,N_11750);
nand U12236 (N_12236,N_11759,N_11985);
xor U12237 (N_12237,N_11874,N_11913);
and U12238 (N_12238,N_11928,N_11661);
or U12239 (N_12239,N_11823,N_11866);
and U12240 (N_12240,N_11668,N_11776);
nand U12241 (N_12241,N_11526,N_11569);
nor U12242 (N_12242,N_11647,N_11519);
nor U12243 (N_12243,N_11792,N_11530);
or U12244 (N_12244,N_11701,N_11708);
nand U12245 (N_12245,N_11853,N_11590);
nor U12246 (N_12246,N_11508,N_11991);
nor U12247 (N_12247,N_11634,N_11954);
or U12248 (N_12248,N_11512,N_11979);
and U12249 (N_12249,N_11871,N_11761);
nand U12250 (N_12250,N_11866,N_11876);
and U12251 (N_12251,N_11633,N_11753);
xnor U12252 (N_12252,N_11832,N_11636);
or U12253 (N_12253,N_11755,N_11743);
nor U12254 (N_12254,N_11626,N_11613);
and U12255 (N_12255,N_11715,N_11630);
and U12256 (N_12256,N_11676,N_11761);
nand U12257 (N_12257,N_11531,N_11752);
and U12258 (N_12258,N_11847,N_11975);
xnor U12259 (N_12259,N_11598,N_11747);
xnor U12260 (N_12260,N_11637,N_11595);
xor U12261 (N_12261,N_11604,N_11691);
or U12262 (N_12262,N_11600,N_11617);
nor U12263 (N_12263,N_11917,N_11525);
nand U12264 (N_12264,N_11697,N_11727);
or U12265 (N_12265,N_11907,N_11756);
or U12266 (N_12266,N_11606,N_11866);
or U12267 (N_12267,N_11614,N_11625);
xnor U12268 (N_12268,N_11848,N_11923);
nand U12269 (N_12269,N_11537,N_11565);
nand U12270 (N_12270,N_11969,N_11583);
and U12271 (N_12271,N_11835,N_11762);
nor U12272 (N_12272,N_11821,N_11558);
or U12273 (N_12273,N_11974,N_11687);
and U12274 (N_12274,N_11883,N_11664);
xnor U12275 (N_12275,N_11577,N_11813);
nor U12276 (N_12276,N_11917,N_11983);
and U12277 (N_12277,N_11803,N_11589);
or U12278 (N_12278,N_11880,N_11577);
or U12279 (N_12279,N_11958,N_11601);
nand U12280 (N_12280,N_11689,N_11571);
nor U12281 (N_12281,N_11882,N_11829);
and U12282 (N_12282,N_11918,N_11775);
nand U12283 (N_12283,N_11510,N_11998);
xor U12284 (N_12284,N_11773,N_11698);
xor U12285 (N_12285,N_11826,N_11691);
nand U12286 (N_12286,N_11998,N_11503);
nand U12287 (N_12287,N_11512,N_11596);
nor U12288 (N_12288,N_11802,N_11562);
xnor U12289 (N_12289,N_11732,N_11765);
xnor U12290 (N_12290,N_11999,N_11978);
nor U12291 (N_12291,N_11789,N_11512);
nor U12292 (N_12292,N_11583,N_11869);
and U12293 (N_12293,N_11788,N_11841);
or U12294 (N_12294,N_11836,N_11540);
xnor U12295 (N_12295,N_11542,N_11838);
nor U12296 (N_12296,N_11853,N_11793);
xnor U12297 (N_12297,N_11671,N_11604);
nand U12298 (N_12298,N_11581,N_11665);
xnor U12299 (N_12299,N_11639,N_11624);
nor U12300 (N_12300,N_11819,N_11505);
xor U12301 (N_12301,N_11874,N_11987);
and U12302 (N_12302,N_11958,N_11840);
xnor U12303 (N_12303,N_11545,N_11853);
xor U12304 (N_12304,N_11695,N_11618);
and U12305 (N_12305,N_11647,N_11701);
xnor U12306 (N_12306,N_11631,N_11783);
xnor U12307 (N_12307,N_11886,N_11821);
xnor U12308 (N_12308,N_11567,N_11762);
nor U12309 (N_12309,N_11951,N_11630);
nor U12310 (N_12310,N_11857,N_11935);
nor U12311 (N_12311,N_11917,N_11945);
and U12312 (N_12312,N_11962,N_11730);
and U12313 (N_12313,N_11643,N_11740);
and U12314 (N_12314,N_11950,N_11586);
nor U12315 (N_12315,N_11692,N_11773);
nand U12316 (N_12316,N_11798,N_11548);
or U12317 (N_12317,N_11842,N_11621);
nand U12318 (N_12318,N_11678,N_11620);
or U12319 (N_12319,N_11885,N_11917);
or U12320 (N_12320,N_11576,N_11504);
xnor U12321 (N_12321,N_11757,N_11912);
xnor U12322 (N_12322,N_11807,N_11500);
or U12323 (N_12323,N_11545,N_11964);
xnor U12324 (N_12324,N_11890,N_11740);
nand U12325 (N_12325,N_11961,N_11660);
or U12326 (N_12326,N_11721,N_11946);
nor U12327 (N_12327,N_11901,N_11870);
nand U12328 (N_12328,N_11952,N_11900);
or U12329 (N_12329,N_11760,N_11851);
nand U12330 (N_12330,N_11635,N_11725);
or U12331 (N_12331,N_11968,N_11554);
and U12332 (N_12332,N_11946,N_11671);
and U12333 (N_12333,N_11917,N_11815);
nor U12334 (N_12334,N_11864,N_11782);
nor U12335 (N_12335,N_11523,N_11570);
and U12336 (N_12336,N_11645,N_11886);
and U12337 (N_12337,N_11875,N_11970);
or U12338 (N_12338,N_11960,N_11844);
xnor U12339 (N_12339,N_11581,N_11854);
or U12340 (N_12340,N_11853,N_11755);
and U12341 (N_12341,N_11647,N_11769);
or U12342 (N_12342,N_11857,N_11968);
and U12343 (N_12343,N_11973,N_11966);
nand U12344 (N_12344,N_11757,N_11529);
and U12345 (N_12345,N_11836,N_11791);
nor U12346 (N_12346,N_11668,N_11883);
nand U12347 (N_12347,N_11723,N_11924);
and U12348 (N_12348,N_11942,N_11915);
and U12349 (N_12349,N_11843,N_11793);
xnor U12350 (N_12350,N_11934,N_11525);
or U12351 (N_12351,N_11672,N_11946);
or U12352 (N_12352,N_11502,N_11901);
and U12353 (N_12353,N_11786,N_11915);
nand U12354 (N_12354,N_11838,N_11839);
nor U12355 (N_12355,N_11839,N_11812);
xnor U12356 (N_12356,N_11527,N_11825);
nand U12357 (N_12357,N_11523,N_11685);
and U12358 (N_12358,N_11679,N_11953);
and U12359 (N_12359,N_11681,N_11955);
and U12360 (N_12360,N_11625,N_11721);
nand U12361 (N_12361,N_11524,N_11960);
nand U12362 (N_12362,N_11538,N_11681);
xor U12363 (N_12363,N_11813,N_11658);
nor U12364 (N_12364,N_11752,N_11994);
or U12365 (N_12365,N_11861,N_11598);
xnor U12366 (N_12366,N_11801,N_11788);
xnor U12367 (N_12367,N_11979,N_11593);
nand U12368 (N_12368,N_11863,N_11868);
nor U12369 (N_12369,N_11538,N_11794);
and U12370 (N_12370,N_11551,N_11926);
xor U12371 (N_12371,N_11590,N_11612);
and U12372 (N_12372,N_11963,N_11627);
xnor U12373 (N_12373,N_11630,N_11547);
and U12374 (N_12374,N_11858,N_11564);
xnor U12375 (N_12375,N_11559,N_11504);
nand U12376 (N_12376,N_11653,N_11858);
or U12377 (N_12377,N_11532,N_11641);
or U12378 (N_12378,N_11974,N_11748);
or U12379 (N_12379,N_11914,N_11736);
or U12380 (N_12380,N_11539,N_11675);
nand U12381 (N_12381,N_11871,N_11782);
xor U12382 (N_12382,N_11769,N_11943);
or U12383 (N_12383,N_11648,N_11612);
nand U12384 (N_12384,N_11879,N_11527);
nand U12385 (N_12385,N_11704,N_11580);
nand U12386 (N_12386,N_11919,N_11630);
xnor U12387 (N_12387,N_11995,N_11857);
nand U12388 (N_12388,N_11619,N_11828);
nor U12389 (N_12389,N_11939,N_11903);
and U12390 (N_12390,N_11955,N_11593);
nand U12391 (N_12391,N_11782,N_11601);
or U12392 (N_12392,N_11855,N_11988);
xnor U12393 (N_12393,N_11606,N_11560);
xor U12394 (N_12394,N_11676,N_11720);
nand U12395 (N_12395,N_11961,N_11600);
nand U12396 (N_12396,N_11637,N_11639);
and U12397 (N_12397,N_11735,N_11803);
nor U12398 (N_12398,N_11757,N_11732);
and U12399 (N_12399,N_11889,N_11579);
xor U12400 (N_12400,N_11932,N_11946);
xor U12401 (N_12401,N_11520,N_11602);
xor U12402 (N_12402,N_11510,N_11756);
and U12403 (N_12403,N_11865,N_11822);
nand U12404 (N_12404,N_11736,N_11522);
or U12405 (N_12405,N_11872,N_11934);
xor U12406 (N_12406,N_11905,N_11729);
nor U12407 (N_12407,N_11662,N_11620);
xor U12408 (N_12408,N_11952,N_11756);
and U12409 (N_12409,N_11537,N_11824);
xor U12410 (N_12410,N_11663,N_11885);
xnor U12411 (N_12411,N_11954,N_11721);
and U12412 (N_12412,N_11891,N_11587);
nand U12413 (N_12413,N_11588,N_11737);
xnor U12414 (N_12414,N_11922,N_11766);
and U12415 (N_12415,N_11944,N_11997);
xor U12416 (N_12416,N_11906,N_11821);
nor U12417 (N_12417,N_11796,N_11777);
and U12418 (N_12418,N_11651,N_11613);
or U12419 (N_12419,N_11508,N_11788);
and U12420 (N_12420,N_11929,N_11511);
or U12421 (N_12421,N_11522,N_11545);
nor U12422 (N_12422,N_11899,N_11961);
and U12423 (N_12423,N_11742,N_11714);
xnor U12424 (N_12424,N_11854,N_11716);
nor U12425 (N_12425,N_11784,N_11601);
or U12426 (N_12426,N_11747,N_11750);
nor U12427 (N_12427,N_11964,N_11775);
xor U12428 (N_12428,N_11709,N_11641);
nor U12429 (N_12429,N_11657,N_11795);
and U12430 (N_12430,N_11910,N_11553);
nand U12431 (N_12431,N_11851,N_11978);
and U12432 (N_12432,N_11856,N_11666);
xnor U12433 (N_12433,N_11753,N_11621);
or U12434 (N_12434,N_11595,N_11799);
xor U12435 (N_12435,N_11819,N_11574);
or U12436 (N_12436,N_11865,N_11534);
or U12437 (N_12437,N_11605,N_11540);
nand U12438 (N_12438,N_11613,N_11994);
and U12439 (N_12439,N_11735,N_11647);
and U12440 (N_12440,N_11758,N_11909);
and U12441 (N_12441,N_11770,N_11965);
nand U12442 (N_12442,N_11758,N_11925);
nand U12443 (N_12443,N_11528,N_11563);
nor U12444 (N_12444,N_11968,N_11810);
xor U12445 (N_12445,N_11698,N_11896);
xor U12446 (N_12446,N_11834,N_11829);
nor U12447 (N_12447,N_11725,N_11738);
nor U12448 (N_12448,N_11847,N_11856);
nor U12449 (N_12449,N_11705,N_11944);
xnor U12450 (N_12450,N_11694,N_11843);
nor U12451 (N_12451,N_11571,N_11784);
xor U12452 (N_12452,N_11695,N_11883);
xor U12453 (N_12453,N_11880,N_11544);
xnor U12454 (N_12454,N_11742,N_11846);
xor U12455 (N_12455,N_11531,N_11611);
xnor U12456 (N_12456,N_11840,N_11993);
and U12457 (N_12457,N_11726,N_11876);
and U12458 (N_12458,N_11567,N_11909);
and U12459 (N_12459,N_11861,N_11761);
or U12460 (N_12460,N_11898,N_11817);
nand U12461 (N_12461,N_11758,N_11715);
and U12462 (N_12462,N_11768,N_11556);
nand U12463 (N_12463,N_11912,N_11960);
nor U12464 (N_12464,N_11642,N_11958);
nand U12465 (N_12465,N_11806,N_11731);
nor U12466 (N_12466,N_11707,N_11913);
or U12467 (N_12467,N_11915,N_11716);
xor U12468 (N_12468,N_11992,N_11863);
nand U12469 (N_12469,N_11794,N_11562);
nand U12470 (N_12470,N_11660,N_11752);
xnor U12471 (N_12471,N_11790,N_11800);
and U12472 (N_12472,N_11712,N_11933);
nand U12473 (N_12473,N_11560,N_11756);
xnor U12474 (N_12474,N_11683,N_11976);
nand U12475 (N_12475,N_11721,N_11898);
and U12476 (N_12476,N_11603,N_11926);
xnor U12477 (N_12477,N_11640,N_11594);
nor U12478 (N_12478,N_11565,N_11784);
xnor U12479 (N_12479,N_11988,N_11688);
nand U12480 (N_12480,N_11779,N_11908);
nand U12481 (N_12481,N_11649,N_11545);
or U12482 (N_12482,N_11758,N_11763);
nand U12483 (N_12483,N_11669,N_11705);
nand U12484 (N_12484,N_11803,N_11892);
and U12485 (N_12485,N_11623,N_11726);
nand U12486 (N_12486,N_11957,N_11929);
xor U12487 (N_12487,N_11594,N_11856);
nor U12488 (N_12488,N_11824,N_11769);
and U12489 (N_12489,N_11703,N_11507);
nand U12490 (N_12490,N_11980,N_11950);
nand U12491 (N_12491,N_11735,N_11555);
xnor U12492 (N_12492,N_11709,N_11919);
xor U12493 (N_12493,N_11660,N_11872);
or U12494 (N_12494,N_11578,N_11769);
nand U12495 (N_12495,N_11695,N_11922);
nor U12496 (N_12496,N_11889,N_11780);
or U12497 (N_12497,N_11679,N_11505);
xor U12498 (N_12498,N_11764,N_11635);
xnor U12499 (N_12499,N_11692,N_11911);
or U12500 (N_12500,N_12067,N_12339);
and U12501 (N_12501,N_12368,N_12159);
and U12502 (N_12502,N_12007,N_12234);
and U12503 (N_12503,N_12393,N_12207);
nor U12504 (N_12504,N_12068,N_12020);
xor U12505 (N_12505,N_12492,N_12484);
or U12506 (N_12506,N_12422,N_12309);
nor U12507 (N_12507,N_12448,N_12366);
nor U12508 (N_12508,N_12015,N_12130);
or U12509 (N_12509,N_12071,N_12299);
and U12510 (N_12510,N_12144,N_12257);
and U12511 (N_12511,N_12146,N_12433);
xnor U12512 (N_12512,N_12218,N_12210);
xnor U12513 (N_12513,N_12051,N_12367);
and U12514 (N_12514,N_12010,N_12415);
or U12515 (N_12515,N_12135,N_12466);
and U12516 (N_12516,N_12246,N_12248);
xnor U12517 (N_12517,N_12410,N_12486);
or U12518 (N_12518,N_12446,N_12385);
nor U12519 (N_12519,N_12495,N_12464);
or U12520 (N_12520,N_12379,N_12077);
nor U12521 (N_12521,N_12217,N_12400);
and U12522 (N_12522,N_12437,N_12178);
nand U12523 (N_12523,N_12037,N_12241);
xor U12524 (N_12524,N_12424,N_12447);
xor U12525 (N_12525,N_12006,N_12046);
xor U12526 (N_12526,N_12341,N_12202);
xor U12527 (N_12527,N_12190,N_12434);
nor U12528 (N_12528,N_12426,N_12087);
and U12529 (N_12529,N_12454,N_12265);
or U12530 (N_12530,N_12014,N_12444);
nand U12531 (N_12531,N_12099,N_12171);
and U12532 (N_12532,N_12009,N_12342);
and U12533 (N_12533,N_12002,N_12222);
and U12534 (N_12534,N_12312,N_12094);
and U12535 (N_12535,N_12462,N_12364);
nand U12536 (N_12536,N_12096,N_12066);
nand U12537 (N_12537,N_12485,N_12028);
or U12538 (N_12538,N_12070,N_12494);
nor U12539 (N_12539,N_12081,N_12295);
nand U12540 (N_12540,N_12329,N_12402);
xor U12541 (N_12541,N_12199,N_12086);
and U12542 (N_12542,N_12291,N_12122);
nor U12543 (N_12543,N_12307,N_12155);
and U12544 (N_12544,N_12269,N_12004);
xor U12545 (N_12545,N_12267,N_12441);
nand U12546 (N_12546,N_12056,N_12397);
and U12547 (N_12547,N_12145,N_12252);
nand U12548 (N_12548,N_12496,N_12074);
nor U12549 (N_12549,N_12351,N_12432);
nand U12550 (N_12550,N_12209,N_12374);
xnor U12551 (N_12551,N_12325,N_12188);
nor U12552 (N_12552,N_12182,N_12132);
xor U12553 (N_12553,N_12301,N_12305);
nor U12554 (N_12554,N_12005,N_12442);
nand U12555 (N_12555,N_12160,N_12230);
nor U12556 (N_12556,N_12233,N_12103);
and U12557 (N_12557,N_12359,N_12224);
xor U12558 (N_12558,N_12438,N_12244);
and U12559 (N_12559,N_12360,N_12034);
xor U12560 (N_12560,N_12197,N_12126);
xor U12561 (N_12561,N_12152,N_12060);
xnor U12562 (N_12562,N_12176,N_12012);
and U12563 (N_12563,N_12475,N_12377);
nor U12564 (N_12564,N_12044,N_12327);
nor U12565 (N_12565,N_12030,N_12451);
or U12566 (N_12566,N_12105,N_12019);
or U12567 (N_12567,N_12247,N_12289);
nand U12568 (N_12568,N_12482,N_12052);
or U12569 (N_12569,N_12361,N_12365);
nor U12570 (N_12570,N_12389,N_12293);
nor U12571 (N_12571,N_12181,N_12065);
or U12572 (N_12572,N_12443,N_12184);
and U12573 (N_12573,N_12064,N_12386);
or U12574 (N_12574,N_12189,N_12287);
or U12575 (N_12575,N_12203,N_12177);
and U12576 (N_12576,N_12027,N_12343);
nor U12577 (N_12577,N_12076,N_12461);
nand U12578 (N_12578,N_12294,N_12480);
nand U12579 (N_12579,N_12399,N_12032);
xnor U12580 (N_12580,N_12084,N_12409);
or U12581 (N_12581,N_12469,N_12185);
nand U12582 (N_12582,N_12430,N_12198);
xor U12583 (N_12583,N_12110,N_12452);
or U12584 (N_12584,N_12137,N_12290);
nand U12585 (N_12585,N_12292,N_12125);
nand U12586 (N_12586,N_12208,N_12211);
xnor U12587 (N_12587,N_12180,N_12196);
xor U12588 (N_12588,N_12420,N_12022);
or U12589 (N_12589,N_12035,N_12033);
or U12590 (N_12590,N_12149,N_12384);
nor U12591 (N_12591,N_12334,N_12322);
or U12592 (N_12592,N_12405,N_12428);
or U12593 (N_12593,N_12375,N_12349);
or U12594 (N_12594,N_12128,N_12314);
nor U12595 (N_12595,N_12062,N_12254);
and U12596 (N_12596,N_12238,N_12416);
xnor U12597 (N_12597,N_12085,N_12371);
nand U12598 (N_12598,N_12091,N_12156);
nand U12599 (N_12599,N_12073,N_12131);
xnor U12600 (N_12600,N_12383,N_12355);
nor U12601 (N_12601,N_12106,N_12088);
or U12602 (N_12602,N_12338,N_12459);
nor U12603 (N_12603,N_12150,N_12281);
xnor U12604 (N_12604,N_12200,N_12258);
nand U12605 (N_12605,N_12411,N_12038);
and U12606 (N_12606,N_12460,N_12001);
nor U12607 (N_12607,N_12205,N_12401);
nand U12608 (N_12608,N_12260,N_12245);
xnor U12609 (N_12609,N_12324,N_12148);
nand U12610 (N_12610,N_12163,N_12332);
nor U12611 (N_12611,N_12192,N_12276);
xnor U12612 (N_12612,N_12382,N_12118);
xnor U12613 (N_12613,N_12151,N_12194);
xor U12614 (N_12614,N_12412,N_12302);
nand U12615 (N_12615,N_12107,N_12288);
nor U12616 (N_12616,N_12278,N_12256);
and U12617 (N_12617,N_12213,N_12483);
nand U12618 (N_12618,N_12271,N_12346);
nand U12619 (N_12619,N_12072,N_12390);
and U12620 (N_12620,N_12057,N_12116);
nand U12621 (N_12621,N_12284,N_12372);
nand U12622 (N_12622,N_12021,N_12493);
nand U12623 (N_12623,N_12311,N_12471);
and U12624 (N_12624,N_12134,N_12303);
or U12625 (N_12625,N_12179,N_12232);
and U12626 (N_12626,N_12499,N_12018);
xor U12627 (N_12627,N_12011,N_12280);
nand U12628 (N_12628,N_12075,N_12221);
nor U12629 (N_12629,N_12223,N_12120);
xnor U12630 (N_12630,N_12488,N_12285);
nand U12631 (N_12631,N_12093,N_12111);
or U12632 (N_12632,N_12440,N_12380);
or U12633 (N_12633,N_12100,N_12138);
nand U12634 (N_12634,N_12490,N_12362);
xnor U12635 (N_12635,N_12348,N_12396);
nand U12636 (N_12636,N_12042,N_12251);
nor U12637 (N_12637,N_12472,N_12392);
xnor U12638 (N_12638,N_12262,N_12369);
nand U12639 (N_12639,N_12083,N_12215);
and U12640 (N_12640,N_12395,N_12175);
xnor U12641 (N_12641,N_12054,N_12336);
nor U12642 (N_12642,N_12363,N_12306);
nand U12643 (N_12643,N_12136,N_12388);
or U12644 (N_12644,N_12310,N_12457);
nand U12645 (N_12645,N_12477,N_12227);
nor U12646 (N_12646,N_12226,N_12425);
nor U12647 (N_12647,N_12450,N_12220);
nand U12648 (N_12648,N_12193,N_12055);
nand U12649 (N_12649,N_12089,N_12268);
nand U12650 (N_12650,N_12167,N_12166);
and U12651 (N_12651,N_12250,N_12406);
and U12652 (N_12652,N_12261,N_12398);
nand U12653 (N_12653,N_12157,N_12162);
or U12654 (N_12654,N_12195,N_12318);
nand U12655 (N_12655,N_12468,N_12139);
or U12656 (N_12656,N_12041,N_12031);
nand U12657 (N_12657,N_12102,N_12029);
nand U12658 (N_12658,N_12259,N_12161);
nor U12659 (N_12659,N_12169,N_12236);
xnor U12660 (N_12660,N_12147,N_12431);
xor U12661 (N_12661,N_12212,N_12242);
nor U12662 (N_12662,N_12376,N_12225);
nand U12663 (N_12663,N_12092,N_12140);
nand U12664 (N_12664,N_12174,N_12117);
or U12665 (N_12665,N_12283,N_12418);
nor U12666 (N_12666,N_12297,N_12344);
nor U12667 (N_12667,N_12404,N_12330);
nand U12668 (N_12668,N_12264,N_12298);
or U12669 (N_12669,N_12273,N_12417);
xnor U12670 (N_12670,N_12481,N_12497);
nand U12671 (N_12671,N_12164,N_12228);
or U12672 (N_12672,N_12082,N_12239);
or U12673 (N_12673,N_12333,N_12063);
or U12674 (N_12674,N_12023,N_12413);
xnor U12675 (N_12675,N_12045,N_12328);
nor U12676 (N_12676,N_12263,N_12394);
and U12677 (N_12677,N_12479,N_12455);
nand U12678 (N_12678,N_12243,N_12079);
xnor U12679 (N_12679,N_12317,N_12331);
nor U12680 (N_12680,N_12097,N_12313);
xnor U12681 (N_12681,N_12121,N_12219);
xor U12682 (N_12682,N_12487,N_12141);
nand U12683 (N_12683,N_12326,N_12000);
xnor U12684 (N_12684,N_12016,N_12143);
nand U12685 (N_12685,N_12498,N_12090);
and U12686 (N_12686,N_12003,N_12489);
xor U12687 (N_12687,N_12323,N_12319);
nand U12688 (N_12688,N_12058,N_12080);
and U12689 (N_12689,N_12115,N_12237);
nor U12690 (N_12690,N_12240,N_12008);
xor U12691 (N_12691,N_12391,N_12059);
nor U12692 (N_12692,N_12049,N_12204);
xnor U12693 (N_12693,N_12119,N_12186);
or U12694 (N_12694,N_12286,N_12114);
nor U12695 (N_12695,N_12229,N_12255);
xnor U12696 (N_12696,N_12275,N_12113);
and U12697 (N_12697,N_12026,N_12463);
nand U12698 (N_12698,N_12474,N_12017);
nor U12699 (N_12699,N_12191,N_12095);
nand U12700 (N_12700,N_12040,N_12345);
and U12701 (N_12701,N_12387,N_12340);
xor U12702 (N_12702,N_12129,N_12353);
and U12703 (N_12703,N_12172,N_12108);
or U12704 (N_12704,N_12036,N_12414);
xnor U12705 (N_12705,N_12216,N_12133);
nand U12706 (N_12706,N_12421,N_12043);
or U12707 (N_12707,N_12347,N_12335);
and U12708 (N_12708,N_12170,N_12025);
or U12709 (N_12709,N_12123,N_12104);
xor U12710 (N_12710,N_12308,N_12453);
and U12711 (N_12711,N_12061,N_12373);
or U12712 (N_12712,N_12439,N_12039);
xor U12713 (N_12713,N_12253,N_12112);
or U12714 (N_12714,N_12249,N_12458);
nand U12715 (N_12715,N_12352,N_12124);
and U12716 (N_12716,N_12435,N_12069);
nor U12717 (N_12717,N_12214,N_12231);
or U12718 (N_12718,N_12053,N_12476);
xor U12719 (N_12719,N_12478,N_12158);
xor U12720 (N_12720,N_12465,N_12473);
and U12721 (N_12721,N_12304,N_12408);
nor U12722 (N_12722,N_12449,N_12357);
nor U12723 (N_12723,N_12337,N_12277);
nand U12724 (N_12724,N_12315,N_12165);
nor U12725 (N_12725,N_12321,N_12320);
and U12726 (N_12726,N_12356,N_12296);
nand U12727 (N_12727,N_12048,N_12013);
nand U12728 (N_12728,N_12378,N_12127);
and U12729 (N_12729,N_12183,N_12419);
and U12730 (N_12730,N_12354,N_12403);
and U12731 (N_12731,N_12350,N_12429);
nand U12732 (N_12732,N_12423,N_12270);
nor U12733 (N_12733,N_12282,N_12358);
and U12734 (N_12734,N_12316,N_12456);
nor U12735 (N_12735,N_12109,N_12445);
nor U12736 (N_12736,N_12206,N_12427);
nand U12737 (N_12737,N_12154,N_12407);
or U12738 (N_12738,N_12491,N_12272);
xor U12739 (N_12739,N_12024,N_12050);
nand U12740 (N_12740,N_12101,N_12300);
or U12741 (N_12741,N_12201,N_12381);
xnor U12742 (N_12742,N_12467,N_12187);
nand U12743 (N_12743,N_12098,N_12279);
and U12744 (N_12744,N_12370,N_12470);
and U12745 (N_12745,N_12235,N_12168);
nand U12746 (N_12746,N_12436,N_12047);
nand U12747 (N_12747,N_12173,N_12153);
xor U12748 (N_12748,N_12274,N_12266);
xnor U12749 (N_12749,N_12142,N_12078);
xnor U12750 (N_12750,N_12163,N_12074);
nand U12751 (N_12751,N_12404,N_12402);
or U12752 (N_12752,N_12497,N_12444);
xnor U12753 (N_12753,N_12268,N_12423);
nor U12754 (N_12754,N_12271,N_12329);
xor U12755 (N_12755,N_12201,N_12258);
and U12756 (N_12756,N_12488,N_12099);
and U12757 (N_12757,N_12095,N_12137);
or U12758 (N_12758,N_12391,N_12333);
nand U12759 (N_12759,N_12157,N_12239);
and U12760 (N_12760,N_12015,N_12429);
xor U12761 (N_12761,N_12162,N_12194);
nand U12762 (N_12762,N_12479,N_12397);
nor U12763 (N_12763,N_12389,N_12186);
and U12764 (N_12764,N_12222,N_12019);
xor U12765 (N_12765,N_12361,N_12125);
xor U12766 (N_12766,N_12173,N_12411);
nor U12767 (N_12767,N_12191,N_12032);
nor U12768 (N_12768,N_12270,N_12477);
and U12769 (N_12769,N_12142,N_12174);
or U12770 (N_12770,N_12092,N_12303);
xnor U12771 (N_12771,N_12153,N_12203);
or U12772 (N_12772,N_12187,N_12200);
or U12773 (N_12773,N_12132,N_12106);
nand U12774 (N_12774,N_12041,N_12262);
or U12775 (N_12775,N_12174,N_12167);
nand U12776 (N_12776,N_12255,N_12069);
nand U12777 (N_12777,N_12219,N_12092);
or U12778 (N_12778,N_12062,N_12070);
or U12779 (N_12779,N_12393,N_12110);
xnor U12780 (N_12780,N_12425,N_12313);
or U12781 (N_12781,N_12025,N_12311);
and U12782 (N_12782,N_12356,N_12246);
nor U12783 (N_12783,N_12338,N_12394);
or U12784 (N_12784,N_12006,N_12169);
nor U12785 (N_12785,N_12112,N_12454);
or U12786 (N_12786,N_12094,N_12114);
nor U12787 (N_12787,N_12371,N_12244);
xor U12788 (N_12788,N_12383,N_12204);
nor U12789 (N_12789,N_12015,N_12306);
nand U12790 (N_12790,N_12335,N_12058);
nor U12791 (N_12791,N_12406,N_12241);
nor U12792 (N_12792,N_12065,N_12147);
nand U12793 (N_12793,N_12358,N_12126);
nor U12794 (N_12794,N_12322,N_12036);
and U12795 (N_12795,N_12204,N_12372);
or U12796 (N_12796,N_12103,N_12462);
nand U12797 (N_12797,N_12351,N_12040);
or U12798 (N_12798,N_12349,N_12187);
nor U12799 (N_12799,N_12043,N_12267);
and U12800 (N_12800,N_12313,N_12261);
and U12801 (N_12801,N_12038,N_12148);
xor U12802 (N_12802,N_12242,N_12013);
xor U12803 (N_12803,N_12165,N_12296);
nor U12804 (N_12804,N_12153,N_12329);
xor U12805 (N_12805,N_12130,N_12099);
and U12806 (N_12806,N_12245,N_12209);
and U12807 (N_12807,N_12021,N_12060);
and U12808 (N_12808,N_12292,N_12306);
nand U12809 (N_12809,N_12217,N_12119);
xor U12810 (N_12810,N_12294,N_12165);
or U12811 (N_12811,N_12431,N_12343);
nand U12812 (N_12812,N_12105,N_12451);
and U12813 (N_12813,N_12160,N_12225);
nor U12814 (N_12814,N_12207,N_12064);
and U12815 (N_12815,N_12347,N_12208);
nand U12816 (N_12816,N_12366,N_12497);
and U12817 (N_12817,N_12315,N_12144);
nand U12818 (N_12818,N_12335,N_12087);
xnor U12819 (N_12819,N_12492,N_12085);
nand U12820 (N_12820,N_12220,N_12169);
nand U12821 (N_12821,N_12006,N_12436);
and U12822 (N_12822,N_12181,N_12380);
nand U12823 (N_12823,N_12263,N_12448);
or U12824 (N_12824,N_12124,N_12152);
xor U12825 (N_12825,N_12362,N_12089);
nand U12826 (N_12826,N_12023,N_12381);
or U12827 (N_12827,N_12179,N_12230);
and U12828 (N_12828,N_12088,N_12162);
and U12829 (N_12829,N_12143,N_12022);
or U12830 (N_12830,N_12234,N_12191);
xor U12831 (N_12831,N_12154,N_12094);
xnor U12832 (N_12832,N_12010,N_12275);
and U12833 (N_12833,N_12066,N_12191);
and U12834 (N_12834,N_12058,N_12065);
nor U12835 (N_12835,N_12022,N_12258);
xor U12836 (N_12836,N_12167,N_12451);
or U12837 (N_12837,N_12221,N_12375);
or U12838 (N_12838,N_12292,N_12091);
or U12839 (N_12839,N_12425,N_12456);
nor U12840 (N_12840,N_12326,N_12280);
xor U12841 (N_12841,N_12197,N_12223);
and U12842 (N_12842,N_12249,N_12497);
nand U12843 (N_12843,N_12374,N_12480);
nand U12844 (N_12844,N_12479,N_12069);
nor U12845 (N_12845,N_12290,N_12172);
nand U12846 (N_12846,N_12366,N_12228);
nand U12847 (N_12847,N_12458,N_12159);
and U12848 (N_12848,N_12084,N_12241);
or U12849 (N_12849,N_12419,N_12116);
nor U12850 (N_12850,N_12402,N_12300);
nor U12851 (N_12851,N_12173,N_12167);
nor U12852 (N_12852,N_12000,N_12164);
nor U12853 (N_12853,N_12226,N_12461);
nor U12854 (N_12854,N_12223,N_12399);
xnor U12855 (N_12855,N_12180,N_12298);
and U12856 (N_12856,N_12043,N_12261);
xnor U12857 (N_12857,N_12329,N_12266);
nor U12858 (N_12858,N_12376,N_12315);
and U12859 (N_12859,N_12258,N_12449);
nor U12860 (N_12860,N_12204,N_12162);
and U12861 (N_12861,N_12090,N_12040);
nand U12862 (N_12862,N_12348,N_12498);
xor U12863 (N_12863,N_12271,N_12289);
nand U12864 (N_12864,N_12008,N_12272);
nand U12865 (N_12865,N_12030,N_12340);
and U12866 (N_12866,N_12234,N_12339);
nand U12867 (N_12867,N_12198,N_12216);
nor U12868 (N_12868,N_12049,N_12017);
xnor U12869 (N_12869,N_12020,N_12311);
or U12870 (N_12870,N_12065,N_12107);
or U12871 (N_12871,N_12170,N_12338);
nand U12872 (N_12872,N_12433,N_12103);
and U12873 (N_12873,N_12420,N_12339);
xor U12874 (N_12874,N_12156,N_12458);
nand U12875 (N_12875,N_12454,N_12120);
nor U12876 (N_12876,N_12341,N_12192);
nand U12877 (N_12877,N_12190,N_12088);
xor U12878 (N_12878,N_12390,N_12315);
or U12879 (N_12879,N_12008,N_12225);
nand U12880 (N_12880,N_12284,N_12002);
nor U12881 (N_12881,N_12227,N_12343);
and U12882 (N_12882,N_12339,N_12392);
nor U12883 (N_12883,N_12148,N_12130);
nand U12884 (N_12884,N_12128,N_12328);
nand U12885 (N_12885,N_12484,N_12010);
or U12886 (N_12886,N_12255,N_12404);
xnor U12887 (N_12887,N_12218,N_12145);
and U12888 (N_12888,N_12445,N_12208);
nand U12889 (N_12889,N_12133,N_12060);
nor U12890 (N_12890,N_12455,N_12480);
or U12891 (N_12891,N_12102,N_12233);
or U12892 (N_12892,N_12133,N_12048);
and U12893 (N_12893,N_12453,N_12374);
nand U12894 (N_12894,N_12452,N_12378);
nand U12895 (N_12895,N_12033,N_12189);
nand U12896 (N_12896,N_12188,N_12048);
nor U12897 (N_12897,N_12203,N_12116);
xor U12898 (N_12898,N_12219,N_12462);
or U12899 (N_12899,N_12399,N_12038);
xor U12900 (N_12900,N_12184,N_12366);
nand U12901 (N_12901,N_12350,N_12259);
nand U12902 (N_12902,N_12315,N_12302);
nand U12903 (N_12903,N_12025,N_12043);
nor U12904 (N_12904,N_12298,N_12318);
or U12905 (N_12905,N_12182,N_12175);
nand U12906 (N_12906,N_12307,N_12344);
nor U12907 (N_12907,N_12450,N_12170);
xnor U12908 (N_12908,N_12090,N_12336);
and U12909 (N_12909,N_12433,N_12443);
nor U12910 (N_12910,N_12112,N_12147);
xnor U12911 (N_12911,N_12416,N_12132);
nand U12912 (N_12912,N_12464,N_12416);
nand U12913 (N_12913,N_12349,N_12439);
xnor U12914 (N_12914,N_12232,N_12164);
nor U12915 (N_12915,N_12175,N_12212);
and U12916 (N_12916,N_12484,N_12224);
and U12917 (N_12917,N_12132,N_12366);
nand U12918 (N_12918,N_12028,N_12176);
or U12919 (N_12919,N_12399,N_12447);
nand U12920 (N_12920,N_12283,N_12415);
and U12921 (N_12921,N_12081,N_12469);
and U12922 (N_12922,N_12264,N_12343);
xor U12923 (N_12923,N_12440,N_12027);
nand U12924 (N_12924,N_12188,N_12115);
or U12925 (N_12925,N_12154,N_12217);
nor U12926 (N_12926,N_12367,N_12289);
nor U12927 (N_12927,N_12391,N_12117);
and U12928 (N_12928,N_12218,N_12158);
or U12929 (N_12929,N_12295,N_12309);
and U12930 (N_12930,N_12470,N_12342);
xnor U12931 (N_12931,N_12130,N_12318);
or U12932 (N_12932,N_12497,N_12479);
nor U12933 (N_12933,N_12272,N_12002);
or U12934 (N_12934,N_12018,N_12257);
xor U12935 (N_12935,N_12254,N_12394);
nand U12936 (N_12936,N_12456,N_12325);
nand U12937 (N_12937,N_12166,N_12371);
and U12938 (N_12938,N_12266,N_12276);
xor U12939 (N_12939,N_12438,N_12037);
xor U12940 (N_12940,N_12120,N_12409);
xnor U12941 (N_12941,N_12007,N_12429);
xnor U12942 (N_12942,N_12121,N_12053);
and U12943 (N_12943,N_12281,N_12213);
nor U12944 (N_12944,N_12356,N_12455);
xor U12945 (N_12945,N_12256,N_12228);
nor U12946 (N_12946,N_12048,N_12385);
and U12947 (N_12947,N_12397,N_12332);
and U12948 (N_12948,N_12028,N_12148);
and U12949 (N_12949,N_12113,N_12265);
or U12950 (N_12950,N_12036,N_12038);
or U12951 (N_12951,N_12307,N_12094);
nor U12952 (N_12952,N_12274,N_12016);
xor U12953 (N_12953,N_12438,N_12177);
or U12954 (N_12954,N_12138,N_12182);
and U12955 (N_12955,N_12364,N_12324);
xnor U12956 (N_12956,N_12451,N_12229);
xor U12957 (N_12957,N_12028,N_12205);
and U12958 (N_12958,N_12228,N_12012);
and U12959 (N_12959,N_12277,N_12494);
xor U12960 (N_12960,N_12046,N_12214);
and U12961 (N_12961,N_12280,N_12123);
xnor U12962 (N_12962,N_12079,N_12351);
xnor U12963 (N_12963,N_12042,N_12440);
xor U12964 (N_12964,N_12175,N_12317);
or U12965 (N_12965,N_12483,N_12463);
nand U12966 (N_12966,N_12491,N_12342);
nor U12967 (N_12967,N_12366,N_12180);
and U12968 (N_12968,N_12225,N_12461);
and U12969 (N_12969,N_12461,N_12126);
nor U12970 (N_12970,N_12381,N_12194);
xor U12971 (N_12971,N_12375,N_12423);
nor U12972 (N_12972,N_12492,N_12008);
or U12973 (N_12973,N_12301,N_12001);
and U12974 (N_12974,N_12164,N_12404);
nor U12975 (N_12975,N_12448,N_12072);
nor U12976 (N_12976,N_12325,N_12043);
nand U12977 (N_12977,N_12077,N_12361);
or U12978 (N_12978,N_12425,N_12180);
nor U12979 (N_12979,N_12338,N_12233);
nor U12980 (N_12980,N_12156,N_12321);
nor U12981 (N_12981,N_12335,N_12153);
or U12982 (N_12982,N_12437,N_12304);
or U12983 (N_12983,N_12048,N_12452);
nor U12984 (N_12984,N_12199,N_12402);
nand U12985 (N_12985,N_12022,N_12279);
nand U12986 (N_12986,N_12266,N_12252);
nor U12987 (N_12987,N_12317,N_12359);
nand U12988 (N_12988,N_12419,N_12404);
xnor U12989 (N_12989,N_12339,N_12229);
xnor U12990 (N_12990,N_12080,N_12362);
xor U12991 (N_12991,N_12312,N_12335);
and U12992 (N_12992,N_12106,N_12141);
nor U12993 (N_12993,N_12359,N_12100);
xor U12994 (N_12994,N_12141,N_12448);
xnor U12995 (N_12995,N_12071,N_12484);
xor U12996 (N_12996,N_12460,N_12350);
nor U12997 (N_12997,N_12283,N_12153);
xor U12998 (N_12998,N_12164,N_12137);
xor U12999 (N_12999,N_12351,N_12489);
and U13000 (N_13000,N_12556,N_12674);
nor U13001 (N_13001,N_12789,N_12708);
xnor U13002 (N_13002,N_12885,N_12914);
nand U13003 (N_13003,N_12593,N_12687);
nor U13004 (N_13004,N_12703,N_12867);
and U13005 (N_13005,N_12531,N_12505);
xor U13006 (N_13006,N_12742,N_12938);
xnor U13007 (N_13007,N_12562,N_12633);
and U13008 (N_13008,N_12585,N_12754);
nand U13009 (N_13009,N_12875,N_12548);
xnor U13010 (N_13010,N_12950,N_12800);
nor U13011 (N_13011,N_12646,N_12919);
or U13012 (N_13012,N_12732,N_12823);
nand U13013 (N_13013,N_12888,N_12761);
nand U13014 (N_13014,N_12921,N_12734);
or U13015 (N_13015,N_12821,N_12838);
nand U13016 (N_13016,N_12760,N_12649);
and U13017 (N_13017,N_12765,N_12965);
nor U13018 (N_13018,N_12715,N_12663);
nor U13019 (N_13019,N_12995,N_12806);
or U13020 (N_13020,N_12826,N_12700);
xor U13021 (N_13021,N_12757,N_12711);
or U13022 (N_13022,N_12980,N_12985);
xnor U13023 (N_13023,N_12746,N_12520);
and U13024 (N_13024,N_12818,N_12848);
nor U13025 (N_13025,N_12790,N_12598);
xor U13026 (N_13026,N_12584,N_12986);
or U13027 (N_13027,N_12517,N_12990);
nand U13028 (N_13028,N_12903,N_12882);
xor U13029 (N_13029,N_12526,N_12997);
and U13030 (N_13030,N_12946,N_12728);
xor U13031 (N_13031,N_12747,N_12776);
and U13032 (N_13032,N_12753,N_12830);
xor U13033 (N_13033,N_12600,N_12840);
nor U13034 (N_13034,N_12973,N_12905);
xor U13035 (N_13035,N_12661,N_12886);
and U13036 (N_13036,N_12542,N_12952);
xnor U13037 (N_13037,N_12524,N_12538);
nor U13038 (N_13038,N_12589,N_12725);
nand U13039 (N_13039,N_12603,N_12942);
nor U13040 (N_13040,N_12839,N_12588);
or U13041 (N_13041,N_12567,N_12772);
and U13042 (N_13042,N_12714,N_12522);
nor U13043 (N_13043,N_12723,N_12509);
nand U13044 (N_13044,N_12716,N_12632);
nor U13045 (N_13045,N_12890,N_12666);
nor U13046 (N_13046,N_12933,N_12705);
and U13047 (N_13047,N_12853,N_12927);
nand U13048 (N_13048,N_12893,N_12523);
or U13049 (N_13049,N_12576,N_12819);
xnor U13050 (N_13050,N_12546,N_12645);
nand U13051 (N_13051,N_12974,N_12502);
nand U13052 (N_13052,N_12932,N_12648);
nor U13053 (N_13053,N_12563,N_12699);
or U13054 (N_13054,N_12810,N_12999);
nor U13055 (N_13055,N_12501,N_12808);
nand U13056 (N_13056,N_12577,N_12904);
nor U13057 (N_13057,N_12718,N_12590);
and U13058 (N_13058,N_12907,N_12792);
nand U13059 (N_13059,N_12749,N_12849);
nor U13060 (N_13060,N_12887,N_12779);
nor U13061 (N_13061,N_12583,N_12636);
and U13062 (N_13062,N_12560,N_12845);
and U13063 (N_13063,N_12870,N_12665);
nor U13064 (N_13064,N_12602,N_12630);
xnor U13065 (N_13065,N_12994,N_12565);
or U13066 (N_13066,N_12859,N_12802);
xnor U13067 (N_13067,N_12568,N_12924);
or U13068 (N_13068,N_12506,N_12956);
or U13069 (N_13069,N_12631,N_12861);
and U13070 (N_13070,N_12774,N_12569);
nor U13071 (N_13071,N_12514,N_12820);
nand U13072 (N_13072,N_12692,N_12672);
nand U13073 (N_13073,N_12954,N_12969);
xnor U13074 (N_13074,N_12793,N_12940);
nor U13075 (N_13075,N_12587,N_12616);
nor U13076 (N_13076,N_12755,N_12635);
and U13077 (N_13077,N_12815,N_12525);
and U13078 (N_13078,N_12876,N_12656);
nor U13079 (N_13079,N_12756,N_12551);
xor U13080 (N_13080,N_12738,N_12961);
and U13081 (N_13081,N_12669,N_12963);
xnor U13082 (N_13082,N_12834,N_12691);
nand U13083 (N_13083,N_12968,N_12827);
and U13084 (N_13084,N_12978,N_12706);
xnor U13085 (N_13085,N_12537,N_12682);
xor U13086 (N_13086,N_12628,N_12564);
nand U13087 (N_13087,N_12852,N_12773);
or U13088 (N_13088,N_12922,N_12608);
nor U13089 (N_13089,N_12730,N_12982);
nor U13090 (N_13090,N_12724,N_12557);
nand U13091 (N_13091,N_12652,N_12580);
nor U13092 (N_13092,N_12612,N_12984);
xnor U13093 (N_13093,N_12987,N_12533);
or U13094 (N_13094,N_12529,N_12637);
or U13095 (N_13095,N_12784,N_12979);
and U13096 (N_13096,N_12872,N_12856);
xor U13097 (N_13097,N_12944,N_12873);
and U13098 (N_13098,N_12748,N_12750);
xnor U13099 (N_13099,N_12998,N_12909);
or U13100 (N_13100,N_12855,N_12770);
and U13101 (N_13101,N_12515,N_12640);
nor U13102 (N_13102,N_12841,N_12739);
nor U13103 (N_13103,N_12992,N_12528);
or U13104 (N_13104,N_12673,N_12555);
and U13105 (N_13105,N_12504,N_12759);
xor U13106 (N_13106,N_12601,N_12824);
nor U13107 (N_13107,N_12783,N_12731);
nor U13108 (N_13108,N_12615,N_12953);
nor U13109 (N_13109,N_12625,N_12662);
nor U13110 (N_13110,N_12923,N_12720);
or U13111 (N_13111,N_12785,N_12690);
nor U13112 (N_13112,N_12717,N_12975);
nor U13113 (N_13113,N_12653,N_12599);
xor U13114 (N_13114,N_12667,N_12796);
nor U13115 (N_13115,N_12655,N_12654);
nor U13116 (N_13116,N_12527,N_12816);
or U13117 (N_13117,N_12573,N_12850);
nand U13118 (N_13118,N_12983,N_12684);
and U13119 (N_13119,N_12869,N_12534);
or U13120 (N_13120,N_12741,N_12912);
or U13121 (N_13121,N_12622,N_12668);
nand U13122 (N_13122,N_12908,N_12638);
xnor U13123 (N_13123,N_12879,N_12833);
nor U13124 (N_13124,N_12670,N_12752);
xor U13125 (N_13125,N_12920,N_12695);
nor U13126 (N_13126,N_12782,N_12701);
nand U13127 (N_13127,N_12581,N_12541);
nand U13128 (N_13128,N_12617,N_12543);
or U13129 (N_13129,N_12644,N_12518);
xor U13130 (N_13130,N_12710,N_12618);
xor U13131 (N_13131,N_12712,N_12647);
nor U13132 (N_13132,N_12610,N_12574);
or U13133 (N_13133,N_12843,N_12788);
or U13134 (N_13134,N_12733,N_12928);
nor U13135 (N_13135,N_12934,N_12916);
nor U13136 (N_13136,N_12609,N_12906);
and U13137 (N_13137,N_12771,N_12804);
xor U13138 (N_13138,N_12862,N_12595);
xnor U13139 (N_13139,N_12769,N_12685);
or U13140 (N_13140,N_12596,N_12678);
nor U13141 (N_13141,N_12947,N_12591);
nor U13142 (N_13142,N_12763,N_12516);
or U13143 (N_13143,N_12863,N_12901);
nor U13144 (N_13144,N_12897,N_12726);
nor U13145 (N_13145,N_12878,N_12858);
or U13146 (N_13146,N_12619,N_12935);
and U13147 (N_13147,N_12536,N_12766);
xor U13148 (N_13148,N_12606,N_12689);
and U13149 (N_13149,N_12966,N_12884);
or U13150 (N_13150,N_12896,N_12962);
nand U13151 (N_13151,N_12677,N_12799);
or U13152 (N_13152,N_12570,N_12623);
and U13153 (N_13153,N_12707,N_12851);
or U13154 (N_13154,N_12605,N_12604);
and U13155 (N_13155,N_12686,N_12976);
xor U13156 (N_13156,N_12795,N_12698);
or U13157 (N_13157,N_12807,N_12917);
or U13158 (N_13158,N_12949,N_12650);
nand U13159 (N_13159,N_12547,N_12575);
and U13160 (N_13160,N_12996,N_12857);
and U13161 (N_13161,N_12696,N_12854);
nand U13162 (N_13162,N_12989,N_12688);
or U13163 (N_13163,N_12880,N_12778);
or U13164 (N_13164,N_12825,N_12764);
or U13165 (N_13165,N_12803,N_12931);
nor U13166 (N_13166,N_12866,N_12967);
nor U13167 (N_13167,N_12642,N_12891);
or U13168 (N_13168,N_12865,N_12500);
or U13169 (N_13169,N_12831,N_12943);
or U13170 (N_13170,N_12626,N_12736);
or U13171 (N_13171,N_12740,N_12955);
nor U13172 (N_13172,N_12939,N_12822);
nand U13173 (N_13173,N_12925,N_12620);
nand U13174 (N_13174,N_12814,N_12768);
nand U13175 (N_13175,N_12828,N_12964);
xor U13176 (N_13176,N_12704,N_12549);
xor U13177 (N_13177,N_12832,N_12675);
nor U13178 (N_13178,N_12797,N_12639);
nand U13179 (N_13179,N_12809,N_12767);
xnor U13180 (N_13180,N_12643,N_12683);
or U13181 (N_13181,N_12558,N_12892);
or U13182 (N_13182,N_12864,N_12657);
nor U13183 (N_13183,N_12811,N_12829);
nand U13184 (N_13184,N_12787,N_12532);
or U13185 (N_13185,N_12729,N_12721);
or U13186 (N_13186,N_12958,N_12511);
nor U13187 (N_13187,N_12813,N_12614);
xor U13188 (N_13188,N_12936,N_12737);
or U13189 (N_13189,N_12719,N_12895);
or U13190 (N_13190,N_12970,N_12868);
and U13191 (N_13191,N_12911,N_12988);
and U13192 (N_13192,N_12572,N_12981);
nor U13193 (N_13193,N_12521,N_12930);
xor U13194 (N_13194,N_12693,N_12812);
and U13195 (N_13195,N_12874,N_12578);
nor U13196 (N_13196,N_12743,N_12805);
nor U13197 (N_13197,N_12842,N_12713);
nand U13198 (N_13198,N_12679,N_12641);
and U13199 (N_13199,N_12651,N_12910);
xor U13200 (N_13200,N_12539,N_12889);
or U13201 (N_13201,N_12676,N_12775);
or U13202 (N_13202,N_12535,N_12550);
xor U13203 (N_13203,N_12624,N_12586);
xor U13204 (N_13204,N_12621,N_12544);
and U13205 (N_13205,N_12709,N_12744);
nor U13206 (N_13206,N_12817,N_12957);
nand U13207 (N_13207,N_12929,N_12745);
and U13208 (N_13208,N_12503,N_12881);
or U13209 (N_13209,N_12900,N_12613);
nor U13210 (N_13210,N_12972,N_12735);
xor U13211 (N_13211,N_12926,N_12960);
and U13212 (N_13212,N_12582,N_12915);
nand U13213 (N_13213,N_12993,N_12545);
or U13214 (N_13214,N_12781,N_12634);
nor U13215 (N_13215,N_12727,N_12553);
nor U13216 (N_13216,N_12627,N_12566);
xor U13217 (N_13217,N_12918,N_12561);
or U13218 (N_13218,N_12894,N_12951);
xnor U13219 (N_13219,N_12552,N_12844);
or U13220 (N_13220,N_12507,N_12877);
or U13221 (N_13221,N_12945,N_12579);
or U13222 (N_13222,N_12780,N_12694);
xor U13223 (N_13223,N_12702,N_12659);
or U13224 (N_13224,N_12899,N_12941);
nand U13225 (N_13225,N_12571,N_12883);
and U13226 (N_13226,N_12629,N_12937);
nor U13227 (N_13227,N_12871,N_12837);
and U13228 (N_13228,N_12898,N_12836);
or U13229 (N_13229,N_12971,N_12794);
or U13230 (N_13230,N_12559,N_12510);
and U13231 (N_13231,N_12959,N_12835);
nand U13232 (N_13232,N_12597,N_12751);
or U13233 (N_13233,N_12611,N_12948);
xnor U13234 (N_13234,N_12681,N_12664);
and U13235 (N_13235,N_12658,N_12594);
xnor U13236 (N_13236,N_12860,N_12791);
nor U13237 (N_13237,N_12512,N_12991);
and U13238 (N_13238,N_12697,N_12913);
nor U13239 (N_13239,N_12540,N_12902);
and U13240 (N_13240,N_12977,N_12762);
xnor U13241 (N_13241,N_12592,N_12847);
nand U13242 (N_13242,N_12680,N_12513);
or U13243 (N_13243,N_12519,N_12777);
nor U13244 (N_13244,N_12798,N_12607);
nand U13245 (N_13245,N_12530,N_12554);
xnor U13246 (N_13246,N_12846,N_12786);
nor U13247 (N_13247,N_12508,N_12722);
nor U13248 (N_13248,N_12660,N_12671);
and U13249 (N_13249,N_12801,N_12758);
or U13250 (N_13250,N_12972,N_12706);
xnor U13251 (N_13251,N_12905,N_12957);
and U13252 (N_13252,N_12934,N_12942);
nand U13253 (N_13253,N_12504,N_12902);
or U13254 (N_13254,N_12822,N_12630);
xnor U13255 (N_13255,N_12531,N_12752);
xor U13256 (N_13256,N_12809,N_12599);
nor U13257 (N_13257,N_12623,N_12991);
xor U13258 (N_13258,N_12912,N_12708);
xnor U13259 (N_13259,N_12987,N_12720);
nand U13260 (N_13260,N_12784,N_12990);
nand U13261 (N_13261,N_12850,N_12780);
nand U13262 (N_13262,N_12734,N_12646);
nand U13263 (N_13263,N_12633,N_12621);
and U13264 (N_13264,N_12757,N_12518);
xnor U13265 (N_13265,N_12743,N_12911);
or U13266 (N_13266,N_12983,N_12789);
xor U13267 (N_13267,N_12828,N_12840);
nor U13268 (N_13268,N_12636,N_12650);
or U13269 (N_13269,N_12950,N_12678);
and U13270 (N_13270,N_12835,N_12518);
xor U13271 (N_13271,N_12613,N_12921);
xnor U13272 (N_13272,N_12921,N_12842);
nor U13273 (N_13273,N_12912,N_12647);
xnor U13274 (N_13274,N_12728,N_12590);
nand U13275 (N_13275,N_12983,N_12718);
nand U13276 (N_13276,N_12657,N_12655);
xor U13277 (N_13277,N_12810,N_12556);
or U13278 (N_13278,N_12785,N_12676);
xor U13279 (N_13279,N_12612,N_12577);
and U13280 (N_13280,N_12700,N_12647);
and U13281 (N_13281,N_12782,N_12558);
nor U13282 (N_13282,N_12841,N_12582);
nand U13283 (N_13283,N_12771,N_12637);
nand U13284 (N_13284,N_12895,N_12671);
nand U13285 (N_13285,N_12591,N_12690);
nand U13286 (N_13286,N_12711,N_12644);
nor U13287 (N_13287,N_12932,N_12755);
nor U13288 (N_13288,N_12745,N_12756);
and U13289 (N_13289,N_12987,N_12912);
nand U13290 (N_13290,N_12785,N_12840);
nand U13291 (N_13291,N_12601,N_12874);
nand U13292 (N_13292,N_12857,N_12657);
xor U13293 (N_13293,N_12597,N_12548);
xnor U13294 (N_13294,N_12533,N_12926);
and U13295 (N_13295,N_12561,N_12593);
nand U13296 (N_13296,N_12737,N_12605);
xnor U13297 (N_13297,N_12548,N_12833);
nand U13298 (N_13298,N_12736,N_12853);
xor U13299 (N_13299,N_12749,N_12641);
nor U13300 (N_13300,N_12538,N_12922);
and U13301 (N_13301,N_12951,N_12736);
and U13302 (N_13302,N_12789,N_12971);
and U13303 (N_13303,N_12979,N_12583);
nand U13304 (N_13304,N_12986,N_12771);
xor U13305 (N_13305,N_12859,N_12651);
xnor U13306 (N_13306,N_12836,N_12686);
xor U13307 (N_13307,N_12634,N_12768);
nor U13308 (N_13308,N_12534,N_12690);
or U13309 (N_13309,N_12894,N_12676);
nor U13310 (N_13310,N_12529,N_12965);
or U13311 (N_13311,N_12511,N_12986);
nor U13312 (N_13312,N_12655,N_12630);
nor U13313 (N_13313,N_12770,N_12648);
nand U13314 (N_13314,N_12747,N_12655);
and U13315 (N_13315,N_12870,N_12720);
xor U13316 (N_13316,N_12515,N_12902);
or U13317 (N_13317,N_12705,N_12641);
xor U13318 (N_13318,N_12867,N_12522);
or U13319 (N_13319,N_12569,N_12897);
nand U13320 (N_13320,N_12930,N_12953);
xor U13321 (N_13321,N_12685,N_12773);
nand U13322 (N_13322,N_12592,N_12981);
xnor U13323 (N_13323,N_12507,N_12651);
xnor U13324 (N_13324,N_12670,N_12572);
nand U13325 (N_13325,N_12708,N_12791);
nor U13326 (N_13326,N_12671,N_12975);
and U13327 (N_13327,N_12565,N_12956);
or U13328 (N_13328,N_12648,N_12647);
or U13329 (N_13329,N_12546,N_12856);
nor U13330 (N_13330,N_12666,N_12879);
xnor U13331 (N_13331,N_12838,N_12945);
nor U13332 (N_13332,N_12905,N_12761);
and U13333 (N_13333,N_12888,N_12900);
and U13334 (N_13334,N_12740,N_12668);
nand U13335 (N_13335,N_12651,N_12972);
or U13336 (N_13336,N_12933,N_12980);
and U13337 (N_13337,N_12758,N_12648);
nand U13338 (N_13338,N_12966,N_12874);
nand U13339 (N_13339,N_12952,N_12895);
and U13340 (N_13340,N_12521,N_12632);
nor U13341 (N_13341,N_12681,N_12849);
xnor U13342 (N_13342,N_12825,N_12812);
nor U13343 (N_13343,N_12678,N_12734);
or U13344 (N_13344,N_12770,N_12879);
nor U13345 (N_13345,N_12883,N_12933);
nand U13346 (N_13346,N_12820,N_12936);
nor U13347 (N_13347,N_12706,N_12814);
nand U13348 (N_13348,N_12532,N_12529);
or U13349 (N_13349,N_12523,N_12920);
or U13350 (N_13350,N_12688,N_12766);
or U13351 (N_13351,N_12839,N_12736);
or U13352 (N_13352,N_12618,N_12879);
nor U13353 (N_13353,N_12631,N_12862);
or U13354 (N_13354,N_12575,N_12720);
and U13355 (N_13355,N_12573,N_12538);
xor U13356 (N_13356,N_12601,N_12644);
or U13357 (N_13357,N_12882,N_12526);
and U13358 (N_13358,N_12802,N_12704);
nor U13359 (N_13359,N_12839,N_12648);
xor U13360 (N_13360,N_12849,N_12619);
or U13361 (N_13361,N_12880,N_12609);
xnor U13362 (N_13362,N_12888,N_12876);
nand U13363 (N_13363,N_12799,N_12526);
nor U13364 (N_13364,N_12855,N_12557);
or U13365 (N_13365,N_12872,N_12888);
or U13366 (N_13366,N_12955,N_12884);
and U13367 (N_13367,N_12506,N_12561);
nor U13368 (N_13368,N_12756,N_12785);
and U13369 (N_13369,N_12661,N_12711);
and U13370 (N_13370,N_12972,N_12787);
nand U13371 (N_13371,N_12552,N_12575);
nor U13372 (N_13372,N_12771,N_12590);
and U13373 (N_13373,N_12628,N_12516);
and U13374 (N_13374,N_12890,N_12687);
nor U13375 (N_13375,N_12671,N_12585);
xnor U13376 (N_13376,N_12614,N_12948);
xnor U13377 (N_13377,N_12650,N_12697);
nand U13378 (N_13378,N_12740,N_12962);
and U13379 (N_13379,N_12578,N_12685);
xnor U13380 (N_13380,N_12778,N_12529);
nor U13381 (N_13381,N_12812,N_12666);
and U13382 (N_13382,N_12949,N_12940);
and U13383 (N_13383,N_12860,N_12622);
nand U13384 (N_13384,N_12916,N_12929);
or U13385 (N_13385,N_12602,N_12838);
nand U13386 (N_13386,N_12888,N_12865);
and U13387 (N_13387,N_12718,N_12777);
nand U13388 (N_13388,N_12700,N_12990);
xnor U13389 (N_13389,N_12514,N_12528);
or U13390 (N_13390,N_12671,N_12930);
nor U13391 (N_13391,N_12536,N_12751);
nor U13392 (N_13392,N_12711,N_12944);
nand U13393 (N_13393,N_12590,N_12925);
nand U13394 (N_13394,N_12988,N_12599);
xnor U13395 (N_13395,N_12872,N_12806);
nor U13396 (N_13396,N_12652,N_12583);
xor U13397 (N_13397,N_12563,N_12767);
or U13398 (N_13398,N_12973,N_12992);
and U13399 (N_13399,N_12922,N_12787);
and U13400 (N_13400,N_12709,N_12575);
or U13401 (N_13401,N_12540,N_12541);
xor U13402 (N_13402,N_12586,N_12606);
nor U13403 (N_13403,N_12612,N_12761);
xor U13404 (N_13404,N_12637,N_12617);
nand U13405 (N_13405,N_12633,N_12567);
xor U13406 (N_13406,N_12985,N_12661);
xor U13407 (N_13407,N_12645,N_12914);
and U13408 (N_13408,N_12896,N_12731);
or U13409 (N_13409,N_12873,N_12975);
xnor U13410 (N_13410,N_12899,N_12597);
xor U13411 (N_13411,N_12921,N_12828);
xor U13412 (N_13412,N_12766,N_12661);
or U13413 (N_13413,N_12914,N_12866);
xor U13414 (N_13414,N_12674,N_12715);
or U13415 (N_13415,N_12953,N_12711);
or U13416 (N_13416,N_12671,N_12715);
nand U13417 (N_13417,N_12590,N_12986);
nand U13418 (N_13418,N_12522,N_12702);
nor U13419 (N_13419,N_12959,N_12518);
or U13420 (N_13420,N_12867,N_12740);
nor U13421 (N_13421,N_12504,N_12664);
or U13422 (N_13422,N_12585,N_12703);
nor U13423 (N_13423,N_12867,N_12722);
or U13424 (N_13424,N_12986,N_12674);
xnor U13425 (N_13425,N_12772,N_12690);
or U13426 (N_13426,N_12520,N_12721);
nand U13427 (N_13427,N_12709,N_12908);
nand U13428 (N_13428,N_12716,N_12908);
nand U13429 (N_13429,N_12778,N_12575);
nor U13430 (N_13430,N_12795,N_12614);
or U13431 (N_13431,N_12971,N_12775);
or U13432 (N_13432,N_12525,N_12858);
and U13433 (N_13433,N_12879,N_12537);
or U13434 (N_13434,N_12530,N_12529);
or U13435 (N_13435,N_12848,N_12815);
and U13436 (N_13436,N_12546,N_12894);
or U13437 (N_13437,N_12746,N_12947);
nand U13438 (N_13438,N_12818,N_12808);
nand U13439 (N_13439,N_12720,N_12867);
xnor U13440 (N_13440,N_12966,N_12659);
nor U13441 (N_13441,N_12684,N_12824);
and U13442 (N_13442,N_12577,N_12984);
nand U13443 (N_13443,N_12902,N_12951);
or U13444 (N_13444,N_12771,N_12889);
and U13445 (N_13445,N_12574,N_12503);
xnor U13446 (N_13446,N_12948,N_12581);
and U13447 (N_13447,N_12791,N_12688);
nor U13448 (N_13448,N_12623,N_12949);
nand U13449 (N_13449,N_12689,N_12854);
nor U13450 (N_13450,N_12721,N_12847);
nor U13451 (N_13451,N_12801,N_12706);
nor U13452 (N_13452,N_12833,N_12930);
nor U13453 (N_13453,N_12913,N_12648);
or U13454 (N_13454,N_12596,N_12919);
or U13455 (N_13455,N_12708,N_12705);
or U13456 (N_13456,N_12981,N_12980);
xnor U13457 (N_13457,N_12703,N_12950);
nor U13458 (N_13458,N_12713,N_12845);
nor U13459 (N_13459,N_12703,N_12740);
nor U13460 (N_13460,N_12773,N_12504);
or U13461 (N_13461,N_12528,N_12878);
nand U13462 (N_13462,N_12703,N_12693);
nor U13463 (N_13463,N_12928,N_12662);
and U13464 (N_13464,N_12848,N_12881);
and U13465 (N_13465,N_12758,N_12875);
nand U13466 (N_13466,N_12539,N_12998);
nand U13467 (N_13467,N_12981,N_12894);
or U13468 (N_13468,N_12850,N_12591);
or U13469 (N_13469,N_12938,N_12880);
nor U13470 (N_13470,N_12868,N_12929);
or U13471 (N_13471,N_12855,N_12730);
nand U13472 (N_13472,N_12834,N_12681);
and U13473 (N_13473,N_12856,N_12616);
xor U13474 (N_13474,N_12586,N_12639);
xor U13475 (N_13475,N_12643,N_12778);
xnor U13476 (N_13476,N_12576,N_12705);
and U13477 (N_13477,N_12769,N_12989);
and U13478 (N_13478,N_12590,N_12824);
nor U13479 (N_13479,N_12653,N_12887);
xor U13480 (N_13480,N_12502,N_12773);
or U13481 (N_13481,N_12553,N_12520);
nor U13482 (N_13482,N_12657,N_12673);
nor U13483 (N_13483,N_12523,N_12790);
nor U13484 (N_13484,N_12979,N_12697);
or U13485 (N_13485,N_12541,N_12914);
or U13486 (N_13486,N_12751,N_12667);
or U13487 (N_13487,N_12866,N_12958);
xnor U13488 (N_13488,N_12543,N_12760);
nand U13489 (N_13489,N_12587,N_12944);
nor U13490 (N_13490,N_12668,N_12938);
xor U13491 (N_13491,N_12727,N_12755);
and U13492 (N_13492,N_12789,N_12993);
nor U13493 (N_13493,N_12738,N_12929);
xor U13494 (N_13494,N_12706,N_12779);
nand U13495 (N_13495,N_12778,N_12939);
or U13496 (N_13496,N_12766,N_12517);
nand U13497 (N_13497,N_12822,N_12882);
nand U13498 (N_13498,N_12721,N_12973);
nor U13499 (N_13499,N_12818,N_12912);
nor U13500 (N_13500,N_13454,N_13306);
nor U13501 (N_13501,N_13399,N_13325);
and U13502 (N_13502,N_13001,N_13056);
nor U13503 (N_13503,N_13096,N_13422);
nand U13504 (N_13504,N_13299,N_13463);
xnor U13505 (N_13505,N_13028,N_13276);
or U13506 (N_13506,N_13457,N_13066);
xnor U13507 (N_13507,N_13054,N_13467);
xnor U13508 (N_13508,N_13197,N_13007);
nor U13509 (N_13509,N_13423,N_13024);
nand U13510 (N_13510,N_13053,N_13067);
and U13511 (N_13511,N_13125,N_13095);
nor U13512 (N_13512,N_13285,N_13492);
or U13513 (N_13513,N_13175,N_13159);
nor U13514 (N_13514,N_13295,N_13397);
nor U13515 (N_13515,N_13392,N_13181);
nand U13516 (N_13516,N_13312,N_13177);
nor U13517 (N_13517,N_13484,N_13390);
or U13518 (N_13518,N_13371,N_13357);
or U13519 (N_13519,N_13241,N_13365);
nor U13520 (N_13520,N_13027,N_13291);
or U13521 (N_13521,N_13078,N_13353);
nor U13522 (N_13522,N_13217,N_13333);
or U13523 (N_13523,N_13219,N_13334);
nand U13524 (N_13524,N_13290,N_13158);
and U13525 (N_13525,N_13267,N_13218);
or U13526 (N_13526,N_13088,N_13465);
or U13527 (N_13527,N_13224,N_13120);
or U13528 (N_13528,N_13081,N_13071);
and U13529 (N_13529,N_13308,N_13037);
xor U13530 (N_13530,N_13242,N_13187);
xnor U13531 (N_13531,N_13494,N_13033);
or U13532 (N_13532,N_13363,N_13246);
xor U13533 (N_13533,N_13212,N_13444);
nand U13534 (N_13534,N_13000,N_13410);
nor U13535 (N_13535,N_13477,N_13336);
nor U13536 (N_13536,N_13247,N_13304);
xor U13537 (N_13537,N_13350,N_13347);
and U13538 (N_13538,N_13155,N_13475);
nand U13539 (N_13539,N_13386,N_13161);
nand U13540 (N_13540,N_13018,N_13442);
xnor U13541 (N_13541,N_13222,N_13493);
nand U13542 (N_13542,N_13145,N_13163);
nor U13543 (N_13543,N_13430,N_13051);
nand U13544 (N_13544,N_13153,N_13164);
or U13545 (N_13545,N_13378,N_13302);
or U13546 (N_13546,N_13329,N_13327);
nor U13547 (N_13547,N_13113,N_13002);
xnor U13548 (N_13548,N_13331,N_13292);
or U13549 (N_13549,N_13394,N_13482);
or U13550 (N_13550,N_13411,N_13045);
or U13551 (N_13551,N_13278,N_13229);
and U13552 (N_13552,N_13006,N_13226);
nor U13553 (N_13553,N_13384,N_13438);
or U13554 (N_13554,N_13070,N_13107);
xor U13555 (N_13555,N_13118,N_13388);
xor U13556 (N_13556,N_13273,N_13449);
nor U13557 (N_13557,N_13473,N_13448);
nor U13558 (N_13558,N_13328,N_13435);
or U13559 (N_13559,N_13244,N_13271);
xor U13560 (N_13560,N_13466,N_13069);
nor U13561 (N_13561,N_13289,N_13373);
and U13562 (N_13562,N_13106,N_13192);
nand U13563 (N_13563,N_13030,N_13205);
nand U13564 (N_13564,N_13134,N_13148);
xor U13565 (N_13565,N_13025,N_13298);
nor U13566 (N_13566,N_13122,N_13166);
nand U13567 (N_13567,N_13049,N_13080);
nor U13568 (N_13568,N_13441,N_13102);
xnor U13569 (N_13569,N_13445,N_13337);
nand U13570 (N_13570,N_13496,N_13468);
and U13571 (N_13571,N_13179,N_13202);
and U13572 (N_13572,N_13180,N_13047);
or U13573 (N_13573,N_13200,N_13446);
nor U13574 (N_13574,N_13128,N_13303);
xnor U13575 (N_13575,N_13479,N_13381);
nand U13576 (N_13576,N_13206,N_13232);
and U13577 (N_13577,N_13287,N_13042);
nand U13578 (N_13578,N_13311,N_13221);
xnor U13579 (N_13579,N_13360,N_13348);
or U13580 (N_13580,N_13048,N_13035);
or U13581 (N_13581,N_13152,N_13238);
or U13582 (N_13582,N_13016,N_13476);
and U13583 (N_13583,N_13346,N_13437);
nor U13584 (N_13584,N_13284,N_13433);
nand U13585 (N_13585,N_13194,N_13117);
and U13586 (N_13586,N_13314,N_13009);
and U13587 (N_13587,N_13352,N_13032);
xor U13588 (N_13588,N_13144,N_13097);
xor U13589 (N_13589,N_13140,N_13379);
xnor U13590 (N_13590,N_13089,N_13338);
or U13591 (N_13591,N_13491,N_13073);
xor U13592 (N_13592,N_13087,N_13021);
xor U13593 (N_13593,N_13447,N_13398);
xnor U13594 (N_13594,N_13077,N_13228);
xnor U13595 (N_13595,N_13204,N_13252);
nor U13596 (N_13596,N_13413,N_13057);
and U13597 (N_13597,N_13227,N_13012);
or U13598 (N_13598,N_13387,N_13074);
nand U13599 (N_13599,N_13110,N_13324);
or U13600 (N_13600,N_13282,N_13436);
or U13601 (N_13601,N_13160,N_13412);
xnor U13602 (N_13602,N_13424,N_13169);
or U13603 (N_13603,N_13198,N_13136);
nand U13604 (N_13604,N_13452,N_13201);
nand U13605 (N_13605,N_13216,N_13139);
xor U13606 (N_13606,N_13039,N_13420);
and U13607 (N_13607,N_13041,N_13429);
nand U13608 (N_13608,N_13450,N_13341);
nor U13609 (N_13609,N_13266,N_13190);
and U13610 (N_13610,N_13279,N_13254);
nand U13611 (N_13611,N_13489,N_13345);
or U13612 (N_13612,N_13320,N_13483);
or U13613 (N_13613,N_13129,N_13258);
and U13614 (N_13614,N_13230,N_13407);
nand U13615 (N_13615,N_13055,N_13093);
nand U13616 (N_13616,N_13130,N_13203);
and U13617 (N_13617,N_13183,N_13419);
nand U13618 (N_13618,N_13374,N_13321);
or U13619 (N_13619,N_13443,N_13355);
nor U13620 (N_13620,N_13456,N_13297);
nor U13621 (N_13621,N_13111,N_13385);
or U13622 (N_13622,N_13309,N_13023);
nor U13623 (N_13623,N_13310,N_13061);
nor U13624 (N_13624,N_13105,N_13370);
and U13625 (N_13625,N_13225,N_13305);
xnor U13626 (N_13626,N_13375,N_13100);
nor U13627 (N_13627,N_13239,N_13235);
xor U13628 (N_13628,N_13060,N_13319);
nor U13629 (N_13629,N_13062,N_13065);
nand U13630 (N_13630,N_13188,N_13135);
and U13631 (N_13631,N_13013,N_13236);
or U13632 (N_13632,N_13059,N_13335);
and U13633 (N_13633,N_13248,N_13277);
and U13634 (N_13634,N_13427,N_13340);
nor U13635 (N_13635,N_13072,N_13004);
xor U13636 (N_13636,N_13404,N_13255);
or U13637 (N_13637,N_13017,N_13418);
and U13638 (N_13638,N_13075,N_13115);
or U13639 (N_13639,N_13498,N_13354);
nand U13640 (N_13640,N_13293,N_13091);
nand U13641 (N_13641,N_13234,N_13112);
xor U13642 (N_13642,N_13326,N_13174);
nand U13643 (N_13643,N_13237,N_13270);
xor U13644 (N_13644,N_13076,N_13036);
or U13645 (N_13645,N_13472,N_13426);
nand U13646 (N_13646,N_13094,N_13401);
and U13647 (N_13647,N_13263,N_13127);
or U13648 (N_13648,N_13461,N_13008);
xor U13649 (N_13649,N_13034,N_13151);
xnor U13650 (N_13650,N_13318,N_13124);
and U13651 (N_13651,N_13356,N_13231);
xor U13652 (N_13652,N_13019,N_13383);
and U13653 (N_13653,N_13275,N_13274);
or U13654 (N_13654,N_13369,N_13020);
and U13655 (N_13655,N_13301,N_13214);
or U13656 (N_13656,N_13090,N_13417);
nor U13657 (N_13657,N_13499,N_13046);
xor U13658 (N_13658,N_13400,N_13063);
or U13659 (N_13659,N_13233,N_13478);
nor U13660 (N_13660,N_13099,N_13439);
nor U13661 (N_13661,N_13487,N_13431);
nor U13662 (N_13662,N_13176,N_13068);
xnor U13663 (N_13663,N_13460,N_13415);
nor U13664 (N_13664,N_13343,N_13349);
xor U13665 (N_13665,N_13167,N_13272);
xor U13666 (N_13666,N_13262,N_13182);
or U13667 (N_13667,N_13215,N_13103);
and U13668 (N_13668,N_13196,N_13126);
nor U13669 (N_13669,N_13114,N_13189);
nor U13670 (N_13670,N_13339,N_13142);
xor U13671 (N_13671,N_13050,N_13014);
nor U13672 (N_13672,N_13086,N_13223);
nor U13673 (N_13673,N_13269,N_13364);
xor U13674 (N_13674,N_13162,N_13405);
nor U13675 (N_13675,N_13141,N_13031);
nor U13676 (N_13676,N_13434,N_13406);
or U13677 (N_13677,N_13245,N_13322);
xor U13678 (N_13678,N_13199,N_13064);
nand U13679 (N_13679,N_13029,N_13119);
nor U13680 (N_13680,N_13083,N_13380);
nor U13681 (N_13681,N_13026,N_13132);
or U13682 (N_13682,N_13010,N_13186);
nor U13683 (N_13683,N_13207,N_13403);
nand U13684 (N_13684,N_13015,N_13358);
nand U13685 (N_13685,N_13082,N_13022);
nor U13686 (N_13686,N_13464,N_13209);
and U13687 (N_13687,N_13300,N_13170);
and U13688 (N_13688,N_13058,N_13391);
xnor U13689 (N_13689,N_13003,N_13480);
xor U13690 (N_13690,N_13313,N_13440);
or U13691 (N_13691,N_13330,N_13372);
and U13692 (N_13692,N_13332,N_13458);
and U13693 (N_13693,N_13286,N_13108);
and U13694 (N_13694,N_13052,N_13432);
and U13695 (N_13695,N_13368,N_13154);
nor U13696 (N_13696,N_13208,N_13395);
nor U13697 (N_13697,N_13408,N_13402);
nor U13698 (N_13698,N_13342,N_13084);
nand U13699 (N_13699,N_13178,N_13143);
xor U13700 (N_13700,N_13495,N_13157);
xnor U13701 (N_13701,N_13146,N_13294);
xor U13702 (N_13702,N_13366,N_13425);
nand U13703 (N_13703,N_13261,N_13085);
xor U13704 (N_13704,N_13362,N_13260);
nand U13705 (N_13705,N_13451,N_13249);
and U13706 (N_13706,N_13121,N_13288);
or U13707 (N_13707,N_13453,N_13389);
or U13708 (N_13708,N_13195,N_13257);
or U13709 (N_13709,N_13101,N_13098);
nand U13710 (N_13710,N_13462,N_13367);
and U13711 (N_13711,N_13210,N_13137);
nor U13712 (N_13712,N_13359,N_13156);
nand U13713 (N_13713,N_13165,N_13393);
or U13714 (N_13714,N_13104,N_13011);
nand U13715 (N_13715,N_13044,N_13109);
and U13716 (N_13716,N_13268,N_13486);
nor U13717 (N_13717,N_13323,N_13043);
and U13718 (N_13718,N_13150,N_13171);
and U13719 (N_13719,N_13079,N_13185);
nand U13720 (N_13720,N_13485,N_13382);
xor U13721 (N_13721,N_13040,N_13471);
nand U13722 (N_13722,N_13168,N_13490);
xnor U13723 (N_13723,N_13184,N_13361);
nor U13724 (N_13724,N_13315,N_13481);
nor U13725 (N_13725,N_13428,N_13488);
or U13726 (N_13726,N_13243,N_13281);
or U13727 (N_13727,N_13421,N_13172);
nor U13728 (N_13728,N_13376,N_13005);
and U13729 (N_13729,N_13149,N_13280);
nor U13730 (N_13730,N_13133,N_13469);
nand U13731 (N_13731,N_13474,N_13251);
xor U13732 (N_13732,N_13193,N_13307);
nor U13733 (N_13733,N_13211,N_13265);
or U13734 (N_13734,N_13253,N_13038);
and U13735 (N_13735,N_13147,N_13259);
nand U13736 (N_13736,N_13416,N_13092);
nor U13737 (N_13737,N_13191,N_13240);
xor U13738 (N_13738,N_13497,N_13409);
and U13739 (N_13739,N_13283,N_13250);
or U13740 (N_13740,N_13316,N_13220);
xnor U13741 (N_13741,N_13470,N_13131);
or U13742 (N_13742,N_13213,N_13256);
and U13743 (N_13743,N_13116,N_13173);
or U13744 (N_13744,N_13264,N_13296);
nand U13745 (N_13745,N_13123,N_13351);
or U13746 (N_13746,N_13396,N_13414);
xnor U13747 (N_13747,N_13317,N_13138);
nor U13748 (N_13748,N_13344,N_13455);
and U13749 (N_13749,N_13459,N_13377);
nor U13750 (N_13750,N_13165,N_13123);
and U13751 (N_13751,N_13352,N_13082);
and U13752 (N_13752,N_13022,N_13490);
or U13753 (N_13753,N_13176,N_13469);
xor U13754 (N_13754,N_13236,N_13440);
xnor U13755 (N_13755,N_13092,N_13033);
nand U13756 (N_13756,N_13131,N_13302);
xnor U13757 (N_13757,N_13179,N_13437);
xnor U13758 (N_13758,N_13469,N_13181);
nor U13759 (N_13759,N_13248,N_13359);
nand U13760 (N_13760,N_13468,N_13295);
xnor U13761 (N_13761,N_13087,N_13442);
and U13762 (N_13762,N_13104,N_13111);
or U13763 (N_13763,N_13026,N_13097);
or U13764 (N_13764,N_13368,N_13157);
nand U13765 (N_13765,N_13197,N_13271);
xor U13766 (N_13766,N_13430,N_13305);
or U13767 (N_13767,N_13467,N_13097);
nand U13768 (N_13768,N_13386,N_13029);
and U13769 (N_13769,N_13327,N_13498);
and U13770 (N_13770,N_13073,N_13036);
nor U13771 (N_13771,N_13195,N_13472);
xnor U13772 (N_13772,N_13034,N_13052);
or U13773 (N_13773,N_13037,N_13020);
nand U13774 (N_13774,N_13144,N_13069);
and U13775 (N_13775,N_13192,N_13181);
nor U13776 (N_13776,N_13414,N_13426);
xnor U13777 (N_13777,N_13138,N_13272);
nor U13778 (N_13778,N_13017,N_13434);
and U13779 (N_13779,N_13094,N_13074);
xnor U13780 (N_13780,N_13123,N_13003);
or U13781 (N_13781,N_13180,N_13315);
nand U13782 (N_13782,N_13390,N_13351);
or U13783 (N_13783,N_13463,N_13192);
xnor U13784 (N_13784,N_13211,N_13296);
and U13785 (N_13785,N_13424,N_13324);
and U13786 (N_13786,N_13486,N_13215);
nor U13787 (N_13787,N_13186,N_13240);
nand U13788 (N_13788,N_13473,N_13488);
and U13789 (N_13789,N_13084,N_13023);
xor U13790 (N_13790,N_13172,N_13334);
nor U13791 (N_13791,N_13128,N_13040);
nand U13792 (N_13792,N_13228,N_13084);
and U13793 (N_13793,N_13272,N_13337);
and U13794 (N_13794,N_13434,N_13261);
or U13795 (N_13795,N_13065,N_13322);
xnor U13796 (N_13796,N_13109,N_13156);
nand U13797 (N_13797,N_13306,N_13401);
and U13798 (N_13798,N_13433,N_13383);
nor U13799 (N_13799,N_13238,N_13141);
nand U13800 (N_13800,N_13185,N_13166);
nor U13801 (N_13801,N_13404,N_13102);
and U13802 (N_13802,N_13222,N_13438);
xnor U13803 (N_13803,N_13373,N_13484);
and U13804 (N_13804,N_13232,N_13072);
nor U13805 (N_13805,N_13016,N_13251);
or U13806 (N_13806,N_13322,N_13058);
nand U13807 (N_13807,N_13443,N_13123);
nand U13808 (N_13808,N_13080,N_13350);
xor U13809 (N_13809,N_13024,N_13416);
or U13810 (N_13810,N_13462,N_13306);
or U13811 (N_13811,N_13076,N_13283);
nor U13812 (N_13812,N_13112,N_13098);
and U13813 (N_13813,N_13088,N_13166);
and U13814 (N_13814,N_13274,N_13488);
or U13815 (N_13815,N_13010,N_13026);
xor U13816 (N_13816,N_13344,N_13191);
nor U13817 (N_13817,N_13369,N_13158);
xnor U13818 (N_13818,N_13437,N_13235);
nor U13819 (N_13819,N_13014,N_13424);
nor U13820 (N_13820,N_13192,N_13366);
nor U13821 (N_13821,N_13283,N_13480);
or U13822 (N_13822,N_13092,N_13396);
or U13823 (N_13823,N_13331,N_13239);
nand U13824 (N_13824,N_13184,N_13388);
and U13825 (N_13825,N_13466,N_13184);
nand U13826 (N_13826,N_13428,N_13166);
nor U13827 (N_13827,N_13255,N_13159);
and U13828 (N_13828,N_13479,N_13455);
xor U13829 (N_13829,N_13115,N_13374);
nor U13830 (N_13830,N_13234,N_13134);
or U13831 (N_13831,N_13450,N_13458);
nand U13832 (N_13832,N_13494,N_13318);
nand U13833 (N_13833,N_13084,N_13240);
xnor U13834 (N_13834,N_13327,N_13148);
xnor U13835 (N_13835,N_13180,N_13289);
nand U13836 (N_13836,N_13294,N_13018);
nor U13837 (N_13837,N_13030,N_13303);
xnor U13838 (N_13838,N_13045,N_13060);
nor U13839 (N_13839,N_13149,N_13212);
and U13840 (N_13840,N_13191,N_13212);
nand U13841 (N_13841,N_13135,N_13499);
and U13842 (N_13842,N_13251,N_13165);
and U13843 (N_13843,N_13461,N_13038);
or U13844 (N_13844,N_13371,N_13378);
nor U13845 (N_13845,N_13455,N_13313);
or U13846 (N_13846,N_13193,N_13471);
nand U13847 (N_13847,N_13320,N_13434);
nand U13848 (N_13848,N_13386,N_13219);
nand U13849 (N_13849,N_13345,N_13497);
xor U13850 (N_13850,N_13019,N_13074);
or U13851 (N_13851,N_13349,N_13265);
nor U13852 (N_13852,N_13264,N_13082);
and U13853 (N_13853,N_13004,N_13443);
and U13854 (N_13854,N_13278,N_13214);
nor U13855 (N_13855,N_13490,N_13149);
and U13856 (N_13856,N_13221,N_13394);
nor U13857 (N_13857,N_13465,N_13235);
and U13858 (N_13858,N_13016,N_13488);
xnor U13859 (N_13859,N_13016,N_13022);
or U13860 (N_13860,N_13347,N_13194);
xor U13861 (N_13861,N_13266,N_13263);
xor U13862 (N_13862,N_13063,N_13179);
nand U13863 (N_13863,N_13435,N_13086);
or U13864 (N_13864,N_13470,N_13297);
and U13865 (N_13865,N_13437,N_13457);
nand U13866 (N_13866,N_13348,N_13165);
and U13867 (N_13867,N_13443,N_13310);
nor U13868 (N_13868,N_13028,N_13003);
and U13869 (N_13869,N_13456,N_13202);
and U13870 (N_13870,N_13026,N_13488);
or U13871 (N_13871,N_13225,N_13456);
nor U13872 (N_13872,N_13087,N_13435);
nand U13873 (N_13873,N_13190,N_13122);
and U13874 (N_13874,N_13346,N_13403);
and U13875 (N_13875,N_13434,N_13154);
nand U13876 (N_13876,N_13095,N_13366);
nand U13877 (N_13877,N_13213,N_13434);
nor U13878 (N_13878,N_13062,N_13395);
nand U13879 (N_13879,N_13488,N_13124);
or U13880 (N_13880,N_13207,N_13230);
nand U13881 (N_13881,N_13279,N_13169);
nand U13882 (N_13882,N_13041,N_13307);
nand U13883 (N_13883,N_13051,N_13324);
and U13884 (N_13884,N_13205,N_13317);
nor U13885 (N_13885,N_13019,N_13031);
nor U13886 (N_13886,N_13476,N_13463);
or U13887 (N_13887,N_13018,N_13420);
or U13888 (N_13888,N_13170,N_13326);
and U13889 (N_13889,N_13365,N_13224);
xor U13890 (N_13890,N_13301,N_13441);
or U13891 (N_13891,N_13181,N_13006);
xor U13892 (N_13892,N_13345,N_13269);
xor U13893 (N_13893,N_13420,N_13068);
nor U13894 (N_13894,N_13133,N_13375);
and U13895 (N_13895,N_13252,N_13237);
xnor U13896 (N_13896,N_13430,N_13362);
and U13897 (N_13897,N_13032,N_13494);
nand U13898 (N_13898,N_13056,N_13194);
nor U13899 (N_13899,N_13189,N_13077);
nand U13900 (N_13900,N_13111,N_13360);
xnor U13901 (N_13901,N_13064,N_13126);
nand U13902 (N_13902,N_13069,N_13060);
nand U13903 (N_13903,N_13403,N_13419);
or U13904 (N_13904,N_13462,N_13318);
and U13905 (N_13905,N_13309,N_13248);
xnor U13906 (N_13906,N_13030,N_13441);
nor U13907 (N_13907,N_13320,N_13448);
and U13908 (N_13908,N_13390,N_13298);
nor U13909 (N_13909,N_13233,N_13118);
nor U13910 (N_13910,N_13421,N_13099);
or U13911 (N_13911,N_13389,N_13408);
and U13912 (N_13912,N_13125,N_13223);
xor U13913 (N_13913,N_13310,N_13230);
xor U13914 (N_13914,N_13140,N_13445);
nand U13915 (N_13915,N_13398,N_13044);
nand U13916 (N_13916,N_13324,N_13061);
nand U13917 (N_13917,N_13010,N_13494);
xnor U13918 (N_13918,N_13030,N_13045);
xnor U13919 (N_13919,N_13335,N_13283);
and U13920 (N_13920,N_13418,N_13123);
xor U13921 (N_13921,N_13010,N_13204);
or U13922 (N_13922,N_13338,N_13211);
nand U13923 (N_13923,N_13207,N_13412);
and U13924 (N_13924,N_13300,N_13270);
and U13925 (N_13925,N_13207,N_13498);
xor U13926 (N_13926,N_13249,N_13196);
nor U13927 (N_13927,N_13341,N_13011);
xor U13928 (N_13928,N_13498,N_13089);
nand U13929 (N_13929,N_13031,N_13431);
nand U13930 (N_13930,N_13235,N_13364);
and U13931 (N_13931,N_13298,N_13196);
or U13932 (N_13932,N_13298,N_13214);
or U13933 (N_13933,N_13117,N_13239);
and U13934 (N_13934,N_13270,N_13415);
xor U13935 (N_13935,N_13093,N_13236);
nor U13936 (N_13936,N_13073,N_13111);
nand U13937 (N_13937,N_13106,N_13035);
nand U13938 (N_13938,N_13300,N_13307);
nand U13939 (N_13939,N_13124,N_13104);
or U13940 (N_13940,N_13303,N_13367);
nor U13941 (N_13941,N_13013,N_13118);
nor U13942 (N_13942,N_13428,N_13142);
and U13943 (N_13943,N_13209,N_13146);
or U13944 (N_13944,N_13258,N_13023);
or U13945 (N_13945,N_13030,N_13237);
xor U13946 (N_13946,N_13430,N_13489);
nor U13947 (N_13947,N_13273,N_13290);
nor U13948 (N_13948,N_13415,N_13123);
or U13949 (N_13949,N_13179,N_13273);
nand U13950 (N_13950,N_13417,N_13049);
xor U13951 (N_13951,N_13365,N_13103);
xnor U13952 (N_13952,N_13090,N_13480);
nor U13953 (N_13953,N_13348,N_13477);
or U13954 (N_13954,N_13221,N_13383);
nand U13955 (N_13955,N_13199,N_13097);
and U13956 (N_13956,N_13346,N_13449);
nor U13957 (N_13957,N_13311,N_13119);
nand U13958 (N_13958,N_13252,N_13192);
and U13959 (N_13959,N_13188,N_13136);
and U13960 (N_13960,N_13086,N_13003);
or U13961 (N_13961,N_13254,N_13053);
or U13962 (N_13962,N_13023,N_13059);
and U13963 (N_13963,N_13314,N_13257);
xor U13964 (N_13964,N_13449,N_13396);
and U13965 (N_13965,N_13280,N_13479);
and U13966 (N_13966,N_13179,N_13060);
and U13967 (N_13967,N_13471,N_13436);
nor U13968 (N_13968,N_13222,N_13194);
nor U13969 (N_13969,N_13397,N_13419);
nand U13970 (N_13970,N_13349,N_13462);
xor U13971 (N_13971,N_13379,N_13341);
xor U13972 (N_13972,N_13012,N_13345);
xor U13973 (N_13973,N_13404,N_13098);
xnor U13974 (N_13974,N_13221,N_13241);
or U13975 (N_13975,N_13372,N_13390);
and U13976 (N_13976,N_13338,N_13402);
or U13977 (N_13977,N_13218,N_13335);
nor U13978 (N_13978,N_13327,N_13182);
xor U13979 (N_13979,N_13149,N_13263);
nand U13980 (N_13980,N_13291,N_13354);
and U13981 (N_13981,N_13082,N_13254);
nand U13982 (N_13982,N_13091,N_13199);
and U13983 (N_13983,N_13133,N_13428);
xnor U13984 (N_13984,N_13103,N_13089);
nor U13985 (N_13985,N_13455,N_13088);
xor U13986 (N_13986,N_13417,N_13002);
or U13987 (N_13987,N_13409,N_13169);
xnor U13988 (N_13988,N_13044,N_13056);
and U13989 (N_13989,N_13314,N_13154);
nand U13990 (N_13990,N_13138,N_13041);
and U13991 (N_13991,N_13355,N_13202);
nand U13992 (N_13992,N_13480,N_13285);
xnor U13993 (N_13993,N_13034,N_13402);
nand U13994 (N_13994,N_13156,N_13206);
nand U13995 (N_13995,N_13377,N_13032);
or U13996 (N_13996,N_13003,N_13025);
xnor U13997 (N_13997,N_13409,N_13090);
nand U13998 (N_13998,N_13406,N_13242);
and U13999 (N_13999,N_13133,N_13251);
and U14000 (N_14000,N_13613,N_13525);
or U14001 (N_14001,N_13767,N_13812);
nor U14002 (N_14002,N_13694,N_13833);
or U14003 (N_14003,N_13878,N_13869);
nor U14004 (N_14004,N_13827,N_13746);
xnor U14005 (N_14005,N_13862,N_13665);
and U14006 (N_14006,N_13765,N_13639);
and U14007 (N_14007,N_13588,N_13944);
or U14008 (N_14008,N_13832,N_13779);
nor U14009 (N_14009,N_13899,N_13573);
and U14010 (N_14010,N_13728,N_13753);
nand U14011 (N_14011,N_13768,N_13824);
nand U14012 (N_14012,N_13763,N_13641);
and U14013 (N_14013,N_13887,N_13582);
or U14014 (N_14014,N_13871,N_13519);
nand U14015 (N_14015,N_13934,N_13638);
nor U14016 (N_14016,N_13806,N_13757);
nand U14017 (N_14017,N_13885,N_13601);
nand U14018 (N_14018,N_13705,N_13707);
xor U14019 (N_14019,N_13595,N_13654);
xor U14020 (N_14020,N_13541,N_13709);
or U14021 (N_14021,N_13546,N_13627);
or U14022 (N_14022,N_13677,N_13791);
nand U14023 (N_14023,N_13984,N_13748);
or U14024 (N_14024,N_13905,N_13852);
nand U14025 (N_14025,N_13835,N_13745);
nor U14026 (N_14026,N_13720,N_13895);
nor U14027 (N_14027,N_13716,N_13931);
nand U14028 (N_14028,N_13772,N_13744);
xnor U14029 (N_14029,N_13840,N_13956);
nor U14030 (N_14030,N_13633,N_13969);
xnor U14031 (N_14031,N_13605,N_13618);
nand U14032 (N_14032,N_13620,N_13859);
nor U14033 (N_14033,N_13894,N_13864);
or U14034 (N_14034,N_13623,N_13794);
nor U14035 (N_14035,N_13922,N_13965);
nor U14036 (N_14036,N_13713,N_13673);
xor U14037 (N_14037,N_13698,N_13567);
or U14038 (N_14038,N_13820,N_13843);
nand U14039 (N_14039,N_13529,N_13955);
and U14040 (N_14040,N_13921,N_13540);
xor U14041 (N_14041,N_13731,N_13509);
or U14042 (N_14042,N_13524,N_13847);
and U14043 (N_14043,N_13874,N_13552);
and U14044 (N_14044,N_13953,N_13930);
nor U14045 (N_14045,N_13981,N_13947);
or U14046 (N_14046,N_13801,N_13816);
and U14047 (N_14047,N_13640,N_13544);
or U14048 (N_14048,N_13932,N_13752);
nand U14049 (N_14049,N_13615,N_13811);
and U14050 (N_14050,N_13534,N_13802);
xor U14051 (N_14051,N_13651,N_13821);
xnor U14052 (N_14052,N_13732,N_13866);
nor U14053 (N_14053,N_13844,N_13590);
nand U14054 (N_14054,N_13635,N_13822);
and U14055 (N_14055,N_13915,N_13626);
nor U14056 (N_14056,N_13780,N_13880);
xor U14057 (N_14057,N_13998,N_13892);
or U14058 (N_14058,N_13838,N_13531);
nand U14059 (N_14059,N_13616,N_13828);
nand U14060 (N_14060,N_13867,N_13689);
or U14061 (N_14061,N_13653,N_13660);
and U14062 (N_14062,N_13942,N_13989);
or U14063 (N_14063,N_13946,N_13789);
xnor U14064 (N_14064,N_13517,N_13991);
nor U14065 (N_14065,N_13629,N_13773);
nor U14066 (N_14066,N_13549,N_13657);
nor U14067 (N_14067,N_13804,N_13542);
nor U14068 (N_14068,N_13697,N_13726);
xnor U14069 (N_14069,N_13670,N_13917);
xor U14070 (N_14070,N_13858,N_13817);
nand U14071 (N_14071,N_13788,N_13888);
or U14072 (N_14072,N_13592,N_13814);
xnor U14073 (N_14073,N_13950,N_13667);
and U14074 (N_14074,N_13987,N_13877);
nor U14075 (N_14075,N_13719,N_13591);
nand U14076 (N_14076,N_13976,N_13703);
or U14077 (N_14077,N_13636,N_13537);
xnor U14078 (N_14078,N_13902,N_13522);
xnor U14079 (N_14079,N_13668,N_13882);
and U14080 (N_14080,N_13586,N_13577);
and U14081 (N_14081,N_13696,N_13557);
xnor U14082 (N_14082,N_13712,N_13523);
or U14083 (N_14083,N_13725,N_13553);
xor U14084 (N_14084,N_13513,N_13808);
nor U14085 (N_14085,N_13711,N_13778);
nor U14086 (N_14086,N_13730,N_13756);
and U14087 (N_14087,N_13505,N_13585);
xnor U14088 (N_14088,N_13996,N_13511);
xnor U14089 (N_14089,N_13680,N_13790);
xnor U14090 (N_14090,N_13960,N_13762);
xor U14091 (N_14091,N_13749,N_13562);
nand U14092 (N_14092,N_13554,N_13611);
xor U14093 (N_14093,N_13920,N_13543);
nor U14094 (N_14094,N_13649,N_13907);
nand U14095 (N_14095,N_13565,N_13970);
or U14096 (N_14096,N_13848,N_13823);
nor U14097 (N_14097,N_13723,N_13959);
xor U14098 (N_14098,N_13760,N_13708);
xnor U14099 (N_14099,N_13584,N_13674);
or U14100 (N_14100,N_13658,N_13928);
and U14101 (N_14101,N_13842,N_13625);
xor U14102 (N_14102,N_13671,N_13691);
nor U14103 (N_14103,N_13906,N_13581);
and U14104 (N_14104,N_13503,N_13643);
xnor U14105 (N_14105,N_13617,N_13722);
or U14106 (N_14106,N_13646,N_13644);
or U14107 (N_14107,N_13770,N_13958);
or U14108 (N_14108,N_13684,N_13837);
nand U14109 (N_14109,N_13841,N_13936);
nor U14110 (N_14110,N_13815,N_13701);
or U14111 (N_14111,N_13632,N_13904);
or U14112 (N_14112,N_13809,N_13662);
xnor U14113 (N_14113,N_13539,N_13783);
xnor U14114 (N_14114,N_13926,N_13851);
or U14115 (N_14115,N_13507,N_13704);
nor U14116 (N_14116,N_13520,N_13807);
and U14117 (N_14117,N_13729,N_13758);
and U14118 (N_14118,N_13900,N_13890);
or U14119 (N_14119,N_13710,N_13571);
xnor U14120 (N_14120,N_13865,N_13576);
or U14121 (N_14121,N_13800,N_13810);
or U14122 (N_14122,N_13980,N_13868);
or U14123 (N_14123,N_13898,N_13533);
nor U14124 (N_14124,N_13631,N_13943);
nand U14125 (N_14125,N_13558,N_13805);
and U14126 (N_14126,N_13737,N_13655);
or U14127 (N_14127,N_13661,N_13974);
and U14128 (N_14128,N_13672,N_13982);
nor U14129 (N_14129,N_13854,N_13594);
nand U14130 (N_14130,N_13938,N_13609);
nand U14131 (N_14131,N_13963,N_13962);
xnor U14132 (N_14132,N_13999,N_13536);
nand U14133 (N_14133,N_13622,N_13574);
xor U14134 (N_14134,N_13836,N_13985);
nand U14135 (N_14135,N_13538,N_13717);
nand U14136 (N_14136,N_13608,N_13714);
or U14137 (N_14137,N_13669,N_13742);
or U14138 (N_14138,N_13939,N_13819);
nor U14139 (N_14139,N_13530,N_13831);
or U14140 (N_14140,N_13604,N_13516);
nor U14141 (N_14141,N_13951,N_13621);
nor U14142 (N_14142,N_13645,N_13897);
xor U14143 (N_14143,N_13515,N_13580);
nand U14144 (N_14144,N_13500,N_13769);
xor U14145 (N_14145,N_13687,N_13518);
or U14146 (N_14146,N_13675,N_13555);
or U14147 (N_14147,N_13872,N_13978);
nor U14148 (N_14148,N_13750,N_13724);
nand U14149 (N_14149,N_13619,N_13508);
and U14150 (N_14150,N_13785,N_13830);
nand U14151 (N_14151,N_13521,N_13688);
or U14152 (N_14152,N_13919,N_13849);
nor U14153 (N_14153,N_13964,N_13966);
nand U14154 (N_14154,N_13940,N_13861);
or U14155 (N_14155,N_13683,N_13600);
nor U14156 (N_14156,N_13875,N_13990);
xor U14157 (N_14157,N_13647,N_13891);
xor U14158 (N_14158,N_13634,N_13781);
nor U14159 (N_14159,N_13776,N_13925);
nor U14160 (N_14160,N_13528,N_13829);
nor U14161 (N_14161,N_13692,N_13826);
nor U14162 (N_14162,N_13702,N_13550);
nor U14163 (N_14163,N_13873,N_13504);
and U14164 (N_14164,N_13918,N_13761);
nor U14165 (N_14165,N_13798,N_13909);
and U14166 (N_14166,N_13648,N_13771);
and U14167 (N_14167,N_13913,N_13889);
xor U14168 (N_14168,N_13563,N_13883);
and U14169 (N_14169,N_13727,N_13997);
nand U14170 (N_14170,N_13568,N_13695);
xor U14171 (N_14171,N_13602,N_13532);
nor U14172 (N_14172,N_13570,N_13579);
and U14173 (N_14173,N_13863,N_13628);
xnor U14174 (N_14174,N_13569,N_13954);
nor U14175 (N_14175,N_13792,N_13656);
and U14176 (N_14176,N_13968,N_13766);
nor U14177 (N_14177,N_13715,N_13652);
and U14178 (N_14178,N_13593,N_13855);
xnor U14179 (N_14179,N_13583,N_13949);
nor U14180 (N_14180,N_13986,N_13948);
and U14181 (N_14181,N_13572,N_13607);
and U14182 (N_14182,N_13912,N_13825);
nor U14183 (N_14183,N_13774,N_13834);
nand U14184 (N_14184,N_13512,N_13735);
xnor U14185 (N_14185,N_13685,N_13911);
xnor U14186 (N_14186,N_13642,N_13977);
nand U14187 (N_14187,N_13856,N_13501);
nand U14188 (N_14188,N_13664,N_13679);
xor U14189 (N_14189,N_13739,N_13681);
and U14190 (N_14190,N_13559,N_13983);
or U14191 (N_14191,N_13957,N_13603);
or U14192 (N_14192,N_13782,N_13850);
and U14193 (N_14193,N_13721,N_13860);
and U14194 (N_14194,N_13933,N_13527);
or U14195 (N_14195,N_13598,N_13736);
nor U14196 (N_14196,N_13813,N_13740);
or U14197 (N_14197,N_13937,N_13799);
or U14198 (N_14198,N_13666,N_13718);
xor U14199 (N_14199,N_13994,N_13548);
nand U14200 (N_14200,N_13857,N_13741);
and U14201 (N_14201,N_13995,N_13846);
xor U14202 (N_14202,N_13693,N_13796);
and U14203 (N_14203,N_13876,N_13733);
xor U14204 (N_14204,N_13514,N_13775);
nor U14205 (N_14205,N_13893,N_13923);
nor U14206 (N_14206,N_13526,N_13614);
and U14207 (N_14207,N_13818,N_13786);
nor U14208 (N_14208,N_13787,N_13993);
or U14209 (N_14209,N_13839,N_13924);
nor U14210 (N_14210,N_13637,N_13908);
nand U14211 (N_14211,N_13564,N_13929);
and U14212 (N_14212,N_13545,N_13886);
xor U14213 (N_14213,N_13663,N_13764);
nor U14214 (N_14214,N_13560,N_13612);
nand U14215 (N_14215,N_13678,N_13927);
nand U14216 (N_14216,N_13979,N_13945);
and U14217 (N_14217,N_13743,N_13578);
and U14218 (N_14218,N_13700,N_13587);
nand U14219 (N_14219,N_13682,N_13597);
nand U14220 (N_14220,N_13575,N_13510);
and U14221 (N_14221,N_13784,N_13734);
or U14222 (N_14222,N_13879,N_13961);
and U14223 (N_14223,N_13676,N_13884);
nor U14224 (N_14224,N_13941,N_13973);
nand U14225 (N_14225,N_13901,N_13738);
and U14226 (N_14226,N_13967,N_13610);
nor U14227 (N_14227,N_13754,N_13975);
nor U14228 (N_14228,N_13755,N_13903);
nor U14229 (N_14229,N_13686,N_13845);
nor U14230 (N_14230,N_13971,N_13795);
and U14231 (N_14231,N_13896,N_13972);
or U14232 (N_14232,N_13777,N_13803);
nand U14233 (N_14233,N_13853,N_13535);
nor U14234 (N_14234,N_13502,N_13910);
xor U14235 (N_14235,N_13506,N_13699);
and U14236 (N_14236,N_13589,N_13596);
nand U14237 (N_14237,N_13747,N_13650);
xnor U14238 (N_14238,N_13659,N_13551);
or U14239 (N_14239,N_13561,N_13599);
or U14240 (N_14240,N_13935,N_13624);
nand U14241 (N_14241,N_13751,N_13952);
nand U14242 (N_14242,N_13759,N_13870);
xor U14243 (N_14243,N_13690,N_13988);
or U14244 (N_14244,N_13793,N_13992);
or U14245 (N_14245,N_13556,N_13547);
xnor U14246 (N_14246,N_13706,N_13606);
nor U14247 (N_14247,N_13566,N_13797);
nand U14248 (N_14248,N_13914,N_13630);
nand U14249 (N_14249,N_13881,N_13916);
xor U14250 (N_14250,N_13710,N_13559);
xor U14251 (N_14251,N_13877,N_13651);
or U14252 (N_14252,N_13824,N_13537);
or U14253 (N_14253,N_13511,N_13517);
and U14254 (N_14254,N_13604,N_13680);
and U14255 (N_14255,N_13591,N_13989);
nor U14256 (N_14256,N_13945,N_13760);
nor U14257 (N_14257,N_13939,N_13705);
nor U14258 (N_14258,N_13541,N_13577);
nor U14259 (N_14259,N_13855,N_13740);
or U14260 (N_14260,N_13542,N_13643);
nor U14261 (N_14261,N_13662,N_13940);
and U14262 (N_14262,N_13504,N_13724);
or U14263 (N_14263,N_13626,N_13639);
or U14264 (N_14264,N_13530,N_13543);
nor U14265 (N_14265,N_13550,N_13903);
nor U14266 (N_14266,N_13896,N_13657);
and U14267 (N_14267,N_13719,N_13712);
nor U14268 (N_14268,N_13963,N_13528);
and U14269 (N_14269,N_13820,N_13631);
or U14270 (N_14270,N_13828,N_13745);
xnor U14271 (N_14271,N_13885,N_13961);
nand U14272 (N_14272,N_13552,N_13540);
nor U14273 (N_14273,N_13709,N_13617);
nor U14274 (N_14274,N_13852,N_13881);
nand U14275 (N_14275,N_13771,N_13573);
xor U14276 (N_14276,N_13722,N_13957);
nor U14277 (N_14277,N_13823,N_13799);
and U14278 (N_14278,N_13846,N_13536);
or U14279 (N_14279,N_13820,N_13796);
nor U14280 (N_14280,N_13954,N_13791);
and U14281 (N_14281,N_13518,N_13985);
nand U14282 (N_14282,N_13666,N_13845);
or U14283 (N_14283,N_13598,N_13519);
nor U14284 (N_14284,N_13854,N_13814);
nand U14285 (N_14285,N_13504,N_13812);
or U14286 (N_14286,N_13521,N_13768);
and U14287 (N_14287,N_13849,N_13710);
nand U14288 (N_14288,N_13970,N_13755);
and U14289 (N_14289,N_13604,N_13901);
or U14290 (N_14290,N_13588,N_13604);
nand U14291 (N_14291,N_13504,N_13959);
xor U14292 (N_14292,N_13904,N_13844);
nor U14293 (N_14293,N_13975,N_13532);
xor U14294 (N_14294,N_13954,N_13574);
nor U14295 (N_14295,N_13747,N_13689);
and U14296 (N_14296,N_13686,N_13642);
and U14297 (N_14297,N_13791,N_13588);
and U14298 (N_14298,N_13604,N_13506);
or U14299 (N_14299,N_13882,N_13767);
xor U14300 (N_14300,N_13649,N_13852);
nand U14301 (N_14301,N_13748,N_13622);
xnor U14302 (N_14302,N_13566,N_13931);
nand U14303 (N_14303,N_13998,N_13648);
xnor U14304 (N_14304,N_13963,N_13517);
nand U14305 (N_14305,N_13641,N_13951);
nand U14306 (N_14306,N_13851,N_13767);
nor U14307 (N_14307,N_13598,N_13594);
and U14308 (N_14308,N_13620,N_13615);
nor U14309 (N_14309,N_13834,N_13728);
nor U14310 (N_14310,N_13559,N_13859);
nand U14311 (N_14311,N_13788,N_13935);
nand U14312 (N_14312,N_13571,N_13717);
nor U14313 (N_14313,N_13940,N_13786);
nor U14314 (N_14314,N_13657,N_13833);
and U14315 (N_14315,N_13838,N_13905);
or U14316 (N_14316,N_13529,N_13905);
xnor U14317 (N_14317,N_13817,N_13518);
nand U14318 (N_14318,N_13797,N_13677);
nor U14319 (N_14319,N_13830,N_13825);
and U14320 (N_14320,N_13658,N_13632);
or U14321 (N_14321,N_13556,N_13786);
nand U14322 (N_14322,N_13945,N_13990);
or U14323 (N_14323,N_13809,N_13617);
and U14324 (N_14324,N_13567,N_13886);
xnor U14325 (N_14325,N_13967,N_13687);
xor U14326 (N_14326,N_13932,N_13808);
xor U14327 (N_14327,N_13516,N_13666);
or U14328 (N_14328,N_13659,N_13785);
or U14329 (N_14329,N_13696,N_13918);
or U14330 (N_14330,N_13823,N_13568);
and U14331 (N_14331,N_13589,N_13772);
or U14332 (N_14332,N_13697,N_13620);
nand U14333 (N_14333,N_13721,N_13995);
xnor U14334 (N_14334,N_13874,N_13522);
nor U14335 (N_14335,N_13682,N_13940);
xor U14336 (N_14336,N_13557,N_13889);
and U14337 (N_14337,N_13689,N_13888);
xor U14338 (N_14338,N_13730,N_13547);
and U14339 (N_14339,N_13850,N_13622);
or U14340 (N_14340,N_13875,N_13515);
xnor U14341 (N_14341,N_13888,N_13824);
and U14342 (N_14342,N_13782,N_13894);
nand U14343 (N_14343,N_13543,N_13690);
nor U14344 (N_14344,N_13735,N_13834);
xnor U14345 (N_14345,N_13975,N_13925);
nand U14346 (N_14346,N_13719,N_13995);
or U14347 (N_14347,N_13614,N_13649);
nor U14348 (N_14348,N_13856,N_13565);
or U14349 (N_14349,N_13614,N_13528);
nor U14350 (N_14350,N_13671,N_13700);
and U14351 (N_14351,N_13954,N_13860);
nor U14352 (N_14352,N_13729,N_13818);
and U14353 (N_14353,N_13869,N_13555);
nand U14354 (N_14354,N_13693,N_13597);
or U14355 (N_14355,N_13771,N_13790);
xor U14356 (N_14356,N_13519,N_13771);
xnor U14357 (N_14357,N_13785,N_13592);
xor U14358 (N_14358,N_13585,N_13617);
nand U14359 (N_14359,N_13870,N_13897);
and U14360 (N_14360,N_13651,N_13887);
and U14361 (N_14361,N_13913,N_13585);
xor U14362 (N_14362,N_13702,N_13647);
xnor U14363 (N_14363,N_13775,N_13926);
nor U14364 (N_14364,N_13659,N_13643);
xnor U14365 (N_14365,N_13749,N_13798);
xnor U14366 (N_14366,N_13500,N_13903);
and U14367 (N_14367,N_13767,N_13623);
and U14368 (N_14368,N_13803,N_13948);
and U14369 (N_14369,N_13564,N_13774);
nor U14370 (N_14370,N_13900,N_13995);
and U14371 (N_14371,N_13577,N_13779);
nor U14372 (N_14372,N_13788,N_13950);
nor U14373 (N_14373,N_13795,N_13714);
xor U14374 (N_14374,N_13902,N_13724);
or U14375 (N_14375,N_13875,N_13910);
and U14376 (N_14376,N_13842,N_13893);
and U14377 (N_14377,N_13647,N_13566);
nand U14378 (N_14378,N_13608,N_13942);
nor U14379 (N_14379,N_13983,N_13991);
and U14380 (N_14380,N_13882,N_13998);
nor U14381 (N_14381,N_13766,N_13555);
nor U14382 (N_14382,N_13669,N_13654);
xnor U14383 (N_14383,N_13849,N_13700);
nand U14384 (N_14384,N_13554,N_13582);
nand U14385 (N_14385,N_13527,N_13886);
and U14386 (N_14386,N_13610,N_13938);
xnor U14387 (N_14387,N_13616,N_13866);
and U14388 (N_14388,N_13688,N_13627);
nand U14389 (N_14389,N_13730,N_13642);
nor U14390 (N_14390,N_13517,N_13976);
or U14391 (N_14391,N_13505,N_13987);
and U14392 (N_14392,N_13609,N_13748);
nor U14393 (N_14393,N_13992,N_13773);
nor U14394 (N_14394,N_13896,N_13631);
nor U14395 (N_14395,N_13623,N_13914);
nor U14396 (N_14396,N_13565,N_13663);
and U14397 (N_14397,N_13983,N_13918);
nand U14398 (N_14398,N_13620,N_13721);
or U14399 (N_14399,N_13675,N_13819);
nor U14400 (N_14400,N_13985,N_13578);
or U14401 (N_14401,N_13608,N_13997);
xnor U14402 (N_14402,N_13799,N_13712);
or U14403 (N_14403,N_13664,N_13803);
nand U14404 (N_14404,N_13767,N_13708);
nand U14405 (N_14405,N_13934,N_13695);
and U14406 (N_14406,N_13874,N_13904);
xnor U14407 (N_14407,N_13731,N_13707);
nor U14408 (N_14408,N_13883,N_13512);
nor U14409 (N_14409,N_13830,N_13828);
xnor U14410 (N_14410,N_13875,N_13743);
xnor U14411 (N_14411,N_13939,N_13842);
and U14412 (N_14412,N_13906,N_13656);
or U14413 (N_14413,N_13681,N_13986);
and U14414 (N_14414,N_13838,N_13520);
and U14415 (N_14415,N_13814,N_13725);
nand U14416 (N_14416,N_13639,N_13501);
xnor U14417 (N_14417,N_13605,N_13523);
xor U14418 (N_14418,N_13962,N_13779);
or U14419 (N_14419,N_13976,N_13832);
xnor U14420 (N_14420,N_13759,N_13850);
nor U14421 (N_14421,N_13722,N_13636);
or U14422 (N_14422,N_13996,N_13924);
and U14423 (N_14423,N_13612,N_13518);
xor U14424 (N_14424,N_13838,N_13791);
or U14425 (N_14425,N_13535,N_13833);
and U14426 (N_14426,N_13750,N_13599);
nor U14427 (N_14427,N_13670,N_13618);
and U14428 (N_14428,N_13980,N_13889);
or U14429 (N_14429,N_13680,N_13949);
nand U14430 (N_14430,N_13734,N_13731);
nand U14431 (N_14431,N_13905,N_13566);
nand U14432 (N_14432,N_13526,N_13503);
and U14433 (N_14433,N_13569,N_13640);
or U14434 (N_14434,N_13629,N_13711);
xor U14435 (N_14435,N_13705,N_13534);
nor U14436 (N_14436,N_13969,N_13921);
nor U14437 (N_14437,N_13768,N_13643);
nand U14438 (N_14438,N_13712,N_13862);
nor U14439 (N_14439,N_13620,N_13851);
xnor U14440 (N_14440,N_13937,N_13639);
nand U14441 (N_14441,N_13543,N_13609);
or U14442 (N_14442,N_13890,N_13954);
nor U14443 (N_14443,N_13831,N_13903);
and U14444 (N_14444,N_13650,N_13716);
nor U14445 (N_14445,N_13693,N_13639);
xnor U14446 (N_14446,N_13844,N_13983);
and U14447 (N_14447,N_13657,N_13683);
or U14448 (N_14448,N_13708,N_13616);
nand U14449 (N_14449,N_13856,N_13728);
nand U14450 (N_14450,N_13579,N_13681);
or U14451 (N_14451,N_13964,N_13948);
xnor U14452 (N_14452,N_13904,N_13756);
nor U14453 (N_14453,N_13621,N_13846);
nor U14454 (N_14454,N_13670,N_13679);
xor U14455 (N_14455,N_13639,N_13851);
and U14456 (N_14456,N_13708,N_13516);
or U14457 (N_14457,N_13982,N_13754);
nand U14458 (N_14458,N_13884,N_13696);
xnor U14459 (N_14459,N_13830,N_13596);
nor U14460 (N_14460,N_13727,N_13951);
nor U14461 (N_14461,N_13769,N_13985);
or U14462 (N_14462,N_13830,N_13728);
xnor U14463 (N_14463,N_13931,N_13682);
and U14464 (N_14464,N_13798,N_13918);
xnor U14465 (N_14465,N_13822,N_13748);
or U14466 (N_14466,N_13964,N_13598);
nor U14467 (N_14467,N_13564,N_13530);
nand U14468 (N_14468,N_13778,N_13526);
xnor U14469 (N_14469,N_13664,N_13866);
xor U14470 (N_14470,N_13567,N_13810);
nand U14471 (N_14471,N_13650,N_13659);
or U14472 (N_14472,N_13684,N_13537);
xnor U14473 (N_14473,N_13855,N_13668);
nor U14474 (N_14474,N_13878,N_13890);
or U14475 (N_14475,N_13798,N_13799);
nand U14476 (N_14476,N_13641,N_13577);
or U14477 (N_14477,N_13712,N_13555);
and U14478 (N_14478,N_13848,N_13775);
or U14479 (N_14479,N_13518,N_13920);
nand U14480 (N_14480,N_13644,N_13715);
nor U14481 (N_14481,N_13856,N_13983);
or U14482 (N_14482,N_13503,N_13604);
and U14483 (N_14483,N_13613,N_13734);
nor U14484 (N_14484,N_13950,N_13922);
nand U14485 (N_14485,N_13748,N_13836);
and U14486 (N_14486,N_13923,N_13731);
or U14487 (N_14487,N_13855,N_13667);
or U14488 (N_14488,N_13981,N_13873);
nor U14489 (N_14489,N_13801,N_13516);
or U14490 (N_14490,N_13580,N_13608);
nand U14491 (N_14491,N_13842,N_13706);
nand U14492 (N_14492,N_13627,N_13540);
xnor U14493 (N_14493,N_13740,N_13880);
nor U14494 (N_14494,N_13947,N_13703);
or U14495 (N_14495,N_13860,N_13760);
nor U14496 (N_14496,N_13599,N_13932);
and U14497 (N_14497,N_13686,N_13637);
and U14498 (N_14498,N_13601,N_13683);
nand U14499 (N_14499,N_13580,N_13987);
xnor U14500 (N_14500,N_14395,N_14323);
xnor U14501 (N_14501,N_14404,N_14451);
nand U14502 (N_14502,N_14016,N_14067);
nor U14503 (N_14503,N_14337,N_14023);
nor U14504 (N_14504,N_14153,N_14454);
or U14505 (N_14505,N_14229,N_14203);
nor U14506 (N_14506,N_14078,N_14358);
nand U14507 (N_14507,N_14316,N_14244);
xor U14508 (N_14508,N_14044,N_14467);
nand U14509 (N_14509,N_14331,N_14371);
nor U14510 (N_14510,N_14264,N_14472);
nor U14511 (N_14511,N_14010,N_14362);
xor U14512 (N_14512,N_14062,N_14150);
nor U14513 (N_14513,N_14131,N_14299);
nor U14514 (N_14514,N_14046,N_14034);
nand U14515 (N_14515,N_14164,N_14145);
or U14516 (N_14516,N_14444,N_14352);
nand U14517 (N_14517,N_14484,N_14367);
or U14518 (N_14518,N_14090,N_14301);
nand U14519 (N_14519,N_14402,N_14054);
nand U14520 (N_14520,N_14155,N_14238);
nand U14521 (N_14521,N_14359,N_14031);
xor U14522 (N_14522,N_14329,N_14220);
xnor U14523 (N_14523,N_14194,N_14324);
and U14524 (N_14524,N_14284,N_14468);
xnor U14525 (N_14525,N_14303,N_14428);
and U14526 (N_14526,N_14386,N_14443);
nand U14527 (N_14527,N_14192,N_14245);
and U14528 (N_14528,N_14388,N_14257);
xnor U14529 (N_14529,N_14374,N_14426);
xor U14530 (N_14530,N_14343,N_14030);
or U14531 (N_14531,N_14469,N_14411);
nor U14532 (N_14532,N_14333,N_14311);
nand U14533 (N_14533,N_14157,N_14247);
nand U14534 (N_14534,N_14189,N_14137);
and U14535 (N_14535,N_14277,N_14384);
nor U14536 (N_14536,N_14136,N_14313);
xor U14537 (N_14537,N_14011,N_14015);
nor U14538 (N_14538,N_14085,N_14409);
nor U14539 (N_14539,N_14278,N_14003);
xor U14540 (N_14540,N_14498,N_14108);
nor U14541 (N_14541,N_14120,N_14250);
nor U14542 (N_14542,N_14349,N_14355);
nor U14543 (N_14543,N_14453,N_14483);
nor U14544 (N_14544,N_14341,N_14289);
and U14545 (N_14545,N_14219,N_14173);
or U14546 (N_14546,N_14288,N_14042);
and U14547 (N_14547,N_14401,N_14394);
or U14548 (N_14548,N_14148,N_14012);
or U14549 (N_14549,N_14475,N_14281);
or U14550 (N_14550,N_14266,N_14061);
xnor U14551 (N_14551,N_14217,N_14246);
and U14552 (N_14552,N_14024,N_14287);
or U14553 (N_14553,N_14378,N_14235);
xor U14554 (N_14554,N_14140,N_14464);
and U14555 (N_14555,N_14332,N_14263);
nand U14556 (N_14556,N_14124,N_14122);
xor U14557 (N_14557,N_14160,N_14424);
and U14558 (N_14558,N_14065,N_14017);
nand U14559 (N_14559,N_14072,N_14013);
xnor U14560 (N_14560,N_14261,N_14115);
or U14561 (N_14561,N_14038,N_14482);
xnor U14562 (N_14562,N_14082,N_14095);
and U14563 (N_14563,N_14066,N_14052);
nand U14564 (N_14564,N_14112,N_14109);
xnor U14565 (N_14565,N_14285,N_14129);
or U14566 (N_14566,N_14460,N_14178);
and U14567 (N_14567,N_14043,N_14369);
or U14568 (N_14568,N_14172,N_14181);
xnor U14569 (N_14569,N_14224,N_14350);
xor U14570 (N_14570,N_14319,N_14166);
and U14571 (N_14571,N_14214,N_14279);
and U14572 (N_14572,N_14184,N_14037);
nor U14573 (N_14573,N_14159,N_14191);
nor U14574 (N_14574,N_14363,N_14373);
nand U14575 (N_14575,N_14312,N_14347);
nand U14576 (N_14576,N_14200,N_14376);
nand U14577 (N_14577,N_14255,N_14199);
xnor U14578 (N_14578,N_14187,N_14293);
xnor U14579 (N_14579,N_14300,N_14274);
or U14580 (N_14580,N_14138,N_14380);
and U14581 (N_14581,N_14391,N_14008);
or U14582 (N_14582,N_14403,N_14215);
nor U14583 (N_14583,N_14387,N_14130);
nor U14584 (N_14584,N_14121,N_14437);
nor U14585 (N_14585,N_14473,N_14465);
and U14586 (N_14586,N_14056,N_14001);
and U14587 (N_14587,N_14190,N_14383);
xor U14588 (N_14588,N_14294,N_14476);
nand U14589 (N_14589,N_14413,N_14055);
and U14590 (N_14590,N_14096,N_14357);
and U14591 (N_14591,N_14099,N_14059);
or U14592 (N_14592,N_14168,N_14417);
and U14593 (N_14593,N_14233,N_14040);
and U14594 (N_14594,N_14158,N_14407);
nor U14595 (N_14595,N_14005,N_14119);
xor U14596 (N_14596,N_14273,N_14009);
nand U14597 (N_14597,N_14340,N_14098);
and U14598 (N_14598,N_14249,N_14075);
or U14599 (N_14599,N_14211,N_14047);
xor U14600 (N_14600,N_14149,N_14458);
nand U14601 (N_14601,N_14182,N_14496);
and U14602 (N_14602,N_14139,N_14039);
nor U14603 (N_14603,N_14268,N_14463);
nand U14604 (N_14604,N_14127,N_14405);
nand U14605 (N_14605,N_14002,N_14156);
nand U14606 (N_14606,N_14448,N_14102);
and U14607 (N_14607,N_14432,N_14161);
nand U14608 (N_14608,N_14133,N_14218);
and U14609 (N_14609,N_14396,N_14125);
xnor U14610 (N_14610,N_14368,N_14076);
nor U14611 (N_14611,N_14495,N_14435);
xor U14612 (N_14612,N_14103,N_14086);
or U14613 (N_14613,N_14207,N_14351);
nor U14614 (N_14614,N_14307,N_14144);
nand U14615 (N_14615,N_14450,N_14101);
xnor U14616 (N_14616,N_14222,N_14068);
or U14617 (N_14617,N_14004,N_14412);
xnor U14618 (N_14618,N_14330,N_14328);
or U14619 (N_14619,N_14489,N_14210);
nor U14620 (N_14620,N_14151,N_14242);
nor U14621 (N_14621,N_14118,N_14456);
and U14622 (N_14622,N_14227,N_14429);
nand U14623 (N_14623,N_14258,N_14026);
nor U14624 (N_14624,N_14425,N_14366);
nor U14625 (N_14625,N_14000,N_14280);
nor U14626 (N_14626,N_14439,N_14298);
nand U14627 (N_14627,N_14389,N_14485);
nor U14628 (N_14628,N_14434,N_14183);
nand U14629 (N_14629,N_14232,N_14310);
or U14630 (N_14630,N_14152,N_14446);
or U14631 (N_14631,N_14142,N_14167);
or U14632 (N_14632,N_14057,N_14237);
nand U14633 (N_14633,N_14419,N_14180);
nand U14634 (N_14634,N_14091,N_14481);
or U14635 (N_14635,N_14364,N_14197);
and U14636 (N_14636,N_14493,N_14006);
xor U14637 (N_14637,N_14077,N_14436);
nand U14638 (N_14638,N_14007,N_14196);
or U14639 (N_14639,N_14259,N_14457);
and U14640 (N_14640,N_14186,N_14486);
or U14641 (N_14641,N_14308,N_14421);
and U14642 (N_14642,N_14491,N_14315);
nor U14643 (N_14643,N_14290,N_14135);
nor U14644 (N_14644,N_14216,N_14423);
or U14645 (N_14645,N_14241,N_14049);
and U14646 (N_14646,N_14382,N_14267);
nand U14647 (N_14647,N_14147,N_14295);
nand U14648 (N_14648,N_14128,N_14276);
and U14649 (N_14649,N_14314,N_14209);
nand U14650 (N_14650,N_14372,N_14175);
and U14651 (N_14651,N_14440,N_14051);
nand U14652 (N_14652,N_14116,N_14195);
and U14653 (N_14653,N_14074,N_14204);
and U14654 (N_14654,N_14336,N_14260);
nor U14655 (N_14655,N_14213,N_14455);
nand U14656 (N_14656,N_14110,N_14397);
xor U14657 (N_14657,N_14063,N_14240);
xor U14658 (N_14658,N_14193,N_14176);
xor U14659 (N_14659,N_14296,N_14418);
nand U14660 (N_14660,N_14275,N_14353);
nand U14661 (N_14661,N_14462,N_14032);
or U14662 (N_14662,N_14014,N_14256);
or U14663 (N_14663,N_14045,N_14375);
xnor U14664 (N_14664,N_14494,N_14079);
nand U14665 (N_14665,N_14080,N_14126);
and U14666 (N_14666,N_14104,N_14479);
nor U14667 (N_14667,N_14459,N_14253);
xnor U14668 (N_14668,N_14445,N_14234);
and U14669 (N_14669,N_14354,N_14338);
and U14670 (N_14670,N_14306,N_14422);
nor U14671 (N_14671,N_14497,N_14179);
or U14672 (N_14672,N_14447,N_14106);
and U14673 (N_14673,N_14239,N_14452);
xnor U14674 (N_14674,N_14018,N_14206);
nand U14675 (N_14675,N_14094,N_14020);
or U14676 (N_14676,N_14365,N_14029);
and U14677 (N_14677,N_14327,N_14438);
xor U14678 (N_14678,N_14262,N_14089);
or U14679 (N_14679,N_14309,N_14348);
xnor U14680 (N_14680,N_14088,N_14248);
and U14681 (N_14681,N_14488,N_14177);
nand U14682 (N_14682,N_14231,N_14113);
and U14683 (N_14683,N_14427,N_14143);
nor U14684 (N_14684,N_14393,N_14304);
and U14685 (N_14685,N_14269,N_14441);
xor U14686 (N_14686,N_14297,N_14198);
and U14687 (N_14687,N_14174,N_14400);
nor U14688 (N_14688,N_14221,N_14302);
nand U14689 (N_14689,N_14228,N_14107);
nand U14690 (N_14690,N_14100,N_14162);
xnor U14691 (N_14691,N_14360,N_14033);
or U14692 (N_14692,N_14025,N_14036);
nand U14693 (N_14693,N_14092,N_14035);
xor U14694 (N_14694,N_14286,N_14202);
and U14695 (N_14695,N_14270,N_14064);
and U14696 (N_14696,N_14339,N_14320);
or U14697 (N_14697,N_14087,N_14392);
xnor U14698 (N_14698,N_14416,N_14361);
nor U14699 (N_14699,N_14069,N_14171);
or U14700 (N_14700,N_14058,N_14430);
nor U14701 (N_14701,N_14117,N_14433);
nor U14702 (N_14702,N_14169,N_14318);
nor U14703 (N_14703,N_14141,N_14381);
nor U14704 (N_14704,N_14053,N_14060);
or U14705 (N_14705,N_14254,N_14325);
and U14706 (N_14706,N_14492,N_14334);
nand U14707 (N_14707,N_14470,N_14070);
and U14708 (N_14708,N_14408,N_14071);
xor U14709 (N_14709,N_14490,N_14272);
nand U14710 (N_14710,N_14084,N_14410);
nor U14711 (N_14711,N_14230,N_14399);
xor U14712 (N_14712,N_14342,N_14048);
and U14713 (N_14713,N_14132,N_14474);
or U14714 (N_14714,N_14165,N_14265);
nand U14715 (N_14715,N_14225,N_14478);
xor U14716 (N_14716,N_14163,N_14134);
xor U14717 (N_14717,N_14499,N_14487);
and U14718 (N_14718,N_14083,N_14022);
or U14719 (N_14719,N_14205,N_14027);
nand U14720 (N_14720,N_14420,N_14345);
or U14721 (N_14721,N_14243,N_14252);
and U14722 (N_14722,N_14414,N_14201);
nand U14723 (N_14723,N_14283,N_14021);
or U14724 (N_14724,N_14081,N_14097);
nand U14725 (N_14725,N_14041,N_14466);
nor U14726 (N_14726,N_14335,N_14326);
or U14727 (N_14727,N_14093,N_14292);
and U14728 (N_14728,N_14212,N_14398);
xor U14729 (N_14729,N_14111,N_14251);
xor U14730 (N_14730,N_14282,N_14370);
nor U14731 (N_14731,N_14385,N_14170);
nand U14732 (N_14732,N_14105,N_14208);
nand U14733 (N_14733,N_14114,N_14321);
nor U14734 (N_14734,N_14344,N_14471);
and U14735 (N_14735,N_14271,N_14346);
and U14736 (N_14736,N_14019,N_14415);
xor U14737 (N_14737,N_14449,N_14050);
and U14738 (N_14738,N_14188,N_14028);
and U14739 (N_14739,N_14322,N_14291);
nor U14740 (N_14740,N_14480,N_14123);
xor U14741 (N_14741,N_14377,N_14379);
and U14742 (N_14742,N_14356,N_14442);
and U14743 (N_14743,N_14236,N_14431);
or U14744 (N_14744,N_14185,N_14477);
nand U14745 (N_14745,N_14305,N_14390);
xnor U14746 (N_14746,N_14154,N_14317);
and U14747 (N_14747,N_14461,N_14226);
xor U14748 (N_14748,N_14073,N_14223);
and U14749 (N_14749,N_14406,N_14146);
xor U14750 (N_14750,N_14158,N_14271);
or U14751 (N_14751,N_14397,N_14287);
nand U14752 (N_14752,N_14195,N_14445);
xnor U14753 (N_14753,N_14176,N_14466);
xor U14754 (N_14754,N_14109,N_14431);
nand U14755 (N_14755,N_14065,N_14227);
nor U14756 (N_14756,N_14069,N_14446);
nand U14757 (N_14757,N_14346,N_14289);
or U14758 (N_14758,N_14498,N_14224);
nand U14759 (N_14759,N_14028,N_14327);
and U14760 (N_14760,N_14100,N_14309);
or U14761 (N_14761,N_14482,N_14117);
and U14762 (N_14762,N_14050,N_14342);
nor U14763 (N_14763,N_14356,N_14365);
xnor U14764 (N_14764,N_14450,N_14093);
and U14765 (N_14765,N_14056,N_14035);
or U14766 (N_14766,N_14318,N_14141);
or U14767 (N_14767,N_14091,N_14154);
xnor U14768 (N_14768,N_14411,N_14492);
nand U14769 (N_14769,N_14227,N_14076);
nor U14770 (N_14770,N_14425,N_14126);
nand U14771 (N_14771,N_14331,N_14337);
nand U14772 (N_14772,N_14363,N_14216);
nor U14773 (N_14773,N_14104,N_14276);
xor U14774 (N_14774,N_14315,N_14125);
nand U14775 (N_14775,N_14238,N_14125);
nand U14776 (N_14776,N_14068,N_14496);
and U14777 (N_14777,N_14313,N_14094);
and U14778 (N_14778,N_14499,N_14231);
nand U14779 (N_14779,N_14452,N_14179);
nand U14780 (N_14780,N_14157,N_14480);
nor U14781 (N_14781,N_14066,N_14430);
or U14782 (N_14782,N_14004,N_14106);
or U14783 (N_14783,N_14354,N_14164);
and U14784 (N_14784,N_14390,N_14043);
or U14785 (N_14785,N_14135,N_14012);
and U14786 (N_14786,N_14425,N_14130);
nor U14787 (N_14787,N_14222,N_14452);
nor U14788 (N_14788,N_14246,N_14403);
xnor U14789 (N_14789,N_14414,N_14465);
xor U14790 (N_14790,N_14357,N_14209);
or U14791 (N_14791,N_14323,N_14067);
nor U14792 (N_14792,N_14392,N_14314);
nor U14793 (N_14793,N_14498,N_14360);
nand U14794 (N_14794,N_14150,N_14325);
nor U14795 (N_14795,N_14251,N_14486);
nand U14796 (N_14796,N_14122,N_14064);
and U14797 (N_14797,N_14253,N_14426);
or U14798 (N_14798,N_14494,N_14445);
and U14799 (N_14799,N_14456,N_14093);
nor U14800 (N_14800,N_14258,N_14389);
xnor U14801 (N_14801,N_14318,N_14480);
xnor U14802 (N_14802,N_14017,N_14144);
xnor U14803 (N_14803,N_14069,N_14434);
or U14804 (N_14804,N_14449,N_14485);
nor U14805 (N_14805,N_14414,N_14330);
xnor U14806 (N_14806,N_14239,N_14493);
nor U14807 (N_14807,N_14138,N_14435);
or U14808 (N_14808,N_14332,N_14373);
nor U14809 (N_14809,N_14270,N_14460);
nand U14810 (N_14810,N_14342,N_14305);
nand U14811 (N_14811,N_14417,N_14109);
and U14812 (N_14812,N_14080,N_14459);
nor U14813 (N_14813,N_14197,N_14094);
nor U14814 (N_14814,N_14161,N_14182);
xor U14815 (N_14815,N_14289,N_14275);
and U14816 (N_14816,N_14149,N_14447);
nand U14817 (N_14817,N_14472,N_14427);
nand U14818 (N_14818,N_14257,N_14083);
and U14819 (N_14819,N_14320,N_14297);
nand U14820 (N_14820,N_14356,N_14378);
nor U14821 (N_14821,N_14036,N_14216);
nor U14822 (N_14822,N_14024,N_14061);
xor U14823 (N_14823,N_14266,N_14386);
or U14824 (N_14824,N_14056,N_14069);
or U14825 (N_14825,N_14001,N_14247);
nor U14826 (N_14826,N_14341,N_14401);
nor U14827 (N_14827,N_14196,N_14337);
and U14828 (N_14828,N_14082,N_14471);
xnor U14829 (N_14829,N_14208,N_14351);
or U14830 (N_14830,N_14292,N_14320);
or U14831 (N_14831,N_14207,N_14283);
nor U14832 (N_14832,N_14411,N_14015);
nand U14833 (N_14833,N_14142,N_14308);
xor U14834 (N_14834,N_14463,N_14038);
xnor U14835 (N_14835,N_14320,N_14232);
nand U14836 (N_14836,N_14239,N_14344);
xor U14837 (N_14837,N_14292,N_14147);
nor U14838 (N_14838,N_14411,N_14152);
nor U14839 (N_14839,N_14407,N_14213);
nand U14840 (N_14840,N_14009,N_14399);
nor U14841 (N_14841,N_14159,N_14495);
nand U14842 (N_14842,N_14013,N_14246);
and U14843 (N_14843,N_14337,N_14183);
nand U14844 (N_14844,N_14306,N_14375);
and U14845 (N_14845,N_14221,N_14443);
nor U14846 (N_14846,N_14253,N_14220);
xor U14847 (N_14847,N_14407,N_14484);
or U14848 (N_14848,N_14038,N_14126);
or U14849 (N_14849,N_14484,N_14340);
nand U14850 (N_14850,N_14077,N_14255);
nand U14851 (N_14851,N_14471,N_14049);
or U14852 (N_14852,N_14236,N_14039);
and U14853 (N_14853,N_14015,N_14122);
nand U14854 (N_14854,N_14468,N_14298);
nand U14855 (N_14855,N_14224,N_14063);
nand U14856 (N_14856,N_14274,N_14265);
nor U14857 (N_14857,N_14425,N_14463);
nor U14858 (N_14858,N_14158,N_14399);
nand U14859 (N_14859,N_14326,N_14142);
nand U14860 (N_14860,N_14091,N_14181);
nand U14861 (N_14861,N_14378,N_14237);
nand U14862 (N_14862,N_14163,N_14226);
nor U14863 (N_14863,N_14225,N_14244);
nand U14864 (N_14864,N_14478,N_14096);
nand U14865 (N_14865,N_14025,N_14379);
or U14866 (N_14866,N_14368,N_14260);
nor U14867 (N_14867,N_14496,N_14439);
and U14868 (N_14868,N_14424,N_14374);
and U14869 (N_14869,N_14250,N_14258);
nor U14870 (N_14870,N_14134,N_14451);
and U14871 (N_14871,N_14085,N_14108);
or U14872 (N_14872,N_14302,N_14232);
or U14873 (N_14873,N_14395,N_14248);
xnor U14874 (N_14874,N_14202,N_14490);
nor U14875 (N_14875,N_14370,N_14266);
nand U14876 (N_14876,N_14113,N_14238);
xor U14877 (N_14877,N_14305,N_14007);
or U14878 (N_14878,N_14109,N_14122);
nor U14879 (N_14879,N_14266,N_14081);
nand U14880 (N_14880,N_14479,N_14189);
and U14881 (N_14881,N_14104,N_14382);
and U14882 (N_14882,N_14253,N_14339);
nor U14883 (N_14883,N_14266,N_14046);
or U14884 (N_14884,N_14335,N_14304);
xnor U14885 (N_14885,N_14004,N_14195);
nand U14886 (N_14886,N_14268,N_14189);
nand U14887 (N_14887,N_14247,N_14168);
nor U14888 (N_14888,N_14068,N_14307);
nand U14889 (N_14889,N_14070,N_14451);
and U14890 (N_14890,N_14461,N_14435);
nor U14891 (N_14891,N_14453,N_14071);
and U14892 (N_14892,N_14154,N_14277);
xnor U14893 (N_14893,N_14191,N_14437);
or U14894 (N_14894,N_14064,N_14460);
nor U14895 (N_14895,N_14280,N_14131);
or U14896 (N_14896,N_14440,N_14115);
nor U14897 (N_14897,N_14251,N_14459);
or U14898 (N_14898,N_14056,N_14020);
or U14899 (N_14899,N_14472,N_14460);
nor U14900 (N_14900,N_14304,N_14055);
xnor U14901 (N_14901,N_14057,N_14368);
nand U14902 (N_14902,N_14263,N_14230);
and U14903 (N_14903,N_14022,N_14115);
or U14904 (N_14904,N_14063,N_14236);
xor U14905 (N_14905,N_14268,N_14158);
or U14906 (N_14906,N_14284,N_14164);
and U14907 (N_14907,N_14447,N_14058);
and U14908 (N_14908,N_14129,N_14207);
and U14909 (N_14909,N_14101,N_14073);
or U14910 (N_14910,N_14146,N_14178);
nor U14911 (N_14911,N_14296,N_14166);
nor U14912 (N_14912,N_14138,N_14419);
nor U14913 (N_14913,N_14352,N_14036);
and U14914 (N_14914,N_14378,N_14007);
nor U14915 (N_14915,N_14180,N_14469);
and U14916 (N_14916,N_14332,N_14226);
or U14917 (N_14917,N_14029,N_14057);
nor U14918 (N_14918,N_14370,N_14397);
nand U14919 (N_14919,N_14332,N_14063);
and U14920 (N_14920,N_14210,N_14190);
nor U14921 (N_14921,N_14077,N_14356);
and U14922 (N_14922,N_14493,N_14213);
and U14923 (N_14923,N_14096,N_14246);
nand U14924 (N_14924,N_14069,N_14124);
or U14925 (N_14925,N_14402,N_14158);
and U14926 (N_14926,N_14377,N_14069);
or U14927 (N_14927,N_14333,N_14008);
nand U14928 (N_14928,N_14347,N_14473);
or U14929 (N_14929,N_14275,N_14003);
or U14930 (N_14930,N_14215,N_14387);
and U14931 (N_14931,N_14466,N_14129);
and U14932 (N_14932,N_14189,N_14423);
nor U14933 (N_14933,N_14173,N_14321);
and U14934 (N_14934,N_14348,N_14283);
and U14935 (N_14935,N_14289,N_14070);
or U14936 (N_14936,N_14127,N_14403);
and U14937 (N_14937,N_14024,N_14115);
or U14938 (N_14938,N_14001,N_14180);
nor U14939 (N_14939,N_14391,N_14496);
nand U14940 (N_14940,N_14360,N_14184);
nor U14941 (N_14941,N_14055,N_14470);
and U14942 (N_14942,N_14051,N_14494);
nor U14943 (N_14943,N_14223,N_14278);
nor U14944 (N_14944,N_14332,N_14108);
nor U14945 (N_14945,N_14312,N_14205);
or U14946 (N_14946,N_14078,N_14261);
and U14947 (N_14947,N_14249,N_14396);
nand U14948 (N_14948,N_14018,N_14204);
xor U14949 (N_14949,N_14383,N_14295);
and U14950 (N_14950,N_14272,N_14025);
or U14951 (N_14951,N_14414,N_14074);
and U14952 (N_14952,N_14167,N_14169);
nand U14953 (N_14953,N_14316,N_14300);
and U14954 (N_14954,N_14140,N_14398);
nor U14955 (N_14955,N_14034,N_14180);
nand U14956 (N_14956,N_14166,N_14339);
nand U14957 (N_14957,N_14004,N_14140);
nor U14958 (N_14958,N_14176,N_14037);
and U14959 (N_14959,N_14426,N_14110);
nor U14960 (N_14960,N_14254,N_14371);
or U14961 (N_14961,N_14458,N_14429);
xnor U14962 (N_14962,N_14308,N_14320);
nand U14963 (N_14963,N_14108,N_14196);
and U14964 (N_14964,N_14263,N_14238);
nor U14965 (N_14965,N_14414,N_14458);
nor U14966 (N_14966,N_14354,N_14043);
and U14967 (N_14967,N_14224,N_14020);
and U14968 (N_14968,N_14297,N_14106);
nand U14969 (N_14969,N_14181,N_14297);
xnor U14970 (N_14970,N_14242,N_14108);
nor U14971 (N_14971,N_14163,N_14312);
or U14972 (N_14972,N_14327,N_14271);
nand U14973 (N_14973,N_14391,N_14481);
and U14974 (N_14974,N_14214,N_14156);
or U14975 (N_14975,N_14210,N_14476);
xnor U14976 (N_14976,N_14434,N_14399);
xnor U14977 (N_14977,N_14008,N_14021);
and U14978 (N_14978,N_14450,N_14102);
xor U14979 (N_14979,N_14359,N_14488);
or U14980 (N_14980,N_14461,N_14381);
nand U14981 (N_14981,N_14219,N_14011);
nor U14982 (N_14982,N_14415,N_14043);
xor U14983 (N_14983,N_14494,N_14107);
and U14984 (N_14984,N_14204,N_14001);
nor U14985 (N_14985,N_14386,N_14130);
nor U14986 (N_14986,N_14349,N_14338);
or U14987 (N_14987,N_14011,N_14036);
nor U14988 (N_14988,N_14153,N_14276);
nand U14989 (N_14989,N_14391,N_14024);
and U14990 (N_14990,N_14268,N_14078);
nand U14991 (N_14991,N_14454,N_14468);
nand U14992 (N_14992,N_14483,N_14267);
and U14993 (N_14993,N_14388,N_14441);
nor U14994 (N_14994,N_14127,N_14074);
nand U14995 (N_14995,N_14000,N_14055);
and U14996 (N_14996,N_14054,N_14489);
nand U14997 (N_14997,N_14053,N_14380);
nand U14998 (N_14998,N_14066,N_14319);
and U14999 (N_14999,N_14277,N_14266);
or UO_0 (O_0,N_14874,N_14899);
nor UO_1 (O_1,N_14764,N_14624);
nand UO_2 (O_2,N_14864,N_14511);
or UO_3 (O_3,N_14691,N_14596);
or UO_4 (O_4,N_14715,N_14922);
and UO_5 (O_5,N_14750,N_14801);
nor UO_6 (O_6,N_14870,N_14723);
xor UO_7 (O_7,N_14600,N_14552);
xnor UO_8 (O_8,N_14857,N_14943);
or UO_9 (O_9,N_14818,N_14805);
xnor UO_10 (O_10,N_14655,N_14911);
nor UO_11 (O_11,N_14665,N_14959);
xor UO_12 (O_12,N_14788,N_14522);
and UO_13 (O_13,N_14734,N_14553);
nor UO_14 (O_14,N_14840,N_14677);
nand UO_15 (O_15,N_14831,N_14937);
nor UO_16 (O_16,N_14848,N_14674);
xor UO_17 (O_17,N_14666,N_14509);
or UO_18 (O_18,N_14693,N_14521);
nor UO_19 (O_19,N_14730,N_14646);
xnor UO_20 (O_20,N_14850,N_14921);
nand UO_21 (O_21,N_14952,N_14751);
or UO_22 (O_22,N_14574,N_14851);
nor UO_23 (O_23,N_14737,N_14664);
nand UO_24 (O_24,N_14705,N_14780);
and UO_25 (O_25,N_14955,N_14580);
xor UO_26 (O_26,N_14732,N_14603);
or UO_27 (O_27,N_14930,N_14692);
nand UO_28 (O_28,N_14740,N_14829);
nand UO_29 (O_29,N_14944,N_14786);
and UO_30 (O_30,N_14636,N_14775);
or UO_31 (O_31,N_14625,N_14556);
nor UO_32 (O_32,N_14961,N_14939);
xnor UO_33 (O_33,N_14929,N_14935);
or UO_34 (O_34,N_14942,N_14814);
nor UO_35 (O_35,N_14611,N_14932);
nand UO_36 (O_36,N_14837,N_14990);
nor UO_37 (O_37,N_14815,N_14680);
or UO_38 (O_38,N_14709,N_14771);
and UO_39 (O_39,N_14845,N_14754);
and UO_40 (O_40,N_14769,N_14650);
and UO_41 (O_41,N_14977,N_14546);
nand UO_42 (O_42,N_14523,N_14773);
xor UO_43 (O_43,N_14638,N_14689);
nor UO_44 (O_44,N_14872,N_14900);
nor UO_45 (O_45,N_14889,N_14895);
nor UO_46 (O_46,N_14980,N_14663);
and UO_47 (O_47,N_14946,N_14909);
nor UO_48 (O_48,N_14746,N_14639);
or UO_49 (O_49,N_14720,N_14513);
nand UO_50 (O_50,N_14634,N_14605);
nor UO_51 (O_51,N_14886,N_14566);
or UO_52 (O_52,N_14994,N_14984);
or UO_53 (O_53,N_14865,N_14936);
or UO_54 (O_54,N_14948,N_14998);
or UO_55 (O_55,N_14954,N_14686);
or UO_56 (O_56,N_14630,N_14969);
nand UO_57 (O_57,N_14827,N_14949);
nor UO_58 (O_58,N_14783,N_14915);
nand UO_59 (O_59,N_14675,N_14687);
nand UO_60 (O_60,N_14503,N_14767);
nor UO_61 (O_61,N_14669,N_14970);
nor UO_62 (O_62,N_14627,N_14789);
and UO_63 (O_63,N_14888,N_14880);
and UO_64 (O_64,N_14619,N_14579);
or UO_65 (O_65,N_14537,N_14867);
or UO_66 (O_66,N_14965,N_14644);
xor UO_67 (O_67,N_14914,N_14702);
or UO_68 (O_68,N_14718,N_14525);
and UO_69 (O_69,N_14933,N_14819);
nor UO_70 (O_70,N_14759,N_14571);
and UO_71 (O_71,N_14685,N_14793);
and UO_72 (O_72,N_14587,N_14810);
or UO_73 (O_73,N_14903,N_14995);
or UO_74 (O_74,N_14877,N_14791);
or UO_75 (O_75,N_14719,N_14821);
nand UO_76 (O_76,N_14881,N_14500);
or UO_77 (O_77,N_14621,N_14530);
and UO_78 (O_78,N_14968,N_14753);
or UO_79 (O_79,N_14904,N_14517);
xnor UO_80 (O_80,N_14802,N_14755);
and UO_81 (O_81,N_14502,N_14906);
and UO_82 (O_82,N_14863,N_14878);
and UO_83 (O_83,N_14510,N_14927);
and UO_84 (O_84,N_14741,N_14823);
xnor UO_85 (O_85,N_14862,N_14806);
or UO_86 (O_86,N_14799,N_14861);
nor UO_87 (O_87,N_14999,N_14598);
and UO_88 (O_88,N_14631,N_14572);
and UO_89 (O_89,N_14544,N_14811);
nand UO_90 (O_90,N_14704,N_14738);
nor UO_91 (O_91,N_14795,N_14698);
and UO_92 (O_92,N_14873,N_14817);
and UO_93 (O_93,N_14992,N_14924);
xor UO_94 (O_94,N_14981,N_14782);
nor UO_95 (O_95,N_14635,N_14642);
nand UO_96 (O_96,N_14550,N_14825);
xnor UO_97 (O_97,N_14830,N_14822);
nor UO_98 (O_98,N_14804,N_14582);
xor UO_99 (O_99,N_14833,N_14604);
nand UO_100 (O_100,N_14542,N_14519);
nand UO_101 (O_101,N_14743,N_14551);
or UO_102 (O_102,N_14694,N_14528);
and UO_103 (O_103,N_14890,N_14725);
and UO_104 (O_104,N_14926,N_14756);
nor UO_105 (O_105,N_14684,N_14671);
xnor UO_106 (O_106,N_14616,N_14785);
xor UO_107 (O_107,N_14853,N_14947);
xor UO_108 (O_108,N_14562,N_14520);
and UO_109 (O_109,N_14991,N_14560);
nor UO_110 (O_110,N_14547,N_14722);
xnor UO_111 (O_111,N_14856,N_14905);
nor UO_112 (O_112,N_14975,N_14748);
xnor UO_113 (O_113,N_14956,N_14798);
nor UO_114 (O_114,N_14727,N_14606);
and UO_115 (O_115,N_14728,N_14855);
or UO_116 (O_116,N_14554,N_14752);
xnor UO_117 (O_117,N_14765,N_14974);
nor UO_118 (O_118,N_14613,N_14539);
xnor UO_119 (O_119,N_14983,N_14907);
or UO_120 (O_120,N_14586,N_14892);
or UO_121 (O_121,N_14614,N_14957);
and UO_122 (O_122,N_14706,N_14920);
xnor UO_123 (O_123,N_14910,N_14667);
nand UO_124 (O_124,N_14569,N_14683);
xor UO_125 (O_125,N_14592,N_14648);
or UO_126 (O_126,N_14717,N_14731);
xnor UO_127 (O_127,N_14615,N_14893);
and UO_128 (O_128,N_14570,N_14966);
or UO_129 (O_129,N_14504,N_14708);
xnor UO_130 (O_130,N_14658,N_14971);
xnor UO_131 (O_131,N_14918,N_14854);
nand UO_132 (O_132,N_14963,N_14637);
nor UO_133 (O_133,N_14938,N_14701);
nor UO_134 (O_134,N_14839,N_14555);
or UO_135 (O_135,N_14973,N_14656);
or UO_136 (O_136,N_14941,N_14897);
and UO_137 (O_137,N_14860,N_14548);
nand UO_138 (O_138,N_14640,N_14797);
nand UO_139 (O_139,N_14573,N_14896);
nor UO_140 (O_140,N_14978,N_14776);
xor UO_141 (O_141,N_14826,N_14505);
nand UO_142 (O_142,N_14527,N_14535);
nor UO_143 (O_143,N_14770,N_14919);
xnor UO_144 (O_144,N_14690,N_14835);
or UO_145 (O_145,N_14997,N_14828);
xnor UO_146 (O_146,N_14917,N_14761);
or UO_147 (O_147,N_14866,N_14545);
nand UO_148 (O_148,N_14711,N_14713);
nor UO_149 (O_149,N_14996,N_14747);
nand UO_150 (O_150,N_14898,N_14678);
and UO_151 (O_151,N_14612,N_14790);
nor UO_152 (O_152,N_14846,N_14697);
or UO_153 (O_153,N_14659,N_14532);
and UO_154 (O_154,N_14875,N_14876);
nor UO_155 (O_155,N_14726,N_14859);
or UO_156 (O_156,N_14595,N_14774);
or UO_157 (O_157,N_14588,N_14602);
nand UO_158 (O_158,N_14882,N_14724);
and UO_159 (O_159,N_14584,N_14591);
or UO_160 (O_160,N_14673,N_14784);
nor UO_161 (O_161,N_14808,N_14565);
xor UO_162 (O_162,N_14609,N_14703);
xor UO_163 (O_163,N_14960,N_14832);
xnor UO_164 (O_164,N_14838,N_14660);
and UO_165 (O_165,N_14950,N_14707);
and UO_166 (O_166,N_14916,N_14958);
or UO_167 (O_167,N_14661,N_14883);
nor UO_168 (O_168,N_14508,N_14651);
nor UO_169 (O_169,N_14590,N_14601);
and UO_170 (O_170,N_14643,N_14986);
nand UO_171 (O_171,N_14581,N_14559);
xor UO_172 (O_172,N_14894,N_14824);
nor UO_173 (O_173,N_14617,N_14836);
nor UO_174 (O_174,N_14744,N_14816);
or UO_175 (O_175,N_14629,N_14695);
xnor UO_176 (O_176,N_14714,N_14632);
and UO_177 (O_177,N_14979,N_14594);
nor UO_178 (O_178,N_14951,N_14514);
nand UO_179 (O_179,N_14803,N_14645);
xor UO_180 (O_180,N_14989,N_14649);
or UO_181 (O_181,N_14869,N_14902);
nor UO_182 (O_182,N_14543,N_14608);
nor UO_183 (O_183,N_14676,N_14820);
xnor UO_184 (O_184,N_14501,N_14540);
nand UO_185 (O_185,N_14976,N_14800);
nor UO_186 (O_186,N_14516,N_14928);
and UO_187 (O_187,N_14842,N_14779);
or UO_188 (O_188,N_14760,N_14716);
or UO_189 (O_189,N_14578,N_14729);
xnor UO_190 (O_190,N_14597,N_14618);
and UO_191 (O_191,N_14940,N_14534);
nand UO_192 (O_192,N_14945,N_14538);
nor UO_193 (O_193,N_14506,N_14735);
or UO_194 (O_194,N_14626,N_14593);
or UO_195 (O_195,N_14982,N_14852);
nand UO_196 (O_196,N_14901,N_14657);
or UO_197 (O_197,N_14699,N_14662);
and UO_198 (O_198,N_14813,N_14844);
nand UO_199 (O_199,N_14843,N_14583);
and UO_200 (O_200,N_14879,N_14633);
nor UO_201 (O_201,N_14515,N_14536);
xor UO_202 (O_202,N_14796,N_14622);
and UO_203 (O_203,N_14512,N_14988);
nand UO_204 (O_204,N_14868,N_14589);
and UO_205 (O_205,N_14847,N_14672);
and UO_206 (O_206,N_14964,N_14912);
and UO_207 (O_207,N_14858,N_14762);
nor UO_208 (O_208,N_14576,N_14529);
xnor UO_209 (O_209,N_14654,N_14679);
nor UO_210 (O_210,N_14871,N_14777);
and UO_211 (O_211,N_14891,N_14757);
or UO_212 (O_212,N_14841,N_14620);
nand UO_213 (O_213,N_14524,N_14768);
nor UO_214 (O_214,N_14577,N_14681);
xor UO_215 (O_215,N_14787,N_14668);
xnor UO_216 (O_216,N_14781,N_14567);
nand UO_217 (O_217,N_14607,N_14908);
or UO_218 (O_218,N_14647,N_14733);
and UO_219 (O_219,N_14533,N_14628);
xnor UO_220 (O_220,N_14794,N_14962);
xnor UO_221 (O_221,N_14561,N_14558);
xor UO_222 (O_222,N_14834,N_14507);
and UO_223 (O_223,N_14652,N_14531);
nand UO_224 (O_224,N_14541,N_14967);
or UO_225 (O_225,N_14623,N_14688);
xnor UO_226 (O_226,N_14549,N_14526);
or UO_227 (O_227,N_14925,N_14985);
or UO_228 (O_228,N_14884,N_14758);
and UO_229 (O_229,N_14653,N_14807);
xnor UO_230 (O_230,N_14696,N_14778);
and UO_231 (O_231,N_14993,N_14742);
xnor UO_232 (O_232,N_14766,N_14953);
and UO_233 (O_233,N_14931,N_14670);
nand UO_234 (O_234,N_14849,N_14568);
xnor UO_235 (O_235,N_14518,N_14812);
nor UO_236 (O_236,N_14923,N_14739);
and UO_237 (O_237,N_14610,N_14682);
nand UO_238 (O_238,N_14763,N_14972);
nand UO_239 (O_239,N_14745,N_14585);
nor UO_240 (O_240,N_14557,N_14721);
nand UO_241 (O_241,N_14887,N_14809);
nand UO_242 (O_242,N_14987,N_14641);
xor UO_243 (O_243,N_14563,N_14700);
xnor UO_244 (O_244,N_14885,N_14575);
nand UO_245 (O_245,N_14772,N_14913);
or UO_246 (O_246,N_14564,N_14792);
nand UO_247 (O_247,N_14712,N_14599);
and UO_248 (O_248,N_14749,N_14736);
and UO_249 (O_249,N_14934,N_14710);
xor UO_250 (O_250,N_14564,N_14830);
or UO_251 (O_251,N_14885,N_14900);
xnor UO_252 (O_252,N_14614,N_14846);
or UO_253 (O_253,N_14905,N_14690);
xor UO_254 (O_254,N_14511,N_14779);
or UO_255 (O_255,N_14545,N_14576);
xnor UO_256 (O_256,N_14631,N_14687);
or UO_257 (O_257,N_14868,N_14984);
nand UO_258 (O_258,N_14654,N_14778);
nor UO_259 (O_259,N_14926,N_14976);
nor UO_260 (O_260,N_14807,N_14594);
nor UO_261 (O_261,N_14799,N_14813);
and UO_262 (O_262,N_14602,N_14728);
nor UO_263 (O_263,N_14839,N_14548);
and UO_264 (O_264,N_14578,N_14500);
nor UO_265 (O_265,N_14602,N_14930);
nand UO_266 (O_266,N_14834,N_14843);
and UO_267 (O_267,N_14867,N_14941);
or UO_268 (O_268,N_14644,N_14563);
xor UO_269 (O_269,N_14517,N_14549);
nand UO_270 (O_270,N_14632,N_14839);
xnor UO_271 (O_271,N_14932,N_14555);
nand UO_272 (O_272,N_14995,N_14875);
xor UO_273 (O_273,N_14827,N_14593);
xor UO_274 (O_274,N_14933,N_14838);
and UO_275 (O_275,N_14777,N_14790);
nor UO_276 (O_276,N_14695,N_14801);
or UO_277 (O_277,N_14773,N_14653);
and UO_278 (O_278,N_14576,N_14632);
or UO_279 (O_279,N_14540,N_14629);
or UO_280 (O_280,N_14552,N_14533);
or UO_281 (O_281,N_14768,N_14979);
xor UO_282 (O_282,N_14536,N_14514);
nand UO_283 (O_283,N_14698,N_14893);
or UO_284 (O_284,N_14593,N_14656);
and UO_285 (O_285,N_14522,N_14565);
nor UO_286 (O_286,N_14692,N_14954);
nor UO_287 (O_287,N_14961,N_14517);
nand UO_288 (O_288,N_14617,N_14613);
or UO_289 (O_289,N_14647,N_14804);
or UO_290 (O_290,N_14923,N_14989);
and UO_291 (O_291,N_14720,N_14676);
or UO_292 (O_292,N_14580,N_14917);
nand UO_293 (O_293,N_14611,N_14822);
and UO_294 (O_294,N_14518,N_14981);
nand UO_295 (O_295,N_14998,N_14641);
nor UO_296 (O_296,N_14695,N_14703);
or UO_297 (O_297,N_14681,N_14593);
or UO_298 (O_298,N_14679,N_14519);
xnor UO_299 (O_299,N_14859,N_14576);
nand UO_300 (O_300,N_14599,N_14618);
or UO_301 (O_301,N_14758,N_14685);
nand UO_302 (O_302,N_14760,N_14723);
and UO_303 (O_303,N_14694,N_14826);
or UO_304 (O_304,N_14688,N_14799);
xnor UO_305 (O_305,N_14679,N_14664);
or UO_306 (O_306,N_14996,N_14500);
xnor UO_307 (O_307,N_14899,N_14945);
nand UO_308 (O_308,N_14766,N_14973);
xor UO_309 (O_309,N_14689,N_14708);
nor UO_310 (O_310,N_14603,N_14970);
or UO_311 (O_311,N_14568,N_14617);
nor UO_312 (O_312,N_14515,N_14537);
or UO_313 (O_313,N_14990,N_14578);
nand UO_314 (O_314,N_14806,N_14932);
nand UO_315 (O_315,N_14518,N_14544);
and UO_316 (O_316,N_14701,N_14959);
xnor UO_317 (O_317,N_14770,N_14772);
and UO_318 (O_318,N_14860,N_14715);
xor UO_319 (O_319,N_14886,N_14877);
xor UO_320 (O_320,N_14798,N_14764);
xor UO_321 (O_321,N_14890,N_14805);
or UO_322 (O_322,N_14589,N_14997);
xnor UO_323 (O_323,N_14528,N_14896);
nand UO_324 (O_324,N_14855,N_14506);
or UO_325 (O_325,N_14726,N_14548);
nor UO_326 (O_326,N_14951,N_14714);
nand UO_327 (O_327,N_14957,N_14620);
nand UO_328 (O_328,N_14983,N_14641);
or UO_329 (O_329,N_14736,N_14591);
nor UO_330 (O_330,N_14786,N_14937);
or UO_331 (O_331,N_14613,N_14656);
xor UO_332 (O_332,N_14765,N_14877);
nor UO_333 (O_333,N_14889,N_14738);
xor UO_334 (O_334,N_14764,N_14828);
and UO_335 (O_335,N_14816,N_14560);
and UO_336 (O_336,N_14938,N_14812);
nand UO_337 (O_337,N_14862,N_14637);
and UO_338 (O_338,N_14986,N_14832);
and UO_339 (O_339,N_14688,N_14900);
nor UO_340 (O_340,N_14957,N_14596);
nand UO_341 (O_341,N_14973,N_14546);
or UO_342 (O_342,N_14744,N_14686);
xor UO_343 (O_343,N_14585,N_14642);
and UO_344 (O_344,N_14606,N_14674);
and UO_345 (O_345,N_14685,N_14958);
or UO_346 (O_346,N_14783,N_14751);
and UO_347 (O_347,N_14667,N_14894);
or UO_348 (O_348,N_14862,N_14957);
nand UO_349 (O_349,N_14785,N_14929);
nor UO_350 (O_350,N_14826,N_14730);
nand UO_351 (O_351,N_14954,N_14614);
or UO_352 (O_352,N_14543,N_14663);
nor UO_353 (O_353,N_14575,N_14856);
and UO_354 (O_354,N_14561,N_14914);
and UO_355 (O_355,N_14742,N_14703);
nand UO_356 (O_356,N_14586,N_14751);
nand UO_357 (O_357,N_14686,N_14982);
or UO_358 (O_358,N_14797,N_14644);
xor UO_359 (O_359,N_14732,N_14546);
xnor UO_360 (O_360,N_14587,N_14814);
or UO_361 (O_361,N_14639,N_14691);
xnor UO_362 (O_362,N_14971,N_14859);
xnor UO_363 (O_363,N_14971,N_14544);
nor UO_364 (O_364,N_14855,N_14842);
nor UO_365 (O_365,N_14700,N_14620);
nand UO_366 (O_366,N_14908,N_14599);
nand UO_367 (O_367,N_14639,N_14690);
nand UO_368 (O_368,N_14749,N_14945);
xor UO_369 (O_369,N_14762,N_14871);
or UO_370 (O_370,N_14781,N_14836);
and UO_371 (O_371,N_14605,N_14756);
nor UO_372 (O_372,N_14571,N_14862);
nand UO_373 (O_373,N_14748,N_14805);
nor UO_374 (O_374,N_14696,N_14557);
and UO_375 (O_375,N_14929,N_14703);
xor UO_376 (O_376,N_14595,N_14855);
nand UO_377 (O_377,N_14670,N_14885);
and UO_378 (O_378,N_14906,N_14817);
nor UO_379 (O_379,N_14991,N_14903);
nor UO_380 (O_380,N_14717,N_14558);
xor UO_381 (O_381,N_14697,N_14512);
nor UO_382 (O_382,N_14674,N_14697);
and UO_383 (O_383,N_14648,N_14562);
and UO_384 (O_384,N_14891,N_14572);
and UO_385 (O_385,N_14683,N_14904);
xor UO_386 (O_386,N_14866,N_14588);
or UO_387 (O_387,N_14913,N_14920);
nor UO_388 (O_388,N_14610,N_14690);
nor UO_389 (O_389,N_14613,N_14926);
and UO_390 (O_390,N_14857,N_14936);
xor UO_391 (O_391,N_14852,N_14689);
or UO_392 (O_392,N_14650,N_14614);
nand UO_393 (O_393,N_14649,N_14868);
and UO_394 (O_394,N_14791,N_14958);
nand UO_395 (O_395,N_14908,N_14857);
and UO_396 (O_396,N_14876,N_14551);
and UO_397 (O_397,N_14522,N_14732);
nand UO_398 (O_398,N_14740,N_14940);
nand UO_399 (O_399,N_14715,N_14664);
and UO_400 (O_400,N_14657,N_14875);
or UO_401 (O_401,N_14849,N_14872);
or UO_402 (O_402,N_14643,N_14733);
xnor UO_403 (O_403,N_14654,N_14707);
nor UO_404 (O_404,N_14539,N_14773);
or UO_405 (O_405,N_14841,N_14763);
nand UO_406 (O_406,N_14892,N_14701);
nor UO_407 (O_407,N_14806,N_14569);
xor UO_408 (O_408,N_14814,N_14708);
nand UO_409 (O_409,N_14759,N_14799);
nor UO_410 (O_410,N_14810,N_14881);
xnor UO_411 (O_411,N_14838,N_14669);
nand UO_412 (O_412,N_14763,N_14888);
nand UO_413 (O_413,N_14949,N_14914);
nor UO_414 (O_414,N_14760,N_14815);
nor UO_415 (O_415,N_14582,N_14624);
xor UO_416 (O_416,N_14899,N_14744);
nor UO_417 (O_417,N_14504,N_14836);
and UO_418 (O_418,N_14606,N_14841);
and UO_419 (O_419,N_14657,N_14601);
nor UO_420 (O_420,N_14938,N_14829);
xor UO_421 (O_421,N_14537,N_14779);
nand UO_422 (O_422,N_14740,N_14790);
nor UO_423 (O_423,N_14560,N_14577);
and UO_424 (O_424,N_14517,N_14604);
xnor UO_425 (O_425,N_14648,N_14528);
or UO_426 (O_426,N_14649,N_14766);
or UO_427 (O_427,N_14712,N_14927);
nor UO_428 (O_428,N_14665,N_14800);
xnor UO_429 (O_429,N_14617,N_14913);
or UO_430 (O_430,N_14623,N_14744);
nor UO_431 (O_431,N_14723,N_14565);
xor UO_432 (O_432,N_14579,N_14627);
or UO_433 (O_433,N_14514,N_14879);
and UO_434 (O_434,N_14638,N_14962);
nor UO_435 (O_435,N_14854,N_14921);
nor UO_436 (O_436,N_14890,N_14664);
nand UO_437 (O_437,N_14768,N_14857);
nand UO_438 (O_438,N_14717,N_14865);
nand UO_439 (O_439,N_14641,N_14740);
and UO_440 (O_440,N_14628,N_14637);
nor UO_441 (O_441,N_14693,N_14695);
nor UO_442 (O_442,N_14984,N_14833);
nor UO_443 (O_443,N_14864,N_14805);
nor UO_444 (O_444,N_14765,N_14951);
and UO_445 (O_445,N_14980,N_14876);
xor UO_446 (O_446,N_14813,N_14556);
and UO_447 (O_447,N_14546,N_14527);
nand UO_448 (O_448,N_14912,N_14836);
or UO_449 (O_449,N_14988,N_14869);
nand UO_450 (O_450,N_14657,N_14980);
nor UO_451 (O_451,N_14905,N_14614);
nor UO_452 (O_452,N_14679,N_14834);
nor UO_453 (O_453,N_14606,N_14987);
nand UO_454 (O_454,N_14605,N_14597);
xnor UO_455 (O_455,N_14564,N_14736);
and UO_456 (O_456,N_14564,N_14846);
nor UO_457 (O_457,N_14925,N_14730);
or UO_458 (O_458,N_14690,N_14724);
or UO_459 (O_459,N_14594,N_14928);
or UO_460 (O_460,N_14785,N_14926);
and UO_461 (O_461,N_14685,N_14586);
or UO_462 (O_462,N_14574,N_14917);
and UO_463 (O_463,N_14914,N_14840);
xnor UO_464 (O_464,N_14945,N_14962);
and UO_465 (O_465,N_14751,N_14565);
xnor UO_466 (O_466,N_14757,N_14614);
or UO_467 (O_467,N_14753,N_14630);
or UO_468 (O_468,N_14787,N_14580);
xor UO_469 (O_469,N_14704,N_14625);
or UO_470 (O_470,N_14993,N_14584);
or UO_471 (O_471,N_14584,N_14831);
nand UO_472 (O_472,N_14943,N_14744);
nand UO_473 (O_473,N_14836,N_14971);
and UO_474 (O_474,N_14748,N_14673);
xnor UO_475 (O_475,N_14508,N_14704);
nand UO_476 (O_476,N_14942,N_14534);
xor UO_477 (O_477,N_14806,N_14741);
xor UO_478 (O_478,N_14946,N_14567);
or UO_479 (O_479,N_14954,N_14947);
and UO_480 (O_480,N_14631,N_14534);
or UO_481 (O_481,N_14559,N_14675);
xnor UO_482 (O_482,N_14934,N_14807);
and UO_483 (O_483,N_14882,N_14944);
nor UO_484 (O_484,N_14905,N_14706);
or UO_485 (O_485,N_14876,N_14538);
and UO_486 (O_486,N_14858,N_14802);
xnor UO_487 (O_487,N_14518,N_14725);
and UO_488 (O_488,N_14810,N_14873);
nor UO_489 (O_489,N_14999,N_14690);
nand UO_490 (O_490,N_14838,N_14807);
nor UO_491 (O_491,N_14776,N_14935);
nor UO_492 (O_492,N_14588,N_14928);
and UO_493 (O_493,N_14731,N_14901);
or UO_494 (O_494,N_14944,N_14827);
nor UO_495 (O_495,N_14700,N_14835);
xnor UO_496 (O_496,N_14736,N_14831);
nor UO_497 (O_497,N_14732,N_14556);
nand UO_498 (O_498,N_14967,N_14626);
nor UO_499 (O_499,N_14518,N_14614);
or UO_500 (O_500,N_14564,N_14504);
nor UO_501 (O_501,N_14618,N_14941);
nand UO_502 (O_502,N_14686,N_14561);
and UO_503 (O_503,N_14857,N_14813);
nand UO_504 (O_504,N_14950,N_14892);
nand UO_505 (O_505,N_14761,N_14620);
and UO_506 (O_506,N_14884,N_14903);
nand UO_507 (O_507,N_14839,N_14641);
xnor UO_508 (O_508,N_14637,N_14545);
xor UO_509 (O_509,N_14997,N_14981);
or UO_510 (O_510,N_14632,N_14723);
or UO_511 (O_511,N_14721,N_14928);
nand UO_512 (O_512,N_14907,N_14951);
xnor UO_513 (O_513,N_14906,N_14709);
xnor UO_514 (O_514,N_14730,N_14745);
or UO_515 (O_515,N_14989,N_14790);
nor UO_516 (O_516,N_14597,N_14633);
nor UO_517 (O_517,N_14908,N_14570);
nand UO_518 (O_518,N_14564,N_14602);
nand UO_519 (O_519,N_14833,N_14963);
xor UO_520 (O_520,N_14777,N_14986);
or UO_521 (O_521,N_14519,N_14550);
nor UO_522 (O_522,N_14857,N_14788);
nand UO_523 (O_523,N_14603,N_14664);
and UO_524 (O_524,N_14879,N_14669);
nor UO_525 (O_525,N_14978,N_14608);
nand UO_526 (O_526,N_14924,N_14995);
nand UO_527 (O_527,N_14649,N_14672);
and UO_528 (O_528,N_14930,N_14849);
xor UO_529 (O_529,N_14634,N_14914);
and UO_530 (O_530,N_14580,N_14661);
nand UO_531 (O_531,N_14803,N_14532);
and UO_532 (O_532,N_14702,N_14947);
xnor UO_533 (O_533,N_14782,N_14629);
xor UO_534 (O_534,N_14802,N_14593);
and UO_535 (O_535,N_14759,N_14585);
xnor UO_536 (O_536,N_14839,N_14925);
nor UO_537 (O_537,N_14528,N_14996);
xor UO_538 (O_538,N_14528,N_14998);
xnor UO_539 (O_539,N_14562,N_14916);
nand UO_540 (O_540,N_14539,N_14662);
and UO_541 (O_541,N_14528,N_14818);
xor UO_542 (O_542,N_14803,N_14979);
xnor UO_543 (O_543,N_14970,N_14871);
xor UO_544 (O_544,N_14606,N_14717);
xor UO_545 (O_545,N_14876,N_14831);
xnor UO_546 (O_546,N_14610,N_14937);
nor UO_547 (O_547,N_14832,N_14708);
and UO_548 (O_548,N_14684,N_14875);
or UO_549 (O_549,N_14550,N_14988);
nand UO_550 (O_550,N_14696,N_14665);
or UO_551 (O_551,N_14534,N_14904);
or UO_552 (O_552,N_14759,N_14565);
and UO_553 (O_553,N_14744,N_14759);
and UO_554 (O_554,N_14799,N_14818);
and UO_555 (O_555,N_14539,N_14684);
and UO_556 (O_556,N_14623,N_14945);
and UO_557 (O_557,N_14679,N_14891);
nor UO_558 (O_558,N_14760,N_14970);
and UO_559 (O_559,N_14806,N_14964);
xor UO_560 (O_560,N_14800,N_14744);
nor UO_561 (O_561,N_14723,N_14743);
nor UO_562 (O_562,N_14544,N_14987);
nand UO_563 (O_563,N_14961,N_14626);
or UO_564 (O_564,N_14597,N_14943);
nand UO_565 (O_565,N_14605,N_14741);
nand UO_566 (O_566,N_14676,N_14894);
and UO_567 (O_567,N_14706,N_14988);
or UO_568 (O_568,N_14625,N_14746);
xnor UO_569 (O_569,N_14534,N_14885);
or UO_570 (O_570,N_14611,N_14933);
nand UO_571 (O_571,N_14804,N_14648);
nand UO_572 (O_572,N_14740,N_14905);
or UO_573 (O_573,N_14818,N_14904);
nand UO_574 (O_574,N_14661,N_14744);
xnor UO_575 (O_575,N_14831,N_14928);
xnor UO_576 (O_576,N_14632,N_14836);
xnor UO_577 (O_577,N_14699,N_14835);
and UO_578 (O_578,N_14918,N_14841);
and UO_579 (O_579,N_14503,N_14736);
xnor UO_580 (O_580,N_14951,N_14999);
xor UO_581 (O_581,N_14685,N_14631);
or UO_582 (O_582,N_14980,N_14624);
xor UO_583 (O_583,N_14979,N_14986);
or UO_584 (O_584,N_14775,N_14629);
nor UO_585 (O_585,N_14733,N_14606);
nor UO_586 (O_586,N_14557,N_14570);
and UO_587 (O_587,N_14739,N_14507);
and UO_588 (O_588,N_14548,N_14515);
xor UO_589 (O_589,N_14760,N_14511);
and UO_590 (O_590,N_14631,N_14666);
nor UO_591 (O_591,N_14925,N_14835);
or UO_592 (O_592,N_14816,N_14856);
or UO_593 (O_593,N_14667,N_14723);
xnor UO_594 (O_594,N_14725,N_14864);
or UO_595 (O_595,N_14598,N_14575);
xnor UO_596 (O_596,N_14667,N_14999);
and UO_597 (O_597,N_14892,N_14534);
nand UO_598 (O_598,N_14799,N_14685);
nor UO_599 (O_599,N_14951,N_14819);
and UO_600 (O_600,N_14708,N_14870);
xor UO_601 (O_601,N_14965,N_14980);
nor UO_602 (O_602,N_14593,N_14638);
nand UO_603 (O_603,N_14622,N_14847);
nand UO_604 (O_604,N_14736,N_14818);
nor UO_605 (O_605,N_14794,N_14863);
nand UO_606 (O_606,N_14637,N_14969);
xnor UO_607 (O_607,N_14862,N_14960);
nor UO_608 (O_608,N_14642,N_14676);
nand UO_609 (O_609,N_14766,N_14656);
nor UO_610 (O_610,N_14914,N_14866);
and UO_611 (O_611,N_14657,N_14935);
or UO_612 (O_612,N_14689,N_14853);
xor UO_613 (O_613,N_14576,N_14693);
nor UO_614 (O_614,N_14939,N_14882);
or UO_615 (O_615,N_14862,N_14827);
nand UO_616 (O_616,N_14657,N_14509);
nand UO_617 (O_617,N_14845,N_14888);
xor UO_618 (O_618,N_14722,N_14758);
nor UO_619 (O_619,N_14612,N_14510);
nor UO_620 (O_620,N_14543,N_14816);
or UO_621 (O_621,N_14764,N_14781);
and UO_622 (O_622,N_14850,N_14863);
nand UO_623 (O_623,N_14961,N_14589);
nand UO_624 (O_624,N_14533,N_14962);
xor UO_625 (O_625,N_14798,N_14965);
and UO_626 (O_626,N_14511,N_14503);
and UO_627 (O_627,N_14689,N_14979);
nand UO_628 (O_628,N_14672,N_14765);
and UO_629 (O_629,N_14747,N_14761);
nand UO_630 (O_630,N_14825,N_14848);
or UO_631 (O_631,N_14708,N_14550);
nand UO_632 (O_632,N_14534,N_14783);
or UO_633 (O_633,N_14816,N_14711);
and UO_634 (O_634,N_14902,N_14507);
and UO_635 (O_635,N_14900,N_14842);
and UO_636 (O_636,N_14682,N_14709);
and UO_637 (O_637,N_14842,N_14576);
and UO_638 (O_638,N_14871,N_14692);
and UO_639 (O_639,N_14923,N_14650);
and UO_640 (O_640,N_14520,N_14551);
xor UO_641 (O_641,N_14999,N_14856);
nor UO_642 (O_642,N_14793,N_14931);
nor UO_643 (O_643,N_14908,N_14675);
or UO_644 (O_644,N_14933,N_14618);
nor UO_645 (O_645,N_14880,N_14635);
nand UO_646 (O_646,N_14535,N_14544);
nor UO_647 (O_647,N_14595,N_14647);
nor UO_648 (O_648,N_14947,N_14768);
xor UO_649 (O_649,N_14980,N_14940);
nor UO_650 (O_650,N_14902,N_14870);
xor UO_651 (O_651,N_14835,N_14512);
nor UO_652 (O_652,N_14778,N_14541);
or UO_653 (O_653,N_14989,N_14719);
nand UO_654 (O_654,N_14773,N_14554);
xnor UO_655 (O_655,N_14871,N_14612);
nor UO_656 (O_656,N_14500,N_14905);
xnor UO_657 (O_657,N_14998,N_14976);
nand UO_658 (O_658,N_14955,N_14587);
xor UO_659 (O_659,N_14861,N_14673);
xnor UO_660 (O_660,N_14742,N_14851);
nor UO_661 (O_661,N_14964,N_14828);
xnor UO_662 (O_662,N_14522,N_14673);
or UO_663 (O_663,N_14530,N_14836);
or UO_664 (O_664,N_14539,N_14792);
or UO_665 (O_665,N_14693,N_14924);
xor UO_666 (O_666,N_14778,N_14547);
xnor UO_667 (O_667,N_14766,N_14967);
nand UO_668 (O_668,N_14700,N_14574);
nor UO_669 (O_669,N_14644,N_14939);
nor UO_670 (O_670,N_14870,N_14743);
or UO_671 (O_671,N_14907,N_14912);
and UO_672 (O_672,N_14663,N_14870);
or UO_673 (O_673,N_14710,N_14587);
xor UO_674 (O_674,N_14948,N_14523);
and UO_675 (O_675,N_14864,N_14944);
and UO_676 (O_676,N_14831,N_14798);
or UO_677 (O_677,N_14549,N_14918);
or UO_678 (O_678,N_14937,N_14782);
xnor UO_679 (O_679,N_14936,N_14891);
nand UO_680 (O_680,N_14599,N_14905);
nor UO_681 (O_681,N_14542,N_14924);
nand UO_682 (O_682,N_14897,N_14860);
nand UO_683 (O_683,N_14849,N_14538);
xor UO_684 (O_684,N_14977,N_14553);
xor UO_685 (O_685,N_14927,N_14854);
or UO_686 (O_686,N_14593,N_14835);
nand UO_687 (O_687,N_14759,N_14838);
or UO_688 (O_688,N_14975,N_14558);
xor UO_689 (O_689,N_14980,N_14553);
nand UO_690 (O_690,N_14570,N_14521);
xor UO_691 (O_691,N_14792,N_14677);
nor UO_692 (O_692,N_14636,N_14607);
nand UO_693 (O_693,N_14882,N_14935);
nor UO_694 (O_694,N_14950,N_14657);
nor UO_695 (O_695,N_14569,N_14921);
nand UO_696 (O_696,N_14819,N_14761);
and UO_697 (O_697,N_14793,N_14914);
nand UO_698 (O_698,N_14786,N_14901);
nand UO_699 (O_699,N_14792,N_14864);
and UO_700 (O_700,N_14565,N_14657);
or UO_701 (O_701,N_14625,N_14878);
nand UO_702 (O_702,N_14716,N_14504);
nand UO_703 (O_703,N_14672,N_14589);
xnor UO_704 (O_704,N_14840,N_14897);
nor UO_705 (O_705,N_14537,N_14557);
nand UO_706 (O_706,N_14961,N_14665);
nand UO_707 (O_707,N_14552,N_14681);
nor UO_708 (O_708,N_14852,N_14882);
nor UO_709 (O_709,N_14993,N_14546);
xor UO_710 (O_710,N_14606,N_14726);
xor UO_711 (O_711,N_14693,N_14861);
or UO_712 (O_712,N_14811,N_14555);
and UO_713 (O_713,N_14848,N_14872);
nand UO_714 (O_714,N_14875,N_14607);
xnor UO_715 (O_715,N_14810,N_14576);
and UO_716 (O_716,N_14563,N_14862);
xor UO_717 (O_717,N_14989,N_14840);
and UO_718 (O_718,N_14954,N_14859);
or UO_719 (O_719,N_14861,N_14795);
nand UO_720 (O_720,N_14957,N_14995);
nor UO_721 (O_721,N_14711,N_14930);
nand UO_722 (O_722,N_14532,N_14811);
and UO_723 (O_723,N_14653,N_14670);
and UO_724 (O_724,N_14645,N_14796);
nand UO_725 (O_725,N_14808,N_14745);
nor UO_726 (O_726,N_14695,N_14956);
xnor UO_727 (O_727,N_14705,N_14810);
nor UO_728 (O_728,N_14865,N_14962);
nor UO_729 (O_729,N_14510,N_14566);
and UO_730 (O_730,N_14660,N_14959);
xor UO_731 (O_731,N_14838,N_14674);
xor UO_732 (O_732,N_14751,N_14727);
or UO_733 (O_733,N_14964,N_14593);
xor UO_734 (O_734,N_14650,N_14537);
and UO_735 (O_735,N_14914,N_14844);
nand UO_736 (O_736,N_14798,N_14914);
xor UO_737 (O_737,N_14788,N_14629);
nand UO_738 (O_738,N_14802,N_14811);
nand UO_739 (O_739,N_14777,N_14646);
or UO_740 (O_740,N_14795,N_14528);
or UO_741 (O_741,N_14695,N_14599);
nand UO_742 (O_742,N_14825,N_14603);
and UO_743 (O_743,N_14900,N_14923);
or UO_744 (O_744,N_14577,N_14987);
nor UO_745 (O_745,N_14708,N_14578);
and UO_746 (O_746,N_14529,N_14785);
and UO_747 (O_747,N_14582,N_14898);
nand UO_748 (O_748,N_14860,N_14811);
nand UO_749 (O_749,N_14791,N_14760);
or UO_750 (O_750,N_14540,N_14561);
or UO_751 (O_751,N_14939,N_14815);
nand UO_752 (O_752,N_14792,N_14727);
nand UO_753 (O_753,N_14882,N_14623);
nand UO_754 (O_754,N_14577,N_14864);
xnor UO_755 (O_755,N_14899,N_14507);
and UO_756 (O_756,N_14814,N_14609);
xnor UO_757 (O_757,N_14682,N_14852);
nand UO_758 (O_758,N_14808,N_14838);
xor UO_759 (O_759,N_14661,N_14662);
nand UO_760 (O_760,N_14957,N_14574);
nand UO_761 (O_761,N_14643,N_14561);
and UO_762 (O_762,N_14659,N_14997);
nand UO_763 (O_763,N_14825,N_14965);
xnor UO_764 (O_764,N_14551,N_14900);
nand UO_765 (O_765,N_14892,N_14755);
or UO_766 (O_766,N_14888,N_14862);
nor UO_767 (O_767,N_14686,N_14503);
or UO_768 (O_768,N_14718,N_14850);
xor UO_769 (O_769,N_14932,N_14549);
or UO_770 (O_770,N_14817,N_14548);
nand UO_771 (O_771,N_14798,N_14931);
nor UO_772 (O_772,N_14848,N_14643);
nor UO_773 (O_773,N_14768,N_14567);
or UO_774 (O_774,N_14640,N_14858);
and UO_775 (O_775,N_14907,N_14835);
and UO_776 (O_776,N_14590,N_14694);
and UO_777 (O_777,N_14716,N_14930);
xor UO_778 (O_778,N_14677,N_14979);
or UO_779 (O_779,N_14918,N_14619);
nand UO_780 (O_780,N_14575,N_14884);
and UO_781 (O_781,N_14608,N_14901);
or UO_782 (O_782,N_14817,N_14899);
and UO_783 (O_783,N_14579,N_14703);
and UO_784 (O_784,N_14966,N_14620);
xnor UO_785 (O_785,N_14651,N_14666);
nor UO_786 (O_786,N_14727,N_14771);
nor UO_787 (O_787,N_14796,N_14699);
nand UO_788 (O_788,N_14829,N_14569);
and UO_789 (O_789,N_14880,N_14953);
and UO_790 (O_790,N_14899,N_14651);
nand UO_791 (O_791,N_14700,N_14970);
xnor UO_792 (O_792,N_14817,N_14783);
nor UO_793 (O_793,N_14630,N_14853);
nor UO_794 (O_794,N_14589,N_14629);
nand UO_795 (O_795,N_14694,N_14625);
and UO_796 (O_796,N_14847,N_14983);
nor UO_797 (O_797,N_14839,N_14892);
nand UO_798 (O_798,N_14736,N_14846);
and UO_799 (O_799,N_14553,N_14874);
or UO_800 (O_800,N_14885,N_14813);
xnor UO_801 (O_801,N_14794,N_14805);
xor UO_802 (O_802,N_14982,N_14516);
or UO_803 (O_803,N_14592,N_14790);
or UO_804 (O_804,N_14584,N_14705);
xor UO_805 (O_805,N_14649,N_14820);
xor UO_806 (O_806,N_14806,N_14807);
xnor UO_807 (O_807,N_14500,N_14976);
xnor UO_808 (O_808,N_14909,N_14613);
xnor UO_809 (O_809,N_14964,N_14632);
and UO_810 (O_810,N_14733,N_14849);
or UO_811 (O_811,N_14908,N_14714);
nor UO_812 (O_812,N_14605,N_14710);
nand UO_813 (O_813,N_14636,N_14699);
and UO_814 (O_814,N_14908,N_14865);
nor UO_815 (O_815,N_14700,N_14587);
nand UO_816 (O_816,N_14795,N_14790);
nor UO_817 (O_817,N_14664,N_14835);
and UO_818 (O_818,N_14562,N_14527);
xnor UO_819 (O_819,N_14503,N_14864);
and UO_820 (O_820,N_14975,N_14695);
nand UO_821 (O_821,N_14833,N_14934);
nor UO_822 (O_822,N_14652,N_14791);
xor UO_823 (O_823,N_14785,N_14962);
xor UO_824 (O_824,N_14613,N_14666);
nand UO_825 (O_825,N_14690,N_14648);
nor UO_826 (O_826,N_14713,N_14997);
and UO_827 (O_827,N_14740,N_14761);
xor UO_828 (O_828,N_14718,N_14909);
or UO_829 (O_829,N_14802,N_14665);
xor UO_830 (O_830,N_14817,N_14871);
nand UO_831 (O_831,N_14500,N_14659);
and UO_832 (O_832,N_14566,N_14703);
and UO_833 (O_833,N_14583,N_14565);
nor UO_834 (O_834,N_14873,N_14623);
or UO_835 (O_835,N_14864,N_14554);
nor UO_836 (O_836,N_14623,N_14839);
nor UO_837 (O_837,N_14509,N_14526);
nor UO_838 (O_838,N_14961,N_14811);
or UO_839 (O_839,N_14788,N_14868);
or UO_840 (O_840,N_14772,N_14587);
nor UO_841 (O_841,N_14857,N_14557);
or UO_842 (O_842,N_14580,N_14599);
nand UO_843 (O_843,N_14943,N_14885);
or UO_844 (O_844,N_14562,N_14624);
nand UO_845 (O_845,N_14686,N_14784);
and UO_846 (O_846,N_14919,N_14860);
xor UO_847 (O_847,N_14774,N_14929);
or UO_848 (O_848,N_14881,N_14753);
xor UO_849 (O_849,N_14847,N_14558);
nor UO_850 (O_850,N_14718,N_14530);
or UO_851 (O_851,N_14519,N_14540);
and UO_852 (O_852,N_14618,N_14515);
or UO_853 (O_853,N_14668,N_14806);
nor UO_854 (O_854,N_14597,N_14664);
nor UO_855 (O_855,N_14716,N_14665);
nor UO_856 (O_856,N_14540,N_14924);
nor UO_857 (O_857,N_14791,N_14787);
xor UO_858 (O_858,N_14774,N_14524);
nand UO_859 (O_859,N_14919,N_14569);
xnor UO_860 (O_860,N_14955,N_14827);
xor UO_861 (O_861,N_14952,N_14672);
nand UO_862 (O_862,N_14668,N_14938);
xor UO_863 (O_863,N_14667,N_14599);
nand UO_864 (O_864,N_14640,N_14695);
nand UO_865 (O_865,N_14958,N_14632);
or UO_866 (O_866,N_14522,N_14526);
and UO_867 (O_867,N_14773,N_14678);
and UO_868 (O_868,N_14996,N_14752);
nand UO_869 (O_869,N_14531,N_14857);
or UO_870 (O_870,N_14564,N_14733);
and UO_871 (O_871,N_14746,N_14741);
xnor UO_872 (O_872,N_14570,N_14864);
xnor UO_873 (O_873,N_14983,N_14839);
and UO_874 (O_874,N_14708,N_14952);
and UO_875 (O_875,N_14620,N_14500);
and UO_876 (O_876,N_14927,N_14910);
xor UO_877 (O_877,N_14894,N_14830);
or UO_878 (O_878,N_14516,N_14504);
and UO_879 (O_879,N_14873,N_14640);
nor UO_880 (O_880,N_14629,N_14686);
or UO_881 (O_881,N_14736,N_14782);
nand UO_882 (O_882,N_14600,N_14522);
nand UO_883 (O_883,N_14585,N_14648);
nor UO_884 (O_884,N_14656,N_14931);
nor UO_885 (O_885,N_14774,N_14888);
xor UO_886 (O_886,N_14674,N_14807);
xnor UO_887 (O_887,N_14805,N_14656);
and UO_888 (O_888,N_14674,N_14580);
nand UO_889 (O_889,N_14627,N_14718);
xnor UO_890 (O_890,N_14553,N_14962);
or UO_891 (O_891,N_14740,N_14805);
or UO_892 (O_892,N_14796,N_14819);
nand UO_893 (O_893,N_14776,N_14795);
nand UO_894 (O_894,N_14790,N_14926);
xor UO_895 (O_895,N_14780,N_14792);
and UO_896 (O_896,N_14837,N_14787);
nor UO_897 (O_897,N_14930,N_14914);
and UO_898 (O_898,N_14971,N_14783);
xor UO_899 (O_899,N_14894,N_14834);
and UO_900 (O_900,N_14939,N_14586);
nand UO_901 (O_901,N_14718,N_14949);
xor UO_902 (O_902,N_14633,N_14805);
xnor UO_903 (O_903,N_14663,N_14749);
nand UO_904 (O_904,N_14589,N_14987);
xnor UO_905 (O_905,N_14778,N_14642);
or UO_906 (O_906,N_14690,N_14923);
nand UO_907 (O_907,N_14998,N_14980);
or UO_908 (O_908,N_14669,N_14960);
or UO_909 (O_909,N_14548,N_14525);
nor UO_910 (O_910,N_14820,N_14609);
xor UO_911 (O_911,N_14804,N_14965);
xor UO_912 (O_912,N_14816,N_14599);
nand UO_913 (O_913,N_14781,N_14669);
nand UO_914 (O_914,N_14939,N_14685);
xor UO_915 (O_915,N_14987,N_14540);
nor UO_916 (O_916,N_14768,N_14599);
nor UO_917 (O_917,N_14939,N_14543);
or UO_918 (O_918,N_14594,N_14837);
nand UO_919 (O_919,N_14978,N_14877);
or UO_920 (O_920,N_14890,N_14556);
and UO_921 (O_921,N_14829,N_14998);
nor UO_922 (O_922,N_14639,N_14804);
nand UO_923 (O_923,N_14529,N_14810);
xnor UO_924 (O_924,N_14888,N_14975);
nand UO_925 (O_925,N_14691,N_14858);
xnor UO_926 (O_926,N_14532,N_14647);
xnor UO_927 (O_927,N_14681,N_14634);
xor UO_928 (O_928,N_14654,N_14733);
and UO_929 (O_929,N_14811,N_14569);
or UO_930 (O_930,N_14909,N_14665);
or UO_931 (O_931,N_14538,N_14553);
xnor UO_932 (O_932,N_14817,N_14847);
nand UO_933 (O_933,N_14920,N_14820);
nor UO_934 (O_934,N_14916,N_14837);
nor UO_935 (O_935,N_14875,N_14666);
nand UO_936 (O_936,N_14532,N_14837);
xor UO_937 (O_937,N_14898,N_14773);
or UO_938 (O_938,N_14872,N_14922);
and UO_939 (O_939,N_14525,N_14505);
and UO_940 (O_940,N_14721,N_14510);
nor UO_941 (O_941,N_14620,N_14664);
nand UO_942 (O_942,N_14873,N_14861);
or UO_943 (O_943,N_14698,N_14910);
nand UO_944 (O_944,N_14726,N_14630);
xor UO_945 (O_945,N_14678,N_14801);
nand UO_946 (O_946,N_14816,N_14815);
or UO_947 (O_947,N_14833,N_14589);
nor UO_948 (O_948,N_14651,N_14610);
xnor UO_949 (O_949,N_14990,N_14543);
nor UO_950 (O_950,N_14812,N_14794);
nor UO_951 (O_951,N_14680,N_14965);
nor UO_952 (O_952,N_14524,N_14796);
or UO_953 (O_953,N_14507,N_14862);
xnor UO_954 (O_954,N_14808,N_14754);
and UO_955 (O_955,N_14715,N_14505);
nand UO_956 (O_956,N_14772,N_14934);
nand UO_957 (O_957,N_14697,N_14780);
and UO_958 (O_958,N_14879,N_14984);
or UO_959 (O_959,N_14783,N_14777);
nand UO_960 (O_960,N_14658,N_14948);
and UO_961 (O_961,N_14687,N_14904);
and UO_962 (O_962,N_14740,N_14868);
nor UO_963 (O_963,N_14629,N_14912);
xor UO_964 (O_964,N_14746,N_14875);
or UO_965 (O_965,N_14529,N_14943);
and UO_966 (O_966,N_14893,N_14991);
nor UO_967 (O_967,N_14601,N_14538);
nor UO_968 (O_968,N_14794,N_14533);
nor UO_969 (O_969,N_14544,N_14594);
or UO_970 (O_970,N_14888,N_14634);
xnor UO_971 (O_971,N_14842,N_14504);
nor UO_972 (O_972,N_14910,N_14771);
nor UO_973 (O_973,N_14776,N_14669);
xor UO_974 (O_974,N_14602,N_14510);
and UO_975 (O_975,N_14730,N_14940);
nor UO_976 (O_976,N_14695,N_14540);
and UO_977 (O_977,N_14539,N_14919);
or UO_978 (O_978,N_14773,N_14956);
nand UO_979 (O_979,N_14697,N_14920);
and UO_980 (O_980,N_14700,N_14956);
or UO_981 (O_981,N_14771,N_14698);
xor UO_982 (O_982,N_14870,N_14634);
nand UO_983 (O_983,N_14505,N_14565);
or UO_984 (O_984,N_14891,N_14846);
and UO_985 (O_985,N_14517,N_14547);
nor UO_986 (O_986,N_14928,N_14551);
nor UO_987 (O_987,N_14683,N_14840);
nor UO_988 (O_988,N_14674,N_14522);
xor UO_989 (O_989,N_14836,N_14816);
nor UO_990 (O_990,N_14702,N_14964);
and UO_991 (O_991,N_14705,N_14646);
and UO_992 (O_992,N_14578,N_14844);
nor UO_993 (O_993,N_14905,N_14814);
nand UO_994 (O_994,N_14749,N_14858);
and UO_995 (O_995,N_14899,N_14505);
xnor UO_996 (O_996,N_14553,N_14672);
nand UO_997 (O_997,N_14566,N_14931);
and UO_998 (O_998,N_14864,N_14538);
nand UO_999 (O_999,N_14518,N_14986);
nand UO_1000 (O_1000,N_14682,N_14560);
nand UO_1001 (O_1001,N_14788,N_14818);
or UO_1002 (O_1002,N_14973,N_14616);
nor UO_1003 (O_1003,N_14796,N_14508);
and UO_1004 (O_1004,N_14691,N_14632);
and UO_1005 (O_1005,N_14917,N_14701);
and UO_1006 (O_1006,N_14678,N_14888);
and UO_1007 (O_1007,N_14537,N_14850);
nor UO_1008 (O_1008,N_14899,N_14536);
xor UO_1009 (O_1009,N_14822,N_14917);
nor UO_1010 (O_1010,N_14581,N_14851);
nor UO_1011 (O_1011,N_14527,N_14637);
nand UO_1012 (O_1012,N_14816,N_14637);
xnor UO_1013 (O_1013,N_14883,N_14726);
and UO_1014 (O_1014,N_14969,N_14787);
nand UO_1015 (O_1015,N_14862,N_14913);
nor UO_1016 (O_1016,N_14585,N_14951);
xnor UO_1017 (O_1017,N_14752,N_14670);
xnor UO_1018 (O_1018,N_14875,N_14588);
or UO_1019 (O_1019,N_14660,N_14903);
xnor UO_1020 (O_1020,N_14522,N_14976);
xor UO_1021 (O_1021,N_14684,N_14740);
or UO_1022 (O_1022,N_14691,N_14630);
xor UO_1023 (O_1023,N_14853,N_14937);
and UO_1024 (O_1024,N_14922,N_14811);
or UO_1025 (O_1025,N_14892,N_14979);
nand UO_1026 (O_1026,N_14992,N_14521);
or UO_1027 (O_1027,N_14973,N_14579);
xor UO_1028 (O_1028,N_14539,N_14747);
and UO_1029 (O_1029,N_14825,N_14538);
nand UO_1030 (O_1030,N_14841,N_14826);
and UO_1031 (O_1031,N_14911,N_14649);
nand UO_1032 (O_1032,N_14514,N_14510);
and UO_1033 (O_1033,N_14587,N_14702);
and UO_1034 (O_1034,N_14930,N_14848);
xnor UO_1035 (O_1035,N_14680,N_14808);
and UO_1036 (O_1036,N_14808,N_14660);
xnor UO_1037 (O_1037,N_14529,N_14989);
and UO_1038 (O_1038,N_14682,N_14618);
or UO_1039 (O_1039,N_14568,N_14895);
nor UO_1040 (O_1040,N_14634,N_14640);
nand UO_1041 (O_1041,N_14965,N_14901);
or UO_1042 (O_1042,N_14932,N_14692);
or UO_1043 (O_1043,N_14993,N_14592);
nand UO_1044 (O_1044,N_14994,N_14773);
nor UO_1045 (O_1045,N_14503,N_14907);
or UO_1046 (O_1046,N_14583,N_14588);
nor UO_1047 (O_1047,N_14765,N_14570);
nand UO_1048 (O_1048,N_14548,N_14505);
and UO_1049 (O_1049,N_14913,N_14852);
and UO_1050 (O_1050,N_14790,N_14623);
or UO_1051 (O_1051,N_14691,N_14716);
or UO_1052 (O_1052,N_14525,N_14835);
xnor UO_1053 (O_1053,N_14869,N_14840);
nand UO_1054 (O_1054,N_14619,N_14812);
or UO_1055 (O_1055,N_14696,N_14636);
and UO_1056 (O_1056,N_14680,N_14971);
xor UO_1057 (O_1057,N_14858,N_14527);
xnor UO_1058 (O_1058,N_14559,N_14549);
nand UO_1059 (O_1059,N_14516,N_14996);
nor UO_1060 (O_1060,N_14759,N_14763);
xnor UO_1061 (O_1061,N_14988,N_14914);
and UO_1062 (O_1062,N_14940,N_14853);
nand UO_1063 (O_1063,N_14642,N_14521);
or UO_1064 (O_1064,N_14713,N_14968);
or UO_1065 (O_1065,N_14591,N_14619);
nor UO_1066 (O_1066,N_14927,N_14706);
xor UO_1067 (O_1067,N_14890,N_14779);
and UO_1068 (O_1068,N_14593,N_14968);
and UO_1069 (O_1069,N_14539,N_14795);
or UO_1070 (O_1070,N_14988,N_14796);
or UO_1071 (O_1071,N_14545,N_14880);
and UO_1072 (O_1072,N_14749,N_14802);
nand UO_1073 (O_1073,N_14763,N_14876);
xor UO_1074 (O_1074,N_14895,N_14528);
xor UO_1075 (O_1075,N_14725,N_14728);
or UO_1076 (O_1076,N_14574,N_14557);
nand UO_1077 (O_1077,N_14922,N_14786);
nor UO_1078 (O_1078,N_14830,N_14922);
and UO_1079 (O_1079,N_14931,N_14813);
or UO_1080 (O_1080,N_14629,N_14666);
and UO_1081 (O_1081,N_14819,N_14750);
nor UO_1082 (O_1082,N_14652,N_14932);
and UO_1083 (O_1083,N_14944,N_14808);
or UO_1084 (O_1084,N_14703,N_14945);
or UO_1085 (O_1085,N_14548,N_14845);
or UO_1086 (O_1086,N_14959,N_14849);
nor UO_1087 (O_1087,N_14820,N_14905);
nor UO_1088 (O_1088,N_14581,N_14710);
nand UO_1089 (O_1089,N_14543,N_14737);
and UO_1090 (O_1090,N_14990,N_14926);
and UO_1091 (O_1091,N_14611,N_14733);
nor UO_1092 (O_1092,N_14626,N_14819);
xnor UO_1093 (O_1093,N_14676,N_14502);
xnor UO_1094 (O_1094,N_14596,N_14950);
nor UO_1095 (O_1095,N_14536,N_14741);
xnor UO_1096 (O_1096,N_14793,N_14780);
nor UO_1097 (O_1097,N_14961,N_14728);
nand UO_1098 (O_1098,N_14873,N_14979);
nor UO_1099 (O_1099,N_14521,N_14697);
nand UO_1100 (O_1100,N_14715,N_14558);
xnor UO_1101 (O_1101,N_14956,N_14874);
nand UO_1102 (O_1102,N_14569,N_14978);
and UO_1103 (O_1103,N_14798,N_14547);
or UO_1104 (O_1104,N_14817,N_14518);
xor UO_1105 (O_1105,N_14947,N_14880);
or UO_1106 (O_1106,N_14963,N_14832);
or UO_1107 (O_1107,N_14795,N_14970);
nor UO_1108 (O_1108,N_14508,N_14683);
and UO_1109 (O_1109,N_14585,N_14717);
nand UO_1110 (O_1110,N_14582,N_14968);
or UO_1111 (O_1111,N_14540,N_14527);
and UO_1112 (O_1112,N_14951,N_14671);
nor UO_1113 (O_1113,N_14799,N_14948);
and UO_1114 (O_1114,N_14854,N_14973);
xnor UO_1115 (O_1115,N_14772,N_14524);
nor UO_1116 (O_1116,N_14921,N_14503);
xnor UO_1117 (O_1117,N_14576,N_14822);
nor UO_1118 (O_1118,N_14910,N_14613);
nor UO_1119 (O_1119,N_14783,N_14813);
nor UO_1120 (O_1120,N_14824,N_14621);
or UO_1121 (O_1121,N_14724,N_14778);
and UO_1122 (O_1122,N_14891,N_14732);
xnor UO_1123 (O_1123,N_14950,N_14994);
or UO_1124 (O_1124,N_14744,N_14980);
xor UO_1125 (O_1125,N_14689,N_14603);
xor UO_1126 (O_1126,N_14996,N_14514);
or UO_1127 (O_1127,N_14632,N_14899);
xor UO_1128 (O_1128,N_14747,N_14858);
or UO_1129 (O_1129,N_14732,N_14788);
nand UO_1130 (O_1130,N_14820,N_14683);
or UO_1131 (O_1131,N_14553,N_14792);
and UO_1132 (O_1132,N_14970,N_14944);
nand UO_1133 (O_1133,N_14809,N_14881);
xnor UO_1134 (O_1134,N_14622,N_14798);
xor UO_1135 (O_1135,N_14967,N_14712);
nand UO_1136 (O_1136,N_14648,N_14764);
xor UO_1137 (O_1137,N_14609,N_14989);
nand UO_1138 (O_1138,N_14703,N_14590);
or UO_1139 (O_1139,N_14568,N_14831);
xor UO_1140 (O_1140,N_14620,N_14796);
and UO_1141 (O_1141,N_14884,N_14529);
nand UO_1142 (O_1142,N_14889,N_14780);
or UO_1143 (O_1143,N_14734,N_14637);
nand UO_1144 (O_1144,N_14640,N_14649);
nand UO_1145 (O_1145,N_14687,N_14934);
and UO_1146 (O_1146,N_14877,N_14958);
or UO_1147 (O_1147,N_14952,N_14922);
and UO_1148 (O_1148,N_14685,N_14773);
and UO_1149 (O_1149,N_14997,N_14597);
xnor UO_1150 (O_1150,N_14625,N_14779);
or UO_1151 (O_1151,N_14549,N_14688);
or UO_1152 (O_1152,N_14504,N_14543);
nand UO_1153 (O_1153,N_14948,N_14638);
xor UO_1154 (O_1154,N_14658,N_14866);
nand UO_1155 (O_1155,N_14520,N_14572);
and UO_1156 (O_1156,N_14586,N_14820);
nor UO_1157 (O_1157,N_14971,N_14526);
xor UO_1158 (O_1158,N_14978,N_14913);
and UO_1159 (O_1159,N_14952,N_14833);
nor UO_1160 (O_1160,N_14889,N_14699);
nor UO_1161 (O_1161,N_14732,N_14956);
or UO_1162 (O_1162,N_14586,N_14984);
nand UO_1163 (O_1163,N_14742,N_14559);
or UO_1164 (O_1164,N_14737,N_14563);
or UO_1165 (O_1165,N_14892,N_14782);
xor UO_1166 (O_1166,N_14534,N_14808);
and UO_1167 (O_1167,N_14869,N_14626);
or UO_1168 (O_1168,N_14634,N_14782);
and UO_1169 (O_1169,N_14672,N_14739);
nor UO_1170 (O_1170,N_14915,N_14807);
or UO_1171 (O_1171,N_14592,N_14501);
nand UO_1172 (O_1172,N_14823,N_14995);
and UO_1173 (O_1173,N_14611,N_14745);
xnor UO_1174 (O_1174,N_14522,N_14745);
or UO_1175 (O_1175,N_14752,N_14723);
or UO_1176 (O_1176,N_14919,N_14575);
xor UO_1177 (O_1177,N_14665,N_14554);
or UO_1178 (O_1178,N_14589,N_14810);
and UO_1179 (O_1179,N_14954,N_14750);
xor UO_1180 (O_1180,N_14980,N_14941);
xnor UO_1181 (O_1181,N_14982,N_14698);
xnor UO_1182 (O_1182,N_14616,N_14981);
or UO_1183 (O_1183,N_14789,N_14538);
nor UO_1184 (O_1184,N_14823,N_14925);
xor UO_1185 (O_1185,N_14962,N_14569);
xnor UO_1186 (O_1186,N_14992,N_14965);
xor UO_1187 (O_1187,N_14693,N_14863);
nor UO_1188 (O_1188,N_14821,N_14563);
xor UO_1189 (O_1189,N_14934,N_14562);
or UO_1190 (O_1190,N_14527,N_14797);
xnor UO_1191 (O_1191,N_14589,N_14959);
and UO_1192 (O_1192,N_14527,N_14742);
nand UO_1193 (O_1193,N_14845,N_14679);
xnor UO_1194 (O_1194,N_14863,N_14807);
nand UO_1195 (O_1195,N_14872,N_14613);
or UO_1196 (O_1196,N_14694,N_14714);
xor UO_1197 (O_1197,N_14966,N_14663);
and UO_1198 (O_1198,N_14918,N_14694);
nor UO_1199 (O_1199,N_14725,N_14819);
nor UO_1200 (O_1200,N_14962,N_14867);
nor UO_1201 (O_1201,N_14549,N_14842);
or UO_1202 (O_1202,N_14597,N_14851);
and UO_1203 (O_1203,N_14708,N_14808);
and UO_1204 (O_1204,N_14781,N_14686);
xnor UO_1205 (O_1205,N_14577,N_14607);
or UO_1206 (O_1206,N_14756,N_14879);
or UO_1207 (O_1207,N_14823,N_14983);
and UO_1208 (O_1208,N_14703,N_14776);
nor UO_1209 (O_1209,N_14639,N_14611);
xnor UO_1210 (O_1210,N_14909,N_14933);
nand UO_1211 (O_1211,N_14817,N_14665);
nand UO_1212 (O_1212,N_14710,N_14726);
nand UO_1213 (O_1213,N_14797,N_14856);
or UO_1214 (O_1214,N_14990,N_14668);
or UO_1215 (O_1215,N_14686,N_14861);
nor UO_1216 (O_1216,N_14903,N_14958);
xor UO_1217 (O_1217,N_14746,N_14819);
xor UO_1218 (O_1218,N_14993,N_14566);
xnor UO_1219 (O_1219,N_14600,N_14855);
xnor UO_1220 (O_1220,N_14628,N_14939);
xor UO_1221 (O_1221,N_14955,N_14600);
nand UO_1222 (O_1222,N_14567,N_14664);
and UO_1223 (O_1223,N_14591,N_14896);
nor UO_1224 (O_1224,N_14874,N_14813);
nand UO_1225 (O_1225,N_14514,N_14686);
and UO_1226 (O_1226,N_14761,N_14611);
or UO_1227 (O_1227,N_14536,N_14511);
and UO_1228 (O_1228,N_14650,N_14903);
xor UO_1229 (O_1229,N_14817,N_14767);
xnor UO_1230 (O_1230,N_14750,N_14687);
nand UO_1231 (O_1231,N_14983,N_14506);
and UO_1232 (O_1232,N_14551,N_14638);
nand UO_1233 (O_1233,N_14944,N_14872);
xor UO_1234 (O_1234,N_14721,N_14816);
or UO_1235 (O_1235,N_14759,N_14916);
nand UO_1236 (O_1236,N_14976,N_14583);
nor UO_1237 (O_1237,N_14603,N_14754);
nand UO_1238 (O_1238,N_14593,N_14995);
nor UO_1239 (O_1239,N_14863,N_14808);
or UO_1240 (O_1240,N_14832,N_14662);
or UO_1241 (O_1241,N_14934,N_14554);
or UO_1242 (O_1242,N_14973,N_14759);
or UO_1243 (O_1243,N_14663,N_14548);
and UO_1244 (O_1244,N_14709,N_14743);
or UO_1245 (O_1245,N_14544,N_14980);
nand UO_1246 (O_1246,N_14896,N_14656);
nor UO_1247 (O_1247,N_14616,N_14727);
xor UO_1248 (O_1248,N_14965,N_14893);
xor UO_1249 (O_1249,N_14584,N_14808);
xnor UO_1250 (O_1250,N_14792,N_14523);
nor UO_1251 (O_1251,N_14724,N_14881);
nand UO_1252 (O_1252,N_14834,N_14728);
nor UO_1253 (O_1253,N_14701,N_14777);
nand UO_1254 (O_1254,N_14850,N_14922);
and UO_1255 (O_1255,N_14934,N_14526);
or UO_1256 (O_1256,N_14598,N_14835);
nor UO_1257 (O_1257,N_14749,N_14906);
nand UO_1258 (O_1258,N_14589,N_14677);
nand UO_1259 (O_1259,N_14764,N_14646);
nand UO_1260 (O_1260,N_14750,N_14880);
nor UO_1261 (O_1261,N_14793,N_14740);
or UO_1262 (O_1262,N_14877,N_14548);
xor UO_1263 (O_1263,N_14773,N_14520);
nor UO_1264 (O_1264,N_14760,N_14508);
nor UO_1265 (O_1265,N_14813,N_14902);
and UO_1266 (O_1266,N_14920,N_14721);
nand UO_1267 (O_1267,N_14987,N_14903);
nor UO_1268 (O_1268,N_14950,N_14688);
and UO_1269 (O_1269,N_14501,N_14574);
xor UO_1270 (O_1270,N_14772,N_14749);
xor UO_1271 (O_1271,N_14655,N_14955);
and UO_1272 (O_1272,N_14754,N_14903);
nor UO_1273 (O_1273,N_14694,N_14594);
or UO_1274 (O_1274,N_14974,N_14963);
nor UO_1275 (O_1275,N_14963,N_14605);
xor UO_1276 (O_1276,N_14974,N_14682);
nor UO_1277 (O_1277,N_14568,N_14734);
and UO_1278 (O_1278,N_14601,N_14864);
nand UO_1279 (O_1279,N_14758,N_14556);
or UO_1280 (O_1280,N_14657,N_14658);
xor UO_1281 (O_1281,N_14833,N_14618);
nand UO_1282 (O_1282,N_14740,N_14941);
and UO_1283 (O_1283,N_14719,N_14937);
and UO_1284 (O_1284,N_14569,N_14531);
and UO_1285 (O_1285,N_14575,N_14771);
nand UO_1286 (O_1286,N_14901,N_14668);
xor UO_1287 (O_1287,N_14758,N_14652);
nor UO_1288 (O_1288,N_14736,N_14972);
or UO_1289 (O_1289,N_14685,N_14718);
nand UO_1290 (O_1290,N_14848,N_14727);
or UO_1291 (O_1291,N_14896,N_14766);
xnor UO_1292 (O_1292,N_14783,N_14719);
xor UO_1293 (O_1293,N_14702,N_14694);
nor UO_1294 (O_1294,N_14822,N_14705);
nor UO_1295 (O_1295,N_14896,N_14847);
nand UO_1296 (O_1296,N_14668,N_14830);
nor UO_1297 (O_1297,N_14988,N_14516);
and UO_1298 (O_1298,N_14776,N_14709);
and UO_1299 (O_1299,N_14893,N_14641);
xor UO_1300 (O_1300,N_14810,N_14877);
xor UO_1301 (O_1301,N_14607,N_14758);
or UO_1302 (O_1302,N_14866,N_14672);
nor UO_1303 (O_1303,N_14583,N_14681);
xnor UO_1304 (O_1304,N_14509,N_14546);
nand UO_1305 (O_1305,N_14635,N_14744);
nor UO_1306 (O_1306,N_14846,N_14588);
nor UO_1307 (O_1307,N_14855,N_14750);
xnor UO_1308 (O_1308,N_14680,N_14888);
and UO_1309 (O_1309,N_14632,N_14927);
nor UO_1310 (O_1310,N_14923,N_14857);
nand UO_1311 (O_1311,N_14850,N_14966);
or UO_1312 (O_1312,N_14883,N_14701);
and UO_1313 (O_1313,N_14970,N_14808);
nand UO_1314 (O_1314,N_14517,N_14801);
nand UO_1315 (O_1315,N_14758,N_14887);
or UO_1316 (O_1316,N_14681,N_14963);
nand UO_1317 (O_1317,N_14953,N_14541);
nor UO_1318 (O_1318,N_14568,N_14930);
xnor UO_1319 (O_1319,N_14523,N_14649);
nor UO_1320 (O_1320,N_14557,N_14860);
nor UO_1321 (O_1321,N_14619,N_14806);
nand UO_1322 (O_1322,N_14641,N_14563);
xnor UO_1323 (O_1323,N_14630,N_14983);
or UO_1324 (O_1324,N_14530,N_14809);
nand UO_1325 (O_1325,N_14928,N_14795);
nand UO_1326 (O_1326,N_14620,N_14800);
nor UO_1327 (O_1327,N_14883,N_14751);
nand UO_1328 (O_1328,N_14868,N_14900);
nor UO_1329 (O_1329,N_14786,N_14832);
and UO_1330 (O_1330,N_14977,N_14648);
xnor UO_1331 (O_1331,N_14603,N_14545);
and UO_1332 (O_1332,N_14579,N_14802);
nand UO_1333 (O_1333,N_14886,N_14641);
nor UO_1334 (O_1334,N_14681,N_14816);
and UO_1335 (O_1335,N_14845,N_14666);
and UO_1336 (O_1336,N_14782,N_14683);
and UO_1337 (O_1337,N_14582,N_14549);
nor UO_1338 (O_1338,N_14947,N_14942);
xnor UO_1339 (O_1339,N_14688,N_14847);
xor UO_1340 (O_1340,N_14752,N_14512);
or UO_1341 (O_1341,N_14500,N_14834);
nor UO_1342 (O_1342,N_14945,N_14827);
nor UO_1343 (O_1343,N_14959,N_14721);
nor UO_1344 (O_1344,N_14847,N_14752);
nand UO_1345 (O_1345,N_14718,N_14746);
and UO_1346 (O_1346,N_14664,N_14730);
and UO_1347 (O_1347,N_14538,N_14581);
nor UO_1348 (O_1348,N_14770,N_14738);
or UO_1349 (O_1349,N_14565,N_14965);
or UO_1350 (O_1350,N_14514,N_14511);
xor UO_1351 (O_1351,N_14969,N_14638);
or UO_1352 (O_1352,N_14510,N_14702);
nor UO_1353 (O_1353,N_14813,N_14569);
or UO_1354 (O_1354,N_14533,N_14949);
xnor UO_1355 (O_1355,N_14732,N_14882);
nor UO_1356 (O_1356,N_14663,N_14559);
or UO_1357 (O_1357,N_14941,N_14641);
xnor UO_1358 (O_1358,N_14658,N_14825);
and UO_1359 (O_1359,N_14966,N_14596);
xor UO_1360 (O_1360,N_14724,N_14626);
xnor UO_1361 (O_1361,N_14678,N_14712);
and UO_1362 (O_1362,N_14868,N_14776);
xnor UO_1363 (O_1363,N_14644,N_14586);
and UO_1364 (O_1364,N_14637,N_14509);
nor UO_1365 (O_1365,N_14605,N_14687);
or UO_1366 (O_1366,N_14731,N_14879);
and UO_1367 (O_1367,N_14791,N_14535);
and UO_1368 (O_1368,N_14621,N_14634);
and UO_1369 (O_1369,N_14595,N_14845);
nor UO_1370 (O_1370,N_14690,N_14800);
and UO_1371 (O_1371,N_14742,N_14775);
xor UO_1372 (O_1372,N_14533,N_14610);
and UO_1373 (O_1373,N_14968,N_14933);
nor UO_1374 (O_1374,N_14822,N_14525);
nand UO_1375 (O_1375,N_14800,N_14619);
nand UO_1376 (O_1376,N_14863,N_14822);
nand UO_1377 (O_1377,N_14733,N_14801);
and UO_1378 (O_1378,N_14869,N_14732);
xor UO_1379 (O_1379,N_14854,N_14549);
or UO_1380 (O_1380,N_14504,N_14577);
and UO_1381 (O_1381,N_14936,N_14592);
nand UO_1382 (O_1382,N_14833,N_14516);
xor UO_1383 (O_1383,N_14524,N_14711);
xnor UO_1384 (O_1384,N_14899,N_14972);
nand UO_1385 (O_1385,N_14765,N_14675);
nor UO_1386 (O_1386,N_14982,N_14572);
and UO_1387 (O_1387,N_14842,N_14711);
or UO_1388 (O_1388,N_14696,N_14544);
or UO_1389 (O_1389,N_14680,N_14532);
xor UO_1390 (O_1390,N_14807,N_14565);
nor UO_1391 (O_1391,N_14861,N_14812);
and UO_1392 (O_1392,N_14980,N_14758);
and UO_1393 (O_1393,N_14698,N_14622);
xor UO_1394 (O_1394,N_14862,N_14891);
nand UO_1395 (O_1395,N_14748,N_14993);
nor UO_1396 (O_1396,N_14970,N_14608);
nand UO_1397 (O_1397,N_14584,N_14944);
nand UO_1398 (O_1398,N_14919,N_14657);
xor UO_1399 (O_1399,N_14911,N_14746);
or UO_1400 (O_1400,N_14555,N_14899);
nand UO_1401 (O_1401,N_14697,N_14713);
and UO_1402 (O_1402,N_14912,N_14966);
and UO_1403 (O_1403,N_14508,N_14555);
and UO_1404 (O_1404,N_14582,N_14633);
and UO_1405 (O_1405,N_14561,N_14666);
or UO_1406 (O_1406,N_14996,N_14529);
xor UO_1407 (O_1407,N_14918,N_14904);
xnor UO_1408 (O_1408,N_14712,N_14770);
xor UO_1409 (O_1409,N_14782,N_14797);
nand UO_1410 (O_1410,N_14791,N_14720);
xor UO_1411 (O_1411,N_14624,N_14777);
nand UO_1412 (O_1412,N_14872,N_14803);
or UO_1413 (O_1413,N_14943,N_14608);
nand UO_1414 (O_1414,N_14662,N_14748);
or UO_1415 (O_1415,N_14799,N_14784);
xnor UO_1416 (O_1416,N_14706,N_14818);
or UO_1417 (O_1417,N_14859,N_14845);
nand UO_1418 (O_1418,N_14688,N_14756);
xnor UO_1419 (O_1419,N_14905,N_14886);
xnor UO_1420 (O_1420,N_14957,N_14907);
and UO_1421 (O_1421,N_14836,N_14829);
nand UO_1422 (O_1422,N_14924,N_14597);
or UO_1423 (O_1423,N_14783,N_14754);
nand UO_1424 (O_1424,N_14821,N_14693);
nand UO_1425 (O_1425,N_14526,N_14713);
nand UO_1426 (O_1426,N_14583,N_14649);
xnor UO_1427 (O_1427,N_14505,N_14869);
or UO_1428 (O_1428,N_14723,N_14640);
nand UO_1429 (O_1429,N_14556,N_14534);
or UO_1430 (O_1430,N_14767,N_14822);
nor UO_1431 (O_1431,N_14738,N_14665);
xor UO_1432 (O_1432,N_14913,N_14611);
xnor UO_1433 (O_1433,N_14699,N_14553);
or UO_1434 (O_1434,N_14786,N_14840);
and UO_1435 (O_1435,N_14789,N_14959);
or UO_1436 (O_1436,N_14887,N_14931);
xnor UO_1437 (O_1437,N_14776,N_14701);
or UO_1438 (O_1438,N_14576,N_14997);
nand UO_1439 (O_1439,N_14653,N_14898);
or UO_1440 (O_1440,N_14556,N_14733);
and UO_1441 (O_1441,N_14887,N_14631);
or UO_1442 (O_1442,N_14906,N_14979);
and UO_1443 (O_1443,N_14851,N_14828);
or UO_1444 (O_1444,N_14638,N_14876);
nor UO_1445 (O_1445,N_14656,N_14830);
nand UO_1446 (O_1446,N_14960,N_14854);
or UO_1447 (O_1447,N_14723,N_14501);
nand UO_1448 (O_1448,N_14597,N_14963);
xor UO_1449 (O_1449,N_14841,N_14571);
nand UO_1450 (O_1450,N_14871,N_14929);
xor UO_1451 (O_1451,N_14687,N_14749);
or UO_1452 (O_1452,N_14790,N_14705);
nor UO_1453 (O_1453,N_14939,N_14718);
or UO_1454 (O_1454,N_14933,N_14916);
xor UO_1455 (O_1455,N_14595,N_14503);
or UO_1456 (O_1456,N_14749,N_14547);
or UO_1457 (O_1457,N_14843,N_14653);
xnor UO_1458 (O_1458,N_14702,N_14946);
nor UO_1459 (O_1459,N_14982,N_14723);
and UO_1460 (O_1460,N_14909,N_14989);
nand UO_1461 (O_1461,N_14968,N_14838);
nor UO_1462 (O_1462,N_14558,N_14500);
nand UO_1463 (O_1463,N_14793,N_14672);
and UO_1464 (O_1464,N_14680,N_14970);
nor UO_1465 (O_1465,N_14890,N_14508);
or UO_1466 (O_1466,N_14590,N_14711);
nor UO_1467 (O_1467,N_14603,N_14583);
and UO_1468 (O_1468,N_14718,N_14711);
xnor UO_1469 (O_1469,N_14966,N_14707);
or UO_1470 (O_1470,N_14664,N_14767);
and UO_1471 (O_1471,N_14827,N_14514);
or UO_1472 (O_1472,N_14714,N_14776);
xor UO_1473 (O_1473,N_14773,N_14905);
nor UO_1474 (O_1474,N_14538,N_14539);
xnor UO_1475 (O_1475,N_14505,N_14545);
nor UO_1476 (O_1476,N_14951,N_14636);
nand UO_1477 (O_1477,N_14589,N_14891);
nor UO_1478 (O_1478,N_14801,N_14682);
and UO_1479 (O_1479,N_14517,N_14869);
nor UO_1480 (O_1480,N_14897,N_14758);
or UO_1481 (O_1481,N_14884,N_14703);
xor UO_1482 (O_1482,N_14613,N_14551);
nor UO_1483 (O_1483,N_14714,N_14636);
or UO_1484 (O_1484,N_14604,N_14600);
xnor UO_1485 (O_1485,N_14992,N_14926);
xnor UO_1486 (O_1486,N_14519,N_14955);
nor UO_1487 (O_1487,N_14978,N_14941);
or UO_1488 (O_1488,N_14953,N_14816);
nand UO_1489 (O_1489,N_14686,N_14690);
or UO_1490 (O_1490,N_14685,N_14501);
nor UO_1491 (O_1491,N_14916,N_14822);
nand UO_1492 (O_1492,N_14914,N_14962);
and UO_1493 (O_1493,N_14559,N_14693);
nand UO_1494 (O_1494,N_14589,N_14738);
nand UO_1495 (O_1495,N_14601,N_14655);
or UO_1496 (O_1496,N_14553,N_14890);
nor UO_1497 (O_1497,N_14812,N_14537);
and UO_1498 (O_1498,N_14713,N_14780);
nand UO_1499 (O_1499,N_14783,N_14968);
nand UO_1500 (O_1500,N_14620,N_14695);
xnor UO_1501 (O_1501,N_14929,N_14975);
and UO_1502 (O_1502,N_14981,N_14794);
and UO_1503 (O_1503,N_14618,N_14792);
nand UO_1504 (O_1504,N_14631,N_14574);
nor UO_1505 (O_1505,N_14990,N_14513);
or UO_1506 (O_1506,N_14771,N_14859);
xor UO_1507 (O_1507,N_14676,N_14742);
nor UO_1508 (O_1508,N_14894,N_14795);
or UO_1509 (O_1509,N_14873,N_14698);
or UO_1510 (O_1510,N_14546,N_14677);
xnor UO_1511 (O_1511,N_14716,N_14610);
or UO_1512 (O_1512,N_14613,N_14855);
or UO_1513 (O_1513,N_14641,N_14727);
nand UO_1514 (O_1514,N_14976,N_14875);
nor UO_1515 (O_1515,N_14599,N_14749);
xnor UO_1516 (O_1516,N_14873,N_14558);
nand UO_1517 (O_1517,N_14886,N_14786);
nand UO_1518 (O_1518,N_14800,N_14514);
and UO_1519 (O_1519,N_14634,N_14764);
nor UO_1520 (O_1520,N_14799,N_14854);
nand UO_1521 (O_1521,N_14840,N_14609);
nor UO_1522 (O_1522,N_14699,N_14735);
or UO_1523 (O_1523,N_14936,N_14909);
or UO_1524 (O_1524,N_14814,N_14953);
or UO_1525 (O_1525,N_14896,N_14897);
and UO_1526 (O_1526,N_14615,N_14534);
nand UO_1527 (O_1527,N_14998,N_14510);
nand UO_1528 (O_1528,N_14747,N_14944);
and UO_1529 (O_1529,N_14905,N_14704);
nand UO_1530 (O_1530,N_14814,N_14930);
or UO_1531 (O_1531,N_14517,N_14875);
nor UO_1532 (O_1532,N_14560,N_14921);
nand UO_1533 (O_1533,N_14708,N_14974);
nor UO_1534 (O_1534,N_14783,N_14878);
nor UO_1535 (O_1535,N_14575,N_14852);
and UO_1536 (O_1536,N_14669,N_14747);
nand UO_1537 (O_1537,N_14938,N_14991);
nor UO_1538 (O_1538,N_14598,N_14828);
nand UO_1539 (O_1539,N_14951,N_14554);
or UO_1540 (O_1540,N_14832,N_14556);
and UO_1541 (O_1541,N_14916,N_14943);
and UO_1542 (O_1542,N_14767,N_14684);
nor UO_1543 (O_1543,N_14641,N_14934);
nor UO_1544 (O_1544,N_14556,N_14557);
nor UO_1545 (O_1545,N_14691,N_14760);
or UO_1546 (O_1546,N_14841,N_14602);
nand UO_1547 (O_1547,N_14902,N_14727);
nand UO_1548 (O_1548,N_14742,N_14636);
nand UO_1549 (O_1549,N_14809,N_14692);
and UO_1550 (O_1550,N_14544,N_14993);
or UO_1551 (O_1551,N_14972,N_14969);
xnor UO_1552 (O_1552,N_14532,N_14865);
nand UO_1553 (O_1553,N_14716,N_14833);
nand UO_1554 (O_1554,N_14734,N_14885);
nor UO_1555 (O_1555,N_14961,N_14897);
xor UO_1556 (O_1556,N_14541,N_14786);
xnor UO_1557 (O_1557,N_14550,N_14776);
xnor UO_1558 (O_1558,N_14575,N_14612);
nand UO_1559 (O_1559,N_14798,N_14579);
xor UO_1560 (O_1560,N_14622,N_14585);
xor UO_1561 (O_1561,N_14775,N_14675);
xnor UO_1562 (O_1562,N_14553,N_14728);
and UO_1563 (O_1563,N_14862,N_14519);
xnor UO_1564 (O_1564,N_14947,N_14744);
or UO_1565 (O_1565,N_14813,N_14505);
and UO_1566 (O_1566,N_14974,N_14789);
and UO_1567 (O_1567,N_14652,N_14803);
nand UO_1568 (O_1568,N_14998,N_14727);
and UO_1569 (O_1569,N_14727,N_14857);
nand UO_1570 (O_1570,N_14880,N_14789);
and UO_1571 (O_1571,N_14511,N_14972);
nand UO_1572 (O_1572,N_14831,N_14932);
or UO_1573 (O_1573,N_14926,N_14670);
and UO_1574 (O_1574,N_14657,N_14740);
xor UO_1575 (O_1575,N_14507,N_14983);
nor UO_1576 (O_1576,N_14631,N_14625);
xnor UO_1577 (O_1577,N_14568,N_14665);
nor UO_1578 (O_1578,N_14906,N_14916);
nor UO_1579 (O_1579,N_14798,N_14746);
and UO_1580 (O_1580,N_14784,N_14512);
or UO_1581 (O_1581,N_14682,N_14639);
nor UO_1582 (O_1582,N_14790,N_14807);
xnor UO_1583 (O_1583,N_14801,N_14731);
nand UO_1584 (O_1584,N_14700,N_14605);
nand UO_1585 (O_1585,N_14567,N_14766);
nor UO_1586 (O_1586,N_14904,N_14981);
xnor UO_1587 (O_1587,N_14842,N_14613);
xor UO_1588 (O_1588,N_14681,N_14614);
xnor UO_1589 (O_1589,N_14572,N_14694);
nand UO_1590 (O_1590,N_14575,N_14585);
xor UO_1591 (O_1591,N_14922,N_14837);
nor UO_1592 (O_1592,N_14571,N_14951);
or UO_1593 (O_1593,N_14857,N_14919);
nand UO_1594 (O_1594,N_14720,N_14553);
and UO_1595 (O_1595,N_14974,N_14898);
nor UO_1596 (O_1596,N_14908,N_14544);
nand UO_1597 (O_1597,N_14976,N_14677);
and UO_1598 (O_1598,N_14908,N_14998);
or UO_1599 (O_1599,N_14892,N_14642);
nor UO_1600 (O_1600,N_14640,N_14884);
nor UO_1601 (O_1601,N_14847,N_14920);
and UO_1602 (O_1602,N_14540,N_14586);
or UO_1603 (O_1603,N_14777,N_14693);
xnor UO_1604 (O_1604,N_14797,N_14825);
and UO_1605 (O_1605,N_14956,N_14518);
nand UO_1606 (O_1606,N_14981,N_14806);
nor UO_1607 (O_1607,N_14839,N_14500);
nand UO_1608 (O_1608,N_14838,N_14852);
nor UO_1609 (O_1609,N_14613,N_14824);
xnor UO_1610 (O_1610,N_14648,N_14569);
or UO_1611 (O_1611,N_14531,N_14894);
and UO_1612 (O_1612,N_14922,N_14598);
and UO_1613 (O_1613,N_14869,N_14819);
nand UO_1614 (O_1614,N_14589,N_14605);
or UO_1615 (O_1615,N_14557,N_14756);
nor UO_1616 (O_1616,N_14822,N_14543);
xor UO_1617 (O_1617,N_14996,N_14741);
nor UO_1618 (O_1618,N_14957,N_14920);
xnor UO_1619 (O_1619,N_14856,N_14762);
nand UO_1620 (O_1620,N_14792,N_14555);
or UO_1621 (O_1621,N_14996,N_14601);
and UO_1622 (O_1622,N_14516,N_14793);
and UO_1623 (O_1623,N_14521,N_14942);
or UO_1624 (O_1624,N_14932,N_14988);
nand UO_1625 (O_1625,N_14926,N_14819);
nor UO_1626 (O_1626,N_14780,N_14727);
and UO_1627 (O_1627,N_14573,N_14606);
xor UO_1628 (O_1628,N_14964,N_14617);
and UO_1629 (O_1629,N_14725,N_14966);
or UO_1630 (O_1630,N_14914,N_14788);
nand UO_1631 (O_1631,N_14769,N_14546);
nor UO_1632 (O_1632,N_14530,N_14617);
and UO_1633 (O_1633,N_14874,N_14542);
xor UO_1634 (O_1634,N_14743,N_14849);
nand UO_1635 (O_1635,N_14807,N_14795);
and UO_1636 (O_1636,N_14708,N_14815);
xnor UO_1637 (O_1637,N_14671,N_14630);
or UO_1638 (O_1638,N_14883,N_14544);
nor UO_1639 (O_1639,N_14618,N_14649);
and UO_1640 (O_1640,N_14901,N_14722);
nand UO_1641 (O_1641,N_14863,N_14830);
nor UO_1642 (O_1642,N_14800,N_14651);
or UO_1643 (O_1643,N_14884,N_14603);
nand UO_1644 (O_1644,N_14901,N_14886);
or UO_1645 (O_1645,N_14781,N_14922);
nand UO_1646 (O_1646,N_14966,N_14623);
or UO_1647 (O_1647,N_14711,N_14890);
and UO_1648 (O_1648,N_14789,N_14643);
nor UO_1649 (O_1649,N_14996,N_14913);
or UO_1650 (O_1650,N_14667,N_14596);
xor UO_1651 (O_1651,N_14993,N_14741);
nor UO_1652 (O_1652,N_14793,N_14840);
xnor UO_1653 (O_1653,N_14642,N_14995);
nand UO_1654 (O_1654,N_14854,N_14529);
or UO_1655 (O_1655,N_14660,N_14831);
and UO_1656 (O_1656,N_14984,N_14907);
and UO_1657 (O_1657,N_14505,N_14843);
nor UO_1658 (O_1658,N_14552,N_14935);
or UO_1659 (O_1659,N_14601,N_14696);
nand UO_1660 (O_1660,N_14778,N_14753);
nand UO_1661 (O_1661,N_14543,N_14750);
and UO_1662 (O_1662,N_14992,N_14694);
and UO_1663 (O_1663,N_14690,N_14782);
nor UO_1664 (O_1664,N_14862,N_14525);
nand UO_1665 (O_1665,N_14765,N_14542);
nand UO_1666 (O_1666,N_14999,N_14751);
nand UO_1667 (O_1667,N_14903,N_14922);
nor UO_1668 (O_1668,N_14735,N_14943);
nand UO_1669 (O_1669,N_14795,N_14796);
or UO_1670 (O_1670,N_14660,N_14601);
nand UO_1671 (O_1671,N_14614,N_14765);
or UO_1672 (O_1672,N_14564,N_14636);
nor UO_1673 (O_1673,N_14696,N_14504);
nor UO_1674 (O_1674,N_14725,N_14652);
nor UO_1675 (O_1675,N_14800,N_14806);
or UO_1676 (O_1676,N_14820,N_14775);
xnor UO_1677 (O_1677,N_14567,N_14502);
and UO_1678 (O_1678,N_14801,N_14946);
nor UO_1679 (O_1679,N_14941,N_14828);
and UO_1680 (O_1680,N_14970,N_14657);
nor UO_1681 (O_1681,N_14659,N_14661);
and UO_1682 (O_1682,N_14687,N_14698);
and UO_1683 (O_1683,N_14866,N_14599);
nand UO_1684 (O_1684,N_14792,N_14675);
nor UO_1685 (O_1685,N_14636,N_14633);
nor UO_1686 (O_1686,N_14935,N_14544);
xor UO_1687 (O_1687,N_14794,N_14517);
or UO_1688 (O_1688,N_14538,N_14528);
and UO_1689 (O_1689,N_14928,N_14917);
nor UO_1690 (O_1690,N_14806,N_14843);
nand UO_1691 (O_1691,N_14658,N_14965);
and UO_1692 (O_1692,N_14722,N_14639);
or UO_1693 (O_1693,N_14527,N_14583);
nor UO_1694 (O_1694,N_14919,N_14935);
or UO_1695 (O_1695,N_14734,N_14556);
nand UO_1696 (O_1696,N_14954,N_14618);
or UO_1697 (O_1697,N_14584,N_14658);
xor UO_1698 (O_1698,N_14590,N_14545);
nand UO_1699 (O_1699,N_14519,N_14836);
nand UO_1700 (O_1700,N_14534,N_14933);
or UO_1701 (O_1701,N_14734,N_14616);
xnor UO_1702 (O_1702,N_14982,N_14954);
and UO_1703 (O_1703,N_14888,N_14599);
xor UO_1704 (O_1704,N_14680,N_14639);
and UO_1705 (O_1705,N_14538,N_14610);
and UO_1706 (O_1706,N_14872,N_14955);
and UO_1707 (O_1707,N_14747,N_14717);
or UO_1708 (O_1708,N_14887,N_14881);
and UO_1709 (O_1709,N_14822,N_14872);
nor UO_1710 (O_1710,N_14621,N_14612);
or UO_1711 (O_1711,N_14617,N_14692);
and UO_1712 (O_1712,N_14947,N_14770);
and UO_1713 (O_1713,N_14609,N_14688);
xnor UO_1714 (O_1714,N_14772,N_14548);
or UO_1715 (O_1715,N_14641,N_14681);
nand UO_1716 (O_1716,N_14544,N_14709);
xor UO_1717 (O_1717,N_14694,N_14835);
xnor UO_1718 (O_1718,N_14926,N_14965);
xnor UO_1719 (O_1719,N_14940,N_14835);
nand UO_1720 (O_1720,N_14977,N_14562);
nor UO_1721 (O_1721,N_14595,N_14622);
nor UO_1722 (O_1722,N_14963,N_14508);
or UO_1723 (O_1723,N_14606,N_14559);
nor UO_1724 (O_1724,N_14825,N_14871);
and UO_1725 (O_1725,N_14793,N_14842);
or UO_1726 (O_1726,N_14834,N_14863);
nor UO_1727 (O_1727,N_14843,N_14740);
nand UO_1728 (O_1728,N_14585,N_14990);
nand UO_1729 (O_1729,N_14891,N_14677);
xnor UO_1730 (O_1730,N_14817,N_14946);
or UO_1731 (O_1731,N_14877,N_14585);
xor UO_1732 (O_1732,N_14592,N_14724);
nor UO_1733 (O_1733,N_14999,N_14699);
nor UO_1734 (O_1734,N_14928,N_14856);
nor UO_1735 (O_1735,N_14533,N_14828);
nor UO_1736 (O_1736,N_14539,N_14738);
and UO_1737 (O_1737,N_14558,N_14697);
nor UO_1738 (O_1738,N_14628,N_14797);
and UO_1739 (O_1739,N_14598,N_14989);
or UO_1740 (O_1740,N_14541,N_14709);
nand UO_1741 (O_1741,N_14854,N_14841);
nand UO_1742 (O_1742,N_14896,N_14514);
xor UO_1743 (O_1743,N_14602,N_14650);
and UO_1744 (O_1744,N_14562,N_14839);
xnor UO_1745 (O_1745,N_14850,N_14686);
xor UO_1746 (O_1746,N_14856,N_14596);
or UO_1747 (O_1747,N_14599,N_14907);
nand UO_1748 (O_1748,N_14628,N_14500);
nor UO_1749 (O_1749,N_14630,N_14767);
nand UO_1750 (O_1750,N_14745,N_14593);
and UO_1751 (O_1751,N_14888,N_14549);
nand UO_1752 (O_1752,N_14591,N_14585);
nand UO_1753 (O_1753,N_14544,N_14644);
nand UO_1754 (O_1754,N_14919,N_14667);
nor UO_1755 (O_1755,N_14648,N_14989);
xnor UO_1756 (O_1756,N_14508,N_14842);
and UO_1757 (O_1757,N_14666,N_14871);
xnor UO_1758 (O_1758,N_14871,N_14966);
nand UO_1759 (O_1759,N_14641,N_14848);
and UO_1760 (O_1760,N_14960,N_14948);
nand UO_1761 (O_1761,N_14718,N_14938);
and UO_1762 (O_1762,N_14710,N_14861);
and UO_1763 (O_1763,N_14774,N_14907);
nor UO_1764 (O_1764,N_14918,N_14798);
and UO_1765 (O_1765,N_14774,N_14747);
and UO_1766 (O_1766,N_14866,N_14611);
xor UO_1767 (O_1767,N_14806,N_14965);
xor UO_1768 (O_1768,N_14924,N_14901);
xnor UO_1769 (O_1769,N_14809,N_14893);
xor UO_1770 (O_1770,N_14572,N_14704);
nor UO_1771 (O_1771,N_14808,N_14916);
nor UO_1772 (O_1772,N_14757,N_14940);
xor UO_1773 (O_1773,N_14706,N_14635);
nor UO_1774 (O_1774,N_14753,N_14880);
or UO_1775 (O_1775,N_14984,N_14716);
nand UO_1776 (O_1776,N_14711,N_14588);
and UO_1777 (O_1777,N_14695,N_14697);
nand UO_1778 (O_1778,N_14971,N_14885);
nand UO_1779 (O_1779,N_14519,N_14788);
xor UO_1780 (O_1780,N_14719,N_14720);
or UO_1781 (O_1781,N_14934,N_14766);
or UO_1782 (O_1782,N_14732,N_14782);
nand UO_1783 (O_1783,N_14704,N_14620);
xnor UO_1784 (O_1784,N_14780,N_14735);
or UO_1785 (O_1785,N_14681,N_14647);
and UO_1786 (O_1786,N_14629,N_14897);
or UO_1787 (O_1787,N_14583,N_14810);
nand UO_1788 (O_1788,N_14509,N_14748);
xnor UO_1789 (O_1789,N_14892,N_14815);
xor UO_1790 (O_1790,N_14899,N_14985);
or UO_1791 (O_1791,N_14894,N_14744);
xor UO_1792 (O_1792,N_14747,N_14821);
or UO_1793 (O_1793,N_14784,N_14586);
and UO_1794 (O_1794,N_14768,N_14598);
and UO_1795 (O_1795,N_14553,N_14878);
and UO_1796 (O_1796,N_14872,N_14675);
xor UO_1797 (O_1797,N_14750,N_14673);
nand UO_1798 (O_1798,N_14968,N_14977);
or UO_1799 (O_1799,N_14725,N_14616);
nand UO_1800 (O_1800,N_14702,N_14863);
and UO_1801 (O_1801,N_14870,N_14784);
or UO_1802 (O_1802,N_14525,N_14760);
or UO_1803 (O_1803,N_14838,N_14983);
and UO_1804 (O_1804,N_14589,N_14992);
or UO_1805 (O_1805,N_14971,N_14558);
nor UO_1806 (O_1806,N_14654,N_14851);
xor UO_1807 (O_1807,N_14575,N_14533);
xnor UO_1808 (O_1808,N_14719,N_14960);
xnor UO_1809 (O_1809,N_14873,N_14970);
and UO_1810 (O_1810,N_14688,N_14692);
nor UO_1811 (O_1811,N_14608,N_14880);
and UO_1812 (O_1812,N_14567,N_14715);
nand UO_1813 (O_1813,N_14832,N_14719);
nor UO_1814 (O_1814,N_14525,N_14579);
or UO_1815 (O_1815,N_14965,N_14996);
nand UO_1816 (O_1816,N_14539,N_14974);
nand UO_1817 (O_1817,N_14866,N_14673);
nor UO_1818 (O_1818,N_14860,N_14925);
nand UO_1819 (O_1819,N_14695,N_14870);
or UO_1820 (O_1820,N_14603,N_14823);
and UO_1821 (O_1821,N_14828,N_14762);
nand UO_1822 (O_1822,N_14632,N_14798);
nand UO_1823 (O_1823,N_14705,N_14620);
and UO_1824 (O_1824,N_14930,N_14823);
nand UO_1825 (O_1825,N_14598,N_14730);
nor UO_1826 (O_1826,N_14527,N_14618);
nor UO_1827 (O_1827,N_14854,N_14508);
or UO_1828 (O_1828,N_14628,N_14615);
nor UO_1829 (O_1829,N_14713,N_14666);
nand UO_1830 (O_1830,N_14828,N_14837);
nand UO_1831 (O_1831,N_14911,N_14520);
nand UO_1832 (O_1832,N_14590,N_14816);
and UO_1833 (O_1833,N_14646,N_14602);
or UO_1834 (O_1834,N_14743,N_14610);
nand UO_1835 (O_1835,N_14523,N_14530);
and UO_1836 (O_1836,N_14697,N_14504);
xor UO_1837 (O_1837,N_14715,N_14897);
or UO_1838 (O_1838,N_14720,N_14770);
xor UO_1839 (O_1839,N_14846,N_14901);
or UO_1840 (O_1840,N_14843,N_14509);
or UO_1841 (O_1841,N_14979,N_14520);
or UO_1842 (O_1842,N_14803,N_14802);
nor UO_1843 (O_1843,N_14949,N_14979);
or UO_1844 (O_1844,N_14749,N_14973);
nor UO_1845 (O_1845,N_14629,N_14713);
nand UO_1846 (O_1846,N_14856,N_14631);
or UO_1847 (O_1847,N_14599,N_14686);
nor UO_1848 (O_1848,N_14842,N_14645);
nand UO_1849 (O_1849,N_14514,N_14722);
and UO_1850 (O_1850,N_14952,N_14747);
xor UO_1851 (O_1851,N_14735,N_14521);
nor UO_1852 (O_1852,N_14718,N_14713);
nor UO_1853 (O_1853,N_14942,N_14608);
xor UO_1854 (O_1854,N_14803,N_14793);
or UO_1855 (O_1855,N_14881,N_14611);
and UO_1856 (O_1856,N_14752,N_14500);
nand UO_1857 (O_1857,N_14685,N_14916);
nor UO_1858 (O_1858,N_14904,N_14844);
xnor UO_1859 (O_1859,N_14991,N_14974);
or UO_1860 (O_1860,N_14888,N_14503);
and UO_1861 (O_1861,N_14731,N_14577);
nor UO_1862 (O_1862,N_14819,N_14547);
xnor UO_1863 (O_1863,N_14710,N_14623);
nand UO_1864 (O_1864,N_14781,N_14933);
and UO_1865 (O_1865,N_14896,N_14931);
nor UO_1866 (O_1866,N_14990,N_14698);
nor UO_1867 (O_1867,N_14837,N_14645);
nor UO_1868 (O_1868,N_14641,N_14796);
xnor UO_1869 (O_1869,N_14995,N_14982);
and UO_1870 (O_1870,N_14903,N_14968);
nor UO_1871 (O_1871,N_14527,N_14612);
or UO_1872 (O_1872,N_14546,N_14752);
or UO_1873 (O_1873,N_14622,N_14839);
xor UO_1874 (O_1874,N_14736,N_14994);
xnor UO_1875 (O_1875,N_14656,N_14816);
xnor UO_1876 (O_1876,N_14715,N_14868);
nor UO_1877 (O_1877,N_14953,N_14975);
and UO_1878 (O_1878,N_14868,N_14624);
nor UO_1879 (O_1879,N_14662,N_14933);
xnor UO_1880 (O_1880,N_14543,N_14713);
and UO_1881 (O_1881,N_14632,N_14806);
or UO_1882 (O_1882,N_14552,N_14712);
xor UO_1883 (O_1883,N_14582,N_14941);
nor UO_1884 (O_1884,N_14955,N_14745);
nand UO_1885 (O_1885,N_14774,N_14911);
xnor UO_1886 (O_1886,N_14908,N_14618);
nor UO_1887 (O_1887,N_14849,N_14759);
and UO_1888 (O_1888,N_14719,N_14884);
xor UO_1889 (O_1889,N_14536,N_14821);
nand UO_1890 (O_1890,N_14559,N_14839);
or UO_1891 (O_1891,N_14799,N_14745);
nor UO_1892 (O_1892,N_14680,N_14540);
nand UO_1893 (O_1893,N_14674,N_14739);
or UO_1894 (O_1894,N_14934,N_14549);
and UO_1895 (O_1895,N_14689,N_14971);
and UO_1896 (O_1896,N_14872,N_14950);
nor UO_1897 (O_1897,N_14786,N_14938);
and UO_1898 (O_1898,N_14993,N_14695);
and UO_1899 (O_1899,N_14570,N_14925);
or UO_1900 (O_1900,N_14610,N_14790);
nor UO_1901 (O_1901,N_14626,N_14512);
nor UO_1902 (O_1902,N_14804,N_14843);
or UO_1903 (O_1903,N_14798,N_14614);
and UO_1904 (O_1904,N_14935,N_14594);
or UO_1905 (O_1905,N_14613,N_14943);
nor UO_1906 (O_1906,N_14725,N_14946);
or UO_1907 (O_1907,N_14640,N_14969);
and UO_1908 (O_1908,N_14961,N_14586);
and UO_1909 (O_1909,N_14569,N_14525);
nand UO_1910 (O_1910,N_14598,N_14939);
nand UO_1911 (O_1911,N_14878,N_14640);
nor UO_1912 (O_1912,N_14884,N_14920);
nand UO_1913 (O_1913,N_14517,N_14841);
nand UO_1914 (O_1914,N_14855,N_14614);
nor UO_1915 (O_1915,N_14601,N_14642);
nor UO_1916 (O_1916,N_14954,N_14654);
or UO_1917 (O_1917,N_14777,N_14654);
or UO_1918 (O_1918,N_14586,N_14702);
and UO_1919 (O_1919,N_14896,N_14743);
xnor UO_1920 (O_1920,N_14597,N_14659);
nand UO_1921 (O_1921,N_14730,N_14557);
nor UO_1922 (O_1922,N_14843,N_14912);
and UO_1923 (O_1923,N_14739,N_14619);
or UO_1924 (O_1924,N_14762,N_14929);
or UO_1925 (O_1925,N_14624,N_14755);
nand UO_1926 (O_1926,N_14688,N_14816);
nor UO_1927 (O_1927,N_14666,N_14764);
and UO_1928 (O_1928,N_14981,N_14548);
or UO_1929 (O_1929,N_14621,N_14684);
and UO_1930 (O_1930,N_14736,N_14595);
xnor UO_1931 (O_1931,N_14547,N_14539);
or UO_1932 (O_1932,N_14971,N_14787);
or UO_1933 (O_1933,N_14748,N_14679);
xor UO_1934 (O_1934,N_14939,N_14594);
nand UO_1935 (O_1935,N_14722,N_14540);
nand UO_1936 (O_1936,N_14577,N_14937);
nor UO_1937 (O_1937,N_14699,N_14571);
xor UO_1938 (O_1938,N_14755,N_14807);
and UO_1939 (O_1939,N_14856,N_14755);
xor UO_1940 (O_1940,N_14534,N_14903);
nand UO_1941 (O_1941,N_14970,N_14780);
xnor UO_1942 (O_1942,N_14612,N_14693);
nor UO_1943 (O_1943,N_14642,N_14926);
or UO_1944 (O_1944,N_14898,N_14752);
or UO_1945 (O_1945,N_14694,N_14959);
nand UO_1946 (O_1946,N_14823,N_14990);
nand UO_1947 (O_1947,N_14767,N_14788);
nand UO_1948 (O_1948,N_14616,N_14730);
and UO_1949 (O_1949,N_14927,N_14972);
or UO_1950 (O_1950,N_14791,N_14898);
nor UO_1951 (O_1951,N_14814,N_14660);
xnor UO_1952 (O_1952,N_14744,N_14871);
xor UO_1953 (O_1953,N_14764,N_14842);
xnor UO_1954 (O_1954,N_14696,N_14526);
or UO_1955 (O_1955,N_14643,N_14899);
and UO_1956 (O_1956,N_14876,N_14742);
and UO_1957 (O_1957,N_14635,N_14569);
and UO_1958 (O_1958,N_14757,N_14889);
nor UO_1959 (O_1959,N_14743,N_14923);
nand UO_1960 (O_1960,N_14845,N_14972);
nand UO_1961 (O_1961,N_14639,N_14909);
or UO_1962 (O_1962,N_14812,N_14874);
nor UO_1963 (O_1963,N_14760,N_14979);
nand UO_1964 (O_1964,N_14872,N_14831);
xor UO_1965 (O_1965,N_14658,N_14998);
nor UO_1966 (O_1966,N_14541,N_14816);
nor UO_1967 (O_1967,N_14691,N_14767);
nand UO_1968 (O_1968,N_14547,N_14873);
xor UO_1969 (O_1969,N_14836,N_14511);
xnor UO_1970 (O_1970,N_14534,N_14874);
xor UO_1971 (O_1971,N_14861,N_14810);
nand UO_1972 (O_1972,N_14969,N_14623);
xor UO_1973 (O_1973,N_14947,N_14884);
nor UO_1974 (O_1974,N_14966,N_14686);
xor UO_1975 (O_1975,N_14750,N_14677);
or UO_1976 (O_1976,N_14560,N_14910);
xor UO_1977 (O_1977,N_14754,N_14583);
nor UO_1978 (O_1978,N_14559,N_14819);
xor UO_1979 (O_1979,N_14524,N_14712);
nor UO_1980 (O_1980,N_14911,N_14788);
xnor UO_1981 (O_1981,N_14864,N_14521);
nor UO_1982 (O_1982,N_14516,N_14574);
or UO_1983 (O_1983,N_14877,N_14868);
xor UO_1984 (O_1984,N_14791,N_14581);
nand UO_1985 (O_1985,N_14733,N_14673);
nand UO_1986 (O_1986,N_14935,N_14728);
nor UO_1987 (O_1987,N_14899,N_14940);
and UO_1988 (O_1988,N_14730,N_14861);
and UO_1989 (O_1989,N_14554,N_14536);
and UO_1990 (O_1990,N_14645,N_14945);
nor UO_1991 (O_1991,N_14905,N_14535);
nor UO_1992 (O_1992,N_14717,N_14513);
and UO_1993 (O_1993,N_14669,N_14525);
or UO_1994 (O_1994,N_14615,N_14504);
nand UO_1995 (O_1995,N_14885,N_14835);
and UO_1996 (O_1996,N_14919,N_14831);
xnor UO_1997 (O_1997,N_14918,N_14575);
nor UO_1998 (O_1998,N_14710,N_14686);
nand UO_1999 (O_1999,N_14829,N_14633);
endmodule