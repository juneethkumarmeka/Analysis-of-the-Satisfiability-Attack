module basic_750_5000_1000_5_levels_2xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nor U0 (N_0,In_254,In_551);
nor U1 (N_1,In_713,In_99);
and U2 (N_2,In_539,In_447);
nor U3 (N_3,In_352,In_624);
or U4 (N_4,In_157,In_143);
nand U5 (N_5,In_717,In_298);
nor U6 (N_6,In_31,In_708);
and U7 (N_7,In_586,In_477);
or U8 (N_8,In_324,In_715);
nand U9 (N_9,In_230,In_608);
nor U10 (N_10,In_361,In_735);
or U11 (N_11,In_236,In_259);
and U12 (N_12,In_538,In_472);
nand U13 (N_13,In_503,In_355);
and U14 (N_14,In_504,In_532);
nor U15 (N_15,In_332,In_674);
xor U16 (N_16,In_574,In_408);
or U17 (N_17,In_556,In_58);
or U18 (N_18,In_493,In_716);
or U19 (N_19,In_393,In_125);
or U20 (N_20,In_321,In_738);
nor U21 (N_21,In_359,In_670);
nand U22 (N_22,In_64,In_225);
or U23 (N_23,In_198,In_304);
and U24 (N_24,In_212,In_579);
or U25 (N_25,In_741,In_368);
nor U26 (N_26,In_244,In_197);
and U27 (N_27,In_592,In_126);
or U28 (N_28,In_686,In_612);
nor U29 (N_29,In_333,In_17);
nor U30 (N_30,In_296,In_326);
and U31 (N_31,In_164,In_475);
and U32 (N_32,In_264,In_168);
and U33 (N_33,In_48,In_144);
and U34 (N_34,In_20,In_505);
nor U35 (N_35,In_680,In_93);
or U36 (N_36,In_522,In_402);
and U37 (N_37,In_367,In_242);
xor U38 (N_38,In_513,In_4);
or U39 (N_39,In_258,In_293);
and U40 (N_40,In_16,In_709);
nor U41 (N_41,In_598,In_620);
nand U42 (N_42,In_691,In_671);
nor U43 (N_43,In_678,In_241);
or U44 (N_44,In_578,In_446);
or U45 (N_45,In_512,In_582);
nand U46 (N_46,In_165,In_481);
and U47 (N_47,In_457,In_497);
nand U48 (N_48,In_452,In_290);
nor U49 (N_49,In_596,In_123);
nor U50 (N_50,In_473,In_737);
nor U51 (N_51,In_181,In_590);
or U52 (N_52,In_461,In_748);
nor U53 (N_53,In_410,In_185);
nor U54 (N_54,In_435,In_414);
nor U55 (N_55,In_372,In_15);
and U56 (N_56,In_621,In_224);
or U57 (N_57,In_138,In_635);
or U58 (N_58,In_378,In_413);
and U59 (N_59,In_279,In_134);
and U60 (N_60,In_26,In_38);
nor U61 (N_61,In_336,In_525);
nor U62 (N_62,In_394,In_456);
nand U63 (N_63,In_191,In_631);
or U64 (N_64,In_733,In_644);
and U65 (N_65,In_662,In_445);
nor U66 (N_66,In_221,In_439);
nand U67 (N_67,In_59,In_309);
xnor U68 (N_68,In_688,In_687);
nor U69 (N_69,In_405,In_195);
and U70 (N_70,In_724,In_711);
nor U71 (N_71,In_348,In_301);
and U72 (N_72,In_178,In_284);
or U73 (N_73,In_365,In_208);
nand U74 (N_74,In_676,In_295);
and U75 (N_75,In_523,In_102);
or U76 (N_76,In_239,In_392);
nand U77 (N_77,In_7,In_28);
or U78 (N_78,In_501,In_223);
nor U79 (N_79,In_700,In_730);
nand U80 (N_80,In_213,In_74);
nor U81 (N_81,In_329,In_147);
and U82 (N_82,In_60,In_369);
and U83 (N_83,In_617,In_331);
nand U84 (N_84,In_101,In_651);
and U85 (N_85,In_633,In_698);
or U86 (N_86,In_739,In_601);
and U87 (N_87,In_266,In_443);
nor U88 (N_88,In_660,In_43);
or U89 (N_89,In_47,In_146);
or U90 (N_90,In_193,In_535);
nand U91 (N_91,In_509,In_299);
or U92 (N_92,In_669,In_82);
xor U93 (N_93,In_434,In_531);
nor U94 (N_94,In_554,In_455);
nand U95 (N_95,In_196,In_575);
and U96 (N_96,In_8,In_81);
and U97 (N_97,In_73,In_702);
and U98 (N_98,In_136,In_474);
and U99 (N_99,In_552,In_561);
and U100 (N_100,In_118,In_749);
or U101 (N_101,In_94,In_720);
nand U102 (N_102,In_694,In_431);
nand U103 (N_103,In_114,In_637);
and U104 (N_104,In_384,In_3);
and U105 (N_105,In_335,In_602);
and U106 (N_106,In_334,In_404);
or U107 (N_107,In_159,In_650);
or U108 (N_108,In_154,In_11);
nand U109 (N_109,In_222,In_35);
or U110 (N_110,In_12,In_486);
or U111 (N_111,In_636,In_565);
nand U112 (N_112,In_453,In_665);
nor U113 (N_113,In_173,In_576);
or U114 (N_114,In_72,In_233);
and U115 (N_115,In_417,In_220);
xnor U116 (N_116,In_206,In_247);
and U117 (N_117,In_706,In_260);
nand U118 (N_118,In_87,In_95);
and U119 (N_119,In_559,In_342);
or U120 (N_120,In_358,In_729);
and U121 (N_121,In_667,In_723);
and U122 (N_122,In_176,In_591);
or U123 (N_123,In_613,In_507);
nor U124 (N_124,In_380,In_619);
nor U125 (N_125,In_25,In_180);
or U126 (N_126,In_628,In_282);
or U127 (N_127,In_75,In_423);
nor U128 (N_128,In_29,In_320);
nand U129 (N_129,In_418,In_179);
nor U130 (N_130,In_252,In_255);
nor U131 (N_131,In_263,In_373);
nor U132 (N_132,In_630,In_366);
nand U133 (N_133,In_106,In_124);
and U134 (N_134,In_177,In_141);
or U135 (N_135,In_1,In_110);
nor U136 (N_136,In_524,In_545);
xnor U137 (N_137,In_683,In_530);
or U138 (N_138,In_495,In_360);
and U139 (N_139,In_42,In_409);
and U140 (N_140,In_302,In_484);
nand U141 (N_141,In_50,In_746);
nor U142 (N_142,In_14,In_675);
nand U143 (N_143,In_657,In_697);
xnor U144 (N_144,In_465,In_257);
and U145 (N_145,In_740,In_448);
nor U146 (N_146,In_696,In_132);
nand U147 (N_147,In_292,In_385);
nor U148 (N_148,In_375,In_133);
nand U149 (N_149,In_214,In_387);
nand U150 (N_150,In_528,In_416);
nor U151 (N_151,In_626,In_376);
xnor U152 (N_152,In_218,In_280);
nor U153 (N_153,In_227,In_459);
nor U154 (N_154,In_422,In_69);
and U155 (N_155,In_45,In_476);
or U156 (N_156,In_322,In_39);
or U157 (N_157,In_661,In_210);
nand U158 (N_158,In_30,In_152);
nor U159 (N_159,In_347,In_605);
nand U160 (N_160,In_703,In_427);
or U161 (N_161,In_122,In_745);
nand U162 (N_162,In_469,In_231);
or U163 (N_163,In_438,In_580);
xnor U164 (N_164,In_21,In_415);
nor U165 (N_165,In_105,In_67);
nand U166 (N_166,In_100,In_389);
nor U167 (N_167,In_468,In_182);
or U168 (N_168,In_491,In_615);
nor U169 (N_169,In_131,In_444);
xnor U170 (N_170,In_253,In_645);
nand U171 (N_171,In_648,In_421);
nand U172 (N_172,In_116,In_340);
or U173 (N_173,In_211,In_719);
nand U174 (N_174,In_692,In_411);
nor U175 (N_175,In_442,In_609);
or U176 (N_176,In_432,In_204);
nor U177 (N_177,In_516,In_640);
nand U178 (N_178,In_151,In_625);
nor U179 (N_179,In_49,In_471);
or U180 (N_180,In_643,In_175);
nor U181 (N_181,In_108,In_510);
nor U182 (N_182,In_117,In_272);
nor U183 (N_183,In_271,In_623);
nor U184 (N_184,In_107,In_364);
nand U185 (N_185,In_502,In_449);
nand U186 (N_186,In_89,In_611);
xnor U187 (N_187,In_500,In_44);
or U188 (N_188,In_357,In_424);
and U189 (N_189,In_76,In_85);
and U190 (N_190,In_649,In_515);
and U191 (N_191,In_462,In_96);
or U192 (N_192,In_287,In_78);
and U193 (N_193,In_62,In_201);
nor U194 (N_194,In_316,In_546);
and U195 (N_195,In_543,In_343);
nor U196 (N_196,In_205,In_184);
nand U197 (N_197,In_341,In_544);
nand U198 (N_198,In_337,In_269);
and U199 (N_199,In_412,In_560);
and U200 (N_200,In_0,In_721);
and U201 (N_201,In_450,In_597);
or U202 (N_202,In_202,In_203);
and U203 (N_203,In_396,In_377);
and U204 (N_204,In_307,In_65);
and U205 (N_205,In_519,In_398);
and U206 (N_206,In_192,In_354);
or U207 (N_207,In_603,In_310);
nand U208 (N_208,In_542,In_306);
or U209 (N_209,In_655,In_112);
nor U210 (N_210,In_514,In_103);
nand U211 (N_211,In_156,In_440);
nor U212 (N_212,In_234,In_186);
nand U213 (N_213,In_92,In_534);
and U214 (N_214,In_485,In_63);
or U215 (N_215,In_18,In_460);
nand U216 (N_216,In_228,In_200);
or U217 (N_217,In_317,In_526);
or U218 (N_218,In_494,In_170);
nand U219 (N_219,In_428,In_441);
or U220 (N_220,In_386,In_267);
nor U221 (N_221,In_672,In_699);
and U222 (N_222,In_172,In_232);
and U223 (N_223,In_437,In_243);
nor U224 (N_224,In_547,In_726);
and U225 (N_225,In_158,In_511);
and U226 (N_226,In_496,In_249);
nand U227 (N_227,In_250,In_506);
and U228 (N_228,In_240,In_32);
or U229 (N_229,In_285,In_315);
nor U230 (N_230,In_382,In_53);
or U231 (N_231,In_685,In_673);
or U232 (N_232,In_283,In_288);
nor U233 (N_233,In_658,In_664);
and U234 (N_234,In_262,In_695);
or U235 (N_235,In_482,In_743);
or U236 (N_236,In_209,In_610);
or U237 (N_237,In_84,In_614);
nand U238 (N_238,In_704,In_548);
nand U239 (N_239,In_479,In_127);
nand U240 (N_240,In_634,In_27);
nor U241 (N_241,In_349,In_97);
or U242 (N_242,In_568,In_451);
nor U243 (N_243,In_150,In_10);
or U244 (N_244,In_55,In_86);
xnor U245 (N_245,In_518,In_275);
or U246 (N_246,In_226,In_115);
or U247 (N_247,In_139,In_109);
or U248 (N_248,In_160,In_594);
and U249 (N_249,In_276,In_480);
nand U250 (N_250,In_140,In_338);
or U251 (N_251,In_571,In_701);
nand U252 (N_252,In_722,In_171);
and U253 (N_253,In_588,In_46);
and U254 (N_254,In_463,In_356);
nand U255 (N_255,In_339,In_52);
nor U256 (N_256,In_346,In_80);
nand U257 (N_257,In_273,In_646);
nand U258 (N_258,In_549,In_83);
nand U259 (N_259,In_142,In_281);
or U260 (N_260,In_167,In_584);
or U261 (N_261,In_642,In_90);
or U262 (N_262,In_587,In_627);
or U263 (N_263,In_128,In_23);
nor U264 (N_264,In_407,In_189);
nor U265 (N_265,In_6,In_153);
and U266 (N_266,In_569,In_216);
or U267 (N_267,In_174,In_572);
nor U268 (N_268,In_155,In_57);
xor U269 (N_269,In_56,In_363);
nand U270 (N_270,In_19,In_61);
and U271 (N_271,In_188,In_488);
nand U272 (N_272,In_583,In_466);
nor U273 (N_273,In_54,In_705);
or U274 (N_274,In_313,In_742);
nand U275 (N_275,In_458,In_235);
and U276 (N_276,In_682,In_647);
nand U277 (N_277,In_51,In_344);
nand U278 (N_278,In_718,In_577);
nor U279 (N_279,In_581,In_727);
and U280 (N_280,In_277,In_419);
nand U281 (N_281,In_300,In_536);
and U282 (N_282,In_37,In_558);
or U283 (N_283,In_731,In_563);
nand U284 (N_284,In_308,In_570);
and U285 (N_285,In_653,In_540);
or U286 (N_286,In_732,In_454);
nor U287 (N_287,In_606,In_345);
nand U288 (N_288,In_268,In_553);
or U289 (N_289,In_291,In_289);
and U290 (N_290,In_681,In_79);
nor U291 (N_291,In_183,In_734);
nand U292 (N_292,In_573,In_248);
or U293 (N_293,In_381,In_521);
or U294 (N_294,In_391,In_566);
nand U295 (N_295,In_677,In_641);
nor U296 (N_296,In_24,In_129);
and U297 (N_297,In_426,In_390);
nor U298 (N_298,In_351,In_595);
and U299 (N_299,In_36,In_728);
nand U300 (N_300,In_490,In_420);
nor U301 (N_301,In_618,In_632);
or U302 (N_302,In_325,In_66);
and U303 (N_303,In_379,In_71);
nand U304 (N_304,In_533,In_425);
and U305 (N_305,In_725,In_604);
nand U306 (N_306,In_684,In_400);
and U307 (N_307,In_564,In_656);
or U308 (N_308,In_219,In_508);
nor U309 (N_309,In_707,In_406);
nand U310 (N_310,In_362,In_589);
or U311 (N_311,In_217,In_199);
and U312 (N_312,In_654,In_666);
and U313 (N_313,In_40,In_330);
nor U314 (N_314,In_88,In_246);
nand U315 (N_315,In_163,In_2);
nor U316 (N_316,In_567,In_371);
and U317 (N_317,In_98,In_712);
nand U318 (N_318,In_207,In_492);
and U319 (N_319,In_555,In_639);
nand U320 (N_320,In_149,In_245);
nand U321 (N_321,In_113,In_397);
and U322 (N_322,In_370,In_467);
nand U323 (N_323,In_541,In_130);
nand U324 (N_324,In_312,In_13);
and U325 (N_325,In_148,In_693);
nand U326 (N_326,In_401,In_187);
or U327 (N_327,In_311,In_120);
and U328 (N_328,In_190,In_256);
or U329 (N_329,In_137,In_470);
nor U330 (N_330,In_265,In_520);
nor U331 (N_331,In_70,In_238);
nand U332 (N_332,In_690,In_747);
and U333 (N_333,In_261,In_557);
and U334 (N_334,In_9,In_395);
nor U335 (N_335,In_600,In_286);
nor U336 (N_336,In_77,In_323);
nand U337 (N_337,In_585,In_319);
nor U338 (N_338,In_305,In_607);
nand U339 (N_339,In_251,In_274);
nand U340 (N_340,In_34,In_22);
or U341 (N_341,In_41,In_483);
and U342 (N_342,In_652,In_328);
nor U343 (N_343,In_194,In_169);
and U344 (N_344,In_314,In_294);
or U345 (N_345,In_303,In_215);
nand U346 (N_346,In_663,In_119);
nand U347 (N_347,In_498,In_714);
nand U348 (N_348,In_430,In_616);
nor U349 (N_349,In_517,In_550);
nand U350 (N_350,In_33,In_350);
nand U351 (N_351,In_622,In_679);
and U352 (N_352,In_599,In_429);
and U353 (N_353,In_270,In_710);
nor U354 (N_354,In_744,In_318);
nand U355 (N_355,In_499,In_638);
nand U356 (N_356,In_489,In_121);
and U357 (N_357,In_433,In_478);
nand U358 (N_358,In_689,In_562);
and U359 (N_359,In_5,In_166);
or U360 (N_360,In_162,In_91);
nand U361 (N_361,In_388,In_629);
or U362 (N_362,In_436,In_229);
and U363 (N_363,In_487,In_403);
nand U364 (N_364,In_135,In_374);
and U365 (N_365,In_668,In_383);
or U366 (N_366,In_297,In_353);
nor U367 (N_367,In_736,In_537);
nand U368 (N_368,In_68,In_464);
nand U369 (N_369,In_527,In_593);
nand U370 (N_370,In_161,In_278);
nand U371 (N_371,In_529,In_145);
or U372 (N_372,In_111,In_659);
nand U373 (N_373,In_237,In_327);
nor U374 (N_374,In_104,In_399);
nand U375 (N_375,In_704,In_458);
or U376 (N_376,In_9,In_221);
nor U377 (N_377,In_452,In_411);
nand U378 (N_378,In_472,In_327);
nand U379 (N_379,In_363,In_577);
nor U380 (N_380,In_363,In_657);
or U381 (N_381,In_638,In_319);
nor U382 (N_382,In_75,In_133);
or U383 (N_383,In_337,In_264);
nand U384 (N_384,In_122,In_364);
and U385 (N_385,In_70,In_504);
nor U386 (N_386,In_145,In_17);
and U387 (N_387,In_578,In_400);
nand U388 (N_388,In_456,In_567);
nor U389 (N_389,In_334,In_448);
nor U390 (N_390,In_472,In_162);
and U391 (N_391,In_21,In_87);
or U392 (N_392,In_650,In_589);
or U393 (N_393,In_329,In_67);
or U394 (N_394,In_707,In_455);
nand U395 (N_395,In_56,In_545);
and U396 (N_396,In_7,In_474);
xor U397 (N_397,In_391,In_370);
or U398 (N_398,In_195,In_323);
or U399 (N_399,In_657,In_84);
or U400 (N_400,In_105,In_14);
and U401 (N_401,In_632,In_82);
and U402 (N_402,In_369,In_301);
nor U403 (N_403,In_505,In_143);
and U404 (N_404,In_597,In_686);
nor U405 (N_405,In_318,In_242);
nand U406 (N_406,In_466,In_217);
or U407 (N_407,In_734,In_258);
or U408 (N_408,In_530,In_658);
or U409 (N_409,In_527,In_322);
nand U410 (N_410,In_291,In_692);
xor U411 (N_411,In_447,In_183);
and U412 (N_412,In_166,In_384);
nor U413 (N_413,In_318,In_262);
or U414 (N_414,In_527,In_96);
nor U415 (N_415,In_170,In_729);
and U416 (N_416,In_124,In_263);
or U417 (N_417,In_242,In_126);
and U418 (N_418,In_101,In_578);
nand U419 (N_419,In_511,In_118);
or U420 (N_420,In_246,In_114);
nand U421 (N_421,In_51,In_616);
or U422 (N_422,In_291,In_101);
xor U423 (N_423,In_358,In_102);
and U424 (N_424,In_57,In_84);
or U425 (N_425,In_651,In_693);
nand U426 (N_426,In_747,In_301);
nand U427 (N_427,In_457,In_436);
and U428 (N_428,In_480,In_622);
and U429 (N_429,In_518,In_662);
nand U430 (N_430,In_170,In_85);
nor U431 (N_431,In_5,In_263);
or U432 (N_432,In_533,In_446);
nand U433 (N_433,In_169,In_702);
nor U434 (N_434,In_360,In_179);
or U435 (N_435,In_189,In_253);
or U436 (N_436,In_375,In_724);
nand U437 (N_437,In_577,In_230);
nor U438 (N_438,In_461,In_127);
or U439 (N_439,In_508,In_53);
and U440 (N_440,In_431,In_19);
or U441 (N_441,In_194,In_183);
or U442 (N_442,In_119,In_360);
nor U443 (N_443,In_17,In_637);
nand U444 (N_444,In_727,In_259);
and U445 (N_445,In_602,In_255);
and U446 (N_446,In_523,In_450);
nand U447 (N_447,In_693,In_448);
nand U448 (N_448,In_489,In_668);
and U449 (N_449,In_117,In_450);
nand U450 (N_450,In_563,In_595);
and U451 (N_451,In_146,In_607);
or U452 (N_452,In_46,In_164);
and U453 (N_453,In_567,In_513);
nand U454 (N_454,In_246,In_397);
nor U455 (N_455,In_234,In_166);
or U456 (N_456,In_204,In_469);
nand U457 (N_457,In_7,In_307);
nand U458 (N_458,In_417,In_721);
and U459 (N_459,In_313,In_221);
and U460 (N_460,In_25,In_583);
or U461 (N_461,In_685,In_387);
xor U462 (N_462,In_252,In_244);
and U463 (N_463,In_539,In_191);
or U464 (N_464,In_16,In_688);
nor U465 (N_465,In_389,In_500);
and U466 (N_466,In_171,In_343);
nor U467 (N_467,In_521,In_361);
or U468 (N_468,In_203,In_527);
nand U469 (N_469,In_525,In_56);
or U470 (N_470,In_441,In_3);
nand U471 (N_471,In_301,In_182);
or U472 (N_472,In_678,In_471);
or U473 (N_473,In_599,In_97);
nor U474 (N_474,In_625,In_476);
and U475 (N_475,In_23,In_252);
nand U476 (N_476,In_21,In_207);
nand U477 (N_477,In_611,In_9);
or U478 (N_478,In_548,In_442);
nor U479 (N_479,In_485,In_744);
nand U480 (N_480,In_257,In_365);
or U481 (N_481,In_38,In_629);
and U482 (N_482,In_333,In_176);
or U483 (N_483,In_420,In_318);
and U484 (N_484,In_323,In_389);
and U485 (N_485,In_650,In_248);
nor U486 (N_486,In_0,In_407);
and U487 (N_487,In_523,In_484);
nand U488 (N_488,In_566,In_563);
and U489 (N_489,In_578,In_735);
or U490 (N_490,In_309,In_640);
and U491 (N_491,In_30,In_185);
and U492 (N_492,In_495,In_6);
and U493 (N_493,In_241,In_567);
nor U494 (N_494,In_279,In_389);
nand U495 (N_495,In_263,In_142);
nand U496 (N_496,In_55,In_252);
nand U497 (N_497,In_212,In_612);
and U498 (N_498,In_321,In_421);
nor U499 (N_499,In_666,In_690);
or U500 (N_500,In_520,In_416);
nand U501 (N_501,In_404,In_462);
nand U502 (N_502,In_397,In_611);
and U503 (N_503,In_355,In_538);
nand U504 (N_504,In_242,In_608);
nand U505 (N_505,In_609,In_337);
and U506 (N_506,In_681,In_564);
nand U507 (N_507,In_610,In_150);
nor U508 (N_508,In_91,In_134);
nor U509 (N_509,In_570,In_255);
and U510 (N_510,In_577,In_426);
nand U511 (N_511,In_402,In_526);
or U512 (N_512,In_676,In_383);
nor U513 (N_513,In_165,In_724);
nand U514 (N_514,In_657,In_99);
and U515 (N_515,In_41,In_417);
nand U516 (N_516,In_428,In_543);
nand U517 (N_517,In_718,In_477);
and U518 (N_518,In_540,In_343);
nor U519 (N_519,In_189,In_435);
or U520 (N_520,In_539,In_271);
xor U521 (N_521,In_348,In_519);
or U522 (N_522,In_195,In_283);
xor U523 (N_523,In_348,In_533);
or U524 (N_524,In_580,In_345);
and U525 (N_525,In_476,In_269);
nor U526 (N_526,In_431,In_311);
xnor U527 (N_527,In_350,In_560);
nor U528 (N_528,In_175,In_664);
or U529 (N_529,In_300,In_297);
or U530 (N_530,In_104,In_448);
or U531 (N_531,In_685,In_674);
nor U532 (N_532,In_527,In_328);
nand U533 (N_533,In_457,In_674);
or U534 (N_534,In_639,In_482);
and U535 (N_535,In_706,In_514);
nor U536 (N_536,In_378,In_227);
nand U537 (N_537,In_560,In_276);
nor U538 (N_538,In_156,In_97);
nand U539 (N_539,In_313,In_553);
or U540 (N_540,In_667,In_205);
or U541 (N_541,In_304,In_602);
nand U542 (N_542,In_303,In_172);
and U543 (N_543,In_161,In_395);
or U544 (N_544,In_188,In_438);
nand U545 (N_545,In_469,In_39);
and U546 (N_546,In_734,In_571);
nor U547 (N_547,In_231,In_433);
nor U548 (N_548,In_151,In_114);
nand U549 (N_549,In_542,In_324);
nor U550 (N_550,In_135,In_262);
and U551 (N_551,In_681,In_554);
nand U552 (N_552,In_735,In_409);
or U553 (N_553,In_406,In_189);
nor U554 (N_554,In_451,In_418);
and U555 (N_555,In_0,In_102);
or U556 (N_556,In_94,In_269);
or U557 (N_557,In_672,In_666);
and U558 (N_558,In_513,In_598);
and U559 (N_559,In_316,In_715);
nor U560 (N_560,In_93,In_249);
nand U561 (N_561,In_241,In_70);
nand U562 (N_562,In_77,In_125);
nand U563 (N_563,In_21,In_105);
nor U564 (N_564,In_211,In_734);
or U565 (N_565,In_439,In_280);
and U566 (N_566,In_38,In_603);
or U567 (N_567,In_721,In_470);
and U568 (N_568,In_494,In_675);
or U569 (N_569,In_525,In_41);
or U570 (N_570,In_115,In_536);
nand U571 (N_571,In_727,In_70);
nand U572 (N_572,In_427,In_21);
and U573 (N_573,In_521,In_581);
or U574 (N_574,In_259,In_66);
or U575 (N_575,In_62,In_174);
nand U576 (N_576,In_536,In_26);
nand U577 (N_577,In_148,In_19);
xnor U578 (N_578,In_36,In_655);
nor U579 (N_579,In_710,In_201);
nand U580 (N_580,In_218,In_100);
or U581 (N_581,In_394,In_678);
or U582 (N_582,In_44,In_160);
and U583 (N_583,In_225,In_19);
or U584 (N_584,In_348,In_312);
nand U585 (N_585,In_730,In_502);
nand U586 (N_586,In_490,In_146);
nor U587 (N_587,In_34,In_594);
nand U588 (N_588,In_11,In_500);
or U589 (N_589,In_229,In_443);
or U590 (N_590,In_727,In_21);
xor U591 (N_591,In_290,In_458);
nor U592 (N_592,In_161,In_121);
nor U593 (N_593,In_632,In_479);
and U594 (N_594,In_73,In_625);
nor U595 (N_595,In_553,In_300);
nand U596 (N_596,In_448,In_717);
and U597 (N_597,In_136,In_643);
and U598 (N_598,In_44,In_116);
nand U599 (N_599,In_525,In_126);
xnor U600 (N_600,In_305,In_292);
or U601 (N_601,In_277,In_395);
or U602 (N_602,In_212,In_124);
nand U603 (N_603,In_409,In_236);
nand U604 (N_604,In_650,In_580);
or U605 (N_605,In_38,In_102);
or U606 (N_606,In_61,In_239);
nand U607 (N_607,In_374,In_651);
nand U608 (N_608,In_288,In_30);
nand U609 (N_609,In_644,In_201);
and U610 (N_610,In_649,In_467);
or U611 (N_611,In_614,In_749);
and U612 (N_612,In_196,In_619);
nor U613 (N_613,In_164,In_227);
and U614 (N_614,In_405,In_39);
nor U615 (N_615,In_470,In_688);
or U616 (N_616,In_160,In_434);
and U617 (N_617,In_58,In_247);
nand U618 (N_618,In_574,In_336);
nor U619 (N_619,In_531,In_356);
or U620 (N_620,In_644,In_330);
and U621 (N_621,In_12,In_11);
and U622 (N_622,In_613,In_544);
nor U623 (N_623,In_336,In_174);
and U624 (N_624,In_558,In_483);
or U625 (N_625,In_408,In_371);
nand U626 (N_626,In_734,In_326);
nand U627 (N_627,In_173,In_68);
nor U628 (N_628,In_454,In_299);
nor U629 (N_629,In_300,In_71);
nand U630 (N_630,In_303,In_179);
and U631 (N_631,In_151,In_233);
nor U632 (N_632,In_562,In_620);
or U633 (N_633,In_205,In_80);
nand U634 (N_634,In_90,In_253);
or U635 (N_635,In_215,In_223);
nor U636 (N_636,In_578,In_238);
nand U637 (N_637,In_133,In_486);
or U638 (N_638,In_300,In_33);
or U639 (N_639,In_680,In_725);
nor U640 (N_640,In_193,In_221);
nand U641 (N_641,In_144,In_515);
and U642 (N_642,In_409,In_722);
xnor U643 (N_643,In_682,In_475);
and U644 (N_644,In_416,In_740);
or U645 (N_645,In_232,In_577);
nor U646 (N_646,In_474,In_713);
and U647 (N_647,In_199,In_80);
and U648 (N_648,In_478,In_214);
or U649 (N_649,In_19,In_104);
and U650 (N_650,In_471,In_575);
nor U651 (N_651,In_115,In_220);
or U652 (N_652,In_660,In_485);
nand U653 (N_653,In_38,In_153);
xnor U654 (N_654,In_170,In_342);
nor U655 (N_655,In_678,In_40);
and U656 (N_656,In_76,In_165);
nor U657 (N_657,In_661,In_712);
or U658 (N_658,In_248,In_473);
nand U659 (N_659,In_346,In_16);
and U660 (N_660,In_27,In_406);
nand U661 (N_661,In_394,In_104);
nand U662 (N_662,In_178,In_660);
or U663 (N_663,In_153,In_276);
nand U664 (N_664,In_733,In_412);
nand U665 (N_665,In_173,In_353);
nor U666 (N_666,In_435,In_36);
nand U667 (N_667,In_716,In_365);
nand U668 (N_668,In_697,In_573);
nand U669 (N_669,In_503,In_172);
or U670 (N_670,In_730,In_325);
or U671 (N_671,In_172,In_731);
nor U672 (N_672,In_656,In_54);
or U673 (N_673,In_463,In_238);
or U674 (N_674,In_365,In_44);
nand U675 (N_675,In_245,In_197);
and U676 (N_676,In_292,In_454);
or U677 (N_677,In_407,In_115);
or U678 (N_678,In_119,In_282);
nand U679 (N_679,In_232,In_548);
and U680 (N_680,In_206,In_666);
or U681 (N_681,In_734,In_46);
and U682 (N_682,In_600,In_503);
and U683 (N_683,In_481,In_735);
or U684 (N_684,In_399,In_89);
nand U685 (N_685,In_521,In_309);
nor U686 (N_686,In_201,In_32);
or U687 (N_687,In_217,In_557);
nand U688 (N_688,In_316,In_161);
and U689 (N_689,In_212,In_239);
or U690 (N_690,In_566,In_389);
nand U691 (N_691,In_540,In_672);
xnor U692 (N_692,In_638,In_250);
nor U693 (N_693,In_209,In_656);
or U694 (N_694,In_562,In_121);
or U695 (N_695,In_516,In_509);
nand U696 (N_696,In_139,In_12);
nand U697 (N_697,In_719,In_218);
nor U698 (N_698,In_562,In_589);
and U699 (N_699,In_598,In_580);
nor U700 (N_700,In_550,In_399);
or U701 (N_701,In_446,In_514);
nand U702 (N_702,In_255,In_334);
and U703 (N_703,In_698,In_449);
nor U704 (N_704,In_57,In_608);
nand U705 (N_705,In_546,In_85);
and U706 (N_706,In_185,In_546);
or U707 (N_707,In_123,In_451);
or U708 (N_708,In_331,In_77);
nand U709 (N_709,In_201,In_571);
xor U710 (N_710,In_491,In_204);
nand U711 (N_711,In_623,In_490);
nand U712 (N_712,In_563,In_592);
nor U713 (N_713,In_460,In_657);
nor U714 (N_714,In_216,In_604);
nor U715 (N_715,In_151,In_562);
nand U716 (N_716,In_469,In_493);
or U717 (N_717,In_693,In_325);
or U718 (N_718,In_31,In_501);
nand U719 (N_719,In_509,In_657);
and U720 (N_720,In_97,In_337);
nor U721 (N_721,In_159,In_674);
nor U722 (N_722,In_481,In_471);
and U723 (N_723,In_582,In_150);
nand U724 (N_724,In_120,In_77);
and U725 (N_725,In_662,In_246);
or U726 (N_726,In_449,In_451);
or U727 (N_727,In_626,In_639);
or U728 (N_728,In_572,In_554);
nand U729 (N_729,In_611,In_483);
and U730 (N_730,In_69,In_626);
nand U731 (N_731,In_593,In_328);
and U732 (N_732,In_638,In_423);
nand U733 (N_733,In_239,In_102);
nor U734 (N_734,In_149,In_381);
or U735 (N_735,In_385,In_216);
and U736 (N_736,In_138,In_695);
and U737 (N_737,In_443,In_391);
nor U738 (N_738,In_101,In_514);
and U739 (N_739,In_311,In_603);
nand U740 (N_740,In_714,In_167);
nor U741 (N_741,In_435,In_310);
or U742 (N_742,In_18,In_40);
and U743 (N_743,In_296,In_531);
and U744 (N_744,In_740,In_357);
xnor U745 (N_745,In_237,In_16);
or U746 (N_746,In_740,In_130);
nor U747 (N_747,In_58,In_167);
xor U748 (N_748,In_548,In_558);
nor U749 (N_749,In_656,In_510);
or U750 (N_750,In_651,In_703);
and U751 (N_751,In_256,In_147);
xnor U752 (N_752,In_37,In_469);
nand U753 (N_753,In_355,In_645);
and U754 (N_754,In_121,In_461);
and U755 (N_755,In_709,In_49);
or U756 (N_756,In_566,In_731);
nand U757 (N_757,In_589,In_598);
nand U758 (N_758,In_370,In_338);
nor U759 (N_759,In_735,In_560);
or U760 (N_760,In_118,In_190);
and U761 (N_761,In_610,In_372);
nor U762 (N_762,In_126,In_577);
or U763 (N_763,In_511,In_391);
nor U764 (N_764,In_618,In_271);
and U765 (N_765,In_190,In_739);
or U766 (N_766,In_127,In_198);
and U767 (N_767,In_118,In_415);
nand U768 (N_768,In_427,In_526);
nand U769 (N_769,In_235,In_640);
nand U770 (N_770,In_91,In_564);
nor U771 (N_771,In_240,In_569);
nand U772 (N_772,In_259,In_550);
and U773 (N_773,In_137,In_405);
nand U774 (N_774,In_333,In_530);
and U775 (N_775,In_343,In_15);
and U776 (N_776,In_670,In_377);
nor U777 (N_777,In_285,In_346);
or U778 (N_778,In_459,In_69);
or U779 (N_779,In_221,In_450);
nor U780 (N_780,In_210,In_165);
and U781 (N_781,In_425,In_267);
nor U782 (N_782,In_36,In_73);
nand U783 (N_783,In_124,In_285);
nand U784 (N_784,In_16,In_534);
nand U785 (N_785,In_712,In_204);
nor U786 (N_786,In_331,In_444);
or U787 (N_787,In_667,In_206);
nand U788 (N_788,In_240,In_344);
nor U789 (N_789,In_320,In_483);
or U790 (N_790,In_312,In_119);
and U791 (N_791,In_471,In_543);
or U792 (N_792,In_719,In_651);
nor U793 (N_793,In_390,In_498);
or U794 (N_794,In_64,In_27);
and U795 (N_795,In_320,In_712);
nand U796 (N_796,In_704,In_64);
nand U797 (N_797,In_583,In_390);
nand U798 (N_798,In_589,In_123);
nand U799 (N_799,In_453,In_134);
or U800 (N_800,In_504,In_695);
and U801 (N_801,In_336,In_213);
nor U802 (N_802,In_650,In_677);
and U803 (N_803,In_41,In_361);
or U804 (N_804,In_558,In_117);
nor U805 (N_805,In_231,In_660);
or U806 (N_806,In_641,In_486);
and U807 (N_807,In_137,In_599);
xor U808 (N_808,In_275,In_567);
or U809 (N_809,In_581,In_199);
or U810 (N_810,In_296,In_422);
nand U811 (N_811,In_75,In_582);
nand U812 (N_812,In_749,In_267);
nor U813 (N_813,In_237,In_532);
nand U814 (N_814,In_72,In_316);
nand U815 (N_815,In_445,In_494);
nand U816 (N_816,In_632,In_463);
xor U817 (N_817,In_310,In_561);
and U818 (N_818,In_671,In_192);
nand U819 (N_819,In_654,In_167);
and U820 (N_820,In_470,In_642);
nand U821 (N_821,In_105,In_82);
and U822 (N_822,In_520,In_448);
nor U823 (N_823,In_475,In_32);
and U824 (N_824,In_611,In_27);
nor U825 (N_825,In_672,In_370);
and U826 (N_826,In_422,In_341);
and U827 (N_827,In_166,In_642);
and U828 (N_828,In_53,In_155);
nand U829 (N_829,In_634,In_622);
nor U830 (N_830,In_440,In_331);
and U831 (N_831,In_341,In_723);
nor U832 (N_832,In_386,In_26);
xor U833 (N_833,In_516,In_694);
nand U834 (N_834,In_357,In_442);
and U835 (N_835,In_259,In_164);
nor U836 (N_836,In_663,In_487);
or U837 (N_837,In_547,In_392);
and U838 (N_838,In_313,In_619);
and U839 (N_839,In_636,In_231);
nor U840 (N_840,In_174,In_417);
nor U841 (N_841,In_349,In_459);
and U842 (N_842,In_517,In_126);
nor U843 (N_843,In_10,In_460);
and U844 (N_844,In_708,In_434);
nor U845 (N_845,In_249,In_404);
nor U846 (N_846,In_580,In_474);
nand U847 (N_847,In_483,In_112);
nand U848 (N_848,In_110,In_585);
nand U849 (N_849,In_12,In_334);
nand U850 (N_850,In_510,In_628);
nand U851 (N_851,In_632,In_357);
nor U852 (N_852,In_427,In_471);
nor U853 (N_853,In_333,In_126);
nor U854 (N_854,In_359,In_461);
or U855 (N_855,In_558,In_329);
and U856 (N_856,In_111,In_576);
or U857 (N_857,In_85,In_393);
and U858 (N_858,In_732,In_198);
nor U859 (N_859,In_459,In_542);
or U860 (N_860,In_128,In_50);
or U861 (N_861,In_729,In_471);
nand U862 (N_862,In_465,In_653);
or U863 (N_863,In_621,In_151);
xor U864 (N_864,In_157,In_309);
nand U865 (N_865,In_305,In_18);
nand U866 (N_866,In_108,In_710);
and U867 (N_867,In_368,In_0);
nand U868 (N_868,In_576,In_337);
nor U869 (N_869,In_82,In_165);
and U870 (N_870,In_586,In_549);
or U871 (N_871,In_4,In_501);
nand U872 (N_872,In_577,In_164);
xor U873 (N_873,In_655,In_718);
and U874 (N_874,In_509,In_385);
nor U875 (N_875,In_248,In_119);
nor U876 (N_876,In_151,In_248);
nor U877 (N_877,In_80,In_351);
nor U878 (N_878,In_254,In_26);
nand U879 (N_879,In_234,In_249);
and U880 (N_880,In_31,In_277);
and U881 (N_881,In_590,In_33);
nor U882 (N_882,In_506,In_46);
nand U883 (N_883,In_142,In_740);
or U884 (N_884,In_480,In_332);
or U885 (N_885,In_615,In_56);
or U886 (N_886,In_393,In_129);
nand U887 (N_887,In_345,In_492);
nor U888 (N_888,In_431,In_115);
or U889 (N_889,In_276,In_453);
nand U890 (N_890,In_482,In_613);
and U891 (N_891,In_733,In_600);
nand U892 (N_892,In_361,In_148);
nand U893 (N_893,In_707,In_712);
or U894 (N_894,In_531,In_602);
nor U895 (N_895,In_641,In_356);
nor U896 (N_896,In_379,In_386);
nor U897 (N_897,In_534,In_126);
or U898 (N_898,In_728,In_618);
or U899 (N_899,In_429,In_731);
and U900 (N_900,In_197,In_9);
and U901 (N_901,In_237,In_215);
or U902 (N_902,In_617,In_304);
nor U903 (N_903,In_61,In_244);
and U904 (N_904,In_289,In_503);
xnor U905 (N_905,In_120,In_573);
and U906 (N_906,In_290,In_219);
nand U907 (N_907,In_265,In_706);
xor U908 (N_908,In_514,In_541);
and U909 (N_909,In_467,In_322);
or U910 (N_910,In_121,In_99);
or U911 (N_911,In_6,In_438);
nor U912 (N_912,In_646,In_267);
and U913 (N_913,In_0,In_247);
nor U914 (N_914,In_195,In_362);
or U915 (N_915,In_210,In_331);
nand U916 (N_916,In_476,In_666);
and U917 (N_917,In_632,In_584);
nor U918 (N_918,In_232,In_468);
nor U919 (N_919,In_74,In_291);
nor U920 (N_920,In_580,In_170);
or U921 (N_921,In_746,In_159);
nor U922 (N_922,In_253,In_141);
and U923 (N_923,In_574,In_530);
and U924 (N_924,In_298,In_535);
nor U925 (N_925,In_746,In_169);
or U926 (N_926,In_404,In_264);
or U927 (N_927,In_221,In_499);
and U928 (N_928,In_550,In_192);
nor U929 (N_929,In_78,In_711);
or U930 (N_930,In_37,In_506);
nor U931 (N_931,In_23,In_62);
nand U932 (N_932,In_194,In_200);
nor U933 (N_933,In_663,In_651);
nor U934 (N_934,In_93,In_241);
nand U935 (N_935,In_738,In_508);
nand U936 (N_936,In_252,In_4);
nand U937 (N_937,In_612,In_670);
nor U938 (N_938,In_453,In_232);
nand U939 (N_939,In_51,In_229);
xor U940 (N_940,In_623,In_202);
or U941 (N_941,In_351,In_219);
nand U942 (N_942,In_35,In_296);
and U943 (N_943,In_327,In_199);
nor U944 (N_944,In_420,In_737);
or U945 (N_945,In_570,In_395);
or U946 (N_946,In_592,In_139);
or U947 (N_947,In_449,In_26);
nand U948 (N_948,In_178,In_203);
nand U949 (N_949,In_631,In_409);
or U950 (N_950,In_500,In_468);
or U951 (N_951,In_31,In_226);
and U952 (N_952,In_695,In_301);
or U953 (N_953,In_547,In_627);
and U954 (N_954,In_202,In_12);
nor U955 (N_955,In_401,In_517);
nor U956 (N_956,In_224,In_72);
nand U957 (N_957,In_75,In_320);
nor U958 (N_958,In_440,In_233);
and U959 (N_959,In_348,In_37);
nor U960 (N_960,In_131,In_467);
nand U961 (N_961,In_302,In_191);
or U962 (N_962,In_410,In_476);
or U963 (N_963,In_626,In_135);
or U964 (N_964,In_376,In_360);
and U965 (N_965,In_59,In_77);
nor U966 (N_966,In_84,In_93);
and U967 (N_967,In_572,In_350);
nor U968 (N_968,In_111,In_498);
and U969 (N_969,In_284,In_161);
nor U970 (N_970,In_360,In_192);
and U971 (N_971,In_727,In_689);
nor U972 (N_972,In_560,In_501);
nor U973 (N_973,In_577,In_593);
nor U974 (N_974,In_157,In_46);
or U975 (N_975,In_392,In_47);
nand U976 (N_976,In_181,In_76);
and U977 (N_977,In_47,In_307);
or U978 (N_978,In_88,In_318);
nand U979 (N_979,In_200,In_119);
nand U980 (N_980,In_600,In_75);
nor U981 (N_981,In_376,In_443);
nor U982 (N_982,In_6,In_149);
nand U983 (N_983,In_519,In_37);
nand U984 (N_984,In_13,In_181);
nand U985 (N_985,In_275,In_529);
or U986 (N_986,In_315,In_548);
nand U987 (N_987,In_261,In_677);
nor U988 (N_988,In_544,In_224);
or U989 (N_989,In_334,In_636);
and U990 (N_990,In_328,In_45);
nand U991 (N_991,In_455,In_265);
nor U992 (N_992,In_394,In_269);
nand U993 (N_993,In_274,In_397);
nor U994 (N_994,In_9,In_468);
nor U995 (N_995,In_216,In_266);
nand U996 (N_996,In_382,In_456);
and U997 (N_997,In_384,In_262);
nand U998 (N_998,In_595,In_362);
and U999 (N_999,In_264,In_600);
and U1000 (N_1000,N_92,N_863);
or U1001 (N_1001,N_500,N_20);
nor U1002 (N_1002,N_621,N_835);
nor U1003 (N_1003,N_821,N_507);
and U1004 (N_1004,N_772,N_257);
nand U1005 (N_1005,N_998,N_258);
or U1006 (N_1006,N_189,N_845);
and U1007 (N_1007,N_607,N_265);
nor U1008 (N_1008,N_634,N_545);
and U1009 (N_1009,N_372,N_771);
nor U1010 (N_1010,N_929,N_622);
nand U1011 (N_1011,N_698,N_39);
nand U1012 (N_1012,N_478,N_994);
nor U1013 (N_1013,N_702,N_591);
nor U1014 (N_1014,N_88,N_530);
nor U1015 (N_1015,N_350,N_367);
nor U1016 (N_1016,N_52,N_949);
nand U1017 (N_1017,N_346,N_36);
and U1018 (N_1018,N_947,N_932);
nand U1019 (N_1019,N_16,N_332);
nor U1020 (N_1020,N_142,N_260);
nor U1021 (N_1021,N_21,N_982);
xor U1022 (N_1022,N_983,N_865);
and U1023 (N_1023,N_503,N_517);
nor U1024 (N_1024,N_104,N_447);
nand U1025 (N_1025,N_944,N_559);
nor U1026 (N_1026,N_717,N_615);
nor U1027 (N_1027,N_709,N_53);
nand U1028 (N_1028,N_329,N_594);
and U1029 (N_1029,N_436,N_651);
nand U1030 (N_1030,N_358,N_619);
nor U1031 (N_1031,N_943,N_66);
nor U1032 (N_1032,N_483,N_223);
and U1033 (N_1033,N_776,N_746);
nor U1034 (N_1034,N_286,N_431);
nand U1035 (N_1035,N_301,N_552);
and U1036 (N_1036,N_800,N_527);
nand U1037 (N_1037,N_981,N_421);
and U1038 (N_1038,N_40,N_577);
and U1039 (N_1039,N_391,N_555);
nor U1040 (N_1040,N_720,N_61);
and U1041 (N_1041,N_830,N_909);
nor U1042 (N_1042,N_586,N_751);
and U1043 (N_1043,N_413,N_650);
and U1044 (N_1044,N_756,N_208);
nand U1045 (N_1045,N_222,N_65);
and U1046 (N_1046,N_846,N_637);
or U1047 (N_1047,N_311,N_597);
nand U1048 (N_1048,N_548,N_339);
nor U1049 (N_1049,N_729,N_697);
and U1050 (N_1050,N_567,N_907);
nand U1051 (N_1051,N_195,N_822);
and U1052 (N_1052,N_374,N_127);
nand U1053 (N_1053,N_658,N_46);
nor U1054 (N_1054,N_762,N_376);
nand U1055 (N_1055,N_921,N_331);
and U1056 (N_1056,N_737,N_216);
or U1057 (N_1057,N_590,N_246);
and U1058 (N_1058,N_533,N_394);
nand U1059 (N_1059,N_494,N_871);
or U1060 (N_1060,N_85,N_589);
nor U1061 (N_1061,N_428,N_707);
xnor U1062 (N_1062,N_814,N_480);
nor U1063 (N_1063,N_758,N_768);
nand U1064 (N_1064,N_973,N_370);
nor U1065 (N_1065,N_302,N_390);
and U1066 (N_1066,N_633,N_701);
nand U1067 (N_1067,N_528,N_749);
or U1068 (N_1068,N_491,N_81);
nor U1069 (N_1069,N_557,N_156);
and U1070 (N_1070,N_902,N_769);
and U1071 (N_1071,N_505,N_726);
or U1072 (N_1072,N_173,N_671);
nor U1073 (N_1073,N_809,N_453);
nand U1074 (N_1074,N_520,N_851);
or U1075 (N_1075,N_522,N_891);
nand U1076 (N_1076,N_963,N_734);
or U1077 (N_1077,N_477,N_427);
nor U1078 (N_1078,N_308,N_688);
and U1079 (N_1079,N_719,N_958);
nand U1080 (N_1080,N_618,N_5);
and U1081 (N_1081,N_109,N_630);
nand U1082 (N_1082,N_916,N_315);
nand U1083 (N_1083,N_914,N_504);
nor U1084 (N_1084,N_324,N_255);
and U1085 (N_1085,N_613,N_248);
nand U1086 (N_1086,N_244,N_291);
or U1087 (N_1087,N_554,N_123);
nand U1088 (N_1088,N_458,N_990);
and U1089 (N_1089,N_913,N_623);
or U1090 (N_1090,N_212,N_672);
nor U1091 (N_1091,N_918,N_653);
nand U1092 (N_1092,N_784,N_899);
xor U1093 (N_1093,N_97,N_514);
nand U1094 (N_1094,N_669,N_160);
and U1095 (N_1095,N_628,N_967);
and U1096 (N_1096,N_384,N_207);
nor U1097 (N_1097,N_885,N_22);
or U1098 (N_1098,N_654,N_64);
nor U1099 (N_1099,N_681,N_12);
nand U1100 (N_1100,N_241,N_873);
xnor U1101 (N_1101,N_656,N_802);
xnor U1102 (N_1102,N_215,N_985);
nor U1103 (N_1103,N_31,N_617);
or U1104 (N_1104,N_366,N_68);
or U1105 (N_1105,N_682,N_282);
or U1106 (N_1106,N_582,N_177);
nand U1107 (N_1107,N_323,N_632);
nand U1108 (N_1108,N_534,N_131);
xor U1109 (N_1109,N_778,N_338);
nand U1110 (N_1110,N_823,N_787);
or U1111 (N_1111,N_939,N_640);
nand U1112 (N_1112,N_472,N_72);
or U1113 (N_1113,N_855,N_462);
nand U1114 (N_1114,N_881,N_411);
nand U1115 (N_1115,N_111,N_306);
nor U1116 (N_1116,N_979,N_463);
nor U1117 (N_1117,N_767,N_174);
nand U1118 (N_1118,N_9,N_203);
nor U1119 (N_1119,N_788,N_412);
and U1120 (N_1120,N_580,N_889);
and U1121 (N_1121,N_437,N_735);
and U1122 (N_1122,N_704,N_793);
and U1123 (N_1123,N_354,N_231);
and U1124 (N_1124,N_599,N_867);
or U1125 (N_1125,N_280,N_598);
or U1126 (N_1126,N_502,N_202);
or U1127 (N_1127,N_908,N_397);
and U1128 (N_1128,N_410,N_158);
or U1129 (N_1129,N_403,N_449);
nand U1130 (N_1130,N_588,N_225);
or U1131 (N_1131,N_314,N_135);
and U1132 (N_1132,N_644,N_550);
and U1133 (N_1133,N_196,N_780);
or U1134 (N_1134,N_538,N_129);
xor U1135 (N_1135,N_581,N_17);
and U1136 (N_1136,N_529,N_100);
nand U1137 (N_1137,N_262,N_708);
nor U1138 (N_1138,N_307,N_465);
nor U1139 (N_1139,N_101,N_815);
or U1140 (N_1140,N_647,N_506);
nand U1141 (N_1141,N_816,N_853);
nand U1142 (N_1142,N_812,N_128);
and U1143 (N_1143,N_952,N_696);
or U1144 (N_1144,N_677,N_831);
and U1145 (N_1145,N_404,N_94);
or U1146 (N_1146,N_897,N_446);
or U1147 (N_1147,N_86,N_381);
nor U1148 (N_1148,N_44,N_89);
nand U1149 (N_1149,N_469,N_32);
or U1150 (N_1150,N_84,N_475);
or U1151 (N_1151,N_214,N_13);
and U1152 (N_1152,N_833,N_743);
nor U1153 (N_1153,N_95,N_6);
or U1154 (N_1154,N_674,N_261);
and U1155 (N_1155,N_245,N_182);
nor U1156 (N_1156,N_572,N_638);
nor U1157 (N_1157,N_206,N_344);
nand U1158 (N_1158,N_984,N_229);
and U1159 (N_1159,N_595,N_98);
nor U1160 (N_1160,N_243,N_515);
and U1161 (N_1161,N_728,N_551);
nor U1162 (N_1162,N_804,N_278);
and U1163 (N_1163,N_740,N_826);
nor U1164 (N_1164,N_711,N_612);
nor U1165 (N_1165,N_721,N_148);
nor U1166 (N_1166,N_976,N_763);
nand U1167 (N_1167,N_145,N_606);
or U1168 (N_1168,N_143,N_236);
or U1169 (N_1169,N_498,N_284);
and U1170 (N_1170,N_636,N_903);
and U1171 (N_1171,N_542,N_93);
and U1172 (N_1172,N_493,N_336);
nand U1173 (N_1173,N_247,N_103);
or U1174 (N_1174,N_836,N_620);
nor U1175 (N_1175,N_635,N_991);
and U1176 (N_1176,N_774,N_348);
and U1177 (N_1177,N_874,N_213);
nand U1178 (N_1178,N_825,N_353);
and U1179 (N_1179,N_604,N_923);
nand U1180 (N_1180,N_194,N_710);
and U1181 (N_1181,N_497,N_954);
or U1182 (N_1182,N_549,N_254);
and U1183 (N_1183,N_789,N_27);
or U1184 (N_1184,N_673,N_797);
nor U1185 (N_1185,N_333,N_11);
nor U1186 (N_1186,N_796,N_54);
nand U1187 (N_1187,N_288,N_912);
nand U1188 (N_1188,N_537,N_235);
and U1189 (N_1189,N_322,N_355);
or U1190 (N_1190,N_883,N_573);
nor U1191 (N_1191,N_226,N_425);
nand U1192 (N_1192,N_365,N_327);
nor U1193 (N_1193,N_553,N_523);
nand U1194 (N_1194,N_648,N_352);
nand U1195 (N_1195,N_794,N_840);
and U1196 (N_1196,N_175,N_924);
nand U1197 (N_1197,N_470,N_441);
nor U1198 (N_1198,N_155,N_316);
xor U1199 (N_1199,N_209,N_509);
or U1200 (N_1200,N_79,N_820);
and U1201 (N_1201,N_313,N_3);
nor U1202 (N_1202,N_201,N_844);
or U1203 (N_1203,N_576,N_592);
nor U1204 (N_1204,N_432,N_198);
nor U1205 (N_1205,N_655,N_218);
and U1206 (N_1206,N_420,N_753);
and U1207 (N_1207,N_687,N_884);
or U1208 (N_1208,N_583,N_666);
nand U1209 (N_1209,N_955,N_798);
nand U1210 (N_1210,N_188,N_661);
and U1211 (N_1211,N_747,N_965);
nor U1212 (N_1212,N_543,N_657);
or U1213 (N_1213,N_91,N_481);
and U1214 (N_1214,N_312,N_186);
and U1215 (N_1215,N_276,N_783);
nand U1216 (N_1216,N_665,N_745);
nand U1217 (N_1217,N_18,N_434);
and U1218 (N_1218,N_414,N_392);
nor U1219 (N_1219,N_678,N_748);
or U1220 (N_1220,N_304,N_340);
and U1221 (N_1221,N_948,N_561);
nor U1222 (N_1222,N_754,N_813);
nor U1223 (N_1223,N_96,N_806);
nor U1224 (N_1224,N_942,N_490);
and U1225 (N_1225,N_41,N_137);
nor U1226 (N_1226,N_405,N_319);
nand U1227 (N_1227,N_968,N_387);
nor U1228 (N_1228,N_759,N_832);
nand U1229 (N_1229,N_80,N_69);
and U1230 (N_1230,N_685,N_722);
nor U1231 (N_1231,N_872,N_87);
or U1232 (N_1232,N_879,N_880);
nor U1233 (N_1233,N_895,N_971);
or U1234 (N_1234,N_922,N_373);
or U1235 (N_1235,N_888,N_102);
or U1236 (N_1236,N_950,N_556);
nand U1237 (N_1237,N_118,N_133);
or U1238 (N_1238,N_0,N_703);
or U1239 (N_1239,N_83,N_892);
nand U1240 (N_1240,N_356,N_911);
or U1241 (N_1241,N_219,N_435);
nand U1242 (N_1242,N_113,N_742);
xor U1243 (N_1243,N_675,N_153);
nor U1244 (N_1244,N_574,N_807);
nor U1245 (N_1245,N_466,N_693);
nor U1246 (N_1246,N_151,N_105);
and U1247 (N_1247,N_570,N_519);
nor U1248 (N_1248,N_876,N_290);
and U1249 (N_1249,N_975,N_579);
nor U1250 (N_1250,N_139,N_303);
or U1251 (N_1251,N_608,N_627);
nor U1252 (N_1252,N_170,N_318);
nor U1253 (N_1253,N_532,N_668);
nor U1254 (N_1254,N_773,N_915);
nand U1255 (N_1255,N_90,N_724);
nand U1256 (N_1256,N_386,N_325);
nand U1257 (N_1257,N_361,N_988);
and U1258 (N_1258,N_77,N_117);
nand U1259 (N_1259,N_602,N_869);
or U1260 (N_1260,N_126,N_275);
nand U1261 (N_1261,N_38,N_416);
nand U1262 (N_1262,N_992,N_919);
nor U1263 (N_1263,N_974,N_70);
and U1264 (N_1264,N_250,N_192);
or U1265 (N_1265,N_646,N_839);
and U1266 (N_1266,N_183,N_861);
and U1267 (N_1267,N_824,N_781);
or U1268 (N_1268,N_566,N_680);
or U1269 (N_1269,N_964,N_371);
or U1270 (N_1270,N_442,N_264);
or U1271 (N_1271,N_289,N_179);
and U1272 (N_1272,N_692,N_396);
and U1273 (N_1273,N_266,N_970);
or U1274 (N_1274,N_766,N_341);
nand U1275 (N_1275,N_438,N_320);
or U1276 (N_1276,N_712,N_511);
and U1277 (N_1277,N_645,N_144);
nand U1278 (N_1278,N_540,N_140);
nand U1279 (N_1279,N_488,N_684);
nand U1280 (N_1280,N_642,N_120);
nor U1281 (N_1281,N_492,N_699);
nor U1282 (N_1282,N_864,N_736);
nand U1283 (N_1283,N_896,N_811);
nand U1284 (N_1284,N_852,N_829);
nand U1285 (N_1285,N_310,N_937);
or U1286 (N_1286,N_78,N_631);
or U1287 (N_1287,N_114,N_799);
or U1288 (N_1288,N_443,N_2);
and U1289 (N_1289,N_546,N_29);
nand U1290 (N_1290,N_14,N_169);
nand U1291 (N_1291,N_450,N_147);
and U1292 (N_1292,N_989,N_960);
or U1293 (N_1293,N_150,N_134);
nor U1294 (N_1294,N_689,N_228);
xor U1295 (N_1295,N_489,N_106);
nand U1296 (N_1296,N_934,N_945);
and U1297 (N_1297,N_525,N_191);
and U1298 (N_1298,N_733,N_168);
or U1299 (N_1299,N_526,N_249);
nor U1300 (N_1300,N_999,N_518);
nand U1301 (N_1301,N_269,N_558);
nor U1302 (N_1302,N_43,N_940);
or U1303 (N_1303,N_423,N_210);
or U1304 (N_1304,N_877,N_461);
or U1305 (N_1305,N_440,N_51);
xor U1306 (N_1306,N_380,N_157);
nand U1307 (N_1307,N_842,N_121);
or U1308 (N_1308,N_35,N_452);
and U1309 (N_1309,N_584,N_775);
nand U1310 (N_1310,N_957,N_565);
and U1311 (N_1311,N_904,N_292);
and U1312 (N_1312,N_395,N_345);
and U1313 (N_1313,N_920,N_433);
and U1314 (N_1314,N_227,N_281);
nor U1315 (N_1315,N_605,N_321);
or U1316 (N_1316,N_459,N_730);
nor U1317 (N_1317,N_424,N_232);
and U1318 (N_1318,N_828,N_136);
nand U1319 (N_1319,N_178,N_905);
xor U1320 (N_1320,N_870,N_299);
nor U1321 (N_1321,N_676,N_987);
and U1322 (N_1322,N_107,N_429);
and U1323 (N_1323,N_337,N_841);
and U1324 (N_1324,N_409,N_808);
nand U1325 (N_1325,N_818,N_856);
nor U1326 (N_1326,N_791,N_415);
nand U1327 (N_1327,N_935,N_455);
xnor U1328 (N_1328,N_242,N_159);
and U1329 (N_1329,N_277,N_110);
xor U1330 (N_1330,N_388,N_351);
xnor U1331 (N_1331,N_611,N_297);
and U1332 (N_1332,N_847,N_801);
and U1333 (N_1333,N_805,N_256);
nand U1334 (N_1334,N_162,N_850);
or U1335 (N_1335,N_473,N_263);
or U1336 (N_1336,N_167,N_639);
nand U1337 (N_1337,N_866,N_616);
and U1338 (N_1338,N_849,N_58);
nand U1339 (N_1339,N_237,N_460);
or U1340 (N_1340,N_283,N_330);
or U1341 (N_1341,N_760,N_230);
and U1342 (N_1342,N_995,N_487);
nor U1343 (N_1343,N_15,N_716);
and U1344 (N_1344,N_238,N_777);
and U1345 (N_1345,N_510,N_50);
or U1346 (N_1346,N_910,N_204);
and U1347 (N_1347,N_977,N_596);
and U1348 (N_1348,N_521,N_695);
nor U1349 (N_1349,N_539,N_670);
and U1350 (N_1350,N_211,N_393);
or U1351 (N_1351,N_71,N_193);
nand U1352 (N_1352,N_400,N_363);
nand U1353 (N_1353,N_936,N_184);
nand U1354 (N_1354,N_785,N_398);
nand U1355 (N_1355,N_927,N_7);
nand U1356 (N_1356,N_854,N_513);
and U1357 (N_1357,N_761,N_34);
nor U1358 (N_1358,N_385,N_270);
or U1359 (N_1359,N_690,N_482);
and U1360 (N_1360,N_399,N_585);
nor U1361 (N_1361,N_593,N_124);
and U1362 (N_1362,N_508,N_660);
nand U1363 (N_1363,N_713,N_300);
and U1364 (N_1364,N_499,N_770);
or U1365 (N_1365,N_817,N_408);
and U1366 (N_1366,N_418,N_221);
or U1367 (N_1367,N_24,N_878);
nor U1368 (N_1368,N_643,N_19);
or U1369 (N_1369,N_146,N_382);
or U1370 (N_1370,N_444,N_486);
or U1371 (N_1371,N_45,N_335);
and U1372 (N_1372,N_894,N_224);
or U1373 (N_1373,N_700,N_900);
nand U1374 (N_1374,N_587,N_63);
or U1375 (N_1375,N_326,N_547);
or U1376 (N_1376,N_739,N_417);
nand U1377 (N_1377,N_959,N_360);
and U1378 (N_1378,N_112,N_890);
xor U1379 (N_1379,N_457,N_317);
xnor U1380 (N_1380,N_217,N_8);
or U1381 (N_1381,N_838,N_233);
nand U1382 (N_1382,N_234,N_1);
nand U1383 (N_1383,N_401,N_171);
and U1384 (N_1384,N_686,N_328);
and U1385 (N_1385,N_536,N_73);
xnor U1386 (N_1386,N_859,N_33);
or U1387 (N_1387,N_10,N_60);
nor U1388 (N_1388,N_454,N_969);
or U1389 (N_1389,N_122,N_274);
nand U1390 (N_1390,N_744,N_205);
nand U1391 (N_1391,N_993,N_868);
and U1392 (N_1392,N_926,N_827);
nor U1393 (N_1393,N_138,N_164);
nand U1394 (N_1394,N_239,N_858);
or U1395 (N_1395,N_163,N_860);
or U1396 (N_1396,N_172,N_149);
or U1397 (N_1397,N_220,N_792);
nand U1398 (N_1398,N_706,N_402);
nand U1399 (N_1399,N_516,N_757);
and U1400 (N_1400,N_917,N_560);
nand U1401 (N_1401,N_715,N_629);
or U1402 (N_1402,N_26,N_512);
xor U1403 (N_1403,N_562,N_378);
and U1404 (N_1404,N_731,N_62);
nor U1405 (N_1405,N_293,N_887);
nor U1406 (N_1406,N_74,N_116);
nor U1407 (N_1407,N_285,N_349);
or U1408 (N_1408,N_82,N_803);
nand U1409 (N_1409,N_741,N_609);
nand U1410 (N_1410,N_875,N_426);
or U1411 (N_1411,N_125,N_28);
nor U1412 (N_1412,N_649,N_364);
and U1413 (N_1413,N_980,N_786);
or U1414 (N_1414,N_610,N_810);
nand U1415 (N_1415,N_819,N_928);
nand U1416 (N_1416,N_925,N_569);
nand U1417 (N_1417,N_42,N_564);
nand U1418 (N_1418,N_176,N_47);
and U1419 (N_1419,N_997,N_99);
and U1420 (N_1420,N_108,N_130);
nand U1421 (N_1421,N_119,N_750);
nor U1422 (N_1422,N_190,N_972);
and U1423 (N_1423,N_563,N_501);
nor U1424 (N_1424,N_898,N_343);
nand U1425 (N_1425,N_886,N_166);
nor U1426 (N_1426,N_342,N_25);
and U1427 (N_1427,N_603,N_451);
nor U1428 (N_1428,N_956,N_614);
xnor U1429 (N_1429,N_694,N_48);
nand U1430 (N_1430,N_966,N_765);
and U1431 (N_1431,N_931,N_795);
nor U1432 (N_1432,N_782,N_714);
and U1433 (N_1433,N_541,N_837);
nand U1434 (N_1434,N_625,N_368);
nand U1435 (N_1435,N_790,N_406);
or U1436 (N_1436,N_571,N_495);
nand U1437 (N_1437,N_601,N_251);
nor U1438 (N_1438,N_377,N_132);
nand U1439 (N_1439,N_524,N_305);
and U1440 (N_1440,N_755,N_468);
and U1441 (N_1441,N_334,N_893);
and U1442 (N_1442,N_389,N_165);
nand U1443 (N_1443,N_115,N_941);
nor U1444 (N_1444,N_930,N_986);
nand U1445 (N_1445,N_496,N_294);
nor U1446 (N_1446,N_267,N_309);
or U1447 (N_1447,N_843,N_578);
or U1448 (N_1448,N_4,N_271);
nor U1449 (N_1449,N_185,N_359);
or U1450 (N_1450,N_422,N_199);
nor U1451 (N_1451,N_933,N_723);
nor U1452 (N_1452,N_448,N_725);
nand U1453 (N_1453,N_600,N_152);
nand U1454 (N_1454,N_764,N_407);
nand U1455 (N_1455,N_383,N_779);
and U1456 (N_1456,N_23,N_961);
nor U1457 (N_1457,N_296,N_272);
xnor U1458 (N_1458,N_347,N_652);
nand U1459 (N_1459,N_882,N_484);
nand U1460 (N_1460,N_57,N_575);
nor U1461 (N_1461,N_626,N_240);
nand U1462 (N_1462,N_951,N_59);
and U1463 (N_1463,N_938,N_568);
or U1464 (N_1464,N_187,N_901);
nor U1465 (N_1465,N_544,N_996);
and U1466 (N_1466,N_268,N_287);
nand U1467 (N_1467,N_379,N_471);
and U1468 (N_1468,N_535,N_181);
and U1469 (N_1469,N_37,N_362);
and U1470 (N_1470,N_705,N_259);
or U1471 (N_1471,N_161,N_834);
or U1472 (N_1472,N_732,N_848);
and U1473 (N_1473,N_485,N_56);
and U1474 (N_1474,N_76,N_727);
nand U1475 (N_1475,N_862,N_445);
nand U1476 (N_1476,N_906,N_197);
nor U1477 (N_1477,N_55,N_479);
and U1478 (N_1478,N_752,N_857);
or U1479 (N_1479,N_279,N_667);
nand U1480 (N_1480,N_467,N_298);
and U1481 (N_1481,N_946,N_456);
or U1482 (N_1482,N_154,N_531);
xor U1483 (N_1483,N_252,N_357);
or U1484 (N_1484,N_659,N_200);
or U1485 (N_1485,N_439,N_738);
or U1486 (N_1486,N_476,N_273);
and U1487 (N_1487,N_664,N_683);
nor U1488 (N_1488,N_962,N_369);
and U1489 (N_1489,N_49,N_464);
or U1490 (N_1490,N_67,N_141);
nor U1491 (N_1491,N_430,N_419);
nor U1492 (N_1492,N_295,N_375);
or U1493 (N_1493,N_679,N_624);
and U1494 (N_1494,N_30,N_253);
nand U1495 (N_1495,N_691,N_953);
and U1496 (N_1496,N_474,N_662);
nor U1497 (N_1497,N_641,N_180);
and U1498 (N_1498,N_718,N_75);
nand U1499 (N_1499,N_978,N_663);
or U1500 (N_1500,N_453,N_291);
nand U1501 (N_1501,N_738,N_615);
or U1502 (N_1502,N_448,N_788);
nand U1503 (N_1503,N_775,N_562);
or U1504 (N_1504,N_75,N_878);
nor U1505 (N_1505,N_450,N_887);
nor U1506 (N_1506,N_448,N_883);
nand U1507 (N_1507,N_685,N_75);
nand U1508 (N_1508,N_953,N_420);
nor U1509 (N_1509,N_759,N_704);
and U1510 (N_1510,N_873,N_789);
or U1511 (N_1511,N_159,N_366);
nor U1512 (N_1512,N_858,N_238);
nand U1513 (N_1513,N_299,N_433);
nand U1514 (N_1514,N_904,N_943);
or U1515 (N_1515,N_620,N_579);
nor U1516 (N_1516,N_451,N_799);
and U1517 (N_1517,N_776,N_969);
nand U1518 (N_1518,N_512,N_579);
nor U1519 (N_1519,N_897,N_485);
nor U1520 (N_1520,N_959,N_308);
nor U1521 (N_1521,N_113,N_278);
nand U1522 (N_1522,N_280,N_427);
nor U1523 (N_1523,N_732,N_233);
nor U1524 (N_1524,N_482,N_561);
and U1525 (N_1525,N_408,N_293);
or U1526 (N_1526,N_771,N_788);
and U1527 (N_1527,N_338,N_322);
nor U1528 (N_1528,N_841,N_813);
nor U1529 (N_1529,N_78,N_379);
xor U1530 (N_1530,N_787,N_839);
nor U1531 (N_1531,N_773,N_753);
and U1532 (N_1532,N_320,N_699);
xor U1533 (N_1533,N_27,N_877);
or U1534 (N_1534,N_279,N_865);
nand U1535 (N_1535,N_33,N_190);
nand U1536 (N_1536,N_806,N_970);
or U1537 (N_1537,N_527,N_808);
or U1538 (N_1538,N_530,N_244);
and U1539 (N_1539,N_936,N_799);
and U1540 (N_1540,N_8,N_369);
nor U1541 (N_1541,N_792,N_519);
nor U1542 (N_1542,N_911,N_759);
nor U1543 (N_1543,N_177,N_837);
and U1544 (N_1544,N_957,N_39);
and U1545 (N_1545,N_344,N_997);
xor U1546 (N_1546,N_859,N_365);
nand U1547 (N_1547,N_406,N_857);
nor U1548 (N_1548,N_429,N_957);
nand U1549 (N_1549,N_978,N_283);
nand U1550 (N_1550,N_61,N_523);
or U1551 (N_1551,N_560,N_840);
nand U1552 (N_1552,N_111,N_56);
nor U1553 (N_1553,N_408,N_401);
nor U1554 (N_1554,N_926,N_13);
nand U1555 (N_1555,N_4,N_217);
nor U1556 (N_1556,N_243,N_897);
and U1557 (N_1557,N_568,N_375);
nor U1558 (N_1558,N_54,N_239);
and U1559 (N_1559,N_721,N_869);
nor U1560 (N_1560,N_737,N_399);
nor U1561 (N_1561,N_694,N_822);
or U1562 (N_1562,N_748,N_659);
and U1563 (N_1563,N_136,N_410);
and U1564 (N_1564,N_441,N_338);
or U1565 (N_1565,N_361,N_871);
nor U1566 (N_1566,N_698,N_303);
nand U1567 (N_1567,N_277,N_159);
or U1568 (N_1568,N_138,N_859);
nor U1569 (N_1569,N_361,N_445);
or U1570 (N_1570,N_193,N_67);
nor U1571 (N_1571,N_478,N_744);
or U1572 (N_1572,N_698,N_67);
nand U1573 (N_1573,N_115,N_396);
and U1574 (N_1574,N_423,N_12);
and U1575 (N_1575,N_64,N_923);
nor U1576 (N_1576,N_882,N_209);
nand U1577 (N_1577,N_923,N_473);
nand U1578 (N_1578,N_660,N_969);
or U1579 (N_1579,N_12,N_139);
nor U1580 (N_1580,N_579,N_672);
or U1581 (N_1581,N_189,N_598);
nand U1582 (N_1582,N_718,N_316);
nand U1583 (N_1583,N_111,N_749);
nand U1584 (N_1584,N_699,N_636);
nand U1585 (N_1585,N_985,N_874);
nand U1586 (N_1586,N_370,N_50);
nor U1587 (N_1587,N_147,N_572);
and U1588 (N_1588,N_213,N_246);
nor U1589 (N_1589,N_272,N_69);
nor U1590 (N_1590,N_55,N_202);
and U1591 (N_1591,N_918,N_865);
nand U1592 (N_1592,N_567,N_974);
or U1593 (N_1593,N_535,N_898);
or U1594 (N_1594,N_174,N_57);
and U1595 (N_1595,N_116,N_691);
and U1596 (N_1596,N_780,N_70);
nand U1597 (N_1597,N_553,N_947);
and U1598 (N_1598,N_102,N_347);
or U1599 (N_1599,N_42,N_675);
or U1600 (N_1600,N_68,N_516);
or U1601 (N_1601,N_797,N_806);
nor U1602 (N_1602,N_482,N_585);
or U1603 (N_1603,N_874,N_458);
or U1604 (N_1604,N_752,N_838);
nor U1605 (N_1605,N_873,N_864);
nand U1606 (N_1606,N_836,N_114);
and U1607 (N_1607,N_132,N_904);
nand U1608 (N_1608,N_511,N_186);
and U1609 (N_1609,N_366,N_725);
or U1610 (N_1610,N_980,N_503);
or U1611 (N_1611,N_46,N_495);
or U1612 (N_1612,N_911,N_993);
nor U1613 (N_1613,N_379,N_695);
and U1614 (N_1614,N_338,N_181);
and U1615 (N_1615,N_112,N_819);
nand U1616 (N_1616,N_864,N_912);
nand U1617 (N_1617,N_45,N_873);
xor U1618 (N_1618,N_726,N_440);
and U1619 (N_1619,N_55,N_623);
and U1620 (N_1620,N_271,N_0);
or U1621 (N_1621,N_696,N_556);
nand U1622 (N_1622,N_581,N_389);
nor U1623 (N_1623,N_494,N_96);
xnor U1624 (N_1624,N_457,N_694);
nor U1625 (N_1625,N_518,N_979);
or U1626 (N_1626,N_526,N_875);
and U1627 (N_1627,N_209,N_772);
or U1628 (N_1628,N_757,N_299);
and U1629 (N_1629,N_862,N_651);
nand U1630 (N_1630,N_157,N_763);
nand U1631 (N_1631,N_45,N_668);
and U1632 (N_1632,N_815,N_201);
nor U1633 (N_1633,N_715,N_589);
nand U1634 (N_1634,N_347,N_611);
nand U1635 (N_1635,N_20,N_632);
nor U1636 (N_1636,N_148,N_792);
nor U1637 (N_1637,N_732,N_960);
and U1638 (N_1638,N_903,N_484);
or U1639 (N_1639,N_824,N_722);
nand U1640 (N_1640,N_497,N_316);
nand U1641 (N_1641,N_42,N_961);
or U1642 (N_1642,N_76,N_797);
or U1643 (N_1643,N_365,N_884);
and U1644 (N_1644,N_742,N_712);
nor U1645 (N_1645,N_801,N_358);
nand U1646 (N_1646,N_938,N_834);
nand U1647 (N_1647,N_681,N_605);
xnor U1648 (N_1648,N_319,N_13);
or U1649 (N_1649,N_503,N_685);
and U1650 (N_1650,N_427,N_696);
and U1651 (N_1651,N_941,N_376);
nand U1652 (N_1652,N_245,N_573);
nor U1653 (N_1653,N_573,N_42);
or U1654 (N_1654,N_926,N_269);
or U1655 (N_1655,N_399,N_992);
nor U1656 (N_1656,N_213,N_328);
nor U1657 (N_1657,N_586,N_795);
nand U1658 (N_1658,N_740,N_477);
nor U1659 (N_1659,N_613,N_722);
nand U1660 (N_1660,N_505,N_924);
or U1661 (N_1661,N_761,N_697);
and U1662 (N_1662,N_551,N_780);
nand U1663 (N_1663,N_474,N_166);
nand U1664 (N_1664,N_817,N_26);
and U1665 (N_1665,N_264,N_516);
and U1666 (N_1666,N_945,N_416);
nor U1667 (N_1667,N_552,N_634);
and U1668 (N_1668,N_718,N_488);
nand U1669 (N_1669,N_813,N_357);
and U1670 (N_1670,N_66,N_342);
and U1671 (N_1671,N_786,N_31);
or U1672 (N_1672,N_475,N_700);
and U1673 (N_1673,N_630,N_548);
or U1674 (N_1674,N_319,N_171);
nor U1675 (N_1675,N_916,N_614);
and U1676 (N_1676,N_759,N_473);
and U1677 (N_1677,N_594,N_784);
nor U1678 (N_1678,N_600,N_673);
nor U1679 (N_1679,N_506,N_765);
nand U1680 (N_1680,N_407,N_261);
and U1681 (N_1681,N_910,N_534);
nor U1682 (N_1682,N_163,N_680);
nand U1683 (N_1683,N_219,N_225);
and U1684 (N_1684,N_530,N_228);
nand U1685 (N_1685,N_923,N_508);
and U1686 (N_1686,N_36,N_576);
nand U1687 (N_1687,N_443,N_415);
nand U1688 (N_1688,N_504,N_231);
xor U1689 (N_1689,N_545,N_94);
nor U1690 (N_1690,N_734,N_355);
nand U1691 (N_1691,N_395,N_182);
or U1692 (N_1692,N_691,N_992);
nor U1693 (N_1693,N_965,N_113);
or U1694 (N_1694,N_690,N_314);
nor U1695 (N_1695,N_67,N_834);
or U1696 (N_1696,N_428,N_246);
and U1697 (N_1697,N_538,N_137);
and U1698 (N_1698,N_559,N_279);
or U1699 (N_1699,N_286,N_177);
nand U1700 (N_1700,N_207,N_996);
and U1701 (N_1701,N_474,N_38);
nor U1702 (N_1702,N_697,N_767);
and U1703 (N_1703,N_145,N_718);
nand U1704 (N_1704,N_875,N_909);
nor U1705 (N_1705,N_39,N_296);
nand U1706 (N_1706,N_75,N_913);
and U1707 (N_1707,N_773,N_848);
or U1708 (N_1708,N_957,N_13);
nand U1709 (N_1709,N_292,N_436);
nor U1710 (N_1710,N_345,N_592);
nand U1711 (N_1711,N_27,N_463);
or U1712 (N_1712,N_859,N_244);
and U1713 (N_1713,N_268,N_81);
and U1714 (N_1714,N_485,N_842);
xnor U1715 (N_1715,N_671,N_195);
or U1716 (N_1716,N_601,N_60);
nand U1717 (N_1717,N_482,N_144);
or U1718 (N_1718,N_916,N_555);
nor U1719 (N_1719,N_336,N_928);
nand U1720 (N_1720,N_914,N_563);
and U1721 (N_1721,N_978,N_949);
and U1722 (N_1722,N_326,N_665);
nor U1723 (N_1723,N_206,N_598);
nor U1724 (N_1724,N_747,N_241);
or U1725 (N_1725,N_517,N_831);
or U1726 (N_1726,N_813,N_756);
nor U1727 (N_1727,N_495,N_250);
and U1728 (N_1728,N_909,N_49);
or U1729 (N_1729,N_944,N_563);
and U1730 (N_1730,N_196,N_39);
and U1731 (N_1731,N_751,N_585);
or U1732 (N_1732,N_416,N_217);
and U1733 (N_1733,N_430,N_353);
nand U1734 (N_1734,N_435,N_304);
nor U1735 (N_1735,N_888,N_494);
or U1736 (N_1736,N_220,N_644);
xnor U1737 (N_1737,N_285,N_62);
nor U1738 (N_1738,N_806,N_163);
and U1739 (N_1739,N_705,N_173);
and U1740 (N_1740,N_636,N_591);
nor U1741 (N_1741,N_893,N_202);
and U1742 (N_1742,N_517,N_586);
and U1743 (N_1743,N_164,N_155);
and U1744 (N_1744,N_364,N_59);
and U1745 (N_1745,N_197,N_179);
nor U1746 (N_1746,N_178,N_999);
and U1747 (N_1747,N_463,N_427);
nand U1748 (N_1748,N_360,N_129);
and U1749 (N_1749,N_242,N_799);
or U1750 (N_1750,N_664,N_202);
nor U1751 (N_1751,N_476,N_810);
or U1752 (N_1752,N_533,N_232);
or U1753 (N_1753,N_642,N_701);
nor U1754 (N_1754,N_206,N_57);
and U1755 (N_1755,N_880,N_718);
and U1756 (N_1756,N_733,N_709);
nor U1757 (N_1757,N_132,N_870);
or U1758 (N_1758,N_299,N_328);
nor U1759 (N_1759,N_34,N_340);
or U1760 (N_1760,N_687,N_529);
and U1761 (N_1761,N_422,N_469);
and U1762 (N_1762,N_372,N_845);
and U1763 (N_1763,N_427,N_579);
xor U1764 (N_1764,N_161,N_382);
and U1765 (N_1765,N_535,N_395);
nand U1766 (N_1766,N_477,N_373);
and U1767 (N_1767,N_991,N_972);
nand U1768 (N_1768,N_730,N_651);
nor U1769 (N_1769,N_82,N_860);
and U1770 (N_1770,N_577,N_136);
nand U1771 (N_1771,N_366,N_404);
nor U1772 (N_1772,N_458,N_168);
and U1773 (N_1773,N_612,N_17);
nor U1774 (N_1774,N_699,N_778);
nor U1775 (N_1775,N_588,N_500);
xor U1776 (N_1776,N_537,N_838);
nand U1777 (N_1777,N_804,N_389);
nor U1778 (N_1778,N_153,N_227);
and U1779 (N_1779,N_165,N_567);
nor U1780 (N_1780,N_843,N_64);
nor U1781 (N_1781,N_873,N_40);
nand U1782 (N_1782,N_219,N_104);
nand U1783 (N_1783,N_227,N_873);
nand U1784 (N_1784,N_258,N_128);
or U1785 (N_1785,N_669,N_759);
and U1786 (N_1786,N_723,N_885);
and U1787 (N_1787,N_235,N_849);
or U1788 (N_1788,N_794,N_952);
nand U1789 (N_1789,N_514,N_660);
or U1790 (N_1790,N_652,N_184);
nand U1791 (N_1791,N_582,N_746);
or U1792 (N_1792,N_338,N_133);
or U1793 (N_1793,N_165,N_299);
nor U1794 (N_1794,N_73,N_724);
or U1795 (N_1795,N_572,N_699);
nor U1796 (N_1796,N_175,N_473);
nor U1797 (N_1797,N_609,N_13);
and U1798 (N_1798,N_908,N_20);
and U1799 (N_1799,N_327,N_127);
nand U1800 (N_1800,N_314,N_806);
nor U1801 (N_1801,N_129,N_413);
nor U1802 (N_1802,N_926,N_141);
xnor U1803 (N_1803,N_130,N_353);
nand U1804 (N_1804,N_310,N_739);
or U1805 (N_1805,N_467,N_286);
nor U1806 (N_1806,N_191,N_425);
or U1807 (N_1807,N_196,N_908);
and U1808 (N_1808,N_357,N_376);
or U1809 (N_1809,N_734,N_617);
and U1810 (N_1810,N_921,N_668);
nor U1811 (N_1811,N_258,N_891);
and U1812 (N_1812,N_97,N_899);
and U1813 (N_1813,N_278,N_536);
nand U1814 (N_1814,N_462,N_814);
nor U1815 (N_1815,N_741,N_481);
nand U1816 (N_1816,N_38,N_197);
or U1817 (N_1817,N_690,N_960);
nand U1818 (N_1818,N_204,N_601);
nor U1819 (N_1819,N_771,N_480);
and U1820 (N_1820,N_867,N_333);
or U1821 (N_1821,N_904,N_47);
nor U1822 (N_1822,N_794,N_662);
and U1823 (N_1823,N_959,N_966);
nor U1824 (N_1824,N_405,N_884);
and U1825 (N_1825,N_280,N_596);
nor U1826 (N_1826,N_174,N_800);
nor U1827 (N_1827,N_544,N_397);
nor U1828 (N_1828,N_116,N_485);
nand U1829 (N_1829,N_726,N_532);
and U1830 (N_1830,N_276,N_939);
nor U1831 (N_1831,N_941,N_174);
nand U1832 (N_1832,N_318,N_923);
or U1833 (N_1833,N_90,N_106);
nand U1834 (N_1834,N_642,N_949);
nor U1835 (N_1835,N_784,N_551);
nand U1836 (N_1836,N_961,N_261);
nor U1837 (N_1837,N_889,N_157);
or U1838 (N_1838,N_833,N_848);
nor U1839 (N_1839,N_187,N_725);
and U1840 (N_1840,N_320,N_963);
nor U1841 (N_1841,N_222,N_132);
nand U1842 (N_1842,N_725,N_757);
or U1843 (N_1843,N_248,N_2);
or U1844 (N_1844,N_846,N_38);
or U1845 (N_1845,N_746,N_679);
nand U1846 (N_1846,N_820,N_81);
and U1847 (N_1847,N_121,N_847);
nor U1848 (N_1848,N_78,N_713);
and U1849 (N_1849,N_328,N_217);
nand U1850 (N_1850,N_71,N_822);
and U1851 (N_1851,N_290,N_936);
xor U1852 (N_1852,N_152,N_130);
xor U1853 (N_1853,N_334,N_227);
or U1854 (N_1854,N_436,N_352);
nand U1855 (N_1855,N_173,N_40);
and U1856 (N_1856,N_473,N_752);
or U1857 (N_1857,N_768,N_547);
or U1858 (N_1858,N_827,N_517);
or U1859 (N_1859,N_999,N_176);
or U1860 (N_1860,N_845,N_529);
or U1861 (N_1861,N_797,N_196);
nand U1862 (N_1862,N_676,N_389);
or U1863 (N_1863,N_312,N_273);
or U1864 (N_1864,N_565,N_777);
or U1865 (N_1865,N_108,N_233);
nor U1866 (N_1866,N_314,N_803);
xnor U1867 (N_1867,N_81,N_256);
nor U1868 (N_1868,N_266,N_978);
nand U1869 (N_1869,N_452,N_45);
nor U1870 (N_1870,N_682,N_151);
nand U1871 (N_1871,N_663,N_901);
or U1872 (N_1872,N_784,N_927);
and U1873 (N_1873,N_846,N_989);
nand U1874 (N_1874,N_700,N_950);
and U1875 (N_1875,N_136,N_688);
or U1876 (N_1876,N_283,N_760);
and U1877 (N_1877,N_804,N_770);
nand U1878 (N_1878,N_698,N_181);
nor U1879 (N_1879,N_506,N_795);
nand U1880 (N_1880,N_590,N_450);
and U1881 (N_1881,N_576,N_795);
nand U1882 (N_1882,N_304,N_545);
and U1883 (N_1883,N_439,N_786);
nand U1884 (N_1884,N_332,N_101);
and U1885 (N_1885,N_787,N_692);
xor U1886 (N_1886,N_104,N_177);
and U1887 (N_1887,N_660,N_336);
nor U1888 (N_1888,N_464,N_54);
nor U1889 (N_1889,N_61,N_508);
and U1890 (N_1890,N_676,N_585);
nor U1891 (N_1891,N_835,N_519);
and U1892 (N_1892,N_240,N_20);
nand U1893 (N_1893,N_889,N_236);
nor U1894 (N_1894,N_440,N_364);
or U1895 (N_1895,N_92,N_112);
and U1896 (N_1896,N_550,N_209);
nor U1897 (N_1897,N_966,N_766);
nand U1898 (N_1898,N_995,N_335);
and U1899 (N_1899,N_144,N_267);
or U1900 (N_1900,N_185,N_5);
or U1901 (N_1901,N_716,N_849);
nand U1902 (N_1902,N_948,N_130);
nand U1903 (N_1903,N_903,N_333);
or U1904 (N_1904,N_104,N_116);
nand U1905 (N_1905,N_704,N_24);
nand U1906 (N_1906,N_571,N_217);
nor U1907 (N_1907,N_646,N_721);
nand U1908 (N_1908,N_975,N_738);
or U1909 (N_1909,N_49,N_264);
or U1910 (N_1910,N_386,N_556);
nand U1911 (N_1911,N_590,N_70);
and U1912 (N_1912,N_826,N_672);
nor U1913 (N_1913,N_147,N_200);
nor U1914 (N_1914,N_337,N_621);
nand U1915 (N_1915,N_882,N_291);
nor U1916 (N_1916,N_643,N_946);
xnor U1917 (N_1917,N_329,N_396);
nor U1918 (N_1918,N_773,N_543);
nand U1919 (N_1919,N_930,N_126);
or U1920 (N_1920,N_260,N_224);
nand U1921 (N_1921,N_763,N_963);
and U1922 (N_1922,N_224,N_890);
nand U1923 (N_1923,N_789,N_803);
and U1924 (N_1924,N_574,N_589);
and U1925 (N_1925,N_10,N_359);
nor U1926 (N_1926,N_630,N_18);
or U1927 (N_1927,N_245,N_526);
nor U1928 (N_1928,N_671,N_168);
or U1929 (N_1929,N_41,N_162);
or U1930 (N_1930,N_426,N_435);
and U1931 (N_1931,N_662,N_765);
or U1932 (N_1932,N_50,N_211);
nand U1933 (N_1933,N_771,N_559);
nor U1934 (N_1934,N_156,N_672);
nor U1935 (N_1935,N_711,N_394);
nand U1936 (N_1936,N_802,N_532);
and U1937 (N_1937,N_799,N_956);
or U1938 (N_1938,N_955,N_908);
and U1939 (N_1939,N_900,N_160);
nor U1940 (N_1940,N_587,N_636);
and U1941 (N_1941,N_839,N_900);
nor U1942 (N_1942,N_215,N_616);
xor U1943 (N_1943,N_976,N_948);
nor U1944 (N_1944,N_108,N_434);
or U1945 (N_1945,N_618,N_168);
nand U1946 (N_1946,N_923,N_167);
nand U1947 (N_1947,N_727,N_383);
nand U1948 (N_1948,N_367,N_649);
or U1949 (N_1949,N_120,N_746);
and U1950 (N_1950,N_952,N_420);
nand U1951 (N_1951,N_15,N_366);
nand U1952 (N_1952,N_121,N_101);
nand U1953 (N_1953,N_406,N_982);
or U1954 (N_1954,N_238,N_746);
nand U1955 (N_1955,N_190,N_282);
nor U1956 (N_1956,N_897,N_332);
and U1957 (N_1957,N_991,N_790);
nand U1958 (N_1958,N_530,N_933);
nand U1959 (N_1959,N_427,N_620);
nand U1960 (N_1960,N_891,N_743);
or U1961 (N_1961,N_16,N_770);
or U1962 (N_1962,N_90,N_122);
nand U1963 (N_1963,N_48,N_518);
and U1964 (N_1964,N_587,N_508);
or U1965 (N_1965,N_44,N_99);
or U1966 (N_1966,N_616,N_491);
nand U1967 (N_1967,N_684,N_161);
nand U1968 (N_1968,N_196,N_128);
or U1969 (N_1969,N_438,N_312);
nor U1970 (N_1970,N_452,N_924);
nand U1971 (N_1971,N_786,N_546);
nand U1972 (N_1972,N_725,N_180);
or U1973 (N_1973,N_794,N_210);
nor U1974 (N_1974,N_932,N_698);
and U1975 (N_1975,N_248,N_941);
nand U1976 (N_1976,N_960,N_767);
nand U1977 (N_1977,N_305,N_774);
nor U1978 (N_1978,N_608,N_506);
or U1979 (N_1979,N_20,N_771);
nor U1980 (N_1980,N_630,N_484);
and U1981 (N_1981,N_621,N_633);
nor U1982 (N_1982,N_394,N_213);
nand U1983 (N_1983,N_272,N_550);
or U1984 (N_1984,N_428,N_342);
nand U1985 (N_1985,N_378,N_202);
and U1986 (N_1986,N_622,N_165);
nor U1987 (N_1987,N_252,N_987);
nor U1988 (N_1988,N_574,N_132);
nor U1989 (N_1989,N_934,N_46);
nor U1990 (N_1990,N_716,N_639);
and U1991 (N_1991,N_970,N_430);
and U1992 (N_1992,N_498,N_130);
and U1993 (N_1993,N_294,N_443);
nor U1994 (N_1994,N_564,N_151);
or U1995 (N_1995,N_696,N_233);
or U1996 (N_1996,N_94,N_795);
nor U1997 (N_1997,N_787,N_746);
nor U1998 (N_1998,N_474,N_603);
nand U1999 (N_1999,N_140,N_121);
or U2000 (N_2000,N_1667,N_1911);
nand U2001 (N_2001,N_1382,N_1362);
or U2002 (N_2002,N_1358,N_1521);
nand U2003 (N_2003,N_1343,N_1914);
or U2004 (N_2004,N_1162,N_1950);
nor U2005 (N_2005,N_1140,N_1683);
and U2006 (N_2006,N_1957,N_1067);
or U2007 (N_2007,N_1388,N_1026);
and U2008 (N_2008,N_1621,N_1841);
xor U2009 (N_2009,N_1701,N_1478);
and U2010 (N_2010,N_1090,N_1978);
or U2011 (N_2011,N_1337,N_1158);
and U2012 (N_2012,N_1271,N_1879);
and U2013 (N_2013,N_1689,N_1627);
or U2014 (N_2014,N_1599,N_1406);
nor U2015 (N_2015,N_1850,N_1589);
nor U2016 (N_2016,N_1348,N_1369);
nor U2017 (N_2017,N_1792,N_1440);
nand U2018 (N_2018,N_1344,N_1138);
and U2019 (N_2019,N_1458,N_1125);
and U2020 (N_2020,N_1577,N_1722);
nor U2021 (N_2021,N_1314,N_1568);
or U2022 (N_2022,N_1353,N_1919);
and U2023 (N_2023,N_1244,N_1432);
nand U2024 (N_2024,N_1112,N_1059);
and U2025 (N_2025,N_1718,N_1964);
nand U2026 (N_2026,N_1329,N_1876);
or U2027 (N_2027,N_1053,N_1756);
nand U2028 (N_2028,N_1601,N_1522);
and U2029 (N_2029,N_1100,N_1130);
and U2030 (N_2030,N_1154,N_1014);
or U2031 (N_2031,N_1468,N_1893);
nor U2032 (N_2032,N_1085,N_1019);
and U2033 (N_2033,N_1632,N_1526);
nand U2034 (N_2034,N_1381,N_1352);
xor U2035 (N_2035,N_1096,N_1205);
or U2036 (N_2036,N_1342,N_1239);
or U2037 (N_2037,N_1598,N_1617);
nor U2038 (N_2038,N_1071,N_1608);
nor U2039 (N_2039,N_1425,N_1646);
nor U2040 (N_2040,N_1098,N_1769);
nor U2041 (N_2041,N_1423,N_1419);
nor U2042 (N_2042,N_1028,N_1603);
and U2043 (N_2043,N_1541,N_1490);
and U2044 (N_2044,N_1538,N_1361);
nand U2045 (N_2045,N_1120,N_1084);
nor U2046 (N_2046,N_1315,N_1954);
nor U2047 (N_2047,N_1637,N_1581);
and U2048 (N_2048,N_1961,N_1414);
or U2049 (N_2049,N_1706,N_1547);
or U2050 (N_2050,N_1629,N_1684);
nand U2051 (N_2051,N_1102,N_1437);
nor U2052 (N_2052,N_1131,N_1234);
nand U2053 (N_2053,N_1256,N_1228);
nor U2054 (N_2054,N_1293,N_1820);
nand U2055 (N_2055,N_1669,N_1346);
and U2056 (N_2056,N_1114,N_1366);
or U2057 (N_2057,N_1695,N_1659);
and U2058 (N_2058,N_1697,N_1472);
nand U2059 (N_2059,N_1106,N_1707);
nor U2060 (N_2060,N_1012,N_1741);
nor U2061 (N_2061,N_1364,N_1363);
or U2062 (N_2062,N_1262,N_1279);
nand U2063 (N_2063,N_1563,N_1980);
nand U2064 (N_2064,N_1874,N_1378);
or U2065 (N_2065,N_1996,N_1811);
or U2066 (N_2066,N_1951,N_1188);
nor U2067 (N_2067,N_1748,N_1123);
nand U2068 (N_2068,N_1595,N_1297);
nand U2069 (N_2069,N_1415,N_1524);
or U2070 (N_2070,N_1967,N_1172);
and U2071 (N_2071,N_1851,N_1430);
nor U2072 (N_2072,N_1405,N_1104);
nor U2073 (N_2073,N_1076,N_1968);
or U2074 (N_2074,N_1576,N_1010);
nor U2075 (N_2075,N_1549,N_1987);
xnor U2076 (N_2076,N_1194,N_1069);
or U2077 (N_2077,N_1909,N_1094);
or U2078 (N_2078,N_1157,N_1221);
nor U2079 (N_2079,N_1605,N_1898);
nand U2080 (N_2080,N_1803,N_1556);
or U2081 (N_2081,N_1530,N_1207);
nor U2082 (N_2082,N_1491,N_1159);
and U2083 (N_2083,N_1034,N_1307);
nor U2084 (N_2084,N_1087,N_1775);
nor U2085 (N_2085,N_1002,N_1716);
nor U2086 (N_2086,N_1270,N_1875);
nor U2087 (N_2087,N_1955,N_1359);
nor U2088 (N_2088,N_1986,N_1141);
or U2089 (N_2089,N_1042,N_1241);
and U2090 (N_2090,N_1108,N_1052);
nand U2091 (N_2091,N_1523,N_1901);
or U2092 (N_2092,N_1011,N_1258);
nor U2093 (N_2093,N_1401,N_1077);
nor U2094 (N_2094,N_1110,N_1449);
nor U2095 (N_2095,N_1509,N_1858);
nor U2096 (N_2096,N_1306,N_1164);
nand U2097 (N_2097,N_1990,N_1135);
and U2098 (N_2098,N_1784,N_1918);
or U2099 (N_2099,N_1804,N_1899);
and U2100 (N_2100,N_1264,N_1673);
or U2101 (N_2101,N_1494,N_1339);
and U2102 (N_2102,N_1450,N_1309);
nand U2103 (N_2103,N_1166,N_1838);
nor U2104 (N_2104,N_1248,N_1025);
or U2105 (N_2105,N_1660,N_1311);
xnor U2106 (N_2106,N_1195,N_1808);
nand U2107 (N_2107,N_1712,N_1585);
and U2108 (N_2108,N_1463,N_1932);
nand U2109 (N_2109,N_1083,N_1249);
nor U2110 (N_2110,N_1906,N_1146);
or U2111 (N_2111,N_1434,N_1190);
or U2112 (N_2112,N_1299,N_1873);
nand U2113 (N_2113,N_1704,N_1007);
nand U2114 (N_2114,N_1261,N_1941);
and U2115 (N_2115,N_1044,N_1461);
nand U2116 (N_2116,N_1799,N_1182);
or U2117 (N_2117,N_1924,N_1615);
or U2118 (N_2118,N_1005,N_1762);
nand U2119 (N_2119,N_1744,N_1355);
nor U2120 (N_2120,N_1152,N_1101);
or U2121 (N_2121,N_1082,N_1252);
nor U2122 (N_2122,N_1760,N_1206);
xor U2123 (N_2123,N_1849,N_1956);
or U2124 (N_2124,N_1181,N_1066);
or U2125 (N_2125,N_1267,N_1230);
and U2126 (N_2126,N_1511,N_1073);
nor U2127 (N_2127,N_1810,N_1685);
or U2128 (N_2128,N_1829,N_1847);
nand U2129 (N_2129,N_1528,N_1481);
or U2130 (N_2130,N_1702,N_1947);
and U2131 (N_2131,N_1525,N_1675);
nor U2132 (N_2132,N_1429,N_1265);
nand U2133 (N_2133,N_1836,N_1935);
nor U2134 (N_2134,N_1086,N_1455);
and U2135 (N_2135,N_1477,N_1142);
and U2136 (N_2136,N_1554,N_1962);
nor U2137 (N_2137,N_1009,N_1859);
or U2138 (N_2138,N_1319,N_1537);
nor U2139 (N_2139,N_1118,N_1246);
nand U2140 (N_2140,N_1119,N_1553);
or U2141 (N_2141,N_1649,N_1211);
nor U2142 (N_2142,N_1180,N_1700);
and U2143 (N_2143,N_1383,N_1322);
nand U2144 (N_2144,N_1232,N_1217);
or U2145 (N_2145,N_1619,N_1604);
nand U2146 (N_2146,N_1767,N_1001);
or U2147 (N_2147,N_1374,N_1313);
nor U2148 (N_2148,N_1325,N_1593);
xnor U2149 (N_2149,N_1237,N_1690);
nand U2150 (N_2150,N_1652,N_1379);
nand U2151 (N_2151,N_1189,N_1668);
nand U2152 (N_2152,N_1122,N_1367);
or U2153 (N_2153,N_1570,N_1393);
and U2154 (N_2154,N_1946,N_1229);
and U2155 (N_2155,N_1451,N_1788);
and U2156 (N_2156,N_1498,N_1193);
and U2157 (N_2157,N_1179,N_1150);
nor U2158 (N_2158,N_1173,N_1630);
nor U2159 (N_2159,N_1433,N_1891);
and U2160 (N_2160,N_1506,N_1976);
nand U2161 (N_2161,N_1817,N_1070);
or U2162 (N_2162,N_1103,N_1269);
nor U2163 (N_2163,N_1726,N_1939);
nor U2164 (N_2164,N_1384,N_1360);
and U2165 (N_2165,N_1116,N_1653);
nor U2166 (N_2166,N_1963,N_1806);
and U2167 (N_2167,N_1705,N_1163);
and U2168 (N_2168,N_1796,N_1880);
nand U2169 (N_2169,N_1222,N_1143);
or U2170 (N_2170,N_1539,N_1895);
nor U2171 (N_2171,N_1065,N_1686);
and U2172 (N_2172,N_1613,N_1749);
and U2173 (N_2173,N_1137,N_1051);
and U2174 (N_2174,N_1959,N_1027);
nand U2175 (N_2175,N_1008,N_1356);
or U2176 (N_2176,N_1018,N_1156);
and U2177 (N_2177,N_1607,N_1949);
nor U2178 (N_2178,N_1520,N_1504);
nand U2179 (N_2179,N_1917,N_1109);
nand U2180 (N_2180,N_1965,N_1624);
and U2181 (N_2181,N_1183,N_1871);
nor U2182 (N_2182,N_1816,N_1291);
or U2183 (N_2183,N_1507,N_1147);
nand U2184 (N_2184,N_1282,N_1719);
and U2185 (N_2185,N_1960,N_1441);
nor U2186 (N_2186,N_1443,N_1212);
and U2187 (N_2187,N_1395,N_1943);
or U2188 (N_2188,N_1136,N_1856);
and U2189 (N_2189,N_1846,N_1715);
xor U2190 (N_2190,N_1663,N_1519);
nand U2191 (N_2191,N_1736,N_1128);
or U2192 (N_2192,N_1742,N_1412);
nand U2193 (N_2193,N_1492,N_1983);
nor U2194 (N_2194,N_1268,N_1371);
nand U2195 (N_2195,N_1679,N_1870);
nor U2196 (N_2196,N_1896,N_1410);
or U2197 (N_2197,N_1915,N_1869);
and U2198 (N_2198,N_1737,N_1835);
or U2199 (N_2199,N_1467,N_1226);
or U2200 (N_2200,N_1113,N_1703);
or U2201 (N_2201,N_1040,N_1332);
or U2202 (N_2202,N_1931,N_1644);
nand U2203 (N_2203,N_1017,N_1985);
nand U2204 (N_2204,N_1236,N_1782);
nor U2205 (N_2205,N_1628,N_1512);
and U2206 (N_2206,N_1739,N_1323);
nor U2207 (N_2207,N_1802,N_1885);
or U2208 (N_2208,N_1699,N_1013);
and U2209 (N_2209,N_1091,N_1370);
nand U2210 (N_2210,N_1828,N_1480);
or U2211 (N_2211,N_1198,N_1310);
nor U2212 (N_2212,N_1609,N_1517);
and U2213 (N_2213,N_1097,N_1584);
nand U2214 (N_2214,N_1691,N_1773);
or U2215 (N_2215,N_1015,N_1284);
and U2216 (N_2216,N_1940,N_1402);
nand U2217 (N_2217,N_1501,N_1709);
and U2218 (N_2218,N_1341,N_1532);
or U2219 (N_2219,N_1174,N_1529);
or U2220 (N_2220,N_1783,N_1151);
or U2221 (N_2221,N_1747,N_1635);
nand U2222 (N_2222,N_1732,N_1155);
nor U2223 (N_2223,N_1493,N_1694);
and U2224 (N_2224,N_1105,N_1555);
nor U2225 (N_2225,N_1698,N_1571);
or U2226 (N_2226,N_1030,N_1724);
nor U2227 (N_2227,N_1231,N_1459);
nand U2228 (N_2228,N_1016,N_1989);
and U2229 (N_2229,N_1175,N_1862);
nand U2230 (N_2230,N_1047,N_1446);
nand U2231 (N_2231,N_1641,N_1813);
nand U2232 (N_2232,N_1243,N_1148);
and U2233 (N_2233,N_1020,N_1385);
and U2234 (N_2234,N_1503,N_1745);
nor U2235 (N_2235,N_1717,N_1565);
nand U2236 (N_2236,N_1778,N_1992);
and U2237 (N_2237,N_1165,N_1647);
nand U2238 (N_2238,N_1942,N_1039);
or U2239 (N_2239,N_1215,N_1210);
or U2240 (N_2240,N_1111,N_1460);
or U2241 (N_2241,N_1734,N_1510);
nand U2242 (N_2242,N_1489,N_1768);
nor U2243 (N_2243,N_1582,N_1400);
nand U2244 (N_2244,N_1214,N_1320);
and U2245 (N_2245,N_1302,N_1305);
nand U2246 (N_2246,N_1822,N_1981);
nand U2247 (N_2247,N_1331,N_1857);
or U2248 (N_2248,N_1597,N_1612);
or U2249 (N_2249,N_1505,N_1833);
nand U2250 (N_2250,N_1024,N_1487);
nand U2251 (N_2251,N_1099,N_1396);
and U2252 (N_2252,N_1907,N_1693);
nor U2253 (N_2253,N_1334,N_1483);
nand U2254 (N_2254,N_1476,N_1250);
xor U2255 (N_2255,N_1304,N_1753);
or U2256 (N_2256,N_1516,N_1473);
or U2257 (N_2257,N_1386,N_1298);
or U2258 (N_2258,N_1133,N_1266);
nand U2259 (N_2259,N_1462,N_1674);
and U2260 (N_2260,N_1794,N_1095);
and U2261 (N_2261,N_1502,N_1966);
nor U2262 (N_2262,N_1764,N_1814);
or U2263 (N_2263,N_1454,N_1561);
nand U2264 (N_2264,N_1276,N_1872);
nand U2265 (N_2265,N_1973,N_1815);
nand U2266 (N_2266,N_1636,N_1390);
or U2267 (N_2267,N_1488,N_1184);
nor U2268 (N_2268,N_1057,N_1991);
and U2269 (N_2269,N_1245,N_1275);
nand U2270 (N_2270,N_1616,N_1448);
or U2271 (N_2271,N_1204,N_1273);
xor U2272 (N_2272,N_1733,N_1347);
and U2273 (N_2273,N_1470,N_1176);
nand U2274 (N_2274,N_1995,N_1678);
nand U2275 (N_2275,N_1912,N_1456);
nor U2276 (N_2276,N_1594,N_1127);
or U2277 (N_2277,N_1642,N_1890);
and U2278 (N_2278,N_1812,N_1727);
nor U2279 (N_2279,N_1830,N_1421);
nand U2280 (N_2280,N_1043,N_1933);
nor U2281 (N_2281,N_1560,N_1916);
nand U2282 (N_2282,N_1970,N_1735);
or U2283 (N_2283,N_1640,N_1575);
or U2284 (N_2284,N_1731,N_1000);
nor U2285 (N_2285,N_1495,N_1422);
or U2286 (N_2286,N_1373,N_1452);
nand U2287 (N_2287,N_1643,N_1786);
or U2288 (N_2288,N_1160,N_1639);
and U2289 (N_2289,N_1377,N_1479);
nor U2290 (N_2290,N_1281,N_1031);
nor U2291 (N_2291,N_1620,N_1790);
nor U2292 (N_2292,N_1787,N_1124);
and U2293 (N_2293,N_1169,N_1247);
and U2294 (N_2294,N_1149,N_1681);
and U2295 (N_2295,N_1417,N_1333);
nand U2296 (N_2296,N_1404,N_1442);
nand U2297 (N_2297,N_1260,N_1910);
or U2298 (N_2298,N_1546,N_1979);
nor U2299 (N_2299,N_1408,N_1327);
and U2300 (N_2300,N_1428,N_1397);
nor U2301 (N_2301,N_1038,N_1625);
or U2302 (N_2302,N_1614,N_1436);
and U2303 (N_2303,N_1394,N_1888);
and U2304 (N_2304,N_1336,N_1626);
or U2305 (N_2305,N_1021,N_1219);
nand U2306 (N_2306,N_1740,N_1825);
nor U2307 (N_2307,N_1721,N_1945);
nor U2308 (N_2308,N_1092,N_1171);
nor U2309 (N_2309,N_1278,N_1864);
nand U2310 (N_2310,N_1235,N_1682);
nand U2311 (N_2311,N_1930,N_1819);
and U2312 (N_2312,N_1426,N_1466);
or U2313 (N_2313,N_1080,N_1789);
and U2314 (N_2314,N_1671,N_1295);
or U2315 (N_2315,N_1781,N_1413);
nand U2316 (N_2316,N_1839,N_1666);
or U2317 (N_2317,N_1048,N_1225);
or U2318 (N_2318,N_1185,N_1167);
or U2319 (N_2319,N_1424,N_1622);
nand U2320 (N_2320,N_1904,N_1564);
or U2321 (N_2321,N_1557,N_1283);
and U2322 (N_2322,N_1062,N_1592);
nor U2323 (N_2323,N_1664,N_1312);
nand U2324 (N_2324,N_1469,N_1288);
nor U2325 (N_2325,N_1255,N_1937);
xor U2326 (N_2326,N_1208,N_1677);
nor U2327 (N_2327,N_1797,N_1178);
nor U2328 (N_2328,N_1944,N_1218);
nor U2329 (N_2329,N_1004,N_1216);
and U2330 (N_2330,N_1921,N_1757);
or U2331 (N_2331,N_1618,N_1848);
and U2332 (N_2332,N_1464,N_1958);
and U2333 (N_2333,N_1407,N_1447);
nand U2334 (N_2334,N_1006,N_1687);
or U2335 (N_2335,N_1316,N_1925);
nand U2336 (N_2336,N_1064,N_1531);
and U2337 (N_2337,N_1984,N_1170);
nand U2338 (N_2338,N_1752,N_1761);
and U2339 (N_2339,N_1894,N_1187);
or U2340 (N_2340,N_1350,N_1600);
nand U2341 (N_2341,N_1497,N_1153);
nor U2342 (N_2342,N_1439,N_1280);
nand U2343 (N_2343,N_1022,N_1903);
and U2344 (N_2344,N_1058,N_1060);
nand U2345 (N_2345,N_1126,N_1061);
and U2346 (N_2346,N_1496,N_1089);
and U2347 (N_2347,N_1380,N_1399);
and U2348 (N_2348,N_1289,N_1758);
and U2349 (N_2349,N_1807,N_1566);
xnor U2350 (N_2350,N_1286,N_1318);
nand U2351 (N_2351,N_1867,N_1431);
and U2352 (N_2352,N_1032,N_1948);
and U2353 (N_2353,N_1438,N_1499);
and U2354 (N_2354,N_1203,N_1777);
and U2355 (N_2355,N_1728,N_1238);
and U2356 (N_2356,N_1908,N_1435);
and U2357 (N_2357,N_1285,N_1661);
or U2358 (N_2358,N_1844,N_1586);
and U2359 (N_2359,N_1088,N_1068);
nor U2360 (N_2360,N_1515,N_1514);
nand U2361 (N_2361,N_1569,N_1486);
nor U2362 (N_2362,N_1036,N_1696);
nand U2363 (N_2363,N_1892,N_1656);
and U2364 (N_2364,N_1863,N_1411);
nand U2365 (N_2365,N_1633,N_1420);
nor U2366 (N_2366,N_1887,N_1121);
and U2367 (N_2367,N_1263,N_1177);
nand U2368 (N_2368,N_1200,N_1920);
or U2369 (N_2369,N_1993,N_1720);
nor U2370 (N_2370,N_1081,N_1793);
nor U2371 (N_2371,N_1834,N_1253);
and U2372 (N_2372,N_1913,N_1301);
and U2373 (N_2373,N_1975,N_1861);
nand U2374 (N_2374,N_1191,N_1711);
or U2375 (N_2375,N_1572,N_1772);
and U2376 (N_2376,N_1409,N_1129);
nor U2377 (N_2377,N_1843,N_1832);
nor U2378 (N_2378,N_1551,N_1453);
nor U2379 (N_2379,N_1115,N_1550);
nand U2380 (N_2380,N_1754,N_1387);
or U2381 (N_2381,N_1602,N_1578);
xnor U2382 (N_2382,N_1050,N_1317);
and U2383 (N_2383,N_1883,N_1227);
nand U2384 (N_2384,N_1886,N_1665);
nand U2385 (N_2385,N_1631,N_1638);
or U2386 (N_2386,N_1513,N_1771);
and U2387 (N_2387,N_1045,N_1465);
and U2388 (N_2388,N_1075,N_1324);
and U2389 (N_2389,N_1750,N_1676);
and U2390 (N_2390,N_1840,N_1054);
nand U2391 (N_2391,N_1199,N_1540);
xnor U2392 (N_2392,N_1596,N_1330);
nor U2393 (N_2393,N_1534,N_1821);
and U2394 (N_2394,N_1845,N_1527);
nand U2395 (N_2395,N_1779,N_1482);
nand U2396 (N_2396,N_1444,N_1934);
nor U2397 (N_2397,N_1938,N_1536);
nand U2398 (N_2398,N_1303,N_1117);
and U2399 (N_2399,N_1340,N_1798);
or U2400 (N_2400,N_1692,N_1795);
or U2401 (N_2401,N_1854,N_1389);
nand U2402 (N_2402,N_1474,N_1860);
or U2403 (N_2403,N_1063,N_1392);
nand U2404 (N_2404,N_1161,N_1606);
nand U2405 (N_2405,N_1257,N_1548);
nand U2406 (N_2406,N_1209,N_1831);
or U2407 (N_2407,N_1672,N_1800);
and U2408 (N_2408,N_1936,N_1651);
nand U2409 (N_2409,N_1823,N_1972);
nor U2410 (N_2410,N_1055,N_1977);
or U2411 (N_2411,N_1192,N_1926);
xor U2412 (N_2412,N_1927,N_1791);
nand U2413 (N_2413,N_1445,N_1372);
or U2414 (N_2414,N_1923,N_1139);
nor U2415 (N_2415,N_1579,N_1662);
nor U2416 (N_2416,N_1023,N_1866);
or U2417 (N_2417,N_1837,N_1457);
or U2418 (N_2418,N_1865,N_1999);
nor U2419 (N_2419,N_1552,N_1994);
nor U2420 (N_2420,N_1558,N_1535);
or U2421 (N_2421,N_1738,N_1645);
or U2422 (N_2422,N_1824,N_1878);
and U2423 (N_2423,N_1375,N_1277);
and U2424 (N_2424,N_1922,N_1544);
nor U2425 (N_2425,N_1475,N_1345);
nand U2426 (N_2426,N_1416,N_1670);
nand U2427 (N_2427,N_1376,N_1897);
or U2428 (N_2428,N_1326,N_1485);
nor U2429 (N_2429,N_1074,N_1533);
and U2430 (N_2430,N_1952,N_1292);
and U2431 (N_2431,N_1144,N_1583);
or U2432 (N_2432,N_1290,N_1902);
nor U2433 (N_2433,N_1623,N_1648);
and U2434 (N_2434,N_1308,N_1776);
nor U2435 (N_2435,N_1251,N_1801);
or U2436 (N_2436,N_1543,N_1971);
or U2437 (N_2437,N_1197,N_1766);
nand U2438 (N_2438,N_1770,N_1877);
nor U2439 (N_2439,N_1708,N_1559);
nand U2440 (N_2440,N_1785,N_1418);
nand U2441 (N_2441,N_1500,N_1805);
or U2442 (N_2442,N_1403,N_1471);
or U2443 (N_2443,N_1321,N_1997);
or U2444 (N_2444,N_1037,N_1328);
nand U2445 (N_2445,N_1714,N_1988);
and U2446 (N_2446,N_1729,N_1591);
nor U2447 (N_2447,N_1368,N_1658);
nor U2448 (N_2448,N_1233,N_1881);
nand U2449 (N_2449,N_1357,N_1855);
and U2450 (N_2450,N_1134,N_1884);
or U2451 (N_2451,N_1590,N_1033);
nor U2452 (N_2452,N_1774,N_1567);
nor U2453 (N_2453,N_1765,N_1562);
nand U2454 (N_2454,N_1780,N_1484);
or U2455 (N_2455,N_1542,N_1610);
nor U2456 (N_2456,N_1427,N_1049);
nand U2457 (N_2457,N_1029,N_1842);
nand U2458 (N_2458,N_1508,N_1391);
nand U2459 (N_2459,N_1518,N_1296);
nand U2460 (N_2460,N_1287,N_1650);
xor U2461 (N_2461,N_1853,N_1168);
nor U2462 (N_2462,N_1634,N_1079);
or U2463 (N_2463,N_1093,N_1035);
nand U2464 (N_2464,N_1611,N_1354);
nor U2465 (N_2465,N_1107,N_1259);
and U2466 (N_2466,N_1713,N_1969);
nor U2467 (N_2467,N_1186,N_1202);
nand U2468 (N_2468,N_1254,N_1349);
nor U2469 (N_2469,N_1294,N_1818);
nand U2470 (N_2470,N_1654,N_1809);
or U2471 (N_2471,N_1224,N_1974);
and U2472 (N_2472,N_1132,N_1827);
and U2473 (N_2473,N_1900,N_1545);
nand U2474 (N_2474,N_1755,N_1240);
nor U2475 (N_2475,N_1220,N_1882);
xnor U2476 (N_2476,N_1587,N_1889);
nand U2477 (N_2477,N_1046,N_1998);
and U2478 (N_2478,N_1398,N_1300);
nor U2479 (N_2479,N_1574,N_1223);
and U2480 (N_2480,N_1953,N_1928);
nand U2481 (N_2481,N_1078,N_1688);
or U2482 (N_2482,N_1201,N_1274);
or U2483 (N_2483,N_1759,N_1335);
or U2484 (N_2484,N_1003,N_1723);
or U2485 (N_2485,N_1730,N_1929);
nor U2486 (N_2486,N_1751,N_1868);
nor U2487 (N_2487,N_1056,N_1213);
nand U2488 (N_2488,N_1580,N_1145);
nand U2489 (N_2489,N_1826,N_1746);
or U2490 (N_2490,N_1072,N_1196);
and U2491 (N_2491,N_1041,N_1351);
nand U2492 (N_2492,N_1743,N_1852);
nor U2493 (N_2493,N_1588,N_1982);
and U2494 (N_2494,N_1725,N_1272);
and U2495 (N_2495,N_1338,N_1710);
and U2496 (N_2496,N_1242,N_1573);
or U2497 (N_2497,N_1680,N_1905);
nand U2498 (N_2498,N_1655,N_1657);
nor U2499 (N_2499,N_1763,N_1365);
and U2500 (N_2500,N_1148,N_1493);
and U2501 (N_2501,N_1416,N_1414);
and U2502 (N_2502,N_1759,N_1480);
nand U2503 (N_2503,N_1415,N_1452);
and U2504 (N_2504,N_1852,N_1818);
nand U2505 (N_2505,N_1621,N_1283);
nor U2506 (N_2506,N_1683,N_1648);
and U2507 (N_2507,N_1707,N_1738);
nor U2508 (N_2508,N_1970,N_1772);
and U2509 (N_2509,N_1090,N_1760);
or U2510 (N_2510,N_1434,N_1973);
and U2511 (N_2511,N_1043,N_1780);
or U2512 (N_2512,N_1627,N_1262);
nor U2513 (N_2513,N_1354,N_1816);
and U2514 (N_2514,N_1892,N_1890);
nand U2515 (N_2515,N_1742,N_1369);
nor U2516 (N_2516,N_1679,N_1700);
nor U2517 (N_2517,N_1989,N_1796);
nand U2518 (N_2518,N_1666,N_1172);
and U2519 (N_2519,N_1886,N_1878);
nand U2520 (N_2520,N_1410,N_1353);
nand U2521 (N_2521,N_1964,N_1970);
and U2522 (N_2522,N_1767,N_1655);
nand U2523 (N_2523,N_1076,N_1794);
nand U2524 (N_2524,N_1344,N_1063);
nand U2525 (N_2525,N_1489,N_1433);
or U2526 (N_2526,N_1524,N_1689);
nand U2527 (N_2527,N_1473,N_1457);
nor U2528 (N_2528,N_1894,N_1712);
nor U2529 (N_2529,N_1049,N_1575);
or U2530 (N_2530,N_1116,N_1447);
nor U2531 (N_2531,N_1081,N_1041);
or U2532 (N_2532,N_1030,N_1623);
and U2533 (N_2533,N_1318,N_1455);
nor U2534 (N_2534,N_1940,N_1174);
or U2535 (N_2535,N_1107,N_1780);
nand U2536 (N_2536,N_1598,N_1237);
and U2537 (N_2537,N_1711,N_1135);
or U2538 (N_2538,N_1182,N_1424);
nor U2539 (N_2539,N_1051,N_1125);
and U2540 (N_2540,N_1607,N_1322);
or U2541 (N_2541,N_1264,N_1179);
nand U2542 (N_2542,N_1488,N_1170);
nand U2543 (N_2543,N_1843,N_1383);
or U2544 (N_2544,N_1086,N_1674);
and U2545 (N_2545,N_1500,N_1352);
nor U2546 (N_2546,N_1309,N_1649);
and U2547 (N_2547,N_1936,N_1949);
nand U2548 (N_2548,N_1876,N_1998);
and U2549 (N_2549,N_1644,N_1664);
and U2550 (N_2550,N_1885,N_1934);
nand U2551 (N_2551,N_1344,N_1022);
and U2552 (N_2552,N_1237,N_1385);
nor U2553 (N_2553,N_1553,N_1008);
nor U2554 (N_2554,N_1996,N_1698);
or U2555 (N_2555,N_1584,N_1819);
or U2556 (N_2556,N_1389,N_1033);
and U2557 (N_2557,N_1694,N_1463);
or U2558 (N_2558,N_1874,N_1200);
nand U2559 (N_2559,N_1454,N_1105);
nor U2560 (N_2560,N_1985,N_1127);
nand U2561 (N_2561,N_1320,N_1326);
and U2562 (N_2562,N_1442,N_1256);
and U2563 (N_2563,N_1522,N_1258);
or U2564 (N_2564,N_1497,N_1719);
nand U2565 (N_2565,N_1230,N_1571);
and U2566 (N_2566,N_1538,N_1113);
or U2567 (N_2567,N_1292,N_1535);
nor U2568 (N_2568,N_1197,N_1190);
nor U2569 (N_2569,N_1408,N_1754);
nand U2570 (N_2570,N_1874,N_1607);
or U2571 (N_2571,N_1543,N_1526);
or U2572 (N_2572,N_1890,N_1922);
nor U2573 (N_2573,N_1886,N_1639);
nand U2574 (N_2574,N_1240,N_1037);
and U2575 (N_2575,N_1028,N_1801);
nor U2576 (N_2576,N_1626,N_1422);
nand U2577 (N_2577,N_1535,N_1534);
and U2578 (N_2578,N_1969,N_1134);
and U2579 (N_2579,N_1061,N_1644);
or U2580 (N_2580,N_1998,N_1085);
or U2581 (N_2581,N_1629,N_1973);
nor U2582 (N_2582,N_1904,N_1766);
or U2583 (N_2583,N_1249,N_1444);
or U2584 (N_2584,N_1866,N_1521);
or U2585 (N_2585,N_1896,N_1926);
nor U2586 (N_2586,N_1251,N_1105);
nand U2587 (N_2587,N_1582,N_1423);
nor U2588 (N_2588,N_1572,N_1233);
xnor U2589 (N_2589,N_1043,N_1276);
or U2590 (N_2590,N_1229,N_1321);
and U2591 (N_2591,N_1626,N_1108);
or U2592 (N_2592,N_1017,N_1516);
nor U2593 (N_2593,N_1371,N_1031);
xor U2594 (N_2594,N_1366,N_1902);
nor U2595 (N_2595,N_1116,N_1578);
nor U2596 (N_2596,N_1628,N_1170);
and U2597 (N_2597,N_1104,N_1023);
nand U2598 (N_2598,N_1127,N_1811);
and U2599 (N_2599,N_1519,N_1322);
nor U2600 (N_2600,N_1856,N_1700);
and U2601 (N_2601,N_1465,N_1795);
and U2602 (N_2602,N_1506,N_1941);
nand U2603 (N_2603,N_1791,N_1251);
nor U2604 (N_2604,N_1328,N_1081);
and U2605 (N_2605,N_1174,N_1647);
and U2606 (N_2606,N_1941,N_1960);
or U2607 (N_2607,N_1963,N_1680);
and U2608 (N_2608,N_1106,N_1256);
and U2609 (N_2609,N_1415,N_1617);
nor U2610 (N_2610,N_1844,N_1765);
nor U2611 (N_2611,N_1190,N_1857);
or U2612 (N_2612,N_1091,N_1673);
and U2613 (N_2613,N_1770,N_1213);
nand U2614 (N_2614,N_1703,N_1382);
nor U2615 (N_2615,N_1147,N_1244);
or U2616 (N_2616,N_1447,N_1048);
nor U2617 (N_2617,N_1400,N_1971);
and U2618 (N_2618,N_1633,N_1724);
nor U2619 (N_2619,N_1410,N_1199);
nor U2620 (N_2620,N_1277,N_1135);
and U2621 (N_2621,N_1647,N_1513);
and U2622 (N_2622,N_1653,N_1835);
nor U2623 (N_2623,N_1408,N_1829);
and U2624 (N_2624,N_1296,N_1433);
nand U2625 (N_2625,N_1062,N_1744);
or U2626 (N_2626,N_1272,N_1116);
nor U2627 (N_2627,N_1352,N_1750);
or U2628 (N_2628,N_1020,N_1806);
nand U2629 (N_2629,N_1762,N_1897);
nand U2630 (N_2630,N_1220,N_1751);
and U2631 (N_2631,N_1801,N_1472);
nor U2632 (N_2632,N_1832,N_1837);
nor U2633 (N_2633,N_1299,N_1521);
or U2634 (N_2634,N_1564,N_1039);
and U2635 (N_2635,N_1180,N_1516);
nand U2636 (N_2636,N_1632,N_1214);
nor U2637 (N_2637,N_1737,N_1405);
nand U2638 (N_2638,N_1372,N_1427);
or U2639 (N_2639,N_1189,N_1870);
nor U2640 (N_2640,N_1119,N_1199);
nand U2641 (N_2641,N_1349,N_1361);
or U2642 (N_2642,N_1147,N_1013);
nor U2643 (N_2643,N_1762,N_1448);
or U2644 (N_2644,N_1175,N_1585);
nor U2645 (N_2645,N_1927,N_1321);
nand U2646 (N_2646,N_1108,N_1615);
nor U2647 (N_2647,N_1284,N_1471);
nand U2648 (N_2648,N_1913,N_1153);
or U2649 (N_2649,N_1683,N_1105);
or U2650 (N_2650,N_1547,N_1691);
or U2651 (N_2651,N_1191,N_1011);
nor U2652 (N_2652,N_1591,N_1886);
or U2653 (N_2653,N_1743,N_1500);
nor U2654 (N_2654,N_1303,N_1052);
nor U2655 (N_2655,N_1948,N_1266);
nor U2656 (N_2656,N_1832,N_1247);
and U2657 (N_2657,N_1548,N_1067);
and U2658 (N_2658,N_1711,N_1998);
nor U2659 (N_2659,N_1293,N_1488);
and U2660 (N_2660,N_1744,N_1374);
nand U2661 (N_2661,N_1246,N_1687);
nand U2662 (N_2662,N_1796,N_1647);
nor U2663 (N_2663,N_1365,N_1401);
and U2664 (N_2664,N_1740,N_1725);
or U2665 (N_2665,N_1486,N_1184);
and U2666 (N_2666,N_1937,N_1399);
and U2667 (N_2667,N_1404,N_1864);
or U2668 (N_2668,N_1382,N_1491);
nor U2669 (N_2669,N_1335,N_1004);
nor U2670 (N_2670,N_1508,N_1283);
nor U2671 (N_2671,N_1312,N_1099);
nor U2672 (N_2672,N_1537,N_1098);
nor U2673 (N_2673,N_1457,N_1682);
nor U2674 (N_2674,N_1901,N_1055);
and U2675 (N_2675,N_1983,N_1524);
and U2676 (N_2676,N_1865,N_1290);
and U2677 (N_2677,N_1635,N_1216);
and U2678 (N_2678,N_1712,N_1685);
or U2679 (N_2679,N_1974,N_1200);
and U2680 (N_2680,N_1205,N_1273);
or U2681 (N_2681,N_1935,N_1114);
nand U2682 (N_2682,N_1216,N_1797);
or U2683 (N_2683,N_1594,N_1705);
nand U2684 (N_2684,N_1822,N_1500);
nor U2685 (N_2685,N_1740,N_1572);
nand U2686 (N_2686,N_1824,N_1640);
nor U2687 (N_2687,N_1448,N_1703);
nor U2688 (N_2688,N_1626,N_1805);
and U2689 (N_2689,N_1029,N_1276);
and U2690 (N_2690,N_1211,N_1486);
or U2691 (N_2691,N_1117,N_1049);
and U2692 (N_2692,N_1591,N_1517);
nand U2693 (N_2693,N_1101,N_1538);
and U2694 (N_2694,N_1128,N_1592);
and U2695 (N_2695,N_1560,N_1584);
or U2696 (N_2696,N_1236,N_1356);
or U2697 (N_2697,N_1494,N_1019);
and U2698 (N_2698,N_1729,N_1077);
nand U2699 (N_2699,N_1847,N_1522);
nor U2700 (N_2700,N_1338,N_1732);
or U2701 (N_2701,N_1615,N_1687);
and U2702 (N_2702,N_1168,N_1236);
nor U2703 (N_2703,N_1642,N_1610);
and U2704 (N_2704,N_1639,N_1175);
or U2705 (N_2705,N_1197,N_1631);
nand U2706 (N_2706,N_1919,N_1844);
and U2707 (N_2707,N_1281,N_1312);
and U2708 (N_2708,N_1566,N_1642);
nor U2709 (N_2709,N_1821,N_1018);
or U2710 (N_2710,N_1025,N_1674);
nor U2711 (N_2711,N_1319,N_1187);
or U2712 (N_2712,N_1842,N_1219);
nand U2713 (N_2713,N_1679,N_1052);
or U2714 (N_2714,N_1441,N_1254);
and U2715 (N_2715,N_1258,N_1075);
nand U2716 (N_2716,N_1619,N_1720);
nand U2717 (N_2717,N_1410,N_1112);
and U2718 (N_2718,N_1605,N_1157);
nand U2719 (N_2719,N_1437,N_1402);
or U2720 (N_2720,N_1629,N_1196);
or U2721 (N_2721,N_1723,N_1001);
nand U2722 (N_2722,N_1895,N_1168);
nor U2723 (N_2723,N_1819,N_1464);
nand U2724 (N_2724,N_1130,N_1941);
or U2725 (N_2725,N_1280,N_1166);
and U2726 (N_2726,N_1351,N_1882);
or U2727 (N_2727,N_1283,N_1660);
or U2728 (N_2728,N_1497,N_1401);
or U2729 (N_2729,N_1469,N_1348);
nand U2730 (N_2730,N_1051,N_1492);
nor U2731 (N_2731,N_1436,N_1114);
nor U2732 (N_2732,N_1076,N_1685);
or U2733 (N_2733,N_1851,N_1717);
or U2734 (N_2734,N_1514,N_1077);
or U2735 (N_2735,N_1078,N_1840);
nand U2736 (N_2736,N_1334,N_1242);
and U2737 (N_2737,N_1776,N_1645);
nand U2738 (N_2738,N_1081,N_1743);
nand U2739 (N_2739,N_1139,N_1451);
nand U2740 (N_2740,N_1748,N_1999);
or U2741 (N_2741,N_1619,N_1504);
nor U2742 (N_2742,N_1860,N_1258);
nand U2743 (N_2743,N_1849,N_1689);
nand U2744 (N_2744,N_1536,N_1892);
or U2745 (N_2745,N_1810,N_1867);
nand U2746 (N_2746,N_1607,N_1618);
or U2747 (N_2747,N_1462,N_1422);
and U2748 (N_2748,N_1273,N_1431);
and U2749 (N_2749,N_1449,N_1012);
nor U2750 (N_2750,N_1458,N_1951);
and U2751 (N_2751,N_1385,N_1067);
nand U2752 (N_2752,N_1118,N_1833);
nand U2753 (N_2753,N_1863,N_1905);
and U2754 (N_2754,N_1398,N_1312);
nand U2755 (N_2755,N_1647,N_1163);
nor U2756 (N_2756,N_1891,N_1602);
and U2757 (N_2757,N_1885,N_1191);
and U2758 (N_2758,N_1646,N_1949);
and U2759 (N_2759,N_1341,N_1138);
or U2760 (N_2760,N_1891,N_1925);
or U2761 (N_2761,N_1118,N_1839);
and U2762 (N_2762,N_1603,N_1616);
nor U2763 (N_2763,N_1852,N_1744);
nor U2764 (N_2764,N_1870,N_1638);
nand U2765 (N_2765,N_1851,N_1895);
or U2766 (N_2766,N_1900,N_1204);
nor U2767 (N_2767,N_1889,N_1532);
or U2768 (N_2768,N_1353,N_1260);
or U2769 (N_2769,N_1323,N_1012);
nand U2770 (N_2770,N_1787,N_1694);
or U2771 (N_2771,N_1772,N_1473);
nor U2772 (N_2772,N_1598,N_1720);
nand U2773 (N_2773,N_1578,N_1933);
and U2774 (N_2774,N_1716,N_1417);
nand U2775 (N_2775,N_1243,N_1308);
nor U2776 (N_2776,N_1201,N_1151);
or U2777 (N_2777,N_1084,N_1570);
nor U2778 (N_2778,N_1592,N_1538);
nand U2779 (N_2779,N_1103,N_1882);
or U2780 (N_2780,N_1184,N_1080);
and U2781 (N_2781,N_1153,N_1109);
or U2782 (N_2782,N_1859,N_1629);
nand U2783 (N_2783,N_1148,N_1217);
or U2784 (N_2784,N_1917,N_1156);
and U2785 (N_2785,N_1456,N_1092);
or U2786 (N_2786,N_1377,N_1670);
and U2787 (N_2787,N_1447,N_1965);
and U2788 (N_2788,N_1908,N_1208);
or U2789 (N_2789,N_1967,N_1512);
nand U2790 (N_2790,N_1425,N_1865);
nand U2791 (N_2791,N_1366,N_1431);
xor U2792 (N_2792,N_1794,N_1672);
and U2793 (N_2793,N_1583,N_1744);
nor U2794 (N_2794,N_1337,N_1258);
nor U2795 (N_2795,N_1211,N_1542);
and U2796 (N_2796,N_1300,N_1392);
nor U2797 (N_2797,N_1928,N_1535);
and U2798 (N_2798,N_1869,N_1751);
or U2799 (N_2799,N_1293,N_1500);
or U2800 (N_2800,N_1770,N_1623);
or U2801 (N_2801,N_1674,N_1657);
nand U2802 (N_2802,N_1758,N_1806);
xor U2803 (N_2803,N_1452,N_1428);
or U2804 (N_2804,N_1476,N_1783);
nor U2805 (N_2805,N_1592,N_1412);
or U2806 (N_2806,N_1133,N_1061);
and U2807 (N_2807,N_1587,N_1500);
nand U2808 (N_2808,N_1741,N_1596);
or U2809 (N_2809,N_1304,N_1615);
nor U2810 (N_2810,N_1072,N_1050);
or U2811 (N_2811,N_1916,N_1334);
or U2812 (N_2812,N_1743,N_1180);
or U2813 (N_2813,N_1812,N_1479);
nand U2814 (N_2814,N_1829,N_1848);
nor U2815 (N_2815,N_1544,N_1595);
or U2816 (N_2816,N_1914,N_1484);
nand U2817 (N_2817,N_1404,N_1893);
or U2818 (N_2818,N_1922,N_1475);
or U2819 (N_2819,N_1100,N_1454);
or U2820 (N_2820,N_1102,N_1999);
or U2821 (N_2821,N_1589,N_1528);
nand U2822 (N_2822,N_1484,N_1117);
nand U2823 (N_2823,N_1365,N_1318);
and U2824 (N_2824,N_1050,N_1427);
nand U2825 (N_2825,N_1290,N_1487);
or U2826 (N_2826,N_1768,N_1883);
and U2827 (N_2827,N_1824,N_1608);
and U2828 (N_2828,N_1964,N_1815);
nand U2829 (N_2829,N_1488,N_1314);
nor U2830 (N_2830,N_1504,N_1828);
or U2831 (N_2831,N_1064,N_1117);
nand U2832 (N_2832,N_1429,N_1995);
xnor U2833 (N_2833,N_1944,N_1574);
and U2834 (N_2834,N_1207,N_1133);
and U2835 (N_2835,N_1919,N_1143);
or U2836 (N_2836,N_1337,N_1722);
and U2837 (N_2837,N_1034,N_1322);
nor U2838 (N_2838,N_1745,N_1281);
and U2839 (N_2839,N_1469,N_1850);
nand U2840 (N_2840,N_1776,N_1893);
or U2841 (N_2841,N_1899,N_1598);
or U2842 (N_2842,N_1619,N_1652);
or U2843 (N_2843,N_1827,N_1957);
nor U2844 (N_2844,N_1407,N_1269);
nand U2845 (N_2845,N_1254,N_1276);
or U2846 (N_2846,N_1881,N_1542);
nand U2847 (N_2847,N_1734,N_1401);
nand U2848 (N_2848,N_1223,N_1035);
and U2849 (N_2849,N_1137,N_1548);
nor U2850 (N_2850,N_1630,N_1113);
nand U2851 (N_2851,N_1564,N_1270);
or U2852 (N_2852,N_1266,N_1722);
and U2853 (N_2853,N_1607,N_1143);
nor U2854 (N_2854,N_1479,N_1046);
nand U2855 (N_2855,N_1949,N_1684);
nand U2856 (N_2856,N_1357,N_1192);
nand U2857 (N_2857,N_1725,N_1414);
or U2858 (N_2858,N_1388,N_1227);
nor U2859 (N_2859,N_1163,N_1516);
nor U2860 (N_2860,N_1013,N_1004);
or U2861 (N_2861,N_1244,N_1853);
and U2862 (N_2862,N_1226,N_1299);
and U2863 (N_2863,N_1345,N_1749);
or U2864 (N_2864,N_1212,N_1318);
or U2865 (N_2865,N_1456,N_1337);
and U2866 (N_2866,N_1998,N_1029);
or U2867 (N_2867,N_1372,N_1522);
nand U2868 (N_2868,N_1073,N_1659);
nor U2869 (N_2869,N_1883,N_1454);
nor U2870 (N_2870,N_1872,N_1415);
nor U2871 (N_2871,N_1184,N_1522);
nor U2872 (N_2872,N_1070,N_1035);
nor U2873 (N_2873,N_1804,N_1117);
or U2874 (N_2874,N_1642,N_1753);
or U2875 (N_2875,N_1522,N_1040);
or U2876 (N_2876,N_1683,N_1435);
or U2877 (N_2877,N_1844,N_1523);
nand U2878 (N_2878,N_1855,N_1581);
or U2879 (N_2879,N_1277,N_1732);
or U2880 (N_2880,N_1975,N_1853);
or U2881 (N_2881,N_1046,N_1607);
nand U2882 (N_2882,N_1797,N_1523);
nand U2883 (N_2883,N_1717,N_1120);
xor U2884 (N_2884,N_1294,N_1507);
nand U2885 (N_2885,N_1264,N_1830);
nand U2886 (N_2886,N_1375,N_1610);
nor U2887 (N_2887,N_1166,N_1026);
nand U2888 (N_2888,N_1161,N_1845);
and U2889 (N_2889,N_1182,N_1133);
nand U2890 (N_2890,N_1271,N_1299);
nor U2891 (N_2891,N_1669,N_1019);
or U2892 (N_2892,N_1438,N_1545);
or U2893 (N_2893,N_1512,N_1076);
nand U2894 (N_2894,N_1742,N_1917);
or U2895 (N_2895,N_1030,N_1755);
nand U2896 (N_2896,N_1359,N_1368);
nand U2897 (N_2897,N_1235,N_1875);
nand U2898 (N_2898,N_1865,N_1112);
or U2899 (N_2899,N_1094,N_1789);
or U2900 (N_2900,N_1963,N_1231);
or U2901 (N_2901,N_1870,N_1635);
nor U2902 (N_2902,N_1419,N_1710);
or U2903 (N_2903,N_1643,N_1057);
nor U2904 (N_2904,N_1205,N_1063);
nand U2905 (N_2905,N_1334,N_1139);
and U2906 (N_2906,N_1094,N_1343);
or U2907 (N_2907,N_1449,N_1080);
nor U2908 (N_2908,N_1029,N_1721);
or U2909 (N_2909,N_1669,N_1821);
nor U2910 (N_2910,N_1187,N_1311);
nor U2911 (N_2911,N_1134,N_1909);
nand U2912 (N_2912,N_1397,N_1062);
nand U2913 (N_2913,N_1101,N_1543);
nor U2914 (N_2914,N_1171,N_1773);
and U2915 (N_2915,N_1015,N_1473);
and U2916 (N_2916,N_1266,N_1393);
nand U2917 (N_2917,N_1452,N_1925);
and U2918 (N_2918,N_1084,N_1891);
or U2919 (N_2919,N_1744,N_1836);
or U2920 (N_2920,N_1140,N_1113);
and U2921 (N_2921,N_1738,N_1392);
nor U2922 (N_2922,N_1190,N_1969);
or U2923 (N_2923,N_1128,N_1067);
nand U2924 (N_2924,N_1205,N_1610);
nor U2925 (N_2925,N_1500,N_1771);
nand U2926 (N_2926,N_1821,N_1535);
and U2927 (N_2927,N_1184,N_1929);
or U2928 (N_2928,N_1556,N_1945);
or U2929 (N_2929,N_1187,N_1033);
and U2930 (N_2930,N_1388,N_1885);
and U2931 (N_2931,N_1301,N_1921);
nor U2932 (N_2932,N_1301,N_1271);
nor U2933 (N_2933,N_1702,N_1398);
nor U2934 (N_2934,N_1544,N_1949);
nand U2935 (N_2935,N_1769,N_1474);
nand U2936 (N_2936,N_1572,N_1520);
or U2937 (N_2937,N_1940,N_1030);
and U2938 (N_2938,N_1584,N_1942);
or U2939 (N_2939,N_1619,N_1033);
nor U2940 (N_2940,N_1632,N_1768);
nand U2941 (N_2941,N_1534,N_1530);
nor U2942 (N_2942,N_1886,N_1226);
or U2943 (N_2943,N_1493,N_1985);
nand U2944 (N_2944,N_1076,N_1212);
nor U2945 (N_2945,N_1264,N_1488);
and U2946 (N_2946,N_1023,N_1244);
and U2947 (N_2947,N_1098,N_1337);
nand U2948 (N_2948,N_1727,N_1591);
nand U2949 (N_2949,N_1497,N_1576);
xnor U2950 (N_2950,N_1205,N_1973);
and U2951 (N_2951,N_1346,N_1624);
and U2952 (N_2952,N_1008,N_1687);
nand U2953 (N_2953,N_1220,N_1118);
nor U2954 (N_2954,N_1977,N_1507);
nand U2955 (N_2955,N_1064,N_1426);
and U2956 (N_2956,N_1251,N_1022);
nand U2957 (N_2957,N_1822,N_1180);
nand U2958 (N_2958,N_1356,N_1859);
and U2959 (N_2959,N_1979,N_1457);
nand U2960 (N_2960,N_1690,N_1293);
and U2961 (N_2961,N_1611,N_1565);
or U2962 (N_2962,N_1402,N_1225);
or U2963 (N_2963,N_1034,N_1677);
nor U2964 (N_2964,N_1065,N_1356);
or U2965 (N_2965,N_1805,N_1284);
and U2966 (N_2966,N_1107,N_1407);
nand U2967 (N_2967,N_1676,N_1536);
and U2968 (N_2968,N_1753,N_1646);
nand U2969 (N_2969,N_1153,N_1589);
nand U2970 (N_2970,N_1824,N_1436);
and U2971 (N_2971,N_1970,N_1523);
or U2972 (N_2972,N_1280,N_1241);
nand U2973 (N_2973,N_1935,N_1269);
or U2974 (N_2974,N_1542,N_1152);
nor U2975 (N_2975,N_1662,N_1694);
nand U2976 (N_2976,N_1675,N_1563);
nor U2977 (N_2977,N_1486,N_1031);
and U2978 (N_2978,N_1040,N_1067);
or U2979 (N_2979,N_1193,N_1588);
nor U2980 (N_2980,N_1791,N_1525);
nor U2981 (N_2981,N_1145,N_1211);
and U2982 (N_2982,N_1281,N_1344);
or U2983 (N_2983,N_1887,N_1168);
nand U2984 (N_2984,N_1551,N_1791);
and U2985 (N_2985,N_1397,N_1345);
and U2986 (N_2986,N_1492,N_1217);
nand U2987 (N_2987,N_1138,N_1133);
and U2988 (N_2988,N_1818,N_1595);
and U2989 (N_2989,N_1403,N_1002);
and U2990 (N_2990,N_1634,N_1763);
nor U2991 (N_2991,N_1143,N_1777);
nor U2992 (N_2992,N_1944,N_1126);
or U2993 (N_2993,N_1235,N_1534);
and U2994 (N_2994,N_1075,N_1995);
or U2995 (N_2995,N_1330,N_1402);
and U2996 (N_2996,N_1743,N_1537);
nor U2997 (N_2997,N_1087,N_1343);
or U2998 (N_2998,N_1767,N_1756);
nand U2999 (N_2999,N_1218,N_1448);
or U3000 (N_3000,N_2455,N_2750);
or U3001 (N_3001,N_2766,N_2183);
and U3002 (N_3002,N_2491,N_2617);
and U3003 (N_3003,N_2136,N_2020);
or U3004 (N_3004,N_2948,N_2248);
nand U3005 (N_3005,N_2919,N_2632);
nand U3006 (N_3006,N_2857,N_2936);
and U3007 (N_3007,N_2541,N_2992);
nand U3008 (N_3008,N_2159,N_2745);
nand U3009 (N_3009,N_2611,N_2677);
and U3010 (N_3010,N_2037,N_2889);
nand U3011 (N_3011,N_2079,N_2867);
nand U3012 (N_3012,N_2916,N_2363);
or U3013 (N_3013,N_2732,N_2240);
and U3014 (N_3014,N_2585,N_2430);
nand U3015 (N_3015,N_2127,N_2665);
or U3016 (N_3016,N_2711,N_2760);
nor U3017 (N_3017,N_2154,N_2879);
nor U3018 (N_3018,N_2554,N_2881);
nand U3019 (N_3019,N_2534,N_2326);
or U3020 (N_3020,N_2654,N_2525);
and U3021 (N_3021,N_2775,N_2187);
nor U3022 (N_3022,N_2519,N_2771);
nor U3023 (N_3023,N_2122,N_2048);
or U3024 (N_3024,N_2040,N_2494);
or U3025 (N_3025,N_2006,N_2345);
nand U3026 (N_3026,N_2113,N_2241);
or U3027 (N_3027,N_2421,N_2153);
and U3028 (N_3028,N_2313,N_2818);
and U3029 (N_3029,N_2386,N_2353);
nand U3030 (N_3030,N_2662,N_2317);
nor U3031 (N_3031,N_2956,N_2843);
and U3032 (N_3032,N_2655,N_2747);
nand U3033 (N_3033,N_2223,N_2328);
nand U3034 (N_3034,N_2870,N_2644);
and U3035 (N_3035,N_2651,N_2939);
and U3036 (N_3036,N_2613,N_2781);
and U3037 (N_3037,N_2051,N_2476);
and U3038 (N_3038,N_2957,N_2266);
nand U3039 (N_3039,N_2707,N_2892);
and U3040 (N_3040,N_2675,N_2145);
xnor U3041 (N_3041,N_2167,N_2319);
or U3042 (N_3042,N_2549,N_2720);
nor U3043 (N_3043,N_2635,N_2898);
and U3044 (N_3044,N_2514,N_2575);
or U3045 (N_3045,N_2785,N_2774);
and U3046 (N_3046,N_2242,N_2931);
or U3047 (N_3047,N_2161,N_2038);
nor U3048 (N_3048,N_2503,N_2551);
nand U3049 (N_3049,N_2042,N_2681);
nor U3050 (N_3050,N_2715,N_2214);
nor U3051 (N_3051,N_2335,N_2330);
xnor U3052 (N_3052,N_2704,N_2258);
nand U3053 (N_3053,N_2521,N_2464);
nand U3054 (N_3054,N_2171,N_2088);
and U3055 (N_3055,N_2095,N_2587);
xor U3056 (N_3056,N_2960,N_2373);
or U3057 (N_3057,N_2968,N_2988);
nand U3058 (N_3058,N_2433,N_2907);
nand U3059 (N_3059,N_2542,N_2506);
xor U3060 (N_3060,N_2350,N_2828);
nor U3061 (N_3061,N_2914,N_2264);
xor U3062 (N_3062,N_2190,N_2897);
or U3063 (N_3063,N_2492,N_2984);
nor U3064 (N_3064,N_2454,N_2073);
and U3065 (N_3065,N_2388,N_2513);
or U3066 (N_3066,N_2323,N_2558);
or U3067 (N_3067,N_2010,N_2666);
or U3068 (N_3068,N_2678,N_2544);
and U3069 (N_3069,N_2356,N_2761);
nor U3070 (N_3070,N_2652,N_2201);
or U3071 (N_3071,N_2653,N_2926);
or U3072 (N_3072,N_2007,N_2615);
or U3073 (N_3073,N_2823,N_2083);
nor U3074 (N_3074,N_2583,N_2450);
nand U3075 (N_3075,N_2708,N_2200);
nor U3076 (N_3076,N_2794,N_2250);
and U3077 (N_3077,N_2211,N_2697);
nand U3078 (N_3078,N_2486,N_2366);
and U3079 (N_3079,N_2289,N_2780);
nor U3080 (N_3080,N_2305,N_2825);
and U3081 (N_3081,N_2621,N_2231);
nand U3082 (N_3082,N_2118,N_2199);
or U3083 (N_3083,N_2149,N_2605);
or U3084 (N_3084,N_2121,N_2470);
nand U3085 (N_3085,N_2721,N_2508);
nand U3086 (N_3086,N_2495,N_2379);
nand U3087 (N_3087,N_2923,N_2813);
and U3088 (N_3088,N_2302,N_2772);
nor U3089 (N_3089,N_2821,N_2873);
nand U3090 (N_3090,N_2413,N_2237);
nor U3091 (N_3091,N_2983,N_2216);
nand U3092 (N_3092,N_2212,N_2487);
nor U3093 (N_3093,N_2570,N_2927);
or U3094 (N_3094,N_2535,N_2522);
and U3095 (N_3095,N_2723,N_2259);
and U3096 (N_3096,N_2973,N_2279);
nor U3097 (N_3097,N_2036,N_2620);
nand U3098 (N_3098,N_2315,N_2303);
xnor U3099 (N_3099,N_2185,N_2922);
nand U3100 (N_3100,N_2601,N_2424);
or U3101 (N_3101,N_2880,N_2545);
or U3102 (N_3102,N_2878,N_2298);
or U3103 (N_3103,N_2148,N_2947);
nor U3104 (N_3104,N_2093,N_2844);
nor U3105 (N_3105,N_2102,N_2540);
nand U3106 (N_3106,N_2504,N_2206);
and U3107 (N_3107,N_2905,N_2566);
nand U3108 (N_3108,N_2461,N_2217);
and U3109 (N_3109,N_2204,N_2233);
nor U3110 (N_3110,N_2589,N_2033);
nand U3111 (N_3111,N_2378,N_2719);
or U3112 (N_3112,N_2131,N_2105);
nand U3113 (N_3113,N_2238,N_2740);
or U3114 (N_3114,N_2229,N_2657);
nor U3115 (N_3115,N_2584,N_2107);
or U3116 (N_3116,N_2498,N_2032);
or U3117 (N_3117,N_2137,N_2580);
nand U3118 (N_3118,N_2224,N_2727);
nand U3119 (N_3119,N_2372,N_2468);
and U3120 (N_3120,N_2518,N_2307);
nand U3121 (N_3121,N_2225,N_2273);
and U3122 (N_3122,N_2855,N_2427);
and U3123 (N_3123,N_2432,N_2344);
or U3124 (N_3124,N_2827,N_2256);
nand U3125 (N_3125,N_2269,N_2779);
nor U3126 (N_3126,N_2529,N_2493);
and U3127 (N_3127,N_2816,N_2451);
and U3128 (N_3128,N_2932,N_2092);
nor U3129 (N_3129,N_2067,N_2347);
nand U3130 (N_3130,N_2861,N_2702);
nor U3131 (N_3131,N_2547,N_2556);
nand U3132 (N_3132,N_2967,N_2146);
xnor U3133 (N_3133,N_2714,N_2478);
or U3134 (N_3134,N_2483,N_2218);
and U3135 (N_3135,N_2375,N_2458);
or U3136 (N_3136,N_2381,N_2044);
nor U3137 (N_3137,N_2890,N_2985);
and U3138 (N_3138,N_2725,N_2467);
and U3139 (N_3139,N_2756,N_2520);
nor U3140 (N_3140,N_2981,N_2955);
nand U3141 (N_3141,N_2156,N_2342);
nor U3142 (N_3142,N_2791,N_2596);
and U3143 (N_3143,N_2134,N_2025);
and U3144 (N_3144,N_2884,N_2619);
nand U3145 (N_3145,N_2856,N_2862);
or U3146 (N_3146,N_2096,N_2920);
nand U3147 (N_3147,N_2784,N_2724);
or U3148 (N_3148,N_2417,N_2624);
nand U3149 (N_3149,N_2263,N_2429);
or U3150 (N_3150,N_2663,N_2274);
nand U3151 (N_3151,N_2989,N_2143);
xnor U3152 (N_3152,N_2202,N_2604);
nor U3153 (N_3153,N_2471,N_2921);
nand U3154 (N_3154,N_2374,N_2236);
nand U3155 (N_3155,N_2453,N_2959);
nor U3156 (N_3156,N_2360,N_2933);
nand U3157 (N_3157,N_2752,N_2170);
and U3158 (N_3158,N_2295,N_2163);
nand U3159 (N_3159,N_2835,N_2401);
nor U3160 (N_3160,N_2845,N_2557);
or U3161 (N_3161,N_2247,N_2160);
and U3162 (N_3162,N_2022,N_2035);
xor U3163 (N_3163,N_2490,N_2533);
nor U3164 (N_3164,N_2408,N_2626);
nand U3165 (N_3165,N_2184,N_2996);
or U3166 (N_3166,N_2039,N_2966);
and U3167 (N_3167,N_2050,N_2339);
and U3168 (N_3168,N_2232,N_2368);
nor U3169 (N_3169,N_2338,N_2552);
nand U3170 (N_3170,N_2078,N_2918);
and U3171 (N_3171,N_2405,N_2400);
or U3172 (N_3172,N_2700,N_2997);
nand U3173 (N_3173,N_2803,N_2142);
nor U3174 (N_3174,N_2327,N_2592);
or U3175 (N_3175,N_2402,N_2442);
nor U3176 (N_3176,N_2348,N_2423);
and U3177 (N_3177,N_2380,N_2838);
and U3178 (N_3178,N_2883,N_2003);
and U3179 (N_3179,N_2833,N_2778);
nand U3180 (N_3180,N_2768,N_2412);
nor U3181 (N_3181,N_2999,N_2151);
nand U3182 (N_3182,N_2925,N_2071);
or U3183 (N_3183,N_2625,N_2910);
nor U3184 (N_3184,N_2638,N_2516);
nand U3185 (N_3185,N_2851,N_2895);
or U3186 (N_3186,N_2640,N_2893);
or U3187 (N_3187,N_2452,N_2527);
and U3188 (N_3188,N_2840,N_2972);
or U3189 (N_3189,N_2776,N_2497);
or U3190 (N_3190,N_2139,N_2019);
nor U3191 (N_3191,N_2859,N_2087);
nor U3192 (N_3192,N_2062,N_2986);
nand U3193 (N_3193,N_2832,N_2739);
nor U3194 (N_3194,N_2065,N_2913);
nor U3195 (N_3195,N_2964,N_2868);
nand U3196 (N_3196,N_2562,N_2712);
nor U3197 (N_3197,N_2684,N_2963);
nand U3198 (N_3198,N_2735,N_2125);
nor U3199 (N_3199,N_2124,N_2710);
nor U3200 (N_3200,N_2705,N_2786);
and U3201 (N_3201,N_2479,N_2757);
xnor U3202 (N_3202,N_2100,N_2063);
nand U3203 (N_3203,N_2055,N_2773);
or U3204 (N_3204,N_2270,N_2299);
and U3205 (N_3205,N_2239,N_2882);
or U3206 (N_3206,N_2340,N_2060);
or U3207 (N_3207,N_2709,N_2568);
nor U3208 (N_3208,N_2886,N_2915);
xnor U3209 (N_3209,N_2523,N_2646);
nand U3210 (N_3210,N_2296,N_2829);
nor U3211 (N_3211,N_2627,N_2449);
and U3212 (N_3212,N_2788,N_2826);
and U3213 (N_3213,N_2945,N_2538);
nand U3214 (N_3214,N_2369,N_2642);
nand U3215 (N_3215,N_2616,N_2436);
nand U3216 (N_3216,N_2607,N_2061);
and U3217 (N_3217,N_2045,N_2820);
nand U3218 (N_3218,N_2252,N_2517);
nor U3219 (N_3219,N_2446,N_2852);
or U3220 (N_3220,N_2942,N_2397);
nor U3221 (N_3221,N_2352,N_2106);
nor U3222 (N_3222,N_2563,N_2489);
or U3223 (N_3223,N_2324,N_2482);
nand U3224 (N_3224,N_2731,N_2415);
or U3225 (N_3225,N_2481,N_2165);
xnor U3226 (N_3226,N_2166,N_2016);
nand U3227 (N_3227,N_2441,N_2975);
or U3228 (N_3228,N_2909,N_2245);
or U3229 (N_3229,N_2126,N_2026);
nand U3230 (N_3230,N_2135,N_2116);
or U3231 (N_3231,N_2080,N_2853);
and U3232 (N_3232,N_2046,N_2311);
nor U3233 (N_3233,N_2089,N_2722);
nor U3234 (N_3234,N_2977,N_2462);
or U3235 (N_3235,N_2141,N_2950);
or U3236 (N_3236,N_2849,N_2595);
or U3237 (N_3237,N_2590,N_2532);
or U3238 (N_3238,N_2800,N_2431);
nand U3239 (N_3239,N_2755,N_2656);
nor U3240 (N_3240,N_2696,N_2475);
and U3241 (N_3241,N_2935,N_2178);
nor U3242 (N_3242,N_2537,N_2924);
or U3243 (N_3243,N_2811,N_2633);
nand U3244 (N_3244,N_2894,N_2075);
nor U3245 (N_3245,N_2804,N_2460);
nor U3246 (N_3246,N_2070,N_2112);
or U3247 (N_3247,N_2014,N_2002);
nand U3248 (N_3248,N_2047,N_2104);
or U3249 (N_3249,N_2896,N_2701);
nand U3250 (N_3250,N_2426,N_2349);
or U3251 (N_3251,N_2140,N_2569);
nor U3252 (N_3252,N_2359,N_2748);
or U3253 (N_3253,N_2371,N_2255);
nor U3254 (N_3254,N_2974,N_2243);
or U3255 (N_3255,N_2117,N_2208);
and U3256 (N_3256,N_2608,N_2797);
nor U3257 (N_3257,N_2980,N_2249);
or U3258 (N_3258,N_2673,N_2744);
xor U3259 (N_3259,N_2157,N_2180);
nand U3260 (N_3260,N_2703,N_2694);
or U3261 (N_3261,N_2899,N_2439);
nor U3262 (N_3262,N_2235,N_2993);
nor U3263 (N_3263,N_2539,N_2734);
and U3264 (N_3264,N_2824,N_2012);
nor U3265 (N_3265,N_2336,N_2836);
or U3266 (N_3266,N_2565,N_2597);
and U3267 (N_3267,N_2129,N_2480);
nor U3268 (N_3268,N_2337,N_2174);
and U3269 (N_3269,N_2422,N_2034);
nor U3270 (N_3270,N_2689,N_2354);
and U3271 (N_3271,N_2409,N_2741);
and U3272 (N_3272,N_2888,N_2528);
and U3273 (N_3273,N_2636,N_2777);
nor U3274 (N_3274,N_2680,N_2995);
nor U3275 (N_3275,N_2837,N_2682);
nor U3276 (N_3276,N_2819,N_2929);
nor U3277 (N_3277,N_2253,N_2874);
and U3278 (N_3278,N_2792,N_2280);
nor U3279 (N_3279,N_2941,N_2979);
nor U3280 (N_3280,N_2806,N_2622);
and U3281 (N_3281,N_2599,N_2282);
and U3282 (N_3282,N_2500,N_2130);
and U3283 (N_3283,N_2579,N_2706);
nand U3284 (N_3284,N_2809,N_2013);
or U3285 (N_3285,N_2937,N_2394);
or U3286 (N_3286,N_2396,N_2733);
and U3287 (N_3287,N_2283,N_2091);
and U3288 (N_3288,N_2203,N_2086);
nand U3289 (N_3289,N_2419,N_2262);
xnor U3290 (N_3290,N_2603,N_2692);
or U3291 (N_3291,N_2132,N_2138);
nor U3292 (N_3292,N_2227,N_2290);
nand U3293 (N_3293,N_2284,N_2213);
nor U3294 (N_3294,N_2854,N_2383);
nand U3295 (N_3295,N_2182,N_2501);
nor U3296 (N_3296,N_2660,N_2376);
nand U3297 (N_3297,N_2278,N_2331);
or U3298 (N_3298,N_2390,N_2195);
or U3299 (N_3299,N_2841,N_2275);
nor U3300 (N_3300,N_2384,N_2578);
nand U3301 (N_3301,N_2312,N_2054);
and U3302 (N_3302,N_2272,N_2787);
and U3303 (N_3303,N_2728,N_2457);
and U3304 (N_3304,N_2308,N_2094);
and U3305 (N_3305,N_2215,N_2097);
nor U3306 (N_3306,N_2940,N_2567);
or U3307 (N_3307,N_2737,N_2164);
nand U3308 (N_3308,N_2023,N_2645);
and U3309 (N_3309,N_2978,N_2699);
and U3310 (N_3310,N_2128,N_2749);
or U3311 (N_3311,N_2260,N_2234);
and U3312 (N_3312,N_2875,N_2021);
nand U3313 (N_3313,N_2526,N_2300);
or U3314 (N_3314,N_2763,N_2198);
nand U3315 (N_3315,N_2944,N_2316);
nand U3316 (N_3316,N_2512,N_2355);
nor U3317 (N_3317,N_2553,N_2357);
and U3318 (N_3318,N_2414,N_2524);
nand U3319 (N_3319,N_2018,N_2648);
nand U3320 (N_3320,N_2814,N_2586);
nor U3321 (N_3321,N_2364,N_2971);
nand U3322 (N_3322,N_2000,N_2609);
nor U3323 (N_3323,N_2158,N_2435);
and U3324 (N_3324,N_2459,N_2812);
nand U3325 (N_3325,N_2110,N_2325);
nor U3326 (N_3326,N_2210,N_2795);
and U3327 (N_3327,N_2762,N_2865);
and U3328 (N_3328,N_2465,N_2954);
nor U3329 (N_3329,N_2005,N_2332);
and U3330 (N_3330,N_2885,N_2822);
or U3331 (N_3331,N_2004,N_2848);
nor U3332 (N_3332,N_2056,N_2420);
and U3333 (N_3333,N_2277,N_2286);
and U3334 (N_3334,N_2858,N_2186);
or U3335 (N_3335,N_2103,N_2831);
nand U3336 (N_3336,N_2686,N_2976);
or U3337 (N_3337,N_2962,N_2389);
or U3338 (N_3338,N_2869,N_2998);
nand U3339 (N_3339,N_2428,N_2798);
and U3340 (N_3340,N_2434,N_2120);
nand U3341 (N_3341,N_2769,N_2098);
nand U3342 (N_3342,N_2416,N_2515);
and U3343 (N_3343,N_2292,N_2181);
nor U3344 (N_3344,N_2499,N_2850);
nand U3345 (N_3345,N_2310,N_2293);
nand U3346 (N_3346,N_2011,N_2099);
nand U3347 (N_3347,N_2801,N_2082);
and U3348 (N_3348,N_2674,N_2876);
nor U3349 (N_3349,N_2267,N_2030);
nand U3350 (N_3350,N_2230,N_2438);
and U3351 (N_3351,N_2029,N_2555);
and U3352 (N_3352,N_2630,N_2069);
nor U3353 (N_3353,N_2144,N_2982);
nand U3354 (N_3354,N_2226,N_2268);
nand U3355 (N_3355,N_2334,N_2008);
nand U3356 (N_3356,N_2698,N_2805);
or U3357 (N_3357,N_2447,N_2934);
nand U3358 (N_3358,N_2842,N_2866);
nand U3359 (N_3359,N_2015,N_2770);
nand U3360 (N_3360,N_2802,N_2437);
nand U3361 (N_3361,N_2891,N_2990);
or U3362 (N_3362,N_2509,N_2536);
or U3363 (N_3363,N_2690,N_2953);
nor U3364 (N_3364,N_2343,N_2058);
nand U3365 (N_3365,N_2864,N_2188);
and U3366 (N_3366,N_2254,N_2670);
nand U3367 (N_3367,N_2602,N_2411);
and U3368 (N_3368,N_2175,N_2507);
and U3369 (N_3369,N_2001,N_2904);
or U3370 (N_3370,N_2228,N_2691);
or U3371 (N_3371,N_2564,N_2716);
nor U3372 (N_3372,N_2387,N_2901);
or U3373 (N_3373,N_2606,N_2028);
and U3374 (N_3374,N_2759,N_2367);
nand U3375 (N_3375,N_2077,N_2115);
nor U3376 (N_3376,N_2808,N_2176);
or U3377 (N_3377,N_2543,N_2938);
nor U3378 (N_3378,N_2560,N_2629);
and U3379 (N_3379,N_2903,N_2659);
nor U3380 (N_3380,N_2729,N_2758);
or U3381 (N_3381,N_2320,N_2318);
and U3382 (N_3382,N_2685,N_2614);
or U3383 (N_3383,N_2197,N_2637);
and U3384 (N_3384,N_2911,N_2746);
nand U3385 (N_3385,N_2783,N_2949);
nand U3386 (N_3386,N_2810,N_2991);
and U3387 (N_3387,N_2610,N_2577);
nor U3388 (N_3388,N_2031,N_2649);
nand U3389 (N_3389,N_2123,N_2496);
nor U3390 (N_3390,N_2650,N_2111);
and U3391 (N_3391,N_2246,N_2908);
xor U3392 (N_3392,N_2561,N_2177);
nand U3393 (N_3393,N_2790,N_2582);
and U3394 (N_3394,N_2667,N_2057);
and U3395 (N_3395,N_2322,N_2477);
nand U3396 (N_3396,N_2017,N_2598);
nand U3397 (N_3397,N_2287,N_2191);
and U3398 (N_3398,N_2398,N_2754);
nand U3399 (N_3399,N_2251,N_2189);
and U3400 (N_3400,N_2119,N_2072);
nand U3401 (N_3401,N_2133,N_2168);
nand U3402 (N_3402,N_2505,N_2391);
or U3403 (N_3403,N_2846,N_2930);
nand U3404 (N_3404,N_2839,N_2917);
and U3405 (N_3405,N_2546,N_2987);
or U3406 (N_3406,N_2162,N_2618);
or U3407 (N_3407,N_2679,N_2049);
nand U3408 (N_3408,N_2362,N_2341);
nand U3409 (N_3409,N_2473,N_2333);
and U3410 (N_3410,N_2445,N_2297);
nor U3411 (N_3411,N_2346,N_2695);
and U3412 (N_3412,N_2764,N_2736);
nor U3413 (N_3413,N_2726,N_2643);
nand U3414 (N_3414,N_2713,N_2571);
nand U3415 (N_3415,N_2150,N_2193);
nand U3416 (N_3416,N_2510,N_2329);
or U3417 (N_3417,N_2594,N_2257);
or U3418 (N_3418,N_2672,N_2600);
or U3419 (N_3419,N_2573,N_2753);
nand U3420 (N_3420,N_2076,N_2782);
or U3421 (N_3421,N_2834,N_2052);
nor U3422 (N_3422,N_2219,N_2276);
xor U3423 (N_3423,N_2074,N_2472);
and U3424 (N_3424,N_2730,N_2906);
nand U3425 (N_3425,N_2502,N_2053);
or U3426 (N_3426,N_2817,N_2403);
nor U3427 (N_3427,N_2304,N_2365);
or U3428 (N_3428,N_2623,N_2440);
nand U3429 (N_3429,N_2550,N_2309);
and U3430 (N_3430,N_2912,N_2951);
nor U3431 (N_3431,N_2294,N_2265);
and U3432 (N_3432,N_2418,N_2474);
nand U3433 (N_3433,N_2043,N_2155);
and U3434 (N_3434,N_2404,N_2220);
or U3435 (N_3435,N_2576,N_2172);
nand U3436 (N_3436,N_2109,N_2410);
and U3437 (N_3437,N_2676,N_2877);
nand U3438 (N_3438,N_2064,N_2207);
nor U3439 (N_3439,N_2205,N_2738);
nor U3440 (N_3440,N_2024,N_2658);
or U3441 (N_3441,N_2081,N_2593);
and U3442 (N_3442,N_2668,N_2306);
or U3443 (N_3443,N_2169,N_2793);
nor U3444 (N_3444,N_2382,N_2221);
nor U3445 (N_3445,N_2271,N_2634);
xnor U3446 (N_3446,N_2196,N_2488);
nand U3447 (N_3447,N_2946,N_2301);
nor U3448 (N_3448,N_2399,N_2574);
and U3449 (N_3449,N_2612,N_2009);
nand U3450 (N_3450,N_2084,N_2377);
or U3451 (N_3451,N_2194,N_2392);
or U3452 (N_3452,N_2358,N_2108);
nor U3453 (N_3453,N_2661,N_2443);
nand U3454 (N_3454,N_2291,N_2530);
or U3455 (N_3455,N_2173,N_2059);
nand U3456 (N_3456,N_2407,N_2041);
and U3457 (N_3457,N_2799,N_2965);
nand U3458 (N_3458,N_2531,N_2321);
nor U3459 (N_3459,N_2222,N_2994);
or U3460 (N_3460,N_2969,N_2872);
nor U3461 (N_3461,N_2209,N_2484);
nand U3462 (N_3462,N_2385,N_2639);
or U3463 (N_3463,N_2900,N_2815);
and U3464 (N_3464,N_2244,N_2581);
or U3465 (N_3465,N_2559,N_2485);
or U3466 (N_3466,N_2147,N_2928);
or U3467 (N_3467,N_2669,N_2027);
nor U3468 (N_3468,N_2847,N_2902);
nor U3469 (N_3469,N_2469,N_2830);
or U3470 (N_3470,N_2463,N_2631);
nand U3471 (N_3471,N_2285,N_2742);
and U3472 (N_3472,N_2370,N_2863);
nor U3473 (N_3473,N_2693,N_2288);
or U3474 (N_3474,N_2628,N_2683);
or U3475 (N_3475,N_2548,N_2511);
nand U3476 (N_3476,N_2085,N_2393);
or U3477 (N_3477,N_2743,N_2572);
nor U3478 (N_3478,N_2466,N_2361);
and U3479 (N_3479,N_2068,N_2192);
nand U3480 (N_3480,N_2887,N_2688);
nor U3481 (N_3481,N_2351,N_2395);
or U3482 (N_3482,N_2718,N_2871);
or U3483 (N_3483,N_2958,N_2456);
nand U3484 (N_3484,N_2767,N_2591);
and U3485 (N_3485,N_2641,N_2114);
nand U3486 (N_3486,N_2647,N_2860);
nand U3487 (N_3487,N_2425,N_2152);
or U3488 (N_3488,N_2066,N_2588);
and U3489 (N_3489,N_2807,N_2687);
nand U3490 (N_3490,N_2952,N_2961);
or U3491 (N_3491,N_2717,N_2970);
and U3492 (N_3492,N_2444,N_2179);
nor U3493 (N_3493,N_2751,N_2090);
and U3494 (N_3494,N_2664,N_2671);
or U3495 (N_3495,N_2314,N_2261);
and U3496 (N_3496,N_2789,N_2281);
nor U3497 (N_3497,N_2406,N_2101);
nand U3498 (N_3498,N_2796,N_2765);
and U3499 (N_3499,N_2448,N_2943);
and U3500 (N_3500,N_2386,N_2159);
or U3501 (N_3501,N_2521,N_2182);
nor U3502 (N_3502,N_2051,N_2594);
and U3503 (N_3503,N_2425,N_2361);
nor U3504 (N_3504,N_2824,N_2223);
and U3505 (N_3505,N_2174,N_2651);
and U3506 (N_3506,N_2268,N_2886);
nor U3507 (N_3507,N_2443,N_2795);
nand U3508 (N_3508,N_2768,N_2242);
nand U3509 (N_3509,N_2565,N_2846);
and U3510 (N_3510,N_2030,N_2593);
nor U3511 (N_3511,N_2630,N_2048);
and U3512 (N_3512,N_2047,N_2103);
and U3513 (N_3513,N_2190,N_2655);
and U3514 (N_3514,N_2902,N_2590);
nand U3515 (N_3515,N_2785,N_2878);
or U3516 (N_3516,N_2796,N_2520);
and U3517 (N_3517,N_2059,N_2455);
nand U3518 (N_3518,N_2975,N_2480);
nand U3519 (N_3519,N_2630,N_2029);
xor U3520 (N_3520,N_2059,N_2065);
nor U3521 (N_3521,N_2478,N_2047);
nand U3522 (N_3522,N_2839,N_2727);
or U3523 (N_3523,N_2633,N_2650);
or U3524 (N_3524,N_2884,N_2038);
and U3525 (N_3525,N_2155,N_2125);
and U3526 (N_3526,N_2037,N_2969);
or U3527 (N_3527,N_2650,N_2140);
nand U3528 (N_3528,N_2076,N_2110);
and U3529 (N_3529,N_2574,N_2248);
and U3530 (N_3530,N_2207,N_2078);
or U3531 (N_3531,N_2746,N_2382);
nand U3532 (N_3532,N_2597,N_2070);
nand U3533 (N_3533,N_2173,N_2409);
and U3534 (N_3534,N_2331,N_2463);
nand U3535 (N_3535,N_2064,N_2617);
and U3536 (N_3536,N_2771,N_2138);
nand U3537 (N_3537,N_2956,N_2688);
nor U3538 (N_3538,N_2170,N_2814);
nand U3539 (N_3539,N_2323,N_2532);
and U3540 (N_3540,N_2889,N_2749);
nand U3541 (N_3541,N_2580,N_2312);
nand U3542 (N_3542,N_2798,N_2427);
or U3543 (N_3543,N_2645,N_2072);
or U3544 (N_3544,N_2808,N_2241);
or U3545 (N_3545,N_2755,N_2440);
or U3546 (N_3546,N_2493,N_2343);
or U3547 (N_3547,N_2557,N_2844);
and U3548 (N_3548,N_2190,N_2769);
and U3549 (N_3549,N_2420,N_2116);
and U3550 (N_3550,N_2978,N_2802);
nor U3551 (N_3551,N_2375,N_2847);
and U3552 (N_3552,N_2355,N_2170);
or U3553 (N_3553,N_2411,N_2321);
nor U3554 (N_3554,N_2605,N_2137);
and U3555 (N_3555,N_2247,N_2421);
nor U3556 (N_3556,N_2924,N_2714);
or U3557 (N_3557,N_2153,N_2619);
nand U3558 (N_3558,N_2297,N_2244);
nor U3559 (N_3559,N_2087,N_2890);
or U3560 (N_3560,N_2298,N_2421);
nand U3561 (N_3561,N_2276,N_2490);
nor U3562 (N_3562,N_2990,N_2122);
nor U3563 (N_3563,N_2290,N_2623);
nand U3564 (N_3564,N_2088,N_2167);
nand U3565 (N_3565,N_2405,N_2106);
nand U3566 (N_3566,N_2714,N_2705);
or U3567 (N_3567,N_2239,N_2401);
nor U3568 (N_3568,N_2299,N_2665);
and U3569 (N_3569,N_2759,N_2632);
nor U3570 (N_3570,N_2788,N_2479);
or U3571 (N_3571,N_2896,N_2717);
xor U3572 (N_3572,N_2438,N_2016);
and U3573 (N_3573,N_2117,N_2417);
nand U3574 (N_3574,N_2408,N_2766);
or U3575 (N_3575,N_2123,N_2250);
and U3576 (N_3576,N_2682,N_2581);
nand U3577 (N_3577,N_2288,N_2965);
or U3578 (N_3578,N_2150,N_2924);
nor U3579 (N_3579,N_2900,N_2185);
or U3580 (N_3580,N_2891,N_2010);
nand U3581 (N_3581,N_2941,N_2899);
or U3582 (N_3582,N_2301,N_2571);
nor U3583 (N_3583,N_2385,N_2766);
or U3584 (N_3584,N_2811,N_2037);
nor U3585 (N_3585,N_2124,N_2433);
and U3586 (N_3586,N_2715,N_2917);
or U3587 (N_3587,N_2265,N_2565);
or U3588 (N_3588,N_2555,N_2799);
nor U3589 (N_3589,N_2534,N_2092);
or U3590 (N_3590,N_2742,N_2736);
or U3591 (N_3591,N_2455,N_2598);
nor U3592 (N_3592,N_2505,N_2342);
nor U3593 (N_3593,N_2691,N_2737);
and U3594 (N_3594,N_2717,N_2224);
nand U3595 (N_3595,N_2442,N_2379);
or U3596 (N_3596,N_2263,N_2336);
and U3597 (N_3597,N_2899,N_2383);
nand U3598 (N_3598,N_2179,N_2723);
nand U3599 (N_3599,N_2475,N_2840);
and U3600 (N_3600,N_2633,N_2470);
nand U3601 (N_3601,N_2459,N_2396);
nand U3602 (N_3602,N_2575,N_2603);
nand U3603 (N_3603,N_2090,N_2184);
nor U3604 (N_3604,N_2707,N_2214);
nor U3605 (N_3605,N_2001,N_2913);
or U3606 (N_3606,N_2877,N_2979);
nor U3607 (N_3607,N_2531,N_2315);
nand U3608 (N_3608,N_2992,N_2751);
xor U3609 (N_3609,N_2124,N_2168);
nand U3610 (N_3610,N_2167,N_2781);
nand U3611 (N_3611,N_2346,N_2941);
or U3612 (N_3612,N_2017,N_2065);
nor U3613 (N_3613,N_2839,N_2668);
or U3614 (N_3614,N_2416,N_2167);
nand U3615 (N_3615,N_2097,N_2944);
nor U3616 (N_3616,N_2399,N_2395);
and U3617 (N_3617,N_2994,N_2503);
or U3618 (N_3618,N_2470,N_2189);
nor U3619 (N_3619,N_2654,N_2426);
and U3620 (N_3620,N_2339,N_2130);
nor U3621 (N_3621,N_2664,N_2137);
nor U3622 (N_3622,N_2697,N_2468);
nand U3623 (N_3623,N_2428,N_2442);
nand U3624 (N_3624,N_2151,N_2918);
and U3625 (N_3625,N_2360,N_2962);
nor U3626 (N_3626,N_2813,N_2568);
nor U3627 (N_3627,N_2954,N_2909);
and U3628 (N_3628,N_2732,N_2382);
nor U3629 (N_3629,N_2551,N_2163);
and U3630 (N_3630,N_2618,N_2643);
or U3631 (N_3631,N_2112,N_2044);
nor U3632 (N_3632,N_2621,N_2225);
or U3633 (N_3633,N_2196,N_2579);
xor U3634 (N_3634,N_2361,N_2881);
and U3635 (N_3635,N_2011,N_2198);
and U3636 (N_3636,N_2423,N_2135);
nand U3637 (N_3637,N_2611,N_2143);
or U3638 (N_3638,N_2257,N_2327);
or U3639 (N_3639,N_2435,N_2076);
nor U3640 (N_3640,N_2969,N_2207);
nand U3641 (N_3641,N_2522,N_2755);
and U3642 (N_3642,N_2589,N_2604);
or U3643 (N_3643,N_2220,N_2443);
and U3644 (N_3644,N_2611,N_2056);
nand U3645 (N_3645,N_2562,N_2637);
or U3646 (N_3646,N_2289,N_2429);
or U3647 (N_3647,N_2246,N_2894);
nand U3648 (N_3648,N_2814,N_2830);
nor U3649 (N_3649,N_2002,N_2736);
nor U3650 (N_3650,N_2425,N_2438);
and U3651 (N_3651,N_2799,N_2372);
nor U3652 (N_3652,N_2279,N_2147);
nand U3653 (N_3653,N_2532,N_2469);
nand U3654 (N_3654,N_2166,N_2342);
or U3655 (N_3655,N_2637,N_2874);
nor U3656 (N_3656,N_2138,N_2802);
nand U3657 (N_3657,N_2208,N_2552);
nor U3658 (N_3658,N_2139,N_2410);
nand U3659 (N_3659,N_2826,N_2190);
or U3660 (N_3660,N_2352,N_2595);
or U3661 (N_3661,N_2798,N_2582);
or U3662 (N_3662,N_2517,N_2795);
or U3663 (N_3663,N_2603,N_2068);
and U3664 (N_3664,N_2872,N_2760);
nand U3665 (N_3665,N_2115,N_2828);
and U3666 (N_3666,N_2939,N_2164);
nor U3667 (N_3667,N_2879,N_2301);
or U3668 (N_3668,N_2722,N_2250);
nand U3669 (N_3669,N_2109,N_2689);
nor U3670 (N_3670,N_2927,N_2521);
or U3671 (N_3671,N_2704,N_2413);
nor U3672 (N_3672,N_2957,N_2022);
nor U3673 (N_3673,N_2285,N_2522);
and U3674 (N_3674,N_2094,N_2549);
and U3675 (N_3675,N_2374,N_2127);
and U3676 (N_3676,N_2393,N_2128);
xor U3677 (N_3677,N_2406,N_2097);
or U3678 (N_3678,N_2709,N_2402);
and U3679 (N_3679,N_2590,N_2472);
or U3680 (N_3680,N_2982,N_2826);
nor U3681 (N_3681,N_2534,N_2176);
nand U3682 (N_3682,N_2919,N_2361);
or U3683 (N_3683,N_2733,N_2039);
and U3684 (N_3684,N_2378,N_2660);
or U3685 (N_3685,N_2806,N_2929);
nand U3686 (N_3686,N_2528,N_2401);
or U3687 (N_3687,N_2936,N_2425);
nand U3688 (N_3688,N_2922,N_2440);
and U3689 (N_3689,N_2147,N_2284);
and U3690 (N_3690,N_2653,N_2174);
or U3691 (N_3691,N_2655,N_2748);
and U3692 (N_3692,N_2989,N_2943);
nor U3693 (N_3693,N_2400,N_2241);
or U3694 (N_3694,N_2516,N_2668);
or U3695 (N_3695,N_2600,N_2572);
or U3696 (N_3696,N_2954,N_2606);
and U3697 (N_3697,N_2564,N_2731);
nand U3698 (N_3698,N_2188,N_2087);
or U3699 (N_3699,N_2756,N_2409);
nor U3700 (N_3700,N_2503,N_2309);
nand U3701 (N_3701,N_2759,N_2928);
nand U3702 (N_3702,N_2106,N_2129);
and U3703 (N_3703,N_2753,N_2211);
nand U3704 (N_3704,N_2320,N_2155);
or U3705 (N_3705,N_2988,N_2819);
nor U3706 (N_3706,N_2967,N_2244);
or U3707 (N_3707,N_2198,N_2807);
nor U3708 (N_3708,N_2454,N_2197);
xnor U3709 (N_3709,N_2368,N_2538);
and U3710 (N_3710,N_2088,N_2070);
and U3711 (N_3711,N_2541,N_2523);
or U3712 (N_3712,N_2844,N_2096);
nand U3713 (N_3713,N_2468,N_2951);
and U3714 (N_3714,N_2176,N_2173);
nor U3715 (N_3715,N_2819,N_2594);
xor U3716 (N_3716,N_2937,N_2974);
or U3717 (N_3717,N_2433,N_2147);
xor U3718 (N_3718,N_2145,N_2081);
and U3719 (N_3719,N_2725,N_2322);
or U3720 (N_3720,N_2461,N_2720);
nand U3721 (N_3721,N_2568,N_2871);
nor U3722 (N_3722,N_2586,N_2801);
nor U3723 (N_3723,N_2939,N_2857);
and U3724 (N_3724,N_2495,N_2604);
or U3725 (N_3725,N_2374,N_2490);
and U3726 (N_3726,N_2050,N_2307);
nand U3727 (N_3727,N_2908,N_2377);
nor U3728 (N_3728,N_2401,N_2423);
nand U3729 (N_3729,N_2843,N_2481);
xor U3730 (N_3730,N_2263,N_2317);
and U3731 (N_3731,N_2624,N_2294);
nor U3732 (N_3732,N_2620,N_2355);
nand U3733 (N_3733,N_2614,N_2997);
nor U3734 (N_3734,N_2996,N_2819);
nand U3735 (N_3735,N_2003,N_2035);
nand U3736 (N_3736,N_2749,N_2629);
and U3737 (N_3737,N_2539,N_2039);
and U3738 (N_3738,N_2304,N_2511);
nor U3739 (N_3739,N_2897,N_2106);
or U3740 (N_3740,N_2859,N_2909);
or U3741 (N_3741,N_2238,N_2678);
nor U3742 (N_3742,N_2798,N_2987);
or U3743 (N_3743,N_2580,N_2905);
and U3744 (N_3744,N_2792,N_2002);
or U3745 (N_3745,N_2268,N_2445);
and U3746 (N_3746,N_2995,N_2301);
nand U3747 (N_3747,N_2189,N_2776);
and U3748 (N_3748,N_2095,N_2773);
nand U3749 (N_3749,N_2445,N_2329);
nand U3750 (N_3750,N_2574,N_2264);
and U3751 (N_3751,N_2384,N_2716);
nor U3752 (N_3752,N_2601,N_2897);
nor U3753 (N_3753,N_2784,N_2311);
nand U3754 (N_3754,N_2127,N_2971);
and U3755 (N_3755,N_2207,N_2323);
and U3756 (N_3756,N_2592,N_2287);
nor U3757 (N_3757,N_2722,N_2958);
nor U3758 (N_3758,N_2091,N_2941);
nand U3759 (N_3759,N_2227,N_2124);
and U3760 (N_3760,N_2798,N_2060);
nand U3761 (N_3761,N_2635,N_2412);
and U3762 (N_3762,N_2987,N_2455);
nand U3763 (N_3763,N_2980,N_2669);
and U3764 (N_3764,N_2280,N_2307);
or U3765 (N_3765,N_2854,N_2171);
and U3766 (N_3766,N_2475,N_2884);
nand U3767 (N_3767,N_2347,N_2074);
or U3768 (N_3768,N_2323,N_2799);
or U3769 (N_3769,N_2691,N_2575);
and U3770 (N_3770,N_2301,N_2482);
nand U3771 (N_3771,N_2585,N_2600);
or U3772 (N_3772,N_2599,N_2064);
nand U3773 (N_3773,N_2638,N_2194);
or U3774 (N_3774,N_2282,N_2561);
nor U3775 (N_3775,N_2338,N_2662);
or U3776 (N_3776,N_2172,N_2999);
or U3777 (N_3777,N_2124,N_2878);
and U3778 (N_3778,N_2382,N_2903);
or U3779 (N_3779,N_2246,N_2729);
nor U3780 (N_3780,N_2932,N_2339);
and U3781 (N_3781,N_2638,N_2402);
nor U3782 (N_3782,N_2763,N_2526);
or U3783 (N_3783,N_2530,N_2783);
and U3784 (N_3784,N_2516,N_2786);
nand U3785 (N_3785,N_2519,N_2884);
and U3786 (N_3786,N_2726,N_2111);
nor U3787 (N_3787,N_2374,N_2323);
nor U3788 (N_3788,N_2137,N_2931);
and U3789 (N_3789,N_2613,N_2143);
nor U3790 (N_3790,N_2843,N_2772);
or U3791 (N_3791,N_2226,N_2307);
and U3792 (N_3792,N_2741,N_2727);
xor U3793 (N_3793,N_2954,N_2495);
nand U3794 (N_3794,N_2011,N_2522);
nand U3795 (N_3795,N_2529,N_2254);
and U3796 (N_3796,N_2528,N_2129);
nand U3797 (N_3797,N_2075,N_2344);
nor U3798 (N_3798,N_2868,N_2077);
nor U3799 (N_3799,N_2809,N_2859);
or U3800 (N_3800,N_2775,N_2689);
or U3801 (N_3801,N_2022,N_2164);
or U3802 (N_3802,N_2535,N_2613);
and U3803 (N_3803,N_2527,N_2598);
or U3804 (N_3804,N_2017,N_2033);
and U3805 (N_3805,N_2964,N_2784);
nor U3806 (N_3806,N_2624,N_2121);
nand U3807 (N_3807,N_2837,N_2451);
nor U3808 (N_3808,N_2457,N_2186);
nand U3809 (N_3809,N_2766,N_2349);
nor U3810 (N_3810,N_2378,N_2976);
or U3811 (N_3811,N_2766,N_2083);
and U3812 (N_3812,N_2567,N_2537);
nand U3813 (N_3813,N_2248,N_2701);
nand U3814 (N_3814,N_2001,N_2170);
and U3815 (N_3815,N_2962,N_2543);
nand U3816 (N_3816,N_2738,N_2174);
nand U3817 (N_3817,N_2998,N_2528);
nand U3818 (N_3818,N_2820,N_2546);
nor U3819 (N_3819,N_2946,N_2708);
or U3820 (N_3820,N_2964,N_2521);
nor U3821 (N_3821,N_2620,N_2095);
and U3822 (N_3822,N_2236,N_2348);
or U3823 (N_3823,N_2445,N_2855);
or U3824 (N_3824,N_2949,N_2182);
nand U3825 (N_3825,N_2228,N_2550);
nand U3826 (N_3826,N_2438,N_2733);
or U3827 (N_3827,N_2522,N_2784);
or U3828 (N_3828,N_2974,N_2129);
and U3829 (N_3829,N_2912,N_2556);
or U3830 (N_3830,N_2093,N_2642);
and U3831 (N_3831,N_2328,N_2756);
nor U3832 (N_3832,N_2312,N_2226);
nand U3833 (N_3833,N_2293,N_2866);
or U3834 (N_3834,N_2762,N_2914);
or U3835 (N_3835,N_2658,N_2072);
or U3836 (N_3836,N_2150,N_2575);
nor U3837 (N_3837,N_2367,N_2557);
nand U3838 (N_3838,N_2615,N_2154);
or U3839 (N_3839,N_2910,N_2494);
nor U3840 (N_3840,N_2717,N_2786);
nor U3841 (N_3841,N_2429,N_2889);
nand U3842 (N_3842,N_2292,N_2981);
nand U3843 (N_3843,N_2160,N_2540);
or U3844 (N_3844,N_2058,N_2889);
nand U3845 (N_3845,N_2018,N_2589);
and U3846 (N_3846,N_2274,N_2433);
nor U3847 (N_3847,N_2711,N_2829);
nand U3848 (N_3848,N_2927,N_2146);
and U3849 (N_3849,N_2655,N_2706);
and U3850 (N_3850,N_2499,N_2988);
xnor U3851 (N_3851,N_2770,N_2087);
and U3852 (N_3852,N_2848,N_2236);
or U3853 (N_3853,N_2557,N_2902);
or U3854 (N_3854,N_2739,N_2939);
nand U3855 (N_3855,N_2504,N_2611);
or U3856 (N_3856,N_2806,N_2812);
and U3857 (N_3857,N_2476,N_2678);
nand U3858 (N_3858,N_2572,N_2066);
nor U3859 (N_3859,N_2166,N_2082);
nand U3860 (N_3860,N_2635,N_2695);
or U3861 (N_3861,N_2213,N_2459);
nand U3862 (N_3862,N_2098,N_2404);
nor U3863 (N_3863,N_2789,N_2930);
or U3864 (N_3864,N_2030,N_2479);
nand U3865 (N_3865,N_2303,N_2819);
and U3866 (N_3866,N_2697,N_2759);
and U3867 (N_3867,N_2985,N_2187);
nand U3868 (N_3868,N_2676,N_2223);
nand U3869 (N_3869,N_2062,N_2322);
nand U3870 (N_3870,N_2203,N_2738);
and U3871 (N_3871,N_2481,N_2105);
nand U3872 (N_3872,N_2668,N_2400);
nand U3873 (N_3873,N_2282,N_2437);
and U3874 (N_3874,N_2395,N_2912);
and U3875 (N_3875,N_2078,N_2786);
and U3876 (N_3876,N_2332,N_2646);
nand U3877 (N_3877,N_2994,N_2271);
nor U3878 (N_3878,N_2507,N_2470);
or U3879 (N_3879,N_2549,N_2695);
nor U3880 (N_3880,N_2388,N_2878);
or U3881 (N_3881,N_2304,N_2748);
xor U3882 (N_3882,N_2645,N_2294);
nand U3883 (N_3883,N_2062,N_2780);
nand U3884 (N_3884,N_2412,N_2872);
nand U3885 (N_3885,N_2504,N_2661);
nand U3886 (N_3886,N_2392,N_2839);
nor U3887 (N_3887,N_2649,N_2964);
nor U3888 (N_3888,N_2413,N_2114);
and U3889 (N_3889,N_2188,N_2971);
nand U3890 (N_3890,N_2878,N_2039);
and U3891 (N_3891,N_2439,N_2607);
and U3892 (N_3892,N_2439,N_2393);
or U3893 (N_3893,N_2145,N_2545);
nor U3894 (N_3894,N_2971,N_2148);
nor U3895 (N_3895,N_2614,N_2216);
or U3896 (N_3896,N_2847,N_2017);
and U3897 (N_3897,N_2424,N_2783);
or U3898 (N_3898,N_2584,N_2015);
and U3899 (N_3899,N_2062,N_2028);
and U3900 (N_3900,N_2826,N_2297);
nand U3901 (N_3901,N_2384,N_2650);
xnor U3902 (N_3902,N_2334,N_2506);
and U3903 (N_3903,N_2738,N_2895);
nor U3904 (N_3904,N_2585,N_2399);
or U3905 (N_3905,N_2619,N_2667);
or U3906 (N_3906,N_2723,N_2993);
nor U3907 (N_3907,N_2878,N_2019);
nor U3908 (N_3908,N_2738,N_2138);
nand U3909 (N_3909,N_2172,N_2289);
nand U3910 (N_3910,N_2101,N_2611);
nor U3911 (N_3911,N_2888,N_2434);
nor U3912 (N_3912,N_2517,N_2974);
nand U3913 (N_3913,N_2034,N_2485);
nand U3914 (N_3914,N_2070,N_2317);
or U3915 (N_3915,N_2017,N_2053);
nor U3916 (N_3916,N_2372,N_2407);
or U3917 (N_3917,N_2663,N_2183);
and U3918 (N_3918,N_2668,N_2330);
nor U3919 (N_3919,N_2671,N_2457);
and U3920 (N_3920,N_2301,N_2559);
or U3921 (N_3921,N_2867,N_2982);
or U3922 (N_3922,N_2385,N_2233);
and U3923 (N_3923,N_2607,N_2823);
nand U3924 (N_3924,N_2507,N_2558);
and U3925 (N_3925,N_2399,N_2516);
and U3926 (N_3926,N_2557,N_2559);
nor U3927 (N_3927,N_2829,N_2054);
nand U3928 (N_3928,N_2103,N_2434);
nor U3929 (N_3929,N_2202,N_2038);
nand U3930 (N_3930,N_2070,N_2328);
and U3931 (N_3931,N_2306,N_2386);
nand U3932 (N_3932,N_2745,N_2276);
nor U3933 (N_3933,N_2546,N_2369);
or U3934 (N_3934,N_2330,N_2069);
nand U3935 (N_3935,N_2852,N_2336);
or U3936 (N_3936,N_2686,N_2747);
nand U3937 (N_3937,N_2004,N_2117);
xnor U3938 (N_3938,N_2291,N_2867);
nand U3939 (N_3939,N_2226,N_2033);
nor U3940 (N_3940,N_2191,N_2491);
nand U3941 (N_3941,N_2842,N_2218);
and U3942 (N_3942,N_2384,N_2222);
nand U3943 (N_3943,N_2926,N_2272);
and U3944 (N_3944,N_2213,N_2203);
nor U3945 (N_3945,N_2546,N_2166);
and U3946 (N_3946,N_2626,N_2544);
or U3947 (N_3947,N_2261,N_2495);
or U3948 (N_3948,N_2140,N_2196);
nor U3949 (N_3949,N_2113,N_2583);
nor U3950 (N_3950,N_2893,N_2259);
nand U3951 (N_3951,N_2526,N_2825);
or U3952 (N_3952,N_2549,N_2657);
nor U3953 (N_3953,N_2847,N_2559);
nor U3954 (N_3954,N_2163,N_2634);
and U3955 (N_3955,N_2715,N_2728);
nand U3956 (N_3956,N_2906,N_2917);
nand U3957 (N_3957,N_2062,N_2288);
or U3958 (N_3958,N_2324,N_2699);
or U3959 (N_3959,N_2087,N_2311);
or U3960 (N_3960,N_2563,N_2706);
or U3961 (N_3961,N_2323,N_2614);
nand U3962 (N_3962,N_2415,N_2516);
xor U3963 (N_3963,N_2394,N_2237);
or U3964 (N_3964,N_2636,N_2393);
nand U3965 (N_3965,N_2021,N_2944);
nand U3966 (N_3966,N_2519,N_2653);
and U3967 (N_3967,N_2168,N_2774);
nor U3968 (N_3968,N_2813,N_2097);
xor U3969 (N_3969,N_2732,N_2390);
and U3970 (N_3970,N_2772,N_2436);
and U3971 (N_3971,N_2153,N_2516);
or U3972 (N_3972,N_2028,N_2868);
or U3973 (N_3973,N_2867,N_2242);
nand U3974 (N_3974,N_2090,N_2012);
nand U3975 (N_3975,N_2957,N_2975);
nor U3976 (N_3976,N_2938,N_2667);
nand U3977 (N_3977,N_2879,N_2967);
and U3978 (N_3978,N_2199,N_2491);
or U3979 (N_3979,N_2094,N_2700);
nand U3980 (N_3980,N_2659,N_2304);
nor U3981 (N_3981,N_2629,N_2665);
or U3982 (N_3982,N_2234,N_2585);
nand U3983 (N_3983,N_2530,N_2504);
or U3984 (N_3984,N_2554,N_2803);
nand U3985 (N_3985,N_2056,N_2732);
xnor U3986 (N_3986,N_2676,N_2120);
or U3987 (N_3987,N_2652,N_2559);
or U3988 (N_3988,N_2370,N_2884);
nand U3989 (N_3989,N_2041,N_2063);
and U3990 (N_3990,N_2500,N_2703);
nor U3991 (N_3991,N_2792,N_2185);
nand U3992 (N_3992,N_2887,N_2616);
and U3993 (N_3993,N_2783,N_2228);
nor U3994 (N_3994,N_2975,N_2131);
nand U3995 (N_3995,N_2245,N_2209);
xor U3996 (N_3996,N_2370,N_2447);
or U3997 (N_3997,N_2280,N_2286);
nand U3998 (N_3998,N_2972,N_2132);
nand U3999 (N_3999,N_2015,N_2437);
nand U4000 (N_4000,N_3302,N_3116);
or U4001 (N_4001,N_3327,N_3576);
nand U4002 (N_4002,N_3352,N_3557);
nor U4003 (N_4003,N_3092,N_3425);
and U4004 (N_4004,N_3065,N_3593);
nand U4005 (N_4005,N_3978,N_3053);
or U4006 (N_4006,N_3742,N_3209);
and U4007 (N_4007,N_3395,N_3825);
or U4008 (N_4008,N_3719,N_3625);
nand U4009 (N_4009,N_3136,N_3312);
and U4010 (N_4010,N_3357,N_3084);
nand U4011 (N_4011,N_3752,N_3566);
or U4012 (N_4012,N_3580,N_3850);
nor U4013 (N_4013,N_3885,N_3358);
nand U4014 (N_4014,N_3161,N_3841);
or U4015 (N_4015,N_3316,N_3474);
and U4016 (N_4016,N_3134,N_3964);
or U4017 (N_4017,N_3293,N_3820);
or U4018 (N_4018,N_3674,N_3149);
or U4019 (N_4019,N_3592,N_3399);
and U4020 (N_4020,N_3659,N_3415);
and U4021 (N_4021,N_3722,N_3520);
nand U4022 (N_4022,N_3485,N_3274);
nor U4023 (N_4023,N_3433,N_3194);
nor U4024 (N_4024,N_3559,N_3087);
nand U4025 (N_4025,N_3698,N_3423);
nand U4026 (N_4026,N_3782,N_3950);
and U4027 (N_4027,N_3914,N_3379);
nor U4028 (N_4028,N_3107,N_3465);
and U4029 (N_4029,N_3029,N_3365);
and U4030 (N_4030,N_3754,N_3522);
and U4031 (N_4031,N_3220,N_3565);
nand U4032 (N_4032,N_3244,N_3085);
nand U4033 (N_4033,N_3102,N_3989);
nand U4034 (N_4034,N_3930,N_3034);
or U4035 (N_4035,N_3180,N_3815);
and U4036 (N_4036,N_3762,N_3119);
and U4037 (N_4037,N_3677,N_3708);
nand U4038 (N_4038,N_3787,N_3957);
or U4039 (N_4039,N_3620,N_3952);
and U4040 (N_4040,N_3819,N_3925);
nor U4041 (N_4041,N_3088,N_3689);
nor U4042 (N_4042,N_3036,N_3456);
xor U4043 (N_4043,N_3880,N_3490);
nand U4044 (N_4044,N_3804,N_3699);
nand U4045 (N_4045,N_3313,N_3486);
and U4046 (N_4046,N_3811,N_3893);
xor U4047 (N_4047,N_3051,N_3290);
nor U4048 (N_4048,N_3303,N_3702);
or U4049 (N_4049,N_3622,N_3460);
or U4050 (N_4050,N_3900,N_3604);
xnor U4051 (N_4051,N_3556,N_3636);
nor U4052 (N_4052,N_3377,N_3340);
nand U4053 (N_4053,N_3586,N_3650);
nand U4054 (N_4054,N_3905,N_3398);
nor U4055 (N_4055,N_3151,N_3493);
or U4056 (N_4056,N_3693,N_3019);
or U4057 (N_4057,N_3382,N_3956);
and U4058 (N_4058,N_3219,N_3928);
and U4059 (N_4059,N_3922,N_3959);
and U4060 (N_4060,N_3389,N_3942);
or U4061 (N_4061,N_3458,N_3550);
nand U4062 (N_4062,N_3401,N_3467);
nand U4063 (N_4063,N_3005,N_3445);
or U4064 (N_4064,N_3546,N_3129);
and U4065 (N_4065,N_3827,N_3201);
nand U4066 (N_4066,N_3795,N_3642);
nand U4067 (N_4067,N_3569,N_3283);
or U4068 (N_4068,N_3561,N_3749);
or U4069 (N_4069,N_3725,N_3282);
or U4070 (N_4070,N_3619,N_3778);
and U4071 (N_4071,N_3391,N_3598);
nand U4072 (N_4072,N_3332,N_3449);
or U4073 (N_4073,N_3344,N_3128);
nor U4074 (N_4074,N_3466,N_3295);
nand U4075 (N_4075,N_3488,N_3632);
nor U4076 (N_4076,N_3881,N_3847);
nand U4077 (N_4077,N_3008,N_3431);
or U4078 (N_4078,N_3127,N_3629);
and U4079 (N_4079,N_3383,N_3206);
or U4080 (N_4080,N_3003,N_3926);
nor U4081 (N_4081,N_3104,N_3857);
or U4082 (N_4082,N_3118,N_3866);
nand U4083 (N_4083,N_3413,N_3765);
and U4084 (N_4084,N_3786,N_3949);
or U4085 (N_4085,N_3788,N_3526);
nand U4086 (N_4086,N_3156,N_3169);
nor U4087 (N_4087,N_3342,N_3328);
or U4088 (N_4088,N_3388,N_3323);
nor U4089 (N_4089,N_3492,N_3061);
and U4090 (N_4090,N_3030,N_3172);
or U4091 (N_4091,N_3571,N_3213);
or U4092 (N_4092,N_3440,N_3020);
nand U4093 (N_4093,N_3977,N_3418);
and U4094 (N_4094,N_3807,N_3444);
or U4095 (N_4095,N_3744,N_3140);
nand U4096 (N_4096,N_3426,N_3867);
or U4097 (N_4097,N_3056,N_3938);
and U4098 (N_4098,N_3767,N_3532);
or U4099 (N_4099,N_3363,N_3774);
nor U4100 (N_4100,N_3835,N_3921);
nand U4101 (N_4101,N_3178,N_3609);
and U4102 (N_4102,N_3370,N_3376);
nand U4103 (N_4103,N_3972,N_3718);
nand U4104 (N_4104,N_3696,N_3549);
nand U4105 (N_4105,N_3270,N_3200);
and U4106 (N_4106,N_3063,N_3606);
nand U4107 (N_4107,N_3904,N_3548);
and U4108 (N_4108,N_3840,N_3975);
and U4109 (N_4109,N_3230,N_3325);
nand U4110 (N_4110,N_3182,N_3760);
nor U4111 (N_4111,N_3464,N_3494);
or U4112 (N_4112,N_3150,N_3160);
or U4113 (N_4113,N_3918,N_3692);
or U4114 (N_4114,N_3732,N_3417);
xor U4115 (N_4115,N_3663,N_3641);
nand U4116 (N_4116,N_3155,N_3145);
and U4117 (N_4117,N_3208,N_3748);
nor U4118 (N_4118,N_3254,N_3015);
or U4119 (N_4119,N_3585,N_3761);
nor U4120 (N_4120,N_3233,N_3753);
or U4121 (N_4121,N_3683,N_3372);
nand U4122 (N_4122,N_3511,N_3540);
and U4123 (N_4123,N_3607,N_3966);
nand U4124 (N_4124,N_3052,N_3876);
nand U4125 (N_4125,N_3125,N_3126);
nor U4126 (N_4126,N_3988,N_3789);
or U4127 (N_4127,N_3644,N_3745);
and U4128 (N_4128,N_3205,N_3064);
or U4129 (N_4129,N_3552,N_3285);
or U4130 (N_4130,N_3231,N_3082);
and U4131 (N_4131,N_3995,N_3454);
nand U4132 (N_4132,N_3680,N_3050);
nor U4133 (N_4133,N_3948,N_3793);
nand U4134 (N_4134,N_3730,N_3943);
nor U4135 (N_4135,N_3798,N_3993);
nand U4136 (N_4136,N_3672,N_3994);
nor U4137 (N_4137,N_3353,N_3971);
nor U4138 (N_4138,N_3953,N_3305);
xnor U4139 (N_4139,N_3378,N_3535);
or U4140 (N_4140,N_3470,N_3734);
nor U4141 (N_4141,N_3865,N_3682);
nand U4142 (N_4142,N_3249,N_3300);
or U4143 (N_4143,N_3211,N_3123);
nand U4144 (N_4144,N_3089,N_3545);
or U4145 (N_4145,N_3530,N_3027);
nor U4146 (N_4146,N_3755,N_3860);
xnor U4147 (N_4147,N_3714,N_3021);
and U4148 (N_4148,N_3864,N_3616);
and U4149 (N_4149,N_3687,N_3210);
xnor U4150 (N_4150,N_3845,N_3738);
nand U4151 (N_4151,N_3472,N_3475);
nor U4152 (N_4152,N_3094,N_3588);
xnor U4153 (N_4153,N_3503,N_3838);
nor U4154 (N_4154,N_3527,N_3414);
nor U4155 (N_4155,N_3255,N_3326);
nor U4156 (N_4156,N_3605,N_3217);
nor U4157 (N_4157,N_3481,N_3601);
and U4158 (N_4158,N_3846,N_3664);
nor U4159 (N_4159,N_3355,N_3531);
nand U4160 (N_4160,N_3074,N_3099);
nor U4161 (N_4161,N_3902,N_3832);
or U4162 (N_4162,N_3276,N_3412);
or U4163 (N_4163,N_3038,N_3842);
nor U4164 (N_4164,N_3035,N_3911);
or U4165 (N_4165,N_3013,N_3041);
nor U4166 (N_4166,N_3941,N_3004);
nor U4167 (N_4167,N_3910,N_3886);
or U4168 (N_4168,N_3157,N_3341);
and U4169 (N_4169,N_3783,N_3132);
nand U4170 (N_4170,N_3856,N_3248);
or U4171 (N_4171,N_3599,N_3017);
or U4172 (N_4172,N_3103,N_3181);
or U4173 (N_4173,N_3110,N_3101);
or U4174 (N_4174,N_3228,N_3534);
or U4175 (N_4175,N_3967,N_3784);
or U4176 (N_4176,N_3875,N_3600);
nor U4177 (N_4177,N_3919,N_3638);
and U4178 (N_4178,N_3721,N_3195);
or U4179 (N_4179,N_3288,N_3188);
nand U4180 (N_4180,N_3296,N_3808);
xnor U4181 (N_4181,N_3899,N_3174);
or U4182 (N_4182,N_3079,N_3309);
and U4183 (N_4183,N_3484,N_3190);
nor U4184 (N_4184,N_3595,N_3555);
and U4185 (N_4185,N_3512,N_3796);
nand U4186 (N_4186,N_3596,N_3521);
nor U4187 (N_4187,N_3429,N_3269);
nand U4188 (N_4188,N_3350,N_3739);
nor U4189 (N_4189,N_3777,N_3317);
and U4190 (N_4190,N_3076,N_3434);
nor U4191 (N_4191,N_3828,N_3311);
and U4192 (N_4192,N_3983,N_3649);
and U4193 (N_4193,N_3614,N_3694);
or U4194 (N_4194,N_3543,N_3558);
xor U4195 (N_4195,N_3315,N_3381);
and U4196 (N_4196,N_3916,N_3046);
and U4197 (N_4197,N_3697,N_3635);
nor U4198 (N_4198,N_3068,N_3772);
nor U4199 (N_4199,N_3896,N_3380);
nand U4200 (N_4200,N_3397,N_3816);
or U4201 (N_4201,N_3356,N_3982);
nor U4202 (N_4202,N_3320,N_3242);
nor U4203 (N_4203,N_3675,N_3997);
or U4204 (N_4204,N_3830,N_3277);
or U4205 (N_4205,N_3322,N_3590);
xor U4206 (N_4206,N_3478,N_3523);
or U4207 (N_4207,N_3022,N_3582);
nand U4208 (N_4208,N_3139,N_3243);
nand U4209 (N_4209,N_3985,N_3669);
nand U4210 (N_4210,N_3333,N_3093);
nand U4211 (N_4211,N_3477,N_3851);
xnor U4212 (N_4212,N_3098,N_3979);
and U4213 (N_4213,N_3268,N_3678);
nor U4214 (N_4214,N_3304,N_3564);
and U4215 (N_4215,N_3045,N_3758);
nor U4216 (N_4216,N_3096,N_3081);
nand U4217 (N_4217,N_3075,N_3498);
or U4218 (N_4218,N_3554,N_3179);
nand U4219 (N_4219,N_3387,N_3280);
or U4220 (N_4220,N_3791,N_3077);
nor U4221 (N_4221,N_3097,N_3373);
and U4222 (N_4222,N_3222,N_3040);
and U4223 (N_4223,N_3792,N_3108);
nor U4224 (N_4224,N_3062,N_3324);
nor U4225 (N_4225,N_3167,N_3023);
nor U4226 (N_4226,N_3501,N_3319);
nor U4227 (N_4227,N_3048,N_3671);
nor U4228 (N_4228,N_3289,N_3236);
xnor U4229 (N_4229,N_3199,N_3007);
nor U4230 (N_4230,N_3025,N_3653);
nand U4231 (N_4231,N_3164,N_3482);
or U4232 (N_4232,N_3516,N_3407);
nand U4233 (N_4233,N_3452,N_3539);
nor U4234 (N_4234,N_3894,N_3766);
and U4235 (N_4235,N_3717,N_3196);
nand U4236 (N_4236,N_3113,N_3281);
nor U4237 (N_4237,N_3651,N_3121);
and U4238 (N_4238,N_3197,N_3861);
and U4239 (N_4239,N_3897,N_3756);
or U4240 (N_4240,N_3901,N_3275);
nand U4241 (N_4241,N_3903,N_3855);
and U4242 (N_4242,N_3733,N_3505);
and U4243 (N_4243,N_3240,N_3623);
nor U4244 (N_4244,N_3541,N_3510);
or U4245 (N_4245,N_3091,N_3594);
or U4246 (N_4246,N_3504,N_3529);
nand U4247 (N_4247,N_3831,N_3170);
nor U4248 (N_4248,N_3043,N_3962);
or U4249 (N_4249,N_3273,N_3042);
nor U4250 (N_4250,N_3335,N_3416);
nor U4251 (N_4251,N_3879,N_3681);
and U4252 (N_4252,N_3495,N_3451);
nand U4253 (N_4253,N_3848,N_3781);
nand U4254 (N_4254,N_3078,N_3430);
nand U4255 (N_4255,N_3610,N_3297);
nor U4256 (N_4256,N_3310,N_3345);
nor U4257 (N_4257,N_3337,N_3567);
nand U4258 (N_4258,N_3822,N_3973);
and U4259 (N_4259,N_3839,N_3990);
nand U4260 (N_4260,N_3266,N_3869);
nand U4261 (N_4261,N_3525,N_3656);
nor U4262 (N_4262,N_3727,N_3386);
nor U4263 (N_4263,N_3006,N_3974);
and U4264 (N_4264,N_3823,N_3611);
or U4265 (N_4265,N_3083,N_3951);
nor U4266 (N_4266,N_3508,N_3216);
nand U4267 (N_4267,N_3260,N_3496);
nor U4268 (N_4268,N_3602,N_3970);
and U4269 (N_4269,N_3801,N_3346);
or U4270 (N_4270,N_3441,N_3028);
nand U4271 (N_4271,N_3471,N_3165);
or U4272 (N_4272,N_3166,N_3716);
nand U4273 (N_4273,N_3907,N_3001);
nand U4274 (N_4274,N_3768,N_3307);
and U4275 (N_4275,N_3238,N_3502);
or U4276 (N_4276,N_3012,N_3575);
and U4277 (N_4277,N_3963,N_3497);
nand U4278 (N_4278,N_3895,N_3059);
nand U4279 (N_4279,N_3929,N_3690);
nand U4280 (N_4280,N_3321,N_3618);
nor U4281 (N_4281,N_3553,N_3259);
nand U4282 (N_4282,N_3154,N_3818);
nand U4283 (N_4283,N_3223,N_3453);
or U4284 (N_4284,N_3873,N_3987);
nand U4285 (N_4285,N_3203,N_3785);
nor U4286 (N_4286,N_3507,N_3400);
nor U4287 (N_4287,N_3250,N_3264);
nand U4288 (N_4288,N_3836,N_3646);
or U4289 (N_4289,N_3267,N_3655);
nand U4290 (N_4290,N_3491,N_3735);
xor U4291 (N_4291,N_3647,N_3991);
nand U4292 (N_4292,N_3999,N_3634);
or U4293 (N_4293,N_3780,N_3359);
nand U4294 (N_4294,N_3701,N_3146);
nand U4295 (N_4295,N_3448,N_3750);
and U4296 (N_4296,N_3331,N_3299);
nand U4297 (N_4297,N_3737,N_3329);
or U4298 (N_4298,N_3863,N_3954);
or U4299 (N_4299,N_3461,N_3192);
nor U4300 (N_4300,N_3877,N_3579);
and U4301 (N_4301,N_3884,N_3821);
and U4302 (N_4302,N_3229,N_3080);
and U4303 (N_4303,N_3292,N_3878);
nor U4304 (N_4304,N_3060,N_3958);
or U4305 (N_4305,N_3723,N_3854);
nor U4306 (N_4306,N_3584,N_3130);
and U4307 (N_4307,N_3731,N_3396);
and U4308 (N_4308,N_3743,N_3067);
nor U4309 (N_4309,N_3660,N_3621);
and U4310 (N_4310,N_3252,N_3524);
or U4311 (N_4311,N_3763,N_3162);
and U4312 (N_4312,N_3237,N_3829);
or U4313 (N_4313,N_3314,N_3256);
or U4314 (N_4314,N_3131,N_3769);
or U4315 (N_4315,N_3891,N_3287);
or U4316 (N_4316,N_3890,N_3436);
nand U4317 (N_4317,N_3446,N_3872);
nand U4318 (N_4318,N_3538,N_3679);
and U4319 (N_4319,N_3898,N_3120);
nand U4320 (N_4320,N_3262,N_3805);
nor U4321 (N_4321,N_3726,N_3403);
and U4322 (N_4322,N_3142,N_3137);
and U4323 (N_4323,N_3667,N_3405);
or U4324 (N_4324,N_3703,N_3562);
or U4325 (N_4325,N_3544,N_3214);
and U4326 (N_4326,N_3057,N_3528);
and U4327 (N_4327,N_3519,N_3318);
nand U4328 (N_4328,N_3463,N_3648);
nor U4329 (N_4329,N_3676,N_3657);
and U4330 (N_4330,N_3643,N_3759);
and U4331 (N_4331,N_3124,N_3133);
nor U4332 (N_4332,N_3257,N_3578);
or U4333 (N_4333,N_3946,N_3058);
or U4334 (N_4334,N_3100,N_3980);
nor U4335 (N_4335,N_3563,N_3171);
nand U4336 (N_4336,N_3360,N_3284);
xor U4337 (N_4337,N_3258,N_3779);
and U4338 (N_4338,N_3207,N_3152);
or U4339 (N_4339,N_3141,N_3961);
and U4340 (N_4340,N_3095,N_3221);
nor U4341 (N_4341,N_3912,N_3707);
nand U4342 (N_4342,N_3039,N_3122);
nand U4343 (N_4343,N_3944,N_3457);
nor U4344 (N_4344,N_3969,N_3711);
and U4345 (N_4345,N_3709,N_3715);
and U4346 (N_4346,N_3603,N_3515);
or U4347 (N_4347,N_3976,N_3551);
nor U4348 (N_4348,N_3392,N_3934);
or U4349 (N_4349,N_3047,N_3802);
nor U4350 (N_4350,N_3408,N_3764);
and U4351 (N_4351,N_3633,N_3371);
nor U4352 (N_4352,N_3591,N_3069);
and U4353 (N_4353,N_3892,N_3746);
nor U4354 (N_4354,N_3343,N_3480);
nor U4355 (N_4355,N_3009,N_3932);
or U4356 (N_4356,N_3741,N_3560);
or U4357 (N_4357,N_3246,N_3695);
nand U4358 (N_4358,N_3513,N_3455);
nand U4359 (N_4359,N_3010,N_3874);
nand U4360 (N_4360,N_3945,N_3018);
nand U4361 (N_4361,N_3394,N_3443);
or U4362 (N_4362,N_3364,N_3105);
nor U4363 (N_4363,N_3837,N_3410);
nand U4364 (N_4364,N_3235,N_3888);
and U4365 (N_4365,N_3913,N_3992);
or U4366 (N_4366,N_3011,N_3700);
nand U4367 (N_4367,N_3826,N_3361);
or U4368 (N_4368,N_3965,N_3114);
nand U4369 (N_4369,N_3462,N_3354);
nor U4370 (N_4370,N_3232,N_3138);
nor U4371 (N_4371,N_3245,N_3797);
or U4372 (N_4372,N_3583,N_3349);
or U4373 (N_4373,N_3112,N_3773);
nand U4374 (N_4374,N_3514,N_3447);
xor U4375 (N_4375,N_3882,N_3577);
and U4376 (N_4376,N_3814,N_3186);
and U4377 (N_4377,N_3049,N_3234);
or U4378 (N_4378,N_3163,N_3198);
and U4379 (N_4379,N_3868,N_3568);
nor U4380 (N_4380,N_3817,N_3608);
and U4381 (N_4381,N_3177,N_3435);
nand U4382 (N_4382,N_3306,N_3574);
nor U4383 (N_4383,N_3986,N_3483);
nand U4384 (N_4384,N_3909,N_3185);
or U4385 (N_4385,N_3573,N_3843);
or U4386 (N_4386,N_3937,N_3627);
nand U4387 (N_4387,N_3261,N_3668);
or U4388 (N_4388,N_3427,N_3032);
or U4389 (N_4389,N_3639,N_3628);
and U4390 (N_4390,N_3686,N_3247);
nor U4391 (N_4391,N_3518,N_3024);
and U4392 (N_4392,N_3547,N_3661);
nor U4393 (N_4393,N_3109,N_3940);
or U4394 (N_4394,N_3000,N_3710);
or U4395 (N_4395,N_3153,N_3645);
nor U4396 (N_4396,N_3747,N_3115);
and U4397 (N_4397,N_3813,N_3450);
or U4398 (N_4398,N_3135,N_3637);
or U4399 (N_4399,N_3158,N_3640);
nor U4400 (N_4400,N_3375,N_3612);
nand U4401 (N_4401,N_3824,N_3241);
nand U4402 (N_4402,N_3889,N_3615);
nor U4403 (N_4403,N_3033,N_3409);
nand U4404 (N_4404,N_3173,N_3368);
xnor U4405 (N_4405,N_3202,N_3442);
or U4406 (N_4406,N_3736,N_3968);
nand U4407 (N_4407,N_3833,N_3626);
and U4408 (N_4408,N_3106,N_3168);
nand U4409 (N_4409,N_3487,N_3298);
and U4410 (N_4410,N_3271,N_3055);
and U4411 (N_4411,N_3887,N_3390);
nor U4412 (N_4412,N_3770,N_3432);
and U4413 (N_4413,N_3111,N_3996);
or U4414 (N_4414,N_3666,N_3479);
and U4415 (N_4415,N_3489,N_3336);
nand U4416 (N_4416,N_3542,N_3175);
nand U4417 (N_4417,N_3706,N_3803);
or U4418 (N_4418,N_3031,N_3421);
and U4419 (N_4419,N_3572,N_3226);
or U4420 (N_4420,N_3927,N_3631);
and U4421 (N_4421,N_3385,N_3920);
nor U4422 (N_4422,N_3799,N_3704);
and U4423 (N_4423,N_3347,N_3037);
and U4424 (N_4424,N_3339,N_3691);
nor U4425 (N_4425,N_3422,N_3844);
nand U4426 (N_4426,N_3251,N_3908);
nand U4427 (N_4427,N_3187,N_3499);
and U4428 (N_4428,N_3367,N_3740);
and U4429 (N_4429,N_3086,N_3054);
and U4430 (N_4430,N_3670,N_3148);
nand U4431 (N_4431,N_3705,N_3939);
nor U4432 (N_4432,N_3026,N_3189);
nand U4433 (N_4433,N_3771,N_3712);
xor U4434 (N_4434,N_3570,N_3215);
and U4435 (N_4435,N_3362,N_3351);
nand U4436 (N_4436,N_3533,N_3665);
nand U4437 (N_4437,N_3286,N_3070);
nand U4438 (N_4438,N_3159,N_3852);
nor U4439 (N_4439,N_3955,N_3853);
nor U4440 (N_4440,N_3419,N_3117);
nor U4441 (N_4441,N_3144,N_3193);
nand U4442 (N_4442,N_3301,N_3366);
nor U4443 (N_4443,N_3473,N_3617);
or U4444 (N_4444,N_3924,N_3834);
and U4445 (N_4445,N_3016,N_3673);
nor U4446 (N_4446,N_3263,N_3800);
nand U4447 (N_4447,N_3775,N_3509);
xnor U4448 (N_4448,N_3662,N_3374);
or U4449 (N_4449,N_3517,N_3859);
or U4450 (N_4450,N_3809,N_3871);
or U4451 (N_4451,N_3581,N_3685);
or U4452 (N_4452,N_3308,N_3072);
and U4453 (N_4453,N_3688,N_3224);
nand U4454 (N_4454,N_3684,N_3729);
or U4455 (N_4455,N_3384,N_3073);
nor U4456 (N_4456,N_3506,N_3143);
and U4457 (N_4457,N_3212,N_3402);
and U4458 (N_4458,N_3652,N_3147);
and U4459 (N_4459,N_3728,N_3984);
nor U4460 (N_4460,N_3066,N_3906);
nand U4461 (N_4461,N_3239,N_3338);
nand U4462 (N_4462,N_3624,N_3776);
and U4463 (N_4463,N_3812,N_3947);
and U4464 (N_4464,N_3044,N_3630);
nand U4465 (N_4465,N_3468,N_3393);
or U4466 (N_4466,N_3183,N_3790);
or U4467 (N_4467,N_3915,N_3176);
nand U4468 (N_4468,N_3935,N_3870);
and U4469 (N_4469,N_3981,N_3654);
nor U4470 (N_4470,N_3428,N_3279);
nor U4471 (N_4471,N_3227,N_3537);
nor U4472 (N_4472,N_3438,N_3757);
or U4473 (N_4473,N_3369,N_3713);
nand U4474 (N_4474,N_3272,N_3294);
nor U4475 (N_4475,N_3420,N_3424);
and U4476 (N_4476,N_3002,N_3348);
or U4477 (N_4477,N_3404,N_3724);
nand U4478 (N_4478,N_3225,N_3794);
nand U4479 (N_4479,N_3658,N_3883);
or U4480 (N_4480,N_3810,N_3936);
and U4481 (N_4481,N_3476,N_3931);
nor U4482 (N_4482,N_3334,N_3253);
nor U4483 (N_4483,N_3960,N_3330);
or U4484 (N_4484,N_3459,N_3437);
nor U4485 (N_4485,N_3014,N_3998);
or U4486 (N_4486,N_3933,N_3406);
or U4487 (N_4487,N_3589,N_3500);
nand U4488 (N_4488,N_3411,N_3858);
nor U4489 (N_4489,N_3917,N_3090);
nand U4490 (N_4490,N_3291,N_3923);
nor U4491 (N_4491,N_3278,N_3849);
nand U4492 (N_4492,N_3469,N_3806);
nand U4493 (N_4493,N_3536,N_3265);
nand U4494 (N_4494,N_3439,N_3204);
nor U4495 (N_4495,N_3862,N_3613);
nand U4496 (N_4496,N_3184,N_3191);
nand U4497 (N_4497,N_3720,N_3587);
nand U4498 (N_4498,N_3597,N_3071);
or U4499 (N_4499,N_3218,N_3751);
or U4500 (N_4500,N_3642,N_3402);
nor U4501 (N_4501,N_3160,N_3229);
nor U4502 (N_4502,N_3832,N_3536);
nand U4503 (N_4503,N_3931,N_3409);
or U4504 (N_4504,N_3092,N_3130);
nand U4505 (N_4505,N_3810,N_3674);
nand U4506 (N_4506,N_3234,N_3137);
xnor U4507 (N_4507,N_3450,N_3909);
nor U4508 (N_4508,N_3472,N_3662);
or U4509 (N_4509,N_3260,N_3070);
and U4510 (N_4510,N_3211,N_3067);
or U4511 (N_4511,N_3391,N_3734);
nand U4512 (N_4512,N_3445,N_3770);
nand U4513 (N_4513,N_3618,N_3311);
nor U4514 (N_4514,N_3050,N_3463);
or U4515 (N_4515,N_3110,N_3959);
nor U4516 (N_4516,N_3679,N_3135);
nor U4517 (N_4517,N_3800,N_3767);
nor U4518 (N_4518,N_3296,N_3955);
nand U4519 (N_4519,N_3969,N_3840);
nand U4520 (N_4520,N_3735,N_3133);
nor U4521 (N_4521,N_3804,N_3924);
nor U4522 (N_4522,N_3708,N_3426);
nand U4523 (N_4523,N_3099,N_3124);
or U4524 (N_4524,N_3225,N_3490);
and U4525 (N_4525,N_3840,N_3309);
or U4526 (N_4526,N_3405,N_3825);
or U4527 (N_4527,N_3340,N_3954);
and U4528 (N_4528,N_3251,N_3056);
or U4529 (N_4529,N_3598,N_3967);
or U4530 (N_4530,N_3180,N_3064);
and U4531 (N_4531,N_3766,N_3071);
or U4532 (N_4532,N_3498,N_3125);
and U4533 (N_4533,N_3067,N_3821);
or U4534 (N_4534,N_3406,N_3630);
and U4535 (N_4535,N_3264,N_3025);
or U4536 (N_4536,N_3314,N_3849);
and U4537 (N_4537,N_3866,N_3102);
nor U4538 (N_4538,N_3233,N_3465);
nor U4539 (N_4539,N_3027,N_3967);
and U4540 (N_4540,N_3393,N_3048);
nand U4541 (N_4541,N_3685,N_3273);
or U4542 (N_4542,N_3526,N_3959);
xnor U4543 (N_4543,N_3283,N_3937);
nor U4544 (N_4544,N_3434,N_3074);
or U4545 (N_4545,N_3041,N_3531);
nand U4546 (N_4546,N_3992,N_3027);
and U4547 (N_4547,N_3590,N_3175);
nor U4548 (N_4548,N_3658,N_3877);
and U4549 (N_4549,N_3646,N_3871);
and U4550 (N_4550,N_3539,N_3777);
nand U4551 (N_4551,N_3226,N_3512);
or U4552 (N_4552,N_3550,N_3936);
and U4553 (N_4553,N_3955,N_3829);
nand U4554 (N_4554,N_3968,N_3274);
nand U4555 (N_4555,N_3142,N_3373);
or U4556 (N_4556,N_3701,N_3655);
nand U4557 (N_4557,N_3976,N_3037);
xor U4558 (N_4558,N_3282,N_3863);
nand U4559 (N_4559,N_3426,N_3935);
or U4560 (N_4560,N_3309,N_3502);
nand U4561 (N_4561,N_3392,N_3243);
and U4562 (N_4562,N_3742,N_3517);
and U4563 (N_4563,N_3061,N_3069);
nor U4564 (N_4564,N_3857,N_3255);
nor U4565 (N_4565,N_3903,N_3128);
nand U4566 (N_4566,N_3244,N_3245);
or U4567 (N_4567,N_3824,N_3640);
and U4568 (N_4568,N_3012,N_3722);
or U4569 (N_4569,N_3903,N_3838);
or U4570 (N_4570,N_3842,N_3461);
nand U4571 (N_4571,N_3850,N_3835);
or U4572 (N_4572,N_3550,N_3885);
nor U4573 (N_4573,N_3193,N_3554);
nand U4574 (N_4574,N_3439,N_3011);
and U4575 (N_4575,N_3515,N_3258);
nand U4576 (N_4576,N_3979,N_3542);
nor U4577 (N_4577,N_3135,N_3393);
nand U4578 (N_4578,N_3406,N_3277);
and U4579 (N_4579,N_3806,N_3541);
and U4580 (N_4580,N_3690,N_3196);
nor U4581 (N_4581,N_3483,N_3634);
or U4582 (N_4582,N_3648,N_3563);
and U4583 (N_4583,N_3928,N_3068);
or U4584 (N_4584,N_3922,N_3650);
nor U4585 (N_4585,N_3389,N_3378);
and U4586 (N_4586,N_3552,N_3764);
nand U4587 (N_4587,N_3756,N_3121);
and U4588 (N_4588,N_3656,N_3515);
or U4589 (N_4589,N_3767,N_3229);
or U4590 (N_4590,N_3492,N_3639);
nor U4591 (N_4591,N_3222,N_3750);
or U4592 (N_4592,N_3423,N_3276);
nor U4593 (N_4593,N_3470,N_3909);
and U4594 (N_4594,N_3987,N_3389);
nor U4595 (N_4595,N_3462,N_3916);
and U4596 (N_4596,N_3867,N_3353);
nor U4597 (N_4597,N_3778,N_3642);
and U4598 (N_4598,N_3506,N_3551);
nand U4599 (N_4599,N_3493,N_3271);
and U4600 (N_4600,N_3427,N_3994);
and U4601 (N_4601,N_3260,N_3689);
xor U4602 (N_4602,N_3705,N_3789);
and U4603 (N_4603,N_3927,N_3247);
nand U4604 (N_4604,N_3386,N_3101);
and U4605 (N_4605,N_3552,N_3187);
nand U4606 (N_4606,N_3055,N_3036);
nand U4607 (N_4607,N_3553,N_3668);
nor U4608 (N_4608,N_3932,N_3854);
and U4609 (N_4609,N_3729,N_3339);
and U4610 (N_4610,N_3986,N_3255);
nor U4611 (N_4611,N_3441,N_3984);
and U4612 (N_4612,N_3048,N_3701);
nor U4613 (N_4613,N_3829,N_3395);
or U4614 (N_4614,N_3030,N_3941);
nand U4615 (N_4615,N_3946,N_3482);
nor U4616 (N_4616,N_3992,N_3970);
and U4617 (N_4617,N_3514,N_3978);
nand U4618 (N_4618,N_3328,N_3337);
and U4619 (N_4619,N_3988,N_3209);
or U4620 (N_4620,N_3730,N_3805);
or U4621 (N_4621,N_3019,N_3647);
nor U4622 (N_4622,N_3192,N_3197);
or U4623 (N_4623,N_3665,N_3418);
nand U4624 (N_4624,N_3276,N_3254);
and U4625 (N_4625,N_3419,N_3696);
and U4626 (N_4626,N_3009,N_3456);
or U4627 (N_4627,N_3769,N_3928);
or U4628 (N_4628,N_3319,N_3555);
xnor U4629 (N_4629,N_3701,N_3355);
and U4630 (N_4630,N_3661,N_3488);
nand U4631 (N_4631,N_3727,N_3779);
and U4632 (N_4632,N_3212,N_3925);
nand U4633 (N_4633,N_3635,N_3525);
and U4634 (N_4634,N_3977,N_3596);
nor U4635 (N_4635,N_3444,N_3590);
nand U4636 (N_4636,N_3293,N_3502);
and U4637 (N_4637,N_3884,N_3983);
or U4638 (N_4638,N_3203,N_3207);
nor U4639 (N_4639,N_3319,N_3945);
or U4640 (N_4640,N_3575,N_3465);
nor U4641 (N_4641,N_3748,N_3432);
nor U4642 (N_4642,N_3633,N_3994);
and U4643 (N_4643,N_3387,N_3351);
nand U4644 (N_4644,N_3880,N_3001);
nand U4645 (N_4645,N_3140,N_3116);
nand U4646 (N_4646,N_3734,N_3788);
or U4647 (N_4647,N_3531,N_3055);
and U4648 (N_4648,N_3894,N_3053);
and U4649 (N_4649,N_3564,N_3107);
or U4650 (N_4650,N_3317,N_3833);
and U4651 (N_4651,N_3244,N_3191);
nor U4652 (N_4652,N_3006,N_3297);
or U4653 (N_4653,N_3636,N_3340);
nor U4654 (N_4654,N_3122,N_3659);
or U4655 (N_4655,N_3013,N_3886);
nor U4656 (N_4656,N_3957,N_3706);
nor U4657 (N_4657,N_3814,N_3741);
or U4658 (N_4658,N_3470,N_3874);
nor U4659 (N_4659,N_3454,N_3125);
nor U4660 (N_4660,N_3336,N_3164);
nand U4661 (N_4661,N_3918,N_3602);
and U4662 (N_4662,N_3251,N_3566);
nor U4663 (N_4663,N_3063,N_3380);
or U4664 (N_4664,N_3477,N_3331);
nand U4665 (N_4665,N_3080,N_3280);
and U4666 (N_4666,N_3690,N_3020);
nor U4667 (N_4667,N_3427,N_3915);
or U4668 (N_4668,N_3474,N_3759);
nand U4669 (N_4669,N_3706,N_3454);
nor U4670 (N_4670,N_3576,N_3498);
nand U4671 (N_4671,N_3769,N_3664);
and U4672 (N_4672,N_3573,N_3756);
or U4673 (N_4673,N_3035,N_3364);
and U4674 (N_4674,N_3118,N_3354);
or U4675 (N_4675,N_3245,N_3863);
xnor U4676 (N_4676,N_3170,N_3077);
and U4677 (N_4677,N_3164,N_3568);
nand U4678 (N_4678,N_3720,N_3634);
xnor U4679 (N_4679,N_3412,N_3640);
nor U4680 (N_4680,N_3391,N_3819);
nor U4681 (N_4681,N_3330,N_3402);
nand U4682 (N_4682,N_3311,N_3288);
and U4683 (N_4683,N_3978,N_3952);
and U4684 (N_4684,N_3062,N_3111);
nor U4685 (N_4685,N_3991,N_3588);
xor U4686 (N_4686,N_3169,N_3736);
nand U4687 (N_4687,N_3047,N_3178);
and U4688 (N_4688,N_3760,N_3159);
nor U4689 (N_4689,N_3463,N_3584);
and U4690 (N_4690,N_3529,N_3846);
nor U4691 (N_4691,N_3119,N_3731);
nor U4692 (N_4692,N_3351,N_3774);
or U4693 (N_4693,N_3423,N_3034);
or U4694 (N_4694,N_3122,N_3521);
and U4695 (N_4695,N_3132,N_3989);
or U4696 (N_4696,N_3671,N_3983);
nand U4697 (N_4697,N_3365,N_3139);
or U4698 (N_4698,N_3473,N_3514);
and U4699 (N_4699,N_3703,N_3054);
and U4700 (N_4700,N_3516,N_3925);
nand U4701 (N_4701,N_3609,N_3598);
nor U4702 (N_4702,N_3864,N_3143);
and U4703 (N_4703,N_3233,N_3361);
nand U4704 (N_4704,N_3612,N_3175);
or U4705 (N_4705,N_3749,N_3083);
nand U4706 (N_4706,N_3977,N_3270);
or U4707 (N_4707,N_3039,N_3202);
xor U4708 (N_4708,N_3572,N_3338);
and U4709 (N_4709,N_3637,N_3581);
nand U4710 (N_4710,N_3519,N_3774);
or U4711 (N_4711,N_3666,N_3952);
and U4712 (N_4712,N_3287,N_3244);
and U4713 (N_4713,N_3601,N_3304);
nand U4714 (N_4714,N_3511,N_3627);
nor U4715 (N_4715,N_3870,N_3599);
or U4716 (N_4716,N_3469,N_3716);
and U4717 (N_4717,N_3837,N_3685);
nand U4718 (N_4718,N_3374,N_3000);
and U4719 (N_4719,N_3373,N_3356);
nor U4720 (N_4720,N_3884,N_3656);
or U4721 (N_4721,N_3428,N_3515);
and U4722 (N_4722,N_3649,N_3214);
and U4723 (N_4723,N_3442,N_3225);
nand U4724 (N_4724,N_3125,N_3250);
nor U4725 (N_4725,N_3166,N_3727);
nand U4726 (N_4726,N_3517,N_3019);
and U4727 (N_4727,N_3911,N_3761);
or U4728 (N_4728,N_3875,N_3102);
nor U4729 (N_4729,N_3947,N_3029);
nand U4730 (N_4730,N_3246,N_3766);
nand U4731 (N_4731,N_3002,N_3103);
nand U4732 (N_4732,N_3650,N_3909);
xnor U4733 (N_4733,N_3316,N_3649);
or U4734 (N_4734,N_3361,N_3609);
and U4735 (N_4735,N_3028,N_3086);
and U4736 (N_4736,N_3809,N_3559);
and U4737 (N_4737,N_3798,N_3931);
and U4738 (N_4738,N_3166,N_3939);
nor U4739 (N_4739,N_3847,N_3761);
nor U4740 (N_4740,N_3409,N_3510);
and U4741 (N_4741,N_3201,N_3984);
nand U4742 (N_4742,N_3709,N_3541);
or U4743 (N_4743,N_3842,N_3144);
nor U4744 (N_4744,N_3531,N_3913);
or U4745 (N_4745,N_3973,N_3611);
or U4746 (N_4746,N_3190,N_3899);
or U4747 (N_4747,N_3515,N_3994);
nor U4748 (N_4748,N_3569,N_3739);
nand U4749 (N_4749,N_3844,N_3228);
and U4750 (N_4750,N_3466,N_3211);
nor U4751 (N_4751,N_3030,N_3773);
and U4752 (N_4752,N_3624,N_3297);
or U4753 (N_4753,N_3062,N_3775);
nor U4754 (N_4754,N_3625,N_3005);
and U4755 (N_4755,N_3390,N_3347);
nand U4756 (N_4756,N_3375,N_3887);
nand U4757 (N_4757,N_3296,N_3494);
or U4758 (N_4758,N_3042,N_3341);
or U4759 (N_4759,N_3223,N_3459);
nand U4760 (N_4760,N_3168,N_3340);
nor U4761 (N_4761,N_3837,N_3306);
or U4762 (N_4762,N_3868,N_3990);
or U4763 (N_4763,N_3341,N_3754);
or U4764 (N_4764,N_3895,N_3681);
and U4765 (N_4765,N_3632,N_3744);
nand U4766 (N_4766,N_3850,N_3623);
or U4767 (N_4767,N_3667,N_3842);
nand U4768 (N_4768,N_3410,N_3392);
xor U4769 (N_4769,N_3966,N_3199);
nand U4770 (N_4770,N_3020,N_3427);
nand U4771 (N_4771,N_3434,N_3803);
nor U4772 (N_4772,N_3632,N_3358);
nor U4773 (N_4773,N_3177,N_3851);
and U4774 (N_4774,N_3174,N_3751);
or U4775 (N_4775,N_3917,N_3875);
nor U4776 (N_4776,N_3100,N_3928);
and U4777 (N_4777,N_3021,N_3371);
nand U4778 (N_4778,N_3486,N_3664);
nand U4779 (N_4779,N_3027,N_3151);
and U4780 (N_4780,N_3177,N_3717);
nand U4781 (N_4781,N_3044,N_3312);
or U4782 (N_4782,N_3475,N_3484);
or U4783 (N_4783,N_3114,N_3314);
or U4784 (N_4784,N_3648,N_3767);
and U4785 (N_4785,N_3265,N_3735);
nor U4786 (N_4786,N_3374,N_3704);
nor U4787 (N_4787,N_3581,N_3743);
and U4788 (N_4788,N_3174,N_3538);
nor U4789 (N_4789,N_3746,N_3778);
xor U4790 (N_4790,N_3438,N_3065);
and U4791 (N_4791,N_3431,N_3187);
nand U4792 (N_4792,N_3825,N_3473);
and U4793 (N_4793,N_3956,N_3243);
and U4794 (N_4794,N_3390,N_3680);
nand U4795 (N_4795,N_3572,N_3277);
and U4796 (N_4796,N_3717,N_3991);
nor U4797 (N_4797,N_3393,N_3507);
nand U4798 (N_4798,N_3650,N_3072);
xor U4799 (N_4799,N_3278,N_3939);
nor U4800 (N_4800,N_3874,N_3193);
and U4801 (N_4801,N_3561,N_3309);
nor U4802 (N_4802,N_3738,N_3790);
nand U4803 (N_4803,N_3345,N_3472);
nand U4804 (N_4804,N_3278,N_3215);
nand U4805 (N_4805,N_3405,N_3159);
nor U4806 (N_4806,N_3547,N_3800);
or U4807 (N_4807,N_3367,N_3994);
nor U4808 (N_4808,N_3339,N_3772);
nand U4809 (N_4809,N_3313,N_3899);
or U4810 (N_4810,N_3030,N_3448);
or U4811 (N_4811,N_3650,N_3099);
nand U4812 (N_4812,N_3757,N_3368);
nor U4813 (N_4813,N_3641,N_3616);
nand U4814 (N_4814,N_3629,N_3849);
nand U4815 (N_4815,N_3705,N_3656);
nand U4816 (N_4816,N_3247,N_3360);
nor U4817 (N_4817,N_3563,N_3145);
nand U4818 (N_4818,N_3574,N_3605);
and U4819 (N_4819,N_3285,N_3916);
xor U4820 (N_4820,N_3661,N_3056);
or U4821 (N_4821,N_3507,N_3917);
or U4822 (N_4822,N_3639,N_3611);
and U4823 (N_4823,N_3235,N_3147);
nand U4824 (N_4824,N_3589,N_3852);
or U4825 (N_4825,N_3678,N_3805);
or U4826 (N_4826,N_3511,N_3958);
or U4827 (N_4827,N_3294,N_3328);
or U4828 (N_4828,N_3173,N_3259);
and U4829 (N_4829,N_3552,N_3037);
nor U4830 (N_4830,N_3527,N_3710);
xnor U4831 (N_4831,N_3305,N_3025);
nor U4832 (N_4832,N_3694,N_3474);
nor U4833 (N_4833,N_3114,N_3110);
nor U4834 (N_4834,N_3342,N_3991);
and U4835 (N_4835,N_3995,N_3839);
or U4836 (N_4836,N_3823,N_3699);
nor U4837 (N_4837,N_3135,N_3774);
or U4838 (N_4838,N_3336,N_3999);
and U4839 (N_4839,N_3957,N_3480);
nor U4840 (N_4840,N_3392,N_3952);
and U4841 (N_4841,N_3453,N_3704);
nand U4842 (N_4842,N_3427,N_3678);
nor U4843 (N_4843,N_3593,N_3206);
nand U4844 (N_4844,N_3493,N_3738);
or U4845 (N_4845,N_3810,N_3063);
nor U4846 (N_4846,N_3020,N_3244);
nand U4847 (N_4847,N_3852,N_3664);
or U4848 (N_4848,N_3683,N_3236);
xor U4849 (N_4849,N_3609,N_3981);
or U4850 (N_4850,N_3290,N_3503);
xor U4851 (N_4851,N_3355,N_3447);
or U4852 (N_4852,N_3428,N_3124);
and U4853 (N_4853,N_3878,N_3552);
nor U4854 (N_4854,N_3264,N_3982);
or U4855 (N_4855,N_3873,N_3456);
nor U4856 (N_4856,N_3154,N_3627);
or U4857 (N_4857,N_3523,N_3059);
and U4858 (N_4858,N_3843,N_3911);
or U4859 (N_4859,N_3940,N_3524);
nand U4860 (N_4860,N_3568,N_3991);
or U4861 (N_4861,N_3396,N_3417);
nand U4862 (N_4862,N_3744,N_3008);
nand U4863 (N_4863,N_3061,N_3604);
nor U4864 (N_4864,N_3536,N_3718);
nand U4865 (N_4865,N_3073,N_3333);
nor U4866 (N_4866,N_3909,N_3490);
nor U4867 (N_4867,N_3328,N_3529);
nand U4868 (N_4868,N_3584,N_3170);
nand U4869 (N_4869,N_3476,N_3422);
and U4870 (N_4870,N_3230,N_3522);
nand U4871 (N_4871,N_3167,N_3014);
or U4872 (N_4872,N_3833,N_3322);
nor U4873 (N_4873,N_3952,N_3684);
nor U4874 (N_4874,N_3856,N_3496);
xor U4875 (N_4875,N_3139,N_3520);
or U4876 (N_4876,N_3361,N_3509);
and U4877 (N_4877,N_3241,N_3328);
or U4878 (N_4878,N_3671,N_3368);
nor U4879 (N_4879,N_3551,N_3663);
and U4880 (N_4880,N_3702,N_3191);
or U4881 (N_4881,N_3361,N_3746);
nand U4882 (N_4882,N_3474,N_3645);
or U4883 (N_4883,N_3604,N_3845);
nor U4884 (N_4884,N_3742,N_3580);
and U4885 (N_4885,N_3304,N_3568);
nor U4886 (N_4886,N_3200,N_3564);
nand U4887 (N_4887,N_3131,N_3023);
and U4888 (N_4888,N_3310,N_3719);
and U4889 (N_4889,N_3594,N_3864);
nor U4890 (N_4890,N_3300,N_3964);
and U4891 (N_4891,N_3463,N_3170);
nand U4892 (N_4892,N_3158,N_3328);
or U4893 (N_4893,N_3745,N_3384);
or U4894 (N_4894,N_3238,N_3345);
or U4895 (N_4895,N_3014,N_3745);
nor U4896 (N_4896,N_3327,N_3480);
or U4897 (N_4897,N_3803,N_3072);
and U4898 (N_4898,N_3114,N_3465);
or U4899 (N_4899,N_3681,N_3311);
nor U4900 (N_4900,N_3403,N_3029);
nand U4901 (N_4901,N_3524,N_3639);
xnor U4902 (N_4902,N_3277,N_3721);
nor U4903 (N_4903,N_3189,N_3418);
nand U4904 (N_4904,N_3532,N_3442);
and U4905 (N_4905,N_3095,N_3945);
nor U4906 (N_4906,N_3523,N_3851);
or U4907 (N_4907,N_3975,N_3990);
nor U4908 (N_4908,N_3863,N_3814);
nand U4909 (N_4909,N_3985,N_3447);
and U4910 (N_4910,N_3823,N_3565);
nor U4911 (N_4911,N_3721,N_3364);
nand U4912 (N_4912,N_3540,N_3698);
and U4913 (N_4913,N_3798,N_3958);
or U4914 (N_4914,N_3301,N_3655);
nor U4915 (N_4915,N_3919,N_3665);
and U4916 (N_4916,N_3308,N_3004);
xnor U4917 (N_4917,N_3806,N_3767);
xnor U4918 (N_4918,N_3065,N_3842);
nand U4919 (N_4919,N_3013,N_3167);
nor U4920 (N_4920,N_3423,N_3995);
nor U4921 (N_4921,N_3561,N_3873);
nor U4922 (N_4922,N_3356,N_3165);
and U4923 (N_4923,N_3228,N_3591);
and U4924 (N_4924,N_3898,N_3626);
or U4925 (N_4925,N_3837,N_3923);
or U4926 (N_4926,N_3738,N_3387);
nand U4927 (N_4927,N_3926,N_3615);
nor U4928 (N_4928,N_3451,N_3235);
or U4929 (N_4929,N_3534,N_3933);
nand U4930 (N_4930,N_3549,N_3075);
nor U4931 (N_4931,N_3975,N_3873);
nand U4932 (N_4932,N_3920,N_3909);
or U4933 (N_4933,N_3239,N_3643);
nor U4934 (N_4934,N_3599,N_3908);
nor U4935 (N_4935,N_3912,N_3524);
nand U4936 (N_4936,N_3131,N_3912);
or U4937 (N_4937,N_3043,N_3605);
nand U4938 (N_4938,N_3696,N_3338);
and U4939 (N_4939,N_3777,N_3388);
or U4940 (N_4940,N_3722,N_3459);
nor U4941 (N_4941,N_3770,N_3497);
or U4942 (N_4942,N_3567,N_3924);
nor U4943 (N_4943,N_3681,N_3153);
and U4944 (N_4944,N_3007,N_3274);
and U4945 (N_4945,N_3548,N_3430);
nor U4946 (N_4946,N_3297,N_3988);
nand U4947 (N_4947,N_3864,N_3091);
nand U4948 (N_4948,N_3169,N_3021);
nand U4949 (N_4949,N_3626,N_3726);
or U4950 (N_4950,N_3301,N_3800);
xnor U4951 (N_4951,N_3374,N_3202);
nand U4952 (N_4952,N_3132,N_3725);
or U4953 (N_4953,N_3835,N_3726);
nor U4954 (N_4954,N_3913,N_3865);
or U4955 (N_4955,N_3408,N_3704);
nor U4956 (N_4956,N_3029,N_3316);
nor U4957 (N_4957,N_3841,N_3252);
nand U4958 (N_4958,N_3952,N_3855);
nand U4959 (N_4959,N_3213,N_3907);
or U4960 (N_4960,N_3987,N_3975);
nand U4961 (N_4961,N_3878,N_3886);
nor U4962 (N_4962,N_3792,N_3853);
nand U4963 (N_4963,N_3787,N_3945);
nand U4964 (N_4964,N_3951,N_3271);
or U4965 (N_4965,N_3785,N_3456);
and U4966 (N_4966,N_3012,N_3119);
nor U4967 (N_4967,N_3478,N_3064);
nor U4968 (N_4968,N_3269,N_3052);
xor U4969 (N_4969,N_3715,N_3681);
and U4970 (N_4970,N_3070,N_3891);
or U4971 (N_4971,N_3314,N_3170);
nand U4972 (N_4972,N_3263,N_3654);
and U4973 (N_4973,N_3337,N_3320);
nor U4974 (N_4974,N_3448,N_3820);
xor U4975 (N_4975,N_3709,N_3058);
nand U4976 (N_4976,N_3672,N_3525);
and U4977 (N_4977,N_3258,N_3709);
and U4978 (N_4978,N_3193,N_3271);
and U4979 (N_4979,N_3170,N_3759);
and U4980 (N_4980,N_3477,N_3894);
and U4981 (N_4981,N_3693,N_3208);
or U4982 (N_4982,N_3707,N_3686);
and U4983 (N_4983,N_3575,N_3321);
and U4984 (N_4984,N_3645,N_3351);
xor U4985 (N_4985,N_3785,N_3902);
or U4986 (N_4986,N_3184,N_3085);
and U4987 (N_4987,N_3006,N_3391);
nand U4988 (N_4988,N_3189,N_3149);
nand U4989 (N_4989,N_3300,N_3774);
and U4990 (N_4990,N_3979,N_3999);
nor U4991 (N_4991,N_3467,N_3066);
nor U4992 (N_4992,N_3224,N_3537);
and U4993 (N_4993,N_3523,N_3981);
nor U4994 (N_4994,N_3668,N_3500);
or U4995 (N_4995,N_3771,N_3722);
and U4996 (N_4996,N_3919,N_3062);
nor U4997 (N_4997,N_3039,N_3435);
nand U4998 (N_4998,N_3918,N_3135);
nor U4999 (N_4999,N_3076,N_3767);
or UO_0 (O_0,N_4309,N_4366);
nand UO_1 (O_1,N_4654,N_4134);
nand UO_2 (O_2,N_4140,N_4641);
or UO_3 (O_3,N_4264,N_4041);
nand UO_4 (O_4,N_4006,N_4777);
or UO_5 (O_5,N_4093,N_4231);
nor UO_6 (O_6,N_4016,N_4298);
nand UO_7 (O_7,N_4084,N_4333);
nand UO_8 (O_8,N_4306,N_4353);
and UO_9 (O_9,N_4574,N_4444);
nand UO_10 (O_10,N_4060,N_4200);
and UO_11 (O_11,N_4845,N_4705);
nand UO_12 (O_12,N_4086,N_4288);
nor UO_13 (O_13,N_4282,N_4014);
nor UO_14 (O_14,N_4431,N_4585);
nand UO_15 (O_15,N_4927,N_4983);
nand UO_16 (O_16,N_4879,N_4092);
nor UO_17 (O_17,N_4906,N_4109);
and UO_18 (O_18,N_4963,N_4580);
nor UO_19 (O_19,N_4368,N_4382);
nand UO_20 (O_20,N_4550,N_4136);
or UO_21 (O_21,N_4937,N_4647);
or UO_22 (O_22,N_4496,N_4481);
nand UO_23 (O_23,N_4950,N_4301);
nand UO_24 (O_24,N_4532,N_4812);
nor UO_25 (O_25,N_4455,N_4988);
nor UO_26 (O_26,N_4024,N_4478);
and UO_27 (O_27,N_4652,N_4113);
and UO_28 (O_28,N_4827,N_4752);
or UO_29 (O_29,N_4671,N_4278);
or UO_30 (O_30,N_4248,N_4543);
and UO_31 (O_31,N_4155,N_4450);
and UO_32 (O_32,N_4596,N_4731);
nand UO_33 (O_33,N_4957,N_4861);
or UO_34 (O_34,N_4074,N_4876);
and UO_35 (O_35,N_4748,N_4848);
and UO_36 (O_36,N_4249,N_4324);
nor UO_37 (O_37,N_4243,N_4501);
nor UO_38 (O_38,N_4164,N_4939);
and UO_39 (O_39,N_4000,N_4530);
and UO_40 (O_40,N_4008,N_4192);
nand UO_41 (O_41,N_4507,N_4296);
and UO_42 (O_42,N_4573,N_4430);
nor UO_43 (O_43,N_4858,N_4975);
nor UO_44 (O_44,N_4290,N_4971);
nor UO_45 (O_45,N_4911,N_4406);
and UO_46 (O_46,N_4807,N_4184);
xnor UO_47 (O_47,N_4468,N_4201);
nor UO_48 (O_48,N_4304,N_4685);
and UO_49 (O_49,N_4106,N_4261);
and UO_50 (O_50,N_4889,N_4300);
nor UO_51 (O_51,N_4629,N_4129);
and UO_52 (O_52,N_4826,N_4271);
nand UO_53 (O_53,N_4133,N_4616);
nand UO_54 (O_54,N_4214,N_4589);
nor UO_55 (O_55,N_4851,N_4797);
and UO_56 (O_56,N_4057,N_4378);
nand UO_57 (O_57,N_4563,N_4438);
nor UO_58 (O_58,N_4757,N_4101);
or UO_59 (O_59,N_4479,N_4972);
xor UO_60 (O_60,N_4979,N_4707);
or UO_61 (O_61,N_4454,N_4985);
and UO_62 (O_62,N_4664,N_4880);
xnor UO_63 (O_63,N_4929,N_4974);
xnor UO_64 (O_64,N_4286,N_4055);
and UO_65 (O_65,N_4349,N_4559);
xnor UO_66 (O_66,N_4970,N_4577);
nand UO_67 (O_67,N_4233,N_4718);
and UO_68 (O_68,N_4095,N_4319);
or UO_69 (O_69,N_4295,N_4066);
or UO_70 (O_70,N_4071,N_4139);
nand UO_71 (O_71,N_4809,N_4330);
or UO_72 (O_72,N_4502,N_4676);
nand UO_73 (O_73,N_4508,N_4512);
nor UO_74 (O_74,N_4383,N_4365);
nor UO_75 (O_75,N_4829,N_4299);
or UO_76 (O_76,N_4036,N_4379);
and UO_77 (O_77,N_4566,N_4535);
nand UO_78 (O_78,N_4599,N_4749);
and UO_79 (O_79,N_4067,N_4254);
or UO_80 (O_80,N_4608,N_4750);
xnor UO_81 (O_81,N_4340,N_4302);
nor UO_82 (O_82,N_4514,N_4400);
nor UO_83 (O_83,N_4766,N_4409);
or UO_84 (O_84,N_4314,N_4740);
and UO_85 (O_85,N_4185,N_4790);
and UO_86 (O_86,N_4989,N_4811);
or UO_87 (O_87,N_4980,N_4097);
nor UO_88 (O_88,N_4619,N_4361);
nand UO_89 (O_89,N_4423,N_4359);
and UO_90 (O_90,N_4061,N_4645);
or UO_91 (O_91,N_4021,N_4449);
and UO_92 (O_92,N_4149,N_4236);
or UO_93 (O_93,N_4914,N_4999);
or UO_94 (O_94,N_4590,N_4403);
nand UO_95 (O_95,N_4064,N_4625);
nor UO_96 (O_96,N_4661,N_4161);
or UO_97 (O_97,N_4334,N_4698);
nand UO_98 (O_98,N_4808,N_4903);
nor UO_99 (O_99,N_4011,N_4251);
nor UO_100 (O_100,N_4904,N_4928);
or UO_101 (O_101,N_4193,N_4742);
and UO_102 (O_102,N_4504,N_4405);
or UO_103 (O_103,N_4572,N_4537);
and UO_104 (O_104,N_4956,N_4273);
nor UO_105 (O_105,N_4246,N_4902);
nand UO_106 (O_106,N_4126,N_4331);
and UO_107 (O_107,N_4962,N_4965);
xnor UO_108 (O_108,N_4156,N_4500);
and UO_109 (O_109,N_4894,N_4402);
and UO_110 (O_110,N_4367,N_4804);
or UO_111 (O_111,N_4217,N_4649);
nor UO_112 (O_112,N_4047,N_4210);
nand UO_113 (O_113,N_4866,N_4491);
nor UO_114 (O_114,N_4469,N_4393);
and UO_115 (O_115,N_4555,N_4706);
nor UO_116 (O_116,N_4597,N_4646);
and UO_117 (O_117,N_4745,N_4801);
nand UO_118 (O_118,N_4639,N_4862);
nand UO_119 (O_119,N_4173,N_4490);
nand UO_120 (O_120,N_4453,N_4044);
nor UO_121 (O_121,N_4341,N_4255);
xnor UO_122 (O_122,N_4396,N_4056);
xnor UO_123 (O_123,N_4815,N_4374);
and UO_124 (O_124,N_4571,N_4798);
or UO_125 (O_125,N_4051,N_4351);
nand UO_126 (O_126,N_4179,N_4096);
or UO_127 (O_127,N_4470,N_4235);
or UO_128 (O_128,N_4819,N_4747);
nor UO_129 (O_129,N_4683,N_4059);
or UO_130 (O_130,N_4289,N_4709);
xor UO_131 (O_131,N_4034,N_4332);
nor UO_132 (O_132,N_4864,N_4763);
or UO_133 (O_133,N_4125,N_4803);
nand UO_134 (O_134,N_4040,N_4792);
or UO_135 (O_135,N_4076,N_4445);
or UO_136 (O_136,N_4699,N_4744);
nor UO_137 (O_137,N_4219,N_4690);
or UO_138 (O_138,N_4420,N_4098);
and UO_139 (O_139,N_4814,N_4380);
and UO_140 (O_140,N_4322,N_4620);
and UO_141 (O_141,N_4369,N_4081);
or UO_142 (O_142,N_4778,N_4020);
or UO_143 (O_143,N_4658,N_4198);
nand UO_144 (O_144,N_4327,N_4544);
xor UO_145 (O_145,N_4528,N_4886);
and UO_146 (O_146,N_4575,N_4952);
or UO_147 (O_147,N_4818,N_4593);
or UO_148 (O_148,N_4693,N_4739);
or UO_149 (O_149,N_4913,N_4499);
xnor UO_150 (O_150,N_4068,N_4591);
or UO_151 (O_151,N_4837,N_4996);
and UO_152 (O_152,N_4472,N_4230);
or UO_153 (O_153,N_4005,N_4517);
and UO_154 (O_154,N_4922,N_4653);
and UO_155 (O_155,N_4460,N_4579);
nand UO_156 (O_156,N_4208,N_4525);
and UO_157 (O_157,N_4700,N_4531);
or UO_158 (O_158,N_4694,N_4515);
nand UO_159 (O_159,N_4119,N_4923);
xnor UO_160 (O_160,N_4428,N_4411);
nor UO_161 (O_161,N_4935,N_4488);
nor UO_162 (O_162,N_4657,N_4174);
nand UO_163 (O_163,N_4849,N_4642);
nand UO_164 (O_164,N_4216,N_4949);
or UO_165 (O_165,N_4211,N_4343);
nor UO_166 (O_166,N_4978,N_4840);
or UO_167 (O_167,N_4542,N_4723);
and UO_168 (O_168,N_4726,N_4142);
nor UO_169 (O_169,N_4900,N_4943);
and UO_170 (O_170,N_4358,N_4838);
nor UO_171 (O_171,N_4162,N_4955);
and UO_172 (O_172,N_4265,N_4905);
and UO_173 (O_173,N_4189,N_4678);
and UO_174 (O_174,N_4408,N_4388);
and UO_175 (O_175,N_4874,N_4519);
or UO_176 (O_176,N_4263,N_4407);
nor UO_177 (O_177,N_4743,N_4222);
and UO_178 (O_178,N_4667,N_4242);
nand UO_179 (O_179,N_4342,N_4973);
and UO_180 (O_180,N_4924,N_4520);
nand UO_181 (O_181,N_4982,N_4634);
nand UO_182 (O_182,N_4822,N_4026);
nor UO_183 (O_183,N_4885,N_4713);
or UO_184 (O_184,N_4839,N_4029);
or UO_185 (O_185,N_4169,N_4780);
and UO_186 (O_186,N_4116,N_4735);
nor UO_187 (O_187,N_4004,N_4268);
or UO_188 (O_188,N_4147,N_4033);
or UO_189 (O_189,N_4651,N_4633);
nor UO_190 (O_190,N_4476,N_4392);
nor UO_191 (O_191,N_4746,N_4830);
nor UO_192 (O_192,N_4285,N_4486);
nor UO_193 (O_193,N_4281,N_4225);
and UO_194 (O_194,N_4387,N_4099);
and UO_195 (O_195,N_4805,N_4677);
nor UO_196 (O_196,N_4613,N_4753);
nand UO_197 (O_197,N_4487,N_4719);
and UO_198 (O_198,N_4480,N_4774);
and UO_199 (O_199,N_4370,N_4650);
or UO_200 (O_200,N_4586,N_4357);
nor UO_201 (O_201,N_4120,N_4931);
nor UO_202 (O_202,N_4053,N_4666);
nand UO_203 (O_203,N_4729,N_4522);
and UO_204 (O_204,N_4461,N_4199);
and UO_205 (O_205,N_4578,N_4776);
nor UO_206 (O_206,N_4262,N_4323);
nor UO_207 (O_207,N_4190,N_4831);
or UO_208 (O_208,N_4562,N_4930);
nor UO_209 (O_209,N_4197,N_4028);
nor UO_210 (O_210,N_4786,N_4648);
and UO_211 (O_211,N_4123,N_4703);
nand UO_212 (O_212,N_4524,N_4631);
nand UO_213 (O_213,N_4277,N_4860);
nand UO_214 (O_214,N_4115,N_4137);
or UO_215 (O_215,N_4817,N_4335);
nor UO_216 (O_216,N_4019,N_4321);
or UO_217 (O_217,N_4172,N_4505);
nor UO_218 (O_218,N_4617,N_4463);
and UO_219 (O_219,N_4088,N_4075);
nor UO_220 (O_220,N_4435,N_4381);
or UO_221 (O_221,N_4283,N_4609);
nor UO_222 (O_222,N_4954,N_4412);
nand UO_223 (O_223,N_4781,N_4362);
and UO_224 (O_224,N_4503,N_4727);
or UO_225 (O_225,N_4439,N_4764);
xnor UO_226 (O_226,N_4390,N_4284);
or UO_227 (O_227,N_4204,N_4738);
nand UO_228 (O_228,N_4857,N_4841);
and UO_229 (O_229,N_4462,N_4576);
nand UO_230 (O_230,N_4269,N_4344);
nand UO_231 (O_231,N_4604,N_4953);
nand UO_232 (O_232,N_4675,N_4176);
and UO_233 (O_233,N_4112,N_4656);
and UO_234 (O_234,N_4663,N_4234);
nor UO_235 (O_235,N_4336,N_4938);
nor UO_236 (O_236,N_4570,N_4104);
nor UO_237 (O_237,N_4910,N_4375);
nand UO_238 (O_238,N_4058,N_4662);
or UO_239 (O_239,N_4846,N_4612);
and UO_240 (O_240,N_4003,N_4784);
or UO_241 (O_241,N_4205,N_4276);
and UO_242 (O_242,N_4884,N_4356);
nor UO_243 (O_243,N_4206,N_4032);
xor UO_244 (O_244,N_4796,N_4847);
xnor UO_245 (O_245,N_4659,N_4135);
nor UO_246 (O_246,N_4384,N_4391);
or UO_247 (O_247,N_4813,N_4087);
or UO_248 (O_248,N_4888,N_4665);
or UO_249 (O_249,N_4511,N_4178);
nand UO_250 (O_250,N_4352,N_4926);
nand UO_251 (O_251,N_4090,N_4548);
or UO_252 (O_252,N_4602,N_4377);
nor UO_253 (O_253,N_4626,N_4867);
or UO_254 (O_254,N_4001,N_4079);
nor UO_255 (O_255,N_4364,N_4668);
or UO_256 (O_256,N_4475,N_4187);
or UO_257 (O_257,N_4315,N_4509);
nand UO_258 (O_258,N_4869,N_4892);
or UO_259 (O_259,N_4681,N_4043);
and UO_260 (O_260,N_4132,N_4958);
nand UO_261 (O_261,N_4794,N_4437);
or UO_262 (O_262,N_4168,N_4583);
nand UO_263 (O_263,N_4760,N_4121);
or UO_264 (O_264,N_4695,N_4761);
nor UO_265 (O_265,N_4877,N_4909);
nor UO_266 (O_266,N_4640,N_4326);
or UO_267 (O_267,N_4027,N_4077);
or UO_268 (O_268,N_4603,N_4799);
and UO_269 (O_269,N_4605,N_4997);
or UO_270 (O_270,N_4751,N_4145);
nand UO_271 (O_271,N_4239,N_4800);
nor UO_272 (O_272,N_4547,N_4130);
nor UO_273 (O_273,N_4274,N_4151);
or UO_274 (O_274,N_4976,N_4795);
or UO_275 (O_275,N_4933,N_4226);
nand UO_276 (O_276,N_4674,N_4373);
nor UO_277 (O_277,N_4218,N_4538);
nor UO_278 (O_278,N_4832,N_4360);
and UO_279 (O_279,N_4477,N_4404);
and UO_280 (O_280,N_4863,N_4539);
xor UO_281 (O_281,N_4714,N_4756);
nor UO_282 (O_282,N_4768,N_4049);
nor UO_283 (O_283,N_4898,N_4635);
or UO_284 (O_284,N_4934,N_4918);
or UO_285 (O_285,N_4836,N_4793);
and UO_286 (O_286,N_4755,N_4990);
nand UO_287 (O_287,N_4679,N_4506);
and UO_288 (O_288,N_4039,N_4701);
nor UO_289 (O_289,N_4157,N_4312);
and UO_290 (O_290,N_4720,N_4941);
and UO_291 (O_291,N_4995,N_4417);
nand UO_292 (O_292,N_4765,N_4587);
and UO_293 (O_293,N_4080,N_4844);
nor UO_294 (O_294,N_4842,N_4399);
nand UO_295 (O_295,N_4146,N_4223);
and UO_296 (O_296,N_4940,N_4891);
nand UO_297 (O_297,N_4536,N_4859);
or UO_298 (O_298,N_4592,N_4181);
nor UO_299 (O_299,N_4546,N_4611);
or UO_300 (O_300,N_4188,N_4452);
nor UO_301 (O_301,N_4177,N_4769);
or UO_302 (O_302,N_4561,N_4521);
nor UO_303 (O_303,N_4883,N_4257);
or UO_304 (O_304,N_4584,N_4144);
xnor UO_305 (O_305,N_4969,N_4318);
or UO_306 (O_306,N_4569,N_4854);
or UO_307 (O_307,N_4946,N_4986);
nor UO_308 (O_308,N_4824,N_4287);
or UO_309 (O_309,N_4948,N_4510);
nand UO_310 (O_310,N_4007,N_4758);
and UO_311 (O_311,N_4091,N_4191);
nand UO_312 (O_312,N_4899,N_4672);
nor UO_313 (O_313,N_4637,N_4473);
or UO_314 (O_314,N_4893,N_4175);
or UO_315 (O_315,N_4457,N_4907);
xnor UO_316 (O_316,N_4912,N_4682);
nor UO_317 (O_317,N_4103,N_4163);
nor UO_318 (O_318,N_4977,N_4686);
nand UO_319 (O_319,N_4991,N_4541);
and UO_320 (O_320,N_4410,N_4426);
xnor UO_321 (O_321,N_4458,N_4467);
xor UO_322 (O_322,N_4644,N_4771);
nand UO_323 (O_323,N_4078,N_4715);
nand UO_324 (O_324,N_4882,N_4256);
or UO_325 (O_325,N_4209,N_4716);
nand UO_326 (O_326,N_4670,N_4887);
nor UO_327 (O_327,N_4878,N_4338);
nor UO_328 (O_328,N_4310,N_4856);
and UO_329 (O_329,N_4712,N_4048);
and UO_330 (O_330,N_4182,N_4582);
or UO_331 (O_331,N_4741,N_4557);
or UO_332 (O_332,N_4691,N_4702);
and UO_333 (O_333,N_4346,N_4456);
or UO_334 (O_334,N_4896,N_4489);
nor UO_335 (O_335,N_4624,N_4916);
nand UO_336 (O_336,N_4855,N_4871);
or UO_337 (O_337,N_4643,N_4260);
or UO_338 (O_338,N_4451,N_4474);
nand UO_339 (O_339,N_4994,N_4529);
nor UO_340 (O_340,N_4221,N_4944);
xnor UO_341 (O_341,N_4967,N_4031);
and UO_342 (O_342,N_4442,N_4237);
and UO_343 (O_343,N_4921,N_4317);
nor UO_344 (O_344,N_4207,N_4238);
and UO_345 (O_345,N_4636,N_4297);
or UO_346 (O_346,N_4037,N_4363);
or UO_347 (O_347,N_4012,N_4728);
nor UO_348 (O_348,N_4416,N_4992);
nand UO_349 (O_349,N_4013,N_4063);
or UO_350 (O_350,N_4919,N_4413);
or UO_351 (O_351,N_4072,N_4783);
or UO_352 (O_352,N_4770,N_4114);
and UO_353 (O_353,N_4865,N_4773);
nand UO_354 (O_354,N_4291,N_4434);
or UO_355 (O_355,N_4419,N_4704);
or UO_356 (O_356,N_4038,N_4152);
nor UO_357 (O_357,N_4117,N_4951);
or UO_358 (O_358,N_4984,N_4482);
or UO_359 (O_359,N_4447,N_4843);
nor UO_360 (O_360,N_4212,N_4901);
or UO_361 (O_361,N_4549,N_4725);
and UO_362 (O_362,N_4881,N_4272);
and UO_363 (O_363,N_4607,N_4788);
or UO_364 (O_364,N_4443,N_4551);
or UO_365 (O_365,N_4228,N_4810);
xnor UO_366 (O_366,N_4229,N_4158);
nor UO_367 (O_367,N_4534,N_4556);
nand UO_368 (O_368,N_4736,N_4166);
nor UO_369 (O_369,N_4429,N_4372);
and UO_370 (O_370,N_4552,N_4960);
nor UO_371 (O_371,N_4545,N_4852);
and UO_372 (O_372,N_4348,N_4968);
and UO_373 (O_373,N_4554,N_4025);
and UO_374 (O_374,N_4385,N_4108);
nor UO_375 (O_375,N_4961,N_4615);
nand UO_376 (O_376,N_4094,N_4945);
nor UO_377 (O_377,N_4835,N_4523);
nor UO_378 (O_378,N_4073,N_4386);
xor UO_379 (O_379,N_4540,N_4823);
nor UO_380 (O_380,N_4244,N_4623);
nand UO_381 (O_381,N_4565,N_4942);
and UO_382 (O_382,N_4621,N_4526);
and UO_383 (O_383,N_4313,N_4932);
nor UO_384 (O_384,N_4292,N_4376);
or UO_385 (O_385,N_4227,N_4567);
nand UO_386 (O_386,N_4062,N_4981);
or UO_387 (O_387,N_4303,N_4240);
nor UO_388 (O_388,N_4015,N_4339);
or UO_389 (O_389,N_4669,N_4131);
xor UO_390 (O_390,N_4280,N_4594);
nor UO_391 (O_391,N_4082,N_4389);
nand UO_392 (O_392,N_4337,N_4733);
or UO_393 (O_393,N_4195,N_4833);
nor UO_394 (O_394,N_4987,N_4558);
nand UO_395 (O_395,N_4070,N_4448);
nand UO_396 (O_396,N_4259,N_4202);
nor UO_397 (O_397,N_4820,N_4107);
or UO_398 (O_398,N_4418,N_4002);
nand UO_399 (O_399,N_4414,N_4085);
and UO_400 (O_400,N_4253,N_4966);
and UO_401 (O_401,N_4203,N_4627);
nor UO_402 (O_402,N_4266,N_4687);
nor UO_403 (O_403,N_4601,N_4010);
nand UO_404 (O_404,N_4688,N_4440);
nor UO_405 (O_405,N_4320,N_4875);
nand UO_406 (O_406,N_4150,N_4754);
nor UO_407 (O_407,N_4908,N_4828);
nand UO_408 (O_408,N_4371,N_4581);
or UO_409 (O_409,N_4915,N_4127);
nand UO_410 (O_410,N_4267,N_4684);
nand UO_411 (O_411,N_4345,N_4279);
or UO_412 (O_412,N_4638,N_4895);
nor UO_413 (O_413,N_4459,N_4495);
nand UO_414 (O_414,N_4632,N_4083);
nand UO_415 (O_415,N_4825,N_4293);
and UO_416 (O_416,N_4308,N_4270);
or UO_417 (O_417,N_4355,N_4610);
or UO_418 (O_418,N_4167,N_4089);
nor UO_419 (O_419,N_4250,N_4446);
and UO_420 (O_420,N_4153,N_4568);
or UO_421 (O_421,N_4936,N_4220);
nand UO_422 (O_422,N_4154,N_4821);
xnor UO_423 (O_423,N_4328,N_4258);
or UO_424 (O_424,N_4050,N_4850);
nor UO_425 (O_425,N_4311,N_4595);
and UO_426 (O_426,N_4433,N_4213);
nand UO_427 (O_427,N_4141,N_4787);
and UO_428 (O_428,N_4425,N_4630);
nand UO_429 (O_429,N_4527,N_4159);
and UO_430 (O_430,N_4959,N_4180);
xnor UO_431 (O_431,N_4102,N_4917);
xnor UO_432 (O_432,N_4588,N_4232);
or UO_433 (O_433,N_4553,N_4516);
nand UO_434 (O_434,N_4680,N_4779);
nor UO_435 (O_435,N_4215,N_4484);
and UO_436 (O_436,N_4465,N_4009);
and UO_437 (O_437,N_4816,N_4100);
or UO_438 (O_438,N_4673,N_4689);
and UO_439 (O_439,N_4294,N_4105);
nand UO_440 (O_440,N_4394,N_4485);
or UO_441 (O_441,N_4325,N_4660);
or UO_442 (O_442,N_4498,N_4247);
and UO_443 (O_443,N_4692,N_4354);
or UO_444 (O_444,N_4998,N_4920);
and UO_445 (O_445,N_4069,N_4186);
nor UO_446 (O_446,N_4427,N_4110);
xnor UO_447 (O_447,N_4993,N_4035);
or UO_448 (O_448,N_4118,N_4853);
or UO_449 (O_449,N_4436,N_4415);
or UO_450 (O_450,N_4802,N_4018);
nand UO_451 (O_451,N_4023,N_4350);
xnor UO_452 (O_452,N_4054,N_4518);
and UO_453 (O_453,N_4697,N_4432);
nor UO_454 (O_454,N_4148,N_4045);
or UO_455 (O_455,N_4772,N_4622);
and UO_456 (O_456,N_4614,N_4492);
nand UO_457 (O_457,N_4165,N_4708);
or UO_458 (O_458,N_4628,N_4897);
and UO_459 (O_459,N_4030,N_4052);
nor UO_460 (O_460,N_4398,N_4759);
and UO_461 (O_461,N_4724,N_4065);
and UO_462 (O_462,N_4128,N_4422);
and UO_463 (O_463,N_4834,N_4710);
or UO_464 (O_464,N_4873,N_4767);
or UO_465 (O_465,N_4722,N_4170);
nand UO_466 (O_466,N_4789,N_4046);
nor UO_467 (O_467,N_4122,N_4483);
and UO_468 (O_468,N_4316,N_4245);
and UO_469 (O_469,N_4868,N_4890);
nand UO_470 (O_470,N_4618,N_4925);
nand UO_471 (O_471,N_4241,N_4964);
or UO_472 (O_472,N_4732,N_4513);
nor UO_473 (O_473,N_4171,N_4947);
nor UO_474 (O_474,N_4497,N_4196);
or UO_475 (O_475,N_4401,N_4307);
nand UO_476 (O_476,N_4600,N_4183);
and UO_477 (O_477,N_4017,N_4421);
nand UO_478 (O_478,N_4791,N_4762);
and UO_479 (O_479,N_4042,N_4252);
nand UO_480 (O_480,N_4655,N_4870);
or UO_481 (O_481,N_4395,N_4022);
and UO_482 (O_482,N_4737,N_4466);
nor UO_483 (O_483,N_4143,N_4194);
nor UO_484 (O_484,N_4606,N_4124);
or UO_485 (O_485,N_4275,N_4734);
and UO_486 (O_486,N_4160,N_4721);
or UO_487 (O_487,N_4397,N_4441);
nor UO_488 (O_488,N_4717,N_4711);
nor UO_489 (O_489,N_4775,N_4471);
or UO_490 (O_490,N_4329,N_4560);
nand UO_491 (O_491,N_4598,N_4533);
nor UO_492 (O_492,N_4493,N_4730);
or UO_493 (O_493,N_4305,N_4347);
nor UO_494 (O_494,N_4494,N_4782);
xnor UO_495 (O_495,N_4138,N_4464);
and UO_496 (O_496,N_4872,N_4564);
and UO_497 (O_497,N_4806,N_4424);
or UO_498 (O_498,N_4696,N_4785);
xor UO_499 (O_499,N_4224,N_4111);
and UO_500 (O_500,N_4804,N_4637);
nor UO_501 (O_501,N_4615,N_4440);
or UO_502 (O_502,N_4935,N_4618);
and UO_503 (O_503,N_4861,N_4377);
and UO_504 (O_504,N_4405,N_4533);
nand UO_505 (O_505,N_4512,N_4087);
or UO_506 (O_506,N_4634,N_4448);
and UO_507 (O_507,N_4552,N_4823);
xnor UO_508 (O_508,N_4420,N_4231);
and UO_509 (O_509,N_4199,N_4640);
nand UO_510 (O_510,N_4085,N_4940);
and UO_511 (O_511,N_4579,N_4464);
and UO_512 (O_512,N_4356,N_4864);
or UO_513 (O_513,N_4980,N_4555);
and UO_514 (O_514,N_4831,N_4040);
nand UO_515 (O_515,N_4211,N_4920);
and UO_516 (O_516,N_4842,N_4257);
or UO_517 (O_517,N_4016,N_4617);
and UO_518 (O_518,N_4342,N_4492);
nand UO_519 (O_519,N_4119,N_4889);
or UO_520 (O_520,N_4530,N_4434);
nor UO_521 (O_521,N_4062,N_4724);
or UO_522 (O_522,N_4835,N_4391);
xor UO_523 (O_523,N_4870,N_4967);
nor UO_524 (O_524,N_4494,N_4080);
xnor UO_525 (O_525,N_4817,N_4911);
nor UO_526 (O_526,N_4123,N_4790);
and UO_527 (O_527,N_4043,N_4606);
or UO_528 (O_528,N_4764,N_4575);
or UO_529 (O_529,N_4806,N_4303);
or UO_530 (O_530,N_4214,N_4185);
nand UO_531 (O_531,N_4635,N_4837);
nor UO_532 (O_532,N_4752,N_4791);
or UO_533 (O_533,N_4741,N_4055);
nor UO_534 (O_534,N_4289,N_4427);
or UO_535 (O_535,N_4397,N_4480);
nand UO_536 (O_536,N_4622,N_4163);
and UO_537 (O_537,N_4527,N_4356);
or UO_538 (O_538,N_4232,N_4571);
nand UO_539 (O_539,N_4876,N_4638);
nor UO_540 (O_540,N_4032,N_4286);
and UO_541 (O_541,N_4914,N_4784);
nand UO_542 (O_542,N_4254,N_4114);
or UO_543 (O_543,N_4053,N_4726);
nand UO_544 (O_544,N_4105,N_4730);
and UO_545 (O_545,N_4663,N_4809);
and UO_546 (O_546,N_4233,N_4736);
nor UO_547 (O_547,N_4556,N_4301);
or UO_548 (O_548,N_4490,N_4958);
or UO_549 (O_549,N_4860,N_4994);
and UO_550 (O_550,N_4600,N_4060);
and UO_551 (O_551,N_4732,N_4232);
xor UO_552 (O_552,N_4450,N_4103);
or UO_553 (O_553,N_4716,N_4778);
and UO_554 (O_554,N_4291,N_4166);
nor UO_555 (O_555,N_4680,N_4972);
and UO_556 (O_556,N_4731,N_4132);
nor UO_557 (O_557,N_4520,N_4309);
nor UO_558 (O_558,N_4681,N_4471);
nor UO_559 (O_559,N_4684,N_4985);
xnor UO_560 (O_560,N_4961,N_4251);
nor UO_561 (O_561,N_4801,N_4933);
nor UO_562 (O_562,N_4600,N_4365);
nand UO_563 (O_563,N_4656,N_4141);
and UO_564 (O_564,N_4862,N_4293);
and UO_565 (O_565,N_4089,N_4018);
and UO_566 (O_566,N_4742,N_4478);
nand UO_567 (O_567,N_4978,N_4564);
or UO_568 (O_568,N_4466,N_4621);
and UO_569 (O_569,N_4569,N_4594);
or UO_570 (O_570,N_4145,N_4277);
or UO_571 (O_571,N_4343,N_4062);
or UO_572 (O_572,N_4565,N_4648);
nand UO_573 (O_573,N_4629,N_4570);
nand UO_574 (O_574,N_4255,N_4631);
nor UO_575 (O_575,N_4238,N_4429);
nand UO_576 (O_576,N_4473,N_4789);
nor UO_577 (O_577,N_4009,N_4742);
and UO_578 (O_578,N_4844,N_4887);
nand UO_579 (O_579,N_4573,N_4052);
nand UO_580 (O_580,N_4601,N_4689);
or UO_581 (O_581,N_4691,N_4816);
nand UO_582 (O_582,N_4533,N_4903);
and UO_583 (O_583,N_4778,N_4759);
nor UO_584 (O_584,N_4676,N_4975);
nand UO_585 (O_585,N_4679,N_4984);
or UO_586 (O_586,N_4672,N_4628);
and UO_587 (O_587,N_4112,N_4405);
xor UO_588 (O_588,N_4866,N_4416);
nand UO_589 (O_589,N_4751,N_4206);
and UO_590 (O_590,N_4283,N_4280);
nor UO_591 (O_591,N_4448,N_4815);
and UO_592 (O_592,N_4390,N_4403);
nor UO_593 (O_593,N_4517,N_4756);
and UO_594 (O_594,N_4345,N_4783);
or UO_595 (O_595,N_4357,N_4864);
or UO_596 (O_596,N_4064,N_4612);
nor UO_597 (O_597,N_4147,N_4901);
and UO_598 (O_598,N_4159,N_4374);
or UO_599 (O_599,N_4805,N_4301);
or UO_600 (O_600,N_4584,N_4419);
and UO_601 (O_601,N_4595,N_4106);
nor UO_602 (O_602,N_4898,N_4529);
and UO_603 (O_603,N_4557,N_4766);
and UO_604 (O_604,N_4387,N_4990);
nor UO_605 (O_605,N_4450,N_4380);
nand UO_606 (O_606,N_4939,N_4851);
nand UO_607 (O_607,N_4970,N_4879);
nand UO_608 (O_608,N_4608,N_4123);
nand UO_609 (O_609,N_4085,N_4534);
nor UO_610 (O_610,N_4788,N_4139);
nand UO_611 (O_611,N_4135,N_4265);
or UO_612 (O_612,N_4330,N_4184);
nor UO_613 (O_613,N_4515,N_4707);
and UO_614 (O_614,N_4400,N_4547);
nor UO_615 (O_615,N_4380,N_4473);
or UO_616 (O_616,N_4115,N_4803);
nor UO_617 (O_617,N_4831,N_4941);
and UO_618 (O_618,N_4685,N_4334);
nand UO_619 (O_619,N_4741,N_4161);
nor UO_620 (O_620,N_4852,N_4296);
nand UO_621 (O_621,N_4036,N_4972);
xor UO_622 (O_622,N_4493,N_4557);
nand UO_623 (O_623,N_4180,N_4513);
or UO_624 (O_624,N_4008,N_4158);
nor UO_625 (O_625,N_4866,N_4396);
nor UO_626 (O_626,N_4489,N_4421);
and UO_627 (O_627,N_4210,N_4135);
or UO_628 (O_628,N_4696,N_4732);
and UO_629 (O_629,N_4542,N_4482);
nand UO_630 (O_630,N_4016,N_4563);
nor UO_631 (O_631,N_4495,N_4470);
nand UO_632 (O_632,N_4616,N_4487);
and UO_633 (O_633,N_4118,N_4495);
and UO_634 (O_634,N_4715,N_4388);
nor UO_635 (O_635,N_4041,N_4753);
and UO_636 (O_636,N_4741,N_4327);
or UO_637 (O_637,N_4285,N_4014);
nor UO_638 (O_638,N_4877,N_4013);
nor UO_639 (O_639,N_4752,N_4383);
and UO_640 (O_640,N_4840,N_4330);
nor UO_641 (O_641,N_4775,N_4792);
nor UO_642 (O_642,N_4811,N_4041);
nand UO_643 (O_643,N_4416,N_4420);
nand UO_644 (O_644,N_4521,N_4458);
nand UO_645 (O_645,N_4410,N_4771);
nand UO_646 (O_646,N_4076,N_4867);
nand UO_647 (O_647,N_4334,N_4216);
or UO_648 (O_648,N_4423,N_4557);
or UO_649 (O_649,N_4279,N_4377);
nand UO_650 (O_650,N_4496,N_4343);
or UO_651 (O_651,N_4158,N_4084);
or UO_652 (O_652,N_4142,N_4036);
nor UO_653 (O_653,N_4495,N_4802);
nand UO_654 (O_654,N_4944,N_4437);
and UO_655 (O_655,N_4194,N_4448);
and UO_656 (O_656,N_4710,N_4454);
nand UO_657 (O_657,N_4510,N_4028);
or UO_658 (O_658,N_4876,N_4575);
nand UO_659 (O_659,N_4542,N_4101);
nor UO_660 (O_660,N_4594,N_4731);
or UO_661 (O_661,N_4119,N_4016);
nor UO_662 (O_662,N_4662,N_4407);
or UO_663 (O_663,N_4744,N_4156);
nand UO_664 (O_664,N_4295,N_4622);
nand UO_665 (O_665,N_4014,N_4099);
or UO_666 (O_666,N_4382,N_4043);
and UO_667 (O_667,N_4666,N_4753);
or UO_668 (O_668,N_4732,N_4852);
and UO_669 (O_669,N_4690,N_4775);
and UO_670 (O_670,N_4560,N_4466);
or UO_671 (O_671,N_4488,N_4302);
and UO_672 (O_672,N_4974,N_4673);
and UO_673 (O_673,N_4296,N_4088);
nor UO_674 (O_674,N_4024,N_4180);
or UO_675 (O_675,N_4832,N_4672);
nor UO_676 (O_676,N_4709,N_4232);
nand UO_677 (O_677,N_4031,N_4860);
and UO_678 (O_678,N_4744,N_4777);
xnor UO_679 (O_679,N_4516,N_4043);
nand UO_680 (O_680,N_4714,N_4367);
and UO_681 (O_681,N_4920,N_4292);
or UO_682 (O_682,N_4536,N_4740);
nand UO_683 (O_683,N_4216,N_4005);
and UO_684 (O_684,N_4339,N_4868);
nor UO_685 (O_685,N_4087,N_4154);
or UO_686 (O_686,N_4623,N_4361);
nor UO_687 (O_687,N_4325,N_4650);
and UO_688 (O_688,N_4995,N_4776);
nand UO_689 (O_689,N_4844,N_4504);
xnor UO_690 (O_690,N_4783,N_4064);
or UO_691 (O_691,N_4780,N_4119);
and UO_692 (O_692,N_4400,N_4175);
nand UO_693 (O_693,N_4723,N_4681);
nand UO_694 (O_694,N_4644,N_4495);
or UO_695 (O_695,N_4116,N_4951);
and UO_696 (O_696,N_4991,N_4144);
nand UO_697 (O_697,N_4566,N_4844);
xnor UO_698 (O_698,N_4382,N_4348);
or UO_699 (O_699,N_4848,N_4320);
or UO_700 (O_700,N_4611,N_4062);
and UO_701 (O_701,N_4996,N_4281);
and UO_702 (O_702,N_4084,N_4917);
nor UO_703 (O_703,N_4581,N_4690);
nand UO_704 (O_704,N_4049,N_4708);
or UO_705 (O_705,N_4370,N_4701);
nand UO_706 (O_706,N_4144,N_4040);
and UO_707 (O_707,N_4162,N_4871);
or UO_708 (O_708,N_4763,N_4382);
and UO_709 (O_709,N_4164,N_4940);
and UO_710 (O_710,N_4375,N_4907);
and UO_711 (O_711,N_4035,N_4567);
nor UO_712 (O_712,N_4350,N_4725);
nand UO_713 (O_713,N_4599,N_4276);
or UO_714 (O_714,N_4773,N_4032);
or UO_715 (O_715,N_4721,N_4667);
nor UO_716 (O_716,N_4050,N_4204);
nor UO_717 (O_717,N_4019,N_4789);
xnor UO_718 (O_718,N_4883,N_4073);
nor UO_719 (O_719,N_4765,N_4502);
xnor UO_720 (O_720,N_4904,N_4215);
xor UO_721 (O_721,N_4378,N_4684);
nand UO_722 (O_722,N_4434,N_4601);
or UO_723 (O_723,N_4677,N_4044);
nor UO_724 (O_724,N_4719,N_4241);
or UO_725 (O_725,N_4070,N_4574);
or UO_726 (O_726,N_4495,N_4604);
nand UO_727 (O_727,N_4096,N_4075);
nor UO_728 (O_728,N_4866,N_4585);
and UO_729 (O_729,N_4810,N_4197);
nor UO_730 (O_730,N_4815,N_4035);
or UO_731 (O_731,N_4510,N_4301);
and UO_732 (O_732,N_4316,N_4005);
nand UO_733 (O_733,N_4823,N_4262);
nor UO_734 (O_734,N_4009,N_4200);
nand UO_735 (O_735,N_4537,N_4926);
nor UO_736 (O_736,N_4867,N_4355);
or UO_737 (O_737,N_4819,N_4813);
nand UO_738 (O_738,N_4905,N_4716);
or UO_739 (O_739,N_4932,N_4271);
nand UO_740 (O_740,N_4074,N_4494);
and UO_741 (O_741,N_4125,N_4906);
or UO_742 (O_742,N_4191,N_4616);
nand UO_743 (O_743,N_4040,N_4501);
nor UO_744 (O_744,N_4044,N_4362);
or UO_745 (O_745,N_4080,N_4138);
or UO_746 (O_746,N_4188,N_4782);
nor UO_747 (O_747,N_4624,N_4588);
nor UO_748 (O_748,N_4359,N_4839);
nand UO_749 (O_749,N_4233,N_4116);
or UO_750 (O_750,N_4183,N_4612);
or UO_751 (O_751,N_4886,N_4080);
nor UO_752 (O_752,N_4811,N_4003);
nand UO_753 (O_753,N_4157,N_4417);
or UO_754 (O_754,N_4147,N_4662);
nor UO_755 (O_755,N_4015,N_4423);
or UO_756 (O_756,N_4206,N_4903);
nand UO_757 (O_757,N_4793,N_4301);
and UO_758 (O_758,N_4750,N_4866);
nor UO_759 (O_759,N_4419,N_4219);
or UO_760 (O_760,N_4637,N_4489);
or UO_761 (O_761,N_4158,N_4608);
nand UO_762 (O_762,N_4059,N_4996);
nor UO_763 (O_763,N_4958,N_4882);
xor UO_764 (O_764,N_4437,N_4233);
nand UO_765 (O_765,N_4449,N_4820);
nand UO_766 (O_766,N_4175,N_4351);
or UO_767 (O_767,N_4396,N_4378);
nor UO_768 (O_768,N_4209,N_4040);
xnor UO_769 (O_769,N_4460,N_4884);
or UO_770 (O_770,N_4833,N_4041);
nor UO_771 (O_771,N_4331,N_4720);
and UO_772 (O_772,N_4190,N_4992);
nor UO_773 (O_773,N_4669,N_4686);
and UO_774 (O_774,N_4281,N_4783);
or UO_775 (O_775,N_4485,N_4376);
nor UO_776 (O_776,N_4788,N_4749);
and UO_777 (O_777,N_4351,N_4496);
nand UO_778 (O_778,N_4269,N_4928);
nor UO_779 (O_779,N_4072,N_4713);
and UO_780 (O_780,N_4568,N_4605);
nand UO_781 (O_781,N_4445,N_4412);
and UO_782 (O_782,N_4742,N_4772);
nand UO_783 (O_783,N_4112,N_4727);
nand UO_784 (O_784,N_4986,N_4210);
or UO_785 (O_785,N_4565,N_4036);
or UO_786 (O_786,N_4418,N_4777);
nor UO_787 (O_787,N_4122,N_4698);
nor UO_788 (O_788,N_4705,N_4500);
and UO_789 (O_789,N_4798,N_4441);
and UO_790 (O_790,N_4693,N_4819);
nand UO_791 (O_791,N_4432,N_4297);
nand UO_792 (O_792,N_4309,N_4958);
or UO_793 (O_793,N_4990,N_4288);
and UO_794 (O_794,N_4298,N_4476);
nand UO_795 (O_795,N_4934,N_4604);
nor UO_796 (O_796,N_4433,N_4339);
nor UO_797 (O_797,N_4285,N_4227);
nand UO_798 (O_798,N_4076,N_4896);
nand UO_799 (O_799,N_4997,N_4143);
and UO_800 (O_800,N_4097,N_4431);
nor UO_801 (O_801,N_4834,N_4547);
nor UO_802 (O_802,N_4545,N_4595);
and UO_803 (O_803,N_4119,N_4171);
or UO_804 (O_804,N_4137,N_4086);
or UO_805 (O_805,N_4304,N_4267);
or UO_806 (O_806,N_4174,N_4265);
nor UO_807 (O_807,N_4506,N_4584);
nor UO_808 (O_808,N_4783,N_4777);
xnor UO_809 (O_809,N_4352,N_4416);
nor UO_810 (O_810,N_4787,N_4169);
or UO_811 (O_811,N_4739,N_4545);
and UO_812 (O_812,N_4922,N_4011);
nor UO_813 (O_813,N_4194,N_4219);
and UO_814 (O_814,N_4965,N_4439);
nand UO_815 (O_815,N_4078,N_4458);
or UO_816 (O_816,N_4972,N_4441);
nor UO_817 (O_817,N_4377,N_4983);
nand UO_818 (O_818,N_4714,N_4447);
nand UO_819 (O_819,N_4183,N_4105);
or UO_820 (O_820,N_4730,N_4402);
and UO_821 (O_821,N_4666,N_4572);
nand UO_822 (O_822,N_4459,N_4466);
or UO_823 (O_823,N_4796,N_4338);
or UO_824 (O_824,N_4727,N_4883);
or UO_825 (O_825,N_4287,N_4358);
nor UO_826 (O_826,N_4391,N_4064);
and UO_827 (O_827,N_4488,N_4872);
nor UO_828 (O_828,N_4723,N_4441);
nor UO_829 (O_829,N_4293,N_4802);
and UO_830 (O_830,N_4823,N_4508);
xor UO_831 (O_831,N_4977,N_4394);
nor UO_832 (O_832,N_4563,N_4433);
nor UO_833 (O_833,N_4677,N_4878);
and UO_834 (O_834,N_4475,N_4140);
or UO_835 (O_835,N_4835,N_4723);
or UO_836 (O_836,N_4677,N_4987);
xnor UO_837 (O_837,N_4587,N_4551);
or UO_838 (O_838,N_4756,N_4154);
nor UO_839 (O_839,N_4330,N_4345);
and UO_840 (O_840,N_4780,N_4534);
nand UO_841 (O_841,N_4749,N_4985);
nand UO_842 (O_842,N_4227,N_4920);
and UO_843 (O_843,N_4625,N_4464);
nand UO_844 (O_844,N_4590,N_4731);
nand UO_845 (O_845,N_4533,N_4449);
or UO_846 (O_846,N_4924,N_4914);
and UO_847 (O_847,N_4452,N_4496);
nor UO_848 (O_848,N_4380,N_4900);
nor UO_849 (O_849,N_4883,N_4867);
nand UO_850 (O_850,N_4852,N_4987);
or UO_851 (O_851,N_4349,N_4498);
and UO_852 (O_852,N_4618,N_4078);
nor UO_853 (O_853,N_4198,N_4358);
nand UO_854 (O_854,N_4238,N_4599);
or UO_855 (O_855,N_4130,N_4181);
nand UO_856 (O_856,N_4512,N_4676);
nand UO_857 (O_857,N_4603,N_4419);
or UO_858 (O_858,N_4088,N_4219);
nand UO_859 (O_859,N_4505,N_4663);
and UO_860 (O_860,N_4946,N_4798);
nand UO_861 (O_861,N_4470,N_4317);
or UO_862 (O_862,N_4125,N_4039);
and UO_863 (O_863,N_4287,N_4567);
nor UO_864 (O_864,N_4395,N_4386);
nor UO_865 (O_865,N_4843,N_4168);
xor UO_866 (O_866,N_4002,N_4215);
xor UO_867 (O_867,N_4932,N_4059);
nand UO_868 (O_868,N_4376,N_4923);
or UO_869 (O_869,N_4231,N_4391);
or UO_870 (O_870,N_4355,N_4841);
nand UO_871 (O_871,N_4617,N_4067);
nor UO_872 (O_872,N_4274,N_4221);
or UO_873 (O_873,N_4223,N_4958);
and UO_874 (O_874,N_4681,N_4301);
or UO_875 (O_875,N_4753,N_4902);
nand UO_876 (O_876,N_4895,N_4210);
nand UO_877 (O_877,N_4767,N_4424);
or UO_878 (O_878,N_4874,N_4036);
or UO_879 (O_879,N_4781,N_4447);
or UO_880 (O_880,N_4695,N_4587);
or UO_881 (O_881,N_4040,N_4070);
nand UO_882 (O_882,N_4464,N_4242);
nand UO_883 (O_883,N_4117,N_4288);
or UO_884 (O_884,N_4507,N_4437);
nand UO_885 (O_885,N_4996,N_4745);
nor UO_886 (O_886,N_4182,N_4539);
nor UO_887 (O_887,N_4780,N_4174);
or UO_888 (O_888,N_4612,N_4391);
and UO_889 (O_889,N_4247,N_4016);
nand UO_890 (O_890,N_4946,N_4011);
nand UO_891 (O_891,N_4504,N_4590);
nor UO_892 (O_892,N_4082,N_4447);
and UO_893 (O_893,N_4855,N_4708);
xor UO_894 (O_894,N_4593,N_4971);
and UO_895 (O_895,N_4695,N_4923);
and UO_896 (O_896,N_4298,N_4083);
and UO_897 (O_897,N_4212,N_4599);
or UO_898 (O_898,N_4944,N_4348);
and UO_899 (O_899,N_4479,N_4405);
or UO_900 (O_900,N_4834,N_4223);
nand UO_901 (O_901,N_4477,N_4858);
and UO_902 (O_902,N_4648,N_4511);
nor UO_903 (O_903,N_4347,N_4968);
or UO_904 (O_904,N_4150,N_4091);
and UO_905 (O_905,N_4283,N_4744);
nand UO_906 (O_906,N_4190,N_4947);
nand UO_907 (O_907,N_4961,N_4255);
nand UO_908 (O_908,N_4283,N_4697);
and UO_909 (O_909,N_4410,N_4844);
xnor UO_910 (O_910,N_4217,N_4418);
nand UO_911 (O_911,N_4728,N_4319);
xor UO_912 (O_912,N_4771,N_4554);
nor UO_913 (O_913,N_4515,N_4431);
nand UO_914 (O_914,N_4328,N_4568);
or UO_915 (O_915,N_4370,N_4338);
or UO_916 (O_916,N_4798,N_4401);
nor UO_917 (O_917,N_4273,N_4331);
or UO_918 (O_918,N_4825,N_4984);
xnor UO_919 (O_919,N_4430,N_4252);
nand UO_920 (O_920,N_4310,N_4804);
xor UO_921 (O_921,N_4125,N_4989);
nor UO_922 (O_922,N_4059,N_4764);
or UO_923 (O_923,N_4891,N_4572);
nor UO_924 (O_924,N_4105,N_4948);
and UO_925 (O_925,N_4909,N_4915);
nor UO_926 (O_926,N_4145,N_4507);
and UO_927 (O_927,N_4558,N_4187);
and UO_928 (O_928,N_4867,N_4793);
nor UO_929 (O_929,N_4260,N_4758);
and UO_930 (O_930,N_4127,N_4843);
nor UO_931 (O_931,N_4405,N_4603);
or UO_932 (O_932,N_4503,N_4695);
or UO_933 (O_933,N_4323,N_4404);
or UO_934 (O_934,N_4577,N_4877);
nor UO_935 (O_935,N_4232,N_4866);
nor UO_936 (O_936,N_4298,N_4012);
nand UO_937 (O_937,N_4635,N_4105);
nand UO_938 (O_938,N_4662,N_4840);
xor UO_939 (O_939,N_4833,N_4196);
nand UO_940 (O_940,N_4869,N_4831);
nand UO_941 (O_941,N_4919,N_4928);
or UO_942 (O_942,N_4439,N_4618);
and UO_943 (O_943,N_4509,N_4333);
xor UO_944 (O_944,N_4755,N_4300);
and UO_945 (O_945,N_4011,N_4311);
or UO_946 (O_946,N_4024,N_4930);
and UO_947 (O_947,N_4998,N_4146);
or UO_948 (O_948,N_4411,N_4890);
and UO_949 (O_949,N_4635,N_4672);
nand UO_950 (O_950,N_4351,N_4229);
and UO_951 (O_951,N_4379,N_4033);
nor UO_952 (O_952,N_4833,N_4776);
or UO_953 (O_953,N_4931,N_4595);
nand UO_954 (O_954,N_4643,N_4530);
nand UO_955 (O_955,N_4946,N_4326);
nand UO_956 (O_956,N_4201,N_4842);
and UO_957 (O_957,N_4038,N_4405);
nor UO_958 (O_958,N_4642,N_4040);
nor UO_959 (O_959,N_4768,N_4719);
or UO_960 (O_960,N_4857,N_4080);
nor UO_961 (O_961,N_4940,N_4194);
nand UO_962 (O_962,N_4757,N_4752);
nand UO_963 (O_963,N_4207,N_4748);
and UO_964 (O_964,N_4026,N_4612);
nor UO_965 (O_965,N_4995,N_4859);
or UO_966 (O_966,N_4051,N_4188);
nand UO_967 (O_967,N_4112,N_4813);
or UO_968 (O_968,N_4929,N_4157);
and UO_969 (O_969,N_4038,N_4882);
and UO_970 (O_970,N_4028,N_4875);
nand UO_971 (O_971,N_4005,N_4171);
and UO_972 (O_972,N_4202,N_4649);
nor UO_973 (O_973,N_4438,N_4920);
nor UO_974 (O_974,N_4622,N_4778);
nand UO_975 (O_975,N_4164,N_4346);
nand UO_976 (O_976,N_4415,N_4338);
nor UO_977 (O_977,N_4359,N_4220);
and UO_978 (O_978,N_4160,N_4484);
nand UO_979 (O_979,N_4143,N_4425);
or UO_980 (O_980,N_4104,N_4627);
and UO_981 (O_981,N_4829,N_4146);
or UO_982 (O_982,N_4348,N_4923);
or UO_983 (O_983,N_4326,N_4647);
nor UO_984 (O_984,N_4092,N_4153);
and UO_985 (O_985,N_4286,N_4145);
nor UO_986 (O_986,N_4090,N_4741);
and UO_987 (O_987,N_4756,N_4832);
nand UO_988 (O_988,N_4417,N_4822);
or UO_989 (O_989,N_4895,N_4689);
or UO_990 (O_990,N_4861,N_4061);
or UO_991 (O_991,N_4807,N_4638);
and UO_992 (O_992,N_4745,N_4272);
and UO_993 (O_993,N_4696,N_4155);
or UO_994 (O_994,N_4073,N_4082);
nor UO_995 (O_995,N_4571,N_4493);
nor UO_996 (O_996,N_4628,N_4890);
nand UO_997 (O_997,N_4045,N_4589);
and UO_998 (O_998,N_4503,N_4368);
and UO_999 (O_999,N_4136,N_4713);
endmodule