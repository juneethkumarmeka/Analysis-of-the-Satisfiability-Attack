module basic_1500_15000_2000_20_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_373,In_781);
xor U1 (N_1,In_148,In_725);
and U2 (N_2,In_1017,In_677);
nor U3 (N_3,In_979,In_60);
xnor U4 (N_4,In_467,In_1199);
nor U5 (N_5,In_594,In_1088);
xnor U6 (N_6,In_574,In_952);
nor U7 (N_7,In_1124,In_716);
and U8 (N_8,In_1268,In_1257);
or U9 (N_9,In_771,In_1173);
nor U10 (N_10,In_109,In_668);
nor U11 (N_11,In_403,In_863);
nor U12 (N_12,In_122,In_1442);
nor U13 (N_13,In_453,In_253);
nor U14 (N_14,In_150,In_675);
xnor U15 (N_15,In_490,In_1115);
nor U16 (N_16,In_515,In_213);
and U17 (N_17,In_182,In_1427);
nand U18 (N_18,In_839,In_123);
nor U19 (N_19,In_57,In_73);
or U20 (N_20,In_942,In_46);
nor U21 (N_21,In_1476,In_522);
xnor U22 (N_22,In_1155,In_422);
nand U23 (N_23,In_1160,In_1215);
and U24 (N_24,In_1242,In_1392);
and U25 (N_25,In_462,In_731);
or U26 (N_26,In_56,In_1052);
xor U27 (N_27,In_1179,In_265);
xnor U28 (N_28,In_1484,In_706);
and U29 (N_29,In_286,In_282);
or U30 (N_30,In_1200,In_164);
or U31 (N_31,In_118,In_1041);
and U32 (N_32,In_824,In_1329);
or U33 (N_33,In_728,In_153);
nand U34 (N_34,In_11,In_380);
and U35 (N_35,In_1248,In_767);
nand U36 (N_36,In_1485,In_1491);
or U37 (N_37,In_24,In_1250);
nor U38 (N_38,In_1411,In_477);
nand U39 (N_39,In_1,In_978);
nor U40 (N_40,In_1496,In_217);
or U41 (N_41,In_919,In_599);
nand U42 (N_42,In_401,In_473);
nand U43 (N_43,In_708,In_1346);
nand U44 (N_44,In_1143,In_267);
xnor U45 (N_45,In_1420,In_87);
xor U46 (N_46,In_1236,In_793);
xor U47 (N_47,In_1459,In_1235);
nand U48 (N_48,In_171,In_529);
nand U49 (N_49,In_353,In_714);
or U50 (N_50,In_397,In_1376);
or U51 (N_51,In_51,In_970);
nor U52 (N_52,In_378,In_816);
nand U53 (N_53,In_748,In_1367);
nor U54 (N_54,In_975,In_658);
nand U55 (N_55,In_62,In_184);
or U56 (N_56,In_654,In_39);
xnor U57 (N_57,In_1312,In_533);
or U58 (N_58,In_1223,In_717);
or U59 (N_59,In_1359,In_877);
and U60 (N_60,In_961,In_275);
and U61 (N_61,In_96,In_832);
xnor U62 (N_62,In_1460,In_660);
xor U63 (N_63,In_279,In_1466);
nand U64 (N_64,In_916,In_216);
nor U65 (N_65,In_928,In_540);
nor U66 (N_66,In_1415,In_923);
nand U67 (N_67,In_91,In_235);
xor U68 (N_68,In_299,In_797);
xor U69 (N_69,In_1071,In_1452);
or U70 (N_70,In_488,In_45);
and U71 (N_71,In_1214,In_944);
xor U72 (N_72,In_493,In_898);
nand U73 (N_73,In_210,In_1313);
or U74 (N_74,In_1123,In_133);
xor U75 (N_75,In_1053,In_517);
nand U76 (N_76,In_1418,In_193);
or U77 (N_77,In_9,In_922);
and U78 (N_78,In_311,In_638);
and U79 (N_79,In_645,In_34);
nor U80 (N_80,In_609,In_390);
nand U81 (N_81,In_111,In_769);
nand U82 (N_82,In_146,In_1049);
and U83 (N_83,In_1399,In_450);
nand U84 (N_84,In_1158,In_1443);
and U85 (N_85,In_419,In_26);
or U86 (N_86,In_284,In_170);
and U87 (N_87,In_243,In_179);
and U88 (N_88,In_445,In_1067);
or U89 (N_89,In_836,In_1401);
xnor U90 (N_90,In_156,In_256);
nand U91 (N_91,In_71,In_200);
and U92 (N_92,In_705,In_1362);
nor U93 (N_93,In_225,In_1328);
and U94 (N_94,In_1077,In_1239);
xor U95 (N_95,In_16,In_242);
and U96 (N_96,In_766,In_692);
and U97 (N_97,In_630,In_1455);
xnor U98 (N_98,In_802,In_701);
nand U99 (N_99,In_1075,In_1438);
or U100 (N_100,In_583,In_365);
xor U101 (N_101,In_943,In_68);
or U102 (N_102,In_1119,In_1243);
xnor U103 (N_103,In_357,In_306);
nand U104 (N_104,In_425,In_976);
nor U105 (N_105,In_1456,In_1152);
and U106 (N_106,In_1187,In_1280);
nor U107 (N_107,In_21,In_196);
or U108 (N_108,In_546,In_508);
xnor U109 (N_109,In_1462,In_573);
nand U110 (N_110,In_869,In_1330);
and U111 (N_111,In_406,In_953);
or U112 (N_112,In_1360,In_1063);
or U113 (N_113,In_211,In_1426);
nor U114 (N_114,In_479,In_212);
xnor U115 (N_115,In_917,In_7);
nor U116 (N_116,In_966,In_288);
nand U117 (N_117,In_1159,In_69);
or U118 (N_118,In_1416,In_1206);
xor U119 (N_119,In_1389,In_1398);
xor U120 (N_120,In_537,In_910);
nand U121 (N_121,In_588,In_786);
or U122 (N_122,In_159,In_1269);
or U123 (N_123,In_399,In_590);
or U124 (N_124,In_1116,In_1073);
or U125 (N_125,In_1373,In_1209);
or U126 (N_126,In_1380,In_1148);
xnor U127 (N_127,In_469,In_729);
nor U128 (N_128,In_1439,In_871);
nor U129 (N_129,In_794,In_1185);
nand U130 (N_130,In_1461,In_998);
nor U131 (N_131,In_834,In_1271);
nand U132 (N_132,In_1180,In_643);
xor U133 (N_133,In_912,In_591);
nor U134 (N_134,In_138,In_957);
nand U135 (N_135,In_228,In_1107);
xnor U136 (N_136,In_787,In_1054);
nand U137 (N_137,In_709,In_199);
nor U138 (N_138,In_1080,In_608);
nand U139 (N_139,In_438,In_1387);
nand U140 (N_140,In_470,In_1393);
and U141 (N_141,In_757,In_1140);
nand U142 (N_142,In_855,In_1388);
nor U143 (N_143,In_1302,In_1232);
xnor U144 (N_144,In_926,In_1228);
nor U145 (N_145,In_1068,In_1081);
or U146 (N_146,In_801,In_856);
nor U147 (N_147,In_1381,In_831);
or U148 (N_148,In_1403,In_1009);
or U149 (N_149,In_1146,In_551);
or U150 (N_150,In_144,In_1246);
xnor U151 (N_151,In_407,In_1386);
xnor U152 (N_152,In_1106,In_328);
or U153 (N_153,In_486,In_1382);
and U154 (N_154,In_894,In_847);
xnor U155 (N_155,In_1413,In_330);
or U156 (N_156,In_1121,In_338);
nor U157 (N_157,In_75,In_690);
or U158 (N_158,In_1221,In_585);
xnor U159 (N_159,In_1400,In_349);
nor U160 (N_160,In_446,In_531);
nor U161 (N_161,In_959,In_99);
xnor U162 (N_162,In_1127,In_804);
xor U163 (N_163,In_968,In_1164);
nor U164 (N_164,In_94,In_730);
and U165 (N_165,In_49,In_119);
or U166 (N_166,In_218,In_644);
nand U167 (N_167,In_1365,In_1434);
xnor U168 (N_168,In_361,In_1024);
nand U169 (N_169,In_1066,In_678);
nor U170 (N_170,In_1495,In_1047);
xnor U171 (N_171,In_575,In_53);
nor U172 (N_172,In_1207,In_335);
xor U173 (N_173,In_185,In_1153);
nor U174 (N_174,In_84,In_232);
or U175 (N_175,In_1277,In_1102);
and U176 (N_176,In_167,In_1499);
nand U177 (N_177,In_688,In_1113);
and U178 (N_178,In_572,In_682);
nand U179 (N_179,In_61,In_1296);
xor U180 (N_180,In_635,In_521);
or U181 (N_181,In_155,In_1421);
nor U182 (N_182,In_798,In_1136);
and U183 (N_183,In_1132,In_261);
or U184 (N_184,In_79,In_319);
nor U185 (N_185,In_874,In_396);
xnor U186 (N_186,In_637,In_1110);
nor U187 (N_187,In_1454,In_954);
and U188 (N_188,In_958,In_647);
and U189 (N_189,In_411,In_1145);
and U190 (N_190,In_441,In_141);
or U191 (N_191,In_168,In_524);
and U192 (N_192,In_1061,In_893);
or U193 (N_193,In_270,In_1020);
and U194 (N_194,In_219,In_905);
xnor U195 (N_195,In_481,In_458);
nand U196 (N_196,In_656,In_784);
or U197 (N_197,In_271,In_761);
or U198 (N_198,In_819,In_121);
xnor U199 (N_199,In_773,In_1193);
and U200 (N_200,In_363,In_1056);
nor U201 (N_201,In_346,In_974);
nor U202 (N_202,In_972,In_13);
nor U203 (N_203,In_809,In_744);
and U204 (N_204,In_1375,In_1394);
or U205 (N_205,In_707,In_1408);
or U206 (N_206,In_240,In_1058);
xor U207 (N_207,In_77,In_358);
nor U208 (N_208,In_1483,In_665);
xor U209 (N_209,In_1135,In_776);
nand U210 (N_210,In_1410,In_828);
xor U211 (N_211,In_605,In_760);
xor U212 (N_212,In_126,In_613);
or U213 (N_213,In_747,In_614);
and U214 (N_214,In_1011,In_710);
nor U215 (N_215,In_864,In_902);
or U216 (N_216,In_1137,In_1266);
and U217 (N_217,In_444,In_694);
nor U218 (N_218,In_1383,In_745);
or U219 (N_219,In_393,In_440);
nor U220 (N_220,In_332,In_1151);
and U221 (N_221,In_431,In_372);
or U222 (N_222,In_553,In_1321);
nor U223 (N_223,In_1314,In_374);
nor U224 (N_224,In_1311,In_595);
nor U225 (N_225,In_806,In_160);
nand U226 (N_226,In_447,In_1497);
nor U227 (N_227,In_104,In_1281);
or U228 (N_228,In_1372,In_619);
nand U229 (N_229,In_1176,In_1170);
nand U230 (N_230,In_377,In_1197);
xnor U231 (N_231,In_296,In_686);
and U232 (N_232,In_618,In_715);
or U233 (N_233,In_738,In_1368);
nor U234 (N_234,In_110,In_339);
or U235 (N_235,In_724,In_1192);
and U236 (N_236,In_592,In_229);
and U237 (N_237,In_195,In_570);
and U238 (N_238,In_751,In_818);
and U239 (N_239,In_1174,In_949);
xnor U240 (N_240,In_937,In_903);
or U241 (N_241,In_835,In_541);
or U242 (N_242,In_1377,In_264);
or U243 (N_243,In_732,In_366);
and U244 (N_244,In_837,In_556);
nand U245 (N_245,In_1062,In_1256);
nand U246 (N_246,In_132,In_161);
xor U247 (N_247,In_1371,In_375);
or U248 (N_248,In_355,In_207);
and U249 (N_249,In_950,In_1051);
nor U250 (N_250,In_512,In_402);
nor U251 (N_251,In_280,In_1078);
nor U252 (N_252,In_495,In_586);
nor U253 (N_253,In_137,In_1251);
and U254 (N_254,In_866,In_1046);
xor U255 (N_255,In_226,In_134);
nand U256 (N_256,In_1288,In_139);
nand U257 (N_257,In_1396,In_1042);
and U258 (N_258,In_1264,In_1304);
xnor U259 (N_259,In_984,In_1308);
or U260 (N_260,In_1072,In_1293);
xor U261 (N_261,In_1402,In_941);
xor U262 (N_262,In_224,In_689);
or U263 (N_263,In_1134,In_1448);
nor U264 (N_264,In_203,In_868);
nand U265 (N_265,In_790,In_78);
and U266 (N_266,In_1275,In_879);
or U267 (N_267,In_1249,In_1282);
nand U268 (N_268,In_1339,In_414);
nand U269 (N_269,In_763,In_532);
or U270 (N_270,In_166,In_933);
and U271 (N_271,In_711,In_28);
and U272 (N_272,In_1366,In_1327);
nand U273 (N_273,In_130,In_97);
xor U274 (N_274,In_1220,In_89);
nor U275 (N_275,In_885,In_308);
nand U276 (N_276,In_530,In_1195);
or U277 (N_277,In_1423,In_1038);
nor U278 (N_278,In_43,In_1098);
nor U279 (N_279,In_965,In_1218);
or U280 (N_280,In_162,In_1338);
xor U281 (N_281,In_1358,In_1441);
nor U282 (N_282,In_260,In_102);
xnor U283 (N_283,In_115,In_254);
nor U284 (N_284,In_499,In_800);
xor U285 (N_285,In_999,In_1326);
and U286 (N_286,In_1165,In_191);
and U287 (N_287,In_258,In_1324);
and U288 (N_288,In_1120,In_1405);
or U289 (N_289,In_257,In_704);
nand U290 (N_290,In_876,In_15);
nor U291 (N_291,In_1322,In_222);
nor U292 (N_292,In_695,In_1087);
nor U293 (N_293,In_65,In_1292);
nand U294 (N_294,In_1108,In_921);
and U295 (N_295,In_1005,In_1231);
or U296 (N_296,In_1198,In_597);
nor U297 (N_297,In_721,In_865);
nor U298 (N_298,In_430,In_873);
nand U299 (N_299,In_4,In_50);
and U300 (N_300,In_221,In_1224);
nor U301 (N_301,In_733,In_1278);
or U302 (N_302,In_904,In_1297);
and U303 (N_303,In_789,In_336);
xor U304 (N_304,In_1070,In_175);
or U305 (N_305,In_813,In_858);
nor U306 (N_306,In_108,In_1361);
xnor U307 (N_307,In_140,In_227);
nor U308 (N_308,In_1008,In_823);
or U309 (N_309,In_606,In_487);
xor U310 (N_310,In_1479,In_973);
nor U311 (N_311,In_796,In_1352);
nor U312 (N_312,In_277,In_31);
and U313 (N_313,In_772,In_1216);
or U314 (N_314,In_343,In_1010);
nand U315 (N_315,In_245,In_989);
nand U316 (N_316,In_1099,In_1303);
nand U317 (N_317,In_1433,In_1182);
nand U318 (N_318,In_1014,In_1229);
xnor U319 (N_319,In_476,In_436);
and U320 (N_320,In_389,In_391);
nor U321 (N_321,In_1348,In_564);
or U322 (N_322,In_333,In_525);
or U323 (N_323,In_1130,In_812);
and U324 (N_324,In_454,In_1138);
nor U325 (N_325,In_421,In_1270);
xor U326 (N_326,In_1480,In_520);
or U327 (N_327,In_63,In_1184);
xor U328 (N_328,In_987,In_699);
and U329 (N_329,In_982,In_803);
or U330 (N_330,In_427,In_1055);
xor U331 (N_331,In_223,In_560);
nor U332 (N_332,In_1203,In_750);
nand U333 (N_333,In_1261,In_1279);
nand U334 (N_334,In_1202,In_603);
nor U335 (N_335,In_100,In_932);
nor U336 (N_336,In_32,In_1337);
nand U337 (N_337,In_755,In_833);
nand U338 (N_338,In_252,In_285);
nor U339 (N_339,In_951,In_309);
nor U340 (N_340,In_1457,In_1161);
or U341 (N_341,In_1186,In_734);
xnor U342 (N_342,In_1019,In_720);
nand U343 (N_343,In_547,In_627);
and U344 (N_344,In_88,In_713);
or U345 (N_345,In_1473,In_888);
nand U346 (N_346,In_151,In_0);
or U347 (N_347,In_693,In_1390);
xor U348 (N_348,In_1175,In_474);
xor U349 (N_349,In_337,In_895);
and U350 (N_350,In_535,In_384);
nand U351 (N_351,In_550,In_1139);
or U352 (N_352,In_817,In_1333);
nand U353 (N_353,In_501,In_661);
xor U354 (N_354,In_1344,In_1118);
and U355 (N_355,In_272,In_14);
xor U356 (N_356,In_281,In_687);
nand U357 (N_357,In_1370,In_983);
nor U358 (N_358,In_909,In_1350);
or U359 (N_359,In_1472,In_914);
nor U360 (N_360,In_20,In_1468);
nand U361 (N_361,In_1318,In_1447);
or U362 (N_362,In_1446,In_415);
nor U363 (N_363,In_852,In_37);
nor U364 (N_364,In_230,In_163);
nor U365 (N_365,In_95,In_1317);
or U366 (N_366,In_329,In_1492);
nor U367 (N_367,In_428,In_405);
xor U368 (N_368,In_341,In_154);
xor U369 (N_369,In_301,In_1050);
or U370 (N_370,In_849,In_187);
nand U371 (N_371,In_192,In_969);
nor U372 (N_372,In_1191,In_1286);
or U373 (N_373,In_369,In_3);
or U374 (N_374,In_679,In_719);
nor U375 (N_375,In_1210,In_418);
nand U376 (N_376,In_886,In_249);
and U377 (N_377,In_1002,In_566);
and U378 (N_378,In_1163,In_1498);
or U379 (N_379,In_1034,In_19);
nor U380 (N_380,In_316,In_360);
nor U381 (N_381,In_602,In_1004);
nor U382 (N_382,In_514,In_1385);
xnor U383 (N_383,In_274,In_194);
or U384 (N_384,In_752,In_680);
or U385 (N_385,In_534,In_1265);
or U386 (N_386,In_669,In_1273);
nand U387 (N_387,In_237,In_189);
and U388 (N_388,In_1252,In_569);
nor U389 (N_389,In_646,In_451);
nor U390 (N_390,In_1428,In_214);
xnor U391 (N_391,In_1272,In_1353);
or U392 (N_392,In_297,In_1222);
or U393 (N_393,In_502,In_649);
xor U394 (N_394,In_859,In_18);
or U395 (N_395,In_484,In_463);
xnor U396 (N_396,In_1431,In_1316);
and U397 (N_397,In_416,In_845);
xnor U398 (N_398,In_936,In_124);
and U399 (N_399,In_536,In_842);
xor U400 (N_400,In_1369,In_259);
nand U401 (N_401,In_511,In_367);
and U402 (N_402,In_593,In_173);
or U403 (N_403,In_209,In_1095);
nand U404 (N_404,In_1409,In_1213);
and U405 (N_405,In_1167,In_145);
nor U406 (N_406,In_1225,In_844);
or U407 (N_407,In_300,In_673);
xor U408 (N_408,In_413,In_549);
nor U409 (N_409,In_558,In_555);
nor U410 (N_410,In_452,In_33);
xnor U411 (N_411,In_636,In_664);
nor U412 (N_412,In_1237,In_1125);
nor U413 (N_413,In_101,In_1478);
nor U414 (N_414,In_578,In_653);
nand U415 (N_415,In_1449,In_1233);
or U416 (N_416,In_1494,In_820);
and U417 (N_417,In_147,In_404);
and U418 (N_418,In_875,In_35);
xor U419 (N_419,In_1306,In_468);
or U420 (N_420,In_351,In_657);
xor U421 (N_421,In_899,In_671);
or U422 (N_422,In_1026,In_727);
xnor U423 (N_423,In_1262,In_1000);
nor U424 (N_424,In_722,In_964);
or U425 (N_425,In_368,In_197);
or U426 (N_426,In_424,In_829);
and U427 (N_427,In_294,In_1065);
and U428 (N_428,In_685,In_456);
or U429 (N_429,In_5,In_726);
nand U430 (N_430,In_58,In_780);
and U431 (N_431,In_1267,In_273);
nor U432 (N_432,In_80,In_1445);
nand U433 (N_433,In_1453,In_552);
nand U434 (N_434,In_125,In_527);
nand U435 (N_435,In_234,In_1097);
and U436 (N_436,In_201,In_1432);
nand U437 (N_437,In_54,In_811);
nand U438 (N_438,In_674,In_1290);
nor U439 (N_439,In_741,In_239);
nand U440 (N_440,In_1319,In_149);
xnor U441 (N_441,In_236,In_52);
or U442 (N_442,In_394,In_12);
nand U443 (N_443,In_1032,In_872);
nor U444 (N_444,In_1301,In_900);
or U445 (N_445,In_483,In_538);
nor U446 (N_446,In_376,In_1196);
nor U447 (N_447,In_1253,In_1240);
and U448 (N_448,In_352,In_700);
nor U449 (N_449,In_610,In_74);
nand U450 (N_450,In_244,In_298);
nand U451 (N_451,In_92,In_1035);
or U452 (N_452,In_290,In_948);
nand U453 (N_453,In_429,In_276);
nor U454 (N_454,In_1458,In_408);
nand U455 (N_455,In_455,In_568);
or U456 (N_456,In_1487,In_1482);
or U457 (N_457,In_482,In_604);
xnor U458 (N_458,In_616,In_310);
xnor U459 (N_459,In_1040,In_417);
or U460 (N_460,In_1168,In_967);
nand U461 (N_461,In_523,In_190);
nand U462 (N_462,In_307,In_510);
or U463 (N_463,In_439,In_1341);
or U464 (N_464,In_882,In_291);
and U465 (N_465,In_157,In_652);
nand U466 (N_466,In_1397,In_626);
and U467 (N_467,In_90,In_841);
and U468 (N_468,In_437,In_1128);
and U469 (N_469,In_683,In_1245);
or U470 (N_470,In_1310,In_927);
nor U471 (N_471,In_1429,In_356);
nor U472 (N_472,In_1486,In_807);
xnor U473 (N_473,In_821,In_67);
xor U474 (N_474,In_1363,In_480);
xor U475 (N_475,In_105,In_906);
or U476 (N_476,In_896,In_205);
and U477 (N_477,In_736,In_840);
nor U478 (N_478,In_471,In_1238);
or U479 (N_479,In_810,In_30);
nand U480 (N_480,In_23,In_1320);
nor U481 (N_481,In_1336,In_387);
nand U482 (N_482,In_930,In_27);
or U483 (N_483,In_448,In_698);
nor U484 (N_484,In_526,In_1043);
xor U485 (N_485,In_1082,In_754);
or U486 (N_486,In_1469,In_774);
and U487 (N_487,In_600,In_131);
and U488 (N_488,In_303,In_116);
or U489 (N_489,In_1181,In_827);
and U490 (N_490,In_545,In_1379);
nor U491 (N_491,In_612,In_127);
nor U492 (N_492,In_881,In_518);
and U493 (N_493,In_1244,In_1156);
or U494 (N_494,In_347,In_313);
nand U495 (N_495,In_443,In_318);
nor U496 (N_496,In_791,In_1294);
xnor U497 (N_497,In_1178,In_601);
nor U498 (N_498,In_334,In_1059);
or U499 (N_499,In_248,In_1424);
or U500 (N_500,In_120,In_826);
or U501 (N_501,In_1157,In_1340);
or U502 (N_502,In_980,In_1255);
and U503 (N_503,In_1094,In_1299);
nand U504 (N_504,In_461,In_519);
xor U505 (N_505,In_98,In_1030);
or U506 (N_506,In_1103,In_615);
xor U507 (N_507,In_676,In_582);
xor U508 (N_508,In_442,In_631);
nor U509 (N_509,In_178,In_1343);
or U510 (N_510,In_231,In_577);
and U511 (N_511,In_862,In_1493);
and U512 (N_512,In_48,In_1006);
and U513 (N_513,In_1114,In_667);
and U514 (N_514,In_666,In_410);
nor U515 (N_515,In_620,In_1259);
nor U516 (N_516,In_740,In_8);
nand U517 (N_517,In_1028,In_1477);
or U518 (N_518,In_843,In_651);
and U519 (N_519,In_475,In_860);
and U520 (N_520,In_312,In_1463);
nand U521 (N_521,In_815,In_25);
and U522 (N_522,In_516,In_174);
nor U523 (N_523,In_1260,In_1033);
nor U524 (N_524,In_768,In_1171);
nor U525 (N_525,In_940,In_1354);
xnor U526 (N_526,In_1489,In_696);
or U527 (N_527,In_639,In_662);
xnor U528 (N_528,In_183,In_1364);
or U529 (N_529,In_304,In_889);
nor U530 (N_530,In_1144,In_1190);
nand U531 (N_531,In_1022,In_1488);
xor U532 (N_532,In_314,In_997);
nor U533 (N_533,In_584,In_543);
or U534 (N_534,In_625,In_246);
nand U535 (N_535,In_489,In_880);
xnor U536 (N_536,In_587,In_1141);
nand U537 (N_537,In_503,In_278);
nor U538 (N_538,In_388,In_792);
nor U539 (N_539,In_924,In_629);
and U540 (N_540,In_255,In_1470);
nand U541 (N_541,In_215,In_409);
or U542 (N_542,In_995,In_1241);
and U543 (N_543,In_1391,In_1332);
xnor U544 (N_544,In_1069,In_188);
nor U545 (N_545,In_1451,In_901);
xor U546 (N_546,In_753,In_322);
and U547 (N_547,In_1349,In_107);
nand U548 (N_548,In_457,In_1189);
and U549 (N_549,In_1287,In_1031);
nand U550 (N_550,In_1258,In_611);
and U551 (N_551,In_1212,In_742);
and U552 (N_552,In_465,In_931);
nor U553 (N_553,In_1417,In_1300);
nand U554 (N_554,In_496,In_775);
nor U555 (N_555,In_1091,In_106);
nand U556 (N_556,In_117,In_702);
and U557 (N_557,In_867,In_1142);
xnor U558 (N_558,In_412,In_1335);
and U559 (N_559,In_1384,In_756);
nor U560 (N_560,In_180,In_1464);
or U561 (N_561,In_2,In_1169);
and U562 (N_562,In_340,In_659);
xnor U563 (N_563,In_1101,In_136);
xnor U564 (N_564,In_655,In_41);
or U565 (N_565,In_321,In_492);
and U566 (N_566,In_6,In_262);
or U567 (N_567,In_345,In_498);
nor U568 (N_568,In_814,In_788);
nand U569 (N_569,In_42,In_268);
and U570 (N_570,In_617,In_44);
nand U571 (N_571,In_350,In_1425);
and U572 (N_572,In_1331,In_10);
nand U573 (N_573,In_1012,In_765);
nor U574 (N_574,In_1406,In_723);
and U575 (N_575,In_670,In_1284);
xor U576 (N_576,In_684,In_364);
or U577 (N_577,In_1436,In_295);
xnor U578 (N_578,In_762,In_233);
and U579 (N_579,In_1234,In_735);
or U580 (N_580,In_66,In_1465);
nor U581 (N_581,In_1204,In_325);
nor U582 (N_582,In_938,In_362);
nor U583 (N_583,In_712,In_81);
and U584 (N_584,In_1126,In_559);
and U585 (N_585,In_977,In_1217);
or U586 (N_586,In_317,In_663);
xnor U587 (N_587,In_947,In_563);
nand U588 (N_588,In_1183,In_971);
or U589 (N_589,In_1323,In_1263);
and U590 (N_590,In_1404,In_1039);
xor U591 (N_591,In_142,In_1219);
nor U592 (N_592,In_934,In_994);
or U593 (N_593,In_929,In_892);
and U594 (N_594,In_779,In_946);
nor U595 (N_595,In_509,In_1422);
nor U596 (N_596,In_420,In_320);
or U597 (N_597,In_491,In_1342);
nor U598 (N_598,In_59,In_581);
or U599 (N_599,In_40,In_1112);
and U600 (N_600,In_287,In_485);
or U601 (N_601,In_1021,In_238);
nor U602 (N_602,In_348,In_38);
or U603 (N_603,In_472,In_1407);
and U604 (N_604,In_825,In_1064);
nand U605 (N_605,In_263,In_1490);
or U606 (N_606,In_642,In_1430);
nand U607 (N_607,In_624,In_382);
nand U608 (N_608,In_623,In_939);
xor U609 (N_609,In_1208,In_996);
or U610 (N_610,In_854,In_460);
xor U611 (N_611,In_1147,In_143);
and U612 (N_612,In_1092,In_925);
xor U613 (N_613,In_1378,In_580);
nor U614 (N_614,In_758,In_991);
nand U615 (N_615,In_513,In_544);
and U616 (N_616,In_1254,In_1090);
xor U617 (N_617,In_778,In_47);
nor U618 (N_618,In_507,In_93);
nand U619 (N_619,In_1057,In_737);
xnor U620 (N_620,In_1188,In_181);
and U621 (N_621,In_1027,In_1395);
or U622 (N_622,In_1315,In_1334);
xnor U623 (N_623,In_114,In_1018);
xor U624 (N_624,In_433,In_423);
nand U625 (N_625,In_135,In_805);
and U626 (N_626,In_1467,In_1015);
nor U627 (N_627,In_1172,In_1309);
nor U628 (N_628,In_293,In_985);
and U629 (N_629,In_641,In_1194);
nor U630 (N_630,In_963,In_434);
nor U631 (N_631,In_177,In_1247);
nor U632 (N_632,In_746,In_1037);
nor U633 (N_633,In_466,In_956);
nand U634 (N_634,In_1111,In_1201);
nor U635 (N_635,In_992,In_1129);
or U636 (N_636,In_449,In_1086);
nor U637 (N_637,In_344,In_1166);
or U638 (N_638,In_165,In_283);
nand U639 (N_639,In_432,In_172);
xnor U640 (N_640,In_64,In_1048);
nor U641 (N_641,In_1440,In_565);
or U642 (N_642,In_799,In_1357);
xnor U643 (N_643,In_1412,In_158);
or U644 (N_644,In_1471,In_557);
and U645 (N_645,In_607,In_186);
or U646 (N_646,In_1083,In_1307);
nor U647 (N_647,In_589,In_920);
nor U648 (N_648,In_851,In_703);
or U649 (N_649,In_85,In_1295);
nand U650 (N_650,In_55,In_435);
nand U651 (N_651,In_506,In_1274);
and U652 (N_652,In_459,In_884);
xnor U653 (N_653,In_628,In_1205);
or U654 (N_654,In_381,In_206);
nand U655 (N_655,In_1230,In_1029);
nand U656 (N_656,In_247,In_935);
or U657 (N_657,In_571,In_241);
or U658 (N_658,In_1226,In_70);
nor U659 (N_659,In_539,In_386);
nand U660 (N_660,In_1084,In_315);
and U661 (N_661,In_198,In_129);
and U662 (N_662,In_22,In_1007);
and U663 (N_663,In_554,In_1177);
or U664 (N_664,In_945,In_331);
nand U665 (N_665,In_305,In_634);
nor U666 (N_666,In_1076,In_567);
or U667 (N_667,In_681,In_883);
nand U668 (N_668,In_718,In_870);
xor U669 (N_669,In_621,In_962);
nor U670 (N_670,In_528,In_1036);
or U671 (N_671,In_1351,In_152);
nand U672 (N_672,In_302,In_1276);
and U673 (N_673,In_579,In_907);
xor U674 (N_674,In_505,In_633);
or U675 (N_675,In_857,In_981);
or U676 (N_676,In_385,In_1045);
nand U677 (N_677,In_324,In_1474);
or U678 (N_678,In_1149,In_887);
or U679 (N_679,In_576,In_640);
and U680 (N_680,In_398,In_908);
nor U681 (N_681,In_76,In_1444);
nand U682 (N_682,In_266,In_1109);
and U683 (N_683,In_878,In_1085);
nor U684 (N_684,In_176,In_395);
xnor U685 (N_685,In_36,In_897);
nor U686 (N_686,In_208,In_1093);
xnor U687 (N_687,In_596,In_292);
nor U688 (N_688,In_1355,In_822);
xnor U689 (N_689,In_17,In_1345);
or U690 (N_690,In_359,In_128);
nor U691 (N_691,In_202,In_743);
and U692 (N_692,In_1414,In_383);
xor U693 (N_693,In_112,In_323);
nand U694 (N_694,In_86,In_1044);
nand U695 (N_695,In_251,In_250);
xnor U696 (N_696,In_478,In_562);
nand U697 (N_697,In_749,In_342);
xor U698 (N_698,In_1347,In_289);
xor U699 (N_699,In_269,In_850);
or U700 (N_700,In_1100,In_72);
nand U701 (N_701,In_622,In_672);
and U702 (N_702,In_785,In_1289);
or U703 (N_703,In_426,In_82);
and U704 (N_704,In_918,In_1154);
or U705 (N_705,In_955,In_777);
xnor U706 (N_706,In_1025,In_1023);
and U707 (N_707,In_392,In_795);
or U708 (N_708,In_29,In_1003);
xor U709 (N_709,In_848,In_915);
nor U710 (N_710,In_83,In_1013);
xnor U711 (N_711,In_759,In_103);
xnor U712 (N_712,In_1089,In_739);
and U713 (N_713,In_1325,In_1079);
and U714 (N_714,In_650,In_846);
nor U715 (N_715,In_354,In_1211);
xnor U716 (N_716,In_379,In_370);
nor U717 (N_717,In_494,In_1374);
xor U718 (N_718,In_1162,In_988);
nand U719 (N_719,In_169,In_1131);
and U720 (N_720,In_371,In_691);
and U721 (N_721,In_1001,In_1305);
and U722 (N_722,In_1096,In_913);
xor U723 (N_723,In_548,In_1150);
nand U724 (N_724,In_500,In_1285);
nor U725 (N_725,In_326,In_1291);
nand U726 (N_726,In_648,In_890);
and U727 (N_727,In_497,In_542);
nand U728 (N_728,In_1016,In_204);
and U729 (N_729,In_561,In_1283);
nor U730 (N_730,In_1074,In_770);
or U731 (N_731,In_1133,In_1356);
or U732 (N_732,In_1419,In_986);
xnor U733 (N_733,In_464,In_990);
or U734 (N_734,In_1105,In_1298);
and U735 (N_735,In_1437,In_891);
nor U736 (N_736,In_1227,In_911);
and U737 (N_737,In_783,In_838);
xor U738 (N_738,In_632,In_861);
and U739 (N_739,In_598,In_1435);
nand U740 (N_740,In_504,In_853);
nand U741 (N_741,In_1122,In_808);
and U742 (N_742,In_220,In_1117);
xor U743 (N_743,In_697,In_830);
xor U744 (N_744,In_400,In_1475);
and U745 (N_745,In_764,In_1104);
or U746 (N_746,In_960,In_327);
nand U747 (N_747,In_782,In_113);
nand U748 (N_748,In_993,In_1481);
or U749 (N_749,In_1450,In_1060);
xnor U750 (N_750,N_245,N_28);
or U751 (N_751,N_636,N_274);
nand U752 (N_752,N_405,N_477);
nand U753 (N_753,N_183,N_241);
nor U754 (N_754,N_239,N_533);
nand U755 (N_755,N_728,N_289);
and U756 (N_756,N_198,N_266);
or U757 (N_757,N_300,N_738);
xor U758 (N_758,N_562,N_427);
xor U759 (N_759,N_362,N_246);
nand U760 (N_760,N_708,N_354);
nor U761 (N_761,N_600,N_80);
and U762 (N_762,N_382,N_473);
nor U763 (N_763,N_70,N_438);
and U764 (N_764,N_171,N_748);
and U765 (N_765,N_309,N_744);
xor U766 (N_766,N_256,N_252);
nor U767 (N_767,N_125,N_459);
or U768 (N_768,N_116,N_574);
nor U769 (N_769,N_567,N_508);
nor U770 (N_770,N_168,N_392);
nor U771 (N_771,N_659,N_527);
xnor U772 (N_772,N_719,N_177);
xor U773 (N_773,N_400,N_419);
and U774 (N_774,N_449,N_740);
nand U775 (N_775,N_337,N_320);
nor U776 (N_776,N_646,N_620);
nand U777 (N_777,N_645,N_683);
nor U778 (N_778,N_155,N_154);
or U779 (N_779,N_501,N_511);
nand U780 (N_780,N_10,N_253);
xor U781 (N_781,N_234,N_514);
nand U782 (N_782,N_356,N_306);
or U783 (N_783,N_684,N_561);
and U784 (N_784,N_524,N_212);
xnor U785 (N_785,N_414,N_553);
or U786 (N_786,N_389,N_330);
and U787 (N_787,N_550,N_394);
and U788 (N_788,N_216,N_662);
xor U789 (N_789,N_675,N_705);
nand U790 (N_790,N_423,N_361);
or U791 (N_791,N_279,N_148);
nand U792 (N_792,N_98,N_209);
or U793 (N_793,N_175,N_404);
and U794 (N_794,N_580,N_677);
and U795 (N_795,N_189,N_29);
xnor U796 (N_796,N_30,N_136);
and U797 (N_797,N_421,N_525);
nor U798 (N_798,N_140,N_44);
xnor U799 (N_799,N_55,N_27);
and U800 (N_800,N_673,N_446);
nor U801 (N_801,N_113,N_416);
or U802 (N_802,N_66,N_386);
nor U803 (N_803,N_488,N_56);
and U804 (N_804,N_326,N_69);
xor U805 (N_805,N_255,N_224);
or U806 (N_806,N_720,N_443);
nor U807 (N_807,N_199,N_624);
nand U808 (N_808,N_313,N_424);
and U809 (N_809,N_547,N_712);
and U810 (N_810,N_471,N_267);
nor U811 (N_811,N_32,N_745);
or U812 (N_812,N_331,N_79);
or U813 (N_813,N_587,N_182);
nand U814 (N_814,N_22,N_538);
and U815 (N_815,N_544,N_340);
nor U816 (N_816,N_240,N_229);
and U817 (N_817,N_259,N_709);
nor U818 (N_818,N_89,N_322);
nor U819 (N_819,N_746,N_717);
nand U820 (N_820,N_11,N_180);
nor U821 (N_821,N_417,N_582);
or U822 (N_822,N_627,N_83);
nor U823 (N_823,N_144,N_702);
xor U824 (N_824,N_96,N_339);
nand U825 (N_825,N_741,N_689);
nor U826 (N_826,N_594,N_53);
or U827 (N_827,N_21,N_733);
and U828 (N_828,N_222,N_455);
xnor U829 (N_829,N_666,N_93);
or U830 (N_830,N_294,N_197);
nor U831 (N_831,N_608,N_505);
or U832 (N_832,N_138,N_433);
nor U833 (N_833,N_130,N_590);
nor U834 (N_834,N_429,N_36);
and U835 (N_835,N_307,N_617);
or U836 (N_836,N_24,N_325);
nand U837 (N_837,N_577,N_163);
xor U838 (N_838,N_679,N_243);
nor U839 (N_839,N_112,N_217);
or U840 (N_840,N_552,N_342);
xor U841 (N_841,N_203,N_515);
or U842 (N_842,N_440,N_6);
and U843 (N_843,N_598,N_468);
nor U844 (N_844,N_609,N_181);
or U845 (N_845,N_506,N_191);
nor U846 (N_846,N_616,N_166);
nand U847 (N_847,N_467,N_640);
or U848 (N_848,N_481,N_201);
nor U849 (N_849,N_535,N_126);
nand U850 (N_850,N_162,N_393);
and U851 (N_851,N_291,N_97);
nand U852 (N_852,N_391,N_678);
or U853 (N_853,N_132,N_491);
xor U854 (N_854,N_41,N_653);
nor U855 (N_855,N_457,N_575);
xor U856 (N_856,N_588,N_583);
xnor U857 (N_857,N_301,N_651);
nor U858 (N_858,N_61,N_244);
nor U859 (N_859,N_411,N_31);
nand U860 (N_860,N_293,N_165);
nor U861 (N_861,N_570,N_38);
and U862 (N_862,N_559,N_335);
nand U863 (N_863,N_176,N_124);
and U864 (N_864,N_435,N_341);
or U865 (N_865,N_42,N_447);
and U866 (N_866,N_304,N_110);
or U867 (N_867,N_334,N_4);
nor U868 (N_868,N_332,N_13);
xnor U869 (N_869,N_188,N_114);
nor U870 (N_870,N_448,N_739);
or U871 (N_871,N_57,N_642);
and U872 (N_872,N_551,N_19);
or U873 (N_873,N_284,N_220);
nand U874 (N_874,N_613,N_84);
or U875 (N_875,N_599,N_548);
xnor U876 (N_876,N_426,N_682);
nand U877 (N_877,N_532,N_311);
and U878 (N_878,N_249,N_466);
nor U879 (N_879,N_157,N_275);
nand U880 (N_880,N_365,N_46);
nor U881 (N_881,N_686,N_206);
and U882 (N_882,N_12,N_494);
nand U883 (N_883,N_196,N_529);
nand U884 (N_884,N_366,N_3);
nand U885 (N_885,N_370,N_167);
nand U886 (N_886,N_282,N_736);
and U887 (N_887,N_692,N_236);
nor U888 (N_888,N_101,N_352);
xor U889 (N_889,N_487,N_480);
nand U890 (N_890,N_102,N_159);
and U891 (N_891,N_727,N_106);
nand U892 (N_892,N_528,N_81);
nand U893 (N_893,N_86,N_169);
or U894 (N_894,N_91,N_564);
nand U895 (N_895,N_621,N_638);
or U896 (N_896,N_498,N_396);
nand U897 (N_897,N_497,N_513);
nor U898 (N_898,N_237,N_611);
nor U899 (N_899,N_399,N_472);
nand U900 (N_900,N_82,N_158);
nand U901 (N_901,N_543,N_78);
and U902 (N_902,N_635,N_699);
xnor U903 (N_903,N_314,N_17);
xnor U904 (N_904,N_1,N_463);
nand U905 (N_905,N_359,N_412);
nor U906 (N_906,N_72,N_633);
nand U907 (N_907,N_310,N_742);
nor U908 (N_908,N_413,N_479);
or U909 (N_909,N_593,N_456);
nor U910 (N_910,N_16,N_374);
and U911 (N_911,N_601,N_554);
nand U912 (N_912,N_418,N_40);
nand U913 (N_913,N_278,N_518);
and U914 (N_914,N_644,N_139);
nor U915 (N_915,N_451,N_401);
nand U916 (N_916,N_725,N_718);
nor U917 (N_917,N_129,N_735);
nand U918 (N_918,N_333,N_441);
xor U919 (N_919,N_663,N_670);
nor U920 (N_920,N_495,N_496);
or U921 (N_921,N_674,N_474);
xnor U922 (N_922,N_76,N_348);
and U923 (N_923,N_484,N_661);
and U924 (N_924,N_704,N_732);
nand U925 (N_925,N_607,N_280);
nand U926 (N_926,N_190,N_485);
nand U927 (N_927,N_214,N_147);
xor U928 (N_928,N_227,N_486);
nor U929 (N_929,N_254,N_460);
and U930 (N_930,N_127,N_195);
or U931 (N_931,N_437,N_25);
and U932 (N_932,N_265,N_161);
or U933 (N_933,N_377,N_226);
xor U934 (N_934,N_403,N_556);
nor U935 (N_935,N_290,N_656);
or U936 (N_936,N_444,N_297);
xnor U937 (N_937,N_749,N_131);
nand U938 (N_938,N_271,N_308);
and U939 (N_939,N_469,N_60);
xnor U940 (N_940,N_235,N_637);
nand U941 (N_941,N_576,N_632);
nor U942 (N_942,N_225,N_650);
or U943 (N_943,N_629,N_298);
xnor U944 (N_944,N_368,N_118);
nor U945 (N_945,N_694,N_184);
nor U946 (N_946,N_18,N_250);
xor U947 (N_947,N_630,N_523);
xor U948 (N_948,N_453,N_422);
and U949 (N_949,N_104,N_315);
xnor U950 (N_950,N_281,N_390);
nand U951 (N_951,N_302,N_39);
xor U952 (N_952,N_586,N_179);
or U953 (N_953,N_431,N_75);
xor U954 (N_954,N_264,N_94);
and U955 (N_955,N_737,N_230);
or U956 (N_956,N_517,N_296);
nand U957 (N_957,N_273,N_672);
xnor U958 (N_958,N_103,N_628);
nand U959 (N_959,N_660,N_489);
or U960 (N_960,N_285,N_350);
and U961 (N_961,N_522,N_261);
nand U962 (N_962,N_572,N_571);
nor U963 (N_963,N_406,N_379);
nand U964 (N_964,N_478,N_316);
nand U965 (N_965,N_597,N_269);
xnor U966 (N_966,N_664,N_251);
nor U967 (N_967,N_671,N_33);
nor U968 (N_968,N_85,N_436);
and U969 (N_969,N_724,N_619);
xor U970 (N_970,N_615,N_64);
xor U971 (N_971,N_693,N_614);
and U972 (N_972,N_648,N_283);
or U973 (N_973,N_384,N_512);
xnor U974 (N_974,N_74,N_430);
nor U975 (N_975,N_346,N_530);
or U976 (N_976,N_408,N_319);
or U977 (N_977,N_634,N_71);
nand U978 (N_978,N_109,N_713);
xnor U979 (N_979,N_50,N_303);
nor U980 (N_980,N_458,N_685);
nor U981 (N_981,N_120,N_160);
or U982 (N_982,N_90,N_626);
nor U983 (N_983,N_321,N_286);
or U984 (N_984,N_462,N_141);
or U985 (N_985,N_48,N_151);
xnor U986 (N_986,N_743,N_707);
or U987 (N_987,N_383,N_37);
nor U988 (N_988,N_351,N_150);
and U989 (N_989,N_465,N_592);
xnor U990 (N_990,N_111,N_218);
nand U991 (N_991,N_247,N_625);
nand U992 (N_992,N_299,N_715);
or U993 (N_993,N_657,N_123);
and U994 (N_994,N_100,N_665);
xnor U995 (N_995,N_730,N_710);
xor U996 (N_996,N_336,N_353);
and U997 (N_997,N_649,N_563);
xnor U998 (N_998,N_65,N_54);
nand U999 (N_999,N_149,N_714);
nor U1000 (N_1000,N_15,N_450);
nor U1001 (N_1001,N_503,N_584);
nand U1002 (N_1002,N_581,N_639);
nand U1003 (N_1003,N_328,N_329);
and U1004 (N_1004,N_541,N_402);
or U1005 (N_1005,N_287,N_606);
nand U1006 (N_1006,N_270,N_729);
nand U1007 (N_1007,N_483,N_122);
nor U1008 (N_1008,N_146,N_45);
and U1009 (N_1009,N_68,N_0);
or U1010 (N_1010,N_612,N_669);
nand U1011 (N_1011,N_119,N_407);
or U1012 (N_1012,N_49,N_680);
nand U1013 (N_1013,N_117,N_360);
nor U1014 (N_1014,N_170,N_697);
xnor U1015 (N_1015,N_691,N_681);
nand U1016 (N_1016,N_73,N_557);
xor U1017 (N_1017,N_312,N_260);
nand U1018 (N_1018,N_442,N_482);
xnor U1019 (N_1019,N_186,N_723);
xnor U1020 (N_1020,N_380,N_569);
xor U1021 (N_1021,N_409,N_654);
or U1022 (N_1022,N_200,N_452);
or U1023 (N_1023,N_263,N_432);
xnor U1024 (N_1024,N_610,N_213);
nor U1025 (N_1025,N_534,N_142);
and U1026 (N_1026,N_215,N_470);
nor U1027 (N_1027,N_231,N_23);
and U1028 (N_1028,N_349,N_115);
nand U1029 (N_1029,N_690,N_204);
nor U1030 (N_1030,N_134,N_500);
and U1031 (N_1031,N_622,N_133);
nor U1032 (N_1032,N_258,N_26);
nand U1033 (N_1033,N_276,N_502);
and U1034 (N_1034,N_652,N_591);
nand U1035 (N_1035,N_476,N_324);
xnor U1036 (N_1036,N_375,N_317);
or U1037 (N_1037,N_493,N_59);
or U1038 (N_1038,N_262,N_565);
nor U1039 (N_1039,N_268,N_135);
nand U1040 (N_1040,N_34,N_381);
or U1041 (N_1041,N_355,N_373);
nand U1042 (N_1042,N_578,N_376);
nor U1043 (N_1043,N_647,N_605);
and U1044 (N_1044,N_420,N_428);
nor U1045 (N_1045,N_153,N_734);
xnor U1046 (N_1046,N_549,N_210);
nand U1047 (N_1047,N_542,N_272);
nor U1048 (N_1048,N_504,N_358);
nor U1049 (N_1049,N_706,N_371);
or U1050 (N_1050,N_604,N_520);
and U1051 (N_1051,N_521,N_499);
nor U1052 (N_1052,N_388,N_105);
nor U1053 (N_1053,N_211,N_192);
nand U1054 (N_1054,N_526,N_14);
nand U1055 (N_1055,N_454,N_676);
nand U1056 (N_1056,N_461,N_248);
nor U1057 (N_1057,N_178,N_716);
and U1058 (N_1058,N_47,N_338);
or U1059 (N_1059,N_43,N_475);
nand U1060 (N_1060,N_579,N_173);
and U1061 (N_1061,N_363,N_128);
or U1062 (N_1062,N_589,N_623);
or U1063 (N_1063,N_367,N_152);
nor U1064 (N_1064,N_35,N_585);
nand U1065 (N_1065,N_107,N_193);
nand U1066 (N_1066,N_143,N_137);
xnor U1067 (N_1067,N_711,N_726);
nor U1068 (N_1068,N_208,N_318);
and U1069 (N_1069,N_108,N_536);
and U1070 (N_1070,N_67,N_667);
or U1071 (N_1071,N_164,N_9);
nor U1072 (N_1072,N_603,N_121);
xor U1073 (N_1073,N_695,N_602);
xor U1074 (N_1074,N_539,N_242);
or U1075 (N_1075,N_658,N_560);
and U1076 (N_1076,N_410,N_747);
xor U1077 (N_1077,N_92,N_385);
or U1078 (N_1078,N_531,N_207);
nor U1079 (N_1079,N_77,N_566);
nor U1080 (N_1080,N_345,N_722);
nor U1081 (N_1081,N_277,N_492);
nand U1082 (N_1082,N_323,N_369);
xor U1083 (N_1083,N_545,N_233);
or U1084 (N_1084,N_688,N_568);
xnor U1085 (N_1085,N_174,N_357);
nand U1086 (N_1086,N_238,N_464);
nand U1087 (N_1087,N_519,N_295);
nor U1088 (N_1088,N_509,N_573);
xor U1089 (N_1089,N_507,N_88);
nor U1090 (N_1090,N_221,N_537);
nand U1091 (N_1091,N_5,N_228);
nor U1092 (N_1092,N_643,N_698);
nor U1093 (N_1093,N_62,N_641);
xor U1094 (N_1094,N_63,N_696);
nor U1095 (N_1095,N_292,N_445);
and U1096 (N_1096,N_344,N_415);
xor U1097 (N_1097,N_701,N_395);
and U1098 (N_1098,N_595,N_700);
nand U1099 (N_1099,N_20,N_194);
nand U1100 (N_1100,N_490,N_434);
xor U1101 (N_1101,N_631,N_95);
nand U1102 (N_1102,N_51,N_618);
nor U1103 (N_1103,N_185,N_347);
nand U1104 (N_1104,N_397,N_439);
nor U1105 (N_1105,N_378,N_425);
nor U1106 (N_1106,N_655,N_668);
xnor U1107 (N_1107,N_219,N_205);
xnor U1108 (N_1108,N_257,N_372);
xnor U1109 (N_1109,N_596,N_223);
or U1110 (N_1110,N_305,N_232);
or U1111 (N_1111,N_387,N_187);
xor U1112 (N_1112,N_58,N_540);
nor U1113 (N_1113,N_172,N_87);
xnor U1114 (N_1114,N_731,N_99);
and U1115 (N_1115,N_703,N_145);
nand U1116 (N_1116,N_398,N_7);
nand U1117 (N_1117,N_510,N_343);
nor U1118 (N_1118,N_555,N_327);
xor U1119 (N_1119,N_516,N_202);
nor U1120 (N_1120,N_288,N_546);
xor U1121 (N_1121,N_2,N_558);
xnor U1122 (N_1122,N_721,N_687);
nor U1123 (N_1123,N_52,N_364);
xor U1124 (N_1124,N_8,N_156);
nand U1125 (N_1125,N_294,N_124);
and U1126 (N_1126,N_627,N_320);
nor U1127 (N_1127,N_306,N_611);
and U1128 (N_1128,N_438,N_680);
xor U1129 (N_1129,N_644,N_499);
or U1130 (N_1130,N_606,N_651);
and U1131 (N_1131,N_179,N_103);
and U1132 (N_1132,N_103,N_74);
nand U1133 (N_1133,N_670,N_487);
nor U1134 (N_1134,N_6,N_514);
nand U1135 (N_1135,N_542,N_4);
and U1136 (N_1136,N_410,N_81);
nor U1137 (N_1137,N_352,N_633);
and U1138 (N_1138,N_315,N_409);
and U1139 (N_1139,N_677,N_4);
nor U1140 (N_1140,N_528,N_648);
and U1141 (N_1141,N_658,N_370);
nand U1142 (N_1142,N_283,N_367);
nor U1143 (N_1143,N_493,N_707);
and U1144 (N_1144,N_419,N_285);
nand U1145 (N_1145,N_700,N_677);
and U1146 (N_1146,N_694,N_227);
and U1147 (N_1147,N_493,N_276);
and U1148 (N_1148,N_116,N_564);
and U1149 (N_1149,N_29,N_349);
and U1150 (N_1150,N_173,N_4);
xor U1151 (N_1151,N_635,N_332);
or U1152 (N_1152,N_451,N_246);
nor U1153 (N_1153,N_144,N_551);
xnor U1154 (N_1154,N_21,N_432);
nor U1155 (N_1155,N_211,N_89);
and U1156 (N_1156,N_532,N_70);
and U1157 (N_1157,N_540,N_92);
xor U1158 (N_1158,N_703,N_346);
and U1159 (N_1159,N_208,N_264);
nand U1160 (N_1160,N_597,N_644);
and U1161 (N_1161,N_332,N_595);
xnor U1162 (N_1162,N_462,N_348);
or U1163 (N_1163,N_399,N_467);
xnor U1164 (N_1164,N_589,N_14);
nand U1165 (N_1165,N_26,N_355);
and U1166 (N_1166,N_364,N_577);
nor U1167 (N_1167,N_462,N_160);
or U1168 (N_1168,N_29,N_680);
and U1169 (N_1169,N_479,N_381);
or U1170 (N_1170,N_375,N_681);
or U1171 (N_1171,N_690,N_47);
xnor U1172 (N_1172,N_227,N_675);
nor U1173 (N_1173,N_707,N_259);
or U1174 (N_1174,N_290,N_406);
or U1175 (N_1175,N_366,N_285);
nor U1176 (N_1176,N_606,N_597);
xnor U1177 (N_1177,N_480,N_153);
nand U1178 (N_1178,N_254,N_586);
nor U1179 (N_1179,N_401,N_188);
nand U1180 (N_1180,N_539,N_518);
nand U1181 (N_1181,N_528,N_222);
and U1182 (N_1182,N_16,N_286);
and U1183 (N_1183,N_458,N_210);
or U1184 (N_1184,N_118,N_502);
and U1185 (N_1185,N_251,N_17);
xor U1186 (N_1186,N_734,N_253);
nor U1187 (N_1187,N_634,N_225);
and U1188 (N_1188,N_5,N_645);
nor U1189 (N_1189,N_674,N_719);
or U1190 (N_1190,N_612,N_712);
or U1191 (N_1191,N_495,N_723);
xor U1192 (N_1192,N_156,N_543);
and U1193 (N_1193,N_700,N_275);
nor U1194 (N_1194,N_570,N_130);
xor U1195 (N_1195,N_446,N_98);
nor U1196 (N_1196,N_350,N_339);
nand U1197 (N_1197,N_488,N_148);
xnor U1198 (N_1198,N_145,N_332);
or U1199 (N_1199,N_680,N_408);
nor U1200 (N_1200,N_203,N_436);
xnor U1201 (N_1201,N_248,N_174);
xor U1202 (N_1202,N_523,N_556);
nand U1203 (N_1203,N_372,N_545);
or U1204 (N_1204,N_335,N_563);
xnor U1205 (N_1205,N_604,N_214);
or U1206 (N_1206,N_306,N_584);
or U1207 (N_1207,N_722,N_236);
or U1208 (N_1208,N_328,N_455);
nor U1209 (N_1209,N_464,N_444);
xor U1210 (N_1210,N_571,N_163);
or U1211 (N_1211,N_202,N_236);
and U1212 (N_1212,N_444,N_257);
xor U1213 (N_1213,N_81,N_1);
xnor U1214 (N_1214,N_369,N_483);
or U1215 (N_1215,N_592,N_400);
nor U1216 (N_1216,N_687,N_564);
or U1217 (N_1217,N_92,N_517);
xor U1218 (N_1218,N_383,N_741);
nand U1219 (N_1219,N_692,N_500);
nor U1220 (N_1220,N_166,N_623);
xnor U1221 (N_1221,N_463,N_416);
and U1222 (N_1222,N_547,N_747);
or U1223 (N_1223,N_376,N_354);
or U1224 (N_1224,N_733,N_5);
nor U1225 (N_1225,N_376,N_687);
nand U1226 (N_1226,N_700,N_734);
nor U1227 (N_1227,N_155,N_310);
nand U1228 (N_1228,N_43,N_487);
nor U1229 (N_1229,N_507,N_430);
and U1230 (N_1230,N_108,N_426);
nor U1231 (N_1231,N_743,N_255);
or U1232 (N_1232,N_708,N_343);
nor U1233 (N_1233,N_356,N_340);
or U1234 (N_1234,N_353,N_169);
nor U1235 (N_1235,N_412,N_136);
nor U1236 (N_1236,N_450,N_310);
nor U1237 (N_1237,N_130,N_227);
and U1238 (N_1238,N_487,N_313);
nor U1239 (N_1239,N_732,N_418);
nor U1240 (N_1240,N_547,N_357);
nor U1241 (N_1241,N_369,N_637);
nor U1242 (N_1242,N_91,N_151);
and U1243 (N_1243,N_80,N_349);
nor U1244 (N_1244,N_599,N_485);
and U1245 (N_1245,N_79,N_376);
xnor U1246 (N_1246,N_504,N_286);
nand U1247 (N_1247,N_307,N_586);
nand U1248 (N_1248,N_204,N_327);
nand U1249 (N_1249,N_17,N_458);
nand U1250 (N_1250,N_462,N_58);
nand U1251 (N_1251,N_209,N_519);
xnor U1252 (N_1252,N_493,N_248);
or U1253 (N_1253,N_50,N_300);
nor U1254 (N_1254,N_334,N_573);
or U1255 (N_1255,N_509,N_148);
nor U1256 (N_1256,N_482,N_264);
xnor U1257 (N_1257,N_225,N_648);
or U1258 (N_1258,N_743,N_528);
nand U1259 (N_1259,N_90,N_270);
xnor U1260 (N_1260,N_746,N_168);
nand U1261 (N_1261,N_248,N_718);
nor U1262 (N_1262,N_249,N_190);
xnor U1263 (N_1263,N_596,N_75);
and U1264 (N_1264,N_279,N_550);
nand U1265 (N_1265,N_595,N_433);
or U1266 (N_1266,N_693,N_250);
or U1267 (N_1267,N_173,N_620);
and U1268 (N_1268,N_12,N_52);
or U1269 (N_1269,N_184,N_68);
or U1270 (N_1270,N_43,N_662);
nand U1271 (N_1271,N_511,N_198);
or U1272 (N_1272,N_331,N_580);
nor U1273 (N_1273,N_233,N_735);
nor U1274 (N_1274,N_530,N_644);
nor U1275 (N_1275,N_157,N_166);
xor U1276 (N_1276,N_268,N_71);
xor U1277 (N_1277,N_641,N_556);
and U1278 (N_1278,N_220,N_421);
nor U1279 (N_1279,N_697,N_235);
nor U1280 (N_1280,N_10,N_673);
or U1281 (N_1281,N_377,N_480);
nand U1282 (N_1282,N_230,N_104);
and U1283 (N_1283,N_229,N_624);
or U1284 (N_1284,N_443,N_154);
nor U1285 (N_1285,N_372,N_341);
nand U1286 (N_1286,N_690,N_148);
xor U1287 (N_1287,N_206,N_408);
or U1288 (N_1288,N_503,N_105);
and U1289 (N_1289,N_343,N_143);
and U1290 (N_1290,N_430,N_451);
or U1291 (N_1291,N_572,N_220);
xor U1292 (N_1292,N_89,N_138);
or U1293 (N_1293,N_716,N_33);
and U1294 (N_1294,N_743,N_542);
or U1295 (N_1295,N_121,N_350);
nor U1296 (N_1296,N_520,N_717);
nand U1297 (N_1297,N_90,N_562);
or U1298 (N_1298,N_683,N_288);
nor U1299 (N_1299,N_100,N_176);
nand U1300 (N_1300,N_644,N_323);
nand U1301 (N_1301,N_607,N_119);
nand U1302 (N_1302,N_101,N_2);
or U1303 (N_1303,N_167,N_514);
or U1304 (N_1304,N_728,N_561);
nor U1305 (N_1305,N_419,N_74);
nor U1306 (N_1306,N_115,N_142);
xor U1307 (N_1307,N_70,N_490);
and U1308 (N_1308,N_81,N_524);
nand U1309 (N_1309,N_319,N_637);
nor U1310 (N_1310,N_601,N_580);
and U1311 (N_1311,N_604,N_743);
or U1312 (N_1312,N_122,N_312);
and U1313 (N_1313,N_164,N_104);
and U1314 (N_1314,N_264,N_206);
xnor U1315 (N_1315,N_294,N_145);
and U1316 (N_1316,N_401,N_347);
nand U1317 (N_1317,N_522,N_200);
xor U1318 (N_1318,N_304,N_239);
or U1319 (N_1319,N_295,N_202);
and U1320 (N_1320,N_633,N_295);
nor U1321 (N_1321,N_738,N_524);
nand U1322 (N_1322,N_404,N_178);
nand U1323 (N_1323,N_733,N_248);
or U1324 (N_1324,N_171,N_24);
xnor U1325 (N_1325,N_663,N_475);
and U1326 (N_1326,N_478,N_266);
xnor U1327 (N_1327,N_570,N_728);
nand U1328 (N_1328,N_38,N_414);
nor U1329 (N_1329,N_113,N_717);
nor U1330 (N_1330,N_591,N_669);
or U1331 (N_1331,N_113,N_380);
and U1332 (N_1332,N_288,N_164);
nand U1333 (N_1333,N_122,N_247);
nand U1334 (N_1334,N_517,N_118);
and U1335 (N_1335,N_385,N_254);
nor U1336 (N_1336,N_460,N_205);
or U1337 (N_1337,N_235,N_99);
and U1338 (N_1338,N_293,N_12);
or U1339 (N_1339,N_266,N_500);
or U1340 (N_1340,N_400,N_312);
or U1341 (N_1341,N_635,N_157);
and U1342 (N_1342,N_627,N_293);
and U1343 (N_1343,N_699,N_71);
or U1344 (N_1344,N_503,N_51);
or U1345 (N_1345,N_523,N_584);
nand U1346 (N_1346,N_384,N_429);
or U1347 (N_1347,N_237,N_577);
and U1348 (N_1348,N_601,N_247);
nand U1349 (N_1349,N_591,N_643);
nor U1350 (N_1350,N_342,N_452);
nand U1351 (N_1351,N_437,N_14);
nand U1352 (N_1352,N_483,N_714);
nand U1353 (N_1353,N_251,N_598);
xnor U1354 (N_1354,N_269,N_331);
nand U1355 (N_1355,N_412,N_625);
or U1356 (N_1356,N_642,N_460);
or U1357 (N_1357,N_510,N_196);
xnor U1358 (N_1358,N_704,N_688);
nand U1359 (N_1359,N_45,N_169);
nor U1360 (N_1360,N_369,N_482);
or U1361 (N_1361,N_482,N_87);
nand U1362 (N_1362,N_632,N_683);
nor U1363 (N_1363,N_606,N_207);
and U1364 (N_1364,N_83,N_256);
or U1365 (N_1365,N_450,N_639);
or U1366 (N_1366,N_733,N_309);
or U1367 (N_1367,N_551,N_464);
nand U1368 (N_1368,N_211,N_567);
nor U1369 (N_1369,N_334,N_43);
nand U1370 (N_1370,N_567,N_185);
xor U1371 (N_1371,N_39,N_308);
and U1372 (N_1372,N_596,N_706);
or U1373 (N_1373,N_29,N_633);
and U1374 (N_1374,N_577,N_100);
xor U1375 (N_1375,N_420,N_301);
xnor U1376 (N_1376,N_49,N_457);
xnor U1377 (N_1377,N_214,N_384);
and U1378 (N_1378,N_661,N_666);
nand U1379 (N_1379,N_147,N_617);
nor U1380 (N_1380,N_724,N_447);
or U1381 (N_1381,N_483,N_367);
nand U1382 (N_1382,N_535,N_273);
nand U1383 (N_1383,N_649,N_43);
nand U1384 (N_1384,N_614,N_340);
or U1385 (N_1385,N_627,N_361);
nand U1386 (N_1386,N_710,N_250);
xor U1387 (N_1387,N_591,N_468);
nand U1388 (N_1388,N_307,N_18);
or U1389 (N_1389,N_241,N_659);
nand U1390 (N_1390,N_657,N_302);
xor U1391 (N_1391,N_656,N_333);
xnor U1392 (N_1392,N_599,N_43);
and U1393 (N_1393,N_15,N_718);
or U1394 (N_1394,N_246,N_577);
or U1395 (N_1395,N_584,N_28);
nand U1396 (N_1396,N_412,N_567);
nand U1397 (N_1397,N_47,N_173);
or U1398 (N_1398,N_262,N_130);
nand U1399 (N_1399,N_630,N_517);
nand U1400 (N_1400,N_175,N_345);
nand U1401 (N_1401,N_185,N_291);
and U1402 (N_1402,N_749,N_477);
or U1403 (N_1403,N_738,N_120);
xnor U1404 (N_1404,N_633,N_472);
nor U1405 (N_1405,N_432,N_370);
nor U1406 (N_1406,N_322,N_69);
or U1407 (N_1407,N_549,N_653);
nor U1408 (N_1408,N_432,N_287);
nor U1409 (N_1409,N_275,N_740);
xnor U1410 (N_1410,N_218,N_646);
and U1411 (N_1411,N_310,N_577);
xor U1412 (N_1412,N_304,N_288);
and U1413 (N_1413,N_317,N_190);
and U1414 (N_1414,N_468,N_510);
xnor U1415 (N_1415,N_605,N_738);
or U1416 (N_1416,N_487,N_602);
or U1417 (N_1417,N_435,N_530);
nand U1418 (N_1418,N_69,N_704);
and U1419 (N_1419,N_139,N_243);
nor U1420 (N_1420,N_222,N_141);
nand U1421 (N_1421,N_427,N_3);
nor U1422 (N_1422,N_383,N_487);
xor U1423 (N_1423,N_678,N_451);
or U1424 (N_1424,N_629,N_0);
xor U1425 (N_1425,N_730,N_647);
xnor U1426 (N_1426,N_539,N_580);
and U1427 (N_1427,N_610,N_316);
nand U1428 (N_1428,N_483,N_279);
and U1429 (N_1429,N_698,N_49);
xnor U1430 (N_1430,N_454,N_702);
and U1431 (N_1431,N_201,N_441);
nor U1432 (N_1432,N_445,N_689);
and U1433 (N_1433,N_88,N_699);
or U1434 (N_1434,N_488,N_109);
nor U1435 (N_1435,N_685,N_220);
nand U1436 (N_1436,N_412,N_713);
or U1437 (N_1437,N_498,N_110);
xor U1438 (N_1438,N_178,N_150);
nand U1439 (N_1439,N_77,N_451);
and U1440 (N_1440,N_131,N_324);
nand U1441 (N_1441,N_263,N_292);
xnor U1442 (N_1442,N_18,N_161);
and U1443 (N_1443,N_425,N_365);
nand U1444 (N_1444,N_447,N_75);
xnor U1445 (N_1445,N_644,N_293);
xor U1446 (N_1446,N_148,N_531);
nor U1447 (N_1447,N_205,N_125);
nor U1448 (N_1448,N_498,N_227);
nor U1449 (N_1449,N_198,N_232);
and U1450 (N_1450,N_448,N_166);
xnor U1451 (N_1451,N_653,N_496);
xor U1452 (N_1452,N_260,N_634);
nand U1453 (N_1453,N_498,N_326);
or U1454 (N_1454,N_597,N_57);
nand U1455 (N_1455,N_165,N_180);
nor U1456 (N_1456,N_88,N_560);
nand U1457 (N_1457,N_661,N_663);
nand U1458 (N_1458,N_449,N_202);
xor U1459 (N_1459,N_382,N_568);
and U1460 (N_1460,N_658,N_504);
nand U1461 (N_1461,N_659,N_117);
xnor U1462 (N_1462,N_702,N_560);
or U1463 (N_1463,N_577,N_556);
nand U1464 (N_1464,N_105,N_382);
and U1465 (N_1465,N_648,N_226);
or U1466 (N_1466,N_462,N_26);
and U1467 (N_1467,N_58,N_178);
nor U1468 (N_1468,N_619,N_394);
nor U1469 (N_1469,N_652,N_516);
or U1470 (N_1470,N_517,N_213);
or U1471 (N_1471,N_658,N_358);
nand U1472 (N_1472,N_468,N_87);
xor U1473 (N_1473,N_186,N_466);
and U1474 (N_1474,N_121,N_352);
nand U1475 (N_1475,N_26,N_393);
and U1476 (N_1476,N_298,N_437);
xnor U1477 (N_1477,N_723,N_549);
nand U1478 (N_1478,N_731,N_502);
and U1479 (N_1479,N_477,N_22);
nor U1480 (N_1480,N_261,N_672);
nand U1481 (N_1481,N_459,N_131);
and U1482 (N_1482,N_639,N_382);
or U1483 (N_1483,N_673,N_229);
xor U1484 (N_1484,N_527,N_20);
and U1485 (N_1485,N_522,N_648);
and U1486 (N_1486,N_436,N_55);
nor U1487 (N_1487,N_64,N_607);
nand U1488 (N_1488,N_20,N_575);
or U1489 (N_1489,N_701,N_182);
or U1490 (N_1490,N_403,N_347);
or U1491 (N_1491,N_679,N_528);
nor U1492 (N_1492,N_617,N_608);
nor U1493 (N_1493,N_269,N_372);
or U1494 (N_1494,N_605,N_98);
and U1495 (N_1495,N_49,N_243);
xor U1496 (N_1496,N_429,N_195);
nor U1497 (N_1497,N_51,N_311);
or U1498 (N_1498,N_12,N_72);
xnor U1499 (N_1499,N_592,N_437);
nor U1500 (N_1500,N_852,N_1159);
nor U1501 (N_1501,N_1380,N_1401);
xor U1502 (N_1502,N_808,N_906);
and U1503 (N_1503,N_1381,N_1126);
or U1504 (N_1504,N_1449,N_787);
nor U1505 (N_1505,N_943,N_1193);
nor U1506 (N_1506,N_866,N_820);
xor U1507 (N_1507,N_1135,N_1090);
nand U1508 (N_1508,N_1254,N_1334);
or U1509 (N_1509,N_809,N_1057);
or U1510 (N_1510,N_1013,N_1215);
and U1511 (N_1511,N_839,N_833);
and U1512 (N_1512,N_991,N_776);
nand U1513 (N_1513,N_1205,N_1197);
or U1514 (N_1514,N_1257,N_1469);
or U1515 (N_1515,N_1294,N_1123);
and U1516 (N_1516,N_1129,N_941);
nand U1517 (N_1517,N_965,N_1041);
nor U1518 (N_1518,N_881,N_816);
and U1519 (N_1519,N_1183,N_929);
or U1520 (N_1520,N_1406,N_1221);
nand U1521 (N_1521,N_1371,N_978);
nor U1522 (N_1522,N_824,N_1244);
nand U1523 (N_1523,N_910,N_757);
or U1524 (N_1524,N_1264,N_1149);
or U1525 (N_1525,N_834,N_1299);
xnor U1526 (N_1526,N_1204,N_1063);
or U1527 (N_1527,N_972,N_1014);
nor U1528 (N_1528,N_952,N_1166);
nor U1529 (N_1529,N_956,N_1341);
xnor U1530 (N_1530,N_781,N_1106);
or U1531 (N_1531,N_1317,N_1258);
or U1532 (N_1532,N_1100,N_803);
and U1533 (N_1533,N_1280,N_913);
nor U1534 (N_1534,N_1496,N_990);
nand U1535 (N_1535,N_1376,N_1297);
xor U1536 (N_1536,N_815,N_926);
and U1537 (N_1537,N_999,N_1411);
xor U1538 (N_1538,N_1404,N_848);
nor U1539 (N_1539,N_765,N_873);
nand U1540 (N_1540,N_1219,N_868);
nor U1541 (N_1541,N_1246,N_1218);
nor U1542 (N_1542,N_1102,N_1421);
nor U1543 (N_1543,N_1316,N_1058);
or U1544 (N_1544,N_1048,N_1473);
xor U1545 (N_1545,N_905,N_1354);
nor U1546 (N_1546,N_1360,N_779);
xor U1547 (N_1547,N_1247,N_1187);
or U1548 (N_1548,N_1277,N_1462);
xor U1549 (N_1549,N_1253,N_1353);
nand U1550 (N_1550,N_1049,N_1038);
nand U1551 (N_1551,N_760,N_751);
or U1552 (N_1552,N_826,N_1429);
or U1553 (N_1553,N_800,N_1452);
and U1554 (N_1554,N_932,N_1260);
xnor U1555 (N_1555,N_789,N_1078);
and U1556 (N_1556,N_992,N_1117);
nor U1557 (N_1557,N_957,N_1263);
nand U1558 (N_1558,N_769,N_752);
or U1559 (N_1559,N_1392,N_1410);
and U1560 (N_1560,N_1298,N_1236);
xnor U1561 (N_1561,N_1111,N_1467);
nor U1562 (N_1562,N_1202,N_1136);
and U1563 (N_1563,N_1201,N_1385);
nor U1564 (N_1564,N_1115,N_1364);
nand U1565 (N_1565,N_1175,N_1143);
and U1566 (N_1566,N_1224,N_1032);
xnor U1567 (N_1567,N_801,N_1080);
and U1568 (N_1568,N_1366,N_1286);
xor U1569 (N_1569,N_1147,N_1110);
or U1570 (N_1570,N_1255,N_1397);
xnor U1571 (N_1571,N_1169,N_1245);
and U1572 (N_1572,N_1284,N_854);
nand U1573 (N_1573,N_1448,N_1016);
and U1574 (N_1574,N_1367,N_918);
nand U1575 (N_1575,N_1271,N_1304);
nor U1576 (N_1576,N_1209,N_1060);
nand U1577 (N_1577,N_1153,N_890);
nand U1578 (N_1578,N_1004,N_1262);
or U1579 (N_1579,N_782,N_1142);
nor U1580 (N_1580,N_1233,N_1389);
xnor U1581 (N_1581,N_1118,N_773);
nand U1582 (N_1582,N_1107,N_1015);
and U1583 (N_1583,N_1116,N_870);
nand U1584 (N_1584,N_1382,N_1195);
nand U1585 (N_1585,N_1140,N_1192);
xnor U1586 (N_1586,N_1039,N_897);
and U1587 (N_1587,N_1177,N_823);
nor U1588 (N_1588,N_1231,N_953);
xnor U1589 (N_1589,N_1009,N_1314);
nor U1590 (N_1590,N_994,N_1082);
nand U1591 (N_1591,N_1040,N_1295);
or U1592 (N_1592,N_1091,N_1127);
and U1593 (N_1593,N_964,N_1340);
nand U1594 (N_1594,N_844,N_963);
xnor U1595 (N_1595,N_1173,N_1083);
nand U1596 (N_1596,N_960,N_1332);
and U1597 (N_1597,N_1076,N_1164);
nor U1598 (N_1598,N_1229,N_850);
or U1599 (N_1599,N_1368,N_1031);
nor U1600 (N_1600,N_777,N_1276);
and U1601 (N_1601,N_1240,N_1268);
nand U1602 (N_1602,N_1120,N_1069);
and U1603 (N_1603,N_1343,N_1388);
nor U1604 (N_1604,N_1045,N_998);
nor U1605 (N_1605,N_1451,N_1266);
nand U1606 (N_1606,N_1480,N_1170);
nor U1607 (N_1607,N_1270,N_1222);
or U1608 (N_1608,N_1497,N_1103);
nand U1609 (N_1609,N_946,N_1121);
nand U1610 (N_1610,N_1182,N_851);
xor U1611 (N_1611,N_1033,N_754);
nor U1612 (N_1612,N_1163,N_967);
xor U1613 (N_1613,N_1042,N_1279);
and U1614 (N_1614,N_970,N_1490);
and U1615 (N_1615,N_1064,N_814);
xor U1616 (N_1616,N_1134,N_898);
nor U1617 (N_1617,N_1035,N_1239);
nand U1618 (N_1618,N_1085,N_1407);
nor U1619 (N_1619,N_1252,N_1450);
xor U1620 (N_1620,N_836,N_786);
and U1621 (N_1621,N_1198,N_971);
xnor U1622 (N_1622,N_841,N_1386);
and U1623 (N_1623,N_908,N_1191);
or U1624 (N_1624,N_778,N_1171);
nand U1625 (N_1625,N_987,N_899);
or U1626 (N_1626,N_1403,N_1384);
and U1627 (N_1627,N_1423,N_1161);
or U1628 (N_1628,N_1321,N_1241);
or U1629 (N_1629,N_853,N_1303);
or U1630 (N_1630,N_1465,N_1089);
and U1631 (N_1631,N_1399,N_1379);
or U1632 (N_1632,N_1178,N_1457);
or U1633 (N_1633,N_822,N_1409);
xor U1634 (N_1634,N_1413,N_1408);
xnor U1635 (N_1635,N_1088,N_1176);
and U1636 (N_1636,N_1318,N_1155);
or U1637 (N_1637,N_1017,N_864);
and U1638 (N_1638,N_849,N_1207);
nor U1639 (N_1639,N_1483,N_1481);
xnor U1640 (N_1640,N_920,N_931);
xnor U1641 (N_1641,N_1055,N_1005);
nand U1642 (N_1642,N_753,N_1075);
and U1643 (N_1643,N_1488,N_1003);
xnor U1644 (N_1644,N_919,N_1212);
nand U1645 (N_1645,N_1156,N_791);
and U1646 (N_1646,N_805,N_1025);
and U1647 (N_1647,N_887,N_966);
nand U1648 (N_1648,N_1211,N_774);
and U1649 (N_1649,N_1044,N_1414);
or U1650 (N_1650,N_1333,N_1351);
or U1651 (N_1651,N_1208,N_1238);
and U1652 (N_1652,N_871,N_1455);
nand U1653 (N_1653,N_955,N_958);
or U1654 (N_1654,N_980,N_792);
or U1655 (N_1655,N_1030,N_817);
or U1656 (N_1656,N_1174,N_889);
nor U1657 (N_1657,N_1307,N_1369);
xnor U1658 (N_1658,N_1348,N_1259);
xor U1659 (N_1659,N_780,N_1227);
and U1660 (N_1660,N_1151,N_1223);
xnor U1661 (N_1661,N_917,N_825);
nand U1662 (N_1662,N_1415,N_1289);
nor U1663 (N_1663,N_790,N_1188);
or U1664 (N_1664,N_856,N_1491);
and U1665 (N_1665,N_1036,N_842);
or U1666 (N_1666,N_1096,N_764);
nor U1667 (N_1667,N_831,N_1475);
nor U1668 (N_1668,N_1027,N_907);
and U1669 (N_1669,N_1137,N_861);
nor U1670 (N_1670,N_1010,N_1417);
and U1671 (N_1671,N_1431,N_1154);
nor U1672 (N_1672,N_1002,N_988);
xor U1673 (N_1673,N_1402,N_1352);
or U1674 (N_1674,N_1056,N_916);
nand U1675 (N_1675,N_968,N_986);
and U1676 (N_1676,N_1337,N_1186);
nor U1677 (N_1677,N_1302,N_1220);
and U1678 (N_1678,N_1290,N_981);
and U1679 (N_1679,N_912,N_896);
nand U1680 (N_1680,N_974,N_1374);
nand U1681 (N_1681,N_894,N_1378);
and U1682 (N_1682,N_1152,N_1052);
nor U1683 (N_1683,N_1144,N_1130);
xnor U1684 (N_1684,N_865,N_1301);
or U1685 (N_1685,N_1439,N_909);
xor U1686 (N_1686,N_797,N_796);
or U1687 (N_1687,N_1288,N_1084);
or U1688 (N_1688,N_1007,N_904);
or U1689 (N_1689,N_1034,N_1489);
nor U1690 (N_1690,N_788,N_1335);
xnor U1691 (N_1691,N_828,N_959);
nand U1692 (N_1692,N_1158,N_1459);
nor U1693 (N_1693,N_1206,N_1495);
and U1694 (N_1694,N_798,N_1037);
or U1695 (N_1695,N_768,N_892);
xor U1696 (N_1696,N_872,N_1420);
or U1697 (N_1697,N_942,N_1319);
xnor U1698 (N_1698,N_1243,N_767);
xnor U1699 (N_1699,N_1365,N_1092);
or U1700 (N_1700,N_883,N_1453);
and U1701 (N_1701,N_1047,N_1426);
xor U1702 (N_1702,N_1165,N_1363);
nor U1703 (N_1703,N_1493,N_1375);
or U1704 (N_1704,N_984,N_1086);
or U1705 (N_1705,N_802,N_880);
and U1706 (N_1706,N_1430,N_1291);
nor U1707 (N_1707,N_1274,N_1425);
nand U1708 (N_1708,N_785,N_1326);
and U1709 (N_1709,N_1168,N_1342);
xor U1710 (N_1710,N_1199,N_1296);
nand U1711 (N_1711,N_1070,N_1235);
or U1712 (N_1712,N_1466,N_1306);
nand U1713 (N_1713,N_840,N_1492);
nand U1714 (N_1714,N_1101,N_1437);
nor U1715 (N_1715,N_1249,N_1396);
nor U1716 (N_1716,N_1418,N_784);
nand U1717 (N_1717,N_879,N_1463);
or U1718 (N_1718,N_921,N_1099);
nor U1719 (N_1719,N_903,N_982);
xor U1720 (N_1720,N_1338,N_1067);
nor U1721 (N_1721,N_930,N_867);
nor U1722 (N_1722,N_1019,N_1000);
or U1723 (N_1723,N_857,N_1441);
or U1724 (N_1724,N_1024,N_1383);
or U1725 (N_1725,N_1398,N_1022);
nor U1726 (N_1726,N_1131,N_821);
or U1727 (N_1727,N_1471,N_933);
and U1728 (N_1728,N_1427,N_975);
nand U1729 (N_1729,N_1146,N_1356);
xnor U1730 (N_1730,N_1324,N_900);
or U1731 (N_1731,N_1028,N_1095);
nand U1732 (N_1732,N_979,N_1395);
and U1733 (N_1733,N_914,N_1109);
nor U1734 (N_1734,N_1065,N_969);
or U1735 (N_1735,N_911,N_1145);
and U1736 (N_1736,N_1355,N_949);
xor U1737 (N_1737,N_924,N_961);
nor U1738 (N_1738,N_1062,N_1237);
nand U1739 (N_1739,N_1460,N_1189);
nor U1740 (N_1740,N_1098,N_995);
or U1741 (N_1741,N_1112,N_838);
and U1742 (N_1742,N_799,N_1203);
and U1743 (N_1743,N_761,N_1446);
nor U1744 (N_1744,N_1432,N_1422);
xnor U1745 (N_1745,N_1454,N_877);
nand U1746 (N_1746,N_1050,N_1292);
nor U1747 (N_1747,N_1468,N_1445);
xor U1748 (N_1748,N_1331,N_1440);
xnor U1749 (N_1749,N_1323,N_1438);
and U1750 (N_1750,N_1357,N_1479);
or U1751 (N_1751,N_1456,N_1272);
or U1752 (N_1752,N_795,N_869);
or U1753 (N_1753,N_1287,N_948);
nor U1754 (N_1754,N_1011,N_1470);
and U1755 (N_1755,N_1234,N_1119);
nor U1756 (N_1756,N_1315,N_1350);
or U1757 (N_1757,N_1248,N_1419);
nor U1758 (N_1758,N_885,N_1486);
nor U1759 (N_1759,N_1128,N_1278);
or U1760 (N_1760,N_1387,N_1059);
nor U1761 (N_1761,N_1458,N_810);
nand U1762 (N_1762,N_886,N_1179);
nand U1763 (N_1763,N_770,N_813);
nor U1764 (N_1764,N_1180,N_1499);
nor U1765 (N_1765,N_1400,N_1461);
xor U1766 (N_1766,N_1074,N_1167);
nand U1767 (N_1767,N_1051,N_771);
nand U1768 (N_1768,N_1442,N_1113);
or U1769 (N_1769,N_750,N_1424);
nand U1770 (N_1770,N_811,N_1225);
or U1771 (N_1771,N_1079,N_1281);
nand U1772 (N_1772,N_1393,N_1097);
or U1773 (N_1773,N_858,N_1018);
nand U1774 (N_1774,N_1066,N_1213);
nor U1775 (N_1775,N_1020,N_1251);
and U1776 (N_1776,N_843,N_1308);
nand U1777 (N_1777,N_1444,N_1447);
and U1778 (N_1778,N_1132,N_1310);
and U1779 (N_1779,N_891,N_862);
nor U1780 (N_1780,N_1217,N_1162);
and U1781 (N_1781,N_1464,N_902);
xnor U1782 (N_1782,N_1072,N_1157);
xnor U1783 (N_1783,N_827,N_818);
or U1784 (N_1784,N_1484,N_775);
nor U1785 (N_1785,N_1122,N_1210);
nor U1786 (N_1786,N_1114,N_1185);
or U1787 (N_1787,N_938,N_1412);
nand U1788 (N_1788,N_1359,N_1196);
nand U1789 (N_1789,N_1327,N_1309);
or U1790 (N_1790,N_882,N_939);
or U1791 (N_1791,N_1023,N_766);
and U1792 (N_1792,N_837,N_951);
or U1793 (N_1793,N_1482,N_1008);
nor U1794 (N_1794,N_1328,N_1347);
xor U1795 (N_1795,N_1269,N_937);
xnor U1796 (N_1796,N_944,N_762);
nor U1797 (N_1797,N_1054,N_863);
xnor U1798 (N_1798,N_1267,N_1250);
or U1799 (N_1799,N_1485,N_1006);
or U1800 (N_1800,N_1133,N_989);
xnor U1801 (N_1801,N_806,N_807);
xnor U1802 (N_1802,N_1391,N_927);
or U1803 (N_1803,N_976,N_874);
nor U1804 (N_1804,N_1394,N_783);
nand U1805 (N_1805,N_993,N_1361);
or U1806 (N_1806,N_1194,N_1329);
nor U1807 (N_1807,N_940,N_1339);
nand U1808 (N_1808,N_1476,N_794);
nor U1809 (N_1809,N_1370,N_835);
or U1810 (N_1810,N_846,N_1434);
and U1811 (N_1811,N_1061,N_1273);
xor U1812 (N_1812,N_985,N_1305);
xor U1813 (N_1813,N_1081,N_1346);
nand U1814 (N_1814,N_855,N_1344);
or U1815 (N_1815,N_1325,N_1428);
nor U1816 (N_1816,N_1275,N_1474);
or U1817 (N_1817,N_830,N_923);
and U1818 (N_1818,N_1181,N_755);
or U1819 (N_1819,N_1265,N_1141);
nand U1820 (N_1820,N_884,N_1172);
nand U1821 (N_1821,N_1256,N_945);
nor U1822 (N_1822,N_1021,N_1472);
nor U1823 (N_1823,N_936,N_895);
or U1824 (N_1824,N_1190,N_1200);
nor U1825 (N_1825,N_1443,N_1077);
nand U1826 (N_1826,N_1026,N_1436);
nand U1827 (N_1827,N_759,N_878);
nand U1828 (N_1828,N_1228,N_1216);
nor U1829 (N_1829,N_977,N_1487);
xor U1830 (N_1830,N_1261,N_1073);
nor U1831 (N_1831,N_1362,N_983);
nor U1832 (N_1832,N_812,N_829);
nor U1833 (N_1833,N_1312,N_1311);
and U1834 (N_1834,N_772,N_1226);
nand U1835 (N_1835,N_947,N_1336);
nor U1836 (N_1836,N_804,N_1282);
xor U1837 (N_1837,N_1150,N_1372);
nor U1838 (N_1838,N_1087,N_1139);
nor U1839 (N_1839,N_996,N_922);
or U1840 (N_1840,N_997,N_1029);
nand U1841 (N_1841,N_1405,N_1138);
xor U1842 (N_1842,N_1320,N_1093);
nor U1843 (N_1843,N_756,N_1433);
and U1844 (N_1844,N_1313,N_888);
or U1845 (N_1845,N_845,N_1498);
nand U1846 (N_1846,N_876,N_934);
nand U1847 (N_1847,N_763,N_819);
nor U1848 (N_1848,N_1390,N_1373);
nor U1849 (N_1849,N_1494,N_1349);
or U1850 (N_1850,N_1068,N_1160);
nand U1851 (N_1851,N_954,N_1105);
nand U1852 (N_1852,N_1108,N_1345);
or U1853 (N_1853,N_1232,N_793);
and U1854 (N_1854,N_1322,N_973);
nor U1855 (N_1855,N_1148,N_1285);
xor U1856 (N_1856,N_1358,N_758);
nand U1857 (N_1857,N_1184,N_915);
or U1858 (N_1858,N_1214,N_893);
xnor U1859 (N_1859,N_950,N_847);
or U1860 (N_1860,N_935,N_1283);
nand U1861 (N_1861,N_1293,N_1124);
nor U1862 (N_1862,N_901,N_1046);
xnor U1863 (N_1863,N_875,N_1300);
or U1864 (N_1864,N_925,N_1012);
nand U1865 (N_1865,N_832,N_1053);
nor U1866 (N_1866,N_1125,N_1330);
and U1867 (N_1867,N_1377,N_1435);
and U1868 (N_1868,N_1001,N_928);
nand U1869 (N_1869,N_1478,N_1242);
nand U1870 (N_1870,N_1477,N_1094);
nor U1871 (N_1871,N_1043,N_1416);
and U1872 (N_1872,N_859,N_1071);
xnor U1873 (N_1873,N_962,N_860);
xor U1874 (N_1874,N_1104,N_1230);
nand U1875 (N_1875,N_979,N_771);
nor U1876 (N_1876,N_900,N_947);
nor U1877 (N_1877,N_979,N_1215);
and U1878 (N_1878,N_1432,N_1220);
xnor U1879 (N_1879,N_879,N_891);
xnor U1880 (N_1880,N_1048,N_814);
nand U1881 (N_1881,N_1368,N_1433);
and U1882 (N_1882,N_1273,N_1092);
or U1883 (N_1883,N_1057,N_1122);
and U1884 (N_1884,N_1004,N_1488);
nand U1885 (N_1885,N_1070,N_1154);
or U1886 (N_1886,N_875,N_820);
and U1887 (N_1887,N_1014,N_1407);
or U1888 (N_1888,N_1361,N_946);
nand U1889 (N_1889,N_1232,N_1395);
xnor U1890 (N_1890,N_1070,N_918);
and U1891 (N_1891,N_1041,N_988);
and U1892 (N_1892,N_1170,N_929);
nor U1893 (N_1893,N_912,N_1428);
and U1894 (N_1894,N_1047,N_840);
or U1895 (N_1895,N_1312,N_858);
and U1896 (N_1896,N_1177,N_1083);
and U1897 (N_1897,N_883,N_1473);
or U1898 (N_1898,N_913,N_906);
or U1899 (N_1899,N_1158,N_930);
nand U1900 (N_1900,N_1486,N_1411);
nand U1901 (N_1901,N_854,N_1009);
nor U1902 (N_1902,N_1204,N_1401);
and U1903 (N_1903,N_1014,N_1021);
xor U1904 (N_1904,N_1488,N_944);
or U1905 (N_1905,N_839,N_919);
or U1906 (N_1906,N_835,N_888);
and U1907 (N_1907,N_1023,N_1226);
nand U1908 (N_1908,N_974,N_1420);
and U1909 (N_1909,N_1206,N_1499);
nand U1910 (N_1910,N_1244,N_1015);
nor U1911 (N_1911,N_824,N_994);
and U1912 (N_1912,N_832,N_1275);
nand U1913 (N_1913,N_817,N_1118);
and U1914 (N_1914,N_1371,N_1318);
xor U1915 (N_1915,N_1439,N_1366);
nand U1916 (N_1916,N_893,N_1345);
nand U1917 (N_1917,N_1191,N_886);
nor U1918 (N_1918,N_1049,N_1302);
and U1919 (N_1919,N_950,N_811);
nor U1920 (N_1920,N_1235,N_1190);
and U1921 (N_1921,N_1266,N_1311);
nand U1922 (N_1922,N_1049,N_1259);
and U1923 (N_1923,N_1351,N_1357);
xnor U1924 (N_1924,N_890,N_1212);
nor U1925 (N_1925,N_1395,N_1241);
xnor U1926 (N_1926,N_1201,N_1331);
nor U1927 (N_1927,N_961,N_818);
and U1928 (N_1928,N_932,N_850);
or U1929 (N_1929,N_823,N_804);
xor U1930 (N_1930,N_872,N_1384);
nand U1931 (N_1931,N_903,N_1017);
nand U1932 (N_1932,N_980,N_1150);
nor U1933 (N_1933,N_1159,N_1452);
and U1934 (N_1934,N_979,N_1156);
nor U1935 (N_1935,N_1462,N_1302);
and U1936 (N_1936,N_1266,N_833);
or U1937 (N_1937,N_997,N_1444);
or U1938 (N_1938,N_930,N_906);
nand U1939 (N_1939,N_1068,N_1125);
or U1940 (N_1940,N_1069,N_1448);
nor U1941 (N_1941,N_1309,N_1449);
or U1942 (N_1942,N_1056,N_877);
xor U1943 (N_1943,N_855,N_996);
and U1944 (N_1944,N_1213,N_1420);
nand U1945 (N_1945,N_770,N_960);
nor U1946 (N_1946,N_1490,N_1447);
and U1947 (N_1947,N_865,N_1171);
xnor U1948 (N_1948,N_1476,N_1068);
nor U1949 (N_1949,N_1450,N_1277);
or U1950 (N_1950,N_1396,N_1269);
xnor U1951 (N_1951,N_1243,N_1003);
xor U1952 (N_1952,N_1407,N_867);
xor U1953 (N_1953,N_934,N_1157);
and U1954 (N_1954,N_928,N_1110);
nand U1955 (N_1955,N_1200,N_1392);
nor U1956 (N_1956,N_947,N_890);
nor U1957 (N_1957,N_824,N_802);
xnor U1958 (N_1958,N_1249,N_917);
and U1959 (N_1959,N_960,N_1120);
nor U1960 (N_1960,N_1489,N_1094);
and U1961 (N_1961,N_929,N_1093);
and U1962 (N_1962,N_1406,N_889);
nand U1963 (N_1963,N_1019,N_1198);
xor U1964 (N_1964,N_1092,N_1268);
nor U1965 (N_1965,N_921,N_1258);
and U1966 (N_1966,N_1267,N_781);
xnor U1967 (N_1967,N_868,N_904);
or U1968 (N_1968,N_839,N_1326);
nand U1969 (N_1969,N_1163,N_1430);
and U1970 (N_1970,N_813,N_1305);
or U1971 (N_1971,N_1061,N_1498);
xor U1972 (N_1972,N_1107,N_913);
nor U1973 (N_1973,N_808,N_940);
nor U1974 (N_1974,N_1185,N_1076);
or U1975 (N_1975,N_1039,N_1191);
nor U1976 (N_1976,N_934,N_845);
or U1977 (N_1977,N_993,N_1056);
nand U1978 (N_1978,N_970,N_1432);
nand U1979 (N_1979,N_1302,N_1340);
xor U1980 (N_1980,N_863,N_1269);
nand U1981 (N_1981,N_1046,N_1214);
and U1982 (N_1982,N_852,N_774);
nand U1983 (N_1983,N_1440,N_969);
nor U1984 (N_1984,N_1378,N_1297);
nand U1985 (N_1985,N_1377,N_981);
nor U1986 (N_1986,N_1428,N_1252);
and U1987 (N_1987,N_1472,N_1469);
or U1988 (N_1988,N_1030,N_1125);
nand U1989 (N_1989,N_783,N_944);
and U1990 (N_1990,N_1243,N_1177);
and U1991 (N_1991,N_1485,N_1041);
or U1992 (N_1992,N_830,N_1127);
nand U1993 (N_1993,N_764,N_1141);
or U1994 (N_1994,N_909,N_1123);
and U1995 (N_1995,N_874,N_925);
xnor U1996 (N_1996,N_786,N_986);
nand U1997 (N_1997,N_1297,N_1159);
or U1998 (N_1998,N_938,N_931);
and U1999 (N_1999,N_1109,N_836);
and U2000 (N_2000,N_918,N_1178);
xor U2001 (N_2001,N_1070,N_781);
or U2002 (N_2002,N_1422,N_888);
xor U2003 (N_2003,N_1273,N_928);
or U2004 (N_2004,N_1332,N_1297);
and U2005 (N_2005,N_790,N_1348);
or U2006 (N_2006,N_1416,N_1271);
nor U2007 (N_2007,N_1203,N_1069);
xnor U2008 (N_2008,N_803,N_1207);
or U2009 (N_2009,N_937,N_873);
nand U2010 (N_2010,N_785,N_1030);
xor U2011 (N_2011,N_973,N_753);
nand U2012 (N_2012,N_1038,N_1400);
or U2013 (N_2013,N_952,N_1305);
nor U2014 (N_2014,N_1218,N_1487);
or U2015 (N_2015,N_1402,N_1448);
or U2016 (N_2016,N_794,N_811);
and U2017 (N_2017,N_908,N_1247);
or U2018 (N_2018,N_1397,N_810);
nor U2019 (N_2019,N_1426,N_1352);
nor U2020 (N_2020,N_1393,N_781);
nor U2021 (N_2021,N_1263,N_1367);
and U2022 (N_2022,N_1111,N_868);
nor U2023 (N_2023,N_1024,N_853);
or U2024 (N_2024,N_1100,N_1382);
nor U2025 (N_2025,N_1278,N_1066);
or U2026 (N_2026,N_1313,N_1215);
nand U2027 (N_2027,N_1123,N_967);
or U2028 (N_2028,N_1287,N_1054);
or U2029 (N_2029,N_882,N_815);
and U2030 (N_2030,N_1220,N_1379);
xnor U2031 (N_2031,N_858,N_1383);
nor U2032 (N_2032,N_990,N_1325);
nand U2033 (N_2033,N_1354,N_1433);
xor U2034 (N_2034,N_1352,N_753);
xnor U2035 (N_2035,N_1236,N_906);
nand U2036 (N_2036,N_1304,N_1094);
and U2037 (N_2037,N_1308,N_1115);
xnor U2038 (N_2038,N_1341,N_966);
nand U2039 (N_2039,N_855,N_1145);
nand U2040 (N_2040,N_1115,N_907);
nand U2041 (N_2041,N_1228,N_902);
nand U2042 (N_2042,N_988,N_1107);
and U2043 (N_2043,N_1368,N_1185);
xnor U2044 (N_2044,N_1314,N_1148);
and U2045 (N_2045,N_1392,N_1216);
or U2046 (N_2046,N_1094,N_1323);
xor U2047 (N_2047,N_1222,N_1122);
xor U2048 (N_2048,N_954,N_921);
nand U2049 (N_2049,N_923,N_850);
or U2050 (N_2050,N_915,N_1486);
nand U2051 (N_2051,N_1147,N_819);
or U2052 (N_2052,N_1052,N_1405);
and U2053 (N_2053,N_1179,N_1356);
nor U2054 (N_2054,N_1318,N_1474);
and U2055 (N_2055,N_785,N_1252);
xor U2056 (N_2056,N_916,N_1163);
nor U2057 (N_2057,N_1123,N_797);
or U2058 (N_2058,N_1261,N_1240);
or U2059 (N_2059,N_811,N_1321);
nand U2060 (N_2060,N_1479,N_864);
or U2061 (N_2061,N_1418,N_1083);
nor U2062 (N_2062,N_833,N_1489);
nand U2063 (N_2063,N_1051,N_838);
xor U2064 (N_2064,N_979,N_1377);
xor U2065 (N_2065,N_1330,N_759);
nor U2066 (N_2066,N_1153,N_837);
nand U2067 (N_2067,N_1364,N_1200);
xnor U2068 (N_2068,N_863,N_1156);
nand U2069 (N_2069,N_1428,N_985);
and U2070 (N_2070,N_1288,N_1428);
nand U2071 (N_2071,N_1094,N_836);
nand U2072 (N_2072,N_1060,N_904);
nor U2073 (N_2073,N_1350,N_986);
or U2074 (N_2074,N_949,N_1116);
nor U2075 (N_2075,N_1016,N_916);
and U2076 (N_2076,N_1276,N_933);
nor U2077 (N_2077,N_1245,N_1417);
nor U2078 (N_2078,N_1418,N_1123);
nor U2079 (N_2079,N_1326,N_1120);
nor U2080 (N_2080,N_1322,N_1185);
and U2081 (N_2081,N_1129,N_1213);
nor U2082 (N_2082,N_1174,N_977);
nor U2083 (N_2083,N_758,N_828);
xnor U2084 (N_2084,N_1273,N_997);
nand U2085 (N_2085,N_1216,N_1297);
and U2086 (N_2086,N_1481,N_1274);
xor U2087 (N_2087,N_1176,N_1240);
or U2088 (N_2088,N_1100,N_785);
nor U2089 (N_2089,N_1135,N_1408);
or U2090 (N_2090,N_758,N_1075);
or U2091 (N_2091,N_1408,N_881);
nand U2092 (N_2092,N_1456,N_971);
xnor U2093 (N_2093,N_1300,N_1414);
nor U2094 (N_2094,N_1098,N_1277);
nor U2095 (N_2095,N_819,N_1105);
nor U2096 (N_2096,N_865,N_1388);
and U2097 (N_2097,N_866,N_1327);
xnor U2098 (N_2098,N_1020,N_1192);
or U2099 (N_2099,N_1349,N_1279);
or U2100 (N_2100,N_858,N_1469);
nand U2101 (N_2101,N_972,N_1191);
xnor U2102 (N_2102,N_1180,N_1282);
or U2103 (N_2103,N_902,N_1310);
nand U2104 (N_2104,N_1105,N_990);
xnor U2105 (N_2105,N_1014,N_862);
or U2106 (N_2106,N_1043,N_1446);
nand U2107 (N_2107,N_1138,N_809);
nand U2108 (N_2108,N_1261,N_1481);
nand U2109 (N_2109,N_1436,N_1325);
and U2110 (N_2110,N_1074,N_1424);
or U2111 (N_2111,N_1320,N_1258);
and U2112 (N_2112,N_1058,N_1154);
nor U2113 (N_2113,N_1015,N_1463);
nand U2114 (N_2114,N_921,N_1214);
nand U2115 (N_2115,N_1371,N_1232);
xnor U2116 (N_2116,N_832,N_1482);
and U2117 (N_2117,N_1113,N_1026);
nand U2118 (N_2118,N_770,N_994);
or U2119 (N_2119,N_1311,N_1025);
nor U2120 (N_2120,N_1112,N_1412);
or U2121 (N_2121,N_1003,N_1056);
and U2122 (N_2122,N_1232,N_1106);
xnor U2123 (N_2123,N_881,N_1400);
xor U2124 (N_2124,N_802,N_980);
and U2125 (N_2125,N_1131,N_1401);
xor U2126 (N_2126,N_1356,N_1105);
and U2127 (N_2127,N_1138,N_1123);
nand U2128 (N_2128,N_1443,N_898);
nor U2129 (N_2129,N_1218,N_923);
or U2130 (N_2130,N_1312,N_1127);
xor U2131 (N_2131,N_1327,N_789);
or U2132 (N_2132,N_885,N_1204);
nor U2133 (N_2133,N_779,N_801);
or U2134 (N_2134,N_1145,N_1091);
or U2135 (N_2135,N_1151,N_935);
or U2136 (N_2136,N_1017,N_1157);
xor U2137 (N_2137,N_956,N_752);
xor U2138 (N_2138,N_794,N_1198);
nand U2139 (N_2139,N_1103,N_1059);
and U2140 (N_2140,N_948,N_829);
nand U2141 (N_2141,N_800,N_1117);
nor U2142 (N_2142,N_1009,N_776);
nand U2143 (N_2143,N_831,N_1362);
nor U2144 (N_2144,N_825,N_1425);
and U2145 (N_2145,N_1032,N_785);
nor U2146 (N_2146,N_1480,N_1128);
nand U2147 (N_2147,N_1057,N_1484);
or U2148 (N_2148,N_1391,N_857);
or U2149 (N_2149,N_1446,N_1435);
nor U2150 (N_2150,N_852,N_956);
or U2151 (N_2151,N_933,N_1042);
or U2152 (N_2152,N_1241,N_1377);
nand U2153 (N_2153,N_1487,N_912);
nand U2154 (N_2154,N_1109,N_1353);
xnor U2155 (N_2155,N_758,N_885);
nor U2156 (N_2156,N_1053,N_817);
nand U2157 (N_2157,N_1190,N_1417);
nor U2158 (N_2158,N_1129,N_872);
and U2159 (N_2159,N_1026,N_1151);
and U2160 (N_2160,N_1157,N_1451);
or U2161 (N_2161,N_1460,N_1083);
nand U2162 (N_2162,N_780,N_1129);
and U2163 (N_2163,N_1422,N_1475);
nand U2164 (N_2164,N_887,N_753);
xor U2165 (N_2165,N_1305,N_1246);
nor U2166 (N_2166,N_1451,N_1163);
nor U2167 (N_2167,N_1322,N_1308);
nor U2168 (N_2168,N_1391,N_1084);
nand U2169 (N_2169,N_1175,N_1356);
nor U2170 (N_2170,N_1464,N_1173);
nand U2171 (N_2171,N_830,N_921);
or U2172 (N_2172,N_826,N_910);
nor U2173 (N_2173,N_1311,N_981);
nor U2174 (N_2174,N_1070,N_774);
nor U2175 (N_2175,N_926,N_789);
nand U2176 (N_2176,N_1484,N_1334);
or U2177 (N_2177,N_1333,N_1353);
xor U2178 (N_2178,N_1387,N_797);
nand U2179 (N_2179,N_856,N_1142);
and U2180 (N_2180,N_1464,N_954);
xor U2181 (N_2181,N_904,N_1427);
and U2182 (N_2182,N_1482,N_850);
nand U2183 (N_2183,N_1319,N_1109);
xor U2184 (N_2184,N_1328,N_867);
xor U2185 (N_2185,N_958,N_1481);
and U2186 (N_2186,N_1414,N_1384);
nand U2187 (N_2187,N_1085,N_1371);
xnor U2188 (N_2188,N_1434,N_1171);
nor U2189 (N_2189,N_1169,N_1058);
xor U2190 (N_2190,N_1181,N_1375);
nor U2191 (N_2191,N_1039,N_1402);
xor U2192 (N_2192,N_1380,N_821);
or U2193 (N_2193,N_1203,N_1053);
nand U2194 (N_2194,N_1499,N_1174);
and U2195 (N_2195,N_1238,N_808);
nand U2196 (N_2196,N_1129,N_1142);
and U2197 (N_2197,N_1199,N_815);
and U2198 (N_2198,N_1240,N_1146);
nor U2199 (N_2199,N_862,N_786);
and U2200 (N_2200,N_1025,N_907);
or U2201 (N_2201,N_793,N_934);
nand U2202 (N_2202,N_916,N_962);
and U2203 (N_2203,N_1266,N_796);
and U2204 (N_2204,N_804,N_800);
nor U2205 (N_2205,N_1149,N_1198);
nor U2206 (N_2206,N_1340,N_983);
xor U2207 (N_2207,N_1291,N_756);
and U2208 (N_2208,N_1094,N_866);
and U2209 (N_2209,N_793,N_941);
nand U2210 (N_2210,N_1148,N_1153);
or U2211 (N_2211,N_1474,N_1261);
xor U2212 (N_2212,N_1069,N_997);
or U2213 (N_2213,N_1155,N_1431);
and U2214 (N_2214,N_1058,N_1049);
and U2215 (N_2215,N_993,N_1140);
and U2216 (N_2216,N_1405,N_1273);
nand U2217 (N_2217,N_1158,N_1472);
and U2218 (N_2218,N_1469,N_871);
xor U2219 (N_2219,N_1035,N_1494);
or U2220 (N_2220,N_1415,N_1320);
and U2221 (N_2221,N_1119,N_1379);
xor U2222 (N_2222,N_1298,N_1158);
xor U2223 (N_2223,N_1270,N_813);
and U2224 (N_2224,N_1060,N_1320);
nand U2225 (N_2225,N_1066,N_924);
and U2226 (N_2226,N_1394,N_969);
nand U2227 (N_2227,N_1196,N_1355);
nand U2228 (N_2228,N_1361,N_778);
nand U2229 (N_2229,N_868,N_768);
nand U2230 (N_2230,N_1147,N_815);
or U2231 (N_2231,N_810,N_916);
nand U2232 (N_2232,N_866,N_1280);
nand U2233 (N_2233,N_853,N_807);
nor U2234 (N_2234,N_995,N_946);
and U2235 (N_2235,N_1072,N_1027);
nand U2236 (N_2236,N_1397,N_1328);
and U2237 (N_2237,N_1182,N_966);
nand U2238 (N_2238,N_1098,N_1128);
nor U2239 (N_2239,N_1129,N_1412);
and U2240 (N_2240,N_1129,N_1400);
or U2241 (N_2241,N_1017,N_1192);
and U2242 (N_2242,N_1167,N_818);
and U2243 (N_2243,N_1264,N_1451);
or U2244 (N_2244,N_1257,N_1443);
nand U2245 (N_2245,N_1080,N_1377);
xnor U2246 (N_2246,N_1491,N_1352);
nor U2247 (N_2247,N_1004,N_1348);
and U2248 (N_2248,N_812,N_814);
and U2249 (N_2249,N_945,N_1370);
xor U2250 (N_2250,N_2201,N_2012);
or U2251 (N_2251,N_2047,N_2074);
and U2252 (N_2252,N_1938,N_1772);
nor U2253 (N_2253,N_2000,N_2243);
and U2254 (N_2254,N_1936,N_2184);
nor U2255 (N_2255,N_1946,N_1578);
and U2256 (N_2256,N_1674,N_1978);
and U2257 (N_2257,N_1547,N_2085);
and U2258 (N_2258,N_1876,N_1802);
or U2259 (N_2259,N_2109,N_2211);
or U2260 (N_2260,N_2023,N_2155);
xnor U2261 (N_2261,N_1859,N_1537);
nand U2262 (N_2262,N_1786,N_1755);
and U2263 (N_2263,N_2081,N_2038);
nand U2264 (N_2264,N_2215,N_1628);
and U2265 (N_2265,N_1751,N_2236);
or U2266 (N_2266,N_1992,N_1903);
nor U2267 (N_2267,N_1892,N_1721);
nand U2268 (N_2268,N_1618,N_1744);
xnor U2269 (N_2269,N_2135,N_2193);
and U2270 (N_2270,N_1826,N_2159);
nor U2271 (N_2271,N_1595,N_1987);
xor U2272 (N_2272,N_1944,N_2098);
nand U2273 (N_2273,N_1838,N_1503);
nor U2274 (N_2274,N_1932,N_2156);
nor U2275 (N_2275,N_2099,N_1644);
or U2276 (N_2276,N_1544,N_1658);
and U2277 (N_2277,N_1779,N_1750);
xor U2278 (N_2278,N_2041,N_1553);
or U2279 (N_2279,N_2249,N_1507);
and U2280 (N_2280,N_1704,N_2051);
xor U2281 (N_2281,N_1919,N_1549);
nand U2282 (N_2282,N_1716,N_1841);
nand U2283 (N_2283,N_2197,N_1860);
xor U2284 (N_2284,N_1734,N_1599);
or U2285 (N_2285,N_2227,N_2210);
or U2286 (N_2286,N_2168,N_1741);
nand U2287 (N_2287,N_1965,N_1848);
and U2288 (N_2288,N_1951,N_1960);
or U2289 (N_2289,N_2108,N_2030);
or U2290 (N_2290,N_1579,N_1823);
nand U2291 (N_2291,N_1693,N_1817);
or U2292 (N_2292,N_1580,N_1761);
xor U2293 (N_2293,N_1527,N_1943);
nand U2294 (N_2294,N_2224,N_1651);
xnor U2295 (N_2295,N_1656,N_2001);
nor U2296 (N_2296,N_1830,N_2175);
and U2297 (N_2297,N_2142,N_1587);
or U2298 (N_2298,N_2191,N_2077);
nor U2299 (N_2299,N_1519,N_1542);
nor U2300 (N_2300,N_2134,N_1552);
xnor U2301 (N_2301,N_1514,N_2082);
nor U2302 (N_2302,N_1945,N_2061);
nand U2303 (N_2303,N_2186,N_1735);
nand U2304 (N_2304,N_2006,N_1783);
nor U2305 (N_2305,N_1767,N_1774);
and U2306 (N_2306,N_1554,N_1954);
nor U2307 (N_2307,N_2036,N_1781);
nand U2308 (N_2308,N_1714,N_1866);
nor U2309 (N_2309,N_1934,N_2127);
nor U2310 (N_2310,N_2054,N_1921);
or U2311 (N_2311,N_2217,N_1760);
nand U2312 (N_2312,N_1849,N_1792);
nand U2313 (N_2313,N_1950,N_2086);
nand U2314 (N_2314,N_2037,N_1613);
nand U2315 (N_2315,N_1728,N_1685);
nor U2316 (N_2316,N_2183,N_2221);
and U2317 (N_2317,N_2160,N_1652);
nand U2318 (N_2318,N_1971,N_1726);
or U2319 (N_2319,N_1602,N_2066);
and U2320 (N_2320,N_2045,N_1785);
and U2321 (N_2321,N_1626,N_1835);
nor U2322 (N_2322,N_2237,N_1521);
nand U2323 (N_2323,N_1898,N_2005);
xnor U2324 (N_2324,N_1679,N_1655);
nand U2325 (N_2325,N_1840,N_1907);
nand U2326 (N_2326,N_1717,N_1829);
and U2327 (N_2327,N_2130,N_1900);
and U2328 (N_2328,N_1536,N_2044);
or U2329 (N_2329,N_1627,N_2122);
and U2330 (N_2330,N_1962,N_1584);
and U2331 (N_2331,N_1530,N_2234);
nor U2332 (N_2332,N_1798,N_1757);
nor U2333 (N_2333,N_1790,N_1766);
or U2334 (N_2334,N_1605,N_1522);
xor U2335 (N_2335,N_1935,N_2091);
or U2336 (N_2336,N_2039,N_2178);
nand U2337 (N_2337,N_2080,N_1706);
or U2338 (N_2338,N_2120,N_2176);
or U2339 (N_2339,N_1740,N_1683);
nand U2340 (N_2340,N_2196,N_1601);
nand U2341 (N_2341,N_1961,N_1861);
nand U2342 (N_2342,N_2188,N_2032);
nand U2343 (N_2343,N_1502,N_2003);
or U2344 (N_2344,N_2131,N_1643);
xnor U2345 (N_2345,N_1681,N_1621);
and U2346 (N_2346,N_2223,N_1723);
or U2347 (N_2347,N_2096,N_1654);
nand U2348 (N_2348,N_2083,N_1880);
nor U2349 (N_2349,N_1756,N_1515);
or U2350 (N_2350,N_1784,N_2248);
xnor U2351 (N_2351,N_1893,N_1869);
or U2352 (N_2352,N_1853,N_1700);
nand U2353 (N_2353,N_1771,N_1668);
nor U2354 (N_2354,N_1851,N_2162);
xor U2355 (N_2355,N_1816,N_1659);
nor U2356 (N_2356,N_1606,N_1702);
nand U2357 (N_2357,N_1752,N_1633);
or U2358 (N_2358,N_2021,N_2218);
nor U2359 (N_2359,N_1671,N_1974);
xor U2360 (N_2360,N_1870,N_1972);
or U2361 (N_2361,N_1805,N_2070);
or U2362 (N_2362,N_1548,N_1812);
xor U2363 (N_2363,N_1822,N_2095);
and U2364 (N_2364,N_2157,N_1525);
and U2365 (N_2365,N_1941,N_1831);
and U2366 (N_2366,N_1885,N_2121);
nor U2367 (N_2367,N_1908,N_1947);
or U2368 (N_2368,N_1603,N_1966);
nand U2369 (N_2369,N_1543,N_1710);
or U2370 (N_2370,N_1517,N_1591);
or U2371 (N_2371,N_1576,N_1730);
nand U2372 (N_2372,N_1669,N_1989);
and U2373 (N_2373,N_2195,N_2239);
nor U2374 (N_2374,N_1864,N_1887);
nor U2375 (N_2375,N_1691,N_2125);
xor U2376 (N_2376,N_1759,N_2008);
xnor U2377 (N_2377,N_2060,N_1984);
nand U2378 (N_2378,N_2164,N_2004);
and U2379 (N_2379,N_1533,N_1589);
xor U2380 (N_2380,N_2203,N_1653);
xnor U2381 (N_2381,N_1964,N_1791);
nand U2382 (N_2382,N_2238,N_2158);
or U2383 (N_2383,N_2059,N_2089);
nand U2384 (N_2384,N_1672,N_1939);
nand U2385 (N_2385,N_2033,N_1650);
or U2386 (N_2386,N_1827,N_1695);
xor U2387 (N_2387,N_1598,N_1854);
xor U2388 (N_2388,N_1923,N_2222);
xor U2389 (N_2389,N_1764,N_2144);
nand U2390 (N_2390,N_2136,N_1857);
nor U2391 (N_2391,N_2140,N_1957);
xnor U2392 (N_2392,N_1940,N_2245);
nor U2393 (N_2393,N_1933,N_2072);
xnor U2394 (N_2394,N_2180,N_1977);
or U2395 (N_2395,N_1556,N_2209);
xnor U2396 (N_2396,N_1564,N_2213);
nand U2397 (N_2397,N_1657,N_1648);
xor U2398 (N_2398,N_1801,N_1696);
nor U2399 (N_2399,N_1809,N_1720);
or U2400 (N_2400,N_2063,N_2212);
or U2401 (N_2401,N_1763,N_1754);
or U2402 (N_2402,N_1673,N_1794);
and U2403 (N_2403,N_2010,N_2040);
nor U2404 (N_2404,N_1862,N_1890);
and U2405 (N_2405,N_1555,N_1660);
nand U2406 (N_2406,N_2171,N_2194);
and U2407 (N_2407,N_1500,N_1776);
or U2408 (N_2408,N_2035,N_1917);
nor U2409 (N_2409,N_1865,N_2152);
nand U2410 (N_2410,N_1540,N_2011);
nand U2411 (N_2411,N_1586,N_1768);
nor U2412 (N_2412,N_1909,N_1937);
xnor U2413 (N_2413,N_2244,N_2106);
nand U2414 (N_2414,N_1562,N_1677);
nor U2415 (N_2415,N_2151,N_1573);
or U2416 (N_2416,N_2019,N_2093);
or U2417 (N_2417,N_1980,N_2123);
nand U2418 (N_2418,N_1528,N_1516);
xnor U2419 (N_2419,N_1998,N_1538);
nand U2420 (N_2420,N_2103,N_2064);
xor U2421 (N_2421,N_2226,N_2124);
or U2422 (N_2422,N_2230,N_2100);
nor U2423 (N_2423,N_1845,N_1739);
and U2424 (N_2424,N_1689,N_1518);
nand U2425 (N_2425,N_2166,N_1906);
nand U2426 (N_2426,N_2220,N_1788);
and U2427 (N_2427,N_2022,N_1623);
or U2428 (N_2428,N_1567,N_1811);
nand U2429 (N_2429,N_2179,N_1748);
or U2430 (N_2430,N_1795,N_2097);
nand U2431 (N_2431,N_1871,N_2014);
nor U2432 (N_2432,N_2116,N_1868);
nor U2433 (N_2433,N_1747,N_1678);
and U2434 (N_2434,N_1534,N_2219);
nor U2435 (N_2435,N_2202,N_1523);
xor U2436 (N_2436,N_1773,N_1993);
or U2437 (N_2437,N_1886,N_1867);
xnor U2438 (N_2438,N_1545,N_1899);
or U2439 (N_2439,N_2007,N_1787);
nor U2440 (N_2440,N_1872,N_1608);
and U2441 (N_2441,N_1762,N_1782);
or U2442 (N_2442,N_1508,N_1699);
or U2443 (N_2443,N_2247,N_1824);
nand U2444 (N_2444,N_1894,N_2182);
and U2445 (N_2445,N_1570,N_2111);
or U2446 (N_2446,N_1749,N_1800);
nor U2447 (N_2447,N_2189,N_1572);
and U2448 (N_2448,N_1577,N_1692);
and U2449 (N_2449,N_1574,N_2207);
and U2450 (N_2450,N_1630,N_2174);
and U2451 (N_2451,N_1910,N_2148);
and U2452 (N_2452,N_2240,N_1922);
nand U2453 (N_2453,N_1828,N_1529);
xnor U2454 (N_2454,N_1732,N_1915);
and U2455 (N_2455,N_1632,N_1709);
and U2456 (N_2456,N_1645,N_1738);
nor U2457 (N_2457,N_1722,N_2062);
and U2458 (N_2458,N_2177,N_1982);
or U2459 (N_2459,N_2084,N_2058);
and U2460 (N_2460,N_1995,N_1511);
nor U2461 (N_2461,N_2112,N_1501);
nor U2462 (N_2462,N_1581,N_1712);
nor U2463 (N_2463,N_1724,N_1888);
nand U2464 (N_2464,N_2065,N_2110);
nor U2465 (N_2465,N_1510,N_1561);
or U2466 (N_2466,N_1955,N_1733);
and U2467 (N_2467,N_2231,N_1996);
xnor U2468 (N_2468,N_2216,N_1970);
and U2469 (N_2469,N_1551,N_2031);
or U2470 (N_2470,N_2192,N_1667);
nor U2471 (N_2471,N_1506,N_2167);
xnor U2472 (N_2472,N_1930,N_1895);
and U2473 (N_2473,N_1610,N_1807);
or U2474 (N_2474,N_1558,N_1789);
nor U2475 (N_2475,N_1560,N_1832);
xor U2476 (N_2476,N_1931,N_1877);
or U2477 (N_2477,N_1575,N_2105);
and U2478 (N_2478,N_1925,N_1825);
nor U2479 (N_2479,N_1793,N_1979);
nand U2480 (N_2480,N_1746,N_2206);
nor U2481 (N_2481,N_1881,N_2055);
nor U2482 (N_2482,N_1617,N_1858);
and U2483 (N_2483,N_1563,N_2024);
and U2484 (N_2484,N_1884,N_2009);
or U2485 (N_2485,N_1620,N_1883);
nor U2486 (N_2486,N_2026,N_1646);
nand U2487 (N_2487,N_1607,N_1916);
nand U2488 (N_2488,N_1981,N_1690);
xnor U2489 (N_2489,N_1566,N_2068);
or U2490 (N_2490,N_2119,N_2233);
nor U2491 (N_2491,N_1873,N_1670);
nand U2492 (N_2492,N_2128,N_1647);
nor U2493 (N_2493,N_2132,N_1804);
nand U2494 (N_2494,N_2088,N_2198);
nand U2495 (N_2495,N_1524,N_1532);
or U2496 (N_2496,N_2200,N_1843);
and U2497 (N_2497,N_2126,N_1808);
or U2498 (N_2498,N_1953,N_1780);
or U2499 (N_2499,N_1926,N_1684);
nor U2500 (N_2500,N_1703,N_1565);
nor U2501 (N_2501,N_1713,N_2020);
nand U2502 (N_2502,N_1636,N_1615);
nand U2503 (N_2503,N_1731,N_2092);
nand U2504 (N_2504,N_1905,N_1625);
nand U2505 (N_2505,N_1985,N_1997);
nor U2506 (N_2506,N_1707,N_1604);
nor U2507 (N_2507,N_1994,N_1663);
or U2508 (N_2508,N_2138,N_1729);
or U2509 (N_2509,N_2165,N_1844);
xnor U2510 (N_2510,N_1896,N_2228);
xnor U2511 (N_2511,N_1541,N_1638);
xnor U2512 (N_2512,N_2117,N_1622);
and U2513 (N_2513,N_2246,N_2028);
nor U2514 (N_2514,N_1639,N_2013);
nand U2515 (N_2515,N_1701,N_2149);
and U2516 (N_2516,N_1513,N_2141);
and U2517 (N_2517,N_1968,N_1836);
nor U2518 (N_2518,N_1509,N_1694);
nor U2519 (N_2519,N_1973,N_1504);
nor U2520 (N_2520,N_1879,N_1775);
and U2521 (N_2521,N_1662,N_1649);
or U2522 (N_2522,N_1818,N_1904);
and U2523 (N_2523,N_1967,N_1637);
xor U2524 (N_2524,N_1863,N_2050);
or U2525 (N_2525,N_1631,N_1594);
xor U2526 (N_2526,N_1846,N_1814);
xnor U2527 (N_2527,N_1855,N_1927);
or U2528 (N_2528,N_1778,N_1642);
nor U2529 (N_2529,N_1535,N_1986);
nor U2530 (N_2530,N_2076,N_2090);
and U2531 (N_2531,N_2046,N_1833);
and U2532 (N_2532,N_1913,N_1520);
or U2533 (N_2533,N_1718,N_1698);
nor U2534 (N_2534,N_2114,N_2027);
and U2535 (N_2535,N_1539,N_1715);
and U2536 (N_2536,N_1593,N_2199);
xor U2537 (N_2537,N_2129,N_2015);
or U2538 (N_2538,N_1634,N_1609);
or U2539 (N_2539,N_2229,N_1988);
nand U2540 (N_2540,N_1874,N_2017);
nor U2541 (N_2541,N_2057,N_2170);
nor U2542 (N_2542,N_1688,N_2172);
xnor U2543 (N_2543,N_2018,N_1675);
nand U2544 (N_2544,N_2147,N_1745);
nor U2545 (N_2545,N_1777,N_1770);
and U2546 (N_2546,N_1850,N_1640);
or U2547 (N_2547,N_1975,N_2094);
nor U2548 (N_2548,N_1839,N_1616);
or U2549 (N_2549,N_1737,N_2187);
or U2550 (N_2550,N_1597,N_1531);
and U2551 (N_2551,N_2146,N_2069);
nand U2552 (N_2552,N_1736,N_1635);
xnor U2553 (N_2553,N_1882,N_1583);
nor U2554 (N_2554,N_2113,N_1765);
and U2555 (N_2555,N_2181,N_1983);
xor U2556 (N_2556,N_2115,N_2205);
or U2557 (N_2557,N_1847,N_1797);
or U2558 (N_2558,N_1819,N_1676);
nor U2559 (N_2559,N_2034,N_1806);
or U2560 (N_2560,N_2079,N_2002);
nand U2561 (N_2561,N_2185,N_2137);
nand U2562 (N_2562,N_1614,N_1911);
nor U2563 (N_2563,N_1920,N_2214);
nand U2564 (N_2564,N_1799,N_1588);
nor U2565 (N_2565,N_2071,N_2087);
or U2566 (N_2566,N_2049,N_1526);
or U2567 (N_2567,N_1557,N_1918);
nand U2568 (N_2568,N_1963,N_2025);
nor U2569 (N_2569,N_2052,N_2208);
nor U2570 (N_2570,N_2150,N_2056);
xor U2571 (N_2571,N_2104,N_2143);
nor U2572 (N_2572,N_2235,N_1842);
nor U2573 (N_2573,N_2107,N_2029);
xor U2574 (N_2574,N_1912,N_1769);
or U2575 (N_2575,N_1837,N_1612);
and U2576 (N_2576,N_1897,N_1661);
and U2577 (N_2577,N_2078,N_2067);
and U2578 (N_2578,N_1942,N_1991);
or U2579 (N_2579,N_1664,N_1705);
and U2580 (N_2580,N_2102,N_1891);
nand U2581 (N_2581,N_1711,N_2016);
xor U2582 (N_2582,N_1687,N_1928);
and U2583 (N_2583,N_1665,N_1959);
nor U2584 (N_2584,N_1948,N_1686);
nor U2585 (N_2585,N_1550,N_2242);
and U2586 (N_2586,N_2139,N_1878);
nand U2587 (N_2587,N_1956,N_1803);
nor U2588 (N_2588,N_1619,N_1889);
nor U2589 (N_2589,N_1582,N_1902);
nor U2590 (N_2590,N_1815,N_1949);
and U2591 (N_2591,N_1680,N_1629);
nor U2592 (N_2592,N_1682,N_2204);
nor U2593 (N_2593,N_1592,N_1590);
or U2594 (N_2594,N_1856,N_1546);
and U2595 (N_2595,N_1990,N_2118);
and U2596 (N_2596,N_1585,N_1725);
nor U2597 (N_2597,N_1924,N_1624);
or U2598 (N_2598,N_1727,N_1600);
xor U2599 (N_2599,N_1901,N_2173);
or U2600 (N_2600,N_1697,N_1914);
and U2601 (N_2601,N_1611,N_2101);
and U2602 (N_2602,N_1813,N_1810);
nand U2603 (N_2603,N_2073,N_1958);
nand U2604 (N_2604,N_1820,N_1743);
xnor U2605 (N_2605,N_2153,N_2133);
nor U2606 (N_2606,N_2145,N_2241);
or U2607 (N_2607,N_2169,N_1719);
and U2608 (N_2608,N_1568,N_1875);
and U2609 (N_2609,N_1834,N_1512);
and U2610 (N_2610,N_1821,N_1852);
nor U2611 (N_2611,N_2232,N_1666);
or U2612 (N_2612,N_2190,N_2053);
nand U2613 (N_2613,N_1596,N_2225);
nor U2614 (N_2614,N_2163,N_1708);
and U2615 (N_2615,N_2048,N_1753);
and U2616 (N_2616,N_1641,N_2042);
or U2617 (N_2617,N_2154,N_1952);
or U2618 (N_2618,N_1976,N_1969);
or U2619 (N_2619,N_1758,N_2075);
or U2620 (N_2620,N_1569,N_1505);
and U2621 (N_2621,N_1999,N_1559);
xor U2622 (N_2622,N_1571,N_1796);
xnor U2623 (N_2623,N_2043,N_2161);
nand U2624 (N_2624,N_1742,N_1929);
or U2625 (N_2625,N_1725,N_1616);
or U2626 (N_2626,N_1595,N_1574);
or U2627 (N_2627,N_2089,N_1612);
nand U2628 (N_2628,N_1856,N_1900);
or U2629 (N_2629,N_1638,N_1753);
nor U2630 (N_2630,N_1708,N_1666);
nor U2631 (N_2631,N_1774,N_1830);
or U2632 (N_2632,N_1908,N_1962);
or U2633 (N_2633,N_1650,N_1660);
nor U2634 (N_2634,N_1631,N_1798);
xor U2635 (N_2635,N_1801,N_2070);
nand U2636 (N_2636,N_1727,N_2116);
nor U2637 (N_2637,N_1581,N_1516);
or U2638 (N_2638,N_2154,N_2247);
nand U2639 (N_2639,N_2123,N_2176);
or U2640 (N_2640,N_2135,N_1944);
nor U2641 (N_2641,N_2064,N_1766);
xnor U2642 (N_2642,N_1869,N_1817);
and U2643 (N_2643,N_2175,N_1884);
xnor U2644 (N_2644,N_1738,N_1634);
and U2645 (N_2645,N_1535,N_1821);
nor U2646 (N_2646,N_2118,N_1946);
nand U2647 (N_2647,N_1942,N_1749);
and U2648 (N_2648,N_1804,N_2214);
and U2649 (N_2649,N_1653,N_1907);
xnor U2650 (N_2650,N_1896,N_1820);
or U2651 (N_2651,N_2137,N_1729);
nor U2652 (N_2652,N_1723,N_1558);
nor U2653 (N_2653,N_1945,N_1906);
and U2654 (N_2654,N_1757,N_1942);
and U2655 (N_2655,N_1698,N_2049);
nor U2656 (N_2656,N_1582,N_1707);
or U2657 (N_2657,N_2098,N_1725);
xnor U2658 (N_2658,N_1883,N_2034);
xor U2659 (N_2659,N_2085,N_1910);
or U2660 (N_2660,N_2065,N_1513);
and U2661 (N_2661,N_1593,N_1504);
nand U2662 (N_2662,N_1677,N_1856);
nor U2663 (N_2663,N_2140,N_2004);
nand U2664 (N_2664,N_2005,N_2031);
or U2665 (N_2665,N_1888,N_1731);
or U2666 (N_2666,N_1848,N_1730);
nor U2667 (N_2667,N_2087,N_1565);
nand U2668 (N_2668,N_1844,N_1765);
nor U2669 (N_2669,N_2016,N_2106);
and U2670 (N_2670,N_1951,N_1515);
xnor U2671 (N_2671,N_2121,N_1749);
nand U2672 (N_2672,N_1785,N_2175);
nand U2673 (N_2673,N_2191,N_1613);
or U2674 (N_2674,N_1906,N_1919);
nand U2675 (N_2675,N_2193,N_1959);
nand U2676 (N_2676,N_1968,N_1653);
xnor U2677 (N_2677,N_2094,N_2045);
nor U2678 (N_2678,N_1997,N_1803);
xnor U2679 (N_2679,N_1862,N_1795);
and U2680 (N_2680,N_2244,N_1940);
and U2681 (N_2681,N_1770,N_1751);
nor U2682 (N_2682,N_1606,N_1595);
nor U2683 (N_2683,N_2176,N_1859);
or U2684 (N_2684,N_1959,N_2206);
nand U2685 (N_2685,N_1747,N_1537);
or U2686 (N_2686,N_2239,N_1641);
or U2687 (N_2687,N_1835,N_2135);
and U2688 (N_2688,N_1785,N_2037);
and U2689 (N_2689,N_1957,N_1718);
and U2690 (N_2690,N_1594,N_1975);
nand U2691 (N_2691,N_2043,N_1702);
nor U2692 (N_2692,N_1558,N_2135);
nand U2693 (N_2693,N_1563,N_2235);
xnor U2694 (N_2694,N_2125,N_1626);
and U2695 (N_2695,N_2228,N_1518);
xnor U2696 (N_2696,N_1774,N_1536);
nor U2697 (N_2697,N_1656,N_1794);
or U2698 (N_2698,N_1518,N_1625);
nor U2699 (N_2699,N_2103,N_2066);
and U2700 (N_2700,N_1575,N_2201);
nand U2701 (N_2701,N_1802,N_2164);
and U2702 (N_2702,N_1610,N_1627);
or U2703 (N_2703,N_2109,N_1733);
nor U2704 (N_2704,N_2222,N_2080);
or U2705 (N_2705,N_1962,N_1865);
and U2706 (N_2706,N_2154,N_2101);
nand U2707 (N_2707,N_1880,N_2222);
xnor U2708 (N_2708,N_2237,N_1517);
and U2709 (N_2709,N_1760,N_1779);
and U2710 (N_2710,N_1870,N_1831);
or U2711 (N_2711,N_2124,N_1521);
nand U2712 (N_2712,N_1856,N_1727);
nor U2713 (N_2713,N_1810,N_2132);
or U2714 (N_2714,N_2145,N_1721);
nor U2715 (N_2715,N_2188,N_1665);
nand U2716 (N_2716,N_2136,N_1845);
nand U2717 (N_2717,N_1664,N_1516);
and U2718 (N_2718,N_1891,N_1574);
xor U2719 (N_2719,N_1623,N_2241);
and U2720 (N_2720,N_1721,N_1929);
nor U2721 (N_2721,N_2063,N_1678);
or U2722 (N_2722,N_2048,N_1684);
nand U2723 (N_2723,N_1604,N_2198);
xnor U2724 (N_2724,N_1677,N_2042);
and U2725 (N_2725,N_2137,N_1920);
nor U2726 (N_2726,N_1512,N_2095);
nor U2727 (N_2727,N_1786,N_1762);
or U2728 (N_2728,N_1857,N_1626);
xor U2729 (N_2729,N_2007,N_2140);
or U2730 (N_2730,N_2038,N_1514);
nor U2731 (N_2731,N_1786,N_1711);
or U2732 (N_2732,N_1955,N_2237);
nor U2733 (N_2733,N_2150,N_1993);
xor U2734 (N_2734,N_1899,N_2088);
or U2735 (N_2735,N_2225,N_1844);
and U2736 (N_2736,N_1829,N_2047);
nor U2737 (N_2737,N_1659,N_1538);
nand U2738 (N_2738,N_1544,N_1609);
xor U2739 (N_2739,N_1670,N_1957);
and U2740 (N_2740,N_2070,N_1751);
xnor U2741 (N_2741,N_1676,N_1552);
nand U2742 (N_2742,N_1805,N_1600);
or U2743 (N_2743,N_1897,N_1949);
nor U2744 (N_2744,N_1809,N_2005);
nand U2745 (N_2745,N_1985,N_2095);
or U2746 (N_2746,N_2041,N_2176);
nor U2747 (N_2747,N_1970,N_1708);
nor U2748 (N_2748,N_1584,N_2162);
and U2749 (N_2749,N_1603,N_1664);
nor U2750 (N_2750,N_1652,N_2206);
xor U2751 (N_2751,N_2206,N_1574);
nor U2752 (N_2752,N_2015,N_2104);
nor U2753 (N_2753,N_1872,N_1914);
nor U2754 (N_2754,N_1515,N_1921);
nor U2755 (N_2755,N_2092,N_2054);
or U2756 (N_2756,N_2174,N_1596);
or U2757 (N_2757,N_2019,N_1544);
or U2758 (N_2758,N_2112,N_2146);
nand U2759 (N_2759,N_2214,N_2091);
nor U2760 (N_2760,N_2105,N_1800);
nor U2761 (N_2761,N_1983,N_1568);
xor U2762 (N_2762,N_1866,N_1762);
and U2763 (N_2763,N_1657,N_1537);
nand U2764 (N_2764,N_2143,N_2049);
nand U2765 (N_2765,N_1930,N_1505);
and U2766 (N_2766,N_1799,N_2219);
and U2767 (N_2767,N_1825,N_1631);
or U2768 (N_2768,N_2041,N_2154);
xnor U2769 (N_2769,N_1699,N_1971);
or U2770 (N_2770,N_2170,N_1558);
nand U2771 (N_2771,N_1516,N_1584);
xor U2772 (N_2772,N_2209,N_2177);
and U2773 (N_2773,N_2240,N_1793);
or U2774 (N_2774,N_2228,N_2185);
nand U2775 (N_2775,N_1698,N_2154);
xor U2776 (N_2776,N_1928,N_1616);
nor U2777 (N_2777,N_1849,N_2176);
nor U2778 (N_2778,N_2201,N_2080);
xor U2779 (N_2779,N_1869,N_1675);
and U2780 (N_2780,N_2099,N_1908);
nor U2781 (N_2781,N_2156,N_1921);
or U2782 (N_2782,N_1716,N_2160);
xnor U2783 (N_2783,N_2094,N_1647);
or U2784 (N_2784,N_1815,N_2000);
nor U2785 (N_2785,N_2065,N_2064);
nor U2786 (N_2786,N_2144,N_1920);
nor U2787 (N_2787,N_1601,N_1755);
or U2788 (N_2788,N_1684,N_2091);
or U2789 (N_2789,N_1657,N_2188);
and U2790 (N_2790,N_1659,N_1542);
nand U2791 (N_2791,N_1854,N_1859);
nor U2792 (N_2792,N_1598,N_1901);
nor U2793 (N_2793,N_1509,N_1897);
and U2794 (N_2794,N_2009,N_1912);
or U2795 (N_2795,N_1712,N_1866);
nor U2796 (N_2796,N_1584,N_2200);
nor U2797 (N_2797,N_2040,N_2202);
nor U2798 (N_2798,N_1638,N_1919);
and U2799 (N_2799,N_2198,N_1761);
or U2800 (N_2800,N_1687,N_2047);
nor U2801 (N_2801,N_1996,N_1561);
nand U2802 (N_2802,N_1893,N_2022);
or U2803 (N_2803,N_2002,N_1885);
and U2804 (N_2804,N_2011,N_1575);
and U2805 (N_2805,N_1942,N_2238);
or U2806 (N_2806,N_2225,N_1894);
nor U2807 (N_2807,N_1929,N_2202);
xnor U2808 (N_2808,N_2210,N_1567);
and U2809 (N_2809,N_1825,N_1848);
nor U2810 (N_2810,N_2000,N_2056);
or U2811 (N_2811,N_2036,N_1666);
nand U2812 (N_2812,N_2148,N_1716);
or U2813 (N_2813,N_1912,N_1674);
xor U2814 (N_2814,N_1861,N_2154);
or U2815 (N_2815,N_2197,N_2143);
or U2816 (N_2816,N_1528,N_1894);
nor U2817 (N_2817,N_2217,N_2245);
and U2818 (N_2818,N_1621,N_2142);
nor U2819 (N_2819,N_1819,N_2052);
or U2820 (N_2820,N_2101,N_1522);
or U2821 (N_2821,N_2163,N_1657);
nand U2822 (N_2822,N_1786,N_1668);
xor U2823 (N_2823,N_1741,N_2102);
xor U2824 (N_2824,N_1576,N_1661);
and U2825 (N_2825,N_1504,N_1913);
xor U2826 (N_2826,N_2086,N_1664);
nand U2827 (N_2827,N_2128,N_1563);
or U2828 (N_2828,N_1990,N_2012);
nand U2829 (N_2829,N_1667,N_2141);
nand U2830 (N_2830,N_1953,N_2205);
nand U2831 (N_2831,N_2126,N_1850);
nand U2832 (N_2832,N_1727,N_1987);
and U2833 (N_2833,N_2198,N_1602);
nand U2834 (N_2834,N_2230,N_2202);
or U2835 (N_2835,N_1907,N_1873);
xnor U2836 (N_2836,N_2181,N_1616);
xnor U2837 (N_2837,N_2000,N_1669);
nor U2838 (N_2838,N_2020,N_2201);
nand U2839 (N_2839,N_2121,N_1776);
or U2840 (N_2840,N_1554,N_1704);
nand U2841 (N_2841,N_1622,N_1565);
nor U2842 (N_2842,N_1549,N_1969);
and U2843 (N_2843,N_1892,N_2219);
or U2844 (N_2844,N_1762,N_1957);
xnor U2845 (N_2845,N_1594,N_1637);
nor U2846 (N_2846,N_1898,N_2244);
nor U2847 (N_2847,N_1832,N_1607);
and U2848 (N_2848,N_1563,N_1625);
xnor U2849 (N_2849,N_2130,N_2143);
or U2850 (N_2850,N_2101,N_1887);
xor U2851 (N_2851,N_1709,N_2212);
nand U2852 (N_2852,N_1694,N_1859);
nand U2853 (N_2853,N_1933,N_1924);
and U2854 (N_2854,N_1984,N_2242);
xor U2855 (N_2855,N_2141,N_2023);
and U2856 (N_2856,N_1995,N_1563);
xor U2857 (N_2857,N_2093,N_1800);
nand U2858 (N_2858,N_1885,N_2113);
nand U2859 (N_2859,N_2091,N_2152);
or U2860 (N_2860,N_1807,N_2003);
nand U2861 (N_2861,N_1844,N_2046);
xor U2862 (N_2862,N_2223,N_2038);
and U2863 (N_2863,N_1648,N_1666);
nor U2864 (N_2864,N_1595,N_1550);
nor U2865 (N_2865,N_1852,N_1624);
xor U2866 (N_2866,N_1631,N_2152);
and U2867 (N_2867,N_1967,N_1995);
nand U2868 (N_2868,N_1931,N_1902);
and U2869 (N_2869,N_1540,N_2151);
nand U2870 (N_2870,N_1780,N_2044);
and U2871 (N_2871,N_1847,N_1859);
nor U2872 (N_2872,N_2139,N_2109);
and U2873 (N_2873,N_1654,N_1879);
or U2874 (N_2874,N_1591,N_2103);
nor U2875 (N_2875,N_2205,N_1713);
nor U2876 (N_2876,N_1913,N_1630);
or U2877 (N_2877,N_1652,N_1892);
nand U2878 (N_2878,N_1838,N_1976);
nand U2879 (N_2879,N_1589,N_1987);
nor U2880 (N_2880,N_1666,N_1597);
and U2881 (N_2881,N_1759,N_2087);
nand U2882 (N_2882,N_1821,N_1866);
and U2883 (N_2883,N_2024,N_1991);
nor U2884 (N_2884,N_1625,N_2191);
nand U2885 (N_2885,N_2137,N_1855);
and U2886 (N_2886,N_2161,N_2174);
nand U2887 (N_2887,N_1918,N_1927);
xnor U2888 (N_2888,N_1829,N_1544);
nand U2889 (N_2889,N_1973,N_1554);
nand U2890 (N_2890,N_1664,N_1992);
nor U2891 (N_2891,N_1916,N_2202);
nor U2892 (N_2892,N_2154,N_1743);
and U2893 (N_2893,N_1979,N_2161);
xor U2894 (N_2894,N_2137,N_2167);
xnor U2895 (N_2895,N_1564,N_1548);
nand U2896 (N_2896,N_2180,N_1735);
xnor U2897 (N_2897,N_2212,N_2065);
xor U2898 (N_2898,N_1912,N_1668);
and U2899 (N_2899,N_2117,N_2005);
and U2900 (N_2900,N_1876,N_2103);
and U2901 (N_2901,N_1970,N_2164);
xor U2902 (N_2902,N_1913,N_2155);
xor U2903 (N_2903,N_2185,N_1937);
nor U2904 (N_2904,N_2020,N_1573);
or U2905 (N_2905,N_2055,N_1738);
and U2906 (N_2906,N_1799,N_1625);
nor U2907 (N_2907,N_1571,N_2066);
and U2908 (N_2908,N_1910,N_1792);
or U2909 (N_2909,N_1902,N_1719);
nand U2910 (N_2910,N_1887,N_2102);
or U2911 (N_2911,N_1558,N_2140);
xor U2912 (N_2912,N_1914,N_2215);
nand U2913 (N_2913,N_2179,N_1978);
nand U2914 (N_2914,N_2076,N_1669);
and U2915 (N_2915,N_1517,N_1978);
xnor U2916 (N_2916,N_1994,N_2212);
and U2917 (N_2917,N_1607,N_1904);
nor U2918 (N_2918,N_1665,N_1919);
or U2919 (N_2919,N_1620,N_1849);
nand U2920 (N_2920,N_2059,N_1904);
nor U2921 (N_2921,N_2121,N_1649);
and U2922 (N_2922,N_1856,N_1924);
nand U2923 (N_2923,N_2244,N_1598);
xor U2924 (N_2924,N_1684,N_1909);
or U2925 (N_2925,N_1648,N_2015);
xor U2926 (N_2926,N_2177,N_1643);
or U2927 (N_2927,N_1890,N_1805);
xnor U2928 (N_2928,N_2139,N_1658);
nor U2929 (N_2929,N_1569,N_2031);
nor U2930 (N_2930,N_1606,N_1960);
nor U2931 (N_2931,N_1581,N_1764);
or U2932 (N_2932,N_1727,N_1973);
or U2933 (N_2933,N_2055,N_2117);
or U2934 (N_2934,N_2189,N_2136);
or U2935 (N_2935,N_1599,N_1556);
nand U2936 (N_2936,N_2091,N_1836);
nand U2937 (N_2937,N_1741,N_1865);
nor U2938 (N_2938,N_1731,N_2177);
xnor U2939 (N_2939,N_1624,N_1799);
nand U2940 (N_2940,N_1865,N_1511);
and U2941 (N_2941,N_1895,N_1822);
xnor U2942 (N_2942,N_1900,N_2115);
nand U2943 (N_2943,N_1770,N_2209);
nand U2944 (N_2944,N_2184,N_2048);
xor U2945 (N_2945,N_1844,N_2239);
nand U2946 (N_2946,N_1911,N_1974);
xor U2947 (N_2947,N_2118,N_1819);
xnor U2948 (N_2948,N_1564,N_2013);
or U2949 (N_2949,N_1518,N_2014);
nand U2950 (N_2950,N_1699,N_2062);
nor U2951 (N_2951,N_1619,N_1738);
nor U2952 (N_2952,N_1541,N_1925);
nand U2953 (N_2953,N_1833,N_2166);
and U2954 (N_2954,N_1528,N_1724);
nor U2955 (N_2955,N_2136,N_2139);
and U2956 (N_2956,N_1841,N_2130);
xor U2957 (N_2957,N_1520,N_2186);
nand U2958 (N_2958,N_2236,N_1658);
nor U2959 (N_2959,N_1643,N_2119);
nor U2960 (N_2960,N_1536,N_1552);
nor U2961 (N_2961,N_2047,N_2142);
nor U2962 (N_2962,N_1503,N_1617);
and U2963 (N_2963,N_2213,N_1663);
xnor U2964 (N_2964,N_1992,N_2143);
and U2965 (N_2965,N_2020,N_1521);
and U2966 (N_2966,N_2033,N_1845);
and U2967 (N_2967,N_1908,N_1652);
or U2968 (N_2968,N_1704,N_1845);
nand U2969 (N_2969,N_2107,N_1889);
and U2970 (N_2970,N_2006,N_1861);
nor U2971 (N_2971,N_2048,N_1559);
or U2972 (N_2972,N_2121,N_2131);
xnor U2973 (N_2973,N_1850,N_1839);
nand U2974 (N_2974,N_2190,N_1842);
nor U2975 (N_2975,N_2183,N_1758);
nand U2976 (N_2976,N_1581,N_2054);
xnor U2977 (N_2977,N_2016,N_2145);
nor U2978 (N_2978,N_2246,N_2041);
nand U2979 (N_2979,N_1806,N_1525);
or U2980 (N_2980,N_2207,N_1897);
nor U2981 (N_2981,N_2116,N_1897);
or U2982 (N_2982,N_1959,N_1607);
xnor U2983 (N_2983,N_2185,N_1680);
xnor U2984 (N_2984,N_2123,N_1881);
or U2985 (N_2985,N_1959,N_1920);
xor U2986 (N_2986,N_2119,N_1611);
xor U2987 (N_2987,N_1613,N_1590);
nand U2988 (N_2988,N_1937,N_2007);
or U2989 (N_2989,N_1663,N_2140);
xor U2990 (N_2990,N_2087,N_1669);
and U2991 (N_2991,N_1792,N_1855);
nor U2992 (N_2992,N_1909,N_2172);
or U2993 (N_2993,N_1581,N_2209);
nor U2994 (N_2994,N_2140,N_1505);
nand U2995 (N_2995,N_1519,N_2019);
xnor U2996 (N_2996,N_1776,N_2242);
xor U2997 (N_2997,N_1610,N_1661);
nand U2998 (N_2998,N_2045,N_2113);
or U2999 (N_2999,N_1551,N_2130);
xnor U3000 (N_3000,N_2597,N_2280);
xor U3001 (N_3001,N_2293,N_2617);
xnor U3002 (N_3002,N_2957,N_2499);
and U3003 (N_3003,N_2685,N_2865);
nor U3004 (N_3004,N_2360,N_2821);
nand U3005 (N_3005,N_2502,N_2457);
or U3006 (N_3006,N_2784,N_2652);
xnor U3007 (N_3007,N_2377,N_2730);
nor U3008 (N_3008,N_2675,N_2447);
nand U3009 (N_3009,N_2943,N_2708);
nand U3010 (N_3010,N_2759,N_2992);
xor U3011 (N_3011,N_2544,N_2479);
or U3012 (N_3012,N_2789,N_2659);
nor U3013 (N_3013,N_2747,N_2611);
nand U3014 (N_3014,N_2576,N_2982);
xor U3015 (N_3015,N_2868,N_2738);
nor U3016 (N_3016,N_2438,N_2507);
and U3017 (N_3017,N_2612,N_2583);
nand U3018 (N_3018,N_2965,N_2669);
xnor U3019 (N_3019,N_2713,N_2250);
and U3020 (N_3020,N_2797,N_2551);
and U3021 (N_3021,N_2431,N_2344);
xnor U3022 (N_3022,N_2814,N_2372);
nand U3023 (N_3023,N_2754,N_2656);
nand U3024 (N_3024,N_2812,N_2462);
nor U3025 (N_3025,N_2774,N_2436);
xor U3026 (N_3026,N_2296,N_2416);
nor U3027 (N_3027,N_2822,N_2853);
nand U3028 (N_3028,N_2843,N_2324);
xor U3029 (N_3029,N_2839,N_2834);
xnor U3030 (N_3030,N_2629,N_2934);
nor U3031 (N_3031,N_2779,N_2847);
and U3032 (N_3032,N_2326,N_2719);
xnor U3033 (N_3033,N_2320,N_2680);
and U3034 (N_3034,N_2552,N_2863);
and U3035 (N_3035,N_2610,N_2516);
and U3036 (N_3036,N_2419,N_2321);
nand U3037 (N_3037,N_2563,N_2949);
nand U3038 (N_3038,N_2527,N_2302);
nor U3039 (N_3039,N_2857,N_2481);
nand U3040 (N_3040,N_2557,N_2442);
xnor U3041 (N_3041,N_2748,N_2978);
nand U3042 (N_3042,N_2867,N_2701);
or U3043 (N_3043,N_2791,N_2271);
xnor U3044 (N_3044,N_2806,N_2422);
and U3045 (N_3045,N_2603,N_2418);
and U3046 (N_3046,N_2590,N_2497);
and U3047 (N_3047,N_2255,N_2412);
nor U3048 (N_3048,N_2714,N_2971);
and U3049 (N_3049,N_2578,N_2564);
xnor U3050 (N_3050,N_2461,N_2953);
nor U3051 (N_3051,N_2985,N_2517);
nor U3052 (N_3052,N_2846,N_2329);
nor U3053 (N_3053,N_2725,N_2705);
nand U3054 (N_3054,N_2633,N_2687);
xnor U3055 (N_3055,N_2694,N_2401);
nand U3056 (N_3056,N_2709,N_2284);
nand U3057 (N_3057,N_2281,N_2459);
nand U3058 (N_3058,N_2671,N_2876);
xnor U3059 (N_3059,N_2448,N_2991);
nor U3060 (N_3060,N_2399,N_2395);
nor U3061 (N_3061,N_2404,N_2451);
nand U3062 (N_3062,N_2877,N_2547);
and U3063 (N_3063,N_2803,N_2618);
xnor U3064 (N_3064,N_2625,N_2627);
xor U3065 (N_3065,N_2327,N_2945);
nand U3066 (N_3066,N_2323,N_2270);
nand U3067 (N_3067,N_2464,N_2542);
and U3068 (N_3068,N_2826,N_2443);
or U3069 (N_3069,N_2406,N_2873);
nor U3070 (N_3070,N_2930,N_2283);
nand U3071 (N_3071,N_2541,N_2682);
nor U3072 (N_3072,N_2550,N_2415);
or U3073 (N_3073,N_2587,N_2653);
nor U3074 (N_3074,N_2702,N_2661);
nand U3075 (N_3075,N_2763,N_2765);
nor U3076 (N_3076,N_2289,N_2456);
nor U3077 (N_3077,N_2900,N_2494);
and U3078 (N_3078,N_2662,N_2695);
nor U3079 (N_3079,N_2535,N_2735);
xor U3080 (N_3080,N_2282,N_2279);
or U3081 (N_3081,N_2974,N_2512);
and U3082 (N_3082,N_2330,N_2673);
nand U3083 (N_3083,N_2514,N_2488);
xor U3084 (N_3084,N_2760,N_2647);
nand U3085 (N_3085,N_2631,N_2836);
xnor U3086 (N_3086,N_2729,N_2704);
or U3087 (N_3087,N_2390,N_2916);
xor U3088 (N_3088,N_2349,N_2785);
nor U3089 (N_3089,N_2919,N_2973);
nor U3090 (N_3090,N_2491,N_2304);
or U3091 (N_3091,N_2484,N_2305);
nor U3092 (N_3092,N_2534,N_2265);
nand U3093 (N_3093,N_2430,N_2411);
nor U3094 (N_3094,N_2638,N_2813);
and U3095 (N_3095,N_2883,N_2427);
or U3096 (N_3096,N_2635,N_2392);
or U3097 (N_3097,N_2988,N_2744);
nand U3098 (N_3098,N_2439,N_2260);
nand U3099 (N_3099,N_2585,N_2852);
and U3100 (N_3100,N_2726,N_2545);
xnor U3101 (N_3101,N_2844,N_2616);
or U3102 (N_3102,N_2913,N_2463);
nand U3103 (N_3103,N_2696,N_2712);
nand U3104 (N_3104,N_2906,N_2799);
nor U3105 (N_3105,N_2926,N_2875);
and U3106 (N_3106,N_2707,N_2605);
or U3107 (N_3107,N_2340,N_2634);
xor U3108 (N_3108,N_2668,N_2571);
or U3109 (N_3109,N_2972,N_2642);
nand U3110 (N_3110,N_2566,N_2804);
or U3111 (N_3111,N_2994,N_2352);
nand U3112 (N_3112,N_2689,N_2721);
xor U3113 (N_3113,N_2278,N_2966);
nand U3114 (N_3114,N_2872,N_2549);
xnor U3115 (N_3115,N_2833,N_2562);
and U3116 (N_3116,N_2465,N_2924);
nand U3117 (N_3117,N_2783,N_2946);
xor U3118 (N_3118,N_2325,N_2999);
or U3119 (N_3119,N_2776,N_2292);
and U3120 (N_3120,N_2891,N_2503);
nand U3121 (N_3121,N_2397,N_2986);
xor U3122 (N_3122,N_2902,N_2267);
nand U3123 (N_3123,N_2414,N_2905);
or U3124 (N_3124,N_2838,N_2435);
or U3125 (N_3125,N_2529,N_2665);
and U3126 (N_3126,N_2276,N_2408);
nand U3127 (N_3127,N_2644,N_2802);
nand U3128 (N_3128,N_2317,N_2958);
or U3129 (N_3129,N_2718,N_2383);
nor U3130 (N_3130,N_2753,N_2300);
or U3131 (N_3131,N_2683,N_2948);
xnor U3132 (N_3132,N_2252,N_2840);
and U3133 (N_3133,N_2519,N_2533);
and U3134 (N_3134,N_2498,N_2658);
or U3135 (N_3135,N_2579,N_2601);
and U3136 (N_3136,N_2609,N_2472);
nor U3137 (N_3137,N_2703,N_2425);
nand U3138 (N_3138,N_2523,N_2676);
nor U3139 (N_3139,N_2710,N_2391);
nand U3140 (N_3140,N_2429,N_2667);
nor U3141 (N_3141,N_2510,N_2921);
xnor U3142 (N_3142,N_2331,N_2871);
or U3143 (N_3143,N_2742,N_2258);
or U3144 (N_3144,N_2896,N_2449);
or U3145 (N_3145,N_2453,N_2739);
xor U3146 (N_3146,N_2341,N_2750);
nand U3147 (N_3147,N_2801,N_2405);
nor U3148 (N_3148,N_2829,N_2678);
or U3149 (N_3149,N_2370,N_2486);
nand U3150 (N_3150,N_2663,N_2778);
nand U3151 (N_3151,N_2630,N_2940);
xnor U3152 (N_3152,N_2699,N_2935);
or U3153 (N_3153,N_2733,N_2385);
and U3154 (N_3154,N_2367,N_2434);
nand U3155 (N_3155,N_2795,N_2310);
and U3156 (N_3156,N_2645,N_2688);
xor U3157 (N_3157,N_2890,N_2577);
xnor U3158 (N_3158,N_2619,N_2927);
and U3159 (N_3159,N_2558,N_2780);
nand U3160 (N_3160,N_2698,N_2664);
xnor U3161 (N_3161,N_2599,N_2918);
xnor U3162 (N_3162,N_2745,N_2396);
and U3163 (N_3163,N_2850,N_2870);
nand U3164 (N_3164,N_2674,N_2777);
and U3165 (N_3165,N_2602,N_2861);
and U3166 (N_3166,N_2641,N_2526);
and U3167 (N_3167,N_2473,N_2963);
nand U3168 (N_3168,N_2720,N_2758);
nor U3169 (N_3169,N_2468,N_2369);
xor U3170 (N_3170,N_2475,N_2591);
nand U3171 (N_3171,N_2257,N_2649);
and U3172 (N_3172,N_2732,N_2622);
or U3173 (N_3173,N_2474,N_2528);
xnor U3174 (N_3174,N_2345,N_2909);
xor U3175 (N_3175,N_2715,N_2899);
xnor U3176 (N_3176,N_2773,N_2318);
and U3177 (N_3177,N_2772,N_2818);
or U3178 (N_3178,N_2987,N_2990);
or U3179 (N_3179,N_2901,N_2467);
nor U3180 (N_3180,N_2820,N_2660);
and U3181 (N_3181,N_2864,N_2606);
and U3182 (N_3182,N_2537,N_2693);
nand U3183 (N_3183,N_2679,N_2637);
nand U3184 (N_3184,N_2460,N_2740);
or U3185 (N_3185,N_2384,N_2621);
nor U3186 (N_3186,N_2856,N_2493);
nor U3187 (N_3187,N_2827,N_2962);
or U3188 (N_3188,N_2954,N_2588);
and U3189 (N_3189,N_2362,N_2614);
nand U3190 (N_3190,N_2446,N_2771);
and U3191 (N_3191,N_2273,N_2291);
and U3192 (N_3192,N_2737,N_2312);
nand U3193 (N_3193,N_2269,N_2375);
or U3194 (N_3194,N_2513,N_2817);
xnor U3195 (N_3195,N_2775,N_2423);
xor U3196 (N_3196,N_2980,N_2309);
nor U3197 (N_3197,N_2595,N_2368);
or U3198 (N_3198,N_2727,N_2811);
nor U3199 (N_3199,N_2388,N_2356);
xor U3200 (N_3200,N_2573,N_2762);
xor U3201 (N_3201,N_2452,N_2261);
and U3202 (N_3202,N_2787,N_2454);
xor U3203 (N_3203,N_2338,N_2931);
nand U3204 (N_3204,N_2301,N_2722);
xnor U3205 (N_3205,N_2997,N_2858);
nor U3206 (N_3206,N_2706,N_2286);
xor U3207 (N_3207,N_2343,N_2879);
and U3208 (N_3208,N_2543,N_2288);
or U3209 (N_3209,N_2572,N_2692);
or U3210 (N_3210,N_2888,N_2350);
and U3211 (N_3211,N_2848,N_2313);
and U3212 (N_3212,N_2677,N_2593);
nand U3213 (N_3213,N_2908,N_2274);
nand U3214 (N_3214,N_2734,N_2939);
xnor U3215 (N_3215,N_2755,N_2624);
and U3216 (N_3216,N_2615,N_2333);
or U3217 (N_3217,N_2342,N_2420);
xnor U3218 (N_3218,N_2793,N_2574);
nand U3219 (N_3219,N_2794,N_2968);
xor U3220 (N_3220,N_2831,N_2371);
xnor U3221 (N_3221,N_2914,N_2928);
xnor U3222 (N_3222,N_2751,N_2790);
or U3223 (N_3223,N_2700,N_2810);
and U3224 (N_3224,N_2582,N_2509);
or U3225 (N_3225,N_2893,N_2376);
or U3226 (N_3226,N_2936,N_2741);
nor U3227 (N_3227,N_2950,N_2929);
nor U3228 (N_3228,N_2849,N_2508);
or U3229 (N_3229,N_2800,N_2361);
nor U3230 (N_3230,N_2964,N_2386);
nand U3231 (N_3231,N_2316,N_2770);
or U3232 (N_3232,N_2311,N_2654);
and U3233 (N_3233,N_2967,N_2522);
nand U3234 (N_3234,N_2830,N_2640);
or U3235 (N_3235,N_2485,N_2568);
or U3236 (N_3236,N_2989,N_2977);
xor U3237 (N_3237,N_2394,N_2903);
nand U3238 (N_3238,N_2277,N_2560);
nor U3239 (N_3239,N_2596,N_2555);
and U3240 (N_3240,N_2942,N_2933);
nor U3241 (N_3241,N_2860,N_2716);
nand U3242 (N_3242,N_2743,N_2952);
nor U3243 (N_3243,N_2938,N_2378);
or U3244 (N_3244,N_2441,N_2445);
or U3245 (N_3245,N_2684,N_2536);
nand U3246 (N_3246,N_2357,N_2353);
or U3247 (N_3247,N_2569,N_2314);
xnor U3248 (N_3248,N_2275,N_2489);
or U3249 (N_3249,N_2969,N_2816);
or U3250 (N_3250,N_2521,N_2254);
nand U3251 (N_3251,N_2648,N_2897);
xnor U3252 (N_3252,N_2922,N_2354);
xor U3253 (N_3253,N_2912,N_2651);
nor U3254 (N_3254,N_2837,N_2981);
and U3255 (N_3255,N_2374,N_2251);
nor U3256 (N_3256,N_2808,N_2728);
or U3257 (N_3257,N_2670,N_2904);
and U3258 (N_3258,N_2364,N_2724);
nand U3259 (N_3259,N_2917,N_2885);
nor U3260 (N_3260,N_2532,N_2490);
or U3261 (N_3261,N_2381,N_2944);
or U3262 (N_3262,N_2554,N_2690);
and U3263 (N_3263,N_2298,N_2306);
nand U3264 (N_3264,N_2862,N_2432);
and U3265 (N_3265,N_2586,N_2539);
and U3266 (N_3266,N_2339,N_2410);
xnor U3267 (N_3267,N_2466,N_2570);
or U3268 (N_3268,N_2347,N_2524);
nor U3269 (N_3269,N_2655,N_2575);
nand U3270 (N_3270,N_2409,N_2697);
nor U3271 (N_3271,N_2805,N_2880);
xnor U3272 (N_3272,N_2650,N_2455);
nand U3273 (N_3273,N_2553,N_2268);
or U3274 (N_3274,N_2482,N_2348);
nor U3275 (N_3275,N_2556,N_2351);
nand U3276 (N_3276,N_2959,N_2628);
nor U3277 (N_3277,N_2538,N_2984);
xor U3278 (N_3278,N_2500,N_2319);
and U3279 (N_3279,N_2444,N_2626);
nor U3280 (N_3280,N_2851,N_2620);
nor U3281 (N_3281,N_2290,N_2253);
xnor U3282 (N_3282,N_2495,N_2623);
and U3283 (N_3283,N_2835,N_2925);
nand U3284 (N_3284,N_2480,N_2681);
and U3285 (N_3285,N_2841,N_2540);
nand U3286 (N_3286,N_2413,N_2608);
xnor U3287 (N_3287,N_2764,N_2607);
nand U3288 (N_3288,N_2882,N_2767);
xnor U3289 (N_3289,N_2308,N_2471);
nor U3290 (N_3290,N_2294,N_2437);
and U3291 (N_3291,N_2285,N_2749);
and U3292 (N_3292,N_2505,N_2960);
xnor U3293 (N_3293,N_2366,N_2786);
and U3294 (N_3294,N_2511,N_2768);
nand U3295 (N_3295,N_2355,N_2332);
or U3296 (N_3296,N_2970,N_2956);
or U3297 (N_3297,N_2382,N_2363);
nand U3298 (N_3298,N_2266,N_2315);
xnor U3299 (N_3299,N_2809,N_2417);
nor U3300 (N_3300,N_2983,N_2428);
or U3301 (N_3301,N_2389,N_2646);
or U3302 (N_3302,N_2478,N_2711);
or U3303 (N_3303,N_2565,N_2335);
nand U3304 (N_3304,N_2525,N_2889);
or U3305 (N_3305,N_2979,N_2782);
or U3306 (N_3306,N_2769,N_2824);
nor U3307 (N_3307,N_2477,N_2504);
and U3308 (N_3308,N_2643,N_2842);
or U3309 (N_3309,N_2400,N_2387);
or U3310 (N_3310,N_2613,N_2272);
xor U3311 (N_3311,N_2878,N_2600);
nor U3312 (N_3312,N_2845,N_2798);
nand U3313 (N_3313,N_2723,N_2975);
or U3314 (N_3314,N_2881,N_2998);
or U3315 (N_3315,N_2520,N_2380);
nand U3316 (N_3316,N_2402,N_2295);
xnor U3317 (N_3317,N_2910,N_2736);
nor U3318 (N_3318,N_2259,N_2336);
nor U3319 (N_3319,N_2756,N_2393);
nand U3320 (N_3320,N_2632,N_2825);
and U3321 (N_3321,N_2746,N_2307);
nand U3322 (N_3322,N_2886,N_2923);
nand U3323 (N_3323,N_2483,N_2515);
or U3324 (N_3324,N_2492,N_2450);
nor U3325 (N_3325,N_2823,N_2757);
or U3326 (N_3326,N_2731,N_2407);
and U3327 (N_3327,N_2932,N_2894);
xnor U3328 (N_3328,N_2854,N_2421);
or U3329 (N_3329,N_2995,N_2639);
xor U3330 (N_3330,N_2961,N_2328);
nor U3331 (N_3331,N_2501,N_2828);
xnor U3332 (N_3332,N_2955,N_2506);
nand U3333 (N_3333,N_2337,N_2469);
nand U3334 (N_3334,N_2996,N_2262);
nor U3335 (N_3335,N_2766,N_2567);
nand U3336 (N_3336,N_2832,N_2548);
xnor U3337 (N_3337,N_2531,N_2373);
or U3338 (N_3338,N_2717,N_2476);
or U3339 (N_3339,N_2781,N_2604);
or U3340 (N_3340,N_2594,N_2287);
xnor U3341 (N_3341,N_2859,N_2359);
nor U3342 (N_3342,N_2433,N_2299);
and U3343 (N_3343,N_2379,N_2691);
and U3344 (N_3344,N_2666,N_2297);
and U3345 (N_3345,N_2892,N_2686);
xor U3346 (N_3346,N_2365,N_2581);
nand U3347 (N_3347,N_2530,N_2884);
nand U3348 (N_3348,N_2941,N_2788);
nor U3349 (N_3349,N_2874,N_2657);
and U3350 (N_3350,N_2807,N_2752);
and U3351 (N_3351,N_2993,N_2915);
nand U3352 (N_3352,N_2580,N_2264);
nand U3353 (N_3353,N_2920,N_2907);
xor U3354 (N_3354,N_2796,N_2869);
xnor U3355 (N_3355,N_2303,N_2815);
or U3356 (N_3356,N_2866,N_2398);
and U3357 (N_3357,N_2334,N_2672);
nand U3358 (N_3358,N_2559,N_2598);
nor U3359 (N_3359,N_2496,N_2761);
xnor U3360 (N_3360,N_2792,N_2951);
xor U3361 (N_3361,N_2518,N_2911);
nor U3362 (N_3362,N_2887,N_2470);
and U3363 (N_3363,N_2426,N_2584);
nand U3364 (N_3364,N_2487,N_2976);
nor U3365 (N_3365,N_2898,N_2263);
xnor U3366 (N_3366,N_2546,N_2256);
nor U3367 (N_3367,N_2895,N_2346);
and U3368 (N_3368,N_2592,N_2424);
nor U3369 (N_3369,N_2458,N_2855);
nand U3370 (N_3370,N_2937,N_2403);
or U3371 (N_3371,N_2947,N_2358);
or U3372 (N_3372,N_2636,N_2440);
nand U3373 (N_3373,N_2322,N_2589);
xnor U3374 (N_3374,N_2819,N_2561);
xor U3375 (N_3375,N_2773,N_2482);
xor U3376 (N_3376,N_2993,N_2263);
nor U3377 (N_3377,N_2315,N_2407);
nor U3378 (N_3378,N_2751,N_2908);
xnor U3379 (N_3379,N_2407,N_2539);
and U3380 (N_3380,N_2405,N_2275);
xnor U3381 (N_3381,N_2289,N_2437);
nor U3382 (N_3382,N_2766,N_2619);
or U3383 (N_3383,N_2492,N_2549);
and U3384 (N_3384,N_2358,N_2483);
or U3385 (N_3385,N_2770,N_2799);
and U3386 (N_3386,N_2783,N_2830);
nand U3387 (N_3387,N_2312,N_2308);
xnor U3388 (N_3388,N_2302,N_2287);
nor U3389 (N_3389,N_2467,N_2884);
or U3390 (N_3390,N_2935,N_2552);
nand U3391 (N_3391,N_2757,N_2510);
or U3392 (N_3392,N_2400,N_2307);
and U3393 (N_3393,N_2815,N_2494);
or U3394 (N_3394,N_2967,N_2546);
xor U3395 (N_3395,N_2548,N_2819);
nand U3396 (N_3396,N_2388,N_2535);
xnor U3397 (N_3397,N_2504,N_2319);
and U3398 (N_3398,N_2252,N_2656);
or U3399 (N_3399,N_2932,N_2669);
or U3400 (N_3400,N_2251,N_2628);
nand U3401 (N_3401,N_2451,N_2601);
xnor U3402 (N_3402,N_2909,N_2762);
nor U3403 (N_3403,N_2561,N_2865);
xor U3404 (N_3404,N_2574,N_2875);
nor U3405 (N_3405,N_2261,N_2945);
nor U3406 (N_3406,N_2581,N_2364);
and U3407 (N_3407,N_2566,N_2581);
xor U3408 (N_3408,N_2647,N_2732);
xor U3409 (N_3409,N_2991,N_2723);
and U3410 (N_3410,N_2766,N_2432);
xnor U3411 (N_3411,N_2968,N_2917);
or U3412 (N_3412,N_2908,N_2838);
or U3413 (N_3413,N_2367,N_2363);
nor U3414 (N_3414,N_2257,N_2878);
and U3415 (N_3415,N_2591,N_2267);
and U3416 (N_3416,N_2403,N_2592);
or U3417 (N_3417,N_2492,N_2856);
nor U3418 (N_3418,N_2290,N_2630);
nand U3419 (N_3419,N_2976,N_2762);
nand U3420 (N_3420,N_2416,N_2868);
nand U3421 (N_3421,N_2609,N_2387);
xnor U3422 (N_3422,N_2497,N_2472);
nand U3423 (N_3423,N_2275,N_2749);
xnor U3424 (N_3424,N_2259,N_2370);
or U3425 (N_3425,N_2833,N_2910);
or U3426 (N_3426,N_2381,N_2542);
or U3427 (N_3427,N_2672,N_2838);
or U3428 (N_3428,N_2315,N_2835);
and U3429 (N_3429,N_2622,N_2531);
nand U3430 (N_3430,N_2958,N_2894);
nor U3431 (N_3431,N_2355,N_2662);
and U3432 (N_3432,N_2789,N_2325);
nand U3433 (N_3433,N_2977,N_2952);
nor U3434 (N_3434,N_2705,N_2914);
nor U3435 (N_3435,N_2626,N_2423);
nand U3436 (N_3436,N_2823,N_2678);
xnor U3437 (N_3437,N_2369,N_2288);
nand U3438 (N_3438,N_2442,N_2348);
nand U3439 (N_3439,N_2775,N_2718);
xor U3440 (N_3440,N_2514,N_2893);
nor U3441 (N_3441,N_2961,N_2570);
xnor U3442 (N_3442,N_2416,N_2656);
nand U3443 (N_3443,N_2511,N_2258);
nor U3444 (N_3444,N_2294,N_2371);
nor U3445 (N_3445,N_2776,N_2284);
nor U3446 (N_3446,N_2879,N_2561);
or U3447 (N_3447,N_2978,N_2403);
or U3448 (N_3448,N_2563,N_2912);
or U3449 (N_3449,N_2308,N_2699);
xor U3450 (N_3450,N_2747,N_2776);
or U3451 (N_3451,N_2381,N_2340);
nand U3452 (N_3452,N_2808,N_2399);
and U3453 (N_3453,N_2571,N_2608);
xnor U3454 (N_3454,N_2925,N_2668);
nor U3455 (N_3455,N_2272,N_2837);
and U3456 (N_3456,N_2673,N_2600);
and U3457 (N_3457,N_2482,N_2791);
xnor U3458 (N_3458,N_2265,N_2761);
or U3459 (N_3459,N_2822,N_2309);
nand U3460 (N_3460,N_2259,N_2720);
nand U3461 (N_3461,N_2902,N_2253);
nand U3462 (N_3462,N_2862,N_2799);
xor U3463 (N_3463,N_2747,N_2337);
nor U3464 (N_3464,N_2641,N_2808);
nor U3465 (N_3465,N_2742,N_2880);
nand U3466 (N_3466,N_2351,N_2638);
nor U3467 (N_3467,N_2453,N_2519);
xnor U3468 (N_3468,N_2269,N_2946);
xnor U3469 (N_3469,N_2298,N_2811);
xnor U3470 (N_3470,N_2419,N_2813);
nand U3471 (N_3471,N_2721,N_2350);
or U3472 (N_3472,N_2747,N_2858);
nor U3473 (N_3473,N_2431,N_2693);
nand U3474 (N_3474,N_2800,N_2957);
xor U3475 (N_3475,N_2535,N_2340);
nor U3476 (N_3476,N_2327,N_2273);
nor U3477 (N_3477,N_2445,N_2588);
and U3478 (N_3478,N_2520,N_2482);
nand U3479 (N_3479,N_2782,N_2777);
nor U3480 (N_3480,N_2965,N_2796);
and U3481 (N_3481,N_2932,N_2723);
nor U3482 (N_3482,N_2701,N_2352);
xor U3483 (N_3483,N_2885,N_2920);
nor U3484 (N_3484,N_2978,N_2753);
nand U3485 (N_3485,N_2399,N_2837);
xnor U3486 (N_3486,N_2486,N_2359);
nor U3487 (N_3487,N_2741,N_2999);
nor U3488 (N_3488,N_2453,N_2329);
and U3489 (N_3489,N_2945,N_2629);
and U3490 (N_3490,N_2590,N_2897);
xnor U3491 (N_3491,N_2875,N_2908);
or U3492 (N_3492,N_2885,N_2891);
nand U3493 (N_3493,N_2949,N_2941);
nor U3494 (N_3494,N_2315,N_2655);
nor U3495 (N_3495,N_2683,N_2461);
and U3496 (N_3496,N_2451,N_2645);
nor U3497 (N_3497,N_2380,N_2637);
and U3498 (N_3498,N_2521,N_2603);
xnor U3499 (N_3499,N_2670,N_2894);
or U3500 (N_3500,N_2541,N_2766);
nor U3501 (N_3501,N_2735,N_2541);
xnor U3502 (N_3502,N_2694,N_2842);
nor U3503 (N_3503,N_2990,N_2463);
and U3504 (N_3504,N_2866,N_2602);
nand U3505 (N_3505,N_2302,N_2379);
xor U3506 (N_3506,N_2724,N_2764);
nor U3507 (N_3507,N_2446,N_2942);
xor U3508 (N_3508,N_2729,N_2635);
nor U3509 (N_3509,N_2399,N_2623);
nor U3510 (N_3510,N_2450,N_2627);
nor U3511 (N_3511,N_2851,N_2819);
nand U3512 (N_3512,N_2302,N_2617);
nand U3513 (N_3513,N_2296,N_2913);
or U3514 (N_3514,N_2360,N_2391);
xor U3515 (N_3515,N_2388,N_2805);
or U3516 (N_3516,N_2621,N_2518);
nor U3517 (N_3517,N_2414,N_2554);
xnor U3518 (N_3518,N_2386,N_2708);
nand U3519 (N_3519,N_2656,N_2545);
nand U3520 (N_3520,N_2823,N_2425);
xnor U3521 (N_3521,N_2817,N_2585);
or U3522 (N_3522,N_2907,N_2698);
nor U3523 (N_3523,N_2322,N_2480);
or U3524 (N_3524,N_2310,N_2911);
or U3525 (N_3525,N_2882,N_2385);
nor U3526 (N_3526,N_2922,N_2725);
and U3527 (N_3527,N_2306,N_2611);
and U3528 (N_3528,N_2404,N_2554);
and U3529 (N_3529,N_2270,N_2872);
xnor U3530 (N_3530,N_2492,N_2668);
nor U3531 (N_3531,N_2577,N_2997);
nor U3532 (N_3532,N_2461,N_2838);
nand U3533 (N_3533,N_2691,N_2656);
or U3534 (N_3534,N_2593,N_2440);
and U3535 (N_3535,N_2468,N_2903);
xor U3536 (N_3536,N_2385,N_2647);
or U3537 (N_3537,N_2315,N_2955);
nand U3538 (N_3538,N_2499,N_2533);
nor U3539 (N_3539,N_2630,N_2864);
and U3540 (N_3540,N_2427,N_2607);
xor U3541 (N_3541,N_2787,N_2636);
or U3542 (N_3542,N_2551,N_2699);
and U3543 (N_3543,N_2457,N_2455);
and U3544 (N_3544,N_2996,N_2467);
xor U3545 (N_3545,N_2348,N_2319);
nand U3546 (N_3546,N_2762,N_2751);
xnor U3547 (N_3547,N_2359,N_2713);
and U3548 (N_3548,N_2848,N_2882);
nand U3549 (N_3549,N_2536,N_2984);
or U3550 (N_3550,N_2358,N_2497);
nand U3551 (N_3551,N_2669,N_2373);
xnor U3552 (N_3552,N_2624,N_2688);
or U3553 (N_3553,N_2786,N_2722);
xor U3554 (N_3554,N_2737,N_2617);
and U3555 (N_3555,N_2585,N_2474);
or U3556 (N_3556,N_2963,N_2820);
xnor U3557 (N_3557,N_2322,N_2474);
xnor U3558 (N_3558,N_2561,N_2282);
nand U3559 (N_3559,N_2282,N_2629);
xor U3560 (N_3560,N_2827,N_2316);
xor U3561 (N_3561,N_2374,N_2959);
and U3562 (N_3562,N_2381,N_2743);
and U3563 (N_3563,N_2567,N_2554);
or U3564 (N_3564,N_2556,N_2519);
xnor U3565 (N_3565,N_2805,N_2384);
nor U3566 (N_3566,N_2935,N_2839);
nand U3567 (N_3567,N_2930,N_2274);
nand U3568 (N_3568,N_2468,N_2705);
or U3569 (N_3569,N_2756,N_2538);
xnor U3570 (N_3570,N_2816,N_2388);
and U3571 (N_3571,N_2408,N_2636);
and U3572 (N_3572,N_2432,N_2350);
nor U3573 (N_3573,N_2997,N_2900);
and U3574 (N_3574,N_2263,N_2315);
nand U3575 (N_3575,N_2555,N_2749);
and U3576 (N_3576,N_2880,N_2732);
or U3577 (N_3577,N_2845,N_2653);
nand U3578 (N_3578,N_2813,N_2344);
nand U3579 (N_3579,N_2390,N_2765);
xor U3580 (N_3580,N_2576,N_2440);
or U3581 (N_3581,N_2918,N_2886);
xor U3582 (N_3582,N_2581,N_2572);
xnor U3583 (N_3583,N_2307,N_2480);
xnor U3584 (N_3584,N_2588,N_2620);
and U3585 (N_3585,N_2351,N_2867);
nand U3586 (N_3586,N_2822,N_2762);
nor U3587 (N_3587,N_2648,N_2508);
nand U3588 (N_3588,N_2926,N_2734);
nand U3589 (N_3589,N_2840,N_2771);
or U3590 (N_3590,N_2959,N_2530);
or U3591 (N_3591,N_2360,N_2739);
nor U3592 (N_3592,N_2698,N_2394);
nor U3593 (N_3593,N_2674,N_2807);
nand U3594 (N_3594,N_2690,N_2766);
nor U3595 (N_3595,N_2305,N_2434);
xor U3596 (N_3596,N_2321,N_2981);
and U3597 (N_3597,N_2988,N_2459);
nor U3598 (N_3598,N_2563,N_2923);
or U3599 (N_3599,N_2706,N_2812);
nor U3600 (N_3600,N_2502,N_2316);
xnor U3601 (N_3601,N_2563,N_2427);
nor U3602 (N_3602,N_2572,N_2987);
and U3603 (N_3603,N_2862,N_2595);
xor U3604 (N_3604,N_2949,N_2718);
nand U3605 (N_3605,N_2543,N_2871);
or U3606 (N_3606,N_2846,N_2540);
nand U3607 (N_3607,N_2525,N_2572);
nor U3608 (N_3608,N_2252,N_2954);
nand U3609 (N_3609,N_2962,N_2517);
or U3610 (N_3610,N_2655,N_2850);
nand U3611 (N_3611,N_2267,N_2559);
nand U3612 (N_3612,N_2332,N_2933);
xnor U3613 (N_3613,N_2578,N_2454);
xnor U3614 (N_3614,N_2727,N_2737);
nor U3615 (N_3615,N_2507,N_2702);
or U3616 (N_3616,N_2599,N_2859);
xnor U3617 (N_3617,N_2934,N_2522);
nand U3618 (N_3618,N_2389,N_2466);
and U3619 (N_3619,N_2793,N_2673);
xnor U3620 (N_3620,N_2696,N_2627);
nand U3621 (N_3621,N_2382,N_2744);
nand U3622 (N_3622,N_2827,N_2284);
or U3623 (N_3623,N_2916,N_2293);
xnor U3624 (N_3624,N_2751,N_2849);
and U3625 (N_3625,N_2589,N_2633);
or U3626 (N_3626,N_2710,N_2902);
or U3627 (N_3627,N_2519,N_2941);
and U3628 (N_3628,N_2295,N_2351);
nor U3629 (N_3629,N_2947,N_2972);
nand U3630 (N_3630,N_2802,N_2573);
or U3631 (N_3631,N_2960,N_2761);
nand U3632 (N_3632,N_2733,N_2785);
nor U3633 (N_3633,N_2646,N_2666);
or U3634 (N_3634,N_2813,N_2880);
xor U3635 (N_3635,N_2439,N_2332);
xnor U3636 (N_3636,N_2265,N_2655);
xor U3637 (N_3637,N_2986,N_2444);
or U3638 (N_3638,N_2496,N_2251);
or U3639 (N_3639,N_2705,N_2767);
and U3640 (N_3640,N_2413,N_2769);
xnor U3641 (N_3641,N_2313,N_2842);
nand U3642 (N_3642,N_2631,N_2274);
xnor U3643 (N_3643,N_2910,N_2816);
nand U3644 (N_3644,N_2472,N_2503);
xor U3645 (N_3645,N_2607,N_2797);
and U3646 (N_3646,N_2774,N_2553);
nand U3647 (N_3647,N_2823,N_2699);
and U3648 (N_3648,N_2326,N_2738);
or U3649 (N_3649,N_2437,N_2398);
nor U3650 (N_3650,N_2915,N_2786);
nor U3651 (N_3651,N_2867,N_2554);
and U3652 (N_3652,N_2943,N_2587);
and U3653 (N_3653,N_2624,N_2922);
nor U3654 (N_3654,N_2443,N_2541);
or U3655 (N_3655,N_2773,N_2361);
nand U3656 (N_3656,N_2417,N_2468);
and U3657 (N_3657,N_2827,N_2804);
nand U3658 (N_3658,N_2356,N_2930);
nor U3659 (N_3659,N_2683,N_2432);
nand U3660 (N_3660,N_2489,N_2334);
or U3661 (N_3661,N_2293,N_2605);
xor U3662 (N_3662,N_2356,N_2331);
nor U3663 (N_3663,N_2889,N_2749);
and U3664 (N_3664,N_2638,N_2551);
nor U3665 (N_3665,N_2664,N_2314);
and U3666 (N_3666,N_2497,N_2827);
nor U3667 (N_3667,N_2880,N_2677);
nor U3668 (N_3668,N_2747,N_2473);
nand U3669 (N_3669,N_2524,N_2335);
and U3670 (N_3670,N_2906,N_2652);
and U3671 (N_3671,N_2362,N_2488);
xnor U3672 (N_3672,N_2487,N_2932);
or U3673 (N_3673,N_2437,N_2629);
or U3674 (N_3674,N_2981,N_2754);
or U3675 (N_3675,N_2457,N_2631);
nand U3676 (N_3676,N_2839,N_2304);
nor U3677 (N_3677,N_2638,N_2324);
xor U3678 (N_3678,N_2915,N_2642);
nand U3679 (N_3679,N_2409,N_2859);
nand U3680 (N_3680,N_2345,N_2293);
nor U3681 (N_3681,N_2440,N_2778);
and U3682 (N_3682,N_2597,N_2849);
nor U3683 (N_3683,N_2960,N_2331);
nand U3684 (N_3684,N_2750,N_2429);
or U3685 (N_3685,N_2750,N_2932);
and U3686 (N_3686,N_2687,N_2327);
or U3687 (N_3687,N_2837,N_2715);
nand U3688 (N_3688,N_2622,N_2614);
and U3689 (N_3689,N_2994,N_2777);
xor U3690 (N_3690,N_2941,N_2650);
or U3691 (N_3691,N_2679,N_2458);
and U3692 (N_3692,N_2286,N_2731);
or U3693 (N_3693,N_2594,N_2597);
or U3694 (N_3694,N_2281,N_2379);
or U3695 (N_3695,N_2712,N_2851);
xor U3696 (N_3696,N_2634,N_2274);
nor U3697 (N_3697,N_2740,N_2685);
and U3698 (N_3698,N_2515,N_2925);
xor U3699 (N_3699,N_2830,N_2386);
or U3700 (N_3700,N_2280,N_2760);
nor U3701 (N_3701,N_2885,N_2323);
nor U3702 (N_3702,N_2655,N_2250);
and U3703 (N_3703,N_2353,N_2768);
nand U3704 (N_3704,N_2645,N_2602);
nor U3705 (N_3705,N_2464,N_2848);
xor U3706 (N_3706,N_2270,N_2268);
xnor U3707 (N_3707,N_2701,N_2866);
nand U3708 (N_3708,N_2349,N_2322);
and U3709 (N_3709,N_2996,N_2797);
nand U3710 (N_3710,N_2903,N_2497);
nand U3711 (N_3711,N_2795,N_2790);
and U3712 (N_3712,N_2758,N_2339);
nor U3713 (N_3713,N_2971,N_2385);
xor U3714 (N_3714,N_2692,N_2982);
or U3715 (N_3715,N_2617,N_2273);
and U3716 (N_3716,N_2520,N_2481);
nor U3717 (N_3717,N_2522,N_2987);
nand U3718 (N_3718,N_2470,N_2483);
nand U3719 (N_3719,N_2925,N_2453);
and U3720 (N_3720,N_2735,N_2767);
and U3721 (N_3721,N_2617,N_2341);
nor U3722 (N_3722,N_2375,N_2752);
and U3723 (N_3723,N_2270,N_2861);
xor U3724 (N_3724,N_2923,N_2733);
and U3725 (N_3725,N_2859,N_2639);
xnor U3726 (N_3726,N_2868,N_2328);
and U3727 (N_3727,N_2906,N_2531);
or U3728 (N_3728,N_2429,N_2726);
nand U3729 (N_3729,N_2538,N_2593);
nor U3730 (N_3730,N_2523,N_2575);
or U3731 (N_3731,N_2693,N_2776);
or U3732 (N_3732,N_2561,N_2934);
and U3733 (N_3733,N_2519,N_2351);
nand U3734 (N_3734,N_2932,N_2646);
and U3735 (N_3735,N_2655,N_2395);
or U3736 (N_3736,N_2859,N_2597);
nand U3737 (N_3737,N_2267,N_2295);
or U3738 (N_3738,N_2419,N_2737);
and U3739 (N_3739,N_2615,N_2800);
nor U3740 (N_3740,N_2465,N_2598);
nor U3741 (N_3741,N_2611,N_2312);
nor U3742 (N_3742,N_2510,N_2908);
nand U3743 (N_3743,N_2968,N_2697);
nor U3744 (N_3744,N_2449,N_2803);
or U3745 (N_3745,N_2959,N_2642);
nand U3746 (N_3746,N_2335,N_2329);
or U3747 (N_3747,N_2311,N_2807);
xnor U3748 (N_3748,N_2478,N_2657);
and U3749 (N_3749,N_2304,N_2805);
xor U3750 (N_3750,N_3040,N_3704);
xor U3751 (N_3751,N_3315,N_3433);
or U3752 (N_3752,N_3193,N_3312);
and U3753 (N_3753,N_3118,N_3403);
or U3754 (N_3754,N_3094,N_3304);
xor U3755 (N_3755,N_3462,N_3502);
xnor U3756 (N_3756,N_3586,N_3420);
or U3757 (N_3757,N_3331,N_3386);
nand U3758 (N_3758,N_3529,N_3722);
xnor U3759 (N_3759,N_3541,N_3680);
nor U3760 (N_3760,N_3229,N_3011);
nor U3761 (N_3761,N_3689,N_3519);
xnor U3762 (N_3762,N_3300,N_3074);
or U3763 (N_3763,N_3327,N_3592);
xnor U3764 (N_3764,N_3188,N_3336);
or U3765 (N_3765,N_3072,N_3309);
and U3766 (N_3766,N_3718,N_3371);
nand U3767 (N_3767,N_3170,N_3091);
or U3768 (N_3768,N_3552,N_3658);
nand U3769 (N_3769,N_3534,N_3046);
nand U3770 (N_3770,N_3267,N_3477);
xnor U3771 (N_3771,N_3104,N_3106);
and U3772 (N_3772,N_3512,N_3626);
nand U3773 (N_3773,N_3014,N_3060);
or U3774 (N_3774,N_3348,N_3044);
xnor U3775 (N_3775,N_3307,N_3232);
xor U3776 (N_3776,N_3634,N_3198);
nor U3777 (N_3777,N_3730,N_3292);
nor U3778 (N_3778,N_3451,N_3489);
xnor U3779 (N_3779,N_3164,N_3306);
xnor U3780 (N_3780,N_3368,N_3153);
nand U3781 (N_3781,N_3676,N_3570);
and U3782 (N_3782,N_3572,N_3700);
or U3783 (N_3783,N_3407,N_3135);
xor U3784 (N_3784,N_3655,N_3602);
or U3785 (N_3785,N_3498,N_3739);
nor U3786 (N_3786,N_3314,N_3644);
or U3787 (N_3787,N_3578,N_3082);
nand U3788 (N_3788,N_3696,N_3562);
and U3789 (N_3789,N_3151,N_3338);
or U3790 (N_3790,N_3733,N_3621);
or U3791 (N_3791,N_3346,N_3487);
nor U3792 (N_3792,N_3027,N_3440);
nand U3793 (N_3793,N_3488,N_3654);
xnor U3794 (N_3794,N_3035,N_3050);
xnor U3795 (N_3795,N_3693,N_3375);
or U3796 (N_3796,N_3390,N_3418);
or U3797 (N_3797,N_3206,N_3140);
xnor U3798 (N_3798,N_3748,N_3001);
xor U3799 (N_3799,N_3464,N_3583);
nand U3800 (N_3800,N_3340,N_3123);
and U3801 (N_3801,N_3731,N_3650);
nand U3802 (N_3802,N_3182,N_3402);
nor U3803 (N_3803,N_3128,N_3246);
nand U3804 (N_3804,N_3162,N_3528);
xor U3805 (N_3805,N_3501,N_3495);
xor U3806 (N_3806,N_3690,N_3516);
or U3807 (N_3807,N_3115,N_3645);
or U3808 (N_3808,N_3593,N_3203);
nand U3809 (N_3809,N_3530,N_3190);
and U3810 (N_3810,N_3152,N_3125);
or U3811 (N_3811,N_3373,N_3486);
xor U3812 (N_3812,N_3185,N_3301);
xor U3813 (N_3813,N_3025,N_3699);
xnor U3814 (N_3814,N_3241,N_3325);
and U3815 (N_3815,N_3132,N_3350);
nand U3816 (N_3816,N_3098,N_3565);
nor U3817 (N_3817,N_3735,N_3414);
and U3818 (N_3818,N_3540,N_3354);
nand U3819 (N_3819,N_3026,N_3558);
nor U3820 (N_3820,N_3449,N_3353);
and U3821 (N_3821,N_3511,N_3308);
or U3822 (N_3822,N_3201,N_3251);
nand U3823 (N_3823,N_3591,N_3417);
and U3824 (N_3824,N_3559,N_3461);
or U3825 (N_3825,N_3083,N_3599);
or U3826 (N_3826,N_3439,N_3223);
xor U3827 (N_3827,N_3169,N_3505);
xnor U3828 (N_3828,N_3159,N_3313);
and U3829 (N_3829,N_3741,N_3727);
nand U3830 (N_3830,N_3380,N_3549);
nor U3831 (N_3831,N_3265,N_3036);
xnor U3832 (N_3832,N_3577,N_3367);
and U3833 (N_3833,N_3701,N_3432);
and U3834 (N_3834,N_3598,N_3250);
xor U3835 (N_3835,N_3023,N_3204);
and U3836 (N_3836,N_3228,N_3149);
and U3837 (N_3837,N_3419,N_3335);
or U3838 (N_3838,N_3446,N_3337);
xor U3839 (N_3839,N_3225,N_3318);
or U3840 (N_3840,N_3343,N_3005);
nand U3841 (N_3841,N_3475,N_3588);
xnor U3842 (N_3842,N_3341,N_3471);
or U3843 (N_3843,N_3714,N_3435);
xor U3844 (N_3844,N_3608,N_3288);
xnor U3845 (N_3845,N_3394,N_3527);
nor U3846 (N_3846,N_3723,N_3345);
nand U3847 (N_3847,N_3127,N_3736);
and U3848 (N_3848,N_3453,N_3479);
or U3849 (N_3849,N_3236,N_3647);
nand U3850 (N_3850,N_3037,N_3352);
xor U3851 (N_3851,N_3580,N_3356);
xnor U3852 (N_3852,N_3103,N_3284);
or U3853 (N_3853,N_3065,N_3737);
or U3854 (N_3854,N_3447,N_3728);
nor U3855 (N_3855,N_3084,N_3016);
or U3856 (N_3856,N_3633,N_3154);
nor U3857 (N_3857,N_3042,N_3450);
nor U3858 (N_3858,N_3444,N_3085);
nor U3859 (N_3859,N_3073,N_3518);
nor U3860 (N_3860,N_3101,N_3454);
and U3861 (N_3861,N_3632,N_3218);
and U3862 (N_3862,N_3076,N_3720);
xor U3863 (N_3863,N_3653,N_3347);
or U3864 (N_3864,N_3155,N_3317);
xor U3865 (N_3865,N_3648,N_3584);
nor U3866 (N_3866,N_3405,N_3499);
or U3867 (N_3867,N_3744,N_3017);
xnor U3868 (N_3868,N_3000,N_3429);
or U3869 (N_3869,N_3176,N_3636);
xor U3870 (N_3870,N_3525,N_3514);
nand U3871 (N_3871,N_3482,N_3247);
nor U3872 (N_3872,N_3706,N_3726);
xnor U3873 (N_3873,N_3209,N_3329);
nor U3874 (N_3874,N_3692,N_3271);
nand U3875 (N_3875,N_3242,N_3561);
and U3876 (N_3876,N_3674,N_3319);
xor U3877 (N_3877,N_3585,N_3551);
nor U3878 (N_3878,N_3532,N_3517);
xor U3879 (N_3879,N_3253,N_3717);
and U3880 (N_3880,N_3493,N_3360);
nor U3881 (N_3881,N_3576,N_3199);
nand U3882 (N_3882,N_3055,N_3434);
xnor U3883 (N_3883,N_3243,N_3651);
xor U3884 (N_3884,N_3497,N_3660);
nand U3885 (N_3885,N_3226,N_3355);
and U3886 (N_3886,N_3630,N_3470);
or U3887 (N_3887,N_3504,N_3202);
nor U3888 (N_3888,N_3178,N_3589);
and U3889 (N_3889,N_3740,N_3535);
or U3890 (N_3890,N_3569,N_3205);
nor U3891 (N_3891,N_3483,N_3705);
or U3892 (N_3892,N_3034,N_3192);
or U3893 (N_3893,N_3274,N_3062);
xor U3894 (N_3894,N_3183,N_3652);
and U3895 (N_3895,N_3332,N_3485);
or U3896 (N_3896,N_3452,N_3460);
xor U3897 (N_3897,N_3078,N_3550);
xnor U3898 (N_3898,N_3066,N_3625);
xor U3899 (N_3899,N_3004,N_3289);
nor U3900 (N_3900,N_3404,N_3372);
nor U3901 (N_3901,N_3184,N_3662);
or U3902 (N_3902,N_3745,N_3045);
nor U3903 (N_3903,N_3048,N_3299);
nor U3904 (N_3904,N_3702,N_3377);
xnor U3905 (N_3905,N_3145,N_3133);
xnor U3906 (N_3906,N_3285,N_3095);
and U3907 (N_3907,N_3472,N_3738);
nand U3908 (N_3908,N_3039,N_3290);
or U3909 (N_3909,N_3665,N_3208);
nand U3910 (N_3910,N_3494,N_3721);
or U3911 (N_3911,N_3234,N_3413);
or U3912 (N_3912,N_3165,N_3713);
xnor U3913 (N_3913,N_3422,N_3694);
nor U3914 (N_3914,N_3112,N_3677);
xor U3915 (N_3915,N_3672,N_3492);
xor U3916 (N_3916,N_3051,N_3138);
nor U3917 (N_3917,N_3544,N_3456);
nand U3918 (N_3918,N_3370,N_3020);
and U3919 (N_3919,N_3607,N_3266);
and U3920 (N_3920,N_3698,N_3294);
nand U3921 (N_3921,N_3620,N_3349);
and U3922 (N_3922,N_3646,N_3216);
or U3923 (N_3923,N_3656,N_3227);
xor U3924 (N_3924,N_3575,N_3622);
nor U3925 (N_3925,N_3533,N_3709);
xnor U3926 (N_3926,N_3379,N_3161);
xnor U3927 (N_3927,N_3508,N_3100);
xnor U3928 (N_3928,N_3590,N_3070);
nand U3929 (N_3929,N_3542,N_3049);
and U3930 (N_3930,N_3120,N_3029);
or U3931 (N_3931,N_3381,N_3515);
nand U3932 (N_3932,N_3171,N_3272);
nor U3933 (N_3933,N_3087,N_3032);
and U3934 (N_3934,N_3015,N_3137);
xnor U3935 (N_3935,N_3522,N_3142);
and U3936 (N_3936,N_3566,N_3129);
nor U3937 (N_3937,N_3261,N_3631);
nor U3938 (N_3938,N_3537,N_3605);
or U3939 (N_3939,N_3316,N_3437);
nand U3940 (N_3940,N_3712,N_3093);
or U3941 (N_3941,N_3415,N_3252);
and U3942 (N_3942,N_3276,N_3238);
nor U3943 (N_3943,N_3640,N_3215);
or U3944 (N_3944,N_3323,N_3742);
or U3945 (N_3945,N_3364,N_3684);
xnor U3946 (N_3946,N_3611,N_3280);
nor U3947 (N_3947,N_3409,N_3695);
nand U3948 (N_3948,N_3330,N_3090);
or U3949 (N_3949,N_3595,N_3028);
xor U3950 (N_3950,N_3510,N_3436);
nor U3951 (N_3951,N_3196,N_3715);
xnor U3952 (N_3952,N_3217,N_3030);
xor U3953 (N_3953,N_3428,N_3716);
or U3954 (N_3954,N_3298,N_3054);
xnor U3955 (N_3955,N_3326,N_3059);
and U3956 (N_3956,N_3222,N_3391);
or U3957 (N_3957,N_3427,N_3211);
nand U3958 (N_3958,N_3099,N_3177);
nand U3959 (N_3959,N_3642,N_3295);
nand U3960 (N_3960,N_3043,N_3121);
nor U3961 (N_3961,N_3233,N_3089);
and U3962 (N_3962,N_3708,N_3457);
nor U3963 (N_3963,N_3130,N_3679);
or U3964 (N_3964,N_3052,N_3606);
xnor U3965 (N_3965,N_3109,N_3675);
xnor U3966 (N_3966,N_3134,N_3594);
xnor U3967 (N_3967,N_3102,N_3003);
or U3968 (N_3968,N_3174,N_3500);
and U3969 (N_3969,N_3412,N_3547);
and U3970 (N_3970,N_3310,N_3546);
or U3971 (N_3971,N_3442,N_3627);
nor U3972 (N_3972,N_3603,N_3264);
or U3973 (N_3973,N_3416,N_3168);
nand U3974 (N_3974,N_3333,N_3568);
nand U3975 (N_3975,N_3061,N_3021);
and U3976 (N_3976,N_3641,N_3081);
or U3977 (N_3977,N_3022,N_3671);
and U3978 (N_3978,N_3615,N_3195);
or U3979 (N_3979,N_3013,N_3673);
nor U3980 (N_3980,N_3273,N_3197);
nand U3981 (N_3981,N_3678,N_3571);
and U3982 (N_3982,N_3448,N_3408);
nand U3983 (N_3983,N_3543,N_3322);
nor U3984 (N_3984,N_3012,N_3053);
xnor U3985 (N_3985,N_3554,N_3459);
or U3986 (N_3986,N_3255,N_3361);
or U3987 (N_3987,N_3351,N_3581);
nand U3988 (N_3988,N_3619,N_3080);
xor U3989 (N_3989,N_3382,N_3220);
nand U3990 (N_3990,N_3269,N_3245);
xor U3991 (N_3991,N_3524,N_3423);
or U3992 (N_3992,N_3038,N_3019);
or U3993 (N_3993,N_3363,N_3659);
xnor U3994 (N_3994,N_3430,N_3231);
or U3995 (N_3995,N_3669,N_3268);
nand U3996 (N_3996,N_3237,N_3111);
and U3997 (N_3997,N_3207,N_3173);
xnor U3998 (N_3998,N_3564,N_3200);
nand U3999 (N_3999,N_3521,N_3263);
nand U4000 (N_4000,N_3638,N_3088);
nand U4001 (N_4001,N_3224,N_3002);
xor U4002 (N_4002,N_3277,N_3139);
nand U4003 (N_4003,N_3710,N_3393);
and U4004 (N_4004,N_3425,N_3063);
xnor U4005 (N_4005,N_3618,N_3555);
nor U4006 (N_4006,N_3548,N_3279);
nand U4007 (N_4007,N_3743,N_3240);
nor U4008 (N_4008,N_3383,N_3661);
or U4009 (N_4009,N_3281,N_3366);
nor U4010 (N_4010,N_3579,N_3136);
nand U4011 (N_4011,N_3041,N_3376);
and U4012 (N_4012,N_3320,N_3126);
and U4013 (N_4013,N_3725,N_3538);
xor U4014 (N_4014,N_3610,N_3270);
or U4015 (N_4015,N_3746,N_3141);
xor U4016 (N_4016,N_3275,N_3324);
xnor U4017 (N_4017,N_3321,N_3010);
nand U4018 (N_4018,N_3328,N_3186);
xor U4019 (N_4019,N_3445,N_3158);
or U4020 (N_4020,N_3406,N_3068);
nor U4021 (N_4021,N_3385,N_3703);
or U4022 (N_4022,N_3374,N_3557);
and U4023 (N_4023,N_3596,N_3431);
xnor U4024 (N_4024,N_3293,N_3635);
or U4025 (N_4025,N_3387,N_3358);
or U4026 (N_4026,N_3210,N_3481);
nand U4027 (N_4027,N_3563,N_3526);
nor U4028 (N_4028,N_3007,N_3567);
and U4029 (N_4029,N_3248,N_3629);
and U4030 (N_4030,N_3399,N_3681);
or U4031 (N_4031,N_3180,N_3480);
nor U4032 (N_4032,N_3249,N_3008);
nand U4033 (N_4033,N_3484,N_3587);
xnor U4034 (N_4034,N_3146,N_3378);
nor U4035 (N_4035,N_3302,N_3262);
and U4036 (N_4036,N_3219,N_3469);
nand U4037 (N_4037,N_3064,N_3221);
xor U4038 (N_4038,N_3296,N_3258);
and U4039 (N_4039,N_3663,N_3212);
or U4040 (N_4040,N_3560,N_3401);
and U4041 (N_4041,N_3411,N_3410);
nand U4042 (N_4042,N_3024,N_3006);
and U4043 (N_4043,N_3697,N_3092);
nor U4044 (N_4044,N_3286,N_3131);
nand U4045 (N_4045,N_3172,N_3667);
xor U4046 (N_4046,N_3079,N_3613);
and U4047 (N_4047,N_3110,N_3597);
nor U4048 (N_4048,N_3235,N_3463);
and U4049 (N_4049,N_3664,N_3144);
nor U4050 (N_4050,N_3707,N_3114);
or U4051 (N_4051,N_3254,N_3283);
or U4052 (N_4052,N_3291,N_3166);
and U4053 (N_4053,N_3637,N_3628);
xor U4054 (N_4054,N_3749,N_3732);
nand U4055 (N_4055,N_3392,N_3574);
and U4056 (N_4056,N_3031,N_3438);
xor U4057 (N_4057,N_3339,N_3069);
nand U4058 (N_4058,N_3476,N_3455);
or U4059 (N_4059,N_3617,N_3124);
xnor U4060 (N_4060,N_3724,N_3282);
nor U4061 (N_4061,N_3513,N_3441);
xor U4062 (N_4062,N_3175,N_3157);
nand U4063 (N_4063,N_3711,N_3604);
or U4064 (N_4064,N_3478,N_3400);
nor U4065 (N_4065,N_3396,N_3311);
and U4066 (N_4066,N_3362,N_3058);
or U4067 (N_4067,N_3458,N_3107);
nor U4068 (N_4068,N_3278,N_3624);
xor U4069 (N_4069,N_3384,N_3682);
nand U4070 (N_4070,N_3729,N_3057);
nor U4071 (N_4071,N_3421,N_3520);
nand U4072 (N_4072,N_3683,N_3213);
nor U4073 (N_4073,N_3342,N_3297);
and U4074 (N_4074,N_3531,N_3056);
nand U4075 (N_4075,N_3097,N_3156);
xnor U4076 (N_4076,N_3389,N_3506);
nor U4077 (N_4077,N_3194,N_3167);
xor U4078 (N_4078,N_3649,N_3719);
nor U4079 (N_4079,N_3067,N_3116);
nand U4080 (N_4080,N_3287,N_3614);
xor U4081 (N_4081,N_3260,N_3473);
or U4082 (N_4082,N_3122,N_3344);
xor U4083 (N_4083,N_3443,N_3147);
nand U4084 (N_4084,N_3179,N_3105);
xor U4085 (N_4085,N_3685,N_3623);
or U4086 (N_4086,N_3490,N_3071);
nand U4087 (N_4087,N_3113,N_3119);
nor U4088 (N_4088,N_3334,N_3686);
nor U4089 (N_4089,N_3303,N_3507);
xor U4090 (N_4090,N_3256,N_3181);
nand U4091 (N_4091,N_3600,N_3369);
nor U4092 (N_4092,N_3474,N_3357);
or U4093 (N_4093,N_3230,N_3668);
xnor U4094 (N_4094,N_3573,N_3747);
and U4095 (N_4095,N_3259,N_3466);
and U4096 (N_4096,N_3305,N_3734);
xor U4097 (N_4097,N_3601,N_3009);
nor U4098 (N_4098,N_3609,N_3657);
and U4099 (N_4099,N_3616,N_3018);
and U4100 (N_4100,N_3397,N_3687);
xnor U4101 (N_4101,N_3424,N_3670);
nor U4102 (N_4102,N_3691,N_3395);
nand U4103 (N_4103,N_3191,N_3148);
xnor U4104 (N_4104,N_3359,N_3639);
xnor U4105 (N_4105,N_3491,N_3143);
nand U4106 (N_4106,N_3465,N_3496);
nand U4107 (N_4107,N_3582,N_3047);
or U4108 (N_4108,N_3545,N_3257);
xor U4109 (N_4109,N_3033,N_3553);
or U4110 (N_4110,N_3077,N_3688);
or U4111 (N_4111,N_3086,N_3503);
and U4112 (N_4112,N_3117,N_3163);
nor U4113 (N_4113,N_3523,N_3426);
nor U4114 (N_4114,N_3556,N_3509);
and U4115 (N_4115,N_3536,N_3187);
nand U4116 (N_4116,N_3398,N_3666);
nor U4117 (N_4117,N_3160,N_3096);
and U4118 (N_4118,N_3075,N_3468);
xor U4119 (N_4119,N_3150,N_3214);
xnor U4120 (N_4120,N_3643,N_3612);
nand U4121 (N_4121,N_3244,N_3365);
xnor U4122 (N_4122,N_3388,N_3189);
nor U4123 (N_4123,N_3239,N_3467);
or U4124 (N_4124,N_3108,N_3539);
nand U4125 (N_4125,N_3325,N_3637);
xnor U4126 (N_4126,N_3241,N_3521);
or U4127 (N_4127,N_3747,N_3639);
and U4128 (N_4128,N_3725,N_3372);
nor U4129 (N_4129,N_3534,N_3539);
nand U4130 (N_4130,N_3272,N_3542);
xnor U4131 (N_4131,N_3540,N_3054);
nand U4132 (N_4132,N_3468,N_3630);
nor U4133 (N_4133,N_3384,N_3575);
nand U4134 (N_4134,N_3065,N_3039);
or U4135 (N_4135,N_3679,N_3052);
nand U4136 (N_4136,N_3514,N_3600);
nor U4137 (N_4137,N_3259,N_3638);
nor U4138 (N_4138,N_3024,N_3437);
nor U4139 (N_4139,N_3116,N_3375);
xnor U4140 (N_4140,N_3364,N_3182);
or U4141 (N_4141,N_3074,N_3710);
nand U4142 (N_4142,N_3136,N_3601);
xnor U4143 (N_4143,N_3667,N_3119);
and U4144 (N_4144,N_3411,N_3723);
and U4145 (N_4145,N_3564,N_3051);
nand U4146 (N_4146,N_3398,N_3174);
and U4147 (N_4147,N_3720,N_3128);
or U4148 (N_4148,N_3474,N_3618);
nand U4149 (N_4149,N_3022,N_3560);
or U4150 (N_4150,N_3077,N_3675);
or U4151 (N_4151,N_3644,N_3247);
xor U4152 (N_4152,N_3195,N_3010);
nand U4153 (N_4153,N_3360,N_3040);
nor U4154 (N_4154,N_3727,N_3551);
nor U4155 (N_4155,N_3743,N_3355);
and U4156 (N_4156,N_3375,N_3481);
or U4157 (N_4157,N_3566,N_3074);
xnor U4158 (N_4158,N_3115,N_3003);
and U4159 (N_4159,N_3730,N_3661);
or U4160 (N_4160,N_3299,N_3733);
or U4161 (N_4161,N_3256,N_3394);
or U4162 (N_4162,N_3432,N_3375);
xnor U4163 (N_4163,N_3426,N_3708);
nand U4164 (N_4164,N_3263,N_3317);
nand U4165 (N_4165,N_3480,N_3478);
xor U4166 (N_4166,N_3522,N_3120);
nor U4167 (N_4167,N_3651,N_3144);
or U4168 (N_4168,N_3598,N_3659);
and U4169 (N_4169,N_3325,N_3175);
or U4170 (N_4170,N_3226,N_3512);
xor U4171 (N_4171,N_3284,N_3244);
xor U4172 (N_4172,N_3437,N_3395);
xnor U4173 (N_4173,N_3467,N_3220);
xor U4174 (N_4174,N_3308,N_3675);
nand U4175 (N_4175,N_3332,N_3636);
and U4176 (N_4176,N_3263,N_3705);
xor U4177 (N_4177,N_3382,N_3132);
or U4178 (N_4178,N_3344,N_3085);
xnor U4179 (N_4179,N_3031,N_3560);
or U4180 (N_4180,N_3438,N_3122);
nor U4181 (N_4181,N_3526,N_3008);
and U4182 (N_4182,N_3331,N_3282);
or U4183 (N_4183,N_3562,N_3744);
xnor U4184 (N_4184,N_3161,N_3528);
nor U4185 (N_4185,N_3434,N_3718);
or U4186 (N_4186,N_3598,N_3022);
and U4187 (N_4187,N_3413,N_3459);
xnor U4188 (N_4188,N_3305,N_3240);
nand U4189 (N_4189,N_3521,N_3157);
xnor U4190 (N_4190,N_3597,N_3699);
nor U4191 (N_4191,N_3335,N_3264);
and U4192 (N_4192,N_3307,N_3143);
and U4193 (N_4193,N_3158,N_3617);
nor U4194 (N_4194,N_3255,N_3081);
nor U4195 (N_4195,N_3139,N_3469);
nand U4196 (N_4196,N_3734,N_3375);
nand U4197 (N_4197,N_3662,N_3658);
nand U4198 (N_4198,N_3354,N_3377);
nor U4199 (N_4199,N_3711,N_3657);
xor U4200 (N_4200,N_3430,N_3535);
xor U4201 (N_4201,N_3217,N_3498);
or U4202 (N_4202,N_3218,N_3133);
or U4203 (N_4203,N_3536,N_3301);
or U4204 (N_4204,N_3362,N_3720);
and U4205 (N_4205,N_3088,N_3242);
nand U4206 (N_4206,N_3096,N_3659);
nand U4207 (N_4207,N_3737,N_3732);
xor U4208 (N_4208,N_3481,N_3239);
nand U4209 (N_4209,N_3735,N_3189);
and U4210 (N_4210,N_3481,N_3685);
xnor U4211 (N_4211,N_3177,N_3047);
and U4212 (N_4212,N_3551,N_3239);
nor U4213 (N_4213,N_3411,N_3339);
xor U4214 (N_4214,N_3745,N_3609);
xor U4215 (N_4215,N_3148,N_3460);
and U4216 (N_4216,N_3129,N_3620);
or U4217 (N_4217,N_3317,N_3451);
and U4218 (N_4218,N_3595,N_3185);
nand U4219 (N_4219,N_3566,N_3200);
nand U4220 (N_4220,N_3383,N_3734);
xnor U4221 (N_4221,N_3230,N_3290);
nor U4222 (N_4222,N_3379,N_3073);
nand U4223 (N_4223,N_3082,N_3197);
xnor U4224 (N_4224,N_3135,N_3535);
nor U4225 (N_4225,N_3682,N_3440);
or U4226 (N_4226,N_3406,N_3528);
nand U4227 (N_4227,N_3409,N_3528);
and U4228 (N_4228,N_3290,N_3239);
nor U4229 (N_4229,N_3469,N_3692);
nor U4230 (N_4230,N_3234,N_3616);
and U4231 (N_4231,N_3539,N_3217);
nand U4232 (N_4232,N_3335,N_3108);
and U4233 (N_4233,N_3702,N_3463);
nand U4234 (N_4234,N_3499,N_3585);
nor U4235 (N_4235,N_3401,N_3203);
xor U4236 (N_4236,N_3267,N_3630);
or U4237 (N_4237,N_3205,N_3164);
or U4238 (N_4238,N_3630,N_3118);
nand U4239 (N_4239,N_3087,N_3666);
and U4240 (N_4240,N_3626,N_3398);
xor U4241 (N_4241,N_3619,N_3379);
nand U4242 (N_4242,N_3659,N_3371);
or U4243 (N_4243,N_3287,N_3361);
nor U4244 (N_4244,N_3389,N_3018);
and U4245 (N_4245,N_3535,N_3641);
or U4246 (N_4246,N_3466,N_3622);
nor U4247 (N_4247,N_3340,N_3389);
or U4248 (N_4248,N_3061,N_3025);
nor U4249 (N_4249,N_3117,N_3194);
and U4250 (N_4250,N_3013,N_3105);
nor U4251 (N_4251,N_3531,N_3351);
nand U4252 (N_4252,N_3506,N_3456);
nor U4253 (N_4253,N_3125,N_3167);
xor U4254 (N_4254,N_3040,N_3162);
nor U4255 (N_4255,N_3693,N_3403);
xor U4256 (N_4256,N_3581,N_3088);
nor U4257 (N_4257,N_3199,N_3519);
and U4258 (N_4258,N_3617,N_3121);
nand U4259 (N_4259,N_3629,N_3161);
nand U4260 (N_4260,N_3653,N_3555);
nor U4261 (N_4261,N_3688,N_3177);
or U4262 (N_4262,N_3532,N_3569);
or U4263 (N_4263,N_3008,N_3728);
and U4264 (N_4264,N_3106,N_3428);
or U4265 (N_4265,N_3721,N_3741);
or U4266 (N_4266,N_3178,N_3211);
xor U4267 (N_4267,N_3548,N_3212);
and U4268 (N_4268,N_3423,N_3634);
xnor U4269 (N_4269,N_3460,N_3380);
or U4270 (N_4270,N_3065,N_3612);
or U4271 (N_4271,N_3711,N_3693);
or U4272 (N_4272,N_3212,N_3109);
xnor U4273 (N_4273,N_3579,N_3301);
and U4274 (N_4274,N_3470,N_3259);
and U4275 (N_4275,N_3083,N_3116);
nor U4276 (N_4276,N_3304,N_3408);
or U4277 (N_4277,N_3180,N_3124);
xnor U4278 (N_4278,N_3129,N_3546);
or U4279 (N_4279,N_3031,N_3316);
and U4280 (N_4280,N_3105,N_3310);
and U4281 (N_4281,N_3057,N_3412);
or U4282 (N_4282,N_3082,N_3344);
and U4283 (N_4283,N_3707,N_3055);
xor U4284 (N_4284,N_3319,N_3436);
or U4285 (N_4285,N_3372,N_3618);
and U4286 (N_4286,N_3398,N_3629);
nand U4287 (N_4287,N_3534,N_3384);
nand U4288 (N_4288,N_3335,N_3462);
xnor U4289 (N_4289,N_3676,N_3443);
xnor U4290 (N_4290,N_3011,N_3285);
xor U4291 (N_4291,N_3226,N_3170);
nand U4292 (N_4292,N_3272,N_3622);
or U4293 (N_4293,N_3011,N_3484);
xnor U4294 (N_4294,N_3141,N_3029);
or U4295 (N_4295,N_3445,N_3317);
and U4296 (N_4296,N_3027,N_3511);
or U4297 (N_4297,N_3111,N_3321);
or U4298 (N_4298,N_3606,N_3628);
and U4299 (N_4299,N_3745,N_3193);
nor U4300 (N_4300,N_3414,N_3008);
nand U4301 (N_4301,N_3397,N_3733);
and U4302 (N_4302,N_3230,N_3373);
and U4303 (N_4303,N_3407,N_3509);
or U4304 (N_4304,N_3714,N_3705);
nand U4305 (N_4305,N_3610,N_3408);
nand U4306 (N_4306,N_3377,N_3272);
and U4307 (N_4307,N_3127,N_3429);
or U4308 (N_4308,N_3211,N_3709);
or U4309 (N_4309,N_3063,N_3246);
and U4310 (N_4310,N_3423,N_3320);
and U4311 (N_4311,N_3558,N_3168);
xor U4312 (N_4312,N_3099,N_3627);
nor U4313 (N_4313,N_3508,N_3473);
xnor U4314 (N_4314,N_3286,N_3350);
nand U4315 (N_4315,N_3579,N_3284);
xor U4316 (N_4316,N_3646,N_3696);
xor U4317 (N_4317,N_3504,N_3145);
or U4318 (N_4318,N_3598,N_3495);
nand U4319 (N_4319,N_3697,N_3400);
or U4320 (N_4320,N_3439,N_3049);
nor U4321 (N_4321,N_3627,N_3397);
or U4322 (N_4322,N_3294,N_3116);
and U4323 (N_4323,N_3717,N_3002);
nand U4324 (N_4324,N_3029,N_3354);
nand U4325 (N_4325,N_3551,N_3722);
xor U4326 (N_4326,N_3381,N_3554);
or U4327 (N_4327,N_3615,N_3522);
nand U4328 (N_4328,N_3533,N_3287);
nor U4329 (N_4329,N_3582,N_3644);
xnor U4330 (N_4330,N_3118,N_3311);
or U4331 (N_4331,N_3494,N_3653);
nand U4332 (N_4332,N_3032,N_3673);
or U4333 (N_4333,N_3543,N_3079);
nor U4334 (N_4334,N_3299,N_3617);
or U4335 (N_4335,N_3659,N_3436);
xnor U4336 (N_4336,N_3412,N_3664);
or U4337 (N_4337,N_3289,N_3325);
nor U4338 (N_4338,N_3317,N_3742);
nand U4339 (N_4339,N_3735,N_3305);
xor U4340 (N_4340,N_3274,N_3408);
and U4341 (N_4341,N_3223,N_3195);
and U4342 (N_4342,N_3038,N_3728);
or U4343 (N_4343,N_3722,N_3215);
and U4344 (N_4344,N_3273,N_3666);
and U4345 (N_4345,N_3076,N_3492);
xor U4346 (N_4346,N_3359,N_3165);
and U4347 (N_4347,N_3708,N_3110);
or U4348 (N_4348,N_3064,N_3629);
nand U4349 (N_4349,N_3399,N_3556);
or U4350 (N_4350,N_3651,N_3171);
or U4351 (N_4351,N_3349,N_3246);
or U4352 (N_4352,N_3705,N_3266);
or U4353 (N_4353,N_3009,N_3480);
and U4354 (N_4354,N_3228,N_3068);
xor U4355 (N_4355,N_3659,N_3546);
or U4356 (N_4356,N_3493,N_3531);
nand U4357 (N_4357,N_3040,N_3242);
or U4358 (N_4358,N_3031,N_3183);
and U4359 (N_4359,N_3195,N_3359);
xor U4360 (N_4360,N_3689,N_3723);
xnor U4361 (N_4361,N_3584,N_3107);
and U4362 (N_4362,N_3608,N_3102);
nor U4363 (N_4363,N_3210,N_3303);
nand U4364 (N_4364,N_3380,N_3508);
and U4365 (N_4365,N_3207,N_3462);
and U4366 (N_4366,N_3429,N_3724);
xor U4367 (N_4367,N_3745,N_3475);
or U4368 (N_4368,N_3354,N_3572);
nor U4369 (N_4369,N_3415,N_3571);
xor U4370 (N_4370,N_3369,N_3116);
and U4371 (N_4371,N_3353,N_3273);
nand U4372 (N_4372,N_3508,N_3049);
nand U4373 (N_4373,N_3324,N_3227);
nand U4374 (N_4374,N_3362,N_3336);
nand U4375 (N_4375,N_3681,N_3726);
nand U4376 (N_4376,N_3625,N_3455);
xor U4377 (N_4377,N_3668,N_3298);
nor U4378 (N_4378,N_3214,N_3301);
nand U4379 (N_4379,N_3482,N_3205);
nor U4380 (N_4380,N_3067,N_3254);
and U4381 (N_4381,N_3468,N_3520);
and U4382 (N_4382,N_3533,N_3045);
or U4383 (N_4383,N_3053,N_3743);
or U4384 (N_4384,N_3098,N_3177);
nor U4385 (N_4385,N_3311,N_3338);
and U4386 (N_4386,N_3054,N_3338);
nor U4387 (N_4387,N_3511,N_3520);
nor U4388 (N_4388,N_3227,N_3599);
nor U4389 (N_4389,N_3634,N_3160);
xnor U4390 (N_4390,N_3479,N_3195);
or U4391 (N_4391,N_3291,N_3150);
or U4392 (N_4392,N_3271,N_3668);
or U4393 (N_4393,N_3476,N_3192);
and U4394 (N_4394,N_3719,N_3357);
xnor U4395 (N_4395,N_3161,N_3439);
nand U4396 (N_4396,N_3027,N_3336);
nor U4397 (N_4397,N_3345,N_3311);
or U4398 (N_4398,N_3103,N_3229);
nand U4399 (N_4399,N_3618,N_3162);
xnor U4400 (N_4400,N_3360,N_3465);
nor U4401 (N_4401,N_3598,N_3415);
nor U4402 (N_4402,N_3530,N_3479);
xor U4403 (N_4403,N_3439,N_3132);
and U4404 (N_4404,N_3604,N_3255);
nor U4405 (N_4405,N_3443,N_3635);
nand U4406 (N_4406,N_3138,N_3184);
and U4407 (N_4407,N_3440,N_3143);
nand U4408 (N_4408,N_3704,N_3159);
and U4409 (N_4409,N_3229,N_3553);
or U4410 (N_4410,N_3477,N_3302);
and U4411 (N_4411,N_3289,N_3486);
xor U4412 (N_4412,N_3097,N_3281);
xor U4413 (N_4413,N_3011,N_3133);
nand U4414 (N_4414,N_3182,N_3379);
nand U4415 (N_4415,N_3110,N_3002);
nor U4416 (N_4416,N_3200,N_3036);
nor U4417 (N_4417,N_3117,N_3056);
xnor U4418 (N_4418,N_3464,N_3636);
nor U4419 (N_4419,N_3584,N_3365);
and U4420 (N_4420,N_3352,N_3082);
and U4421 (N_4421,N_3713,N_3016);
or U4422 (N_4422,N_3390,N_3132);
and U4423 (N_4423,N_3508,N_3343);
xnor U4424 (N_4424,N_3386,N_3325);
nand U4425 (N_4425,N_3055,N_3607);
and U4426 (N_4426,N_3404,N_3238);
nor U4427 (N_4427,N_3370,N_3330);
nand U4428 (N_4428,N_3594,N_3686);
nand U4429 (N_4429,N_3095,N_3685);
xor U4430 (N_4430,N_3344,N_3157);
or U4431 (N_4431,N_3662,N_3618);
or U4432 (N_4432,N_3670,N_3017);
or U4433 (N_4433,N_3673,N_3589);
and U4434 (N_4434,N_3708,N_3564);
xnor U4435 (N_4435,N_3553,N_3115);
xnor U4436 (N_4436,N_3615,N_3167);
xor U4437 (N_4437,N_3136,N_3060);
nand U4438 (N_4438,N_3251,N_3170);
or U4439 (N_4439,N_3294,N_3202);
or U4440 (N_4440,N_3055,N_3204);
xnor U4441 (N_4441,N_3539,N_3694);
nand U4442 (N_4442,N_3071,N_3257);
nor U4443 (N_4443,N_3551,N_3740);
nor U4444 (N_4444,N_3319,N_3363);
and U4445 (N_4445,N_3320,N_3341);
xnor U4446 (N_4446,N_3104,N_3484);
and U4447 (N_4447,N_3491,N_3444);
and U4448 (N_4448,N_3389,N_3297);
nand U4449 (N_4449,N_3302,N_3460);
nor U4450 (N_4450,N_3080,N_3435);
or U4451 (N_4451,N_3466,N_3628);
and U4452 (N_4452,N_3466,N_3680);
nor U4453 (N_4453,N_3286,N_3576);
and U4454 (N_4454,N_3242,N_3572);
or U4455 (N_4455,N_3084,N_3298);
nor U4456 (N_4456,N_3437,N_3366);
nor U4457 (N_4457,N_3275,N_3616);
nor U4458 (N_4458,N_3743,N_3376);
and U4459 (N_4459,N_3015,N_3344);
nor U4460 (N_4460,N_3368,N_3530);
nor U4461 (N_4461,N_3397,N_3629);
nor U4462 (N_4462,N_3609,N_3328);
or U4463 (N_4463,N_3225,N_3297);
and U4464 (N_4464,N_3537,N_3052);
nor U4465 (N_4465,N_3027,N_3134);
or U4466 (N_4466,N_3689,N_3012);
nand U4467 (N_4467,N_3676,N_3060);
and U4468 (N_4468,N_3262,N_3249);
xor U4469 (N_4469,N_3242,N_3146);
xnor U4470 (N_4470,N_3521,N_3579);
and U4471 (N_4471,N_3300,N_3136);
xor U4472 (N_4472,N_3609,N_3058);
or U4473 (N_4473,N_3713,N_3714);
or U4474 (N_4474,N_3533,N_3627);
and U4475 (N_4475,N_3233,N_3584);
or U4476 (N_4476,N_3023,N_3746);
nor U4477 (N_4477,N_3692,N_3353);
and U4478 (N_4478,N_3648,N_3410);
nand U4479 (N_4479,N_3415,N_3391);
xnor U4480 (N_4480,N_3176,N_3746);
nand U4481 (N_4481,N_3174,N_3016);
or U4482 (N_4482,N_3084,N_3433);
nor U4483 (N_4483,N_3583,N_3724);
nand U4484 (N_4484,N_3497,N_3474);
nor U4485 (N_4485,N_3055,N_3737);
nor U4486 (N_4486,N_3323,N_3723);
and U4487 (N_4487,N_3270,N_3039);
and U4488 (N_4488,N_3155,N_3499);
xnor U4489 (N_4489,N_3055,N_3161);
and U4490 (N_4490,N_3506,N_3701);
or U4491 (N_4491,N_3528,N_3627);
nand U4492 (N_4492,N_3012,N_3682);
and U4493 (N_4493,N_3090,N_3031);
and U4494 (N_4494,N_3650,N_3519);
nand U4495 (N_4495,N_3103,N_3172);
nor U4496 (N_4496,N_3539,N_3014);
nor U4497 (N_4497,N_3698,N_3604);
xor U4498 (N_4498,N_3017,N_3103);
and U4499 (N_4499,N_3639,N_3036);
nor U4500 (N_4500,N_4369,N_4336);
and U4501 (N_4501,N_4117,N_4448);
and U4502 (N_4502,N_3855,N_4390);
or U4503 (N_4503,N_4212,N_3889);
and U4504 (N_4504,N_4127,N_4047);
nand U4505 (N_4505,N_4303,N_3963);
nor U4506 (N_4506,N_4149,N_4193);
nor U4507 (N_4507,N_4175,N_3822);
or U4508 (N_4508,N_4292,N_3977);
or U4509 (N_4509,N_4492,N_3898);
and U4510 (N_4510,N_4133,N_3955);
xor U4511 (N_4511,N_4027,N_4194);
and U4512 (N_4512,N_4498,N_3878);
nand U4513 (N_4513,N_3958,N_3887);
nor U4514 (N_4514,N_4228,N_4024);
nand U4515 (N_4515,N_4397,N_4005);
or U4516 (N_4516,N_4355,N_3847);
xor U4517 (N_4517,N_4293,N_4053);
and U4518 (N_4518,N_4152,N_3750);
and U4519 (N_4519,N_3919,N_4497);
nor U4520 (N_4520,N_3814,N_3986);
xor U4521 (N_4521,N_3781,N_3988);
and U4522 (N_4522,N_4209,N_4368);
xor U4523 (N_4523,N_3992,N_3996);
and U4524 (N_4524,N_4314,N_4210);
xor U4525 (N_4525,N_3852,N_4002);
nor U4526 (N_4526,N_3888,N_4404);
nor U4527 (N_4527,N_4185,N_4250);
nor U4528 (N_4528,N_3901,N_4284);
and U4529 (N_4529,N_4089,N_4499);
and U4530 (N_4530,N_4331,N_4003);
nor U4531 (N_4531,N_4052,N_4470);
nand U4532 (N_4532,N_3941,N_4103);
or U4533 (N_4533,N_4416,N_3776);
xor U4534 (N_4534,N_4333,N_3985);
nor U4535 (N_4535,N_4291,N_3864);
xnor U4536 (N_4536,N_4189,N_4160);
or U4537 (N_4537,N_3960,N_4028);
or U4538 (N_4538,N_4482,N_4255);
nand U4539 (N_4539,N_4281,N_3880);
xnor U4540 (N_4540,N_3928,N_4297);
or U4541 (N_4541,N_4261,N_4258);
nand U4542 (N_4542,N_3845,N_4370);
and U4543 (N_4543,N_3990,N_3982);
xnor U4544 (N_4544,N_4231,N_4265);
nor U4545 (N_4545,N_3789,N_3956);
nor U4546 (N_4546,N_4018,N_4299);
and U4547 (N_4547,N_3932,N_3872);
nor U4548 (N_4548,N_4061,N_3907);
and U4549 (N_4549,N_4062,N_4073);
nand U4550 (N_4550,N_3821,N_3873);
nor U4551 (N_4551,N_4112,N_3858);
nand U4552 (N_4552,N_4049,N_4478);
nor U4553 (N_4553,N_3792,N_4480);
nand U4554 (N_4554,N_3800,N_4268);
or U4555 (N_4555,N_4409,N_4494);
and U4556 (N_4556,N_4392,N_3766);
nor U4557 (N_4557,N_3940,N_4318);
or U4558 (N_4558,N_4286,N_4226);
xnor U4559 (N_4559,N_3937,N_4214);
xnor U4560 (N_4560,N_3882,N_3823);
or U4561 (N_4561,N_3899,N_4420);
xnor U4562 (N_4562,N_3809,N_3819);
and U4563 (N_4563,N_4118,N_4344);
xnor U4564 (N_4564,N_4207,N_3818);
xor U4565 (N_4565,N_4432,N_3836);
xor U4566 (N_4566,N_4013,N_3862);
nand U4567 (N_4567,N_3943,N_4031);
nand U4568 (N_4568,N_4009,N_4307);
or U4569 (N_4569,N_4317,N_4245);
nand U4570 (N_4570,N_4464,N_4247);
nor U4571 (N_4571,N_3846,N_3929);
nor U4572 (N_4572,N_4223,N_3891);
xor U4573 (N_4573,N_4316,N_4056);
nor U4574 (N_4574,N_3951,N_3914);
or U4575 (N_4575,N_3912,N_4235);
nor U4576 (N_4576,N_4387,N_4034);
nand U4577 (N_4577,N_4166,N_4434);
nor U4578 (N_4578,N_4184,N_3752);
nor U4579 (N_4579,N_4467,N_4406);
nor U4580 (N_4580,N_3806,N_3810);
xnor U4581 (N_4581,N_3868,N_4290);
nand U4582 (N_4582,N_4156,N_4102);
or U4583 (N_4583,N_4086,N_4093);
or U4584 (N_4584,N_3915,N_4383);
xor U4585 (N_4585,N_4407,N_4234);
nand U4586 (N_4586,N_4094,N_4449);
and U4587 (N_4587,N_4302,N_4081);
nor U4588 (N_4588,N_4423,N_4341);
and U4589 (N_4589,N_4075,N_3867);
or U4590 (N_4590,N_3825,N_4371);
nor U4591 (N_4591,N_4058,N_4270);
or U4592 (N_4592,N_4008,N_4429);
nor U4593 (N_4593,N_4376,N_4147);
nor U4594 (N_4594,N_4378,N_4298);
and U4595 (N_4595,N_3900,N_3885);
nand U4596 (N_4596,N_3892,N_4437);
nor U4597 (N_4597,N_4114,N_4394);
and U4598 (N_4598,N_3763,N_4266);
nand U4599 (N_4599,N_4459,N_4202);
nor U4600 (N_4600,N_3859,N_3774);
and U4601 (N_4601,N_3777,N_4203);
xnor U4602 (N_4602,N_4040,N_4208);
and U4603 (N_4603,N_4195,N_3854);
or U4604 (N_4604,N_3798,N_4060);
or U4605 (N_4605,N_4413,N_3770);
and U4606 (N_4606,N_4090,N_4431);
nor U4607 (N_4607,N_4236,N_3952);
xor U4608 (N_4608,N_4155,N_4391);
xnor U4609 (N_4609,N_3906,N_4415);
xnor U4610 (N_4610,N_3861,N_4232);
and U4611 (N_4611,N_4430,N_3786);
nand U4612 (N_4612,N_3942,N_4385);
and U4613 (N_4613,N_4072,N_3771);
and U4614 (N_4614,N_4446,N_3835);
nor U4615 (N_4615,N_3920,N_3883);
and U4616 (N_4616,N_4322,N_4338);
or U4617 (N_4617,N_3933,N_4219);
nand U4618 (N_4618,N_3950,N_4453);
and U4619 (N_4619,N_4182,N_4461);
xor U4620 (N_4620,N_4486,N_4412);
and U4621 (N_4621,N_3946,N_3791);
and U4622 (N_4622,N_3954,N_4148);
nand U4623 (N_4623,N_3981,N_3830);
and U4624 (N_4624,N_4334,N_4483);
nor U4625 (N_4625,N_4411,N_4352);
nand U4626 (N_4626,N_4023,N_4457);
nor U4627 (N_4627,N_4279,N_3875);
and U4628 (N_4628,N_4248,N_3833);
or U4629 (N_4629,N_4490,N_4206);
xor U4630 (N_4630,N_4224,N_4264);
nor U4631 (N_4631,N_3793,N_4064);
nand U4632 (N_4632,N_4382,N_4039);
and U4633 (N_4633,N_4222,N_4071);
nand U4634 (N_4634,N_4309,N_4315);
nor U4635 (N_4635,N_3828,N_3790);
nor U4636 (N_4636,N_3820,N_3831);
xnor U4637 (N_4637,N_3797,N_4495);
and U4638 (N_4638,N_3799,N_4400);
nor U4639 (N_4639,N_4204,N_4289);
or U4640 (N_4640,N_4085,N_4358);
xnor U4641 (N_4641,N_4375,N_4115);
and U4642 (N_4642,N_4312,N_4433);
nor U4643 (N_4643,N_3755,N_4424);
and U4644 (N_4644,N_4259,N_3815);
or U4645 (N_4645,N_3778,N_4143);
or U4646 (N_4646,N_4421,N_4325);
and U4647 (N_4647,N_4043,N_4218);
and U4648 (N_4648,N_3964,N_4229);
nand U4649 (N_4649,N_4131,N_4273);
nand U4650 (N_4650,N_4201,N_4489);
and U4651 (N_4651,N_4109,N_3993);
nor U4652 (N_4652,N_4035,N_4374);
and U4653 (N_4653,N_4335,N_3984);
nor U4654 (N_4654,N_4138,N_4283);
nor U4655 (N_4655,N_4227,N_4068);
and U4656 (N_4656,N_3865,N_4097);
or U4657 (N_4657,N_3895,N_4256);
or U4658 (N_4658,N_4381,N_3874);
nand U4659 (N_4659,N_4340,N_4481);
and U4660 (N_4660,N_4479,N_4471);
or U4661 (N_4661,N_3921,N_3893);
and U4662 (N_4662,N_4176,N_4301);
nor U4663 (N_4663,N_4142,N_4183);
nor U4664 (N_4664,N_4139,N_4396);
or U4665 (N_4665,N_3761,N_4083);
nand U4666 (N_4666,N_4285,N_4215);
xnor U4667 (N_4667,N_4244,N_4405);
nor U4668 (N_4668,N_4393,N_3827);
nand U4669 (N_4669,N_3753,N_4168);
and U4670 (N_4670,N_4006,N_4343);
nand U4671 (N_4671,N_4124,N_4123);
and U4672 (N_4672,N_4153,N_4398);
or U4673 (N_4673,N_4144,N_4050);
nor U4674 (N_4674,N_4496,N_4472);
and U4675 (N_4675,N_4197,N_3849);
nor U4676 (N_4676,N_3866,N_4108);
nor U4677 (N_4677,N_3787,N_4037);
xor U4678 (N_4678,N_4158,N_4278);
and U4679 (N_4679,N_4036,N_4020);
nor U4680 (N_4680,N_4107,N_4087);
nor U4681 (N_4681,N_4059,N_4069);
and U4682 (N_4682,N_4096,N_3795);
xnor U4683 (N_4683,N_4065,N_4362);
xnor U4684 (N_4684,N_4414,N_4125);
nand U4685 (N_4685,N_4441,N_4187);
xnor U4686 (N_4686,N_4296,N_3812);
nor U4687 (N_4687,N_4451,N_4252);
nor U4688 (N_4688,N_3911,N_3939);
xor U4689 (N_4689,N_3876,N_4242);
nand U4690 (N_4690,N_4363,N_3877);
nand U4691 (N_4691,N_3974,N_3896);
nand U4692 (N_4692,N_4092,N_4078);
nor U4693 (N_4693,N_3968,N_3934);
and U4694 (N_4694,N_4014,N_4110);
nor U4695 (N_4695,N_4427,N_3917);
or U4696 (N_4696,N_4134,N_4001);
or U4697 (N_4697,N_4349,N_4136);
and U4698 (N_4698,N_4379,N_4051);
xnor U4699 (N_4699,N_4417,N_4044);
xnor U4700 (N_4700,N_3813,N_3913);
nor U4701 (N_4701,N_4269,N_4276);
or U4702 (N_4702,N_4326,N_4076);
nand U4703 (N_4703,N_3909,N_3935);
xnor U4704 (N_4704,N_3923,N_3775);
xor U4705 (N_4705,N_4443,N_4128);
xnor U4706 (N_4706,N_4140,N_4257);
nand U4707 (N_4707,N_3754,N_4122);
nand U4708 (N_4708,N_4100,N_4239);
or U4709 (N_4709,N_3930,N_4330);
nand U4710 (N_4710,N_3773,N_3871);
nor U4711 (N_4711,N_3837,N_4493);
and U4712 (N_4712,N_4458,N_4026);
or U4713 (N_4713,N_4473,N_4260);
and U4714 (N_4714,N_3894,N_4169);
or U4715 (N_4715,N_3785,N_3918);
nand U4716 (N_4716,N_4025,N_4254);
nor U4717 (N_4717,N_4205,N_4164);
xnor U4718 (N_4718,N_4011,N_3805);
and U4719 (N_4719,N_3824,N_3788);
nor U4720 (N_4720,N_3991,N_4384);
and U4721 (N_4721,N_4237,N_3848);
or U4722 (N_4722,N_4084,N_4113);
or U4723 (N_4723,N_4007,N_4313);
nor U4724 (N_4724,N_4141,N_3751);
nor U4725 (N_4725,N_4342,N_3969);
nor U4726 (N_4726,N_3772,N_3979);
or U4727 (N_4727,N_4196,N_4365);
and U4728 (N_4728,N_4033,N_4484);
nor U4729 (N_4729,N_4466,N_4263);
xor U4730 (N_4730,N_3784,N_4366);
xnor U4731 (N_4731,N_3860,N_3857);
nand U4732 (N_4732,N_3840,N_4332);
nand U4733 (N_4733,N_4225,N_4095);
xnor U4734 (N_4734,N_3756,N_3925);
or U4735 (N_4735,N_3948,N_4029);
or U4736 (N_4736,N_4287,N_4249);
nand U4737 (N_4737,N_3936,N_3881);
xnor U4738 (N_4738,N_3760,N_4057);
nand U4739 (N_4739,N_4462,N_4137);
or U4740 (N_4740,N_4132,N_4067);
nor U4741 (N_4741,N_4163,N_4348);
nor U4742 (N_4742,N_4399,N_4190);
nor U4743 (N_4743,N_3980,N_3832);
nor U4744 (N_4744,N_4041,N_4012);
xnor U4745 (N_4745,N_4328,N_3851);
and U4746 (N_4746,N_4386,N_4477);
nand U4747 (N_4747,N_3927,N_4488);
xnor U4748 (N_4748,N_3890,N_3801);
or U4749 (N_4749,N_4272,N_4350);
nor U4750 (N_4750,N_4380,N_4419);
xor U4751 (N_4751,N_4181,N_3966);
nor U4752 (N_4752,N_4474,N_4079);
nor U4753 (N_4753,N_4460,N_3922);
or U4754 (N_4754,N_4346,N_3869);
nor U4755 (N_4755,N_4154,N_4267);
xor U4756 (N_4756,N_4172,N_4324);
and U4757 (N_4757,N_3762,N_4487);
and U4758 (N_4758,N_3764,N_4454);
or U4759 (N_4759,N_4428,N_3886);
or U4760 (N_4760,N_4280,N_4306);
nand U4761 (N_4761,N_4357,N_4373);
nor U4762 (N_4762,N_4135,N_4162);
and U4763 (N_4763,N_4233,N_3902);
xor U4764 (N_4764,N_3816,N_4403);
nand U4765 (N_4765,N_3924,N_4251);
nor U4766 (N_4766,N_4177,N_4319);
and U4767 (N_4767,N_3998,N_3931);
nand U4768 (N_4768,N_3945,N_3961);
nand U4769 (N_4769,N_3926,N_3802);
nor U4770 (N_4770,N_4091,N_4104);
nand U4771 (N_4771,N_4356,N_4321);
nand U4772 (N_4772,N_3938,N_4145);
or U4773 (N_4773,N_3959,N_3947);
xor U4774 (N_4774,N_4116,N_3794);
or U4775 (N_4775,N_4191,N_4019);
and U4776 (N_4776,N_3970,N_4450);
or U4777 (N_4777,N_4444,N_4216);
or U4778 (N_4778,N_4361,N_4129);
xnor U4779 (N_4779,N_3903,N_3965);
and U4780 (N_4780,N_4021,N_3779);
xor U4781 (N_4781,N_3994,N_4440);
nand U4782 (N_4782,N_4401,N_4192);
xor U4783 (N_4783,N_3976,N_4485);
or U4784 (N_4784,N_4010,N_4179);
nor U4785 (N_4785,N_4074,N_3967);
and U4786 (N_4786,N_3826,N_3870);
xnor U4787 (N_4787,N_4353,N_3843);
nand U4788 (N_4788,N_4295,N_4308);
nor U4789 (N_4789,N_4238,N_3971);
and U4790 (N_4790,N_3944,N_4098);
or U4791 (N_4791,N_4300,N_3972);
xnor U4792 (N_4792,N_4159,N_4048);
nand U4793 (N_4793,N_4188,N_4046);
and U4794 (N_4794,N_4452,N_4082);
or U4795 (N_4795,N_3850,N_4294);
nand U4796 (N_4796,N_4271,N_3765);
nand U4797 (N_4797,N_4425,N_4000);
xnor U4798 (N_4798,N_3983,N_4469);
xnor U4799 (N_4799,N_4305,N_4173);
or U4800 (N_4800,N_4388,N_3973);
nor U4801 (N_4801,N_4220,N_4119);
xor U4802 (N_4802,N_4359,N_4186);
nand U4803 (N_4803,N_4422,N_3910);
or U4804 (N_4804,N_4015,N_4111);
nand U4805 (N_4805,N_4455,N_4447);
nor U4806 (N_4806,N_4161,N_4157);
or U4807 (N_4807,N_3803,N_4475);
xnor U4808 (N_4808,N_4199,N_3834);
xor U4809 (N_4809,N_4246,N_4121);
and U4810 (N_4810,N_3989,N_3796);
and U4811 (N_4811,N_3817,N_4491);
or U4812 (N_4812,N_4146,N_4004);
nand U4813 (N_4813,N_3908,N_4311);
nand U4814 (N_4814,N_4126,N_3808);
nand U4815 (N_4815,N_4288,N_4241);
xor U4816 (N_4816,N_3841,N_4174);
xnor U4817 (N_4817,N_4217,N_4274);
nor U4818 (N_4818,N_4151,N_3879);
nand U4819 (N_4819,N_3916,N_4106);
xor U4820 (N_4820,N_4468,N_3975);
or U4821 (N_4821,N_4337,N_4130);
or U4822 (N_4822,N_3757,N_3884);
or U4823 (N_4823,N_4327,N_4066);
or U4824 (N_4824,N_3838,N_4054);
xnor U4825 (N_4825,N_4347,N_4367);
nor U4826 (N_4826,N_4310,N_4070);
xnor U4827 (N_4827,N_4354,N_4055);
or U4828 (N_4828,N_3842,N_4439);
or U4829 (N_4829,N_4178,N_4389);
nor U4830 (N_4830,N_4277,N_3829);
nand U4831 (N_4831,N_3780,N_4063);
and U4832 (N_4832,N_4329,N_4213);
nand U4833 (N_4833,N_4167,N_4364);
xor U4834 (N_4834,N_4476,N_4410);
xor U4835 (N_4835,N_4320,N_3905);
nor U4836 (N_4836,N_4017,N_4211);
xnor U4837 (N_4837,N_4395,N_3987);
and U4838 (N_4838,N_4402,N_4282);
and U4839 (N_4839,N_3962,N_3999);
and U4840 (N_4840,N_3957,N_4170);
nand U4841 (N_4841,N_4171,N_4408);
nand U4842 (N_4842,N_3767,N_4120);
and U4843 (N_4843,N_3897,N_3863);
nand U4844 (N_4844,N_4032,N_3997);
xnor U4845 (N_4845,N_4101,N_4445);
nor U4846 (N_4846,N_4045,N_4088);
xnor U4847 (N_4847,N_4438,N_4198);
nand U4848 (N_4848,N_4275,N_4442);
and U4849 (N_4849,N_4230,N_3949);
xor U4850 (N_4850,N_3758,N_3978);
and U4851 (N_4851,N_3995,N_4418);
xnor U4852 (N_4852,N_4105,N_3844);
nor U4853 (N_4853,N_4077,N_3853);
nand U4854 (N_4854,N_4463,N_4372);
nor U4855 (N_4855,N_4221,N_3804);
nand U4856 (N_4856,N_4435,N_4022);
nor U4857 (N_4857,N_3839,N_4016);
nor U4858 (N_4858,N_4339,N_4304);
and U4859 (N_4859,N_4465,N_4360);
xnor U4860 (N_4860,N_4042,N_4180);
nor U4861 (N_4861,N_4243,N_3769);
or U4862 (N_4862,N_4165,N_4456);
nand U4863 (N_4863,N_3782,N_3811);
nor U4864 (N_4864,N_3783,N_4030);
nor U4865 (N_4865,N_3759,N_4377);
or U4866 (N_4866,N_3856,N_3904);
xnor U4867 (N_4867,N_3953,N_4351);
nor U4868 (N_4868,N_4080,N_4436);
nand U4869 (N_4869,N_4345,N_3807);
and U4870 (N_4870,N_4240,N_4253);
and U4871 (N_4871,N_4200,N_4323);
xnor U4872 (N_4872,N_4038,N_4099);
nor U4873 (N_4873,N_4150,N_4262);
xnor U4874 (N_4874,N_3768,N_4426);
nor U4875 (N_4875,N_4232,N_3863);
xnor U4876 (N_4876,N_4200,N_3966);
nand U4877 (N_4877,N_4191,N_4301);
nand U4878 (N_4878,N_4022,N_4185);
nor U4879 (N_4879,N_3969,N_3759);
nand U4880 (N_4880,N_3783,N_3867);
or U4881 (N_4881,N_3979,N_4005);
xor U4882 (N_4882,N_3937,N_3826);
nor U4883 (N_4883,N_4243,N_4331);
or U4884 (N_4884,N_3824,N_3922);
nor U4885 (N_4885,N_3945,N_3901);
xor U4886 (N_4886,N_3922,N_4128);
and U4887 (N_4887,N_4077,N_3789);
or U4888 (N_4888,N_3980,N_4414);
nand U4889 (N_4889,N_4177,N_3921);
and U4890 (N_4890,N_3895,N_4088);
xor U4891 (N_4891,N_4438,N_3875);
nand U4892 (N_4892,N_3905,N_4190);
nand U4893 (N_4893,N_4448,N_3890);
and U4894 (N_4894,N_4136,N_4209);
nor U4895 (N_4895,N_3867,N_3981);
nand U4896 (N_4896,N_3878,N_4156);
nand U4897 (N_4897,N_4248,N_4348);
nor U4898 (N_4898,N_4356,N_4189);
or U4899 (N_4899,N_4210,N_4469);
xor U4900 (N_4900,N_3904,N_4057);
nor U4901 (N_4901,N_4322,N_4182);
nand U4902 (N_4902,N_3916,N_4334);
nor U4903 (N_4903,N_4394,N_4473);
xnor U4904 (N_4904,N_3762,N_4140);
nor U4905 (N_4905,N_3978,N_4306);
or U4906 (N_4906,N_4464,N_4263);
nand U4907 (N_4907,N_4089,N_4068);
or U4908 (N_4908,N_4246,N_4016);
nor U4909 (N_4909,N_4286,N_3866);
nor U4910 (N_4910,N_3814,N_4170);
or U4911 (N_4911,N_4078,N_4217);
or U4912 (N_4912,N_3784,N_3845);
nor U4913 (N_4913,N_4241,N_4317);
and U4914 (N_4914,N_4412,N_4469);
or U4915 (N_4915,N_3844,N_4324);
xnor U4916 (N_4916,N_4136,N_4334);
nor U4917 (N_4917,N_4224,N_4118);
nand U4918 (N_4918,N_3816,N_3750);
nand U4919 (N_4919,N_4198,N_4429);
xor U4920 (N_4920,N_4356,N_4078);
xnor U4921 (N_4921,N_4361,N_4209);
nand U4922 (N_4922,N_4018,N_4467);
nand U4923 (N_4923,N_4441,N_3966);
xnor U4924 (N_4924,N_4100,N_3828);
and U4925 (N_4925,N_4262,N_4287);
nand U4926 (N_4926,N_3940,N_3760);
or U4927 (N_4927,N_4232,N_4194);
xor U4928 (N_4928,N_4446,N_3989);
or U4929 (N_4929,N_3859,N_4125);
nand U4930 (N_4930,N_4337,N_4389);
nand U4931 (N_4931,N_4258,N_4314);
nor U4932 (N_4932,N_4421,N_3808);
nand U4933 (N_4933,N_4147,N_4126);
nor U4934 (N_4934,N_4451,N_3894);
or U4935 (N_4935,N_3791,N_4056);
and U4936 (N_4936,N_4253,N_3965);
xor U4937 (N_4937,N_3979,N_3794);
nor U4938 (N_4938,N_4130,N_3988);
xor U4939 (N_4939,N_3939,N_4443);
nand U4940 (N_4940,N_3937,N_3775);
and U4941 (N_4941,N_4149,N_4185);
xor U4942 (N_4942,N_4221,N_4453);
and U4943 (N_4943,N_4448,N_4441);
and U4944 (N_4944,N_4138,N_3806);
nand U4945 (N_4945,N_4193,N_3869);
and U4946 (N_4946,N_4357,N_4342);
and U4947 (N_4947,N_4482,N_4476);
nand U4948 (N_4948,N_3924,N_3925);
and U4949 (N_4949,N_3799,N_3973);
nand U4950 (N_4950,N_3927,N_4463);
and U4951 (N_4951,N_4278,N_3899);
or U4952 (N_4952,N_4224,N_4091);
nand U4953 (N_4953,N_4434,N_4277);
nor U4954 (N_4954,N_3795,N_3845);
and U4955 (N_4955,N_4422,N_4437);
and U4956 (N_4956,N_4329,N_4320);
xnor U4957 (N_4957,N_3968,N_4254);
nand U4958 (N_4958,N_3979,N_4268);
and U4959 (N_4959,N_4111,N_4469);
nand U4960 (N_4960,N_3971,N_4461);
nand U4961 (N_4961,N_3926,N_4358);
and U4962 (N_4962,N_4155,N_4170);
nand U4963 (N_4963,N_4258,N_4004);
xor U4964 (N_4964,N_4478,N_4018);
and U4965 (N_4965,N_4098,N_4102);
nor U4966 (N_4966,N_4335,N_3758);
and U4967 (N_4967,N_3904,N_4202);
nor U4968 (N_4968,N_4360,N_4155);
and U4969 (N_4969,N_3790,N_4271);
and U4970 (N_4970,N_4311,N_4241);
nand U4971 (N_4971,N_4226,N_4326);
and U4972 (N_4972,N_3994,N_4460);
nand U4973 (N_4973,N_4227,N_4471);
and U4974 (N_4974,N_4416,N_4247);
and U4975 (N_4975,N_4153,N_4355);
nand U4976 (N_4976,N_4234,N_4414);
or U4977 (N_4977,N_3751,N_3869);
nand U4978 (N_4978,N_4251,N_4352);
nor U4979 (N_4979,N_4387,N_4243);
xnor U4980 (N_4980,N_4175,N_4328);
nand U4981 (N_4981,N_3991,N_3866);
xnor U4982 (N_4982,N_4028,N_4082);
nor U4983 (N_4983,N_4218,N_4109);
and U4984 (N_4984,N_4120,N_4308);
and U4985 (N_4985,N_4337,N_4046);
nor U4986 (N_4986,N_4429,N_3963);
nand U4987 (N_4987,N_4189,N_4419);
xor U4988 (N_4988,N_4487,N_3772);
nor U4989 (N_4989,N_3904,N_3962);
and U4990 (N_4990,N_4337,N_3774);
nand U4991 (N_4991,N_4200,N_4379);
and U4992 (N_4992,N_4396,N_4318);
nor U4993 (N_4993,N_4399,N_3961);
or U4994 (N_4994,N_4384,N_4264);
or U4995 (N_4995,N_3911,N_3894);
nand U4996 (N_4996,N_3961,N_3955);
nand U4997 (N_4997,N_4394,N_3933);
or U4998 (N_4998,N_3939,N_3973);
nand U4999 (N_4999,N_4023,N_4331);
nand U5000 (N_5000,N_4117,N_4143);
nor U5001 (N_5001,N_4099,N_4405);
nand U5002 (N_5002,N_4237,N_4354);
nor U5003 (N_5003,N_4479,N_4236);
or U5004 (N_5004,N_4106,N_4359);
or U5005 (N_5005,N_3847,N_4089);
nor U5006 (N_5006,N_4134,N_4075);
nor U5007 (N_5007,N_4127,N_4121);
and U5008 (N_5008,N_3914,N_4426);
nand U5009 (N_5009,N_3835,N_3870);
or U5010 (N_5010,N_4072,N_4096);
and U5011 (N_5011,N_4395,N_4488);
xor U5012 (N_5012,N_4259,N_3854);
xor U5013 (N_5013,N_4130,N_4439);
nand U5014 (N_5014,N_4008,N_3879);
or U5015 (N_5015,N_3763,N_4460);
nor U5016 (N_5016,N_4421,N_3770);
nand U5017 (N_5017,N_4367,N_4273);
nand U5018 (N_5018,N_4050,N_3756);
xnor U5019 (N_5019,N_4300,N_4073);
nor U5020 (N_5020,N_4312,N_4071);
nor U5021 (N_5021,N_4481,N_3837);
nor U5022 (N_5022,N_3930,N_4225);
nor U5023 (N_5023,N_4092,N_4440);
nor U5024 (N_5024,N_4326,N_3859);
nor U5025 (N_5025,N_3988,N_4437);
nor U5026 (N_5026,N_4229,N_4268);
and U5027 (N_5027,N_3774,N_3861);
xnor U5028 (N_5028,N_4082,N_4239);
xnor U5029 (N_5029,N_3956,N_3819);
nor U5030 (N_5030,N_4483,N_4413);
and U5031 (N_5031,N_4448,N_4246);
nor U5032 (N_5032,N_3754,N_3820);
xor U5033 (N_5033,N_4244,N_4039);
nor U5034 (N_5034,N_4478,N_4109);
or U5035 (N_5035,N_4082,N_4399);
xnor U5036 (N_5036,N_3778,N_4129);
and U5037 (N_5037,N_4054,N_4353);
or U5038 (N_5038,N_4098,N_4108);
nand U5039 (N_5039,N_4320,N_3997);
nor U5040 (N_5040,N_3785,N_3845);
xor U5041 (N_5041,N_4270,N_4242);
nor U5042 (N_5042,N_4004,N_4315);
xnor U5043 (N_5043,N_4256,N_3981);
and U5044 (N_5044,N_4320,N_3786);
nand U5045 (N_5045,N_4402,N_4108);
and U5046 (N_5046,N_4444,N_4380);
xnor U5047 (N_5047,N_4066,N_3863);
or U5048 (N_5048,N_4132,N_4095);
nand U5049 (N_5049,N_4374,N_4053);
and U5050 (N_5050,N_4069,N_4260);
nor U5051 (N_5051,N_4342,N_4168);
nor U5052 (N_5052,N_3840,N_4037);
nand U5053 (N_5053,N_4237,N_4159);
xor U5054 (N_5054,N_4288,N_4274);
xor U5055 (N_5055,N_3982,N_3946);
xnor U5056 (N_5056,N_4391,N_4036);
nor U5057 (N_5057,N_4224,N_3774);
and U5058 (N_5058,N_4093,N_3992);
nor U5059 (N_5059,N_3788,N_4475);
xnor U5060 (N_5060,N_4091,N_4026);
nor U5061 (N_5061,N_4353,N_3765);
or U5062 (N_5062,N_3969,N_3827);
and U5063 (N_5063,N_4390,N_3978);
xor U5064 (N_5064,N_4139,N_3988);
or U5065 (N_5065,N_3945,N_4176);
and U5066 (N_5066,N_4208,N_4403);
or U5067 (N_5067,N_4427,N_4105);
or U5068 (N_5068,N_4006,N_3974);
or U5069 (N_5069,N_4166,N_4051);
or U5070 (N_5070,N_4299,N_3974);
nor U5071 (N_5071,N_4359,N_4340);
and U5072 (N_5072,N_4039,N_4091);
or U5073 (N_5073,N_4261,N_4148);
nor U5074 (N_5074,N_3849,N_4432);
or U5075 (N_5075,N_4402,N_4144);
xor U5076 (N_5076,N_4405,N_4122);
xnor U5077 (N_5077,N_4020,N_4214);
xnor U5078 (N_5078,N_4156,N_4282);
or U5079 (N_5079,N_4205,N_4087);
nand U5080 (N_5080,N_4317,N_3810);
and U5081 (N_5081,N_4334,N_4455);
xor U5082 (N_5082,N_4173,N_4131);
nor U5083 (N_5083,N_4209,N_4132);
and U5084 (N_5084,N_3838,N_4324);
nand U5085 (N_5085,N_3989,N_3907);
and U5086 (N_5086,N_4376,N_4004);
and U5087 (N_5087,N_3872,N_4023);
nand U5088 (N_5088,N_3901,N_3900);
or U5089 (N_5089,N_4169,N_4476);
nor U5090 (N_5090,N_4311,N_4102);
and U5091 (N_5091,N_3929,N_3950);
and U5092 (N_5092,N_3771,N_4417);
xor U5093 (N_5093,N_4067,N_3951);
nor U5094 (N_5094,N_4255,N_4371);
nand U5095 (N_5095,N_3841,N_3844);
nand U5096 (N_5096,N_3980,N_4132);
or U5097 (N_5097,N_4059,N_4131);
nor U5098 (N_5098,N_4188,N_4038);
or U5099 (N_5099,N_3762,N_4415);
nor U5100 (N_5100,N_3964,N_4291);
nor U5101 (N_5101,N_4335,N_4089);
or U5102 (N_5102,N_4116,N_4108);
nor U5103 (N_5103,N_3766,N_4353);
or U5104 (N_5104,N_4169,N_4320);
and U5105 (N_5105,N_3950,N_4486);
xnor U5106 (N_5106,N_3873,N_3880);
and U5107 (N_5107,N_3865,N_3825);
or U5108 (N_5108,N_4350,N_4484);
xor U5109 (N_5109,N_4378,N_4135);
nor U5110 (N_5110,N_4488,N_4048);
xnor U5111 (N_5111,N_4362,N_4438);
xor U5112 (N_5112,N_3974,N_4025);
xnor U5113 (N_5113,N_3989,N_4038);
and U5114 (N_5114,N_4278,N_3938);
xnor U5115 (N_5115,N_4282,N_3991);
or U5116 (N_5116,N_4065,N_4024);
and U5117 (N_5117,N_3815,N_4456);
nor U5118 (N_5118,N_3798,N_3826);
xnor U5119 (N_5119,N_4203,N_3920);
xor U5120 (N_5120,N_4309,N_3977);
and U5121 (N_5121,N_4340,N_4318);
nor U5122 (N_5122,N_4068,N_4130);
nor U5123 (N_5123,N_4401,N_3943);
or U5124 (N_5124,N_3795,N_3848);
nor U5125 (N_5125,N_4453,N_4304);
and U5126 (N_5126,N_3980,N_4073);
or U5127 (N_5127,N_4096,N_4265);
and U5128 (N_5128,N_4090,N_4088);
and U5129 (N_5129,N_3981,N_3933);
or U5130 (N_5130,N_4059,N_3868);
xor U5131 (N_5131,N_4135,N_3789);
nand U5132 (N_5132,N_4330,N_4168);
nor U5133 (N_5133,N_4151,N_4354);
xnor U5134 (N_5134,N_4478,N_4458);
and U5135 (N_5135,N_4306,N_3766);
xor U5136 (N_5136,N_4151,N_4441);
nor U5137 (N_5137,N_3848,N_4392);
and U5138 (N_5138,N_3903,N_4455);
xnor U5139 (N_5139,N_3967,N_4053);
xnor U5140 (N_5140,N_3829,N_4099);
and U5141 (N_5141,N_3865,N_4129);
nand U5142 (N_5142,N_4251,N_4241);
nand U5143 (N_5143,N_4450,N_4201);
nor U5144 (N_5144,N_3761,N_4493);
and U5145 (N_5145,N_4328,N_4173);
or U5146 (N_5146,N_4454,N_4189);
or U5147 (N_5147,N_4275,N_4437);
nand U5148 (N_5148,N_4479,N_4308);
or U5149 (N_5149,N_4401,N_4220);
or U5150 (N_5150,N_3756,N_3770);
or U5151 (N_5151,N_4407,N_3765);
or U5152 (N_5152,N_3908,N_3936);
nand U5153 (N_5153,N_4320,N_4252);
or U5154 (N_5154,N_4075,N_4008);
nand U5155 (N_5155,N_3994,N_4022);
nor U5156 (N_5156,N_3783,N_4118);
nand U5157 (N_5157,N_4100,N_3786);
or U5158 (N_5158,N_4341,N_3899);
nor U5159 (N_5159,N_4074,N_4458);
xor U5160 (N_5160,N_4044,N_4127);
and U5161 (N_5161,N_3754,N_4178);
xor U5162 (N_5162,N_4339,N_4238);
xor U5163 (N_5163,N_3922,N_4146);
nor U5164 (N_5164,N_4346,N_3761);
nor U5165 (N_5165,N_3859,N_4230);
or U5166 (N_5166,N_4418,N_4203);
xor U5167 (N_5167,N_4016,N_3786);
and U5168 (N_5168,N_4145,N_4400);
and U5169 (N_5169,N_4248,N_3798);
nand U5170 (N_5170,N_4462,N_3762);
or U5171 (N_5171,N_4171,N_4313);
nor U5172 (N_5172,N_4415,N_4370);
nand U5173 (N_5173,N_3826,N_3785);
xnor U5174 (N_5174,N_4264,N_3949);
nand U5175 (N_5175,N_4231,N_4363);
or U5176 (N_5176,N_4118,N_4159);
or U5177 (N_5177,N_4107,N_3913);
xnor U5178 (N_5178,N_4076,N_4497);
or U5179 (N_5179,N_4049,N_4195);
nand U5180 (N_5180,N_3754,N_3868);
xnor U5181 (N_5181,N_3821,N_3965);
or U5182 (N_5182,N_4472,N_3796);
xor U5183 (N_5183,N_4151,N_3866);
nand U5184 (N_5184,N_3835,N_4360);
nand U5185 (N_5185,N_4289,N_4060);
xnor U5186 (N_5186,N_4461,N_4064);
and U5187 (N_5187,N_4019,N_4307);
xnor U5188 (N_5188,N_4430,N_3751);
or U5189 (N_5189,N_4088,N_3877);
nand U5190 (N_5190,N_4259,N_4439);
or U5191 (N_5191,N_4222,N_4240);
nand U5192 (N_5192,N_3793,N_3951);
nor U5193 (N_5193,N_3944,N_3849);
nand U5194 (N_5194,N_3945,N_4417);
or U5195 (N_5195,N_4396,N_4070);
xor U5196 (N_5196,N_3780,N_4195);
nor U5197 (N_5197,N_4144,N_4067);
or U5198 (N_5198,N_4339,N_4384);
xor U5199 (N_5199,N_4064,N_3787);
or U5200 (N_5200,N_4319,N_3830);
xor U5201 (N_5201,N_4121,N_4343);
nor U5202 (N_5202,N_4423,N_4039);
or U5203 (N_5203,N_4155,N_4241);
and U5204 (N_5204,N_4237,N_4423);
nand U5205 (N_5205,N_3969,N_3842);
or U5206 (N_5206,N_4090,N_4456);
nand U5207 (N_5207,N_4384,N_3812);
or U5208 (N_5208,N_4307,N_4121);
nor U5209 (N_5209,N_4477,N_4300);
xor U5210 (N_5210,N_4127,N_3889);
or U5211 (N_5211,N_3891,N_4492);
nor U5212 (N_5212,N_3852,N_3821);
nand U5213 (N_5213,N_3810,N_4462);
nor U5214 (N_5214,N_4442,N_4390);
nor U5215 (N_5215,N_4332,N_4137);
nand U5216 (N_5216,N_3758,N_4249);
and U5217 (N_5217,N_3821,N_4275);
and U5218 (N_5218,N_4053,N_3970);
nand U5219 (N_5219,N_4153,N_4464);
nor U5220 (N_5220,N_4366,N_3962);
xor U5221 (N_5221,N_4451,N_4357);
nand U5222 (N_5222,N_4039,N_4486);
and U5223 (N_5223,N_4234,N_4496);
and U5224 (N_5224,N_4156,N_4050);
xnor U5225 (N_5225,N_4485,N_3822);
or U5226 (N_5226,N_3832,N_4039);
nand U5227 (N_5227,N_4480,N_4322);
nand U5228 (N_5228,N_4124,N_4313);
nand U5229 (N_5229,N_3980,N_4432);
or U5230 (N_5230,N_3935,N_4432);
or U5231 (N_5231,N_3951,N_3903);
nand U5232 (N_5232,N_3807,N_4032);
xor U5233 (N_5233,N_3952,N_4260);
or U5234 (N_5234,N_4000,N_4012);
xor U5235 (N_5235,N_3792,N_3768);
nor U5236 (N_5236,N_4053,N_4331);
nand U5237 (N_5237,N_4371,N_4479);
and U5238 (N_5238,N_3920,N_3756);
or U5239 (N_5239,N_4138,N_3794);
nor U5240 (N_5240,N_4186,N_3754);
nor U5241 (N_5241,N_3758,N_4005);
nand U5242 (N_5242,N_4445,N_4374);
nand U5243 (N_5243,N_4125,N_4370);
nand U5244 (N_5244,N_3840,N_4315);
nor U5245 (N_5245,N_3921,N_4451);
or U5246 (N_5246,N_4264,N_4458);
and U5247 (N_5247,N_3897,N_3861);
nand U5248 (N_5248,N_3903,N_4327);
or U5249 (N_5249,N_4256,N_3770);
nand U5250 (N_5250,N_5207,N_4883);
nand U5251 (N_5251,N_5033,N_5082);
xnor U5252 (N_5252,N_4754,N_4742);
nor U5253 (N_5253,N_5108,N_5170);
nand U5254 (N_5254,N_4522,N_4562);
nand U5255 (N_5255,N_4857,N_4518);
nor U5256 (N_5256,N_4550,N_4700);
nor U5257 (N_5257,N_5019,N_4651);
nor U5258 (N_5258,N_4644,N_4971);
or U5259 (N_5259,N_4567,N_5162);
nor U5260 (N_5260,N_5185,N_4619);
xnor U5261 (N_5261,N_5113,N_4759);
and U5262 (N_5262,N_5102,N_5199);
and U5263 (N_5263,N_4652,N_4691);
and U5264 (N_5264,N_4991,N_5234);
nor U5265 (N_5265,N_4812,N_5178);
or U5266 (N_5266,N_4726,N_4616);
and U5267 (N_5267,N_4540,N_5213);
nor U5268 (N_5268,N_4571,N_4875);
nand U5269 (N_5269,N_4687,N_4906);
or U5270 (N_5270,N_4785,N_4859);
and U5271 (N_5271,N_5202,N_4608);
nor U5272 (N_5272,N_5134,N_4879);
or U5273 (N_5273,N_5133,N_5235);
and U5274 (N_5274,N_4880,N_4783);
and U5275 (N_5275,N_4503,N_4966);
or U5276 (N_5276,N_4814,N_4506);
nand U5277 (N_5277,N_4582,N_4909);
nor U5278 (N_5278,N_4579,N_4622);
nor U5279 (N_5279,N_4850,N_4747);
and U5280 (N_5280,N_5231,N_4639);
nand U5281 (N_5281,N_4744,N_4753);
nand U5282 (N_5282,N_4786,N_5237);
xor U5283 (N_5283,N_4757,N_4716);
and U5284 (N_5284,N_4603,N_4830);
or U5285 (N_5285,N_5059,N_4845);
xor U5286 (N_5286,N_4988,N_5174);
or U5287 (N_5287,N_5001,N_5017);
xor U5288 (N_5288,N_5192,N_4671);
or U5289 (N_5289,N_4669,N_4999);
nor U5290 (N_5290,N_4646,N_4807);
nor U5291 (N_5291,N_5233,N_4561);
and U5292 (N_5292,N_4680,N_4728);
nor U5293 (N_5293,N_4575,N_5236);
nand U5294 (N_5294,N_4730,N_4573);
xor U5295 (N_5295,N_4898,N_5000);
nor U5296 (N_5296,N_5028,N_4713);
or U5297 (N_5297,N_4678,N_4935);
or U5298 (N_5298,N_4718,N_5163);
and U5299 (N_5299,N_4572,N_4668);
nor U5300 (N_5300,N_5043,N_4596);
and U5301 (N_5301,N_4655,N_4925);
or U5302 (N_5302,N_5227,N_4665);
nor U5303 (N_5303,N_4510,N_4856);
or U5304 (N_5304,N_4722,N_5049);
or U5305 (N_5305,N_5062,N_4515);
nor U5306 (N_5306,N_5166,N_4922);
nand U5307 (N_5307,N_4610,N_4895);
or U5308 (N_5308,N_4502,N_5022);
nor U5309 (N_5309,N_4541,N_4693);
and U5310 (N_5310,N_4684,N_4926);
and U5311 (N_5311,N_4595,N_4683);
xor U5312 (N_5312,N_5140,N_5160);
and U5313 (N_5313,N_4640,N_5116);
nor U5314 (N_5314,N_5136,N_4558);
and U5315 (N_5315,N_4914,N_4873);
nand U5316 (N_5316,N_4645,N_5002);
nand U5317 (N_5317,N_4954,N_4591);
xnor U5318 (N_5318,N_4779,N_4949);
or U5319 (N_5319,N_5123,N_4772);
or U5320 (N_5320,N_4577,N_4704);
and U5321 (N_5321,N_4863,N_5040);
nand U5322 (N_5322,N_5074,N_4699);
xor U5323 (N_5323,N_5076,N_4546);
nand U5324 (N_5324,N_5183,N_5030);
xor U5325 (N_5325,N_4604,N_4794);
or U5326 (N_5326,N_4536,N_4947);
nor U5327 (N_5327,N_4968,N_4956);
and U5328 (N_5328,N_5057,N_5125);
nand U5329 (N_5329,N_5018,N_4871);
nand U5330 (N_5330,N_4686,N_4641);
and U5331 (N_5331,N_4696,N_4735);
or U5332 (N_5332,N_4594,N_5189);
nor U5333 (N_5333,N_4841,N_4874);
nor U5334 (N_5334,N_4505,N_4525);
nand U5335 (N_5335,N_5119,N_4643);
xnor U5336 (N_5336,N_4725,N_4521);
nor U5337 (N_5337,N_4962,N_4973);
nor U5338 (N_5338,N_4937,N_5181);
and U5339 (N_5339,N_5068,N_5045);
nor U5340 (N_5340,N_4948,N_5055);
nand U5341 (N_5341,N_5054,N_4840);
and U5342 (N_5342,N_4832,N_4800);
or U5343 (N_5343,N_4715,N_4995);
or U5344 (N_5344,N_5249,N_4958);
and U5345 (N_5345,N_5077,N_5099);
nor U5346 (N_5346,N_5010,N_4707);
or U5347 (N_5347,N_4679,N_5241);
and U5348 (N_5348,N_5071,N_5004);
xnor U5349 (N_5349,N_4690,N_4590);
nand U5350 (N_5350,N_4924,N_4819);
nor U5351 (N_5351,N_4854,N_4944);
and U5352 (N_5352,N_4893,N_5135);
or U5353 (N_5353,N_4959,N_4517);
and U5354 (N_5354,N_4773,N_4927);
nand U5355 (N_5355,N_4870,N_5239);
nor U5356 (N_5356,N_5215,N_4588);
nor U5357 (N_5357,N_4580,N_4852);
and U5358 (N_5358,N_4957,N_4817);
and U5359 (N_5359,N_4654,N_4533);
or U5360 (N_5360,N_5141,N_5131);
nand U5361 (N_5361,N_4771,N_4993);
nand U5362 (N_5362,N_4969,N_5031);
nor U5363 (N_5363,N_4736,N_5154);
and U5364 (N_5364,N_5095,N_4711);
nand U5365 (N_5365,N_5075,N_4630);
nor U5366 (N_5366,N_4939,N_4789);
and U5367 (N_5367,N_5220,N_5041);
and U5368 (N_5368,N_4755,N_4627);
and U5369 (N_5369,N_5006,N_4769);
xnor U5370 (N_5370,N_4501,N_5186);
and U5371 (N_5371,N_4647,N_4587);
or U5372 (N_5372,N_4770,N_5052);
or U5373 (N_5373,N_5224,N_4509);
xnor U5374 (N_5374,N_4554,N_4869);
nand U5375 (N_5375,N_4774,N_4638);
nand U5376 (N_5376,N_5219,N_5100);
xnor U5377 (N_5377,N_4945,N_5206);
or U5378 (N_5378,N_4551,N_4681);
and U5379 (N_5379,N_4581,N_4904);
nand U5380 (N_5380,N_4531,N_5156);
nand U5381 (N_5381,N_5122,N_4829);
and U5382 (N_5382,N_5021,N_4583);
xor U5383 (N_5383,N_4805,N_4825);
or U5384 (N_5384,N_4631,N_4996);
or U5385 (N_5385,N_5047,N_4853);
nor U5386 (N_5386,N_5132,N_4712);
nand U5387 (N_5387,N_4940,N_4649);
nand U5388 (N_5388,N_4598,N_4976);
and U5389 (N_5389,N_4936,N_4559);
nor U5390 (N_5390,N_5194,N_4793);
xnor U5391 (N_5391,N_5117,N_4862);
xnor U5392 (N_5392,N_4851,N_4972);
and U5393 (N_5393,N_5155,N_4806);
or U5394 (N_5394,N_4963,N_5026);
nand U5395 (N_5395,N_5078,N_4692);
and U5396 (N_5396,N_5216,N_5051);
nor U5397 (N_5397,N_5101,N_4822);
nand U5398 (N_5398,N_4612,N_4667);
nand U5399 (N_5399,N_4910,N_4877);
or U5400 (N_5400,N_4979,N_5145);
nor U5401 (N_5401,N_4565,N_4743);
or U5402 (N_5402,N_4513,N_5005);
nand U5403 (N_5403,N_4706,N_5245);
nand U5404 (N_5404,N_4688,N_4768);
nand U5405 (N_5405,N_5087,N_5009);
nor U5406 (N_5406,N_4986,N_4808);
and U5407 (N_5407,N_4983,N_4659);
nor U5408 (N_5408,N_5152,N_4710);
and U5409 (N_5409,N_4602,N_4842);
nor U5410 (N_5410,N_5190,N_5214);
nand U5411 (N_5411,N_4763,N_5247);
nor U5412 (N_5412,N_4560,N_5007);
or U5413 (N_5413,N_5187,N_5208);
or U5414 (N_5414,N_4532,N_4760);
xnor U5415 (N_5415,N_4912,N_4865);
xor U5416 (N_5416,N_5063,N_5126);
nor U5417 (N_5417,N_5015,N_4614);
xnor U5418 (N_5418,N_4574,N_4951);
or U5419 (N_5419,N_4738,N_5173);
nand U5420 (N_5420,N_4992,N_5048);
and U5421 (N_5421,N_4766,N_5105);
nor U5422 (N_5422,N_4885,N_5230);
and U5423 (N_5423,N_4504,N_5024);
nor U5424 (N_5424,N_4896,N_4508);
and U5425 (N_5425,N_4882,N_4923);
or U5426 (N_5426,N_4795,N_4682);
or U5427 (N_5427,N_5193,N_4836);
nand U5428 (N_5428,N_4750,N_4586);
or U5429 (N_5429,N_4767,N_4809);
and U5430 (N_5430,N_5085,N_5226);
or U5431 (N_5431,N_4994,N_5060);
nor U5432 (N_5432,N_4818,N_4797);
and U5433 (N_5433,N_5081,N_5203);
and U5434 (N_5434,N_5027,N_5104);
and U5435 (N_5435,N_4828,N_4975);
or U5436 (N_5436,N_4552,N_4650);
nand U5437 (N_5437,N_4867,N_5091);
xor U5438 (N_5438,N_4516,N_5147);
nand U5439 (N_5439,N_4703,N_5032);
xor U5440 (N_5440,N_4907,N_5139);
nand U5441 (N_5441,N_4601,N_5210);
and U5442 (N_5442,N_5110,N_4891);
nor U5443 (N_5443,N_5061,N_4593);
or U5444 (N_5444,N_4816,N_4843);
nand U5445 (N_5445,N_5064,N_4529);
nand U5446 (N_5446,N_4632,N_4672);
or U5447 (N_5447,N_5106,N_4765);
nor U5448 (N_5448,N_4556,N_5164);
xor U5449 (N_5449,N_4978,N_4917);
nor U5450 (N_5450,N_4666,N_4634);
nand U5451 (N_5451,N_4905,N_4899);
xnor U5452 (N_5452,N_4538,N_4539);
nand U5453 (N_5453,N_4670,N_4846);
or U5454 (N_5454,N_4844,N_4578);
or U5455 (N_5455,N_5179,N_5176);
nand U5456 (N_5456,N_5083,N_5121);
and U5457 (N_5457,N_5223,N_5103);
or U5458 (N_5458,N_4613,N_4676);
xor U5459 (N_5459,N_4911,N_4542);
or U5460 (N_5460,N_4903,N_4908);
or U5461 (N_5461,N_4511,N_4648);
xor U5462 (N_5462,N_4900,N_4952);
and U5463 (N_5463,N_4894,N_4543);
nand U5464 (N_5464,N_4702,N_4928);
nor U5465 (N_5465,N_4720,N_4860);
nand U5466 (N_5466,N_5036,N_4820);
nand U5467 (N_5467,N_4855,N_4568);
nor U5468 (N_5468,N_4620,N_5029);
nand U5469 (N_5469,N_4694,N_5070);
nor U5470 (N_5470,N_4549,N_4605);
xor U5471 (N_5471,N_4942,N_4727);
xnor U5472 (N_5472,N_5138,N_4803);
or U5473 (N_5473,N_5058,N_4987);
nor U5474 (N_5474,N_4500,N_5014);
xor U5475 (N_5475,N_5056,N_4835);
and U5476 (N_5476,N_5240,N_4555);
xnor U5477 (N_5477,N_5080,N_4915);
nor U5478 (N_5478,N_5137,N_4980);
nand U5479 (N_5479,N_4781,N_5130);
and U5480 (N_5480,N_4734,N_4848);
and U5481 (N_5481,N_5209,N_4758);
or U5482 (N_5482,N_4920,N_4790);
and U5483 (N_5483,N_5184,N_4931);
or U5484 (N_5484,N_5243,N_5034);
and U5485 (N_5485,N_5196,N_4801);
xnor U5486 (N_5486,N_4827,N_4982);
or U5487 (N_5487,N_4625,N_5109);
or U5488 (N_5488,N_4967,N_4685);
nand U5489 (N_5489,N_4823,N_4756);
or U5490 (N_5490,N_4989,N_4733);
or U5491 (N_5491,N_4752,N_4934);
and U5492 (N_5492,N_4737,N_4674);
nor U5493 (N_5493,N_4675,N_4833);
and U5494 (N_5494,N_5044,N_4938);
nor U5495 (N_5495,N_5157,N_4745);
nand U5496 (N_5496,N_5225,N_4890);
nor U5497 (N_5497,N_4761,N_5142);
xor U5498 (N_5498,N_5232,N_4545);
nand U5499 (N_5499,N_5013,N_5003);
or U5500 (N_5500,N_5107,N_4705);
and U5501 (N_5501,N_4974,N_5090);
or U5502 (N_5502,N_5198,N_4660);
nand U5503 (N_5503,N_4618,N_5180);
or U5504 (N_5504,N_4762,N_5158);
or U5505 (N_5505,N_4740,N_4837);
nor U5506 (N_5506,N_5079,N_4858);
nand U5507 (N_5507,N_4749,N_5248);
nor U5508 (N_5508,N_4732,N_4519);
and U5509 (N_5509,N_4872,N_4585);
or U5510 (N_5510,N_4941,N_4961);
and U5511 (N_5511,N_5195,N_4778);
xor U5512 (N_5512,N_4617,N_5159);
and U5513 (N_5513,N_4592,N_4788);
xor U5514 (N_5514,N_4985,N_4965);
and U5515 (N_5515,N_5144,N_5120);
nor U5516 (N_5516,N_4953,N_4698);
nor U5517 (N_5517,N_4802,N_5050);
nand U5518 (N_5518,N_5149,N_5182);
nor U5519 (N_5519,N_4597,N_5012);
nor U5520 (N_5520,N_4847,N_4977);
and U5521 (N_5521,N_4729,N_4813);
nor U5522 (N_5522,N_4723,N_4607);
nor U5523 (N_5523,N_4791,N_4964);
nand U5524 (N_5524,N_4689,N_5084);
xor U5525 (N_5525,N_5150,N_4826);
nand U5526 (N_5526,N_5042,N_5218);
or U5527 (N_5527,N_5114,N_4628);
nand U5528 (N_5528,N_4599,N_4751);
and U5529 (N_5529,N_4776,N_4623);
and U5530 (N_5530,N_5038,N_4932);
and U5531 (N_5531,N_4701,N_5171);
xor U5532 (N_5532,N_5093,N_5118);
or U5533 (N_5533,N_4714,N_5175);
or U5534 (N_5534,N_4950,N_4635);
or U5535 (N_5535,N_4537,N_4629);
nor U5536 (N_5536,N_5096,N_5200);
and U5537 (N_5537,N_4804,N_5008);
xor U5538 (N_5538,N_4955,N_4878);
and U5539 (N_5539,N_4792,N_5023);
nor U5540 (N_5540,N_5221,N_4810);
nand U5541 (N_5541,N_4798,N_4564);
xnor U5542 (N_5542,N_5072,N_5153);
xnor U5543 (N_5543,N_4748,N_4662);
or U5544 (N_5544,N_5148,N_5086);
and U5545 (N_5545,N_5112,N_5127);
xor U5546 (N_5546,N_4876,N_5217);
and U5547 (N_5547,N_4921,N_4918);
nor U5548 (N_5548,N_4764,N_4998);
xnor U5549 (N_5549,N_4520,N_4902);
xor U5550 (N_5550,N_4775,N_4849);
nand U5551 (N_5551,N_4868,N_4709);
nor U5552 (N_5552,N_5169,N_5067);
nand U5553 (N_5553,N_4930,N_4884);
xor U5554 (N_5554,N_4657,N_4615);
or U5555 (N_5555,N_5115,N_4796);
or U5556 (N_5556,N_5167,N_4563);
and U5557 (N_5557,N_5143,N_5168);
and U5558 (N_5558,N_5238,N_5092);
or U5559 (N_5559,N_4881,N_4864);
or U5560 (N_5560,N_4697,N_4782);
and U5561 (N_5561,N_4787,N_5244);
or U5562 (N_5562,N_4811,N_4784);
nand U5563 (N_5563,N_4901,N_5098);
or U5564 (N_5564,N_4717,N_5111);
nand U5565 (N_5565,N_4919,N_4527);
xor U5566 (N_5566,N_4892,N_4626);
nand U5567 (N_5567,N_5204,N_4838);
xor U5568 (N_5568,N_5229,N_4663);
nand U5569 (N_5569,N_4547,N_4741);
xor U5570 (N_5570,N_4637,N_4621);
or U5571 (N_5571,N_5124,N_5094);
nand U5572 (N_5572,N_4528,N_4570);
and U5573 (N_5573,N_4514,N_5066);
nand U5574 (N_5574,N_4523,N_5016);
nand U5575 (N_5575,N_4834,N_4724);
nor U5576 (N_5576,N_4721,N_4990);
nand U5577 (N_5577,N_4653,N_4557);
or U5578 (N_5578,N_4708,N_5037);
and U5579 (N_5579,N_4606,N_4889);
nor U5580 (N_5580,N_4600,N_4824);
and U5581 (N_5581,N_4731,N_4780);
and U5582 (N_5582,N_4677,N_5165);
xor U5583 (N_5583,N_4566,N_4661);
nand U5584 (N_5584,N_4929,N_5172);
and U5585 (N_5585,N_5188,N_5065);
and U5586 (N_5586,N_5205,N_5161);
nand U5587 (N_5587,N_5039,N_4624);
xor U5588 (N_5588,N_4960,N_4970);
nor U5589 (N_5589,N_4609,N_5246);
and U5590 (N_5590,N_5128,N_4584);
nand U5591 (N_5591,N_4739,N_4997);
or U5592 (N_5592,N_4777,N_4831);
or U5593 (N_5593,N_4887,N_4746);
xnor U5594 (N_5594,N_4576,N_4673);
nand U5595 (N_5595,N_4507,N_4642);
nand U5596 (N_5596,N_5201,N_5177);
xnor U5597 (N_5597,N_4530,N_5035);
or U5598 (N_5598,N_4861,N_4815);
xnor U5599 (N_5599,N_4821,N_4633);
nand U5600 (N_5600,N_4534,N_4946);
or U5601 (N_5601,N_4524,N_4719);
nor U5602 (N_5602,N_5073,N_5212);
nor U5603 (N_5603,N_4664,N_5211);
nor U5604 (N_5604,N_4548,N_4636);
and U5605 (N_5605,N_5197,N_5020);
or U5606 (N_5606,N_5191,N_4897);
nor U5607 (N_5607,N_4589,N_4839);
nand U5608 (N_5608,N_5222,N_4656);
and U5609 (N_5609,N_4553,N_5097);
nand U5610 (N_5610,N_5011,N_4981);
and U5611 (N_5611,N_4984,N_4886);
xor U5612 (N_5612,N_4695,N_4916);
nand U5613 (N_5613,N_4512,N_5046);
nand U5614 (N_5614,N_5129,N_4569);
nor U5615 (N_5615,N_4544,N_4799);
nor U5616 (N_5616,N_4658,N_4535);
nand U5617 (N_5617,N_4913,N_4943);
nor U5618 (N_5618,N_4888,N_5025);
or U5619 (N_5619,N_5053,N_4526);
nor U5620 (N_5620,N_5069,N_5146);
xor U5621 (N_5621,N_5089,N_5088);
and U5622 (N_5622,N_4611,N_5228);
xor U5623 (N_5623,N_5242,N_4866);
or U5624 (N_5624,N_5151,N_4933);
and U5625 (N_5625,N_5016,N_4570);
nor U5626 (N_5626,N_4529,N_5026);
and U5627 (N_5627,N_4527,N_4871);
nor U5628 (N_5628,N_5162,N_4510);
nand U5629 (N_5629,N_4996,N_4893);
or U5630 (N_5630,N_4809,N_4981);
nand U5631 (N_5631,N_4820,N_4673);
and U5632 (N_5632,N_4857,N_5013);
or U5633 (N_5633,N_5205,N_4814);
nand U5634 (N_5634,N_4901,N_5171);
or U5635 (N_5635,N_4990,N_4738);
nor U5636 (N_5636,N_4907,N_4622);
nor U5637 (N_5637,N_4629,N_4764);
or U5638 (N_5638,N_4682,N_5237);
and U5639 (N_5639,N_4931,N_4899);
or U5640 (N_5640,N_4840,N_5210);
and U5641 (N_5641,N_4725,N_4941);
nand U5642 (N_5642,N_4711,N_4621);
or U5643 (N_5643,N_5056,N_4848);
xnor U5644 (N_5644,N_5032,N_4596);
and U5645 (N_5645,N_4555,N_4685);
nand U5646 (N_5646,N_5064,N_4808);
xor U5647 (N_5647,N_4789,N_5089);
nand U5648 (N_5648,N_4512,N_4850);
nor U5649 (N_5649,N_4945,N_4507);
and U5650 (N_5650,N_4604,N_4882);
and U5651 (N_5651,N_4965,N_4974);
or U5652 (N_5652,N_5146,N_5193);
nand U5653 (N_5653,N_5189,N_4773);
nand U5654 (N_5654,N_4676,N_5157);
xnor U5655 (N_5655,N_4982,N_4612);
nor U5656 (N_5656,N_4754,N_4590);
nor U5657 (N_5657,N_4633,N_5225);
nor U5658 (N_5658,N_5094,N_4547);
nor U5659 (N_5659,N_4826,N_4707);
or U5660 (N_5660,N_5022,N_4929);
and U5661 (N_5661,N_5165,N_4958);
or U5662 (N_5662,N_4991,N_4616);
and U5663 (N_5663,N_4734,N_4565);
xor U5664 (N_5664,N_4816,N_5031);
xor U5665 (N_5665,N_4732,N_4855);
or U5666 (N_5666,N_5112,N_5217);
nand U5667 (N_5667,N_5005,N_4885);
and U5668 (N_5668,N_4780,N_4602);
or U5669 (N_5669,N_5219,N_4505);
nor U5670 (N_5670,N_4695,N_5161);
nand U5671 (N_5671,N_5122,N_5178);
and U5672 (N_5672,N_5205,N_4810);
nand U5673 (N_5673,N_4659,N_4873);
xnor U5674 (N_5674,N_5072,N_4824);
nand U5675 (N_5675,N_4703,N_4679);
xnor U5676 (N_5676,N_5082,N_4943);
or U5677 (N_5677,N_4555,N_4779);
xnor U5678 (N_5678,N_4538,N_4632);
or U5679 (N_5679,N_4604,N_4904);
or U5680 (N_5680,N_5121,N_5210);
or U5681 (N_5681,N_4595,N_4964);
or U5682 (N_5682,N_5082,N_5085);
and U5683 (N_5683,N_5086,N_5005);
xor U5684 (N_5684,N_5054,N_5188);
xor U5685 (N_5685,N_5222,N_4975);
or U5686 (N_5686,N_4880,N_4796);
or U5687 (N_5687,N_4836,N_5094);
and U5688 (N_5688,N_4793,N_4851);
xor U5689 (N_5689,N_4500,N_4684);
and U5690 (N_5690,N_4667,N_4715);
nand U5691 (N_5691,N_5031,N_4504);
or U5692 (N_5692,N_4779,N_5013);
nor U5693 (N_5693,N_5085,N_4605);
xnor U5694 (N_5694,N_5148,N_4674);
or U5695 (N_5695,N_4898,N_5037);
nand U5696 (N_5696,N_4874,N_4744);
nor U5697 (N_5697,N_5021,N_5194);
xnor U5698 (N_5698,N_4540,N_4941);
nor U5699 (N_5699,N_4619,N_4978);
nor U5700 (N_5700,N_5108,N_4892);
nor U5701 (N_5701,N_4817,N_4784);
or U5702 (N_5702,N_5081,N_4945);
and U5703 (N_5703,N_5158,N_4966);
nand U5704 (N_5704,N_5107,N_4769);
nand U5705 (N_5705,N_5136,N_4648);
and U5706 (N_5706,N_4570,N_5244);
nor U5707 (N_5707,N_5102,N_5122);
or U5708 (N_5708,N_4658,N_4712);
xnor U5709 (N_5709,N_5140,N_4588);
xnor U5710 (N_5710,N_4693,N_5074);
nand U5711 (N_5711,N_5117,N_4997);
xor U5712 (N_5712,N_5187,N_4616);
nor U5713 (N_5713,N_4960,N_4988);
or U5714 (N_5714,N_4628,N_4991);
nand U5715 (N_5715,N_4811,N_4857);
nand U5716 (N_5716,N_5160,N_5030);
xnor U5717 (N_5717,N_5172,N_5045);
or U5718 (N_5718,N_4701,N_5227);
nor U5719 (N_5719,N_4807,N_4676);
xnor U5720 (N_5720,N_5075,N_4523);
or U5721 (N_5721,N_4655,N_5244);
xor U5722 (N_5722,N_4599,N_5183);
and U5723 (N_5723,N_5150,N_4723);
nand U5724 (N_5724,N_4966,N_4926);
or U5725 (N_5725,N_4533,N_4949);
and U5726 (N_5726,N_4809,N_5044);
or U5727 (N_5727,N_4790,N_4906);
and U5728 (N_5728,N_4913,N_4910);
nand U5729 (N_5729,N_4584,N_4539);
or U5730 (N_5730,N_5189,N_5051);
or U5731 (N_5731,N_5168,N_4898);
xor U5732 (N_5732,N_5248,N_5217);
xor U5733 (N_5733,N_5097,N_4540);
nand U5734 (N_5734,N_4630,N_4617);
or U5735 (N_5735,N_4655,N_4858);
nand U5736 (N_5736,N_5103,N_5129);
and U5737 (N_5737,N_4533,N_4868);
or U5738 (N_5738,N_4933,N_4576);
and U5739 (N_5739,N_5210,N_5196);
xor U5740 (N_5740,N_4577,N_4775);
and U5741 (N_5741,N_5149,N_5082);
nor U5742 (N_5742,N_4993,N_5100);
xnor U5743 (N_5743,N_4579,N_4915);
nand U5744 (N_5744,N_5110,N_5200);
nor U5745 (N_5745,N_4591,N_4960);
nand U5746 (N_5746,N_5147,N_4902);
nor U5747 (N_5747,N_5011,N_4903);
and U5748 (N_5748,N_4927,N_5174);
xor U5749 (N_5749,N_5084,N_4918);
nand U5750 (N_5750,N_5108,N_4672);
or U5751 (N_5751,N_4842,N_4618);
xor U5752 (N_5752,N_4558,N_4646);
and U5753 (N_5753,N_4574,N_5112);
xor U5754 (N_5754,N_4918,N_4627);
nor U5755 (N_5755,N_5120,N_4677);
and U5756 (N_5756,N_4646,N_4836);
xor U5757 (N_5757,N_5044,N_4699);
or U5758 (N_5758,N_4971,N_4828);
or U5759 (N_5759,N_4601,N_5048);
xnor U5760 (N_5760,N_4576,N_4932);
xnor U5761 (N_5761,N_4621,N_4597);
xor U5762 (N_5762,N_5082,N_4509);
nor U5763 (N_5763,N_5170,N_4869);
nor U5764 (N_5764,N_5188,N_5089);
nand U5765 (N_5765,N_4647,N_5002);
nor U5766 (N_5766,N_4845,N_4830);
and U5767 (N_5767,N_4812,N_5249);
and U5768 (N_5768,N_5150,N_4722);
nand U5769 (N_5769,N_4697,N_4708);
xor U5770 (N_5770,N_5021,N_5189);
nand U5771 (N_5771,N_4946,N_4902);
or U5772 (N_5772,N_5189,N_4595);
nand U5773 (N_5773,N_4850,N_5121);
or U5774 (N_5774,N_4991,N_4795);
xnor U5775 (N_5775,N_4846,N_4941);
and U5776 (N_5776,N_4632,N_4936);
nand U5777 (N_5777,N_5023,N_4820);
nor U5778 (N_5778,N_5105,N_5011);
nor U5779 (N_5779,N_4504,N_4701);
or U5780 (N_5780,N_4750,N_5064);
nand U5781 (N_5781,N_5173,N_4864);
or U5782 (N_5782,N_4740,N_4783);
and U5783 (N_5783,N_5108,N_4545);
and U5784 (N_5784,N_4881,N_4948);
or U5785 (N_5785,N_4752,N_4655);
xnor U5786 (N_5786,N_5030,N_4825);
and U5787 (N_5787,N_4869,N_4786);
xor U5788 (N_5788,N_4681,N_5235);
or U5789 (N_5789,N_5126,N_5163);
or U5790 (N_5790,N_4999,N_5111);
nor U5791 (N_5791,N_5156,N_5099);
nor U5792 (N_5792,N_4714,N_4793);
and U5793 (N_5793,N_5121,N_4529);
xnor U5794 (N_5794,N_5040,N_5207);
nand U5795 (N_5795,N_4809,N_4909);
nor U5796 (N_5796,N_5223,N_4734);
or U5797 (N_5797,N_4936,N_5100);
and U5798 (N_5798,N_5152,N_5186);
and U5799 (N_5799,N_4932,N_5205);
nand U5800 (N_5800,N_4990,N_4982);
xor U5801 (N_5801,N_5138,N_5172);
nor U5802 (N_5802,N_4766,N_5223);
and U5803 (N_5803,N_5082,N_4584);
nand U5804 (N_5804,N_5119,N_4508);
or U5805 (N_5805,N_5061,N_4878);
xnor U5806 (N_5806,N_4747,N_4633);
and U5807 (N_5807,N_4964,N_4609);
and U5808 (N_5808,N_5130,N_4773);
or U5809 (N_5809,N_4743,N_5033);
nand U5810 (N_5810,N_5078,N_5077);
or U5811 (N_5811,N_5144,N_4754);
nor U5812 (N_5812,N_5225,N_4965);
and U5813 (N_5813,N_4545,N_4980);
and U5814 (N_5814,N_5220,N_4780);
or U5815 (N_5815,N_4804,N_4663);
and U5816 (N_5816,N_4992,N_4719);
xnor U5817 (N_5817,N_4642,N_4918);
nand U5818 (N_5818,N_4510,N_4746);
or U5819 (N_5819,N_5141,N_4549);
and U5820 (N_5820,N_4580,N_4619);
nor U5821 (N_5821,N_5143,N_5117);
xnor U5822 (N_5822,N_4941,N_4688);
and U5823 (N_5823,N_5045,N_4641);
nor U5824 (N_5824,N_4765,N_4634);
xnor U5825 (N_5825,N_4835,N_4676);
and U5826 (N_5826,N_5032,N_4511);
and U5827 (N_5827,N_4838,N_4789);
nand U5828 (N_5828,N_5158,N_4919);
nor U5829 (N_5829,N_4595,N_4587);
nor U5830 (N_5830,N_4738,N_4959);
nand U5831 (N_5831,N_4525,N_4527);
xnor U5832 (N_5832,N_4684,N_4915);
and U5833 (N_5833,N_4922,N_4667);
nand U5834 (N_5834,N_4695,N_4712);
nor U5835 (N_5835,N_4920,N_4901);
or U5836 (N_5836,N_4750,N_4864);
and U5837 (N_5837,N_4756,N_5054);
xnor U5838 (N_5838,N_5108,N_4599);
or U5839 (N_5839,N_4854,N_5127);
and U5840 (N_5840,N_4690,N_4763);
xor U5841 (N_5841,N_5104,N_4906);
nor U5842 (N_5842,N_4910,N_5070);
xnor U5843 (N_5843,N_4673,N_5111);
and U5844 (N_5844,N_4716,N_4547);
and U5845 (N_5845,N_4655,N_4820);
xor U5846 (N_5846,N_4874,N_5047);
and U5847 (N_5847,N_4869,N_5024);
nor U5848 (N_5848,N_5022,N_5142);
and U5849 (N_5849,N_4993,N_4629);
or U5850 (N_5850,N_4629,N_5228);
or U5851 (N_5851,N_4566,N_4533);
nand U5852 (N_5852,N_4838,N_5178);
xnor U5853 (N_5853,N_5164,N_4884);
and U5854 (N_5854,N_5007,N_4820);
nor U5855 (N_5855,N_4732,N_4972);
nor U5856 (N_5856,N_4538,N_4918);
and U5857 (N_5857,N_5113,N_5116);
and U5858 (N_5858,N_4888,N_4552);
nor U5859 (N_5859,N_4965,N_4907);
xnor U5860 (N_5860,N_4803,N_5158);
nand U5861 (N_5861,N_5144,N_5142);
nor U5862 (N_5862,N_4573,N_4684);
and U5863 (N_5863,N_4916,N_5068);
nor U5864 (N_5864,N_4795,N_4720);
nand U5865 (N_5865,N_4883,N_4756);
nand U5866 (N_5866,N_4793,N_4510);
nand U5867 (N_5867,N_5196,N_4908);
xor U5868 (N_5868,N_4737,N_4862);
xor U5869 (N_5869,N_4913,N_5020);
or U5870 (N_5870,N_5186,N_4970);
and U5871 (N_5871,N_5145,N_4832);
nor U5872 (N_5872,N_5189,N_4984);
xor U5873 (N_5873,N_5032,N_4650);
xnor U5874 (N_5874,N_4732,N_5046);
and U5875 (N_5875,N_4896,N_4502);
nor U5876 (N_5876,N_5176,N_5169);
and U5877 (N_5877,N_4643,N_5137);
nand U5878 (N_5878,N_4707,N_4571);
nand U5879 (N_5879,N_4668,N_4916);
or U5880 (N_5880,N_5081,N_5195);
nor U5881 (N_5881,N_5135,N_5149);
or U5882 (N_5882,N_5039,N_5220);
and U5883 (N_5883,N_4829,N_4549);
nor U5884 (N_5884,N_4738,N_4755);
or U5885 (N_5885,N_4828,N_4622);
or U5886 (N_5886,N_4818,N_4518);
nand U5887 (N_5887,N_4511,N_5020);
and U5888 (N_5888,N_4955,N_4512);
xnor U5889 (N_5889,N_5190,N_5159);
or U5890 (N_5890,N_4763,N_4999);
nand U5891 (N_5891,N_4620,N_5178);
nand U5892 (N_5892,N_5017,N_4952);
and U5893 (N_5893,N_5197,N_4965);
and U5894 (N_5894,N_4563,N_4567);
nor U5895 (N_5895,N_5193,N_5163);
and U5896 (N_5896,N_4759,N_4510);
xnor U5897 (N_5897,N_4641,N_5058);
nor U5898 (N_5898,N_5222,N_4988);
nor U5899 (N_5899,N_4712,N_5170);
nor U5900 (N_5900,N_4656,N_4635);
nor U5901 (N_5901,N_5214,N_5122);
nor U5902 (N_5902,N_5041,N_5027);
and U5903 (N_5903,N_5026,N_4942);
nand U5904 (N_5904,N_4716,N_4679);
xor U5905 (N_5905,N_5023,N_4958);
or U5906 (N_5906,N_4671,N_5030);
nor U5907 (N_5907,N_4660,N_5232);
and U5908 (N_5908,N_5097,N_4933);
nand U5909 (N_5909,N_5210,N_4714);
or U5910 (N_5910,N_4963,N_4624);
nor U5911 (N_5911,N_5046,N_5237);
xor U5912 (N_5912,N_4728,N_5198);
or U5913 (N_5913,N_5058,N_4517);
nor U5914 (N_5914,N_5065,N_4542);
nor U5915 (N_5915,N_5089,N_4838);
nand U5916 (N_5916,N_4867,N_4899);
xnor U5917 (N_5917,N_5137,N_5134);
and U5918 (N_5918,N_5095,N_5105);
or U5919 (N_5919,N_4600,N_5059);
xor U5920 (N_5920,N_5175,N_5164);
xnor U5921 (N_5921,N_4990,N_4937);
xor U5922 (N_5922,N_5030,N_4965);
nand U5923 (N_5923,N_5103,N_5219);
nand U5924 (N_5924,N_4977,N_5059);
or U5925 (N_5925,N_4945,N_5005);
nand U5926 (N_5926,N_4587,N_4942);
or U5927 (N_5927,N_5132,N_5072);
xor U5928 (N_5928,N_4767,N_4536);
nand U5929 (N_5929,N_5243,N_4536);
xor U5930 (N_5930,N_4770,N_5023);
nand U5931 (N_5931,N_4931,N_4716);
and U5932 (N_5932,N_4736,N_4592);
nand U5933 (N_5933,N_4816,N_4852);
nand U5934 (N_5934,N_4607,N_4988);
and U5935 (N_5935,N_4756,N_4853);
xnor U5936 (N_5936,N_4726,N_5137);
and U5937 (N_5937,N_4863,N_4762);
nor U5938 (N_5938,N_4886,N_4991);
or U5939 (N_5939,N_4551,N_4533);
or U5940 (N_5940,N_4890,N_4549);
and U5941 (N_5941,N_5137,N_4841);
and U5942 (N_5942,N_4950,N_4609);
xor U5943 (N_5943,N_4620,N_5233);
and U5944 (N_5944,N_5003,N_5148);
nor U5945 (N_5945,N_5052,N_4993);
or U5946 (N_5946,N_5107,N_5212);
nor U5947 (N_5947,N_5125,N_4852);
or U5948 (N_5948,N_5131,N_4888);
or U5949 (N_5949,N_4646,N_4913);
and U5950 (N_5950,N_4750,N_5088);
or U5951 (N_5951,N_4994,N_4650);
nor U5952 (N_5952,N_5124,N_5036);
nand U5953 (N_5953,N_4540,N_4828);
or U5954 (N_5954,N_4902,N_4687);
nor U5955 (N_5955,N_4912,N_5231);
xor U5956 (N_5956,N_5186,N_4527);
or U5957 (N_5957,N_4771,N_4551);
and U5958 (N_5958,N_5086,N_4635);
nand U5959 (N_5959,N_5121,N_5221);
nand U5960 (N_5960,N_4518,N_5154);
and U5961 (N_5961,N_4904,N_5141);
nand U5962 (N_5962,N_4591,N_5147);
nor U5963 (N_5963,N_5036,N_5244);
and U5964 (N_5964,N_4803,N_4629);
xor U5965 (N_5965,N_4891,N_5034);
xnor U5966 (N_5966,N_4717,N_4718);
nor U5967 (N_5967,N_4714,N_4871);
nor U5968 (N_5968,N_4972,N_5068);
and U5969 (N_5969,N_5019,N_5048);
or U5970 (N_5970,N_4785,N_4610);
and U5971 (N_5971,N_5025,N_4720);
or U5972 (N_5972,N_4718,N_5016);
nand U5973 (N_5973,N_4620,N_4831);
or U5974 (N_5974,N_4515,N_4718);
nor U5975 (N_5975,N_5031,N_4565);
xor U5976 (N_5976,N_5224,N_4871);
xor U5977 (N_5977,N_5013,N_5058);
or U5978 (N_5978,N_5218,N_5101);
and U5979 (N_5979,N_5158,N_4952);
or U5980 (N_5980,N_4740,N_4878);
nand U5981 (N_5981,N_4800,N_4790);
or U5982 (N_5982,N_4519,N_4913);
and U5983 (N_5983,N_4806,N_5093);
xnor U5984 (N_5984,N_5102,N_5157);
nor U5985 (N_5985,N_4953,N_5189);
xnor U5986 (N_5986,N_4647,N_4713);
nand U5987 (N_5987,N_4917,N_5215);
xnor U5988 (N_5988,N_5017,N_5210);
nor U5989 (N_5989,N_5005,N_5207);
or U5990 (N_5990,N_5162,N_4683);
or U5991 (N_5991,N_4742,N_4794);
or U5992 (N_5992,N_4530,N_5095);
or U5993 (N_5993,N_5230,N_5233);
nand U5994 (N_5994,N_5017,N_5011);
xor U5995 (N_5995,N_5219,N_4923);
and U5996 (N_5996,N_4627,N_4702);
or U5997 (N_5997,N_5083,N_4943);
or U5998 (N_5998,N_4927,N_4829);
xnor U5999 (N_5999,N_5103,N_4667);
xor U6000 (N_6000,N_5319,N_5369);
and U6001 (N_6001,N_5255,N_5742);
or U6002 (N_6002,N_5648,N_5499);
xnor U6003 (N_6003,N_5437,N_5746);
and U6004 (N_6004,N_5630,N_5681);
and U6005 (N_6005,N_5784,N_5416);
or U6006 (N_6006,N_5414,N_5675);
xnor U6007 (N_6007,N_5881,N_5834);
and U6008 (N_6008,N_5374,N_5388);
or U6009 (N_6009,N_5835,N_5649);
or U6010 (N_6010,N_5712,N_5926);
or U6011 (N_6011,N_5811,N_5729);
and U6012 (N_6012,N_5776,N_5673);
or U6013 (N_6013,N_5798,N_5534);
xor U6014 (N_6014,N_5274,N_5686);
or U6015 (N_6015,N_5262,N_5544);
and U6016 (N_6016,N_5528,N_5423);
and U6017 (N_6017,N_5894,N_5480);
nor U6018 (N_6018,N_5945,N_5833);
nor U6019 (N_6019,N_5713,N_5587);
nand U6020 (N_6020,N_5783,N_5396);
and U6021 (N_6021,N_5638,N_5506);
or U6022 (N_6022,N_5925,N_5965);
and U6023 (N_6023,N_5955,N_5984);
and U6024 (N_6024,N_5782,N_5699);
xnor U6025 (N_6025,N_5564,N_5901);
nand U6026 (N_6026,N_5879,N_5560);
nand U6027 (N_6027,N_5357,N_5330);
and U6028 (N_6028,N_5379,N_5496);
or U6029 (N_6029,N_5359,N_5497);
or U6030 (N_6030,N_5584,N_5820);
and U6031 (N_6031,N_5709,N_5943);
or U6032 (N_6032,N_5823,N_5424);
xor U6033 (N_6033,N_5633,N_5324);
xnor U6034 (N_6034,N_5458,N_5483);
and U6035 (N_6035,N_5973,N_5397);
xnor U6036 (N_6036,N_5794,N_5860);
nor U6037 (N_6037,N_5609,N_5615);
nor U6038 (N_6038,N_5356,N_5789);
or U6039 (N_6039,N_5949,N_5484);
xnor U6040 (N_6040,N_5392,N_5705);
nand U6041 (N_6041,N_5663,N_5460);
or U6042 (N_6042,N_5567,N_5991);
and U6043 (N_6043,N_5632,N_5969);
xnor U6044 (N_6044,N_5736,N_5817);
or U6045 (N_6045,N_5352,N_5399);
nand U6046 (N_6046,N_5909,N_5539);
nor U6047 (N_6047,N_5536,N_5850);
and U6048 (N_6048,N_5815,N_5596);
xor U6049 (N_6049,N_5474,N_5853);
nor U6050 (N_6050,N_5692,N_5915);
xnor U6051 (N_6051,N_5889,N_5689);
nor U6052 (N_6052,N_5337,N_5515);
xnor U6053 (N_6053,N_5895,N_5946);
and U6054 (N_6054,N_5660,N_5407);
or U6055 (N_6055,N_5883,N_5293);
nor U6056 (N_6056,N_5252,N_5309);
nand U6057 (N_6057,N_5842,N_5321);
nand U6058 (N_6058,N_5655,N_5888);
nand U6059 (N_6059,N_5934,N_5808);
or U6060 (N_6060,N_5485,N_5737);
or U6061 (N_6061,N_5482,N_5758);
nor U6062 (N_6062,N_5932,N_5754);
or U6063 (N_6063,N_5862,N_5875);
or U6064 (N_6064,N_5780,N_5401);
xor U6065 (N_6065,N_5521,N_5732);
nor U6066 (N_6066,N_5626,N_5781);
xnor U6067 (N_6067,N_5362,N_5948);
or U6068 (N_6068,N_5791,N_5899);
or U6069 (N_6069,N_5579,N_5266);
and U6070 (N_6070,N_5878,N_5297);
and U6071 (N_6071,N_5923,N_5511);
or U6072 (N_6072,N_5777,N_5939);
or U6073 (N_6073,N_5565,N_5719);
and U6074 (N_6074,N_5577,N_5892);
and U6075 (N_6075,N_5828,N_5523);
or U6076 (N_6076,N_5725,N_5857);
or U6077 (N_6077,N_5877,N_5957);
xnor U6078 (N_6078,N_5900,N_5651);
xor U6079 (N_6079,N_5890,N_5639);
or U6080 (N_6080,N_5708,N_5300);
nand U6081 (N_6081,N_5740,N_5277);
nand U6082 (N_6082,N_5674,N_5507);
nor U6083 (N_6083,N_5322,N_5592);
xnor U6084 (N_6084,N_5345,N_5287);
nand U6085 (N_6085,N_5799,N_5967);
or U6086 (N_6086,N_5332,N_5444);
or U6087 (N_6087,N_5625,N_5690);
xnor U6088 (N_6088,N_5411,N_5911);
nor U6089 (N_6089,N_5617,N_5271);
nor U6090 (N_6090,N_5968,N_5349);
or U6091 (N_6091,N_5624,N_5953);
nor U6092 (N_6092,N_5541,N_5306);
nand U6093 (N_6093,N_5279,N_5514);
or U6094 (N_6094,N_5961,N_5433);
nor U6095 (N_6095,N_5779,N_5537);
or U6096 (N_6096,N_5825,N_5263);
and U6097 (N_6097,N_5555,N_5446);
nor U6098 (N_6098,N_5891,N_5886);
or U6099 (N_6099,N_5364,N_5677);
nand U6100 (N_6100,N_5477,N_5488);
and U6101 (N_6101,N_5752,N_5320);
nand U6102 (N_6102,N_5302,N_5270);
nor U6103 (N_6103,N_5786,N_5504);
and U6104 (N_6104,N_5486,N_5492);
nor U6105 (N_6105,N_5576,N_5329);
nor U6106 (N_6106,N_5475,N_5394);
or U6107 (N_6107,N_5865,N_5600);
nand U6108 (N_6108,N_5990,N_5869);
and U6109 (N_6109,N_5972,N_5513);
nor U6110 (N_6110,N_5696,N_5643);
xnor U6111 (N_6111,N_5261,N_5406);
or U6112 (N_6112,N_5734,N_5680);
xor U6113 (N_6113,N_5771,N_5415);
nand U6114 (N_6114,N_5461,N_5882);
or U6115 (N_6115,N_5658,N_5826);
nor U6116 (N_6116,N_5375,N_5597);
nand U6117 (N_6117,N_5743,N_5710);
xor U6118 (N_6118,N_5750,N_5970);
nand U6119 (N_6119,N_5898,N_5435);
or U6120 (N_6120,N_5269,N_5525);
nor U6121 (N_6121,N_5520,N_5256);
or U6122 (N_6122,N_5652,N_5490);
or U6123 (N_6123,N_5467,N_5501);
or U6124 (N_6124,N_5298,N_5769);
nand U6125 (N_6125,N_5347,N_5304);
nor U6126 (N_6126,N_5518,N_5914);
nor U6127 (N_6127,N_5805,N_5383);
nor U6128 (N_6128,N_5334,N_5545);
xor U6129 (N_6129,N_5569,N_5711);
nor U6130 (N_6130,N_5801,N_5589);
xor U6131 (N_6131,N_5454,N_5735);
nand U6132 (N_6132,N_5373,N_5434);
or U6133 (N_6133,N_5519,N_5682);
nand U6134 (N_6134,N_5595,N_5469);
nand U6135 (N_6135,N_5951,N_5532);
nor U6136 (N_6136,N_5818,N_5568);
nor U6137 (N_6137,N_5289,N_5348);
or U6138 (N_6138,N_5547,N_5714);
and U6139 (N_6139,N_5331,N_5494);
nand U6140 (N_6140,N_5463,N_5893);
and U6141 (N_6141,N_5453,N_5402);
nor U6142 (N_6142,N_5275,N_5549);
xnor U6143 (N_6143,N_5295,N_5870);
nand U6144 (N_6144,N_5761,N_5646);
nand U6145 (N_6145,N_5614,N_5429);
or U6146 (N_6146,N_5420,N_5443);
nand U6147 (N_6147,N_5941,N_5913);
xnor U6148 (N_6148,N_5728,N_5802);
or U6149 (N_6149,N_5940,N_5887);
and U6150 (N_6150,N_5693,N_5384);
xor U6151 (N_6151,N_5822,N_5809);
xnor U6152 (N_6152,N_5753,N_5723);
and U6153 (N_6153,N_5366,N_5880);
or U6154 (N_6154,N_5276,N_5668);
nor U6155 (N_6155,N_5785,N_5398);
and U6156 (N_6156,N_5744,N_5325);
xor U6157 (N_6157,N_5981,N_5773);
and U6158 (N_6158,N_5363,N_5989);
or U6159 (N_6159,N_5721,N_5351);
and U6160 (N_6160,N_5790,N_5258);
nor U6161 (N_6161,N_5422,N_5376);
and U6162 (N_6162,N_5472,N_5290);
or U6163 (N_6163,N_5389,N_5727);
xnor U6164 (N_6164,N_5959,N_5730);
nand U6165 (N_6165,N_5907,N_5253);
nand U6166 (N_6166,N_5535,N_5999);
or U6167 (N_6167,N_5487,N_5573);
nor U6168 (N_6168,N_5816,N_5640);
and U6169 (N_6169,N_5694,N_5338);
or U6170 (N_6170,N_5554,N_5748);
nor U6171 (N_6171,N_5938,N_5430);
xor U6172 (N_6172,N_5698,N_5585);
or U6173 (N_6173,N_5529,N_5910);
nand U6174 (N_6174,N_5599,N_5548);
nand U6175 (N_6175,N_5839,N_5508);
or U6176 (N_6176,N_5662,N_5350);
or U6177 (N_6177,N_5985,N_5629);
nor U6178 (N_6178,N_5647,N_5718);
and U6179 (N_6179,N_5944,N_5905);
xnor U6180 (N_6180,N_5272,N_5445);
and U6181 (N_6181,N_5966,N_5608);
or U6182 (N_6182,N_5566,N_5700);
nand U6183 (N_6183,N_5716,N_5788);
and U6184 (N_6184,N_5301,N_5512);
xor U6185 (N_6185,N_5903,N_5264);
xor U6186 (N_6186,N_5294,N_5653);
or U6187 (N_6187,N_5847,N_5841);
and U6188 (N_6188,N_5303,N_5755);
nand U6189 (N_6189,N_5361,N_5971);
and U6190 (N_6190,N_5912,N_5412);
nand U6191 (N_6191,N_5558,N_5308);
and U6192 (N_6192,N_5333,N_5542);
and U6193 (N_6193,N_5387,N_5343);
xnor U6194 (N_6194,N_5311,N_5747);
xor U6195 (N_6195,N_5456,N_5618);
or U6196 (N_6196,N_5533,N_5421);
and U6197 (N_6197,N_5503,N_5390);
xor U6198 (N_6198,N_5678,N_5977);
and U6199 (N_6199,N_5688,N_5468);
nand U6200 (N_6200,N_5960,N_5738);
nand U6201 (N_6201,N_5621,N_5278);
nand U6202 (N_6202,N_5635,N_5667);
nand U6203 (N_6203,N_5676,N_5449);
nor U6204 (N_6204,N_5336,N_5268);
or U6205 (N_6205,N_5543,N_5495);
xor U6206 (N_6206,N_5593,N_5812);
xnor U6207 (N_6207,N_5381,N_5551);
nor U6208 (N_6208,N_5843,N_5836);
xor U6209 (N_6209,N_5760,N_5344);
nor U6210 (N_6210,N_5382,N_5832);
nor U6211 (N_6211,N_5958,N_5522);
and U6212 (N_6212,N_5282,N_5413);
or U6213 (N_6213,N_5284,N_5904);
or U6214 (N_6214,N_5530,N_5764);
and U6215 (N_6215,N_5774,N_5441);
and U6216 (N_6216,N_5385,N_5642);
xor U6217 (N_6217,N_5697,N_5299);
or U6218 (N_6218,N_5286,N_5792);
nor U6219 (N_6219,N_5556,N_5603);
nand U6220 (N_6220,N_5408,N_5393);
nand U6221 (N_6221,N_5918,N_5419);
nor U6222 (N_6222,N_5706,N_5717);
or U6223 (N_6223,N_5315,N_5296);
and U6224 (N_6224,N_5645,N_5813);
xnor U6225 (N_6225,N_5563,N_5447);
nor U6226 (N_6226,N_5502,N_5858);
and U6227 (N_6227,N_5583,N_5620);
xor U6228 (N_6228,N_5341,N_5720);
nor U6229 (N_6229,N_5722,N_5606);
and U6230 (N_6230,N_5531,N_5627);
nand U6231 (N_6231,N_5561,N_5980);
or U6232 (N_6232,N_5749,N_5745);
nand U6233 (N_6233,N_5580,N_5793);
xnor U6234 (N_6234,N_5864,N_5993);
xor U6235 (N_6235,N_5481,N_5634);
nor U6236 (N_6236,N_5616,N_5427);
and U6237 (N_6237,N_5679,N_5669);
nor U6238 (N_6238,N_5613,N_5251);
xor U6239 (N_6239,N_5281,N_5465);
xnor U6240 (N_6240,N_5637,N_5259);
nand U6241 (N_6241,N_5916,N_5707);
nor U6242 (N_6242,N_5470,N_5292);
xnor U6243 (N_6243,N_5378,N_5605);
or U6244 (N_6244,N_5731,N_5317);
or U6245 (N_6245,N_5767,N_5510);
nand U6246 (N_6246,N_5810,N_5756);
nand U6247 (N_6247,N_5715,N_5450);
and U6248 (N_6248,N_5974,N_5775);
nor U6249 (N_6249,N_5623,N_5628);
nand U6250 (N_6250,N_5619,N_5844);
nand U6251 (N_6251,N_5814,N_5952);
nand U6252 (N_6252,N_5265,N_5254);
nor U6253 (N_6253,N_5260,N_5803);
nor U6254 (N_6254,N_5919,N_5305);
xnor U6255 (N_6255,N_5500,N_5804);
xnor U6256 (N_6256,N_5695,N_5762);
nand U6257 (N_6257,N_5931,N_5867);
or U6258 (N_6258,N_5451,N_5326);
nand U6259 (N_6259,N_5838,N_5661);
or U6260 (N_6260,N_5796,N_5982);
and U6261 (N_6261,N_5346,N_5726);
nand U6262 (N_6262,N_5307,N_5439);
nand U6263 (N_6263,N_5975,N_5751);
nand U6264 (N_6264,N_5795,N_5436);
nand U6265 (N_6265,N_5610,N_5310);
nand U6266 (N_6266,N_5612,N_5996);
nand U6267 (N_6267,N_5868,N_5340);
nand U6268 (N_6268,N_5323,N_5409);
nor U6269 (N_6269,N_5312,N_5733);
nor U6270 (N_6270,N_5848,N_5947);
or U6271 (N_6271,N_5489,N_5691);
or U6272 (N_6272,N_5493,N_5950);
nor U6273 (N_6273,N_5866,N_5906);
nor U6274 (N_6274,N_5840,N_5942);
nor U6275 (N_6275,N_5557,N_5425);
nor U6276 (N_6276,N_5759,N_5354);
or U6277 (N_6277,N_5594,N_5983);
and U6278 (N_6278,N_5462,N_5819);
or U6279 (N_6279,N_5358,N_5778);
and U6280 (N_6280,N_5391,N_5377);
and U6281 (N_6281,N_5978,N_5831);
or U6282 (N_6282,N_5591,N_5659);
and U6283 (N_6283,N_5479,N_5273);
nand U6284 (N_6284,N_5863,N_5902);
xnor U6285 (N_6285,N_5559,N_5871);
xor U6286 (N_6286,N_5601,N_5355);
nand U6287 (N_6287,N_5339,N_5267);
and U6288 (N_6288,N_5920,N_5448);
xor U6289 (N_6289,N_5874,N_5371);
nor U6290 (N_6290,N_5859,N_5464);
nor U6291 (N_6291,N_5403,N_5829);
xor U6292 (N_6292,N_5852,N_5426);
xor U6293 (N_6293,N_5405,N_5765);
and U6294 (N_6294,N_5553,N_5763);
nor U6295 (N_6295,N_5517,N_5672);
or U6296 (N_6296,N_5739,N_5417);
or U6297 (N_6297,N_5861,N_5571);
or U6298 (N_6298,N_5575,N_5665);
and U6299 (N_6299,N_5928,N_5428);
nand U6300 (N_6300,N_5431,N_5849);
nor U6301 (N_6301,N_5636,N_5288);
or U6302 (N_6302,N_5526,N_5703);
or U6303 (N_6303,N_5418,N_5884);
nand U6304 (N_6304,N_5400,N_5581);
nor U6305 (N_6305,N_5478,N_5318);
nor U6306 (N_6306,N_5438,N_5671);
nand U6307 (N_6307,N_5574,N_5768);
or U6308 (N_6308,N_5684,N_5590);
nand U6309 (N_6309,N_5922,N_5466);
nor U6310 (N_6310,N_5562,N_5685);
and U6311 (N_6311,N_5876,N_5550);
xnor U6312 (N_6312,N_5367,N_5963);
or U6313 (N_6313,N_5937,N_5365);
and U6314 (N_6314,N_5524,N_5654);
nand U6315 (N_6315,N_5787,N_5995);
and U6316 (N_6316,N_5250,N_5757);
xor U6317 (N_6317,N_5410,N_5578);
or U6318 (N_6318,N_5724,N_5602);
nor U6319 (N_6319,N_5687,N_5452);
xnor U6320 (N_6320,N_5540,N_5442);
or U6321 (N_6321,N_5285,N_5992);
nor U6322 (N_6322,N_5806,N_5935);
nand U6323 (N_6323,N_5824,N_5770);
nand U6324 (N_6324,N_5459,N_5921);
nand U6325 (N_6325,N_5586,N_5473);
and U6326 (N_6326,N_5631,N_5664);
xnor U6327 (N_6327,N_5516,N_5854);
or U6328 (N_6328,N_5986,N_5316);
and U6329 (N_6329,N_5701,N_5476);
xor U6330 (N_6330,N_5872,N_5598);
nor U6331 (N_6331,N_5704,N_5327);
xnor U6332 (N_6332,N_5670,N_5650);
nor U6333 (N_6333,N_5837,N_5588);
nand U6334 (N_6334,N_5976,N_5611);
xnor U6335 (N_6335,N_5370,N_5582);
and U6336 (N_6336,N_5933,N_5845);
nand U6337 (N_6337,N_5457,N_5641);
and U6338 (N_6338,N_5741,N_5505);
nor U6339 (N_6339,N_5360,N_5929);
xor U6340 (N_6340,N_5395,N_5908);
xor U6341 (N_6341,N_5821,N_5924);
or U6342 (N_6342,N_5604,N_5280);
nor U6343 (N_6343,N_5807,N_5353);
or U6344 (N_6344,N_5997,N_5314);
or U6345 (N_6345,N_5440,N_5498);
nor U6346 (N_6346,N_5546,N_5856);
and U6347 (N_6347,N_5335,N_5855);
nand U6348 (N_6348,N_5607,N_5800);
xor U6349 (N_6349,N_5917,N_5386);
nand U6350 (N_6350,N_5994,N_5873);
nand U6351 (N_6351,N_5987,N_5851);
or U6352 (N_6352,N_5432,N_5372);
and U6353 (N_6353,N_5527,N_5827);
and U6354 (N_6354,N_5657,N_5656);
xor U6355 (N_6355,N_5702,N_5552);
xor U6356 (N_6356,N_5936,N_5885);
and U6357 (N_6357,N_5998,N_5283);
nand U6358 (N_6358,N_5257,N_5979);
or U6359 (N_6359,N_5830,N_5954);
nor U6360 (N_6360,N_5291,N_5368);
or U6361 (N_6361,N_5930,N_5964);
nor U6362 (N_6362,N_5455,N_5683);
nor U6363 (N_6363,N_5538,N_5313);
xnor U6364 (N_6364,N_5570,N_5846);
nor U6365 (N_6365,N_5896,N_5797);
nor U6366 (N_6366,N_5927,N_5491);
nor U6367 (N_6367,N_5404,N_5772);
nor U6368 (N_6368,N_5509,N_5644);
nor U6369 (N_6369,N_5622,N_5988);
xnor U6370 (N_6370,N_5897,N_5962);
xnor U6371 (N_6371,N_5380,N_5342);
nand U6372 (N_6372,N_5956,N_5572);
nor U6373 (N_6373,N_5666,N_5328);
nor U6374 (N_6374,N_5766,N_5471);
xor U6375 (N_6375,N_5938,N_5567);
nand U6376 (N_6376,N_5364,N_5960);
nor U6377 (N_6377,N_5316,N_5500);
xor U6378 (N_6378,N_5679,N_5273);
and U6379 (N_6379,N_5267,N_5867);
nand U6380 (N_6380,N_5676,N_5297);
or U6381 (N_6381,N_5914,N_5778);
and U6382 (N_6382,N_5722,N_5729);
or U6383 (N_6383,N_5871,N_5519);
nor U6384 (N_6384,N_5915,N_5746);
nand U6385 (N_6385,N_5679,N_5341);
and U6386 (N_6386,N_5847,N_5862);
or U6387 (N_6387,N_5433,N_5298);
nand U6388 (N_6388,N_5508,N_5754);
xor U6389 (N_6389,N_5341,N_5538);
or U6390 (N_6390,N_5482,N_5475);
xor U6391 (N_6391,N_5295,N_5261);
or U6392 (N_6392,N_5521,N_5580);
and U6393 (N_6393,N_5612,N_5508);
and U6394 (N_6394,N_5274,N_5370);
nor U6395 (N_6395,N_5437,N_5928);
nand U6396 (N_6396,N_5712,N_5715);
nand U6397 (N_6397,N_5665,N_5359);
or U6398 (N_6398,N_5849,N_5570);
xnor U6399 (N_6399,N_5621,N_5397);
xnor U6400 (N_6400,N_5839,N_5491);
nand U6401 (N_6401,N_5749,N_5460);
or U6402 (N_6402,N_5314,N_5484);
or U6403 (N_6403,N_5308,N_5937);
nor U6404 (N_6404,N_5449,N_5923);
nor U6405 (N_6405,N_5324,N_5941);
or U6406 (N_6406,N_5533,N_5462);
nor U6407 (N_6407,N_5933,N_5769);
or U6408 (N_6408,N_5853,N_5550);
nand U6409 (N_6409,N_5817,N_5603);
nand U6410 (N_6410,N_5933,N_5740);
nor U6411 (N_6411,N_5539,N_5703);
or U6412 (N_6412,N_5919,N_5526);
nand U6413 (N_6413,N_5800,N_5924);
or U6414 (N_6414,N_5974,N_5825);
nand U6415 (N_6415,N_5427,N_5334);
or U6416 (N_6416,N_5491,N_5320);
and U6417 (N_6417,N_5643,N_5867);
and U6418 (N_6418,N_5343,N_5686);
or U6419 (N_6419,N_5849,N_5691);
or U6420 (N_6420,N_5266,N_5624);
xnor U6421 (N_6421,N_5531,N_5847);
and U6422 (N_6422,N_5743,N_5484);
xnor U6423 (N_6423,N_5756,N_5906);
nand U6424 (N_6424,N_5808,N_5632);
nor U6425 (N_6425,N_5624,N_5626);
nand U6426 (N_6426,N_5609,N_5577);
xnor U6427 (N_6427,N_5938,N_5794);
xor U6428 (N_6428,N_5476,N_5455);
nand U6429 (N_6429,N_5617,N_5357);
nand U6430 (N_6430,N_5383,N_5970);
nand U6431 (N_6431,N_5438,N_5813);
xor U6432 (N_6432,N_5757,N_5536);
nor U6433 (N_6433,N_5400,N_5324);
or U6434 (N_6434,N_5425,N_5373);
and U6435 (N_6435,N_5366,N_5788);
nand U6436 (N_6436,N_5486,N_5732);
or U6437 (N_6437,N_5281,N_5912);
and U6438 (N_6438,N_5986,N_5729);
xnor U6439 (N_6439,N_5608,N_5967);
or U6440 (N_6440,N_5729,N_5615);
nor U6441 (N_6441,N_5719,N_5496);
xor U6442 (N_6442,N_5487,N_5824);
nand U6443 (N_6443,N_5955,N_5827);
nand U6444 (N_6444,N_5672,N_5860);
or U6445 (N_6445,N_5722,N_5900);
xnor U6446 (N_6446,N_5503,N_5492);
xnor U6447 (N_6447,N_5754,N_5582);
or U6448 (N_6448,N_5266,N_5510);
or U6449 (N_6449,N_5529,N_5462);
and U6450 (N_6450,N_5478,N_5403);
nand U6451 (N_6451,N_5574,N_5816);
nor U6452 (N_6452,N_5897,N_5837);
or U6453 (N_6453,N_5624,N_5341);
and U6454 (N_6454,N_5612,N_5686);
nor U6455 (N_6455,N_5541,N_5372);
and U6456 (N_6456,N_5362,N_5744);
nor U6457 (N_6457,N_5326,N_5400);
nor U6458 (N_6458,N_5598,N_5745);
xor U6459 (N_6459,N_5698,N_5545);
or U6460 (N_6460,N_5949,N_5253);
nand U6461 (N_6461,N_5947,N_5276);
nor U6462 (N_6462,N_5786,N_5450);
nor U6463 (N_6463,N_5962,N_5833);
nand U6464 (N_6464,N_5628,N_5665);
or U6465 (N_6465,N_5770,N_5455);
and U6466 (N_6466,N_5975,N_5977);
nor U6467 (N_6467,N_5532,N_5654);
xnor U6468 (N_6468,N_5561,N_5429);
and U6469 (N_6469,N_5693,N_5720);
nand U6470 (N_6470,N_5913,N_5462);
or U6471 (N_6471,N_5367,N_5456);
nand U6472 (N_6472,N_5825,N_5854);
xnor U6473 (N_6473,N_5598,N_5813);
and U6474 (N_6474,N_5917,N_5851);
nand U6475 (N_6475,N_5597,N_5719);
xnor U6476 (N_6476,N_5633,N_5819);
and U6477 (N_6477,N_5449,N_5533);
nand U6478 (N_6478,N_5292,N_5546);
xnor U6479 (N_6479,N_5822,N_5265);
or U6480 (N_6480,N_5699,N_5920);
or U6481 (N_6481,N_5974,N_5641);
and U6482 (N_6482,N_5267,N_5859);
xor U6483 (N_6483,N_5937,N_5610);
nand U6484 (N_6484,N_5922,N_5880);
nor U6485 (N_6485,N_5418,N_5989);
or U6486 (N_6486,N_5304,N_5385);
or U6487 (N_6487,N_5846,N_5848);
nand U6488 (N_6488,N_5348,N_5733);
or U6489 (N_6489,N_5705,N_5887);
nor U6490 (N_6490,N_5483,N_5835);
nand U6491 (N_6491,N_5698,N_5921);
or U6492 (N_6492,N_5985,N_5815);
or U6493 (N_6493,N_5965,N_5901);
nor U6494 (N_6494,N_5690,N_5383);
nor U6495 (N_6495,N_5715,N_5417);
nand U6496 (N_6496,N_5913,N_5729);
or U6497 (N_6497,N_5783,N_5476);
or U6498 (N_6498,N_5882,N_5565);
nor U6499 (N_6499,N_5398,N_5671);
nand U6500 (N_6500,N_5681,N_5896);
nand U6501 (N_6501,N_5356,N_5282);
xnor U6502 (N_6502,N_5766,N_5846);
and U6503 (N_6503,N_5286,N_5469);
xnor U6504 (N_6504,N_5310,N_5867);
nor U6505 (N_6505,N_5472,N_5639);
nand U6506 (N_6506,N_5646,N_5778);
or U6507 (N_6507,N_5943,N_5359);
and U6508 (N_6508,N_5790,N_5387);
xnor U6509 (N_6509,N_5664,N_5365);
or U6510 (N_6510,N_5530,N_5828);
and U6511 (N_6511,N_5490,N_5455);
and U6512 (N_6512,N_5807,N_5512);
and U6513 (N_6513,N_5424,N_5820);
or U6514 (N_6514,N_5881,N_5469);
xnor U6515 (N_6515,N_5672,N_5748);
xor U6516 (N_6516,N_5576,N_5338);
nor U6517 (N_6517,N_5484,N_5406);
nand U6518 (N_6518,N_5798,N_5832);
xnor U6519 (N_6519,N_5807,N_5267);
or U6520 (N_6520,N_5268,N_5913);
or U6521 (N_6521,N_5441,N_5812);
nand U6522 (N_6522,N_5785,N_5386);
xnor U6523 (N_6523,N_5502,N_5633);
and U6524 (N_6524,N_5894,N_5671);
xnor U6525 (N_6525,N_5658,N_5814);
xor U6526 (N_6526,N_5859,N_5801);
xnor U6527 (N_6527,N_5446,N_5399);
nand U6528 (N_6528,N_5877,N_5906);
nand U6529 (N_6529,N_5886,N_5670);
nand U6530 (N_6530,N_5554,N_5683);
xor U6531 (N_6531,N_5837,N_5900);
or U6532 (N_6532,N_5271,N_5533);
xor U6533 (N_6533,N_5465,N_5815);
or U6534 (N_6534,N_5355,N_5768);
nand U6535 (N_6535,N_5316,N_5388);
and U6536 (N_6536,N_5801,N_5810);
xor U6537 (N_6537,N_5599,N_5520);
nor U6538 (N_6538,N_5342,N_5984);
nor U6539 (N_6539,N_5952,N_5934);
or U6540 (N_6540,N_5666,N_5850);
nand U6541 (N_6541,N_5874,N_5345);
nor U6542 (N_6542,N_5667,N_5304);
and U6543 (N_6543,N_5655,N_5420);
or U6544 (N_6544,N_5662,N_5571);
nor U6545 (N_6545,N_5771,N_5528);
nor U6546 (N_6546,N_5882,N_5785);
nand U6547 (N_6547,N_5472,N_5274);
xnor U6548 (N_6548,N_5864,N_5640);
xor U6549 (N_6549,N_5714,N_5444);
xor U6550 (N_6550,N_5759,N_5864);
nor U6551 (N_6551,N_5526,N_5866);
nand U6552 (N_6552,N_5672,N_5438);
and U6553 (N_6553,N_5392,N_5374);
and U6554 (N_6554,N_5918,N_5487);
and U6555 (N_6555,N_5659,N_5810);
nor U6556 (N_6556,N_5921,N_5326);
nor U6557 (N_6557,N_5794,N_5500);
nor U6558 (N_6558,N_5760,N_5516);
nand U6559 (N_6559,N_5467,N_5860);
and U6560 (N_6560,N_5885,N_5310);
or U6561 (N_6561,N_5529,N_5389);
nor U6562 (N_6562,N_5365,N_5597);
nand U6563 (N_6563,N_5499,N_5342);
or U6564 (N_6564,N_5724,N_5945);
nand U6565 (N_6565,N_5262,N_5630);
xor U6566 (N_6566,N_5642,N_5752);
or U6567 (N_6567,N_5545,N_5613);
nand U6568 (N_6568,N_5846,N_5268);
nand U6569 (N_6569,N_5970,N_5615);
xor U6570 (N_6570,N_5917,N_5501);
or U6571 (N_6571,N_5270,N_5869);
nand U6572 (N_6572,N_5806,N_5596);
or U6573 (N_6573,N_5781,N_5684);
xnor U6574 (N_6574,N_5790,N_5992);
nor U6575 (N_6575,N_5285,N_5640);
nand U6576 (N_6576,N_5393,N_5854);
xnor U6577 (N_6577,N_5357,N_5650);
nor U6578 (N_6578,N_5300,N_5416);
nor U6579 (N_6579,N_5640,N_5532);
xor U6580 (N_6580,N_5669,N_5693);
nor U6581 (N_6581,N_5461,N_5587);
and U6582 (N_6582,N_5988,N_5507);
nor U6583 (N_6583,N_5645,N_5796);
nor U6584 (N_6584,N_5996,N_5608);
nor U6585 (N_6585,N_5926,N_5805);
or U6586 (N_6586,N_5299,N_5294);
or U6587 (N_6587,N_5644,N_5517);
xnor U6588 (N_6588,N_5897,N_5417);
or U6589 (N_6589,N_5655,N_5257);
or U6590 (N_6590,N_5824,N_5829);
or U6591 (N_6591,N_5300,N_5483);
and U6592 (N_6592,N_5591,N_5442);
nor U6593 (N_6593,N_5553,N_5410);
xnor U6594 (N_6594,N_5419,N_5988);
xnor U6595 (N_6595,N_5785,N_5966);
nand U6596 (N_6596,N_5912,N_5366);
nand U6597 (N_6597,N_5570,N_5719);
or U6598 (N_6598,N_5757,N_5559);
or U6599 (N_6599,N_5344,N_5828);
nor U6600 (N_6600,N_5944,N_5725);
xor U6601 (N_6601,N_5521,N_5377);
and U6602 (N_6602,N_5933,N_5288);
nand U6603 (N_6603,N_5410,N_5564);
or U6604 (N_6604,N_5606,N_5729);
nand U6605 (N_6605,N_5587,N_5697);
nor U6606 (N_6606,N_5881,N_5947);
or U6607 (N_6607,N_5769,N_5881);
and U6608 (N_6608,N_5594,N_5685);
nor U6609 (N_6609,N_5355,N_5585);
nor U6610 (N_6610,N_5331,N_5905);
nor U6611 (N_6611,N_5447,N_5270);
or U6612 (N_6612,N_5709,N_5951);
or U6613 (N_6613,N_5388,N_5763);
and U6614 (N_6614,N_5425,N_5759);
or U6615 (N_6615,N_5984,N_5897);
nor U6616 (N_6616,N_5261,N_5411);
nor U6617 (N_6617,N_5504,N_5433);
xor U6618 (N_6618,N_5549,N_5637);
or U6619 (N_6619,N_5683,N_5970);
nor U6620 (N_6620,N_5814,N_5601);
nand U6621 (N_6621,N_5714,N_5304);
xnor U6622 (N_6622,N_5463,N_5668);
nand U6623 (N_6623,N_5632,N_5932);
nand U6624 (N_6624,N_5940,N_5522);
xnor U6625 (N_6625,N_5970,N_5753);
xor U6626 (N_6626,N_5792,N_5892);
and U6627 (N_6627,N_5765,N_5468);
nor U6628 (N_6628,N_5251,N_5559);
and U6629 (N_6629,N_5717,N_5571);
or U6630 (N_6630,N_5860,N_5266);
nor U6631 (N_6631,N_5279,N_5567);
nand U6632 (N_6632,N_5433,N_5712);
or U6633 (N_6633,N_5949,N_5724);
nand U6634 (N_6634,N_5953,N_5763);
nor U6635 (N_6635,N_5434,N_5787);
nor U6636 (N_6636,N_5605,N_5930);
and U6637 (N_6637,N_5511,N_5615);
and U6638 (N_6638,N_5733,N_5583);
nor U6639 (N_6639,N_5986,N_5828);
nor U6640 (N_6640,N_5649,N_5581);
xnor U6641 (N_6641,N_5932,N_5267);
and U6642 (N_6642,N_5262,N_5474);
nand U6643 (N_6643,N_5902,N_5843);
nand U6644 (N_6644,N_5619,N_5639);
nand U6645 (N_6645,N_5609,N_5606);
nor U6646 (N_6646,N_5903,N_5791);
nand U6647 (N_6647,N_5900,N_5786);
xor U6648 (N_6648,N_5512,N_5896);
and U6649 (N_6649,N_5310,N_5909);
nand U6650 (N_6650,N_5282,N_5467);
nor U6651 (N_6651,N_5938,N_5782);
or U6652 (N_6652,N_5759,N_5849);
or U6653 (N_6653,N_5475,N_5911);
and U6654 (N_6654,N_5990,N_5536);
nor U6655 (N_6655,N_5566,N_5260);
xnor U6656 (N_6656,N_5270,N_5653);
nor U6657 (N_6657,N_5917,N_5579);
nand U6658 (N_6658,N_5265,N_5251);
xor U6659 (N_6659,N_5975,N_5394);
nand U6660 (N_6660,N_5650,N_5641);
nor U6661 (N_6661,N_5642,N_5506);
nor U6662 (N_6662,N_5797,N_5633);
nor U6663 (N_6663,N_5711,N_5615);
nand U6664 (N_6664,N_5799,N_5685);
nor U6665 (N_6665,N_5524,N_5462);
xor U6666 (N_6666,N_5503,N_5565);
nor U6667 (N_6667,N_5370,N_5368);
and U6668 (N_6668,N_5691,N_5811);
and U6669 (N_6669,N_5474,N_5761);
nand U6670 (N_6670,N_5901,N_5789);
nor U6671 (N_6671,N_5970,N_5910);
xnor U6672 (N_6672,N_5626,N_5588);
nor U6673 (N_6673,N_5729,N_5590);
xor U6674 (N_6674,N_5426,N_5646);
xnor U6675 (N_6675,N_5771,N_5396);
and U6676 (N_6676,N_5342,N_5533);
nand U6677 (N_6677,N_5954,N_5706);
and U6678 (N_6678,N_5619,N_5491);
and U6679 (N_6679,N_5809,N_5919);
and U6680 (N_6680,N_5647,N_5284);
xor U6681 (N_6681,N_5645,N_5493);
nor U6682 (N_6682,N_5960,N_5388);
and U6683 (N_6683,N_5328,N_5329);
nand U6684 (N_6684,N_5518,N_5467);
xor U6685 (N_6685,N_5839,N_5812);
nor U6686 (N_6686,N_5696,N_5779);
and U6687 (N_6687,N_5379,N_5502);
or U6688 (N_6688,N_5802,N_5948);
or U6689 (N_6689,N_5347,N_5772);
or U6690 (N_6690,N_5611,N_5480);
or U6691 (N_6691,N_5817,N_5554);
xnor U6692 (N_6692,N_5607,N_5403);
nand U6693 (N_6693,N_5426,N_5544);
and U6694 (N_6694,N_5475,N_5613);
nor U6695 (N_6695,N_5874,N_5508);
and U6696 (N_6696,N_5838,N_5853);
xor U6697 (N_6697,N_5977,N_5398);
xnor U6698 (N_6698,N_5483,N_5290);
xor U6699 (N_6699,N_5682,N_5395);
or U6700 (N_6700,N_5433,N_5528);
xor U6701 (N_6701,N_5675,N_5362);
xnor U6702 (N_6702,N_5497,N_5406);
and U6703 (N_6703,N_5952,N_5514);
xor U6704 (N_6704,N_5371,N_5284);
nor U6705 (N_6705,N_5662,N_5585);
nand U6706 (N_6706,N_5940,N_5645);
nor U6707 (N_6707,N_5644,N_5481);
or U6708 (N_6708,N_5581,N_5604);
nor U6709 (N_6709,N_5519,N_5284);
or U6710 (N_6710,N_5321,N_5389);
nor U6711 (N_6711,N_5953,N_5259);
nand U6712 (N_6712,N_5867,N_5742);
nor U6713 (N_6713,N_5967,N_5654);
and U6714 (N_6714,N_5956,N_5547);
nor U6715 (N_6715,N_5550,N_5404);
xnor U6716 (N_6716,N_5780,N_5502);
nand U6717 (N_6717,N_5788,N_5912);
and U6718 (N_6718,N_5352,N_5329);
and U6719 (N_6719,N_5914,N_5912);
or U6720 (N_6720,N_5496,N_5890);
or U6721 (N_6721,N_5481,N_5254);
xor U6722 (N_6722,N_5720,N_5749);
or U6723 (N_6723,N_5702,N_5765);
or U6724 (N_6724,N_5345,N_5334);
and U6725 (N_6725,N_5499,N_5445);
xnor U6726 (N_6726,N_5842,N_5528);
nand U6727 (N_6727,N_5533,N_5566);
nand U6728 (N_6728,N_5250,N_5791);
xor U6729 (N_6729,N_5697,N_5938);
xor U6730 (N_6730,N_5558,N_5968);
xnor U6731 (N_6731,N_5593,N_5266);
or U6732 (N_6732,N_5255,N_5407);
nor U6733 (N_6733,N_5565,N_5872);
nor U6734 (N_6734,N_5739,N_5284);
or U6735 (N_6735,N_5573,N_5742);
xor U6736 (N_6736,N_5853,N_5261);
or U6737 (N_6737,N_5712,N_5482);
xor U6738 (N_6738,N_5724,N_5474);
nor U6739 (N_6739,N_5537,N_5668);
xnor U6740 (N_6740,N_5460,N_5846);
or U6741 (N_6741,N_5277,N_5701);
or U6742 (N_6742,N_5355,N_5689);
nor U6743 (N_6743,N_5462,N_5372);
or U6744 (N_6744,N_5928,N_5622);
or U6745 (N_6745,N_5560,N_5998);
nand U6746 (N_6746,N_5605,N_5414);
nor U6747 (N_6747,N_5527,N_5617);
nor U6748 (N_6748,N_5727,N_5398);
and U6749 (N_6749,N_5713,N_5763);
nor U6750 (N_6750,N_6602,N_6146);
or U6751 (N_6751,N_6411,N_6154);
or U6752 (N_6752,N_6649,N_6669);
and U6753 (N_6753,N_6662,N_6706);
nand U6754 (N_6754,N_6027,N_6538);
xor U6755 (N_6755,N_6358,N_6524);
xor U6756 (N_6756,N_6223,N_6641);
or U6757 (N_6757,N_6244,N_6242);
xnor U6758 (N_6758,N_6118,N_6640);
nand U6759 (N_6759,N_6420,N_6664);
and U6760 (N_6760,N_6733,N_6627);
nor U6761 (N_6761,N_6167,N_6594);
and U6762 (N_6762,N_6066,N_6291);
nand U6763 (N_6763,N_6261,N_6425);
or U6764 (N_6764,N_6743,N_6209);
nand U6765 (N_6765,N_6233,N_6406);
xor U6766 (N_6766,N_6289,N_6330);
or U6767 (N_6767,N_6060,N_6539);
nor U6768 (N_6768,N_6587,N_6408);
nor U6769 (N_6769,N_6034,N_6676);
nor U6770 (N_6770,N_6413,N_6115);
xnor U6771 (N_6771,N_6647,N_6482);
nor U6772 (N_6772,N_6504,N_6432);
and U6773 (N_6773,N_6131,N_6045);
xor U6774 (N_6774,N_6449,N_6452);
nor U6775 (N_6775,N_6389,N_6635);
nor U6776 (N_6776,N_6438,N_6596);
nor U6777 (N_6777,N_6100,N_6734);
nand U6778 (N_6778,N_6347,N_6345);
xor U6779 (N_6779,N_6410,N_6670);
and U6780 (N_6780,N_6056,N_6469);
and U6781 (N_6781,N_6334,N_6580);
and U6782 (N_6782,N_6570,N_6661);
nor U6783 (N_6783,N_6283,N_6072);
or U6784 (N_6784,N_6310,N_6551);
xor U6785 (N_6785,N_6695,N_6514);
nand U6786 (N_6786,N_6621,N_6412);
xor U6787 (N_6787,N_6387,N_6161);
or U6788 (N_6788,N_6386,N_6375);
or U6789 (N_6789,N_6337,N_6571);
xor U6790 (N_6790,N_6404,N_6303);
nor U6791 (N_6791,N_6267,N_6014);
and U6792 (N_6792,N_6035,N_6294);
nand U6793 (N_6793,N_6644,N_6129);
nand U6794 (N_6794,N_6363,N_6663);
nand U6795 (N_6795,N_6077,N_6295);
nand U6796 (N_6796,N_6660,N_6119);
xnor U6797 (N_6797,N_6466,N_6665);
nand U6798 (N_6798,N_6147,N_6331);
and U6799 (N_6799,N_6284,N_6276);
or U6800 (N_6800,N_6201,N_6431);
or U6801 (N_6801,N_6632,N_6318);
or U6802 (N_6802,N_6062,N_6455);
xor U6803 (N_6803,N_6237,N_6280);
nor U6804 (N_6804,N_6374,N_6747);
nand U6805 (N_6805,N_6473,N_6262);
xnor U6806 (N_6806,N_6332,N_6155);
and U6807 (N_6807,N_6478,N_6654);
and U6808 (N_6808,N_6107,N_6122);
nand U6809 (N_6809,N_6707,N_6400);
nor U6810 (N_6810,N_6216,N_6137);
nand U6811 (N_6811,N_6275,N_6217);
nor U6812 (N_6812,N_6206,N_6057);
or U6813 (N_6813,N_6555,N_6023);
xor U6814 (N_6814,N_6719,N_6436);
or U6815 (N_6815,N_6177,N_6189);
xor U6816 (N_6816,N_6102,N_6204);
or U6817 (N_6817,N_6203,N_6456);
and U6818 (N_6818,N_6577,N_6317);
or U6819 (N_6819,N_6439,N_6424);
and U6820 (N_6820,N_6191,N_6166);
nand U6821 (N_6821,N_6272,N_6357);
and U6822 (N_6822,N_6705,N_6569);
and U6823 (N_6823,N_6058,N_6630);
nor U6824 (N_6824,N_6396,N_6017);
and U6825 (N_6825,N_6689,N_6721);
nand U6826 (N_6826,N_6239,N_6629);
nand U6827 (N_6827,N_6612,N_6697);
nand U6828 (N_6828,N_6528,N_6433);
xnor U6829 (N_6829,N_6497,N_6659);
or U6830 (N_6830,N_6574,N_6324);
and U6831 (N_6831,N_6454,N_6255);
nand U6832 (N_6832,N_6043,N_6013);
and U6833 (N_6833,N_6590,N_6732);
or U6834 (N_6834,N_6311,N_6414);
and U6835 (N_6835,N_6299,N_6579);
nand U6836 (N_6836,N_6749,N_6366);
or U6837 (N_6837,N_6278,N_6376);
or U6838 (N_6838,N_6200,N_6249);
xor U6839 (N_6839,N_6467,N_6541);
nand U6840 (N_6840,N_6053,N_6365);
and U6841 (N_6841,N_6518,N_6675);
and U6842 (N_6842,N_6002,N_6476);
xnor U6843 (N_6843,N_6111,N_6063);
xnor U6844 (N_6844,N_6718,N_6254);
or U6845 (N_6845,N_6008,N_6051);
xor U6846 (N_6846,N_6407,N_6195);
nand U6847 (N_6847,N_6133,N_6336);
or U6848 (N_6848,N_6353,N_6715);
xnor U6849 (N_6849,N_6625,N_6428);
nand U6850 (N_6850,N_6339,N_6231);
xnor U6851 (N_6851,N_6548,N_6540);
or U6852 (N_6852,N_6495,N_6575);
nor U6853 (N_6853,N_6724,N_6050);
xnor U6854 (N_6854,N_6517,N_6543);
or U6855 (N_6855,N_6595,N_6270);
xor U6856 (N_6856,N_6342,N_6544);
or U6857 (N_6857,N_6487,N_6722);
or U6858 (N_6858,N_6698,N_6636);
xnor U6859 (N_6859,N_6522,N_6315);
nand U6860 (N_6860,N_6713,N_6156);
or U6861 (N_6861,N_6598,N_6246);
nand U6862 (N_6862,N_6116,N_6714);
xnor U6863 (N_6863,N_6513,N_6222);
nand U6864 (N_6864,N_6304,N_6639);
and U6865 (N_6865,N_6308,N_6091);
nand U6866 (N_6866,N_6003,N_6181);
and U6867 (N_6867,N_6461,N_6490);
xnor U6868 (N_6868,N_6323,N_6069);
xnor U6869 (N_6869,N_6033,N_6576);
nor U6870 (N_6870,N_6188,N_6020);
nand U6871 (N_6871,N_6550,N_6282);
and U6872 (N_6872,N_6638,N_6251);
or U6873 (N_6873,N_6109,N_6441);
nor U6874 (N_6874,N_6486,N_6464);
xor U6875 (N_6875,N_6125,N_6593);
nand U6876 (N_6876,N_6040,N_6263);
xnor U6877 (N_6877,N_6578,N_6730);
xor U6878 (N_6878,N_6235,N_6321);
or U6879 (N_6879,N_6509,N_6148);
nor U6880 (N_6880,N_6668,N_6301);
or U6881 (N_6881,N_6187,N_6742);
xor U6882 (N_6882,N_6226,N_6494);
and U6883 (N_6883,N_6159,N_6613);
or U6884 (N_6884,N_6700,N_6309);
nand U6885 (N_6885,N_6736,N_6185);
and U6886 (N_6886,N_6606,N_6319);
xor U6887 (N_6887,N_6150,N_6442);
or U6888 (N_6888,N_6637,N_6238);
or U6889 (N_6889,N_6471,N_6483);
xor U6890 (N_6890,N_6437,N_6610);
and U6891 (N_6891,N_6620,N_6564);
nand U6892 (N_6892,N_6004,N_6470);
nand U6893 (N_6893,N_6197,N_6545);
xnor U6894 (N_6894,N_6170,N_6274);
xor U6895 (N_6895,N_6059,N_6520);
xnor U6896 (N_6896,N_6126,N_6288);
nand U6897 (N_6897,N_6219,N_6287);
or U6898 (N_6898,N_6371,N_6333);
nand U6899 (N_6899,N_6502,N_6601);
xor U6900 (N_6900,N_6380,N_6247);
and U6901 (N_6901,N_6446,N_6085);
or U6902 (N_6902,N_6190,N_6015);
xnor U6903 (N_6903,N_6515,N_6562);
xor U6904 (N_6904,N_6329,N_6307);
or U6905 (N_6905,N_6523,N_6563);
and U6906 (N_6906,N_6508,N_6068);
or U6907 (N_6907,N_6549,N_6395);
nand U6908 (N_6908,N_6526,N_6163);
nor U6909 (N_6909,N_6740,N_6300);
and U6910 (N_6910,N_6584,N_6152);
and U6911 (N_6911,N_6393,N_6082);
nand U6912 (N_6912,N_6305,N_6101);
nand U6913 (N_6913,N_6653,N_6658);
nor U6914 (N_6914,N_6273,N_6685);
nor U6915 (N_6915,N_6018,N_6440);
nand U6916 (N_6916,N_6343,N_6416);
and U6917 (N_6917,N_6123,N_6546);
nor U6918 (N_6918,N_6113,N_6568);
xor U6919 (N_6919,N_6566,N_6506);
nor U6920 (N_6920,N_6480,N_6535);
xnor U6921 (N_6921,N_6739,N_6046);
or U6922 (N_6922,N_6616,N_6415);
and U6923 (N_6923,N_6007,N_6344);
nand U6924 (N_6924,N_6402,N_6117);
and U6925 (N_6925,N_6348,N_6302);
or U6926 (N_6926,N_6199,N_6748);
nor U6927 (N_6927,N_6565,N_6373);
or U6928 (N_6928,N_6090,N_6481);
nor U6929 (N_6929,N_6392,N_6362);
nand U6930 (N_6930,N_6022,N_6368);
nand U6931 (N_6931,N_6269,N_6656);
xnor U6932 (N_6932,N_6558,N_6006);
nand U6933 (N_6933,N_6145,N_6445);
or U6934 (N_6934,N_6005,N_6037);
or U6935 (N_6935,N_6600,N_6691);
nor U6936 (N_6936,N_6552,N_6361);
or U6937 (N_6937,N_6248,N_6720);
and U6938 (N_6938,N_6328,N_6143);
or U6939 (N_6939,N_6423,N_6080);
nand U6940 (N_6940,N_6174,N_6001);
and U6941 (N_6941,N_6048,N_6626);
and U6942 (N_6942,N_6207,N_6493);
nor U6943 (N_6943,N_6028,N_6384);
and U6944 (N_6944,N_6088,N_6218);
nand U6945 (N_6945,N_6712,N_6265);
or U6946 (N_6946,N_6196,N_6553);
nand U6947 (N_6947,N_6671,N_6643);
and U6948 (N_6948,N_6205,N_6099);
or U6949 (N_6949,N_6175,N_6128);
nand U6950 (N_6950,N_6614,N_6475);
xnor U6951 (N_6951,N_6044,N_6220);
nor U6952 (N_6952,N_6227,N_6687);
or U6953 (N_6953,N_6316,N_6709);
or U6954 (N_6954,N_6746,N_6019);
nand U6955 (N_6955,N_6106,N_6460);
xnor U6956 (N_6956,N_6078,N_6211);
nor U6957 (N_6957,N_6176,N_6474);
nand U6958 (N_6958,N_6529,N_6492);
and U6959 (N_6959,N_6427,N_6041);
or U6960 (N_6960,N_6186,N_6448);
nor U6961 (N_6961,N_6607,N_6266);
xor U6962 (N_6962,N_6184,N_6096);
and U6963 (N_6963,N_6049,N_6067);
xor U6964 (N_6964,N_6516,N_6030);
xnor U6965 (N_6965,N_6443,N_6326);
xor U6966 (N_6966,N_6479,N_6491);
or U6967 (N_6967,N_6723,N_6042);
xor U6968 (N_6968,N_6631,N_6694);
nand U6969 (N_6969,N_6055,N_6025);
nand U6970 (N_6970,N_6338,N_6230);
xnor U6971 (N_6971,N_6292,N_6378);
xnor U6972 (N_6972,N_6547,N_6253);
or U6973 (N_6973,N_6104,N_6617);
or U6974 (N_6974,N_6604,N_6560);
nor U6975 (N_6975,N_6245,N_6696);
and U6976 (N_6976,N_6026,N_6277);
xor U6977 (N_6977,N_6016,N_6704);
or U6978 (N_6978,N_6735,N_6716);
nor U6979 (N_6979,N_6390,N_6141);
and U6980 (N_6980,N_6110,N_6369);
xor U6981 (N_6981,N_6744,N_6214);
nor U6982 (N_6982,N_6652,N_6450);
and U6983 (N_6983,N_6367,N_6252);
nor U6984 (N_6984,N_6194,N_6000);
or U6985 (N_6985,N_6711,N_6421);
nand U6986 (N_6986,N_6674,N_6701);
and U6987 (N_6987,N_6071,N_6619);
nor U6988 (N_6988,N_6359,N_6298);
nor U6989 (N_6989,N_6325,N_6618);
and U6990 (N_6990,N_6038,N_6710);
xnor U6991 (N_6991,N_6592,N_6160);
nand U6992 (N_6992,N_6212,N_6312);
and U6993 (N_6993,N_6457,N_6228);
xor U6994 (N_6994,N_6398,N_6105);
or U6995 (N_6995,N_6095,N_6605);
nand U6996 (N_6996,N_6745,N_6335);
or U6997 (N_6997,N_6597,N_6271);
or U6998 (N_6998,N_6135,N_6165);
xnor U6999 (N_6999,N_6702,N_6532);
nor U7000 (N_7000,N_6134,N_6079);
and U7001 (N_7001,N_6405,N_6634);
and U7002 (N_7002,N_6561,N_6542);
and U7003 (N_7003,N_6098,N_6192);
nand U7004 (N_7004,N_6703,N_6388);
or U7005 (N_7005,N_6285,N_6477);
or U7006 (N_7006,N_6666,N_6628);
or U7007 (N_7007,N_6236,N_6484);
and U7008 (N_7008,N_6472,N_6435);
nor U7009 (N_7009,N_6401,N_6505);
xor U7010 (N_7010,N_6281,N_6171);
nor U7011 (N_7011,N_6036,N_6573);
or U7012 (N_7012,N_6708,N_6340);
xnor U7013 (N_7013,N_6264,N_6667);
xnor U7014 (N_7014,N_6232,N_6519);
and U7015 (N_7015,N_6064,N_6651);
xor U7016 (N_7016,N_6417,N_6009);
nand U7017 (N_7017,N_6447,N_6453);
nand U7018 (N_7018,N_6097,N_6142);
nand U7019 (N_7019,N_6260,N_6286);
or U7020 (N_7020,N_6729,N_6582);
xnor U7021 (N_7021,N_6136,N_6451);
or U7022 (N_7022,N_6021,N_6121);
nor U7023 (N_7023,N_6372,N_6213);
and U7024 (N_7024,N_6379,N_6609);
or U7025 (N_7025,N_6370,N_6683);
nand U7026 (N_7026,N_6503,N_6583);
nand U7027 (N_7027,N_6256,N_6149);
nand U7028 (N_7028,N_6157,N_6559);
nor U7029 (N_7029,N_6717,N_6633);
nand U7030 (N_7030,N_6728,N_6693);
nor U7031 (N_7031,N_6180,N_6500);
and U7032 (N_7032,N_6385,N_6243);
xor U7033 (N_7033,N_6164,N_6397);
nor U7034 (N_7034,N_6293,N_6527);
and U7035 (N_7035,N_6418,N_6350);
xnor U7036 (N_7036,N_6250,N_6151);
or U7037 (N_7037,N_6429,N_6692);
xor U7038 (N_7038,N_6341,N_6556);
xnor U7039 (N_7039,N_6144,N_6726);
xnor U7040 (N_7040,N_6737,N_6258);
and U7041 (N_7041,N_6202,N_6496);
xor U7042 (N_7042,N_6224,N_6383);
nand U7043 (N_7043,N_6534,N_6130);
nor U7044 (N_7044,N_6168,N_6684);
and U7045 (N_7045,N_6081,N_6586);
nand U7046 (N_7046,N_6738,N_6531);
and U7047 (N_7047,N_6622,N_6198);
nor U7048 (N_7048,N_6382,N_6179);
xor U7049 (N_7049,N_6591,N_6221);
nor U7050 (N_7050,N_6585,N_6327);
and U7051 (N_7051,N_6377,N_6525);
xnor U7052 (N_7052,N_6306,N_6349);
or U7053 (N_7053,N_6409,N_6391);
and U7054 (N_7054,N_6032,N_6462);
nor U7055 (N_7055,N_6533,N_6047);
and U7056 (N_7056,N_6677,N_6094);
nand U7057 (N_7057,N_6229,N_6089);
or U7058 (N_7058,N_6065,N_6741);
or U7059 (N_7059,N_6183,N_6076);
and U7060 (N_7060,N_6646,N_6193);
xnor U7061 (N_7061,N_6010,N_6182);
xor U7062 (N_7062,N_6364,N_6498);
and U7063 (N_7063,N_6029,N_6039);
and U7064 (N_7064,N_6208,N_6536);
nor U7065 (N_7065,N_6158,N_6680);
and U7066 (N_7066,N_6011,N_6173);
nor U7067 (N_7067,N_6132,N_6314);
and U7068 (N_7068,N_6012,N_6690);
and U7069 (N_7069,N_6599,N_6240);
nand U7070 (N_7070,N_6162,N_6611);
or U7071 (N_7071,N_6727,N_6673);
or U7072 (N_7072,N_6521,N_6061);
and U7073 (N_7073,N_6103,N_6346);
nor U7074 (N_7074,N_6268,N_6083);
and U7075 (N_7075,N_6093,N_6031);
nand U7076 (N_7076,N_6725,N_6655);
nand U7077 (N_7077,N_6603,N_6394);
nor U7078 (N_7078,N_6468,N_6086);
or U7079 (N_7079,N_6322,N_6178);
nor U7080 (N_7080,N_6169,N_6124);
and U7081 (N_7081,N_6686,N_6114);
and U7082 (N_7082,N_6399,N_6485);
xor U7083 (N_7083,N_6225,N_6108);
xor U7084 (N_7084,N_6672,N_6112);
nand U7085 (N_7085,N_6444,N_6215);
nor U7086 (N_7086,N_6297,N_6731);
xor U7087 (N_7087,N_6355,N_6074);
nor U7088 (N_7088,N_6645,N_6352);
nor U7089 (N_7089,N_6422,N_6489);
nand U7090 (N_7090,N_6279,N_6140);
xnor U7091 (N_7091,N_6530,N_6501);
nand U7092 (N_7092,N_6507,N_6678);
and U7093 (N_7093,N_6463,N_6234);
nand U7094 (N_7094,N_6434,N_6120);
nand U7095 (N_7095,N_6581,N_6679);
nor U7096 (N_7096,N_6459,N_6465);
and U7097 (N_7097,N_6360,N_6087);
xnor U7098 (N_7098,N_6084,N_6588);
and U7099 (N_7099,N_6259,N_6511);
nand U7100 (N_7100,N_6313,N_6615);
nor U7101 (N_7101,N_6024,N_6642);
or U7102 (N_7102,N_6092,N_6296);
or U7103 (N_7103,N_6070,N_6241);
nor U7104 (N_7104,N_6127,N_6172);
nor U7105 (N_7105,N_6624,N_6512);
and U7106 (N_7106,N_6210,N_6537);
nor U7107 (N_7107,N_6682,N_6657);
nand U7108 (N_7108,N_6510,N_6290);
or U7109 (N_7109,N_6688,N_6426);
nor U7110 (N_7110,N_6403,N_6458);
or U7111 (N_7111,N_6320,N_6153);
nor U7112 (N_7112,N_6499,N_6554);
and U7113 (N_7113,N_6075,N_6650);
nor U7114 (N_7114,N_6354,N_6648);
and U7115 (N_7115,N_6419,N_6381);
and U7116 (N_7116,N_6589,N_6052);
nand U7117 (N_7117,N_6699,N_6138);
or U7118 (N_7118,N_6073,N_6681);
nand U7119 (N_7119,N_6488,N_6257);
nand U7120 (N_7120,N_6608,N_6623);
or U7121 (N_7121,N_6139,N_6572);
xor U7122 (N_7122,N_6567,N_6356);
nor U7123 (N_7123,N_6054,N_6557);
or U7124 (N_7124,N_6430,N_6351);
and U7125 (N_7125,N_6237,N_6566);
nor U7126 (N_7126,N_6430,N_6177);
nand U7127 (N_7127,N_6052,N_6543);
nand U7128 (N_7128,N_6241,N_6449);
nor U7129 (N_7129,N_6021,N_6132);
nor U7130 (N_7130,N_6177,N_6048);
nand U7131 (N_7131,N_6608,N_6596);
or U7132 (N_7132,N_6708,N_6424);
nand U7133 (N_7133,N_6720,N_6517);
or U7134 (N_7134,N_6674,N_6677);
nor U7135 (N_7135,N_6204,N_6028);
and U7136 (N_7136,N_6420,N_6559);
or U7137 (N_7137,N_6110,N_6313);
nor U7138 (N_7138,N_6152,N_6629);
or U7139 (N_7139,N_6697,N_6180);
xnor U7140 (N_7140,N_6264,N_6137);
nand U7141 (N_7141,N_6482,N_6725);
or U7142 (N_7142,N_6287,N_6183);
nand U7143 (N_7143,N_6054,N_6208);
nand U7144 (N_7144,N_6030,N_6502);
nor U7145 (N_7145,N_6723,N_6506);
or U7146 (N_7146,N_6442,N_6406);
and U7147 (N_7147,N_6207,N_6599);
nand U7148 (N_7148,N_6728,N_6376);
nor U7149 (N_7149,N_6340,N_6261);
xnor U7150 (N_7150,N_6322,N_6732);
or U7151 (N_7151,N_6302,N_6643);
xor U7152 (N_7152,N_6104,N_6173);
nor U7153 (N_7153,N_6217,N_6117);
nor U7154 (N_7154,N_6346,N_6395);
nand U7155 (N_7155,N_6020,N_6100);
nor U7156 (N_7156,N_6423,N_6394);
and U7157 (N_7157,N_6687,N_6406);
nor U7158 (N_7158,N_6068,N_6384);
nor U7159 (N_7159,N_6744,N_6345);
nor U7160 (N_7160,N_6656,N_6712);
xor U7161 (N_7161,N_6387,N_6116);
nand U7162 (N_7162,N_6540,N_6316);
xnor U7163 (N_7163,N_6076,N_6060);
xor U7164 (N_7164,N_6660,N_6169);
nand U7165 (N_7165,N_6120,N_6431);
xor U7166 (N_7166,N_6644,N_6464);
or U7167 (N_7167,N_6323,N_6693);
or U7168 (N_7168,N_6224,N_6465);
xor U7169 (N_7169,N_6093,N_6317);
and U7170 (N_7170,N_6219,N_6489);
nor U7171 (N_7171,N_6035,N_6480);
nand U7172 (N_7172,N_6580,N_6132);
nor U7173 (N_7173,N_6477,N_6435);
nor U7174 (N_7174,N_6519,N_6456);
nor U7175 (N_7175,N_6703,N_6397);
and U7176 (N_7176,N_6664,N_6676);
nand U7177 (N_7177,N_6053,N_6459);
nand U7178 (N_7178,N_6500,N_6362);
or U7179 (N_7179,N_6375,N_6153);
and U7180 (N_7180,N_6392,N_6565);
or U7181 (N_7181,N_6315,N_6228);
xnor U7182 (N_7182,N_6730,N_6267);
or U7183 (N_7183,N_6520,N_6742);
xor U7184 (N_7184,N_6370,N_6244);
nor U7185 (N_7185,N_6288,N_6688);
and U7186 (N_7186,N_6340,N_6112);
nor U7187 (N_7187,N_6537,N_6533);
nor U7188 (N_7188,N_6028,N_6717);
and U7189 (N_7189,N_6454,N_6590);
and U7190 (N_7190,N_6251,N_6345);
nand U7191 (N_7191,N_6688,N_6324);
nand U7192 (N_7192,N_6361,N_6093);
xnor U7193 (N_7193,N_6200,N_6689);
nor U7194 (N_7194,N_6018,N_6603);
or U7195 (N_7195,N_6551,N_6698);
and U7196 (N_7196,N_6061,N_6096);
nand U7197 (N_7197,N_6005,N_6639);
and U7198 (N_7198,N_6690,N_6383);
or U7199 (N_7199,N_6071,N_6088);
or U7200 (N_7200,N_6475,N_6447);
or U7201 (N_7201,N_6092,N_6338);
nand U7202 (N_7202,N_6061,N_6093);
and U7203 (N_7203,N_6479,N_6001);
nor U7204 (N_7204,N_6182,N_6463);
and U7205 (N_7205,N_6035,N_6188);
or U7206 (N_7206,N_6605,N_6547);
nor U7207 (N_7207,N_6662,N_6327);
or U7208 (N_7208,N_6197,N_6351);
nor U7209 (N_7209,N_6572,N_6317);
or U7210 (N_7210,N_6600,N_6166);
nand U7211 (N_7211,N_6378,N_6676);
nor U7212 (N_7212,N_6388,N_6185);
and U7213 (N_7213,N_6073,N_6129);
nor U7214 (N_7214,N_6422,N_6430);
xor U7215 (N_7215,N_6171,N_6525);
or U7216 (N_7216,N_6708,N_6600);
xnor U7217 (N_7217,N_6519,N_6260);
nor U7218 (N_7218,N_6715,N_6198);
or U7219 (N_7219,N_6170,N_6353);
nor U7220 (N_7220,N_6168,N_6022);
nand U7221 (N_7221,N_6727,N_6155);
or U7222 (N_7222,N_6698,N_6102);
or U7223 (N_7223,N_6000,N_6563);
nand U7224 (N_7224,N_6134,N_6159);
xnor U7225 (N_7225,N_6464,N_6570);
xnor U7226 (N_7226,N_6159,N_6471);
and U7227 (N_7227,N_6261,N_6532);
xnor U7228 (N_7228,N_6627,N_6164);
or U7229 (N_7229,N_6378,N_6246);
and U7230 (N_7230,N_6130,N_6681);
nor U7231 (N_7231,N_6717,N_6447);
or U7232 (N_7232,N_6114,N_6510);
nand U7233 (N_7233,N_6224,N_6062);
or U7234 (N_7234,N_6682,N_6000);
or U7235 (N_7235,N_6240,N_6014);
nor U7236 (N_7236,N_6691,N_6427);
and U7237 (N_7237,N_6170,N_6565);
nor U7238 (N_7238,N_6117,N_6449);
xor U7239 (N_7239,N_6045,N_6552);
and U7240 (N_7240,N_6533,N_6666);
nor U7241 (N_7241,N_6243,N_6599);
nand U7242 (N_7242,N_6509,N_6054);
xnor U7243 (N_7243,N_6653,N_6738);
xnor U7244 (N_7244,N_6295,N_6408);
nand U7245 (N_7245,N_6626,N_6217);
nand U7246 (N_7246,N_6678,N_6355);
or U7247 (N_7247,N_6115,N_6186);
nor U7248 (N_7248,N_6085,N_6053);
or U7249 (N_7249,N_6262,N_6043);
nand U7250 (N_7250,N_6347,N_6690);
nor U7251 (N_7251,N_6270,N_6600);
xor U7252 (N_7252,N_6254,N_6744);
and U7253 (N_7253,N_6370,N_6235);
xnor U7254 (N_7254,N_6495,N_6322);
nor U7255 (N_7255,N_6563,N_6527);
nor U7256 (N_7256,N_6745,N_6479);
nand U7257 (N_7257,N_6362,N_6638);
xor U7258 (N_7258,N_6631,N_6318);
nor U7259 (N_7259,N_6401,N_6309);
or U7260 (N_7260,N_6398,N_6060);
xnor U7261 (N_7261,N_6610,N_6031);
or U7262 (N_7262,N_6639,N_6135);
and U7263 (N_7263,N_6742,N_6541);
nor U7264 (N_7264,N_6512,N_6378);
and U7265 (N_7265,N_6181,N_6408);
xnor U7266 (N_7266,N_6042,N_6173);
xor U7267 (N_7267,N_6708,N_6407);
nor U7268 (N_7268,N_6343,N_6531);
or U7269 (N_7269,N_6527,N_6648);
and U7270 (N_7270,N_6515,N_6020);
and U7271 (N_7271,N_6121,N_6056);
nand U7272 (N_7272,N_6099,N_6275);
nand U7273 (N_7273,N_6309,N_6258);
xnor U7274 (N_7274,N_6698,N_6281);
nand U7275 (N_7275,N_6416,N_6460);
nand U7276 (N_7276,N_6093,N_6482);
xnor U7277 (N_7277,N_6609,N_6682);
nand U7278 (N_7278,N_6008,N_6325);
or U7279 (N_7279,N_6400,N_6120);
nand U7280 (N_7280,N_6745,N_6653);
and U7281 (N_7281,N_6292,N_6354);
nor U7282 (N_7282,N_6627,N_6089);
nand U7283 (N_7283,N_6051,N_6316);
or U7284 (N_7284,N_6471,N_6401);
and U7285 (N_7285,N_6002,N_6435);
and U7286 (N_7286,N_6741,N_6696);
and U7287 (N_7287,N_6285,N_6267);
xor U7288 (N_7288,N_6254,N_6553);
and U7289 (N_7289,N_6399,N_6528);
nor U7290 (N_7290,N_6521,N_6548);
xnor U7291 (N_7291,N_6005,N_6506);
and U7292 (N_7292,N_6434,N_6335);
xnor U7293 (N_7293,N_6051,N_6574);
nor U7294 (N_7294,N_6442,N_6623);
nor U7295 (N_7295,N_6736,N_6365);
nor U7296 (N_7296,N_6727,N_6413);
nand U7297 (N_7297,N_6469,N_6047);
xor U7298 (N_7298,N_6530,N_6337);
and U7299 (N_7299,N_6088,N_6670);
or U7300 (N_7300,N_6295,N_6061);
nor U7301 (N_7301,N_6045,N_6604);
or U7302 (N_7302,N_6284,N_6084);
and U7303 (N_7303,N_6132,N_6103);
nor U7304 (N_7304,N_6407,N_6326);
xnor U7305 (N_7305,N_6660,N_6639);
and U7306 (N_7306,N_6293,N_6449);
and U7307 (N_7307,N_6489,N_6234);
xor U7308 (N_7308,N_6615,N_6377);
and U7309 (N_7309,N_6559,N_6497);
nand U7310 (N_7310,N_6716,N_6360);
or U7311 (N_7311,N_6037,N_6068);
nand U7312 (N_7312,N_6296,N_6577);
nand U7313 (N_7313,N_6595,N_6333);
nor U7314 (N_7314,N_6267,N_6374);
or U7315 (N_7315,N_6643,N_6402);
nand U7316 (N_7316,N_6540,N_6198);
nor U7317 (N_7317,N_6316,N_6389);
and U7318 (N_7318,N_6061,N_6348);
nor U7319 (N_7319,N_6295,N_6531);
nor U7320 (N_7320,N_6026,N_6136);
and U7321 (N_7321,N_6111,N_6208);
xor U7322 (N_7322,N_6505,N_6543);
xor U7323 (N_7323,N_6646,N_6534);
or U7324 (N_7324,N_6172,N_6583);
or U7325 (N_7325,N_6346,N_6106);
nand U7326 (N_7326,N_6213,N_6578);
xor U7327 (N_7327,N_6741,N_6309);
nand U7328 (N_7328,N_6362,N_6653);
xnor U7329 (N_7329,N_6110,N_6732);
nor U7330 (N_7330,N_6133,N_6735);
xnor U7331 (N_7331,N_6677,N_6457);
and U7332 (N_7332,N_6209,N_6701);
nand U7333 (N_7333,N_6714,N_6596);
and U7334 (N_7334,N_6374,N_6499);
and U7335 (N_7335,N_6503,N_6420);
xnor U7336 (N_7336,N_6073,N_6032);
nand U7337 (N_7337,N_6580,N_6320);
nor U7338 (N_7338,N_6091,N_6036);
or U7339 (N_7339,N_6643,N_6099);
nand U7340 (N_7340,N_6734,N_6582);
or U7341 (N_7341,N_6247,N_6180);
xor U7342 (N_7342,N_6250,N_6215);
xor U7343 (N_7343,N_6519,N_6402);
and U7344 (N_7344,N_6601,N_6546);
nor U7345 (N_7345,N_6734,N_6175);
and U7346 (N_7346,N_6660,N_6178);
nor U7347 (N_7347,N_6545,N_6639);
xnor U7348 (N_7348,N_6546,N_6292);
nor U7349 (N_7349,N_6548,N_6535);
nor U7350 (N_7350,N_6462,N_6055);
xor U7351 (N_7351,N_6019,N_6133);
and U7352 (N_7352,N_6618,N_6711);
and U7353 (N_7353,N_6532,N_6060);
or U7354 (N_7354,N_6281,N_6213);
nor U7355 (N_7355,N_6291,N_6232);
xor U7356 (N_7356,N_6355,N_6128);
nand U7357 (N_7357,N_6261,N_6500);
or U7358 (N_7358,N_6603,N_6439);
nor U7359 (N_7359,N_6403,N_6179);
xor U7360 (N_7360,N_6626,N_6128);
xnor U7361 (N_7361,N_6117,N_6204);
and U7362 (N_7362,N_6576,N_6182);
and U7363 (N_7363,N_6328,N_6558);
and U7364 (N_7364,N_6679,N_6626);
nand U7365 (N_7365,N_6051,N_6689);
nand U7366 (N_7366,N_6221,N_6464);
or U7367 (N_7367,N_6603,N_6007);
nor U7368 (N_7368,N_6365,N_6443);
nor U7369 (N_7369,N_6284,N_6302);
nand U7370 (N_7370,N_6717,N_6274);
or U7371 (N_7371,N_6457,N_6595);
xor U7372 (N_7372,N_6522,N_6265);
xor U7373 (N_7373,N_6096,N_6419);
xor U7374 (N_7374,N_6412,N_6047);
nand U7375 (N_7375,N_6621,N_6633);
or U7376 (N_7376,N_6574,N_6077);
xnor U7377 (N_7377,N_6209,N_6511);
xnor U7378 (N_7378,N_6727,N_6478);
nor U7379 (N_7379,N_6315,N_6677);
nand U7380 (N_7380,N_6716,N_6061);
nand U7381 (N_7381,N_6421,N_6295);
nand U7382 (N_7382,N_6151,N_6136);
and U7383 (N_7383,N_6727,N_6635);
nand U7384 (N_7384,N_6252,N_6690);
nor U7385 (N_7385,N_6615,N_6306);
xor U7386 (N_7386,N_6669,N_6360);
and U7387 (N_7387,N_6671,N_6706);
xor U7388 (N_7388,N_6204,N_6416);
nand U7389 (N_7389,N_6216,N_6377);
xnor U7390 (N_7390,N_6247,N_6432);
and U7391 (N_7391,N_6501,N_6280);
xnor U7392 (N_7392,N_6434,N_6263);
or U7393 (N_7393,N_6219,N_6001);
xor U7394 (N_7394,N_6171,N_6052);
xor U7395 (N_7395,N_6218,N_6312);
nor U7396 (N_7396,N_6185,N_6214);
nor U7397 (N_7397,N_6424,N_6376);
or U7398 (N_7398,N_6408,N_6305);
and U7399 (N_7399,N_6393,N_6297);
and U7400 (N_7400,N_6065,N_6558);
nor U7401 (N_7401,N_6114,N_6197);
or U7402 (N_7402,N_6729,N_6382);
or U7403 (N_7403,N_6533,N_6294);
xor U7404 (N_7404,N_6368,N_6167);
xnor U7405 (N_7405,N_6412,N_6749);
nor U7406 (N_7406,N_6189,N_6546);
and U7407 (N_7407,N_6205,N_6569);
nand U7408 (N_7408,N_6012,N_6117);
xor U7409 (N_7409,N_6475,N_6385);
or U7410 (N_7410,N_6637,N_6255);
nand U7411 (N_7411,N_6477,N_6469);
nor U7412 (N_7412,N_6521,N_6016);
nand U7413 (N_7413,N_6245,N_6633);
and U7414 (N_7414,N_6395,N_6662);
or U7415 (N_7415,N_6336,N_6552);
xor U7416 (N_7416,N_6563,N_6543);
nand U7417 (N_7417,N_6443,N_6461);
nor U7418 (N_7418,N_6198,N_6360);
and U7419 (N_7419,N_6386,N_6189);
nor U7420 (N_7420,N_6672,N_6744);
and U7421 (N_7421,N_6610,N_6403);
nor U7422 (N_7422,N_6341,N_6535);
and U7423 (N_7423,N_6582,N_6151);
xnor U7424 (N_7424,N_6679,N_6499);
nor U7425 (N_7425,N_6279,N_6677);
nor U7426 (N_7426,N_6403,N_6031);
nor U7427 (N_7427,N_6152,N_6340);
or U7428 (N_7428,N_6044,N_6615);
and U7429 (N_7429,N_6027,N_6224);
nand U7430 (N_7430,N_6480,N_6104);
nor U7431 (N_7431,N_6223,N_6032);
nand U7432 (N_7432,N_6479,N_6579);
or U7433 (N_7433,N_6133,N_6731);
or U7434 (N_7434,N_6235,N_6022);
and U7435 (N_7435,N_6362,N_6548);
or U7436 (N_7436,N_6668,N_6648);
xnor U7437 (N_7437,N_6378,N_6113);
nand U7438 (N_7438,N_6215,N_6219);
nor U7439 (N_7439,N_6021,N_6031);
nand U7440 (N_7440,N_6170,N_6485);
and U7441 (N_7441,N_6295,N_6680);
or U7442 (N_7442,N_6252,N_6626);
and U7443 (N_7443,N_6669,N_6280);
nand U7444 (N_7444,N_6096,N_6744);
or U7445 (N_7445,N_6204,N_6470);
xor U7446 (N_7446,N_6748,N_6471);
and U7447 (N_7447,N_6362,N_6506);
xor U7448 (N_7448,N_6073,N_6573);
nor U7449 (N_7449,N_6409,N_6034);
or U7450 (N_7450,N_6342,N_6398);
nand U7451 (N_7451,N_6457,N_6052);
or U7452 (N_7452,N_6294,N_6692);
nand U7453 (N_7453,N_6245,N_6499);
nand U7454 (N_7454,N_6345,N_6666);
nand U7455 (N_7455,N_6471,N_6615);
nand U7456 (N_7456,N_6111,N_6706);
or U7457 (N_7457,N_6407,N_6404);
or U7458 (N_7458,N_6302,N_6219);
nand U7459 (N_7459,N_6238,N_6740);
and U7460 (N_7460,N_6422,N_6499);
nand U7461 (N_7461,N_6556,N_6452);
nand U7462 (N_7462,N_6294,N_6437);
xnor U7463 (N_7463,N_6587,N_6217);
or U7464 (N_7464,N_6331,N_6171);
nor U7465 (N_7465,N_6065,N_6582);
nand U7466 (N_7466,N_6471,N_6550);
and U7467 (N_7467,N_6671,N_6470);
or U7468 (N_7468,N_6524,N_6298);
nor U7469 (N_7469,N_6073,N_6436);
or U7470 (N_7470,N_6604,N_6509);
nand U7471 (N_7471,N_6369,N_6079);
nand U7472 (N_7472,N_6376,N_6487);
or U7473 (N_7473,N_6042,N_6269);
and U7474 (N_7474,N_6353,N_6472);
xor U7475 (N_7475,N_6202,N_6512);
or U7476 (N_7476,N_6690,N_6375);
nor U7477 (N_7477,N_6573,N_6140);
nand U7478 (N_7478,N_6283,N_6394);
nand U7479 (N_7479,N_6214,N_6641);
nand U7480 (N_7480,N_6575,N_6112);
or U7481 (N_7481,N_6435,N_6042);
nand U7482 (N_7482,N_6419,N_6205);
or U7483 (N_7483,N_6435,N_6068);
nor U7484 (N_7484,N_6229,N_6743);
nand U7485 (N_7485,N_6397,N_6376);
or U7486 (N_7486,N_6255,N_6731);
and U7487 (N_7487,N_6074,N_6427);
and U7488 (N_7488,N_6554,N_6004);
and U7489 (N_7489,N_6068,N_6344);
nor U7490 (N_7490,N_6408,N_6446);
and U7491 (N_7491,N_6575,N_6680);
nand U7492 (N_7492,N_6275,N_6131);
nor U7493 (N_7493,N_6314,N_6406);
or U7494 (N_7494,N_6031,N_6602);
nor U7495 (N_7495,N_6250,N_6565);
or U7496 (N_7496,N_6722,N_6716);
nor U7497 (N_7497,N_6092,N_6283);
nand U7498 (N_7498,N_6331,N_6261);
nor U7499 (N_7499,N_6562,N_6370);
nor U7500 (N_7500,N_7128,N_7143);
xnor U7501 (N_7501,N_7482,N_7302);
and U7502 (N_7502,N_7353,N_7154);
xor U7503 (N_7503,N_7312,N_6990);
nand U7504 (N_7504,N_7110,N_6885);
or U7505 (N_7505,N_7291,N_7084);
or U7506 (N_7506,N_7308,N_7321);
nand U7507 (N_7507,N_7034,N_6894);
and U7508 (N_7508,N_6944,N_7421);
nor U7509 (N_7509,N_6821,N_7236);
and U7510 (N_7510,N_6959,N_7419);
nor U7511 (N_7511,N_7495,N_6788);
nand U7512 (N_7512,N_7371,N_6785);
nor U7513 (N_7513,N_7455,N_7422);
or U7514 (N_7514,N_6943,N_7095);
and U7515 (N_7515,N_7314,N_6983);
xnor U7516 (N_7516,N_7377,N_6856);
or U7517 (N_7517,N_7113,N_6763);
nor U7518 (N_7518,N_7465,N_7029);
xnor U7519 (N_7519,N_7165,N_7124);
nor U7520 (N_7520,N_6799,N_6797);
or U7521 (N_7521,N_7105,N_7187);
or U7522 (N_7522,N_7348,N_7116);
xor U7523 (N_7523,N_6978,N_7394);
nand U7524 (N_7524,N_7446,N_7013);
nor U7525 (N_7525,N_7266,N_7259);
nor U7526 (N_7526,N_6964,N_7052);
nand U7527 (N_7527,N_7317,N_6813);
xor U7528 (N_7528,N_6926,N_6918);
nand U7529 (N_7529,N_6792,N_7180);
xor U7530 (N_7530,N_7145,N_6776);
and U7531 (N_7531,N_6778,N_7218);
and U7532 (N_7532,N_7020,N_6989);
and U7533 (N_7533,N_7149,N_6857);
nand U7534 (N_7534,N_7347,N_7359);
xnor U7535 (N_7535,N_6979,N_7466);
nor U7536 (N_7536,N_7192,N_6953);
nor U7537 (N_7537,N_7489,N_7063);
xnor U7538 (N_7538,N_7244,N_7204);
nor U7539 (N_7539,N_6909,N_6787);
nand U7540 (N_7540,N_6817,N_7431);
nor U7541 (N_7541,N_7185,N_7329);
xnor U7542 (N_7542,N_7328,N_7173);
nor U7543 (N_7543,N_6951,N_7332);
nand U7544 (N_7544,N_6958,N_6783);
nor U7545 (N_7545,N_7471,N_7033);
xor U7546 (N_7546,N_7207,N_7158);
and U7547 (N_7547,N_7378,N_7086);
nor U7548 (N_7548,N_7415,N_7282);
or U7549 (N_7549,N_7385,N_7146);
xor U7550 (N_7550,N_7433,N_7475);
nor U7551 (N_7551,N_6831,N_7133);
and U7552 (N_7552,N_7309,N_7358);
nor U7553 (N_7553,N_6931,N_7074);
nand U7554 (N_7554,N_7168,N_7243);
nor U7555 (N_7555,N_6846,N_7252);
or U7556 (N_7556,N_6955,N_7093);
or U7557 (N_7557,N_6830,N_7193);
nand U7558 (N_7558,N_7306,N_7324);
nand U7559 (N_7559,N_7337,N_7088);
nand U7560 (N_7560,N_7384,N_6913);
and U7561 (N_7561,N_7191,N_7281);
xnor U7562 (N_7562,N_7101,N_6832);
nor U7563 (N_7563,N_7258,N_7263);
nand U7564 (N_7564,N_6908,N_6858);
and U7565 (N_7565,N_7229,N_7411);
nor U7566 (N_7566,N_7225,N_7190);
and U7567 (N_7567,N_7226,N_7296);
and U7568 (N_7568,N_6991,N_7094);
nand U7569 (N_7569,N_7138,N_7107);
or U7570 (N_7570,N_7355,N_7099);
nor U7571 (N_7571,N_7026,N_6896);
and U7572 (N_7572,N_7071,N_7183);
nor U7573 (N_7573,N_7249,N_7382);
or U7574 (N_7574,N_7188,N_7174);
and U7575 (N_7575,N_7399,N_7051);
nand U7576 (N_7576,N_6782,N_6756);
nand U7577 (N_7577,N_7125,N_7354);
nand U7578 (N_7578,N_7268,N_7132);
nor U7579 (N_7579,N_7469,N_6891);
xor U7580 (N_7580,N_7025,N_7265);
and U7581 (N_7581,N_7301,N_7120);
and U7582 (N_7582,N_7459,N_6864);
and U7583 (N_7583,N_6867,N_6895);
xor U7584 (N_7584,N_6934,N_7460);
and U7585 (N_7585,N_7290,N_7420);
nand U7586 (N_7586,N_7085,N_6942);
or U7587 (N_7587,N_7041,N_6967);
xor U7588 (N_7588,N_7269,N_7136);
or U7589 (N_7589,N_7288,N_7068);
nand U7590 (N_7590,N_7184,N_6923);
and U7591 (N_7591,N_6892,N_7498);
and U7592 (N_7592,N_7260,N_6935);
and U7593 (N_7593,N_7059,N_6969);
nand U7594 (N_7594,N_7209,N_7053);
nor U7595 (N_7595,N_7098,N_7346);
or U7596 (N_7596,N_6767,N_7280);
xor U7597 (N_7597,N_6786,N_6835);
and U7598 (N_7598,N_7388,N_7144);
nand U7599 (N_7599,N_7112,N_7039);
or U7600 (N_7600,N_7343,N_6884);
or U7601 (N_7601,N_6876,N_6875);
or U7602 (N_7602,N_7396,N_7267);
or U7603 (N_7603,N_7089,N_7123);
xnor U7604 (N_7604,N_7303,N_7368);
nand U7605 (N_7605,N_7299,N_6865);
xor U7606 (N_7606,N_7040,N_7054);
and U7607 (N_7607,N_6924,N_7151);
and U7608 (N_7608,N_7427,N_7230);
nor U7609 (N_7609,N_7104,N_6781);
or U7610 (N_7610,N_7070,N_7177);
xor U7611 (N_7611,N_7450,N_6998);
xor U7612 (N_7612,N_6780,N_7170);
nand U7613 (N_7613,N_7161,N_6871);
and U7614 (N_7614,N_7087,N_7221);
nand U7615 (N_7615,N_7497,N_7108);
nor U7616 (N_7616,N_7272,N_6950);
xnor U7617 (N_7617,N_7253,N_6771);
and U7618 (N_7618,N_7367,N_7387);
xnor U7619 (N_7619,N_7406,N_7122);
xnor U7620 (N_7620,N_7484,N_6828);
or U7621 (N_7621,N_7076,N_6754);
xor U7622 (N_7622,N_7066,N_7067);
nor U7623 (N_7623,N_7365,N_6842);
or U7624 (N_7624,N_6805,N_7449);
nand U7625 (N_7625,N_7287,N_6854);
and U7626 (N_7626,N_7333,N_7326);
nand U7627 (N_7627,N_7330,N_7492);
or U7628 (N_7628,N_7391,N_6838);
xnor U7629 (N_7629,N_6907,N_6928);
or U7630 (N_7630,N_7235,N_7134);
nor U7631 (N_7631,N_7362,N_6921);
nor U7632 (N_7632,N_6758,N_7380);
nor U7633 (N_7633,N_6889,N_6755);
nand U7634 (N_7634,N_7171,N_7201);
and U7635 (N_7635,N_7486,N_7176);
and U7636 (N_7636,N_7140,N_7247);
xor U7637 (N_7637,N_7361,N_7227);
nand U7638 (N_7638,N_7426,N_6870);
nand U7639 (N_7639,N_7441,N_6766);
and U7640 (N_7640,N_7219,N_7022);
nor U7641 (N_7641,N_7363,N_7445);
or U7642 (N_7642,N_6880,N_6804);
nand U7643 (N_7643,N_7251,N_7157);
nand U7644 (N_7644,N_7454,N_6878);
or U7645 (N_7645,N_7264,N_7091);
xor U7646 (N_7646,N_6966,N_6970);
xor U7647 (N_7647,N_7478,N_7250);
xnor U7648 (N_7648,N_6988,N_6937);
or U7649 (N_7649,N_6903,N_6848);
nor U7650 (N_7650,N_7181,N_7438);
xor U7651 (N_7651,N_6974,N_7077);
nor U7652 (N_7652,N_7083,N_7325);
xor U7653 (N_7653,N_7057,N_6902);
nand U7654 (N_7654,N_7234,N_7163);
nor U7655 (N_7655,N_7414,N_7200);
nor U7656 (N_7656,N_6825,N_7458);
nand U7657 (N_7657,N_6890,N_7019);
xor U7658 (N_7658,N_6794,N_6852);
nand U7659 (N_7659,N_6861,N_6956);
nand U7660 (N_7660,N_7437,N_7480);
or U7661 (N_7661,N_6843,N_6769);
xnor U7662 (N_7662,N_7350,N_6938);
nand U7663 (N_7663,N_6940,N_7389);
nor U7664 (N_7664,N_6985,N_7064);
nor U7665 (N_7665,N_6980,N_6962);
nand U7666 (N_7666,N_7023,N_6922);
nor U7667 (N_7667,N_6936,N_7400);
nand U7668 (N_7668,N_7126,N_7311);
xnor U7669 (N_7669,N_7277,N_7294);
and U7670 (N_7670,N_7494,N_7114);
nand U7671 (N_7671,N_7429,N_6800);
nor U7672 (N_7672,N_6765,N_7404);
or U7673 (N_7673,N_7182,N_6752);
nand U7674 (N_7674,N_6774,N_6806);
xor U7675 (N_7675,N_7351,N_7442);
or U7676 (N_7676,N_7339,N_7295);
or U7677 (N_7677,N_6791,N_6773);
or U7678 (N_7678,N_7405,N_7030);
and U7679 (N_7679,N_6866,N_7049);
or U7680 (N_7680,N_7307,N_6824);
or U7681 (N_7681,N_7255,N_6809);
and U7682 (N_7682,N_7194,N_7135);
nand U7683 (N_7683,N_7100,N_7369);
or U7684 (N_7684,N_7024,N_7018);
xnor U7685 (N_7685,N_7044,N_7476);
nor U7686 (N_7686,N_7440,N_6784);
or U7687 (N_7687,N_7078,N_7357);
and U7688 (N_7688,N_7477,N_7403);
nand U7689 (N_7689,N_7103,N_7042);
nand U7690 (N_7690,N_7461,N_7096);
and U7691 (N_7691,N_7220,N_7313);
and U7692 (N_7692,N_6948,N_7383);
nor U7693 (N_7693,N_6872,N_6883);
xnor U7694 (N_7694,N_7210,N_7416);
or U7695 (N_7695,N_7164,N_7485);
xnor U7696 (N_7696,N_6772,N_7360);
and U7697 (N_7697,N_6977,N_7424);
and U7698 (N_7698,N_6952,N_7334);
nor U7699 (N_7699,N_7257,N_6845);
nand U7700 (N_7700,N_7293,N_7233);
or U7701 (N_7701,N_7046,N_7069);
and U7702 (N_7702,N_7408,N_6963);
nand U7703 (N_7703,N_6789,N_6798);
nand U7704 (N_7704,N_7254,N_7160);
and U7705 (N_7705,N_7242,N_7409);
or U7706 (N_7706,N_7111,N_6897);
nor U7707 (N_7707,N_7016,N_7139);
nand U7708 (N_7708,N_6790,N_6996);
xor U7709 (N_7709,N_7315,N_7496);
or U7710 (N_7710,N_7278,N_6853);
nand U7711 (N_7711,N_7212,N_6834);
nor U7712 (N_7712,N_7276,N_6862);
or U7713 (N_7713,N_6768,N_7331);
nor U7714 (N_7714,N_6973,N_7222);
xnor U7715 (N_7715,N_7004,N_7488);
nand U7716 (N_7716,N_7213,N_6793);
nor U7717 (N_7717,N_6820,N_6911);
and U7718 (N_7718,N_6823,N_7292);
and U7719 (N_7719,N_6987,N_6816);
nor U7720 (N_7720,N_7434,N_7131);
xnor U7721 (N_7721,N_7402,N_6869);
xor U7722 (N_7722,N_7345,N_6919);
or U7723 (N_7723,N_6995,N_7444);
xnor U7724 (N_7724,N_7468,N_6819);
nor U7725 (N_7725,N_6927,N_6912);
and U7726 (N_7726,N_6860,N_7152);
nand U7727 (N_7727,N_7379,N_6982);
and U7728 (N_7728,N_6837,N_7356);
nor U7729 (N_7729,N_6863,N_7055);
or U7730 (N_7730,N_7119,N_7178);
nor U7731 (N_7731,N_7032,N_7027);
nand U7732 (N_7732,N_7453,N_7189);
nand U7733 (N_7733,N_6930,N_6851);
nand U7734 (N_7734,N_7381,N_6920);
or U7735 (N_7735,N_7239,N_6906);
nand U7736 (N_7736,N_6887,N_6900);
nor U7737 (N_7737,N_7109,N_6932);
nand U7738 (N_7738,N_6873,N_7150);
and U7739 (N_7739,N_7467,N_7428);
and U7740 (N_7740,N_7490,N_7447);
xnor U7741 (N_7741,N_6877,N_6992);
nor U7742 (N_7742,N_7375,N_7456);
nand U7743 (N_7743,N_7208,N_6836);
xor U7744 (N_7744,N_7275,N_7092);
and U7745 (N_7745,N_6886,N_7017);
nand U7746 (N_7746,N_7102,N_6779);
nor U7747 (N_7747,N_7240,N_7398);
nand U7748 (N_7748,N_7097,N_7246);
and U7749 (N_7749,N_7197,N_7436);
xnor U7750 (N_7750,N_7432,N_7003);
nand U7751 (N_7751,N_7001,N_7217);
and U7752 (N_7752,N_6847,N_6829);
nand U7753 (N_7753,N_7223,N_7117);
nor U7754 (N_7754,N_6811,N_6925);
and U7755 (N_7755,N_7448,N_7279);
nor U7756 (N_7756,N_7499,N_6947);
or U7757 (N_7757,N_6961,N_7370);
nand U7758 (N_7758,N_7338,N_7142);
xor U7759 (N_7759,N_7021,N_6840);
xnor U7760 (N_7760,N_7155,N_7479);
xnor U7761 (N_7761,N_6917,N_7273);
nor U7762 (N_7762,N_6818,N_7430);
nand U7763 (N_7763,N_7470,N_6762);
xor U7764 (N_7764,N_7386,N_7401);
nor U7765 (N_7765,N_6796,N_6881);
or U7766 (N_7766,N_7079,N_6827);
xnor U7767 (N_7767,N_6975,N_7062);
nand U7768 (N_7768,N_6803,N_7425);
or U7769 (N_7769,N_6957,N_7007);
xnor U7770 (N_7770,N_6888,N_7462);
nand U7771 (N_7771,N_7344,N_7215);
nand U7772 (N_7772,N_7241,N_7153);
nand U7773 (N_7773,N_7452,N_7284);
nor U7774 (N_7774,N_7392,N_6999);
nor U7775 (N_7775,N_7374,N_7127);
and U7776 (N_7776,N_7319,N_7075);
and U7777 (N_7777,N_7349,N_7376);
xnor U7778 (N_7778,N_7310,N_6833);
nand U7779 (N_7779,N_7412,N_7028);
xor U7780 (N_7780,N_7129,N_6753);
or U7781 (N_7781,N_7196,N_7179);
nand U7782 (N_7782,N_7148,N_7245);
nand U7783 (N_7783,N_6826,N_7014);
nand U7784 (N_7784,N_7493,N_7286);
and U7785 (N_7785,N_7336,N_7464);
and U7786 (N_7786,N_7010,N_6849);
or U7787 (N_7787,N_7166,N_7271);
nor U7788 (N_7788,N_7342,N_6984);
or U7789 (N_7789,N_7393,N_7202);
and U7790 (N_7790,N_7335,N_6839);
nor U7791 (N_7791,N_6939,N_6968);
xor U7792 (N_7792,N_7256,N_6814);
and U7793 (N_7793,N_7037,N_6879);
nor U7794 (N_7794,N_7056,N_7372);
or U7795 (N_7795,N_6899,N_6981);
nor U7796 (N_7796,N_7000,N_6960);
nor U7797 (N_7797,N_6764,N_7082);
nor U7798 (N_7798,N_7248,N_7297);
xnor U7799 (N_7799,N_6933,N_7320);
or U7800 (N_7800,N_7011,N_7352);
and U7801 (N_7801,N_7472,N_6822);
nand U7802 (N_7802,N_6976,N_6882);
nor U7803 (N_7803,N_7232,N_7159);
nor U7804 (N_7804,N_6859,N_6915);
nand U7805 (N_7805,N_7130,N_7487);
xor U7806 (N_7806,N_7298,N_7300);
xnor U7807 (N_7807,N_7373,N_7228);
nand U7808 (N_7808,N_7304,N_7006);
nor U7809 (N_7809,N_7121,N_7214);
and U7810 (N_7810,N_6844,N_6905);
nor U7811 (N_7811,N_7061,N_7439);
nand U7812 (N_7812,N_7316,N_6802);
nor U7813 (N_7813,N_7043,N_7366);
nand U7814 (N_7814,N_6971,N_7073);
nor U7815 (N_7815,N_7186,N_7473);
nand U7816 (N_7816,N_7009,N_6904);
xnor U7817 (N_7817,N_7036,N_7048);
nand U7818 (N_7818,N_7118,N_7457);
xor U7819 (N_7819,N_6807,N_7397);
and U7820 (N_7820,N_7169,N_7015);
nor U7821 (N_7821,N_7072,N_7491);
and U7822 (N_7822,N_7008,N_7318);
nor U7823 (N_7823,N_7141,N_7322);
nor U7824 (N_7824,N_7172,N_7224);
nand U7825 (N_7825,N_7012,N_7407);
nor U7826 (N_7826,N_7364,N_7203);
and U7827 (N_7827,N_7060,N_6777);
or U7828 (N_7828,N_6751,N_6757);
nor U7829 (N_7829,N_6815,N_6795);
nand U7830 (N_7830,N_7305,N_7047);
xnor U7831 (N_7831,N_7090,N_6914);
or U7832 (N_7832,N_6946,N_7065);
xnor U7833 (N_7833,N_6901,N_7261);
nor U7834 (N_7834,N_7395,N_7106);
or U7835 (N_7835,N_6850,N_6898);
xnor U7836 (N_7836,N_6759,N_6910);
nand U7837 (N_7837,N_7002,N_7031);
and U7838 (N_7838,N_7481,N_6949);
xnor U7839 (N_7839,N_6810,N_7038);
nor U7840 (N_7840,N_6893,N_7390);
nand U7841 (N_7841,N_6868,N_7115);
and U7842 (N_7842,N_7289,N_6855);
and U7843 (N_7843,N_7418,N_7156);
or U7844 (N_7844,N_7274,N_6808);
and U7845 (N_7845,N_7199,N_7327);
nor U7846 (N_7846,N_7206,N_7483);
nor U7847 (N_7847,N_7045,N_6965);
or U7848 (N_7848,N_6954,N_7283);
nor U7849 (N_7849,N_6993,N_7058);
nor U7850 (N_7850,N_6760,N_6874);
xnor U7851 (N_7851,N_7463,N_7080);
xor U7852 (N_7852,N_7341,N_6997);
nand U7853 (N_7853,N_7423,N_7237);
or U7854 (N_7854,N_6761,N_7005);
nor U7855 (N_7855,N_6972,N_6770);
and U7856 (N_7856,N_7323,N_7451);
xnor U7857 (N_7857,N_6775,N_7081);
nor U7858 (N_7858,N_7050,N_7262);
or U7859 (N_7859,N_7162,N_6986);
and U7860 (N_7860,N_7216,N_7211);
xor U7861 (N_7861,N_6916,N_7285);
nand U7862 (N_7862,N_6812,N_6994);
nor U7863 (N_7863,N_7035,N_7238);
nor U7864 (N_7864,N_6929,N_7413);
or U7865 (N_7865,N_7137,N_7340);
xor U7866 (N_7866,N_6941,N_7198);
xor U7867 (N_7867,N_7175,N_6801);
xor U7868 (N_7868,N_7147,N_7417);
xnor U7869 (N_7869,N_6945,N_7443);
nor U7870 (N_7870,N_7270,N_7205);
nand U7871 (N_7871,N_6750,N_7195);
nand U7872 (N_7872,N_7231,N_7474);
and U7873 (N_7873,N_7410,N_7435);
nand U7874 (N_7874,N_7167,N_6841);
xor U7875 (N_7875,N_7183,N_7331);
and U7876 (N_7876,N_7148,N_7141);
or U7877 (N_7877,N_6788,N_7475);
xor U7878 (N_7878,N_6857,N_6954);
xnor U7879 (N_7879,N_6819,N_7088);
xnor U7880 (N_7880,N_7019,N_7370);
and U7881 (N_7881,N_7470,N_7444);
nor U7882 (N_7882,N_7350,N_7147);
or U7883 (N_7883,N_7341,N_7162);
and U7884 (N_7884,N_7036,N_7044);
or U7885 (N_7885,N_7240,N_7354);
xnor U7886 (N_7886,N_7155,N_7190);
xnor U7887 (N_7887,N_6772,N_7421);
xnor U7888 (N_7888,N_7048,N_7356);
or U7889 (N_7889,N_7103,N_7218);
nand U7890 (N_7890,N_6779,N_7013);
or U7891 (N_7891,N_6758,N_7149);
xnor U7892 (N_7892,N_7228,N_6952);
nand U7893 (N_7893,N_6937,N_7485);
or U7894 (N_7894,N_7001,N_7411);
or U7895 (N_7895,N_6782,N_7297);
xnor U7896 (N_7896,N_7249,N_6933);
xor U7897 (N_7897,N_6823,N_7103);
xor U7898 (N_7898,N_6847,N_7121);
or U7899 (N_7899,N_7030,N_6812);
xnor U7900 (N_7900,N_7255,N_6815);
nor U7901 (N_7901,N_7146,N_6980);
xnor U7902 (N_7902,N_7119,N_6797);
and U7903 (N_7903,N_6902,N_7463);
nand U7904 (N_7904,N_6954,N_7322);
and U7905 (N_7905,N_7072,N_7302);
nand U7906 (N_7906,N_7033,N_7288);
or U7907 (N_7907,N_6818,N_7112);
or U7908 (N_7908,N_7382,N_6937);
nor U7909 (N_7909,N_7377,N_7170);
and U7910 (N_7910,N_6918,N_7339);
nand U7911 (N_7911,N_6979,N_7438);
nor U7912 (N_7912,N_7454,N_7350);
xnor U7913 (N_7913,N_7283,N_7128);
xnor U7914 (N_7914,N_6974,N_7177);
or U7915 (N_7915,N_7493,N_7105);
nor U7916 (N_7916,N_7094,N_7009);
xor U7917 (N_7917,N_7153,N_7268);
nand U7918 (N_7918,N_6949,N_7228);
and U7919 (N_7919,N_7397,N_7024);
xnor U7920 (N_7920,N_7146,N_6922);
nand U7921 (N_7921,N_7469,N_6933);
or U7922 (N_7922,N_6910,N_7143);
and U7923 (N_7923,N_6897,N_7303);
nor U7924 (N_7924,N_7018,N_7308);
and U7925 (N_7925,N_6961,N_7264);
or U7926 (N_7926,N_7349,N_7313);
xor U7927 (N_7927,N_7030,N_6929);
nor U7928 (N_7928,N_7327,N_6873);
and U7929 (N_7929,N_6825,N_7340);
or U7930 (N_7930,N_7115,N_6810);
nor U7931 (N_7931,N_6906,N_6931);
nand U7932 (N_7932,N_7323,N_7147);
and U7933 (N_7933,N_7254,N_7065);
xor U7934 (N_7934,N_6788,N_6995);
and U7935 (N_7935,N_7137,N_7219);
nand U7936 (N_7936,N_7197,N_7131);
or U7937 (N_7937,N_6972,N_7042);
and U7938 (N_7938,N_6996,N_7390);
and U7939 (N_7939,N_7232,N_6828);
nor U7940 (N_7940,N_6778,N_7117);
xnor U7941 (N_7941,N_6825,N_7491);
nand U7942 (N_7942,N_7369,N_7011);
nor U7943 (N_7943,N_7143,N_7469);
or U7944 (N_7944,N_7331,N_7365);
xnor U7945 (N_7945,N_7358,N_6958);
nand U7946 (N_7946,N_7496,N_7475);
or U7947 (N_7947,N_7153,N_6757);
nand U7948 (N_7948,N_7014,N_6750);
and U7949 (N_7949,N_7205,N_7289);
nand U7950 (N_7950,N_7481,N_7245);
xnor U7951 (N_7951,N_7237,N_7129);
nand U7952 (N_7952,N_7256,N_7322);
and U7953 (N_7953,N_7262,N_7013);
nand U7954 (N_7954,N_7456,N_6904);
and U7955 (N_7955,N_7013,N_7040);
xor U7956 (N_7956,N_7290,N_7067);
nor U7957 (N_7957,N_7059,N_7388);
or U7958 (N_7958,N_7113,N_7368);
nand U7959 (N_7959,N_7387,N_6847);
xor U7960 (N_7960,N_7470,N_6881);
and U7961 (N_7961,N_6764,N_7447);
xnor U7962 (N_7962,N_6944,N_7477);
nor U7963 (N_7963,N_6933,N_6949);
nand U7964 (N_7964,N_7369,N_7496);
xnor U7965 (N_7965,N_7219,N_6877);
xor U7966 (N_7966,N_7309,N_6977);
or U7967 (N_7967,N_7258,N_7159);
and U7968 (N_7968,N_7031,N_7238);
and U7969 (N_7969,N_6997,N_7307);
nand U7970 (N_7970,N_7275,N_7324);
or U7971 (N_7971,N_6994,N_7457);
nor U7972 (N_7972,N_7032,N_7117);
or U7973 (N_7973,N_7310,N_7383);
or U7974 (N_7974,N_6797,N_7219);
nor U7975 (N_7975,N_7035,N_6870);
or U7976 (N_7976,N_6976,N_7353);
or U7977 (N_7977,N_6790,N_7217);
and U7978 (N_7978,N_7331,N_7085);
xnor U7979 (N_7979,N_6991,N_7300);
nor U7980 (N_7980,N_7286,N_7360);
nand U7981 (N_7981,N_7138,N_6953);
and U7982 (N_7982,N_6860,N_7193);
and U7983 (N_7983,N_6829,N_6919);
nor U7984 (N_7984,N_6839,N_6870);
nand U7985 (N_7985,N_7360,N_6920);
or U7986 (N_7986,N_6773,N_7455);
nor U7987 (N_7987,N_7475,N_6923);
nor U7988 (N_7988,N_6808,N_6805);
nand U7989 (N_7989,N_7467,N_6803);
or U7990 (N_7990,N_7091,N_7499);
nand U7991 (N_7991,N_6787,N_6911);
or U7992 (N_7992,N_7194,N_7211);
and U7993 (N_7993,N_7015,N_7337);
nor U7994 (N_7994,N_7209,N_7173);
or U7995 (N_7995,N_6788,N_7062);
or U7996 (N_7996,N_6875,N_7219);
and U7997 (N_7997,N_7493,N_7166);
and U7998 (N_7998,N_6950,N_6782);
nor U7999 (N_7999,N_6840,N_6849);
or U8000 (N_8000,N_7031,N_7130);
nor U8001 (N_8001,N_7358,N_7429);
and U8002 (N_8002,N_6756,N_7094);
and U8003 (N_8003,N_6787,N_7463);
nand U8004 (N_8004,N_6933,N_6961);
xnor U8005 (N_8005,N_6993,N_7321);
xor U8006 (N_8006,N_6800,N_7337);
nor U8007 (N_8007,N_7484,N_7196);
and U8008 (N_8008,N_6788,N_7155);
nand U8009 (N_8009,N_7360,N_7494);
nor U8010 (N_8010,N_7493,N_6768);
or U8011 (N_8011,N_7092,N_6811);
and U8012 (N_8012,N_7273,N_6816);
nand U8013 (N_8013,N_7180,N_7158);
and U8014 (N_8014,N_7035,N_7348);
nor U8015 (N_8015,N_7361,N_7490);
or U8016 (N_8016,N_7049,N_7079);
or U8017 (N_8017,N_6772,N_7358);
and U8018 (N_8018,N_7208,N_6843);
and U8019 (N_8019,N_7225,N_7099);
nor U8020 (N_8020,N_6879,N_7299);
nand U8021 (N_8021,N_7304,N_7050);
nor U8022 (N_8022,N_6905,N_7387);
nand U8023 (N_8023,N_7408,N_7482);
nor U8024 (N_8024,N_7262,N_7191);
or U8025 (N_8025,N_7102,N_7004);
and U8026 (N_8026,N_7369,N_6983);
and U8027 (N_8027,N_7331,N_6797);
nand U8028 (N_8028,N_7027,N_6956);
nor U8029 (N_8029,N_7314,N_7046);
nor U8030 (N_8030,N_6967,N_7023);
or U8031 (N_8031,N_6880,N_7059);
xnor U8032 (N_8032,N_6987,N_7079);
and U8033 (N_8033,N_7298,N_7092);
and U8034 (N_8034,N_7307,N_6835);
or U8035 (N_8035,N_7204,N_7073);
nand U8036 (N_8036,N_7215,N_7290);
or U8037 (N_8037,N_7181,N_6974);
xor U8038 (N_8038,N_7120,N_6991);
xor U8039 (N_8039,N_7450,N_6863);
xor U8040 (N_8040,N_6818,N_6996);
or U8041 (N_8041,N_7249,N_6976);
nand U8042 (N_8042,N_6903,N_7033);
or U8043 (N_8043,N_6751,N_6896);
nor U8044 (N_8044,N_7351,N_7445);
nor U8045 (N_8045,N_7327,N_7418);
or U8046 (N_8046,N_6914,N_7107);
or U8047 (N_8047,N_6753,N_7104);
nand U8048 (N_8048,N_6957,N_7173);
and U8049 (N_8049,N_7092,N_6813);
nand U8050 (N_8050,N_7441,N_7273);
xor U8051 (N_8051,N_7487,N_7442);
nand U8052 (N_8052,N_6773,N_7352);
xnor U8053 (N_8053,N_6840,N_7130);
xnor U8054 (N_8054,N_7260,N_7307);
nand U8055 (N_8055,N_7345,N_6942);
nand U8056 (N_8056,N_7236,N_6974);
nand U8057 (N_8057,N_6818,N_7120);
and U8058 (N_8058,N_7159,N_6937);
and U8059 (N_8059,N_7331,N_6791);
nand U8060 (N_8060,N_7460,N_7074);
xnor U8061 (N_8061,N_6977,N_7482);
xor U8062 (N_8062,N_6978,N_6945);
xor U8063 (N_8063,N_7058,N_7405);
nand U8064 (N_8064,N_7306,N_6955);
nand U8065 (N_8065,N_7424,N_7472);
or U8066 (N_8066,N_6882,N_6941);
xnor U8067 (N_8067,N_7200,N_7190);
nor U8068 (N_8068,N_7145,N_7259);
xor U8069 (N_8069,N_7378,N_7209);
xnor U8070 (N_8070,N_7339,N_7287);
nor U8071 (N_8071,N_7189,N_7138);
nor U8072 (N_8072,N_6913,N_6952);
xor U8073 (N_8073,N_6761,N_6860);
and U8074 (N_8074,N_7496,N_6752);
nor U8075 (N_8075,N_6770,N_7188);
or U8076 (N_8076,N_7165,N_7299);
nand U8077 (N_8077,N_7270,N_7002);
nand U8078 (N_8078,N_6958,N_7218);
nor U8079 (N_8079,N_7379,N_7007);
nand U8080 (N_8080,N_7332,N_7360);
and U8081 (N_8081,N_6858,N_7456);
and U8082 (N_8082,N_7337,N_6854);
nand U8083 (N_8083,N_7488,N_6867);
or U8084 (N_8084,N_6762,N_6893);
and U8085 (N_8085,N_7148,N_7191);
xor U8086 (N_8086,N_7313,N_7414);
xor U8087 (N_8087,N_6907,N_6798);
xnor U8088 (N_8088,N_6913,N_6897);
nor U8089 (N_8089,N_7005,N_7149);
nand U8090 (N_8090,N_7461,N_7273);
nand U8091 (N_8091,N_7203,N_6898);
nor U8092 (N_8092,N_7121,N_6801);
xnor U8093 (N_8093,N_7138,N_7417);
and U8094 (N_8094,N_7010,N_7171);
or U8095 (N_8095,N_6847,N_7200);
or U8096 (N_8096,N_7404,N_7167);
xnor U8097 (N_8097,N_7166,N_6874);
nor U8098 (N_8098,N_7157,N_6792);
or U8099 (N_8099,N_7267,N_6799);
nand U8100 (N_8100,N_6842,N_7480);
nor U8101 (N_8101,N_7223,N_6895);
nand U8102 (N_8102,N_7315,N_6778);
xnor U8103 (N_8103,N_7241,N_7222);
and U8104 (N_8104,N_7051,N_7230);
nor U8105 (N_8105,N_6779,N_7251);
or U8106 (N_8106,N_6762,N_7265);
and U8107 (N_8107,N_7187,N_6795);
nor U8108 (N_8108,N_7405,N_7027);
nor U8109 (N_8109,N_7368,N_7103);
xnor U8110 (N_8110,N_6864,N_7377);
nor U8111 (N_8111,N_7190,N_7240);
nor U8112 (N_8112,N_6884,N_6760);
xnor U8113 (N_8113,N_7048,N_7187);
nor U8114 (N_8114,N_7221,N_6860);
nand U8115 (N_8115,N_6756,N_7213);
nand U8116 (N_8116,N_6871,N_7033);
nand U8117 (N_8117,N_6847,N_7331);
xnor U8118 (N_8118,N_7015,N_7298);
and U8119 (N_8119,N_7058,N_7346);
xor U8120 (N_8120,N_7164,N_6826);
xnor U8121 (N_8121,N_7289,N_6802);
nand U8122 (N_8122,N_7405,N_6992);
xnor U8123 (N_8123,N_7483,N_6892);
nand U8124 (N_8124,N_7429,N_7371);
or U8125 (N_8125,N_6848,N_7446);
and U8126 (N_8126,N_7475,N_6934);
and U8127 (N_8127,N_7297,N_6903);
nand U8128 (N_8128,N_7106,N_6825);
nand U8129 (N_8129,N_7441,N_6901);
nand U8130 (N_8130,N_7360,N_6895);
and U8131 (N_8131,N_6955,N_7290);
and U8132 (N_8132,N_6922,N_7422);
xor U8133 (N_8133,N_7310,N_7381);
or U8134 (N_8134,N_6941,N_6872);
or U8135 (N_8135,N_7196,N_7174);
xor U8136 (N_8136,N_6791,N_7144);
xnor U8137 (N_8137,N_6844,N_7430);
and U8138 (N_8138,N_6785,N_7369);
xor U8139 (N_8139,N_7408,N_6965);
nand U8140 (N_8140,N_6750,N_6828);
nand U8141 (N_8141,N_6845,N_6911);
xor U8142 (N_8142,N_7045,N_6987);
and U8143 (N_8143,N_6818,N_7010);
nand U8144 (N_8144,N_7388,N_7051);
and U8145 (N_8145,N_6846,N_7136);
and U8146 (N_8146,N_7143,N_7026);
and U8147 (N_8147,N_7378,N_6977);
or U8148 (N_8148,N_7095,N_7482);
xnor U8149 (N_8149,N_6833,N_7030);
and U8150 (N_8150,N_7007,N_7437);
and U8151 (N_8151,N_6926,N_6988);
xor U8152 (N_8152,N_7183,N_7185);
and U8153 (N_8153,N_7434,N_7127);
nor U8154 (N_8154,N_7499,N_7051);
nand U8155 (N_8155,N_7037,N_6793);
nand U8156 (N_8156,N_7410,N_7497);
and U8157 (N_8157,N_7448,N_6825);
or U8158 (N_8158,N_7343,N_6961);
nand U8159 (N_8159,N_7111,N_7154);
and U8160 (N_8160,N_6973,N_7399);
and U8161 (N_8161,N_7216,N_6781);
nor U8162 (N_8162,N_6778,N_7489);
xor U8163 (N_8163,N_6828,N_6790);
and U8164 (N_8164,N_6997,N_7338);
or U8165 (N_8165,N_6995,N_6987);
nand U8166 (N_8166,N_6797,N_7036);
nor U8167 (N_8167,N_7276,N_6949);
or U8168 (N_8168,N_7246,N_7031);
and U8169 (N_8169,N_7171,N_6848);
nor U8170 (N_8170,N_7489,N_6851);
nor U8171 (N_8171,N_7059,N_6876);
nand U8172 (N_8172,N_7120,N_7041);
or U8173 (N_8173,N_6979,N_7259);
xor U8174 (N_8174,N_6879,N_6983);
or U8175 (N_8175,N_7257,N_7162);
xnor U8176 (N_8176,N_6761,N_6807);
nor U8177 (N_8177,N_7267,N_7400);
nor U8178 (N_8178,N_7090,N_7212);
and U8179 (N_8179,N_7083,N_7351);
and U8180 (N_8180,N_7214,N_7261);
and U8181 (N_8181,N_6771,N_6925);
nor U8182 (N_8182,N_7088,N_7065);
nand U8183 (N_8183,N_7437,N_7040);
and U8184 (N_8184,N_7289,N_7086);
nand U8185 (N_8185,N_6989,N_7036);
nand U8186 (N_8186,N_6913,N_6934);
nand U8187 (N_8187,N_6880,N_7106);
xnor U8188 (N_8188,N_6809,N_7041);
nand U8189 (N_8189,N_7297,N_7339);
nand U8190 (N_8190,N_7265,N_7088);
xor U8191 (N_8191,N_7126,N_6825);
nor U8192 (N_8192,N_7421,N_7151);
or U8193 (N_8193,N_7468,N_7296);
and U8194 (N_8194,N_7126,N_6753);
nor U8195 (N_8195,N_7368,N_6793);
or U8196 (N_8196,N_6761,N_6850);
nand U8197 (N_8197,N_7298,N_7430);
and U8198 (N_8198,N_7013,N_7081);
and U8199 (N_8199,N_7023,N_7480);
nand U8200 (N_8200,N_7034,N_6975);
nor U8201 (N_8201,N_7426,N_7276);
nand U8202 (N_8202,N_7428,N_7204);
nor U8203 (N_8203,N_6975,N_7383);
or U8204 (N_8204,N_7111,N_7476);
and U8205 (N_8205,N_7300,N_7407);
or U8206 (N_8206,N_7127,N_7108);
nor U8207 (N_8207,N_7134,N_7480);
nor U8208 (N_8208,N_7167,N_6816);
or U8209 (N_8209,N_6948,N_7382);
or U8210 (N_8210,N_6995,N_7001);
nor U8211 (N_8211,N_7348,N_7154);
nor U8212 (N_8212,N_6782,N_6913);
xnor U8213 (N_8213,N_7265,N_6828);
and U8214 (N_8214,N_7484,N_7476);
and U8215 (N_8215,N_7343,N_7068);
or U8216 (N_8216,N_7250,N_7296);
or U8217 (N_8217,N_7481,N_7043);
and U8218 (N_8218,N_6885,N_6937);
nor U8219 (N_8219,N_7013,N_7327);
xor U8220 (N_8220,N_6964,N_7364);
or U8221 (N_8221,N_7324,N_6995);
xnor U8222 (N_8222,N_7185,N_6924);
or U8223 (N_8223,N_6963,N_7077);
xor U8224 (N_8224,N_7415,N_7202);
or U8225 (N_8225,N_7487,N_6857);
and U8226 (N_8226,N_7171,N_7427);
or U8227 (N_8227,N_7130,N_7184);
and U8228 (N_8228,N_6995,N_7352);
or U8229 (N_8229,N_6831,N_6909);
or U8230 (N_8230,N_7478,N_7153);
and U8231 (N_8231,N_7489,N_7371);
nand U8232 (N_8232,N_7122,N_6795);
and U8233 (N_8233,N_7202,N_6921);
nand U8234 (N_8234,N_6795,N_6859);
or U8235 (N_8235,N_7476,N_6915);
xnor U8236 (N_8236,N_7373,N_7145);
xnor U8237 (N_8237,N_7106,N_7463);
nor U8238 (N_8238,N_7164,N_7239);
xor U8239 (N_8239,N_6887,N_7335);
and U8240 (N_8240,N_7223,N_7221);
xnor U8241 (N_8241,N_6760,N_7321);
xnor U8242 (N_8242,N_7298,N_6863);
or U8243 (N_8243,N_7310,N_6859);
nor U8244 (N_8244,N_7125,N_7325);
xnor U8245 (N_8245,N_6882,N_6804);
nand U8246 (N_8246,N_7126,N_6772);
or U8247 (N_8247,N_7195,N_7005);
nor U8248 (N_8248,N_6778,N_6852);
nor U8249 (N_8249,N_7098,N_7005);
nand U8250 (N_8250,N_8075,N_7701);
nand U8251 (N_8251,N_8232,N_7987);
or U8252 (N_8252,N_8097,N_7738);
nand U8253 (N_8253,N_7525,N_8082);
nand U8254 (N_8254,N_8059,N_8036);
nor U8255 (N_8255,N_7782,N_8246);
and U8256 (N_8256,N_8127,N_8115);
and U8257 (N_8257,N_7893,N_7875);
and U8258 (N_8258,N_7789,N_8028);
xor U8259 (N_8259,N_7592,N_7857);
nor U8260 (N_8260,N_7953,N_8234);
and U8261 (N_8261,N_7980,N_8033);
and U8262 (N_8262,N_7575,N_7684);
nor U8263 (N_8263,N_7785,N_7669);
and U8264 (N_8264,N_7905,N_8219);
nor U8265 (N_8265,N_8190,N_7708);
xnor U8266 (N_8266,N_8169,N_7871);
and U8267 (N_8267,N_7947,N_7619);
xnor U8268 (N_8268,N_8151,N_8236);
xor U8269 (N_8269,N_7555,N_7858);
and U8270 (N_8270,N_8118,N_7724);
nor U8271 (N_8271,N_8024,N_7897);
and U8272 (N_8272,N_8021,N_7595);
xor U8273 (N_8273,N_8098,N_7794);
or U8274 (N_8274,N_7502,N_7921);
nand U8275 (N_8275,N_7859,N_8144);
nand U8276 (N_8276,N_7550,N_7851);
or U8277 (N_8277,N_8068,N_7647);
and U8278 (N_8278,N_7621,N_8215);
and U8279 (N_8279,N_7951,N_7566);
xnor U8280 (N_8280,N_7615,N_7558);
and U8281 (N_8281,N_8218,N_8119);
and U8282 (N_8282,N_8030,N_7725);
or U8283 (N_8283,N_7998,N_8062);
and U8284 (N_8284,N_7802,N_7690);
xor U8285 (N_8285,N_7672,N_7836);
nand U8286 (N_8286,N_7777,N_8240);
or U8287 (N_8287,N_7767,N_8243);
xnor U8288 (N_8288,N_7878,N_7553);
nand U8289 (N_8289,N_7907,N_7677);
xnor U8290 (N_8290,N_7913,N_7806);
nor U8291 (N_8291,N_7624,N_7706);
nand U8292 (N_8292,N_7795,N_7854);
and U8293 (N_8293,N_7713,N_8235);
and U8294 (N_8294,N_7920,N_7877);
xnor U8295 (N_8295,N_8106,N_8136);
nor U8296 (N_8296,N_8084,N_7526);
nand U8297 (N_8297,N_7779,N_7509);
and U8298 (N_8298,N_8195,N_7564);
nand U8299 (N_8299,N_8147,N_7975);
nor U8300 (N_8300,N_7818,N_8081);
or U8301 (N_8301,N_8100,N_8242);
xnor U8302 (N_8302,N_7830,N_8227);
and U8303 (N_8303,N_8079,N_8006);
nand U8304 (N_8304,N_8065,N_7801);
and U8305 (N_8305,N_7579,N_7589);
nor U8306 (N_8306,N_7629,N_7780);
nand U8307 (N_8307,N_8025,N_8086);
xnor U8308 (N_8308,N_8198,N_8070);
xnor U8309 (N_8309,N_8249,N_7847);
or U8310 (N_8310,N_7899,N_7600);
nor U8311 (N_8311,N_7510,N_7511);
nor U8312 (N_8312,N_8206,N_8095);
nor U8313 (N_8313,N_7872,N_7903);
xor U8314 (N_8314,N_8183,N_8090);
nand U8315 (N_8315,N_7852,N_8055);
and U8316 (N_8316,N_7954,N_8103);
nand U8317 (N_8317,N_7741,N_7915);
and U8318 (N_8318,N_8133,N_7770);
nor U8319 (N_8319,N_8108,N_8110);
or U8320 (N_8320,N_7786,N_7973);
nor U8321 (N_8321,N_7939,N_8132);
and U8322 (N_8322,N_7582,N_7693);
xor U8323 (N_8323,N_7517,N_8117);
and U8324 (N_8324,N_7839,N_7529);
nand U8325 (N_8325,N_8238,N_8157);
xnor U8326 (N_8326,N_7565,N_8176);
nor U8327 (N_8327,N_8137,N_7856);
xnor U8328 (N_8328,N_7761,N_7750);
nand U8329 (N_8329,N_7923,N_7606);
nor U8330 (N_8330,N_7810,N_7547);
nand U8331 (N_8331,N_8091,N_7758);
xnor U8332 (N_8332,N_8208,N_7784);
nor U8333 (N_8333,N_7844,N_7640);
or U8334 (N_8334,N_8221,N_7747);
xor U8335 (N_8335,N_7949,N_7571);
and U8336 (N_8336,N_8085,N_7709);
xnor U8337 (N_8337,N_7500,N_8120);
or U8338 (N_8338,N_7632,N_8032);
nor U8339 (N_8339,N_7674,N_8201);
or U8340 (N_8340,N_7503,N_7874);
or U8341 (N_8341,N_8166,N_7756);
and U8342 (N_8342,N_7804,N_7710);
and U8343 (N_8343,N_7599,N_7530);
and U8344 (N_8344,N_7653,N_8066);
nor U8345 (N_8345,N_8116,N_8224);
and U8346 (N_8346,N_7745,N_7753);
xnor U8347 (N_8347,N_8057,N_7838);
xor U8348 (N_8348,N_8016,N_7612);
xor U8349 (N_8349,N_7772,N_7976);
xnor U8350 (N_8350,N_7751,N_7528);
or U8351 (N_8351,N_7937,N_7828);
xor U8352 (N_8352,N_8229,N_7654);
xnor U8353 (N_8353,N_7989,N_7749);
xnor U8354 (N_8354,N_7603,N_8138);
xnor U8355 (N_8355,N_7679,N_7814);
or U8356 (N_8356,N_7630,N_7918);
xnor U8357 (N_8357,N_8245,N_8019);
nand U8358 (N_8358,N_7744,N_7666);
or U8359 (N_8359,N_7723,N_8143);
and U8360 (N_8360,N_8087,N_7800);
and U8361 (N_8361,N_8193,N_7574);
nand U8362 (N_8362,N_8153,N_7812);
or U8363 (N_8363,N_7898,N_8010);
nand U8364 (N_8364,N_7917,N_7730);
and U8365 (N_8365,N_7896,N_7676);
nor U8366 (N_8366,N_7675,N_8156);
and U8367 (N_8367,N_7831,N_8172);
and U8368 (N_8368,N_8017,N_7885);
nand U8369 (N_8369,N_7737,N_7729);
xor U8370 (N_8370,N_7644,N_7864);
or U8371 (N_8371,N_8128,N_7527);
xnor U8372 (N_8372,N_8222,N_8060);
and U8373 (N_8373,N_7734,N_7646);
and U8374 (N_8374,N_7966,N_7576);
nor U8375 (N_8375,N_7557,N_7657);
and U8376 (N_8376,N_7775,N_7799);
and U8377 (N_8377,N_8163,N_7754);
nand U8378 (N_8378,N_7561,N_7938);
nand U8379 (N_8379,N_7720,N_7868);
nor U8380 (N_8380,N_8158,N_8211);
xnor U8381 (N_8381,N_8225,N_8113);
and U8382 (N_8382,N_7820,N_7585);
or U8383 (N_8383,N_7835,N_7608);
or U8384 (N_8384,N_7583,N_7964);
or U8385 (N_8385,N_7546,N_7959);
and U8386 (N_8386,N_7886,N_8063);
nand U8387 (N_8387,N_8135,N_7922);
xor U8388 (N_8388,N_7656,N_7781);
and U8389 (N_8389,N_7876,N_8165);
nor U8390 (N_8390,N_7648,N_8023);
xnor U8391 (N_8391,N_7670,N_7650);
nor U8392 (N_8392,N_7787,N_7687);
nor U8393 (N_8393,N_8054,N_7727);
nor U8394 (N_8394,N_7521,N_8223);
and U8395 (N_8395,N_7620,N_7933);
and U8396 (N_8396,N_7819,N_8022);
nand U8397 (N_8397,N_8121,N_8209);
nand U8398 (N_8398,N_8125,N_7540);
or U8399 (N_8399,N_7531,N_7642);
xor U8400 (N_8400,N_7807,N_8168);
nand U8401 (N_8401,N_7793,N_7904);
nand U8402 (N_8402,N_7604,N_8126);
and U8403 (N_8403,N_7759,N_8226);
xnor U8404 (N_8404,N_8067,N_7614);
nand U8405 (N_8405,N_8058,N_7637);
nor U8406 (N_8406,N_8196,N_7680);
xnor U8407 (N_8407,N_7635,N_8044);
or U8408 (N_8408,N_7909,N_7813);
nand U8409 (N_8409,N_7548,N_8192);
or U8410 (N_8410,N_7972,N_7570);
or U8411 (N_8411,N_8146,N_8189);
nand U8412 (N_8412,N_7587,N_8233);
nor U8413 (N_8413,N_7934,N_7631);
nand U8414 (N_8414,N_7884,N_7829);
or U8415 (N_8415,N_7969,N_7978);
or U8416 (N_8416,N_7613,N_7742);
nor U8417 (N_8417,N_7662,N_7541);
or U8418 (N_8418,N_8074,N_7661);
nand U8419 (N_8419,N_7816,N_7971);
nand U8420 (N_8420,N_8186,N_7522);
xor U8421 (N_8421,N_7977,N_8034);
nand U8422 (N_8422,N_7707,N_8145);
or U8423 (N_8423,N_8161,N_7883);
xor U8424 (N_8424,N_7771,N_7873);
nand U8425 (N_8425,N_7736,N_7982);
nor U8426 (N_8426,N_7992,N_7968);
nor U8427 (N_8427,N_8105,N_7728);
xnor U8428 (N_8428,N_8013,N_7542);
xnor U8429 (N_8429,N_7688,N_8173);
or U8430 (N_8430,N_8080,N_7649);
or U8431 (N_8431,N_7912,N_7983);
and U8432 (N_8432,N_7501,N_7593);
and U8433 (N_8433,N_7590,N_8042);
and U8434 (N_8434,N_7869,N_7792);
nor U8435 (N_8435,N_8099,N_7961);
or U8436 (N_8436,N_8204,N_7967);
or U8437 (N_8437,N_8139,N_7948);
nor U8438 (N_8438,N_7714,N_7523);
nor U8439 (N_8439,N_7718,N_7958);
and U8440 (N_8440,N_7910,N_7834);
and U8441 (N_8441,N_7837,N_8009);
nand U8442 (N_8442,N_7651,N_8007);
nand U8443 (N_8443,N_8191,N_7733);
nand U8444 (N_8444,N_7732,N_7683);
and U8445 (N_8445,N_8152,N_7860);
nor U8446 (N_8446,N_7658,N_7768);
nand U8447 (N_8447,N_8029,N_7735);
or U8448 (N_8448,N_7508,N_7705);
nand U8449 (N_8449,N_7914,N_7848);
nor U8450 (N_8450,N_7625,N_7569);
and U8451 (N_8451,N_7927,N_7908);
and U8452 (N_8452,N_7668,N_7962);
or U8453 (N_8453,N_7673,N_7929);
nand U8454 (N_8454,N_8045,N_7699);
or U8455 (N_8455,N_8247,N_7586);
xor U8456 (N_8456,N_7892,N_7752);
nor U8457 (N_8457,N_7634,N_7638);
nand U8458 (N_8458,N_7941,N_7827);
or U8459 (N_8459,N_7974,N_7950);
and U8460 (N_8460,N_7660,N_8051);
nor U8461 (N_8461,N_7757,N_8202);
and U8462 (N_8462,N_8162,N_8076);
xor U8463 (N_8463,N_8216,N_7945);
xor U8464 (N_8464,N_7610,N_7686);
and U8465 (N_8465,N_7861,N_8140);
nand U8466 (N_8466,N_8041,N_8171);
nor U8467 (N_8467,N_7957,N_7639);
nand U8468 (N_8468,N_7946,N_7891);
and U8469 (N_8469,N_7715,N_7822);
and U8470 (N_8470,N_7930,N_8154);
and U8471 (N_8471,N_7623,N_8170);
nor U8472 (N_8472,N_7731,N_8150);
and U8473 (N_8473,N_7943,N_8038);
nand U8474 (N_8474,N_7766,N_8122);
xor U8475 (N_8475,N_7549,N_8071);
nand U8476 (N_8476,N_7740,N_8129);
xnor U8477 (N_8477,N_8187,N_7598);
or U8478 (N_8478,N_7524,N_7539);
nand U8479 (N_8479,N_8130,N_8160);
and U8480 (N_8480,N_8047,N_7817);
or U8481 (N_8481,N_8089,N_7901);
xor U8482 (N_8482,N_7988,N_7769);
or U8483 (N_8483,N_7536,N_8230);
nand U8484 (N_8484,N_7984,N_7833);
nand U8485 (N_8485,N_7931,N_7534);
xnor U8486 (N_8486,N_7597,N_7717);
nor U8487 (N_8487,N_8210,N_7652);
nor U8488 (N_8488,N_7694,N_8014);
nand U8489 (N_8489,N_8248,N_7504);
nand U8490 (N_8490,N_7726,N_8181);
nor U8491 (N_8491,N_8175,N_8214);
xnor U8492 (N_8492,N_8123,N_7963);
xor U8493 (N_8493,N_7562,N_8037);
and U8494 (N_8494,N_7849,N_7618);
and U8495 (N_8495,N_7895,N_8102);
and U8496 (N_8496,N_8109,N_7790);
xnor U8497 (N_8497,N_7952,N_7843);
and U8498 (N_8498,N_7823,N_7664);
or U8499 (N_8499,N_7986,N_8124);
nor U8500 (N_8500,N_7870,N_7889);
nor U8501 (N_8501,N_8179,N_8184);
nor U8502 (N_8502,N_8053,N_7783);
or U8503 (N_8503,N_7743,N_7712);
and U8504 (N_8504,N_8008,N_7513);
nor U8505 (N_8505,N_8069,N_8178);
or U8506 (N_8506,N_7826,N_8011);
xor U8507 (N_8507,N_7805,N_7846);
or U8508 (N_8508,N_8049,N_8003);
nand U8509 (N_8509,N_8180,N_7655);
nand U8510 (N_8510,N_7554,N_7567);
nor U8511 (N_8511,N_8056,N_7935);
xor U8512 (N_8512,N_8148,N_7695);
or U8513 (N_8513,N_8188,N_7760);
or U8514 (N_8514,N_7532,N_7545);
and U8515 (N_8515,N_7956,N_8185);
nand U8516 (N_8516,N_8043,N_7719);
nor U8517 (N_8517,N_7588,N_7515);
or U8518 (N_8518,N_7867,N_7681);
or U8519 (N_8519,N_8134,N_7552);
xor U8520 (N_8520,N_7773,N_7824);
or U8521 (N_8521,N_8159,N_8104);
and U8522 (N_8522,N_7538,N_7512);
or U8523 (N_8523,N_8094,N_7568);
xnor U8524 (N_8524,N_8182,N_7890);
nor U8525 (N_8525,N_7739,N_7888);
or U8526 (N_8526,N_7797,N_8239);
and U8527 (N_8527,N_7911,N_8174);
nor U8528 (N_8528,N_7641,N_7533);
or U8529 (N_8529,N_7560,N_7840);
and U8530 (N_8530,N_8207,N_8228);
xor U8531 (N_8531,N_7559,N_7796);
or U8532 (N_8532,N_8237,N_7936);
xnor U8533 (N_8533,N_7605,N_8112);
xnor U8534 (N_8534,N_7821,N_7841);
and U8535 (N_8535,N_7622,N_7979);
xnor U8536 (N_8536,N_8142,N_7996);
or U8537 (N_8537,N_8027,N_7584);
nor U8538 (N_8538,N_7716,N_7685);
nand U8539 (N_8539,N_7985,N_7572);
xnor U8540 (N_8540,N_8167,N_7645);
or U8541 (N_8541,N_7765,N_7762);
nor U8542 (N_8542,N_7711,N_8052);
or U8543 (N_8543,N_7906,N_7879);
xnor U8544 (N_8544,N_7696,N_8073);
and U8545 (N_8545,N_8131,N_7940);
or U8546 (N_8546,N_7722,N_7591);
and U8547 (N_8547,N_7698,N_7932);
nor U8548 (N_8548,N_7863,N_8203);
and U8549 (N_8549,N_8220,N_7809);
xor U8550 (N_8550,N_8088,N_8061);
xor U8551 (N_8551,N_7520,N_8205);
xor U8552 (N_8552,N_7850,N_7689);
or U8553 (N_8553,N_8026,N_7700);
or U8554 (N_8554,N_7556,N_8194);
and U8555 (N_8555,N_8018,N_7551);
and U8556 (N_8556,N_7580,N_7815);
or U8557 (N_8557,N_7633,N_8149);
and U8558 (N_8558,N_8231,N_7791);
or U8559 (N_8559,N_8004,N_7507);
nand U8560 (N_8560,N_7506,N_7755);
and U8561 (N_8561,N_8217,N_7990);
xor U8562 (N_8562,N_7894,N_8093);
xor U8563 (N_8563,N_7981,N_7900);
nor U8564 (N_8564,N_7702,N_7960);
or U8565 (N_8565,N_8199,N_7519);
xnor U8566 (N_8566,N_7577,N_7926);
nand U8567 (N_8567,N_8107,N_8241);
or U8568 (N_8568,N_7671,N_7609);
xor U8569 (N_8569,N_7682,N_8111);
nor U8570 (N_8570,N_7616,N_7667);
xnor U8571 (N_8571,N_7774,N_7881);
nand U8572 (N_8572,N_8164,N_7803);
nand U8573 (N_8573,N_8035,N_7665);
and U8574 (N_8574,N_8040,N_7928);
xor U8575 (N_8575,N_7997,N_7970);
nor U8576 (N_8576,N_7607,N_7994);
or U8577 (N_8577,N_7721,N_8002);
nand U8578 (N_8578,N_7535,N_7505);
or U8579 (N_8579,N_7643,N_7788);
and U8580 (N_8580,N_7594,N_7543);
nand U8581 (N_8581,N_7866,N_7581);
nand U8582 (N_8582,N_7865,N_8092);
xnor U8583 (N_8583,N_7544,N_7627);
xnor U8584 (N_8584,N_7611,N_7617);
nand U8585 (N_8585,N_7811,N_8077);
and U8586 (N_8586,N_7902,N_7748);
xnor U8587 (N_8587,N_7602,N_7746);
or U8588 (N_8588,N_8213,N_7955);
nand U8589 (N_8589,N_8096,N_8050);
or U8590 (N_8590,N_7999,N_7991);
xnor U8591 (N_8591,N_7916,N_7887);
xnor U8592 (N_8592,N_7516,N_7995);
xor U8593 (N_8593,N_7563,N_7626);
nand U8594 (N_8594,N_7704,N_7596);
nor U8595 (N_8595,N_8048,N_8031);
nor U8596 (N_8596,N_7763,N_8244);
nor U8597 (N_8597,N_8012,N_7697);
nand U8598 (N_8598,N_7944,N_7993);
and U8599 (N_8599,N_8064,N_7601);
or U8600 (N_8600,N_8005,N_8114);
nor U8601 (N_8601,N_7842,N_8200);
nand U8602 (N_8602,N_7845,N_8155);
or U8603 (N_8603,N_7518,N_7663);
or U8604 (N_8604,N_7798,N_7691);
xnor U8605 (N_8605,N_7808,N_7925);
and U8606 (N_8606,N_8001,N_7924);
nand U8607 (N_8607,N_8141,N_7778);
nand U8608 (N_8608,N_7514,N_8083);
and U8609 (N_8609,N_8072,N_7764);
nand U8610 (N_8610,N_7628,N_7537);
nor U8611 (N_8611,N_7659,N_7855);
nor U8612 (N_8612,N_8039,N_7703);
nor U8613 (N_8613,N_8177,N_8015);
or U8614 (N_8614,N_8212,N_7880);
nor U8615 (N_8615,N_7573,N_7919);
or U8616 (N_8616,N_7832,N_8000);
nand U8617 (N_8617,N_7578,N_7942);
xnor U8618 (N_8618,N_8101,N_8046);
nand U8619 (N_8619,N_7825,N_7636);
nor U8620 (N_8620,N_7965,N_7776);
nand U8621 (N_8621,N_8197,N_7678);
nand U8622 (N_8622,N_7692,N_7853);
nand U8623 (N_8623,N_7882,N_7862);
or U8624 (N_8624,N_8078,N_8020);
and U8625 (N_8625,N_7823,N_7668);
nor U8626 (N_8626,N_7938,N_7550);
nand U8627 (N_8627,N_7675,N_7597);
xor U8628 (N_8628,N_7962,N_7552);
nor U8629 (N_8629,N_8169,N_7863);
xor U8630 (N_8630,N_8239,N_7959);
nor U8631 (N_8631,N_7519,N_7639);
xor U8632 (N_8632,N_8212,N_7803);
or U8633 (N_8633,N_7904,N_7525);
nor U8634 (N_8634,N_7600,N_8027);
nor U8635 (N_8635,N_7706,N_8182);
xnor U8636 (N_8636,N_8044,N_7852);
and U8637 (N_8637,N_8110,N_7958);
nor U8638 (N_8638,N_7595,N_7871);
and U8639 (N_8639,N_7512,N_7581);
and U8640 (N_8640,N_8067,N_7689);
xor U8641 (N_8641,N_8060,N_7718);
and U8642 (N_8642,N_7782,N_8189);
nand U8643 (N_8643,N_7999,N_7972);
and U8644 (N_8644,N_7645,N_7541);
nor U8645 (N_8645,N_7746,N_7852);
or U8646 (N_8646,N_7985,N_7688);
or U8647 (N_8647,N_7809,N_7614);
and U8648 (N_8648,N_8048,N_7876);
and U8649 (N_8649,N_7770,N_7827);
and U8650 (N_8650,N_7675,N_8138);
nand U8651 (N_8651,N_7839,N_8215);
xnor U8652 (N_8652,N_7939,N_7864);
nor U8653 (N_8653,N_7867,N_7860);
and U8654 (N_8654,N_7863,N_7771);
nor U8655 (N_8655,N_7534,N_7741);
nor U8656 (N_8656,N_8046,N_8024);
or U8657 (N_8657,N_7655,N_7771);
nor U8658 (N_8658,N_7881,N_7605);
nand U8659 (N_8659,N_7727,N_7857);
and U8660 (N_8660,N_7979,N_7976);
xor U8661 (N_8661,N_7616,N_8007);
nand U8662 (N_8662,N_7722,N_8134);
and U8663 (N_8663,N_8082,N_7828);
xor U8664 (N_8664,N_7600,N_7957);
nor U8665 (N_8665,N_7596,N_8040);
xor U8666 (N_8666,N_7763,N_8065);
nand U8667 (N_8667,N_7517,N_8170);
nor U8668 (N_8668,N_7923,N_8092);
nor U8669 (N_8669,N_7985,N_7648);
nand U8670 (N_8670,N_7567,N_7525);
nand U8671 (N_8671,N_7594,N_8015);
xnor U8672 (N_8672,N_7916,N_8188);
nor U8673 (N_8673,N_7619,N_7513);
nor U8674 (N_8674,N_7928,N_7672);
xnor U8675 (N_8675,N_7500,N_7953);
or U8676 (N_8676,N_8095,N_8023);
and U8677 (N_8677,N_7635,N_7651);
nand U8678 (N_8678,N_7603,N_7855);
nor U8679 (N_8679,N_8076,N_8059);
and U8680 (N_8680,N_7929,N_7549);
nand U8681 (N_8681,N_8035,N_7635);
and U8682 (N_8682,N_7670,N_7790);
and U8683 (N_8683,N_8032,N_7809);
or U8684 (N_8684,N_7802,N_7812);
nand U8685 (N_8685,N_7861,N_8036);
xor U8686 (N_8686,N_8167,N_7872);
and U8687 (N_8687,N_8118,N_8066);
nand U8688 (N_8688,N_8182,N_8027);
and U8689 (N_8689,N_7918,N_7792);
or U8690 (N_8690,N_7705,N_7833);
nand U8691 (N_8691,N_7737,N_8169);
xnor U8692 (N_8692,N_8048,N_7959);
xnor U8693 (N_8693,N_7543,N_8132);
xor U8694 (N_8694,N_8125,N_7825);
xnor U8695 (N_8695,N_8223,N_8211);
nand U8696 (N_8696,N_8079,N_7675);
and U8697 (N_8697,N_7647,N_7657);
nor U8698 (N_8698,N_7912,N_7772);
xnor U8699 (N_8699,N_7930,N_8152);
xnor U8700 (N_8700,N_7641,N_7885);
nor U8701 (N_8701,N_8074,N_7924);
nor U8702 (N_8702,N_7756,N_7779);
or U8703 (N_8703,N_8245,N_7643);
nor U8704 (N_8704,N_7836,N_8182);
nand U8705 (N_8705,N_7514,N_8186);
and U8706 (N_8706,N_7756,N_8215);
xnor U8707 (N_8707,N_7741,N_7887);
nand U8708 (N_8708,N_8231,N_8040);
or U8709 (N_8709,N_7746,N_7764);
xnor U8710 (N_8710,N_7510,N_7520);
or U8711 (N_8711,N_8096,N_7730);
xnor U8712 (N_8712,N_7748,N_7904);
and U8713 (N_8713,N_8121,N_7885);
nor U8714 (N_8714,N_8047,N_8065);
nor U8715 (N_8715,N_8036,N_7662);
nor U8716 (N_8716,N_7932,N_7542);
and U8717 (N_8717,N_7590,N_8022);
and U8718 (N_8718,N_7963,N_7536);
or U8719 (N_8719,N_7551,N_7732);
nor U8720 (N_8720,N_8091,N_7930);
nand U8721 (N_8721,N_7698,N_8067);
nor U8722 (N_8722,N_7976,N_7813);
nand U8723 (N_8723,N_7969,N_7913);
nand U8724 (N_8724,N_7953,N_7802);
xor U8725 (N_8725,N_7924,N_7736);
nor U8726 (N_8726,N_7832,N_7586);
nand U8727 (N_8727,N_7831,N_8208);
nand U8728 (N_8728,N_7706,N_7891);
or U8729 (N_8729,N_7794,N_8043);
xor U8730 (N_8730,N_8231,N_7770);
nand U8731 (N_8731,N_7925,N_8044);
nand U8732 (N_8732,N_7610,N_8111);
nor U8733 (N_8733,N_8086,N_7771);
or U8734 (N_8734,N_8198,N_7575);
nor U8735 (N_8735,N_7725,N_8228);
xor U8736 (N_8736,N_7680,N_7772);
xor U8737 (N_8737,N_8059,N_7942);
and U8738 (N_8738,N_8121,N_8190);
xnor U8739 (N_8739,N_7547,N_7692);
xor U8740 (N_8740,N_8211,N_7968);
or U8741 (N_8741,N_7948,N_7650);
nand U8742 (N_8742,N_7866,N_7697);
xor U8743 (N_8743,N_7873,N_7762);
and U8744 (N_8744,N_7727,N_7785);
xor U8745 (N_8745,N_7518,N_7857);
or U8746 (N_8746,N_8146,N_7698);
xor U8747 (N_8747,N_8198,N_8136);
nand U8748 (N_8748,N_8118,N_8009);
xnor U8749 (N_8749,N_8013,N_7513);
or U8750 (N_8750,N_8192,N_8058);
xor U8751 (N_8751,N_7547,N_8121);
nor U8752 (N_8752,N_7723,N_8136);
and U8753 (N_8753,N_8005,N_7734);
xor U8754 (N_8754,N_7798,N_7779);
nand U8755 (N_8755,N_8232,N_7914);
nor U8756 (N_8756,N_7681,N_8082);
nand U8757 (N_8757,N_8089,N_8179);
nand U8758 (N_8758,N_7582,N_7545);
and U8759 (N_8759,N_8236,N_7952);
and U8760 (N_8760,N_8029,N_7678);
and U8761 (N_8761,N_8084,N_7676);
nor U8762 (N_8762,N_7728,N_8187);
nand U8763 (N_8763,N_7794,N_7795);
nand U8764 (N_8764,N_7795,N_7579);
xor U8765 (N_8765,N_8216,N_7561);
nand U8766 (N_8766,N_8002,N_7555);
nor U8767 (N_8767,N_8230,N_7579);
or U8768 (N_8768,N_7935,N_7741);
nor U8769 (N_8769,N_8161,N_7737);
or U8770 (N_8770,N_8154,N_7640);
nor U8771 (N_8771,N_7566,N_7511);
nor U8772 (N_8772,N_7809,N_7707);
xor U8773 (N_8773,N_7637,N_8240);
xor U8774 (N_8774,N_7872,N_7512);
or U8775 (N_8775,N_7798,N_7828);
nor U8776 (N_8776,N_7742,N_7906);
xor U8777 (N_8777,N_7807,N_8107);
xnor U8778 (N_8778,N_7515,N_7854);
xnor U8779 (N_8779,N_7790,N_7608);
and U8780 (N_8780,N_8084,N_8116);
nor U8781 (N_8781,N_8111,N_7753);
and U8782 (N_8782,N_7925,N_7727);
or U8783 (N_8783,N_7899,N_7921);
xor U8784 (N_8784,N_7727,N_7511);
or U8785 (N_8785,N_8121,N_7946);
xnor U8786 (N_8786,N_7518,N_7938);
nor U8787 (N_8787,N_7999,N_7599);
nor U8788 (N_8788,N_8126,N_8137);
nand U8789 (N_8789,N_7663,N_7843);
or U8790 (N_8790,N_7981,N_8168);
nor U8791 (N_8791,N_7767,N_7743);
and U8792 (N_8792,N_7902,N_8227);
nand U8793 (N_8793,N_7576,N_7579);
xnor U8794 (N_8794,N_7803,N_7731);
or U8795 (N_8795,N_8071,N_7967);
or U8796 (N_8796,N_7945,N_8144);
nand U8797 (N_8797,N_7589,N_7658);
nand U8798 (N_8798,N_7537,N_7633);
or U8799 (N_8799,N_8181,N_7582);
nand U8800 (N_8800,N_7794,N_7917);
nand U8801 (N_8801,N_7581,N_7823);
or U8802 (N_8802,N_8176,N_7837);
nor U8803 (N_8803,N_7882,N_7675);
xor U8804 (N_8804,N_8111,N_7847);
xor U8805 (N_8805,N_7500,N_7886);
xnor U8806 (N_8806,N_7994,N_8088);
nor U8807 (N_8807,N_8074,N_7846);
nand U8808 (N_8808,N_7756,N_7760);
nor U8809 (N_8809,N_8070,N_7872);
or U8810 (N_8810,N_7787,N_7878);
nand U8811 (N_8811,N_8175,N_7716);
xnor U8812 (N_8812,N_7509,N_8065);
nand U8813 (N_8813,N_7961,N_8218);
or U8814 (N_8814,N_7824,N_8162);
nand U8815 (N_8815,N_8090,N_7501);
nor U8816 (N_8816,N_7932,N_8139);
nor U8817 (N_8817,N_7745,N_8087);
nor U8818 (N_8818,N_8130,N_7568);
nand U8819 (N_8819,N_8191,N_7692);
nor U8820 (N_8820,N_7599,N_7644);
nand U8821 (N_8821,N_7719,N_7881);
xnor U8822 (N_8822,N_8166,N_8241);
and U8823 (N_8823,N_7977,N_7670);
xor U8824 (N_8824,N_8068,N_7685);
or U8825 (N_8825,N_7724,N_7555);
xnor U8826 (N_8826,N_7745,N_7936);
nand U8827 (N_8827,N_7753,N_7621);
nor U8828 (N_8828,N_7978,N_7571);
nor U8829 (N_8829,N_7924,N_7947);
nor U8830 (N_8830,N_8049,N_7578);
or U8831 (N_8831,N_7734,N_8111);
xor U8832 (N_8832,N_8170,N_8085);
or U8833 (N_8833,N_7850,N_7755);
or U8834 (N_8834,N_8102,N_8238);
or U8835 (N_8835,N_8075,N_7802);
nand U8836 (N_8836,N_7510,N_8040);
nor U8837 (N_8837,N_7611,N_8120);
or U8838 (N_8838,N_7666,N_7686);
nand U8839 (N_8839,N_8089,N_8147);
and U8840 (N_8840,N_7650,N_7667);
or U8841 (N_8841,N_7792,N_8117);
or U8842 (N_8842,N_7579,N_7930);
xor U8843 (N_8843,N_8211,N_8081);
nand U8844 (N_8844,N_8015,N_7523);
nand U8845 (N_8845,N_7868,N_7786);
or U8846 (N_8846,N_7980,N_8231);
and U8847 (N_8847,N_7634,N_8130);
and U8848 (N_8848,N_7918,N_7773);
nand U8849 (N_8849,N_7941,N_7927);
xor U8850 (N_8850,N_8226,N_8124);
nand U8851 (N_8851,N_7790,N_7965);
xor U8852 (N_8852,N_8134,N_8062);
or U8853 (N_8853,N_8093,N_8066);
or U8854 (N_8854,N_7958,N_7780);
or U8855 (N_8855,N_7875,N_7951);
nand U8856 (N_8856,N_8025,N_7649);
nand U8857 (N_8857,N_8246,N_7879);
and U8858 (N_8858,N_8244,N_7789);
and U8859 (N_8859,N_8200,N_7665);
and U8860 (N_8860,N_7521,N_8107);
nor U8861 (N_8861,N_7514,N_8114);
xor U8862 (N_8862,N_7618,N_7968);
and U8863 (N_8863,N_8065,N_8142);
and U8864 (N_8864,N_7552,N_8139);
xnor U8865 (N_8865,N_8053,N_7639);
xor U8866 (N_8866,N_7540,N_7547);
or U8867 (N_8867,N_7732,N_8184);
nand U8868 (N_8868,N_8045,N_7725);
nor U8869 (N_8869,N_7863,N_7798);
nor U8870 (N_8870,N_7519,N_8040);
nor U8871 (N_8871,N_7536,N_8090);
nor U8872 (N_8872,N_7816,N_7593);
nand U8873 (N_8873,N_7639,N_7890);
nor U8874 (N_8874,N_7606,N_7694);
or U8875 (N_8875,N_7592,N_8171);
xor U8876 (N_8876,N_7820,N_7580);
nand U8877 (N_8877,N_8000,N_8089);
or U8878 (N_8878,N_8019,N_7986);
and U8879 (N_8879,N_7579,N_7671);
nor U8880 (N_8880,N_7872,N_7675);
nand U8881 (N_8881,N_7597,N_7637);
xor U8882 (N_8882,N_7741,N_8171);
or U8883 (N_8883,N_7938,N_8150);
nor U8884 (N_8884,N_7515,N_7682);
nand U8885 (N_8885,N_7804,N_7785);
nand U8886 (N_8886,N_7628,N_7503);
xor U8887 (N_8887,N_7955,N_7523);
and U8888 (N_8888,N_7943,N_7933);
xor U8889 (N_8889,N_8045,N_7949);
xnor U8890 (N_8890,N_8099,N_7897);
and U8891 (N_8891,N_7768,N_7509);
nor U8892 (N_8892,N_8073,N_7964);
nor U8893 (N_8893,N_7975,N_7694);
nand U8894 (N_8894,N_8243,N_7790);
or U8895 (N_8895,N_7620,N_7799);
and U8896 (N_8896,N_7899,N_7768);
nor U8897 (N_8897,N_7597,N_7590);
xor U8898 (N_8898,N_7664,N_8015);
and U8899 (N_8899,N_7726,N_7639);
or U8900 (N_8900,N_7858,N_7982);
or U8901 (N_8901,N_8005,N_8115);
xnor U8902 (N_8902,N_7933,N_8150);
and U8903 (N_8903,N_7941,N_7543);
xor U8904 (N_8904,N_8064,N_8120);
nand U8905 (N_8905,N_8193,N_8195);
or U8906 (N_8906,N_7964,N_8084);
nand U8907 (N_8907,N_7882,N_7948);
or U8908 (N_8908,N_8191,N_7759);
nor U8909 (N_8909,N_7599,N_8057);
and U8910 (N_8910,N_8201,N_8063);
nor U8911 (N_8911,N_7672,N_8117);
nand U8912 (N_8912,N_7858,N_8022);
or U8913 (N_8913,N_8116,N_8131);
and U8914 (N_8914,N_7626,N_7846);
nor U8915 (N_8915,N_7552,N_7932);
nand U8916 (N_8916,N_7517,N_8113);
xor U8917 (N_8917,N_7918,N_7821);
nor U8918 (N_8918,N_7902,N_8133);
nor U8919 (N_8919,N_8106,N_7820);
xnor U8920 (N_8920,N_7919,N_7784);
nand U8921 (N_8921,N_8237,N_7530);
and U8922 (N_8922,N_7548,N_7794);
or U8923 (N_8923,N_7722,N_7916);
xnor U8924 (N_8924,N_8212,N_7776);
or U8925 (N_8925,N_8092,N_7606);
nor U8926 (N_8926,N_7970,N_7739);
or U8927 (N_8927,N_8008,N_7893);
and U8928 (N_8928,N_7787,N_7954);
nor U8929 (N_8929,N_8120,N_7543);
and U8930 (N_8930,N_7890,N_7566);
and U8931 (N_8931,N_7799,N_8083);
or U8932 (N_8932,N_7677,N_8186);
xnor U8933 (N_8933,N_7794,N_8031);
nand U8934 (N_8934,N_7926,N_8208);
and U8935 (N_8935,N_8144,N_7925);
xnor U8936 (N_8936,N_7836,N_7899);
nor U8937 (N_8937,N_7505,N_7956);
and U8938 (N_8938,N_8008,N_8128);
or U8939 (N_8939,N_7966,N_8067);
nand U8940 (N_8940,N_8236,N_7718);
or U8941 (N_8941,N_8233,N_7982);
nor U8942 (N_8942,N_7668,N_7660);
or U8943 (N_8943,N_8072,N_7613);
nand U8944 (N_8944,N_7593,N_7652);
nor U8945 (N_8945,N_7592,N_7900);
or U8946 (N_8946,N_7795,N_7759);
or U8947 (N_8947,N_7778,N_7788);
nor U8948 (N_8948,N_8171,N_8077);
nand U8949 (N_8949,N_8044,N_7730);
xnor U8950 (N_8950,N_8217,N_8224);
and U8951 (N_8951,N_8220,N_7784);
nor U8952 (N_8952,N_8226,N_7688);
nand U8953 (N_8953,N_7824,N_7913);
nor U8954 (N_8954,N_8126,N_7674);
or U8955 (N_8955,N_7587,N_7560);
xor U8956 (N_8956,N_7897,N_7975);
or U8957 (N_8957,N_7627,N_8239);
xor U8958 (N_8958,N_7823,N_8121);
or U8959 (N_8959,N_8047,N_7678);
nand U8960 (N_8960,N_7669,N_8002);
xor U8961 (N_8961,N_7807,N_7524);
nor U8962 (N_8962,N_7513,N_7501);
xnor U8963 (N_8963,N_8105,N_8232);
or U8964 (N_8964,N_7551,N_7836);
and U8965 (N_8965,N_8064,N_7746);
xor U8966 (N_8966,N_7797,N_8154);
and U8967 (N_8967,N_7917,N_7716);
nand U8968 (N_8968,N_7927,N_8127);
xor U8969 (N_8969,N_7553,N_7818);
or U8970 (N_8970,N_7509,N_7950);
and U8971 (N_8971,N_7694,N_8032);
and U8972 (N_8972,N_8081,N_8207);
nand U8973 (N_8973,N_7796,N_8055);
and U8974 (N_8974,N_8033,N_7630);
and U8975 (N_8975,N_8063,N_8034);
and U8976 (N_8976,N_7523,N_8074);
nor U8977 (N_8977,N_8155,N_8026);
and U8978 (N_8978,N_8021,N_7633);
and U8979 (N_8979,N_7747,N_7631);
or U8980 (N_8980,N_7934,N_7588);
xnor U8981 (N_8981,N_7997,N_7740);
xnor U8982 (N_8982,N_8170,N_7842);
and U8983 (N_8983,N_8121,N_7855);
or U8984 (N_8984,N_8193,N_7631);
xor U8985 (N_8985,N_7887,N_7522);
or U8986 (N_8986,N_7504,N_7624);
nor U8987 (N_8987,N_7622,N_8024);
nor U8988 (N_8988,N_8085,N_8058);
nor U8989 (N_8989,N_7803,N_7734);
or U8990 (N_8990,N_7779,N_7508);
and U8991 (N_8991,N_7979,N_7664);
nor U8992 (N_8992,N_7654,N_7997);
and U8993 (N_8993,N_8212,N_8192);
nor U8994 (N_8994,N_7921,N_8070);
xnor U8995 (N_8995,N_7907,N_7861);
xor U8996 (N_8996,N_7967,N_7647);
or U8997 (N_8997,N_7577,N_7550);
and U8998 (N_8998,N_7953,N_7898);
nor U8999 (N_8999,N_8178,N_7739);
nand U9000 (N_9000,N_8809,N_8368);
nand U9001 (N_9001,N_8489,N_8847);
or U9002 (N_9002,N_8909,N_8933);
and U9003 (N_9003,N_8363,N_8356);
nand U9004 (N_9004,N_8409,N_8423);
nor U9005 (N_9005,N_8448,N_8360);
and U9006 (N_9006,N_8281,N_8561);
and U9007 (N_9007,N_8577,N_8879);
nor U9008 (N_9008,N_8829,N_8650);
nor U9009 (N_9009,N_8928,N_8585);
and U9010 (N_9010,N_8957,N_8992);
xor U9011 (N_9011,N_8627,N_8660);
or U9012 (N_9012,N_8674,N_8497);
nand U9013 (N_9013,N_8366,N_8835);
xor U9014 (N_9014,N_8420,N_8995);
nor U9015 (N_9015,N_8542,N_8944);
nand U9016 (N_9016,N_8527,N_8776);
and U9017 (N_9017,N_8442,N_8440);
nor U9018 (N_9018,N_8738,N_8739);
nand U9019 (N_9019,N_8945,N_8595);
xnor U9020 (N_9020,N_8669,N_8330);
and U9021 (N_9021,N_8289,N_8837);
and U9022 (N_9022,N_8437,N_8586);
or U9023 (N_9023,N_8814,N_8544);
xnor U9024 (N_9024,N_8500,N_8400);
and U9025 (N_9025,N_8433,N_8887);
and U9026 (N_9026,N_8372,N_8275);
and U9027 (N_9027,N_8850,N_8834);
or U9028 (N_9028,N_8301,N_8720);
nor U9029 (N_9029,N_8274,N_8846);
xor U9030 (N_9030,N_8937,N_8284);
nand U9031 (N_9031,N_8564,N_8656);
nand U9032 (N_9032,N_8996,N_8287);
nand U9033 (N_9033,N_8278,N_8751);
and U9034 (N_9034,N_8839,N_8815);
or U9035 (N_9035,N_8292,N_8371);
and U9036 (N_9036,N_8302,N_8419);
nor U9037 (N_9037,N_8294,N_8477);
nor U9038 (N_9038,N_8759,N_8454);
and U9039 (N_9039,N_8304,N_8820);
xor U9040 (N_9040,N_8606,N_8646);
nand U9041 (N_9041,N_8798,N_8900);
nor U9042 (N_9042,N_8745,N_8699);
xor U9043 (N_9043,N_8563,N_8482);
nand U9044 (N_9044,N_8971,N_8723);
xor U9045 (N_9045,N_8282,N_8469);
and U9046 (N_9046,N_8668,N_8279);
and U9047 (N_9047,N_8936,N_8300);
nand U9048 (N_9048,N_8303,N_8889);
and U9049 (N_9049,N_8805,N_8509);
xnor U9050 (N_9050,N_8393,N_8633);
xor U9051 (N_9051,N_8915,N_8793);
nand U9052 (N_9052,N_8886,N_8685);
nand U9053 (N_9053,N_8891,N_8298);
nor U9054 (N_9054,N_8731,N_8744);
nand U9055 (N_9055,N_8781,N_8286);
nor U9056 (N_9056,N_8600,N_8620);
nand U9057 (N_9057,N_8441,N_8692);
nor U9058 (N_9058,N_8569,N_8686);
xnor U9059 (N_9059,N_8852,N_8696);
and U9060 (N_9060,N_8940,N_8431);
nor U9061 (N_9061,N_8460,N_8474);
nand U9062 (N_9062,N_8794,N_8567);
nand U9063 (N_9063,N_8402,N_8775);
and U9064 (N_9064,N_8664,N_8713);
or U9065 (N_9065,N_8276,N_8521);
nand U9066 (N_9066,N_8753,N_8718);
xnor U9067 (N_9067,N_8908,N_8432);
nor U9068 (N_9068,N_8967,N_8350);
or U9069 (N_9069,N_8817,N_8895);
nand U9070 (N_9070,N_8415,N_8740);
xnor U9071 (N_9071,N_8533,N_8640);
and U9072 (N_9072,N_8486,N_8898);
nor U9073 (N_9073,N_8314,N_8765);
xor U9074 (N_9074,N_8516,N_8288);
and U9075 (N_9075,N_8355,N_8362);
xnor U9076 (N_9076,N_8743,N_8969);
nor U9077 (N_9077,N_8758,N_8466);
or U9078 (N_9078,N_8271,N_8614);
nand U9079 (N_9079,N_8580,N_8926);
xnor U9080 (N_9080,N_8783,N_8306);
or U9081 (N_9081,N_8608,N_8536);
and U9082 (N_9082,N_8724,N_8851);
nand U9083 (N_9083,N_8800,N_8755);
nand U9084 (N_9084,N_8760,N_8719);
xnor U9085 (N_9085,N_8418,N_8872);
or U9086 (N_9086,N_8747,N_8546);
xnor U9087 (N_9087,N_8920,N_8435);
nor U9088 (N_9088,N_8436,N_8568);
xnor U9089 (N_9089,N_8796,N_8924);
nand U9090 (N_9090,N_8260,N_8559);
xnor U9091 (N_9091,N_8667,N_8311);
or U9092 (N_9092,N_8407,N_8451);
and U9093 (N_9093,N_8315,N_8736);
xor U9094 (N_9094,N_8259,N_8804);
and U9095 (N_9095,N_8923,N_8532);
nor U9096 (N_9096,N_8985,N_8327);
xnor U9097 (N_9097,N_8921,N_8914);
nand U9098 (N_9098,N_8677,N_8273);
xor U9099 (N_9099,N_8896,N_8251);
xnor U9100 (N_9100,N_8772,N_8617);
nor U9101 (N_9101,N_8445,N_8866);
nor U9102 (N_9102,N_8263,N_8390);
or U9103 (N_9103,N_8771,N_8575);
or U9104 (N_9104,N_8974,N_8426);
nor U9105 (N_9105,N_8679,N_8512);
nor U9106 (N_9106,N_8396,N_8658);
xor U9107 (N_9107,N_8405,N_8748);
nor U9108 (N_9108,N_8966,N_8652);
or U9109 (N_9109,N_8865,N_8553);
and U9110 (N_9110,N_8810,N_8874);
nor U9111 (N_9111,N_8507,N_8663);
or U9112 (N_9112,N_8792,N_8603);
or U9113 (N_9113,N_8361,N_8571);
nor U9114 (N_9114,N_8429,N_8391);
or U9115 (N_9115,N_8700,N_8636);
or U9116 (N_9116,N_8806,N_8853);
nand U9117 (N_9117,N_8791,N_8681);
and U9118 (N_9118,N_8828,N_8358);
nor U9119 (N_9119,N_8994,N_8905);
nor U9120 (N_9120,N_8819,N_8680);
or U9121 (N_9121,N_8399,N_8897);
and U9122 (N_9122,N_8989,N_8671);
and U9123 (N_9123,N_8919,N_8344);
xor U9124 (N_9124,N_8757,N_8875);
nor U9125 (N_9125,N_8635,N_8709);
nor U9126 (N_9126,N_8557,N_8517);
and U9127 (N_9127,N_8539,N_8843);
and U9128 (N_9128,N_8737,N_8638);
and U9129 (N_9129,N_8458,N_8666);
xnor U9130 (N_9130,N_8822,N_8935);
and U9131 (N_9131,N_8922,N_8811);
xor U9132 (N_9132,N_8647,N_8428);
nand U9133 (N_9133,N_8854,N_8716);
xnor U9134 (N_9134,N_8708,N_8845);
nor U9135 (N_9135,N_8902,N_8778);
nor U9136 (N_9136,N_8756,N_8763);
and U9137 (N_9137,N_8918,N_8857);
nand U9138 (N_9138,N_8998,N_8714);
nor U9139 (N_9139,N_8882,N_8654);
and U9140 (N_9140,N_8554,N_8392);
xnor U9141 (N_9141,N_8593,N_8977);
xor U9142 (N_9142,N_8750,N_8883);
xnor U9143 (N_9143,N_8425,N_8616);
or U9144 (N_9144,N_8495,N_8450);
nor U9145 (N_9145,N_8774,N_8842);
nor U9146 (N_9146,N_8907,N_8528);
nor U9147 (N_9147,N_8421,N_8297);
xor U9148 (N_9148,N_8324,N_8754);
nor U9149 (N_9149,N_8816,N_8256);
and U9150 (N_9150,N_8523,N_8988);
xor U9151 (N_9151,N_8767,N_8867);
xnor U9152 (N_9152,N_8332,N_8480);
nor U9153 (N_9153,N_8272,N_8351);
nor U9154 (N_9154,N_8964,N_8732);
or U9155 (N_9155,N_8683,N_8978);
and U9156 (N_9156,N_8370,N_8548);
and U9157 (N_9157,N_8628,N_8773);
nor U9158 (N_9158,N_8325,N_8932);
and U9159 (N_9159,N_8508,N_8901);
xor U9160 (N_9160,N_8269,N_8946);
nand U9161 (N_9161,N_8629,N_8515);
and U9162 (N_9162,N_8841,N_8795);
nand U9163 (N_9163,N_8594,N_8782);
nand U9164 (N_9164,N_8849,N_8406);
nor U9165 (N_9165,N_8343,N_8576);
xnor U9166 (N_9166,N_8444,N_8510);
and U9167 (N_9167,N_8910,N_8927);
xor U9168 (N_9168,N_8524,N_8547);
and U9169 (N_9169,N_8698,N_8844);
nor U9170 (N_9170,N_8439,N_8305);
nand U9171 (N_9171,N_8549,N_8651);
nor U9172 (N_9172,N_8825,N_8999);
and U9173 (N_9173,N_8769,N_8255);
xor U9174 (N_9174,N_8701,N_8912);
nand U9175 (N_9175,N_8856,N_8352);
xnor U9176 (N_9176,N_8592,N_8943);
and U9177 (N_9177,N_8871,N_8560);
or U9178 (N_9178,N_8704,N_8438);
nand U9179 (N_9179,N_8764,N_8965);
xor U9180 (N_9180,N_8505,N_8947);
nand U9181 (N_9181,N_8803,N_8729);
xnor U9182 (N_9182,N_8383,N_8317);
and U9183 (N_9183,N_8499,N_8550);
or U9184 (N_9184,N_8726,N_8631);
nand U9185 (N_9185,N_8833,N_8987);
and U9186 (N_9186,N_8641,N_8869);
nand U9187 (N_9187,N_8596,N_8687);
nand U9188 (N_9188,N_8963,N_8789);
and U9189 (N_9189,N_8644,N_8838);
nor U9190 (N_9190,N_8457,N_8648);
or U9191 (N_9191,N_8788,N_8503);
xor U9192 (N_9192,N_8813,N_8376);
or U9193 (N_9193,N_8335,N_8802);
xnor U9194 (N_9194,N_8894,N_8582);
xor U9195 (N_9195,N_8630,N_8490);
xnor U9196 (N_9196,N_8341,N_8684);
or U9197 (N_9197,N_8348,N_8868);
xor U9198 (N_9198,N_8878,N_8715);
nor U9199 (N_9199,N_8401,N_8388);
or U9200 (N_9200,N_8917,N_8414);
or U9201 (N_9201,N_8456,N_8742);
nor U9202 (N_9202,N_8379,N_8607);
xnor U9203 (N_9203,N_8855,N_8545);
nand U9204 (N_9204,N_8291,N_8446);
and U9205 (N_9205,N_8583,N_8252);
xnor U9206 (N_9206,N_8707,N_8541);
or U9207 (N_9207,N_8934,N_8321);
nor U9208 (N_9208,N_8254,N_8359);
nand U9209 (N_9209,N_8787,N_8519);
xor U9210 (N_9210,N_8377,N_8903);
nand U9211 (N_9211,N_8290,N_8562);
nor U9212 (N_9212,N_8973,N_8821);
xor U9213 (N_9213,N_8530,N_8982);
nand U9214 (N_9214,N_8380,N_8955);
nand U9215 (N_9215,N_8981,N_8369);
nor U9216 (N_9216,N_8960,N_8502);
nor U9217 (N_9217,N_8318,N_8676);
or U9218 (N_9218,N_8329,N_8312);
nor U9219 (N_9219,N_8899,N_8340);
nor U9220 (N_9220,N_8342,N_8398);
and U9221 (N_9221,N_8345,N_8411);
xor U9222 (N_9222,N_8862,N_8552);
xor U9223 (N_9223,N_8752,N_8602);
nand U9224 (N_9224,N_8331,N_8830);
and U9225 (N_9225,N_8534,N_8639);
or U9226 (N_9226,N_8522,N_8797);
nor U9227 (N_9227,N_8991,N_8483);
or U9228 (N_9228,N_8334,N_8501);
xnor U9229 (N_9229,N_8597,N_8690);
xnor U9230 (N_9230,N_8277,N_8378);
xnor U9231 (N_9231,N_8395,N_8790);
nand U9232 (N_9232,N_8962,N_8703);
and U9233 (N_9233,N_8827,N_8632);
nand U9234 (N_9234,N_8566,N_8610);
nor U9235 (N_9235,N_8320,N_8386);
xnor U9236 (N_9236,N_8518,N_8970);
or U9237 (N_9237,N_8467,N_8367);
nor U9238 (N_9238,N_8471,N_8925);
or U9239 (N_9239,N_8473,N_8643);
nor U9240 (N_9240,N_8824,N_8389);
or U9241 (N_9241,N_8434,N_8478);
nor U9242 (N_9242,N_8893,N_8702);
or U9243 (N_9243,N_8826,N_8950);
and U9244 (N_9244,N_8884,N_8514);
nor U9245 (N_9245,N_8462,N_8622);
nand U9246 (N_9246,N_8976,N_8717);
nor U9247 (N_9247,N_8659,N_8464);
nand U9248 (N_9248,N_8859,N_8374);
or U9249 (N_9249,N_8730,N_8961);
and U9250 (N_9250,N_8556,N_8836);
or U9251 (N_9251,N_8721,N_8615);
xnor U9252 (N_9252,N_8385,N_8734);
nand U9253 (N_9253,N_8506,N_8476);
nor U9254 (N_9254,N_8397,N_8525);
and U9255 (N_9255,N_8258,N_8354);
nand U9256 (N_9256,N_8877,N_8682);
xnor U9257 (N_9257,N_8712,N_8689);
or U9258 (N_9258,N_8888,N_8766);
or U9259 (N_9259,N_8916,N_8537);
and U9260 (N_9260,N_8293,N_8799);
nand U9261 (N_9261,N_8860,N_8558);
xnor U9262 (N_9262,N_8468,N_8410);
xnor U9263 (N_9263,N_8319,N_8349);
xor U9264 (N_9264,N_8316,N_8941);
or U9265 (N_9265,N_8858,N_8487);
nor U9266 (N_9266,N_8812,N_8417);
and U9267 (N_9267,N_8601,N_8831);
xnor U9268 (N_9268,N_8430,N_8453);
or U9269 (N_9269,N_8770,N_8590);
nand U9270 (N_9270,N_8496,N_8939);
nand U9271 (N_9271,N_8675,N_8688);
or U9272 (N_9272,N_8694,N_8840);
xor U9273 (N_9273,N_8322,N_8997);
or U9274 (N_9274,N_8535,N_8818);
xnor U9275 (N_9275,N_8746,N_8339);
xnor U9276 (N_9276,N_8705,N_8672);
and U9277 (N_9277,N_8848,N_8634);
xor U9278 (N_9278,N_8779,N_8832);
nand U9279 (N_9279,N_8513,N_8262);
nor U9280 (N_9280,N_8484,N_8491);
xor U9281 (N_9281,N_8619,N_8954);
and U9282 (N_9282,N_8265,N_8538);
nand U9283 (N_9283,N_8481,N_8861);
nor U9284 (N_9284,N_8381,N_8949);
nor U9285 (N_9285,N_8777,N_8983);
xnor U9286 (N_9286,N_8543,N_8531);
or U9287 (N_9287,N_8975,N_8266);
or U9288 (N_9288,N_8413,N_8412);
nand U9289 (N_9289,N_8447,N_8336);
or U9290 (N_9290,N_8365,N_8749);
and U9291 (N_9291,N_8261,N_8885);
nor U9292 (N_9292,N_8710,N_8599);
and U9293 (N_9293,N_8403,N_8588);
nand U9294 (N_9294,N_8364,N_8959);
and U9295 (N_9295,N_8299,N_8357);
nand U9296 (N_9296,N_8823,N_8493);
nand U9297 (N_9297,N_8711,N_8253);
nand U9298 (N_9298,N_8626,N_8931);
nor U9299 (N_9299,N_8725,N_8881);
or U9300 (N_9300,N_8979,N_8876);
and U9301 (N_9301,N_8761,N_8578);
or U9302 (N_9302,N_8511,N_8670);
and U9303 (N_9303,N_8873,N_8906);
and U9304 (N_9304,N_8598,N_8980);
nand U9305 (N_9305,N_8526,N_8661);
xnor U9306 (N_9306,N_8416,N_8972);
nor U9307 (N_9307,N_8488,N_8613);
xor U9308 (N_9308,N_8455,N_8498);
and U9309 (N_9309,N_8581,N_8695);
xnor U9310 (N_9310,N_8863,N_8727);
xnor U9311 (N_9311,N_8573,N_8485);
and U9312 (N_9312,N_8465,N_8786);
xnor U9313 (N_9313,N_8986,N_8952);
or U9314 (N_9314,N_8930,N_8459);
nand U9315 (N_9315,N_8449,N_8382);
nor U9316 (N_9316,N_8384,N_8611);
xor U9317 (N_9317,N_8993,N_8741);
nor U9318 (N_9318,N_8285,N_8653);
and U9319 (N_9319,N_8733,N_8310);
and U9320 (N_9320,N_8475,N_8948);
nor U9321 (N_9321,N_8589,N_8250);
nor U9322 (N_9322,N_8373,N_8904);
xor U9323 (N_9323,N_8264,N_8308);
nor U9324 (N_9324,N_8333,N_8870);
and U9325 (N_9325,N_8693,N_8990);
nand U9326 (N_9326,N_8492,N_8624);
and U9327 (N_9327,N_8645,N_8612);
nor U9328 (N_9328,N_8323,N_8911);
and U9329 (N_9329,N_8280,N_8604);
xor U9330 (N_9330,N_8938,N_8579);
nand U9331 (N_9331,N_8609,N_8587);
xnor U9332 (N_9332,N_8623,N_8649);
xnor U9333 (N_9333,N_8662,N_8504);
and U9334 (N_9334,N_8665,N_8313);
nand U9335 (N_9335,N_8953,N_8422);
nand U9336 (N_9336,N_8642,N_8618);
or U9337 (N_9337,N_8942,N_8387);
nor U9338 (N_9338,N_8892,N_8762);
nor U9339 (N_9339,N_8295,N_8309);
nand U9340 (N_9340,N_8807,N_8637);
nor U9341 (N_9341,N_8565,N_8574);
or U9342 (N_9342,N_8968,N_8808);
nor U9343 (N_9343,N_8570,N_8890);
and U9344 (N_9344,N_8801,N_8984);
xor U9345 (N_9345,N_8768,N_8472);
xnor U9346 (N_9346,N_8338,N_8929);
xnor U9347 (N_9347,N_8551,N_8555);
nor U9348 (N_9348,N_8328,N_8268);
nor U9349 (N_9349,N_8691,N_8267);
nand U9350 (N_9350,N_8470,N_8706);
xor U9351 (N_9351,N_8283,N_8591);
nor U9352 (N_9352,N_8520,N_8326);
and U9353 (N_9353,N_8443,N_8864);
xnor U9354 (N_9354,N_8394,N_8452);
nand U9355 (N_9355,N_8337,N_8958);
and U9356 (N_9356,N_8404,N_8408);
nor U9357 (N_9357,N_8346,N_8347);
nor U9358 (N_9358,N_8621,N_8913);
nor U9359 (N_9359,N_8307,N_8427);
xor U9360 (N_9360,N_8572,N_8673);
nand U9361 (N_9361,N_8780,N_8951);
or U9362 (N_9362,N_8657,N_8605);
nor U9363 (N_9363,N_8880,N_8270);
nand U9364 (N_9364,N_8296,N_8424);
nor U9365 (N_9365,N_8540,N_8353);
or U9366 (N_9366,N_8529,N_8463);
nand U9367 (N_9367,N_8257,N_8697);
nand U9368 (N_9368,N_8461,N_8728);
nand U9369 (N_9369,N_8625,N_8494);
xnor U9370 (N_9370,N_8655,N_8956);
xnor U9371 (N_9371,N_8735,N_8784);
nor U9372 (N_9372,N_8785,N_8375);
nand U9373 (N_9373,N_8584,N_8678);
or U9374 (N_9374,N_8722,N_8479);
and U9375 (N_9375,N_8708,N_8474);
nor U9376 (N_9376,N_8510,N_8392);
nand U9377 (N_9377,N_8534,N_8861);
or U9378 (N_9378,N_8848,N_8780);
xor U9379 (N_9379,N_8309,N_8808);
xnor U9380 (N_9380,N_8330,N_8963);
nor U9381 (N_9381,N_8662,N_8385);
nand U9382 (N_9382,N_8372,N_8799);
or U9383 (N_9383,N_8417,N_8333);
or U9384 (N_9384,N_8341,N_8782);
or U9385 (N_9385,N_8589,N_8769);
nand U9386 (N_9386,N_8428,N_8429);
nor U9387 (N_9387,N_8986,N_8390);
or U9388 (N_9388,N_8581,N_8403);
and U9389 (N_9389,N_8702,N_8716);
nor U9390 (N_9390,N_8543,N_8583);
and U9391 (N_9391,N_8597,N_8899);
and U9392 (N_9392,N_8961,N_8645);
and U9393 (N_9393,N_8441,N_8724);
xnor U9394 (N_9394,N_8346,N_8619);
xnor U9395 (N_9395,N_8829,N_8812);
and U9396 (N_9396,N_8272,N_8346);
nor U9397 (N_9397,N_8497,N_8694);
or U9398 (N_9398,N_8847,N_8270);
nor U9399 (N_9399,N_8550,N_8570);
and U9400 (N_9400,N_8423,N_8573);
nor U9401 (N_9401,N_8675,N_8972);
nand U9402 (N_9402,N_8386,N_8993);
xor U9403 (N_9403,N_8759,N_8865);
or U9404 (N_9404,N_8317,N_8977);
nand U9405 (N_9405,N_8471,N_8614);
xnor U9406 (N_9406,N_8305,N_8384);
and U9407 (N_9407,N_8562,N_8649);
xor U9408 (N_9408,N_8754,N_8347);
nand U9409 (N_9409,N_8257,N_8375);
nor U9410 (N_9410,N_8830,N_8665);
or U9411 (N_9411,N_8493,N_8880);
xnor U9412 (N_9412,N_8608,N_8272);
xnor U9413 (N_9413,N_8373,N_8493);
nand U9414 (N_9414,N_8623,N_8928);
nor U9415 (N_9415,N_8587,N_8519);
nor U9416 (N_9416,N_8951,N_8877);
or U9417 (N_9417,N_8992,N_8548);
xor U9418 (N_9418,N_8291,N_8753);
nor U9419 (N_9419,N_8779,N_8878);
or U9420 (N_9420,N_8933,N_8886);
nor U9421 (N_9421,N_8952,N_8922);
nor U9422 (N_9422,N_8659,N_8764);
nand U9423 (N_9423,N_8472,N_8493);
and U9424 (N_9424,N_8873,N_8855);
nand U9425 (N_9425,N_8983,N_8746);
nand U9426 (N_9426,N_8723,N_8481);
and U9427 (N_9427,N_8384,N_8841);
and U9428 (N_9428,N_8319,N_8820);
and U9429 (N_9429,N_8531,N_8629);
nand U9430 (N_9430,N_8254,N_8990);
and U9431 (N_9431,N_8576,N_8713);
and U9432 (N_9432,N_8985,N_8651);
nand U9433 (N_9433,N_8495,N_8856);
nand U9434 (N_9434,N_8835,N_8359);
xnor U9435 (N_9435,N_8614,N_8446);
or U9436 (N_9436,N_8667,N_8885);
and U9437 (N_9437,N_8750,N_8321);
and U9438 (N_9438,N_8625,N_8836);
or U9439 (N_9439,N_8797,N_8956);
and U9440 (N_9440,N_8695,N_8943);
and U9441 (N_9441,N_8469,N_8778);
nand U9442 (N_9442,N_8254,N_8888);
or U9443 (N_9443,N_8977,N_8929);
xnor U9444 (N_9444,N_8875,N_8648);
nor U9445 (N_9445,N_8659,N_8971);
nor U9446 (N_9446,N_8555,N_8774);
nor U9447 (N_9447,N_8331,N_8470);
nor U9448 (N_9448,N_8522,N_8446);
and U9449 (N_9449,N_8582,N_8494);
and U9450 (N_9450,N_8480,N_8797);
or U9451 (N_9451,N_8896,N_8526);
nor U9452 (N_9452,N_8963,N_8474);
or U9453 (N_9453,N_8742,N_8903);
or U9454 (N_9454,N_8798,N_8710);
xnor U9455 (N_9455,N_8352,N_8251);
and U9456 (N_9456,N_8888,N_8739);
and U9457 (N_9457,N_8907,N_8943);
or U9458 (N_9458,N_8747,N_8899);
nand U9459 (N_9459,N_8506,N_8437);
or U9460 (N_9460,N_8821,N_8376);
nand U9461 (N_9461,N_8854,N_8996);
nor U9462 (N_9462,N_8692,N_8644);
nor U9463 (N_9463,N_8524,N_8799);
xor U9464 (N_9464,N_8948,N_8451);
nand U9465 (N_9465,N_8821,N_8731);
xor U9466 (N_9466,N_8564,N_8607);
xor U9467 (N_9467,N_8733,N_8388);
nor U9468 (N_9468,N_8977,N_8982);
nand U9469 (N_9469,N_8377,N_8715);
or U9470 (N_9470,N_8551,N_8930);
xor U9471 (N_9471,N_8597,N_8506);
nand U9472 (N_9472,N_8624,N_8917);
xor U9473 (N_9473,N_8394,N_8789);
nand U9474 (N_9474,N_8480,N_8763);
nor U9475 (N_9475,N_8883,N_8259);
and U9476 (N_9476,N_8992,N_8848);
xnor U9477 (N_9477,N_8494,N_8452);
and U9478 (N_9478,N_8984,N_8653);
or U9479 (N_9479,N_8863,N_8352);
and U9480 (N_9480,N_8262,N_8700);
or U9481 (N_9481,N_8729,N_8977);
or U9482 (N_9482,N_8910,N_8622);
nor U9483 (N_9483,N_8975,N_8982);
or U9484 (N_9484,N_8400,N_8579);
nor U9485 (N_9485,N_8717,N_8485);
nand U9486 (N_9486,N_8318,N_8906);
nand U9487 (N_9487,N_8523,N_8319);
or U9488 (N_9488,N_8604,N_8450);
nand U9489 (N_9489,N_8389,N_8641);
and U9490 (N_9490,N_8590,N_8926);
and U9491 (N_9491,N_8360,N_8372);
nor U9492 (N_9492,N_8727,N_8558);
or U9493 (N_9493,N_8758,N_8599);
nand U9494 (N_9494,N_8665,N_8361);
xnor U9495 (N_9495,N_8932,N_8287);
nand U9496 (N_9496,N_8691,N_8900);
nand U9497 (N_9497,N_8463,N_8859);
xnor U9498 (N_9498,N_8647,N_8502);
nor U9499 (N_9499,N_8973,N_8915);
nor U9500 (N_9500,N_8432,N_8440);
nand U9501 (N_9501,N_8584,N_8727);
nand U9502 (N_9502,N_8339,N_8787);
or U9503 (N_9503,N_8874,N_8364);
xnor U9504 (N_9504,N_8789,N_8871);
nor U9505 (N_9505,N_8958,N_8477);
xnor U9506 (N_9506,N_8547,N_8755);
xnor U9507 (N_9507,N_8897,N_8888);
nand U9508 (N_9508,N_8591,N_8689);
nand U9509 (N_9509,N_8421,N_8381);
xor U9510 (N_9510,N_8392,N_8878);
and U9511 (N_9511,N_8545,N_8290);
or U9512 (N_9512,N_8400,N_8268);
or U9513 (N_9513,N_8792,N_8808);
nand U9514 (N_9514,N_8880,N_8422);
or U9515 (N_9515,N_8345,N_8427);
and U9516 (N_9516,N_8558,N_8765);
or U9517 (N_9517,N_8875,N_8657);
or U9518 (N_9518,N_8646,N_8644);
and U9519 (N_9519,N_8901,N_8291);
xnor U9520 (N_9520,N_8336,N_8340);
nand U9521 (N_9521,N_8483,N_8519);
xnor U9522 (N_9522,N_8303,N_8542);
nand U9523 (N_9523,N_8293,N_8457);
nor U9524 (N_9524,N_8415,N_8833);
and U9525 (N_9525,N_8970,N_8531);
or U9526 (N_9526,N_8702,N_8335);
and U9527 (N_9527,N_8705,N_8746);
xor U9528 (N_9528,N_8578,N_8770);
nand U9529 (N_9529,N_8462,N_8635);
or U9530 (N_9530,N_8573,N_8807);
xnor U9531 (N_9531,N_8296,N_8506);
xnor U9532 (N_9532,N_8397,N_8888);
and U9533 (N_9533,N_8332,N_8678);
nand U9534 (N_9534,N_8696,N_8941);
nand U9535 (N_9535,N_8361,N_8629);
or U9536 (N_9536,N_8620,N_8434);
xor U9537 (N_9537,N_8946,N_8288);
or U9538 (N_9538,N_8278,N_8433);
nand U9539 (N_9539,N_8494,N_8332);
and U9540 (N_9540,N_8620,N_8951);
nand U9541 (N_9541,N_8587,N_8949);
nand U9542 (N_9542,N_8642,N_8369);
nand U9543 (N_9543,N_8987,N_8345);
and U9544 (N_9544,N_8891,N_8771);
or U9545 (N_9545,N_8865,N_8455);
or U9546 (N_9546,N_8461,N_8560);
nor U9547 (N_9547,N_8273,N_8439);
or U9548 (N_9548,N_8635,N_8976);
nor U9549 (N_9549,N_8800,N_8841);
or U9550 (N_9550,N_8866,N_8734);
xor U9551 (N_9551,N_8919,N_8772);
or U9552 (N_9552,N_8587,N_8600);
nor U9553 (N_9553,N_8283,N_8484);
nand U9554 (N_9554,N_8911,N_8532);
or U9555 (N_9555,N_8636,N_8468);
and U9556 (N_9556,N_8292,N_8831);
nand U9557 (N_9557,N_8605,N_8830);
or U9558 (N_9558,N_8952,N_8426);
nor U9559 (N_9559,N_8955,N_8573);
nor U9560 (N_9560,N_8870,N_8565);
xor U9561 (N_9561,N_8384,N_8404);
or U9562 (N_9562,N_8440,N_8276);
nand U9563 (N_9563,N_8384,N_8511);
nor U9564 (N_9564,N_8985,N_8946);
or U9565 (N_9565,N_8688,N_8484);
and U9566 (N_9566,N_8763,N_8365);
and U9567 (N_9567,N_8581,N_8639);
nand U9568 (N_9568,N_8753,N_8749);
and U9569 (N_9569,N_8864,N_8398);
nand U9570 (N_9570,N_8844,N_8732);
nand U9571 (N_9571,N_8291,N_8768);
and U9572 (N_9572,N_8862,N_8759);
and U9573 (N_9573,N_8893,N_8272);
xor U9574 (N_9574,N_8480,N_8652);
xnor U9575 (N_9575,N_8454,N_8389);
nand U9576 (N_9576,N_8873,N_8468);
and U9577 (N_9577,N_8256,N_8324);
or U9578 (N_9578,N_8798,N_8353);
and U9579 (N_9579,N_8302,N_8730);
nor U9580 (N_9580,N_8973,N_8719);
nand U9581 (N_9581,N_8788,N_8500);
nand U9582 (N_9582,N_8924,N_8351);
nand U9583 (N_9583,N_8606,N_8857);
nor U9584 (N_9584,N_8312,N_8808);
nand U9585 (N_9585,N_8943,N_8701);
nand U9586 (N_9586,N_8559,N_8814);
nor U9587 (N_9587,N_8979,N_8259);
nor U9588 (N_9588,N_8459,N_8615);
nand U9589 (N_9589,N_8482,N_8411);
nand U9590 (N_9590,N_8816,N_8482);
nor U9591 (N_9591,N_8547,N_8922);
or U9592 (N_9592,N_8653,N_8670);
and U9593 (N_9593,N_8991,N_8657);
nand U9594 (N_9594,N_8502,N_8751);
xnor U9595 (N_9595,N_8876,N_8528);
and U9596 (N_9596,N_8651,N_8561);
and U9597 (N_9597,N_8948,N_8813);
or U9598 (N_9598,N_8685,N_8783);
xor U9599 (N_9599,N_8553,N_8693);
nand U9600 (N_9600,N_8870,N_8379);
nor U9601 (N_9601,N_8364,N_8415);
and U9602 (N_9602,N_8519,N_8380);
and U9603 (N_9603,N_8846,N_8823);
nand U9604 (N_9604,N_8654,N_8458);
or U9605 (N_9605,N_8343,N_8503);
xor U9606 (N_9606,N_8414,N_8993);
xor U9607 (N_9607,N_8777,N_8920);
nor U9608 (N_9608,N_8366,N_8915);
or U9609 (N_9609,N_8604,N_8568);
and U9610 (N_9610,N_8460,N_8885);
xor U9611 (N_9611,N_8470,N_8948);
nor U9612 (N_9612,N_8564,N_8776);
and U9613 (N_9613,N_8893,N_8681);
and U9614 (N_9614,N_8647,N_8741);
and U9615 (N_9615,N_8756,N_8789);
xnor U9616 (N_9616,N_8765,N_8550);
or U9617 (N_9617,N_8792,N_8578);
xor U9618 (N_9618,N_8522,N_8493);
nor U9619 (N_9619,N_8575,N_8665);
xor U9620 (N_9620,N_8822,N_8556);
nor U9621 (N_9621,N_8600,N_8714);
nand U9622 (N_9622,N_8617,N_8261);
xnor U9623 (N_9623,N_8618,N_8447);
nand U9624 (N_9624,N_8456,N_8452);
and U9625 (N_9625,N_8966,N_8295);
nand U9626 (N_9626,N_8449,N_8560);
nand U9627 (N_9627,N_8913,N_8354);
and U9628 (N_9628,N_8374,N_8366);
or U9629 (N_9629,N_8788,N_8767);
nand U9630 (N_9630,N_8793,N_8818);
or U9631 (N_9631,N_8995,N_8515);
xor U9632 (N_9632,N_8854,N_8380);
nor U9633 (N_9633,N_8651,N_8383);
xnor U9634 (N_9634,N_8561,N_8965);
xnor U9635 (N_9635,N_8683,N_8496);
or U9636 (N_9636,N_8680,N_8861);
nand U9637 (N_9637,N_8868,N_8959);
xor U9638 (N_9638,N_8731,N_8386);
nand U9639 (N_9639,N_8922,N_8264);
nor U9640 (N_9640,N_8519,N_8534);
or U9641 (N_9641,N_8621,N_8946);
nand U9642 (N_9642,N_8923,N_8483);
nand U9643 (N_9643,N_8401,N_8602);
nor U9644 (N_9644,N_8906,N_8620);
or U9645 (N_9645,N_8517,N_8328);
or U9646 (N_9646,N_8804,N_8294);
or U9647 (N_9647,N_8936,N_8897);
nor U9648 (N_9648,N_8597,N_8751);
nor U9649 (N_9649,N_8712,N_8769);
and U9650 (N_9650,N_8502,N_8999);
or U9651 (N_9651,N_8496,N_8848);
and U9652 (N_9652,N_8684,N_8305);
nor U9653 (N_9653,N_8833,N_8843);
nand U9654 (N_9654,N_8254,N_8569);
or U9655 (N_9655,N_8846,N_8475);
and U9656 (N_9656,N_8417,N_8955);
xor U9657 (N_9657,N_8932,N_8587);
nor U9658 (N_9658,N_8894,N_8985);
or U9659 (N_9659,N_8446,N_8596);
or U9660 (N_9660,N_8809,N_8535);
or U9661 (N_9661,N_8873,N_8874);
and U9662 (N_9662,N_8649,N_8736);
and U9663 (N_9663,N_8912,N_8810);
nor U9664 (N_9664,N_8539,N_8266);
and U9665 (N_9665,N_8255,N_8871);
xor U9666 (N_9666,N_8389,N_8812);
nand U9667 (N_9667,N_8259,N_8398);
or U9668 (N_9668,N_8740,N_8865);
nand U9669 (N_9669,N_8427,N_8486);
or U9670 (N_9670,N_8541,N_8672);
or U9671 (N_9671,N_8267,N_8407);
nor U9672 (N_9672,N_8511,N_8289);
nor U9673 (N_9673,N_8913,N_8916);
xor U9674 (N_9674,N_8939,N_8682);
nand U9675 (N_9675,N_8913,N_8526);
nand U9676 (N_9676,N_8413,N_8880);
nand U9677 (N_9677,N_8503,N_8623);
or U9678 (N_9678,N_8902,N_8514);
nor U9679 (N_9679,N_8724,N_8710);
nand U9680 (N_9680,N_8377,N_8599);
and U9681 (N_9681,N_8795,N_8760);
nor U9682 (N_9682,N_8729,N_8456);
nor U9683 (N_9683,N_8730,N_8867);
xor U9684 (N_9684,N_8882,N_8479);
nand U9685 (N_9685,N_8322,N_8422);
nor U9686 (N_9686,N_8583,N_8330);
nand U9687 (N_9687,N_8260,N_8775);
xor U9688 (N_9688,N_8542,N_8345);
nor U9689 (N_9689,N_8420,N_8534);
and U9690 (N_9690,N_8799,N_8272);
or U9691 (N_9691,N_8277,N_8939);
nor U9692 (N_9692,N_8519,N_8326);
nand U9693 (N_9693,N_8829,N_8531);
or U9694 (N_9694,N_8733,N_8655);
nor U9695 (N_9695,N_8673,N_8791);
and U9696 (N_9696,N_8697,N_8446);
or U9697 (N_9697,N_8588,N_8459);
nor U9698 (N_9698,N_8560,N_8339);
or U9699 (N_9699,N_8402,N_8642);
or U9700 (N_9700,N_8312,N_8701);
nand U9701 (N_9701,N_8851,N_8312);
nor U9702 (N_9702,N_8758,N_8632);
xnor U9703 (N_9703,N_8304,N_8574);
nor U9704 (N_9704,N_8642,N_8448);
and U9705 (N_9705,N_8739,N_8729);
xnor U9706 (N_9706,N_8936,N_8416);
nor U9707 (N_9707,N_8412,N_8835);
xor U9708 (N_9708,N_8547,N_8790);
and U9709 (N_9709,N_8395,N_8253);
xor U9710 (N_9710,N_8749,N_8973);
or U9711 (N_9711,N_8996,N_8556);
and U9712 (N_9712,N_8862,N_8669);
nand U9713 (N_9713,N_8381,N_8583);
nor U9714 (N_9714,N_8707,N_8551);
or U9715 (N_9715,N_8593,N_8789);
xor U9716 (N_9716,N_8879,N_8361);
nor U9717 (N_9717,N_8556,N_8656);
and U9718 (N_9718,N_8786,N_8589);
nand U9719 (N_9719,N_8715,N_8708);
and U9720 (N_9720,N_8545,N_8694);
nor U9721 (N_9721,N_8560,N_8572);
nor U9722 (N_9722,N_8674,N_8252);
and U9723 (N_9723,N_8260,N_8432);
nor U9724 (N_9724,N_8375,N_8639);
or U9725 (N_9725,N_8283,N_8574);
xor U9726 (N_9726,N_8440,N_8807);
nor U9727 (N_9727,N_8280,N_8464);
nand U9728 (N_9728,N_8786,N_8945);
xor U9729 (N_9729,N_8793,N_8805);
nand U9730 (N_9730,N_8350,N_8985);
or U9731 (N_9731,N_8461,N_8589);
nor U9732 (N_9732,N_8502,N_8393);
nand U9733 (N_9733,N_8364,N_8605);
and U9734 (N_9734,N_8613,N_8324);
xor U9735 (N_9735,N_8323,N_8561);
or U9736 (N_9736,N_8946,N_8954);
xor U9737 (N_9737,N_8350,N_8919);
nor U9738 (N_9738,N_8315,N_8262);
xnor U9739 (N_9739,N_8726,N_8502);
and U9740 (N_9740,N_8849,N_8473);
and U9741 (N_9741,N_8498,N_8699);
nand U9742 (N_9742,N_8603,N_8754);
and U9743 (N_9743,N_8478,N_8659);
nor U9744 (N_9744,N_8488,N_8674);
or U9745 (N_9745,N_8583,N_8644);
nor U9746 (N_9746,N_8844,N_8564);
or U9747 (N_9747,N_8550,N_8484);
nor U9748 (N_9748,N_8430,N_8669);
xor U9749 (N_9749,N_8843,N_8993);
nor U9750 (N_9750,N_9020,N_9592);
xor U9751 (N_9751,N_9030,N_9299);
or U9752 (N_9752,N_9194,N_9025);
nand U9753 (N_9753,N_9217,N_9174);
nor U9754 (N_9754,N_9094,N_9287);
xnor U9755 (N_9755,N_9080,N_9333);
nand U9756 (N_9756,N_9379,N_9008);
nand U9757 (N_9757,N_9411,N_9554);
nand U9758 (N_9758,N_9338,N_9571);
nand U9759 (N_9759,N_9405,N_9152);
and U9760 (N_9760,N_9532,N_9588);
and U9761 (N_9761,N_9419,N_9097);
nor U9762 (N_9762,N_9543,N_9691);
and U9763 (N_9763,N_9474,N_9160);
nor U9764 (N_9764,N_9440,N_9614);
or U9765 (N_9765,N_9507,N_9682);
or U9766 (N_9766,N_9205,N_9130);
nand U9767 (N_9767,N_9671,N_9118);
and U9768 (N_9768,N_9336,N_9653);
nand U9769 (N_9769,N_9086,N_9043);
nand U9770 (N_9770,N_9033,N_9500);
nor U9771 (N_9771,N_9222,N_9083);
or U9772 (N_9772,N_9428,N_9469);
xor U9773 (N_9773,N_9173,N_9503);
nand U9774 (N_9774,N_9393,N_9281);
xnor U9775 (N_9775,N_9465,N_9067);
nand U9776 (N_9776,N_9272,N_9321);
xor U9777 (N_9777,N_9505,N_9572);
xor U9778 (N_9778,N_9215,N_9334);
nor U9779 (N_9779,N_9446,N_9749);
nand U9780 (N_9780,N_9061,N_9093);
xor U9781 (N_9781,N_9212,N_9525);
nor U9782 (N_9782,N_9259,N_9734);
xor U9783 (N_9783,N_9323,N_9736);
or U9784 (N_9784,N_9109,N_9641);
xor U9785 (N_9785,N_9000,N_9552);
xor U9786 (N_9786,N_9280,N_9501);
nor U9787 (N_9787,N_9066,N_9024);
or U9788 (N_9788,N_9581,N_9385);
and U9789 (N_9789,N_9556,N_9089);
or U9790 (N_9790,N_9075,N_9575);
xnor U9791 (N_9791,N_9286,N_9538);
nand U9792 (N_9792,N_9463,N_9680);
xor U9793 (N_9793,N_9392,N_9598);
and U9794 (N_9794,N_9284,N_9052);
nor U9795 (N_9795,N_9417,N_9345);
nand U9796 (N_9796,N_9633,N_9491);
nand U9797 (N_9797,N_9748,N_9161);
and U9798 (N_9798,N_9712,N_9063);
nor U9799 (N_9799,N_9535,N_9143);
xor U9800 (N_9800,N_9518,N_9408);
nor U9801 (N_9801,N_9029,N_9149);
xnor U9802 (N_9802,N_9273,N_9478);
or U9803 (N_9803,N_9156,N_9056);
nor U9804 (N_9804,N_9241,N_9663);
xnor U9805 (N_9805,N_9206,N_9459);
xor U9806 (N_9806,N_9594,N_9434);
or U9807 (N_9807,N_9637,N_9542);
or U9808 (N_9808,N_9528,N_9632);
nand U9809 (N_9809,N_9693,N_9555);
xnor U9810 (N_9810,N_9486,N_9176);
nor U9811 (N_9811,N_9580,N_9074);
nor U9812 (N_9812,N_9037,N_9233);
nand U9813 (N_9813,N_9116,N_9510);
nand U9814 (N_9814,N_9125,N_9017);
nand U9815 (N_9815,N_9353,N_9366);
or U9816 (N_9816,N_9514,N_9047);
nor U9817 (N_9817,N_9689,N_9131);
nand U9818 (N_9818,N_9107,N_9108);
nand U9819 (N_9819,N_9639,N_9007);
xnor U9820 (N_9820,N_9375,N_9512);
nand U9821 (N_9821,N_9307,N_9560);
xor U9822 (N_9822,N_9140,N_9416);
or U9823 (N_9823,N_9620,N_9328);
and U9824 (N_9824,N_9231,N_9714);
and U9825 (N_9825,N_9187,N_9715);
and U9826 (N_9826,N_9103,N_9425);
nand U9827 (N_9827,N_9404,N_9488);
nand U9828 (N_9828,N_9487,N_9230);
nor U9829 (N_9829,N_9022,N_9256);
nor U9830 (N_9830,N_9679,N_9481);
nor U9831 (N_9831,N_9717,N_9648);
nand U9832 (N_9832,N_9036,N_9646);
xor U9833 (N_9833,N_9558,N_9211);
or U9834 (N_9834,N_9263,N_9498);
and U9835 (N_9835,N_9618,N_9248);
nand U9836 (N_9836,N_9119,N_9302);
nor U9837 (N_9837,N_9700,N_9027);
or U9838 (N_9838,N_9662,N_9190);
xor U9839 (N_9839,N_9124,N_9313);
nor U9840 (N_9840,N_9329,N_9562);
nand U9841 (N_9841,N_9553,N_9489);
nand U9842 (N_9842,N_9186,N_9331);
xnor U9843 (N_9843,N_9466,N_9378);
nor U9844 (N_9844,N_9049,N_9236);
xor U9845 (N_9845,N_9519,N_9189);
nand U9846 (N_9846,N_9681,N_9112);
xnor U9847 (N_9847,N_9249,N_9269);
xor U9848 (N_9848,N_9708,N_9227);
and U9849 (N_9849,N_9670,N_9062);
nand U9850 (N_9850,N_9358,N_9545);
or U9851 (N_9851,N_9615,N_9026);
and U9852 (N_9852,N_9628,N_9134);
xnor U9853 (N_9853,N_9669,N_9362);
nor U9854 (N_9854,N_9136,N_9595);
and U9855 (N_9855,N_9247,N_9617);
xnor U9856 (N_9856,N_9676,N_9101);
and U9857 (N_9857,N_9461,N_9407);
nand U9858 (N_9858,N_9665,N_9583);
and U9859 (N_9859,N_9630,N_9208);
nand U9860 (N_9860,N_9088,N_9198);
xnor U9861 (N_9861,N_9352,N_9442);
nor U9862 (N_9862,N_9373,N_9209);
nor U9863 (N_9863,N_9327,N_9707);
xnor U9864 (N_9864,N_9421,N_9695);
and U9865 (N_9865,N_9589,N_9141);
and U9866 (N_9866,N_9432,N_9306);
or U9867 (N_9867,N_9497,N_9480);
and U9868 (N_9868,N_9453,N_9292);
and U9869 (N_9869,N_9138,N_9744);
nand U9870 (N_9870,N_9418,N_9422);
or U9871 (N_9871,N_9485,N_9433);
and U9872 (N_9872,N_9339,N_9098);
nand U9873 (N_9873,N_9578,N_9710);
nand U9874 (N_9874,N_9087,N_9406);
nand U9875 (N_9875,N_9423,N_9511);
nand U9876 (N_9876,N_9585,N_9678);
and U9877 (N_9877,N_9424,N_9398);
and U9878 (N_9878,N_9252,N_9193);
nor U9879 (N_9879,N_9439,N_9240);
xnor U9880 (N_9880,N_9342,N_9283);
xnor U9881 (N_9881,N_9547,N_9105);
and U9882 (N_9882,N_9133,N_9364);
nor U9883 (N_9883,N_9636,N_9316);
nor U9884 (N_9884,N_9625,N_9733);
nor U9885 (N_9885,N_9300,N_9564);
nand U9886 (N_9886,N_9599,N_9294);
nor U9887 (N_9887,N_9743,N_9044);
xnor U9888 (N_9888,N_9386,N_9154);
nor U9889 (N_9889,N_9531,N_9719);
xnor U9890 (N_9890,N_9383,N_9644);
nor U9891 (N_9891,N_9735,N_9367);
or U9892 (N_9892,N_9242,N_9262);
or U9893 (N_9893,N_9293,N_9285);
nand U9894 (N_9894,N_9357,N_9218);
or U9895 (N_9895,N_9675,N_9310);
nand U9896 (N_9896,N_9182,N_9687);
or U9897 (N_9897,N_9229,N_9462);
or U9898 (N_9898,N_9110,N_9275);
nand U9899 (N_9899,N_9035,N_9397);
nand U9900 (N_9900,N_9596,N_9091);
nor U9901 (N_9901,N_9317,N_9072);
nor U9902 (N_9902,N_9725,N_9351);
and U9903 (N_9903,N_9251,N_9267);
xnor U9904 (N_9904,N_9232,N_9239);
nand U9905 (N_9905,N_9548,N_9169);
xor U9906 (N_9906,N_9468,N_9069);
nor U9907 (N_9907,N_9237,N_9612);
xor U9908 (N_9908,N_9115,N_9579);
nor U9909 (N_9909,N_9235,N_9477);
and U9910 (N_9910,N_9655,N_9048);
and U9911 (N_9911,N_9559,N_9586);
nand U9912 (N_9912,N_9390,N_9460);
or U9913 (N_9913,N_9410,N_9245);
xor U9914 (N_9914,N_9246,N_9151);
nand U9915 (N_9915,N_9309,N_9696);
xnor U9916 (N_9916,N_9202,N_9121);
nor U9917 (N_9917,N_9255,N_9738);
or U9918 (N_9918,N_9565,N_9574);
nor U9919 (N_9919,N_9041,N_9381);
or U9920 (N_9920,N_9684,N_9348);
or U9921 (N_9921,N_9346,N_9631);
or U9922 (N_9922,N_9034,N_9128);
xnor U9923 (N_9923,N_9685,N_9060);
nor U9924 (N_9924,N_9312,N_9195);
nor U9925 (N_9925,N_9464,N_9225);
or U9926 (N_9926,N_9650,N_9104);
and U9927 (N_9927,N_9219,N_9551);
or U9928 (N_9928,N_9203,N_9199);
and U9929 (N_9929,N_9085,N_9002);
xnor U9930 (N_9930,N_9039,N_9730);
or U9931 (N_9931,N_9028,N_9204);
nand U9932 (N_9932,N_9661,N_9569);
and U9933 (N_9933,N_9145,N_9254);
and U9934 (N_9934,N_9183,N_9742);
xor U9935 (N_9935,N_9303,N_9702);
or U9936 (N_9936,N_9012,N_9593);
nand U9937 (N_9937,N_9537,N_9168);
or U9938 (N_9938,N_9355,N_9181);
nor U9939 (N_9939,N_9698,N_9613);
nor U9940 (N_9940,N_9172,N_9705);
and U9941 (N_9941,N_9111,N_9371);
nor U9942 (N_9942,N_9142,N_9577);
nand U9943 (N_9943,N_9298,N_9456);
xnor U9944 (N_9944,N_9277,N_9260);
nor U9945 (N_9945,N_9360,N_9207);
and U9946 (N_9946,N_9045,N_9016);
nand U9947 (N_9947,N_9057,N_9213);
and U9948 (N_9948,N_9319,N_9668);
nor U9949 (N_9949,N_9332,N_9566);
or U9950 (N_9950,N_9516,N_9006);
nor U9951 (N_9951,N_9436,N_9677);
or U9952 (N_9952,N_9643,N_9584);
nand U9953 (N_9953,N_9533,N_9605);
nand U9954 (N_9954,N_9472,N_9003);
nor U9955 (N_9955,N_9611,N_9413);
or U9956 (N_9956,N_9420,N_9621);
or U9957 (N_9957,N_9090,N_9368);
and U9958 (N_9958,N_9709,N_9137);
nand U9959 (N_9959,N_9496,N_9064);
xor U9960 (N_9960,N_9502,N_9015);
xnor U9961 (N_9961,N_9311,N_9356);
nand U9962 (N_9962,N_9096,N_9314);
and U9963 (N_9963,N_9377,N_9672);
nor U9964 (N_9964,N_9640,N_9117);
xor U9965 (N_9965,N_9645,N_9659);
xor U9966 (N_9966,N_9324,N_9165);
nand U9967 (N_9967,N_9270,N_9171);
nor U9968 (N_9968,N_9610,N_9221);
or U9969 (N_9969,N_9330,N_9114);
nor U9970 (N_9970,N_9475,N_9253);
nand U9971 (N_9971,N_9737,N_9320);
and U9972 (N_9972,N_9508,N_9102);
nand U9973 (N_9973,N_9447,N_9369);
and U9974 (N_9974,N_9278,N_9257);
nor U9975 (N_9975,N_9721,N_9304);
xnor U9976 (N_9976,N_9515,N_9723);
xor U9977 (N_9977,N_9120,N_9170);
nor U9978 (N_9978,N_9546,N_9079);
or U9979 (N_9979,N_9673,N_9455);
or U9980 (N_9980,N_9726,N_9522);
and U9981 (N_9981,N_9540,N_9290);
or U9982 (N_9982,N_9438,N_9454);
xnor U9983 (N_9983,N_9718,N_9396);
and U9984 (N_9984,N_9527,N_9344);
nand U9985 (N_9985,N_9132,N_9296);
and U9986 (N_9986,N_9155,N_9051);
xnor U9987 (N_9987,N_9506,N_9536);
nor U9988 (N_9988,N_9354,N_9651);
and U9989 (N_9989,N_9224,N_9244);
nor U9990 (N_9990,N_9389,N_9341);
nor U9991 (N_9991,N_9009,N_9656);
nor U9992 (N_9992,N_9520,N_9308);
and U9993 (N_9993,N_9746,N_9082);
and U9994 (N_9994,N_9157,N_9178);
and U9995 (N_9995,N_9164,N_9401);
and U9996 (N_9996,N_9055,N_9731);
or U9997 (N_9997,N_9638,N_9739);
and U9998 (N_9998,N_9166,N_9100);
or U9999 (N_9999,N_9435,N_9380);
and U10000 (N_10000,N_9078,N_9600);
xor U10001 (N_10001,N_9667,N_9184);
or U10002 (N_10002,N_9387,N_9013);
nor U10003 (N_10003,N_9180,N_9622);
or U10004 (N_10004,N_9437,N_9274);
and U10005 (N_10005,N_9409,N_9604);
or U10006 (N_10006,N_9582,N_9590);
or U10007 (N_10007,N_9391,N_9732);
or U10008 (N_10008,N_9429,N_9544);
nand U10009 (N_10009,N_9361,N_9315);
nor U10010 (N_10010,N_9153,N_9363);
nor U10011 (N_10011,N_9196,N_9228);
xnor U10012 (N_10012,N_9517,N_9609);
xnor U10013 (N_10013,N_9146,N_9509);
nor U10014 (N_10014,N_9688,N_9266);
nor U10015 (N_10015,N_9470,N_9443);
xnor U10016 (N_10016,N_9150,N_9076);
and U10017 (N_10017,N_9214,N_9135);
nor U10018 (N_10018,N_9557,N_9549);
nor U10019 (N_10019,N_9724,N_9550);
nand U10020 (N_10020,N_9703,N_9322);
and U10021 (N_10021,N_9701,N_9179);
xnor U10022 (N_10022,N_9697,N_9649);
xnor U10023 (N_10023,N_9426,N_9606);
xor U10024 (N_10024,N_9326,N_9384);
and U10025 (N_10025,N_9226,N_9494);
nand U10026 (N_10026,N_9652,N_9394);
xor U10027 (N_10027,N_9660,N_9728);
and U10028 (N_10028,N_9095,N_9162);
or U10029 (N_10029,N_9713,N_9706);
or U10030 (N_10030,N_9513,N_9335);
or U10031 (N_10031,N_9745,N_9647);
and U10032 (N_10032,N_9018,N_9616);
or U10033 (N_10033,N_9318,N_9042);
nand U10034 (N_10034,N_9521,N_9458);
and U10035 (N_10035,N_9340,N_9046);
nand U10036 (N_10036,N_9674,N_9467);
nor U10037 (N_10037,N_9291,N_9482);
nand U10038 (N_10038,N_9449,N_9059);
and U10039 (N_10039,N_9065,N_9561);
nor U10040 (N_10040,N_9699,N_9359);
xnor U10041 (N_10041,N_9210,N_9019);
and U10042 (N_10042,N_9268,N_9343);
or U10043 (N_10043,N_9587,N_9010);
nand U10044 (N_10044,N_9476,N_9694);
xnor U10045 (N_10045,N_9570,N_9129);
nand U10046 (N_10046,N_9070,N_9539);
and U10047 (N_10047,N_9388,N_9711);
or U10048 (N_10048,N_9167,N_9452);
nor U10049 (N_10049,N_9415,N_9163);
nor U10050 (N_10050,N_9504,N_9740);
or U10051 (N_10051,N_9716,N_9634);
or U10052 (N_10052,N_9021,N_9238);
nand U10053 (N_10053,N_9139,N_9722);
and U10054 (N_10054,N_9258,N_9451);
nand U10055 (N_10055,N_9297,N_9261);
or U10056 (N_10056,N_9372,N_9747);
nor U10057 (N_10057,N_9692,N_9541);
or U10058 (N_10058,N_9608,N_9271);
nand U10059 (N_10059,N_9431,N_9402);
xor U10060 (N_10060,N_9159,N_9603);
xnor U10061 (N_10061,N_9113,N_9288);
nor U10062 (N_10062,N_9664,N_9081);
and U10063 (N_10063,N_9395,N_9492);
or U10064 (N_10064,N_9704,N_9177);
nand U10065 (N_10065,N_9690,N_9077);
and U10066 (N_10066,N_9175,N_9032);
nor U10067 (N_10067,N_9127,N_9192);
nor U10068 (N_10068,N_9399,N_9282);
xnor U10069 (N_10069,N_9727,N_9627);
nor U10070 (N_10070,N_9265,N_9635);
or U10071 (N_10071,N_9720,N_9337);
xnor U10072 (N_10072,N_9050,N_9092);
or U10073 (N_10073,N_9683,N_9126);
nand U10074 (N_10074,N_9530,N_9004);
and U10075 (N_10075,N_9144,N_9490);
or U10076 (N_10076,N_9123,N_9382);
nor U10077 (N_10077,N_9099,N_9325);
xnor U10078 (N_10078,N_9053,N_9279);
and U10079 (N_10079,N_9441,N_9295);
nand U10080 (N_10080,N_9014,N_9524);
xor U10081 (N_10081,N_9666,N_9054);
nor U10082 (N_10082,N_9347,N_9445);
nor U10083 (N_10083,N_9403,N_9427);
xnor U10084 (N_10084,N_9658,N_9457);
or U10085 (N_10085,N_9534,N_9642);
and U10086 (N_10086,N_9106,N_9216);
and U10087 (N_10087,N_9473,N_9349);
xor U10088 (N_10088,N_9243,N_9305);
and U10089 (N_10089,N_9071,N_9529);
xor U10090 (N_10090,N_9414,N_9301);
nand U10091 (N_10091,N_9223,N_9448);
nor U10092 (N_10092,N_9654,N_9040);
and U10093 (N_10093,N_9220,N_9289);
and U10094 (N_10094,N_9741,N_9201);
nand U10095 (N_10095,N_9234,N_9038);
nand U10096 (N_10096,N_9573,N_9479);
xnor U10097 (N_10097,N_9400,N_9629);
and U10098 (N_10098,N_9374,N_9370);
xor U10099 (N_10099,N_9376,N_9350);
or U10100 (N_10100,N_9568,N_9430);
xnor U10101 (N_10101,N_9499,N_9197);
nand U10102 (N_10102,N_9495,N_9188);
or U10103 (N_10103,N_9483,N_9001);
or U10104 (N_10104,N_9250,N_9450);
nor U10105 (N_10105,N_9122,N_9412);
or U10106 (N_10106,N_9686,N_9444);
or U10107 (N_10107,N_9523,N_9058);
nor U10108 (N_10108,N_9597,N_9276);
nand U10109 (N_10109,N_9471,N_9147);
nor U10110 (N_10110,N_9084,N_9624);
nand U10111 (N_10111,N_9602,N_9068);
nand U10112 (N_10112,N_9626,N_9148);
and U10113 (N_10113,N_9567,N_9623);
or U10114 (N_10114,N_9657,N_9031);
xor U10115 (N_10115,N_9607,N_9619);
nor U10116 (N_10116,N_9729,N_9264);
and U10117 (N_10117,N_9005,N_9591);
xnor U10118 (N_10118,N_9601,N_9073);
nor U10119 (N_10119,N_9526,N_9185);
xor U10120 (N_10120,N_9484,N_9365);
or U10121 (N_10121,N_9158,N_9011);
or U10122 (N_10122,N_9563,N_9023);
or U10123 (N_10123,N_9493,N_9576);
nor U10124 (N_10124,N_9191,N_9200);
and U10125 (N_10125,N_9235,N_9280);
and U10126 (N_10126,N_9021,N_9638);
and U10127 (N_10127,N_9546,N_9051);
nor U10128 (N_10128,N_9356,N_9501);
nor U10129 (N_10129,N_9079,N_9748);
or U10130 (N_10130,N_9599,N_9279);
nor U10131 (N_10131,N_9179,N_9649);
nor U10132 (N_10132,N_9616,N_9343);
xnor U10133 (N_10133,N_9240,N_9670);
or U10134 (N_10134,N_9483,N_9008);
and U10135 (N_10135,N_9510,N_9064);
nor U10136 (N_10136,N_9535,N_9676);
and U10137 (N_10137,N_9188,N_9654);
nor U10138 (N_10138,N_9634,N_9215);
xor U10139 (N_10139,N_9606,N_9257);
xor U10140 (N_10140,N_9328,N_9422);
nor U10141 (N_10141,N_9271,N_9187);
or U10142 (N_10142,N_9100,N_9496);
and U10143 (N_10143,N_9601,N_9499);
and U10144 (N_10144,N_9657,N_9012);
nor U10145 (N_10145,N_9344,N_9580);
nand U10146 (N_10146,N_9212,N_9350);
nor U10147 (N_10147,N_9458,N_9630);
nand U10148 (N_10148,N_9690,N_9362);
and U10149 (N_10149,N_9203,N_9106);
nor U10150 (N_10150,N_9006,N_9434);
and U10151 (N_10151,N_9474,N_9634);
nand U10152 (N_10152,N_9507,N_9405);
xnor U10153 (N_10153,N_9590,N_9462);
and U10154 (N_10154,N_9403,N_9277);
nor U10155 (N_10155,N_9074,N_9564);
and U10156 (N_10156,N_9519,N_9613);
or U10157 (N_10157,N_9452,N_9357);
and U10158 (N_10158,N_9243,N_9589);
and U10159 (N_10159,N_9685,N_9160);
or U10160 (N_10160,N_9480,N_9624);
xnor U10161 (N_10161,N_9312,N_9191);
or U10162 (N_10162,N_9249,N_9296);
or U10163 (N_10163,N_9170,N_9455);
nor U10164 (N_10164,N_9369,N_9078);
or U10165 (N_10165,N_9078,N_9453);
or U10166 (N_10166,N_9202,N_9683);
nor U10167 (N_10167,N_9293,N_9325);
xnor U10168 (N_10168,N_9646,N_9597);
or U10169 (N_10169,N_9609,N_9339);
nor U10170 (N_10170,N_9645,N_9697);
or U10171 (N_10171,N_9655,N_9031);
and U10172 (N_10172,N_9458,N_9520);
nor U10173 (N_10173,N_9195,N_9046);
or U10174 (N_10174,N_9356,N_9577);
and U10175 (N_10175,N_9227,N_9055);
nor U10176 (N_10176,N_9271,N_9299);
nand U10177 (N_10177,N_9099,N_9704);
nor U10178 (N_10178,N_9187,N_9667);
xor U10179 (N_10179,N_9650,N_9153);
nor U10180 (N_10180,N_9689,N_9635);
and U10181 (N_10181,N_9007,N_9745);
nand U10182 (N_10182,N_9130,N_9246);
nor U10183 (N_10183,N_9511,N_9451);
nor U10184 (N_10184,N_9689,N_9721);
nor U10185 (N_10185,N_9406,N_9125);
xor U10186 (N_10186,N_9339,N_9447);
or U10187 (N_10187,N_9340,N_9460);
or U10188 (N_10188,N_9189,N_9074);
and U10189 (N_10189,N_9284,N_9034);
xnor U10190 (N_10190,N_9749,N_9131);
and U10191 (N_10191,N_9184,N_9278);
or U10192 (N_10192,N_9028,N_9666);
or U10193 (N_10193,N_9029,N_9436);
nand U10194 (N_10194,N_9649,N_9293);
or U10195 (N_10195,N_9444,N_9397);
and U10196 (N_10196,N_9123,N_9404);
nand U10197 (N_10197,N_9452,N_9500);
xor U10198 (N_10198,N_9505,N_9162);
xnor U10199 (N_10199,N_9575,N_9166);
or U10200 (N_10200,N_9116,N_9439);
or U10201 (N_10201,N_9626,N_9742);
and U10202 (N_10202,N_9056,N_9677);
or U10203 (N_10203,N_9433,N_9047);
and U10204 (N_10204,N_9611,N_9074);
or U10205 (N_10205,N_9749,N_9673);
or U10206 (N_10206,N_9734,N_9183);
or U10207 (N_10207,N_9432,N_9331);
or U10208 (N_10208,N_9673,N_9618);
nor U10209 (N_10209,N_9593,N_9616);
xnor U10210 (N_10210,N_9569,N_9545);
nand U10211 (N_10211,N_9195,N_9040);
and U10212 (N_10212,N_9684,N_9557);
or U10213 (N_10213,N_9335,N_9547);
and U10214 (N_10214,N_9705,N_9427);
nor U10215 (N_10215,N_9530,N_9194);
nand U10216 (N_10216,N_9679,N_9050);
or U10217 (N_10217,N_9000,N_9633);
nor U10218 (N_10218,N_9032,N_9582);
or U10219 (N_10219,N_9697,N_9091);
or U10220 (N_10220,N_9268,N_9368);
and U10221 (N_10221,N_9134,N_9518);
xnor U10222 (N_10222,N_9128,N_9642);
xor U10223 (N_10223,N_9191,N_9375);
xnor U10224 (N_10224,N_9180,N_9359);
nand U10225 (N_10225,N_9097,N_9194);
or U10226 (N_10226,N_9519,N_9693);
nand U10227 (N_10227,N_9573,N_9728);
and U10228 (N_10228,N_9518,N_9748);
or U10229 (N_10229,N_9245,N_9336);
or U10230 (N_10230,N_9486,N_9530);
nand U10231 (N_10231,N_9206,N_9740);
or U10232 (N_10232,N_9345,N_9597);
xor U10233 (N_10233,N_9375,N_9367);
nand U10234 (N_10234,N_9423,N_9339);
or U10235 (N_10235,N_9333,N_9082);
nand U10236 (N_10236,N_9494,N_9063);
xor U10237 (N_10237,N_9676,N_9544);
or U10238 (N_10238,N_9349,N_9228);
xor U10239 (N_10239,N_9178,N_9058);
xor U10240 (N_10240,N_9564,N_9056);
and U10241 (N_10241,N_9301,N_9122);
nor U10242 (N_10242,N_9534,N_9726);
and U10243 (N_10243,N_9410,N_9495);
and U10244 (N_10244,N_9371,N_9692);
nand U10245 (N_10245,N_9049,N_9552);
xor U10246 (N_10246,N_9746,N_9069);
and U10247 (N_10247,N_9393,N_9285);
and U10248 (N_10248,N_9371,N_9595);
xor U10249 (N_10249,N_9427,N_9627);
nand U10250 (N_10250,N_9035,N_9707);
xor U10251 (N_10251,N_9748,N_9738);
or U10252 (N_10252,N_9091,N_9649);
nor U10253 (N_10253,N_9474,N_9697);
nand U10254 (N_10254,N_9527,N_9599);
or U10255 (N_10255,N_9748,N_9530);
nor U10256 (N_10256,N_9059,N_9140);
and U10257 (N_10257,N_9173,N_9004);
and U10258 (N_10258,N_9730,N_9038);
nand U10259 (N_10259,N_9093,N_9168);
nor U10260 (N_10260,N_9264,N_9267);
xnor U10261 (N_10261,N_9273,N_9234);
and U10262 (N_10262,N_9590,N_9718);
xnor U10263 (N_10263,N_9154,N_9063);
nand U10264 (N_10264,N_9681,N_9245);
or U10265 (N_10265,N_9364,N_9069);
xnor U10266 (N_10266,N_9329,N_9525);
or U10267 (N_10267,N_9207,N_9745);
or U10268 (N_10268,N_9569,N_9139);
nor U10269 (N_10269,N_9470,N_9480);
xnor U10270 (N_10270,N_9385,N_9549);
and U10271 (N_10271,N_9579,N_9169);
or U10272 (N_10272,N_9099,N_9214);
and U10273 (N_10273,N_9240,N_9644);
or U10274 (N_10274,N_9666,N_9366);
and U10275 (N_10275,N_9224,N_9148);
and U10276 (N_10276,N_9401,N_9340);
nand U10277 (N_10277,N_9321,N_9676);
nor U10278 (N_10278,N_9065,N_9047);
and U10279 (N_10279,N_9724,N_9002);
nand U10280 (N_10280,N_9151,N_9653);
xor U10281 (N_10281,N_9139,N_9429);
and U10282 (N_10282,N_9094,N_9260);
xnor U10283 (N_10283,N_9511,N_9444);
xor U10284 (N_10284,N_9411,N_9662);
and U10285 (N_10285,N_9292,N_9687);
and U10286 (N_10286,N_9320,N_9547);
and U10287 (N_10287,N_9356,N_9323);
nor U10288 (N_10288,N_9310,N_9676);
nor U10289 (N_10289,N_9143,N_9131);
xnor U10290 (N_10290,N_9153,N_9057);
or U10291 (N_10291,N_9522,N_9228);
xnor U10292 (N_10292,N_9664,N_9673);
nor U10293 (N_10293,N_9748,N_9697);
and U10294 (N_10294,N_9304,N_9185);
and U10295 (N_10295,N_9321,N_9165);
or U10296 (N_10296,N_9092,N_9354);
or U10297 (N_10297,N_9040,N_9380);
nand U10298 (N_10298,N_9118,N_9574);
xor U10299 (N_10299,N_9131,N_9235);
nor U10300 (N_10300,N_9060,N_9433);
nand U10301 (N_10301,N_9049,N_9656);
xnor U10302 (N_10302,N_9263,N_9270);
nand U10303 (N_10303,N_9449,N_9570);
or U10304 (N_10304,N_9617,N_9028);
xnor U10305 (N_10305,N_9319,N_9330);
xnor U10306 (N_10306,N_9029,N_9080);
or U10307 (N_10307,N_9302,N_9744);
nor U10308 (N_10308,N_9229,N_9201);
or U10309 (N_10309,N_9519,N_9537);
nand U10310 (N_10310,N_9487,N_9472);
nor U10311 (N_10311,N_9012,N_9037);
or U10312 (N_10312,N_9176,N_9060);
and U10313 (N_10313,N_9299,N_9456);
xor U10314 (N_10314,N_9443,N_9681);
nand U10315 (N_10315,N_9208,N_9384);
nor U10316 (N_10316,N_9087,N_9318);
nor U10317 (N_10317,N_9541,N_9368);
xnor U10318 (N_10318,N_9749,N_9534);
and U10319 (N_10319,N_9043,N_9475);
nand U10320 (N_10320,N_9306,N_9704);
and U10321 (N_10321,N_9705,N_9220);
and U10322 (N_10322,N_9551,N_9431);
nor U10323 (N_10323,N_9165,N_9221);
nand U10324 (N_10324,N_9520,N_9287);
or U10325 (N_10325,N_9428,N_9021);
nor U10326 (N_10326,N_9592,N_9101);
and U10327 (N_10327,N_9294,N_9407);
or U10328 (N_10328,N_9234,N_9422);
or U10329 (N_10329,N_9664,N_9176);
nand U10330 (N_10330,N_9442,N_9060);
or U10331 (N_10331,N_9556,N_9383);
nand U10332 (N_10332,N_9725,N_9236);
and U10333 (N_10333,N_9060,N_9347);
nor U10334 (N_10334,N_9433,N_9655);
nand U10335 (N_10335,N_9158,N_9615);
nor U10336 (N_10336,N_9415,N_9649);
or U10337 (N_10337,N_9543,N_9707);
or U10338 (N_10338,N_9627,N_9092);
nand U10339 (N_10339,N_9731,N_9095);
xor U10340 (N_10340,N_9633,N_9261);
xnor U10341 (N_10341,N_9702,N_9572);
nand U10342 (N_10342,N_9130,N_9747);
and U10343 (N_10343,N_9445,N_9253);
and U10344 (N_10344,N_9253,N_9352);
xor U10345 (N_10345,N_9266,N_9006);
xnor U10346 (N_10346,N_9062,N_9550);
or U10347 (N_10347,N_9461,N_9174);
nor U10348 (N_10348,N_9206,N_9281);
nand U10349 (N_10349,N_9284,N_9638);
or U10350 (N_10350,N_9215,N_9309);
nor U10351 (N_10351,N_9656,N_9120);
nand U10352 (N_10352,N_9399,N_9333);
nor U10353 (N_10353,N_9415,N_9319);
or U10354 (N_10354,N_9451,N_9118);
or U10355 (N_10355,N_9698,N_9557);
and U10356 (N_10356,N_9435,N_9731);
nand U10357 (N_10357,N_9539,N_9352);
or U10358 (N_10358,N_9104,N_9251);
or U10359 (N_10359,N_9145,N_9481);
and U10360 (N_10360,N_9228,N_9724);
nor U10361 (N_10361,N_9662,N_9436);
xor U10362 (N_10362,N_9077,N_9719);
nand U10363 (N_10363,N_9186,N_9087);
and U10364 (N_10364,N_9426,N_9008);
xor U10365 (N_10365,N_9072,N_9467);
nor U10366 (N_10366,N_9192,N_9341);
or U10367 (N_10367,N_9140,N_9075);
and U10368 (N_10368,N_9453,N_9135);
xor U10369 (N_10369,N_9654,N_9128);
or U10370 (N_10370,N_9265,N_9197);
xnor U10371 (N_10371,N_9700,N_9521);
nand U10372 (N_10372,N_9095,N_9268);
nor U10373 (N_10373,N_9514,N_9395);
nand U10374 (N_10374,N_9453,N_9286);
nand U10375 (N_10375,N_9187,N_9332);
xnor U10376 (N_10376,N_9431,N_9076);
or U10377 (N_10377,N_9598,N_9514);
and U10378 (N_10378,N_9343,N_9685);
or U10379 (N_10379,N_9082,N_9121);
nand U10380 (N_10380,N_9020,N_9645);
nand U10381 (N_10381,N_9244,N_9678);
xnor U10382 (N_10382,N_9741,N_9023);
nor U10383 (N_10383,N_9283,N_9138);
xor U10384 (N_10384,N_9170,N_9040);
or U10385 (N_10385,N_9122,N_9286);
or U10386 (N_10386,N_9391,N_9589);
and U10387 (N_10387,N_9557,N_9235);
nand U10388 (N_10388,N_9626,N_9238);
nand U10389 (N_10389,N_9566,N_9432);
nor U10390 (N_10390,N_9136,N_9614);
nand U10391 (N_10391,N_9088,N_9537);
nand U10392 (N_10392,N_9655,N_9314);
xnor U10393 (N_10393,N_9639,N_9568);
nand U10394 (N_10394,N_9398,N_9137);
or U10395 (N_10395,N_9542,N_9409);
xor U10396 (N_10396,N_9440,N_9687);
or U10397 (N_10397,N_9535,N_9163);
and U10398 (N_10398,N_9030,N_9471);
nand U10399 (N_10399,N_9566,N_9666);
nand U10400 (N_10400,N_9217,N_9602);
nand U10401 (N_10401,N_9473,N_9308);
nor U10402 (N_10402,N_9723,N_9676);
nor U10403 (N_10403,N_9496,N_9462);
nand U10404 (N_10404,N_9502,N_9437);
xor U10405 (N_10405,N_9375,N_9456);
nor U10406 (N_10406,N_9595,N_9627);
and U10407 (N_10407,N_9627,N_9606);
xor U10408 (N_10408,N_9701,N_9153);
nor U10409 (N_10409,N_9309,N_9221);
nand U10410 (N_10410,N_9626,N_9361);
and U10411 (N_10411,N_9360,N_9447);
nand U10412 (N_10412,N_9524,N_9747);
and U10413 (N_10413,N_9365,N_9253);
nor U10414 (N_10414,N_9460,N_9608);
or U10415 (N_10415,N_9304,N_9361);
or U10416 (N_10416,N_9724,N_9306);
or U10417 (N_10417,N_9177,N_9093);
and U10418 (N_10418,N_9176,N_9526);
nor U10419 (N_10419,N_9165,N_9408);
and U10420 (N_10420,N_9656,N_9269);
or U10421 (N_10421,N_9380,N_9534);
and U10422 (N_10422,N_9230,N_9584);
and U10423 (N_10423,N_9644,N_9536);
xor U10424 (N_10424,N_9205,N_9229);
and U10425 (N_10425,N_9230,N_9672);
xor U10426 (N_10426,N_9210,N_9087);
xor U10427 (N_10427,N_9520,N_9341);
nand U10428 (N_10428,N_9114,N_9384);
nand U10429 (N_10429,N_9437,N_9689);
nor U10430 (N_10430,N_9204,N_9093);
nor U10431 (N_10431,N_9640,N_9108);
xnor U10432 (N_10432,N_9435,N_9584);
nor U10433 (N_10433,N_9744,N_9499);
and U10434 (N_10434,N_9251,N_9342);
or U10435 (N_10435,N_9400,N_9320);
xor U10436 (N_10436,N_9076,N_9718);
nor U10437 (N_10437,N_9472,N_9502);
nand U10438 (N_10438,N_9290,N_9719);
xnor U10439 (N_10439,N_9315,N_9683);
nand U10440 (N_10440,N_9705,N_9649);
nand U10441 (N_10441,N_9722,N_9239);
nor U10442 (N_10442,N_9142,N_9655);
xnor U10443 (N_10443,N_9288,N_9061);
and U10444 (N_10444,N_9323,N_9339);
xnor U10445 (N_10445,N_9258,N_9216);
xor U10446 (N_10446,N_9196,N_9389);
and U10447 (N_10447,N_9635,N_9734);
nand U10448 (N_10448,N_9160,N_9496);
nor U10449 (N_10449,N_9055,N_9385);
or U10450 (N_10450,N_9402,N_9667);
or U10451 (N_10451,N_9304,N_9109);
or U10452 (N_10452,N_9320,N_9254);
nor U10453 (N_10453,N_9345,N_9294);
nor U10454 (N_10454,N_9604,N_9023);
or U10455 (N_10455,N_9568,N_9124);
xor U10456 (N_10456,N_9055,N_9450);
xnor U10457 (N_10457,N_9720,N_9400);
nor U10458 (N_10458,N_9065,N_9148);
or U10459 (N_10459,N_9309,N_9041);
nand U10460 (N_10460,N_9114,N_9569);
xnor U10461 (N_10461,N_9216,N_9310);
xnor U10462 (N_10462,N_9500,N_9545);
xor U10463 (N_10463,N_9052,N_9414);
xor U10464 (N_10464,N_9049,N_9370);
or U10465 (N_10465,N_9434,N_9214);
and U10466 (N_10466,N_9247,N_9056);
xor U10467 (N_10467,N_9324,N_9433);
and U10468 (N_10468,N_9234,N_9209);
nand U10469 (N_10469,N_9651,N_9664);
or U10470 (N_10470,N_9469,N_9535);
or U10471 (N_10471,N_9287,N_9669);
nor U10472 (N_10472,N_9676,N_9691);
and U10473 (N_10473,N_9031,N_9237);
nand U10474 (N_10474,N_9711,N_9286);
xor U10475 (N_10475,N_9588,N_9645);
nand U10476 (N_10476,N_9365,N_9093);
xor U10477 (N_10477,N_9178,N_9429);
or U10478 (N_10478,N_9342,N_9180);
nor U10479 (N_10479,N_9149,N_9092);
nor U10480 (N_10480,N_9380,N_9577);
nand U10481 (N_10481,N_9267,N_9283);
and U10482 (N_10482,N_9184,N_9107);
and U10483 (N_10483,N_9513,N_9101);
xnor U10484 (N_10484,N_9383,N_9439);
nand U10485 (N_10485,N_9003,N_9636);
nor U10486 (N_10486,N_9563,N_9159);
nand U10487 (N_10487,N_9096,N_9582);
and U10488 (N_10488,N_9454,N_9742);
nor U10489 (N_10489,N_9043,N_9280);
xnor U10490 (N_10490,N_9159,N_9574);
xnor U10491 (N_10491,N_9454,N_9551);
xor U10492 (N_10492,N_9464,N_9361);
nand U10493 (N_10493,N_9299,N_9412);
or U10494 (N_10494,N_9745,N_9706);
xor U10495 (N_10495,N_9736,N_9324);
xnor U10496 (N_10496,N_9614,N_9150);
and U10497 (N_10497,N_9282,N_9129);
xor U10498 (N_10498,N_9104,N_9246);
and U10499 (N_10499,N_9717,N_9106);
xnor U10500 (N_10500,N_9799,N_9855);
and U10501 (N_10501,N_10408,N_9870);
xnor U10502 (N_10502,N_10456,N_10046);
or U10503 (N_10503,N_10334,N_10471);
xnor U10504 (N_10504,N_10433,N_10427);
and U10505 (N_10505,N_10116,N_9754);
or U10506 (N_10506,N_9859,N_9965);
and U10507 (N_10507,N_10093,N_10118);
nand U10508 (N_10508,N_9789,N_9922);
and U10509 (N_10509,N_9876,N_10249);
or U10510 (N_10510,N_10054,N_10250);
and U10511 (N_10511,N_9982,N_9814);
nor U10512 (N_10512,N_10404,N_9984);
or U10513 (N_10513,N_10181,N_10104);
nor U10514 (N_10514,N_9832,N_10322);
nor U10515 (N_10515,N_10102,N_10390);
xor U10516 (N_10516,N_10360,N_10470);
and U10517 (N_10517,N_10119,N_10167);
xnor U10518 (N_10518,N_10414,N_10256);
nor U10519 (N_10519,N_10371,N_9875);
and U10520 (N_10520,N_9867,N_9810);
or U10521 (N_10521,N_10124,N_10420);
and U10522 (N_10522,N_10346,N_10154);
nand U10523 (N_10523,N_9800,N_9844);
nor U10524 (N_10524,N_9991,N_10342);
or U10525 (N_10525,N_10105,N_10171);
or U10526 (N_10526,N_10425,N_10444);
xor U10527 (N_10527,N_10279,N_10278);
or U10528 (N_10528,N_10143,N_10228);
or U10529 (N_10529,N_10293,N_10125);
or U10530 (N_10530,N_10035,N_9757);
xnor U10531 (N_10531,N_9807,N_9999);
or U10532 (N_10532,N_9821,N_10103);
and U10533 (N_10533,N_9798,N_10101);
or U10534 (N_10534,N_10262,N_10029);
or U10535 (N_10535,N_9804,N_9981);
or U10536 (N_10536,N_10336,N_10384);
or U10537 (N_10537,N_9938,N_9921);
nand U10538 (N_10538,N_10198,N_10481);
nor U10539 (N_10539,N_10255,N_9934);
and U10540 (N_10540,N_9881,N_9928);
or U10541 (N_10541,N_9911,N_10237);
and U10542 (N_10542,N_9899,N_10146);
nand U10543 (N_10543,N_10277,N_10373);
and U10544 (N_10544,N_10487,N_10350);
or U10545 (N_10545,N_9978,N_9846);
or U10546 (N_10546,N_10288,N_9910);
and U10547 (N_10547,N_9772,N_10396);
nor U10548 (N_10548,N_10012,N_10276);
nor U10549 (N_10549,N_10151,N_10202);
xor U10550 (N_10550,N_10023,N_9949);
nor U10551 (N_10551,N_10068,N_10362);
nand U10552 (N_10552,N_9963,N_10159);
and U10553 (N_10553,N_10494,N_10193);
and U10554 (N_10554,N_10061,N_9823);
nor U10555 (N_10555,N_10482,N_9880);
and U10556 (N_10556,N_10285,N_10324);
nor U10557 (N_10557,N_10440,N_10439);
nor U10558 (N_10558,N_10331,N_9847);
or U10559 (N_10559,N_10127,N_10109);
and U10560 (N_10560,N_9784,N_9979);
nand U10561 (N_10561,N_10473,N_9780);
or U10562 (N_10562,N_9883,N_9926);
xor U10563 (N_10563,N_10480,N_10370);
nand U10564 (N_10564,N_10187,N_10260);
or U10565 (N_10565,N_9851,N_10015);
and U10566 (N_10566,N_9994,N_10131);
xor U10567 (N_10567,N_10424,N_9761);
nand U10568 (N_10568,N_10483,N_9808);
or U10569 (N_10569,N_10095,N_10436);
or U10570 (N_10570,N_10087,N_9861);
nor U10571 (N_10571,N_10156,N_10295);
and U10572 (N_10572,N_10066,N_10382);
xnor U10573 (N_10573,N_9886,N_10098);
or U10574 (N_10574,N_10429,N_10273);
xor U10575 (N_10575,N_10168,N_9763);
or U10576 (N_10576,N_10438,N_10174);
nor U10577 (N_10577,N_10430,N_10451);
or U10578 (N_10578,N_9774,N_10311);
and U10579 (N_10579,N_9948,N_10008);
nor U10580 (N_10580,N_10137,N_10050);
nor U10581 (N_10581,N_10217,N_10020);
nand U10582 (N_10582,N_10327,N_9898);
and U10583 (N_10583,N_10234,N_10345);
or U10584 (N_10584,N_9888,N_10163);
xnor U10585 (N_10585,N_9900,N_10166);
nand U10586 (N_10586,N_10199,N_9819);
or U10587 (N_10587,N_10180,N_9970);
nor U10588 (N_10588,N_10085,N_10075);
or U10589 (N_10589,N_9782,N_10107);
nand U10590 (N_10590,N_10259,N_10343);
nand U10591 (N_10591,N_10405,N_9767);
nand U10592 (N_10592,N_10441,N_9751);
and U10593 (N_10593,N_10197,N_10465);
xor U10594 (N_10594,N_10325,N_9943);
or U10595 (N_10595,N_10333,N_10056);
and U10596 (N_10596,N_9904,N_10241);
nor U10597 (N_10597,N_10129,N_9936);
nor U10598 (N_10598,N_9818,N_9887);
or U10599 (N_10599,N_9929,N_10375);
nand U10600 (N_10600,N_9765,N_10144);
nand U10601 (N_10601,N_10263,N_9750);
or U10602 (N_10602,N_10200,N_9903);
xor U10603 (N_10603,N_10286,N_10491);
nor U10604 (N_10604,N_9897,N_10296);
xor U10605 (N_10605,N_10120,N_10352);
and U10606 (N_10606,N_10062,N_10123);
nor U10607 (N_10607,N_10211,N_9977);
xor U10608 (N_10608,N_10460,N_10178);
or U10609 (N_10609,N_10128,N_10317);
nand U10610 (N_10610,N_10206,N_10496);
nor U10611 (N_10611,N_10314,N_9985);
xnor U10612 (N_10612,N_10358,N_10052);
nand U10613 (N_10613,N_10431,N_10133);
nor U10614 (N_10614,N_9838,N_10138);
xor U10615 (N_10615,N_10416,N_9918);
nand U10616 (N_10616,N_9996,N_10157);
nand U10617 (N_10617,N_9775,N_10239);
and U10618 (N_10618,N_9895,N_10114);
nor U10619 (N_10619,N_9891,N_9988);
or U10620 (N_10620,N_9873,N_9783);
nand U10621 (N_10621,N_10215,N_10274);
and U10622 (N_10622,N_10039,N_9995);
xor U10623 (N_10623,N_9860,N_9872);
and U10624 (N_10624,N_10303,N_10486);
or U10625 (N_10625,N_10339,N_10022);
nor U10626 (N_10626,N_9840,N_9952);
nand U10627 (N_10627,N_10484,N_9796);
nand U10628 (N_10628,N_9762,N_9964);
nor U10629 (N_10629,N_10363,N_10057);
xnor U10630 (N_10630,N_10415,N_10300);
or U10631 (N_10631,N_10089,N_10380);
nand U10632 (N_10632,N_9935,N_10160);
xnor U10633 (N_10633,N_9809,N_9769);
and U10634 (N_10634,N_10025,N_10489);
nor U10635 (N_10635,N_10446,N_9824);
and U10636 (N_10636,N_10086,N_10383);
and U10637 (N_10637,N_10495,N_10071);
xor U10638 (N_10638,N_10080,N_10208);
and U10639 (N_10639,N_10267,N_10017);
nor U10640 (N_10640,N_9924,N_9941);
or U10641 (N_10641,N_9820,N_10145);
and U10642 (N_10642,N_9785,N_9885);
xor U10643 (N_10643,N_10497,N_9892);
or U10644 (N_10644,N_9925,N_10176);
xnor U10645 (N_10645,N_9986,N_10328);
or U10646 (N_10646,N_9972,N_10078);
nand U10647 (N_10647,N_10185,N_10379);
nor U10648 (N_10648,N_10353,N_9779);
and U10649 (N_10649,N_10310,N_10398);
nor U10650 (N_10650,N_10281,N_9768);
nand U10651 (N_10651,N_10329,N_10388);
and U10652 (N_10652,N_10448,N_10304);
and U10653 (N_10653,N_9753,N_10203);
xnor U10654 (N_10654,N_10077,N_10407);
and U10655 (N_10655,N_10361,N_10065);
nor U10656 (N_10656,N_10338,N_9912);
xnor U10657 (N_10657,N_10306,N_10014);
or U10658 (N_10658,N_10209,N_10240);
or U10659 (N_10659,N_10115,N_10266);
and U10660 (N_10660,N_10347,N_10386);
nand U10661 (N_10661,N_10401,N_10148);
or U10662 (N_10662,N_9795,N_9976);
nand U10663 (N_10663,N_10063,N_10437);
and U10664 (N_10664,N_10009,N_10454);
or U10665 (N_10665,N_10140,N_10399);
xor U10666 (N_10666,N_10195,N_10011);
or U10667 (N_10667,N_10218,N_10091);
or U10668 (N_10668,N_10452,N_10447);
nand U10669 (N_10669,N_10485,N_9901);
or U10670 (N_10670,N_10330,N_10257);
nor U10671 (N_10671,N_9955,N_9961);
nand U10672 (N_10672,N_10368,N_10292);
and U10673 (N_10673,N_10397,N_9940);
and U10674 (N_10674,N_9834,N_10268);
nand U10675 (N_10675,N_10254,N_10376);
and U10676 (N_10676,N_10030,N_10182);
and U10677 (N_10677,N_10130,N_10337);
and U10678 (N_10678,N_10214,N_10088);
nor U10679 (N_10679,N_9833,N_10003);
and U10680 (N_10680,N_9848,N_9869);
nor U10681 (N_10681,N_9945,N_10313);
nand U10682 (N_10682,N_10097,N_10391);
xor U10683 (N_10683,N_10179,N_10122);
nor U10684 (N_10684,N_10172,N_9917);
or U10685 (N_10685,N_10434,N_10142);
nand U10686 (N_10686,N_10018,N_10196);
or U10687 (N_10687,N_10323,N_9905);
xnor U10688 (N_10688,N_9954,N_10192);
nand U10689 (N_10689,N_10301,N_9831);
or U10690 (N_10690,N_10287,N_10340);
nor U10691 (N_10691,N_10139,N_10040);
xnor U10692 (N_10692,N_10402,N_9865);
xnor U10693 (N_10693,N_10016,N_10147);
or U10694 (N_10694,N_10070,N_9813);
nand U10695 (N_10695,N_9790,N_10344);
xor U10696 (N_10696,N_10406,N_9990);
and U10697 (N_10697,N_10058,N_10302);
xnor U10698 (N_10698,N_10479,N_10270);
and U10699 (N_10699,N_10422,N_10466);
xor U10700 (N_10700,N_10072,N_10136);
xnor U10701 (N_10701,N_10213,N_10175);
nor U10702 (N_10702,N_9882,N_10341);
nor U10703 (N_10703,N_10449,N_10488);
xor U10704 (N_10704,N_10162,N_10069);
nand U10705 (N_10705,N_9956,N_10001);
nand U10706 (N_10706,N_9778,N_9946);
and U10707 (N_10707,N_10443,N_9913);
and U10708 (N_10708,N_10442,N_9871);
and U10709 (N_10709,N_9967,N_10423);
or U10710 (N_10710,N_9817,N_10111);
and U10711 (N_10711,N_10280,N_10335);
and U10712 (N_10712,N_10126,N_10045);
nor U10713 (N_10713,N_10076,N_9792);
and U10714 (N_10714,N_10041,N_10221);
nand U10715 (N_10715,N_10364,N_9927);
and U10716 (N_10716,N_10477,N_10369);
and U10717 (N_10717,N_9770,N_10232);
xnor U10718 (N_10718,N_9787,N_10271);
xnor U10719 (N_10719,N_9957,N_10283);
nor U10720 (N_10720,N_10113,N_10026);
nand U10721 (N_10721,N_10349,N_10393);
or U10722 (N_10722,N_10201,N_9966);
and U10723 (N_10723,N_10356,N_10251);
xor U10724 (N_10724,N_9829,N_10064);
nor U10725 (N_10725,N_9802,N_9879);
nor U10726 (N_10726,N_10037,N_10319);
or U10727 (N_10727,N_10298,N_9975);
nor U10728 (N_10728,N_10028,N_10223);
or U10729 (N_10729,N_10153,N_10297);
or U10730 (N_10730,N_9777,N_9858);
and U10731 (N_10731,N_10365,N_9850);
nand U10732 (N_10732,N_9974,N_10212);
nand U10733 (N_10733,N_10459,N_10242);
nand U10734 (N_10734,N_9791,N_10048);
or U10735 (N_10735,N_9868,N_9835);
and U10736 (N_10736,N_10135,N_10269);
nand U10737 (N_10737,N_9878,N_9993);
xor U10738 (N_10738,N_9815,N_10264);
nor U10739 (N_10739,N_10246,N_10258);
and U10740 (N_10740,N_9839,N_9915);
or U10741 (N_10741,N_10235,N_10222);
nand U10742 (N_10742,N_9771,N_10253);
or U10743 (N_10743,N_10161,N_10013);
or U10744 (N_10744,N_10210,N_9786);
nand U10745 (N_10745,N_9801,N_9837);
or U10746 (N_10746,N_9805,N_10117);
nand U10747 (N_10747,N_10073,N_10244);
xor U10748 (N_10748,N_10354,N_10307);
nand U10749 (N_10749,N_9916,N_10165);
nand U10750 (N_10750,N_10252,N_9950);
and U10751 (N_10751,N_10461,N_10445);
xor U10752 (N_10752,N_10121,N_9854);
nand U10753 (N_10753,N_10134,N_10387);
nor U10754 (N_10754,N_9937,N_10090);
nor U10755 (N_10755,N_9960,N_9864);
xnor U10756 (N_10756,N_9797,N_9788);
xnor U10757 (N_10757,N_10469,N_10106);
or U10758 (N_10758,N_10476,N_10261);
and U10759 (N_10759,N_10305,N_9877);
or U10760 (N_10760,N_10010,N_10173);
and U10761 (N_10761,N_10309,N_10410);
nand U10762 (N_10762,N_10315,N_9997);
xnor U10763 (N_10763,N_10395,N_10004);
nor U10764 (N_10764,N_10188,N_10299);
xor U10765 (N_10765,N_10381,N_10060);
nor U10766 (N_10766,N_9793,N_10099);
xor U10767 (N_10767,N_10194,N_9980);
nor U10768 (N_10768,N_10318,N_9755);
nand U10769 (N_10769,N_9842,N_10275);
and U10770 (N_10770,N_10031,N_9983);
nor U10771 (N_10771,N_10458,N_10191);
xor U10772 (N_10772,N_9992,N_10220);
and U10773 (N_10773,N_9914,N_10428);
and U10774 (N_10774,N_9806,N_9825);
and U10775 (N_10775,N_9909,N_10348);
or U10776 (N_10776,N_10049,N_9989);
and U10777 (N_10777,N_9906,N_10006);
nand U10778 (N_10778,N_10230,N_10389);
nand U10779 (N_10779,N_10413,N_9759);
or U10780 (N_10780,N_10282,N_10038);
xor U10781 (N_10781,N_10385,N_10284);
nand U10782 (N_10782,N_10231,N_10411);
nor U10783 (N_10783,N_10499,N_9933);
nor U10784 (N_10784,N_10478,N_9863);
nor U10785 (N_10785,N_10378,N_10094);
xnor U10786 (N_10786,N_10183,N_10490);
xor U10787 (N_10787,N_9845,N_10177);
xor U10788 (N_10788,N_10189,N_9907);
xor U10789 (N_10789,N_10216,N_10034);
or U10790 (N_10790,N_9930,N_9760);
xor U10791 (N_10791,N_9998,N_10374);
or U10792 (N_10792,N_9893,N_9919);
and U10793 (N_10793,N_9920,N_10229);
nand U10794 (N_10794,N_9766,N_10419);
xnor U10795 (N_10795,N_10186,N_10079);
xnor U10796 (N_10796,N_10248,N_9969);
and U10797 (N_10797,N_9781,N_10498);
xor U10798 (N_10798,N_10289,N_10450);
xnor U10799 (N_10799,N_10096,N_9894);
xor U10800 (N_10800,N_10366,N_10108);
and U10801 (N_10801,N_9853,N_9962);
xnor U10802 (N_10802,N_10418,N_10462);
nor U10803 (N_10803,N_9822,N_10372);
nor U10804 (N_10804,N_10455,N_9947);
nor U10805 (N_10805,N_10236,N_10326);
and U10806 (N_10806,N_10081,N_10412);
and U10807 (N_10807,N_9866,N_9902);
nand U10808 (N_10808,N_10021,N_10475);
or U10809 (N_10809,N_10051,N_9828);
nand U10810 (N_10810,N_10463,N_10047);
or U10811 (N_10811,N_10472,N_10074);
nor U10812 (N_10812,N_10320,N_10112);
or U10813 (N_10813,N_10042,N_10019);
or U10814 (N_10814,N_9841,N_9951);
or U10815 (N_10815,N_10272,N_9776);
or U10816 (N_10816,N_9896,N_10492);
nand U10817 (N_10817,N_10150,N_10059);
xor U10818 (N_10818,N_10468,N_10247);
nor U10819 (N_10819,N_10141,N_10421);
xor U10820 (N_10820,N_10357,N_10149);
and U10821 (N_10821,N_9764,N_10392);
and U10822 (N_10822,N_9923,N_9874);
nand U10823 (N_10823,N_9852,N_9890);
nor U10824 (N_10824,N_10243,N_10245);
nand U10825 (N_10825,N_9968,N_10155);
or U10826 (N_10826,N_10053,N_10493);
or U10827 (N_10827,N_10351,N_9884);
xnor U10828 (N_10828,N_10067,N_10294);
nand U10829 (N_10829,N_9987,N_10224);
nand U10830 (N_10830,N_10083,N_10377);
nand U10831 (N_10831,N_10024,N_9752);
or U10832 (N_10832,N_9811,N_9836);
xor U10833 (N_10833,N_10308,N_10238);
xnor U10834 (N_10834,N_9803,N_10227);
nand U10835 (N_10835,N_9856,N_10044);
or U10836 (N_10836,N_10457,N_9889);
nand U10837 (N_10837,N_9830,N_9849);
nand U10838 (N_10838,N_9932,N_9758);
and U10839 (N_10839,N_10409,N_10453);
nand U10840 (N_10840,N_9958,N_9812);
nor U10841 (N_10841,N_10007,N_9942);
xnor U10842 (N_10842,N_10005,N_10082);
and U10843 (N_10843,N_9756,N_9857);
and U10844 (N_10844,N_9862,N_9794);
xnor U10845 (N_10845,N_9908,N_10219);
nand U10846 (N_10846,N_10265,N_10158);
xor U10847 (N_10847,N_10027,N_10132);
xor U10848 (N_10848,N_9931,N_9959);
nor U10849 (N_10849,N_10164,N_10316);
nor U10850 (N_10850,N_10474,N_10055);
xor U10851 (N_10851,N_9826,N_10169);
and U10852 (N_10852,N_10432,N_10225);
xnor U10853 (N_10853,N_10092,N_10036);
xor U10854 (N_10854,N_10207,N_10435);
and U10855 (N_10855,N_9953,N_10170);
xor U10856 (N_10856,N_10002,N_10332);
nand U10857 (N_10857,N_10226,N_10403);
xor U10858 (N_10858,N_9827,N_10290);
or U10859 (N_10859,N_10190,N_9939);
nor U10860 (N_10860,N_9944,N_9971);
and U10861 (N_10861,N_10367,N_10394);
xnor U10862 (N_10862,N_10321,N_10400);
and U10863 (N_10863,N_10464,N_10205);
nor U10864 (N_10864,N_10355,N_10467);
or U10865 (N_10865,N_10233,N_10110);
nor U10866 (N_10866,N_10043,N_10359);
xor U10867 (N_10867,N_10417,N_10000);
or U10868 (N_10868,N_9973,N_9773);
or U10869 (N_10869,N_10032,N_10152);
xor U10870 (N_10870,N_10312,N_10291);
and U10871 (N_10871,N_9816,N_10426);
or U10872 (N_10872,N_10100,N_10033);
or U10873 (N_10873,N_10204,N_10184);
xnor U10874 (N_10874,N_10084,N_9843);
and U10875 (N_10875,N_9971,N_10436);
nor U10876 (N_10876,N_10401,N_10024);
and U10877 (N_10877,N_9804,N_9915);
xor U10878 (N_10878,N_10223,N_10123);
xor U10879 (N_10879,N_10214,N_10374);
nand U10880 (N_10880,N_10045,N_10395);
and U10881 (N_10881,N_10203,N_10190);
and U10882 (N_10882,N_10453,N_10242);
or U10883 (N_10883,N_9818,N_10486);
xnor U10884 (N_10884,N_10312,N_10405);
or U10885 (N_10885,N_10499,N_10215);
and U10886 (N_10886,N_10493,N_10266);
xor U10887 (N_10887,N_10004,N_10075);
xnor U10888 (N_10888,N_10195,N_9962);
and U10889 (N_10889,N_10479,N_10247);
xor U10890 (N_10890,N_9978,N_9921);
nor U10891 (N_10891,N_10169,N_10134);
and U10892 (N_10892,N_9961,N_10407);
and U10893 (N_10893,N_9908,N_10450);
nor U10894 (N_10894,N_9858,N_10167);
nand U10895 (N_10895,N_10219,N_10047);
or U10896 (N_10896,N_10204,N_9970);
and U10897 (N_10897,N_10290,N_9944);
nand U10898 (N_10898,N_9938,N_10000);
xnor U10899 (N_10899,N_10004,N_10215);
xor U10900 (N_10900,N_9854,N_10478);
xor U10901 (N_10901,N_10464,N_9946);
or U10902 (N_10902,N_10328,N_10447);
nand U10903 (N_10903,N_10265,N_10410);
and U10904 (N_10904,N_9864,N_10359);
or U10905 (N_10905,N_10085,N_10015);
or U10906 (N_10906,N_9766,N_9916);
nor U10907 (N_10907,N_10148,N_10166);
or U10908 (N_10908,N_10135,N_10231);
xnor U10909 (N_10909,N_9960,N_10103);
xnor U10910 (N_10910,N_10392,N_10139);
or U10911 (N_10911,N_10159,N_9875);
xnor U10912 (N_10912,N_10281,N_10056);
nand U10913 (N_10913,N_10114,N_10356);
and U10914 (N_10914,N_9982,N_9809);
and U10915 (N_10915,N_10153,N_10274);
or U10916 (N_10916,N_10393,N_10004);
xnor U10917 (N_10917,N_10480,N_9907);
nand U10918 (N_10918,N_9838,N_10095);
nand U10919 (N_10919,N_9784,N_10212);
nand U10920 (N_10920,N_10153,N_9930);
nor U10921 (N_10921,N_10098,N_9820);
nand U10922 (N_10922,N_10263,N_10334);
nand U10923 (N_10923,N_9913,N_10325);
and U10924 (N_10924,N_10498,N_10132);
or U10925 (N_10925,N_10331,N_10287);
nand U10926 (N_10926,N_10313,N_10207);
and U10927 (N_10927,N_9789,N_10159);
nor U10928 (N_10928,N_10376,N_9934);
and U10929 (N_10929,N_9819,N_10079);
nand U10930 (N_10930,N_10008,N_10486);
and U10931 (N_10931,N_10387,N_10390);
nor U10932 (N_10932,N_10098,N_10368);
nor U10933 (N_10933,N_9970,N_9782);
nand U10934 (N_10934,N_10124,N_10070);
nand U10935 (N_10935,N_9866,N_10388);
and U10936 (N_10936,N_10066,N_10394);
or U10937 (N_10937,N_9932,N_10339);
nor U10938 (N_10938,N_9928,N_9998);
xor U10939 (N_10939,N_9971,N_10397);
xnor U10940 (N_10940,N_10137,N_9764);
nor U10941 (N_10941,N_10314,N_10380);
xnor U10942 (N_10942,N_10156,N_10238);
and U10943 (N_10943,N_9975,N_10067);
and U10944 (N_10944,N_10180,N_10081);
xor U10945 (N_10945,N_10148,N_10344);
or U10946 (N_10946,N_10119,N_9920);
and U10947 (N_10947,N_9774,N_10329);
xnor U10948 (N_10948,N_10077,N_10266);
nand U10949 (N_10949,N_10309,N_10202);
nand U10950 (N_10950,N_10173,N_10323);
and U10951 (N_10951,N_10089,N_9774);
nor U10952 (N_10952,N_10317,N_10346);
nand U10953 (N_10953,N_10014,N_9883);
or U10954 (N_10954,N_10440,N_9973);
or U10955 (N_10955,N_10110,N_10063);
or U10956 (N_10956,N_10043,N_10257);
nor U10957 (N_10957,N_10018,N_9803);
or U10958 (N_10958,N_10493,N_10134);
xor U10959 (N_10959,N_10358,N_9772);
xor U10960 (N_10960,N_10065,N_10122);
nor U10961 (N_10961,N_10497,N_10037);
nor U10962 (N_10962,N_10387,N_9789);
and U10963 (N_10963,N_10374,N_9789);
xor U10964 (N_10964,N_10405,N_10145);
xor U10965 (N_10965,N_9986,N_10011);
nor U10966 (N_10966,N_10404,N_10478);
nor U10967 (N_10967,N_10284,N_10384);
nand U10968 (N_10968,N_10413,N_9873);
and U10969 (N_10969,N_10485,N_9763);
xnor U10970 (N_10970,N_10142,N_10043);
nand U10971 (N_10971,N_9861,N_10184);
and U10972 (N_10972,N_9978,N_10266);
nand U10973 (N_10973,N_9883,N_9836);
xor U10974 (N_10974,N_9951,N_10240);
xor U10975 (N_10975,N_9862,N_10174);
nand U10976 (N_10976,N_10487,N_10084);
and U10977 (N_10977,N_10050,N_9955);
xnor U10978 (N_10978,N_10360,N_10265);
and U10979 (N_10979,N_10146,N_10374);
xnor U10980 (N_10980,N_10311,N_10385);
xnor U10981 (N_10981,N_10141,N_9839);
nand U10982 (N_10982,N_9902,N_9825);
and U10983 (N_10983,N_10313,N_10219);
or U10984 (N_10984,N_10241,N_10435);
and U10985 (N_10985,N_10248,N_10198);
and U10986 (N_10986,N_9894,N_10422);
nor U10987 (N_10987,N_10085,N_10491);
and U10988 (N_10988,N_9752,N_10204);
and U10989 (N_10989,N_10052,N_10038);
or U10990 (N_10990,N_10226,N_10023);
nor U10991 (N_10991,N_10078,N_10104);
and U10992 (N_10992,N_10396,N_10224);
or U10993 (N_10993,N_10082,N_10399);
or U10994 (N_10994,N_10020,N_10174);
and U10995 (N_10995,N_10271,N_9923);
and U10996 (N_10996,N_10368,N_9931);
and U10997 (N_10997,N_10410,N_10108);
and U10998 (N_10998,N_10074,N_9779);
xor U10999 (N_10999,N_10471,N_9903);
xor U11000 (N_11000,N_10297,N_10088);
and U11001 (N_11001,N_10119,N_9849);
nand U11002 (N_11002,N_10474,N_10417);
and U11003 (N_11003,N_10217,N_10367);
xor U11004 (N_11004,N_9903,N_10107);
nand U11005 (N_11005,N_9811,N_10310);
or U11006 (N_11006,N_10415,N_10153);
nand U11007 (N_11007,N_10379,N_9989);
xor U11008 (N_11008,N_10152,N_10066);
nor U11009 (N_11009,N_9977,N_10288);
xor U11010 (N_11010,N_10149,N_10330);
nand U11011 (N_11011,N_10427,N_10487);
xnor U11012 (N_11012,N_10471,N_10040);
nand U11013 (N_11013,N_9771,N_10429);
xor U11014 (N_11014,N_10231,N_10038);
nand U11015 (N_11015,N_10059,N_10056);
nor U11016 (N_11016,N_10151,N_10031);
nand U11017 (N_11017,N_10251,N_10185);
or U11018 (N_11018,N_10236,N_10153);
nand U11019 (N_11019,N_10445,N_10426);
and U11020 (N_11020,N_10461,N_10251);
and U11021 (N_11021,N_10123,N_9796);
xnor U11022 (N_11022,N_9757,N_9893);
nand U11023 (N_11023,N_10126,N_10290);
and U11024 (N_11024,N_10465,N_9994);
nor U11025 (N_11025,N_9921,N_10278);
or U11026 (N_11026,N_10101,N_10179);
and U11027 (N_11027,N_10203,N_10065);
or U11028 (N_11028,N_9841,N_10196);
nand U11029 (N_11029,N_9867,N_10423);
nor U11030 (N_11030,N_9987,N_10307);
nand U11031 (N_11031,N_9944,N_10095);
xor U11032 (N_11032,N_10346,N_9998);
and U11033 (N_11033,N_9867,N_10099);
nor U11034 (N_11034,N_10152,N_10457);
nor U11035 (N_11035,N_10066,N_9869);
xor U11036 (N_11036,N_10326,N_10244);
or U11037 (N_11037,N_10394,N_10334);
and U11038 (N_11038,N_10402,N_9963);
nor U11039 (N_11039,N_10194,N_9954);
or U11040 (N_11040,N_10273,N_10120);
and U11041 (N_11041,N_10022,N_10411);
nor U11042 (N_11042,N_10219,N_9912);
and U11043 (N_11043,N_9898,N_10042);
and U11044 (N_11044,N_9816,N_10147);
or U11045 (N_11045,N_10051,N_10430);
nor U11046 (N_11046,N_10338,N_10303);
nor U11047 (N_11047,N_9782,N_10454);
nand U11048 (N_11048,N_10429,N_10319);
nor U11049 (N_11049,N_10215,N_10376);
xor U11050 (N_11050,N_10109,N_9816);
xor U11051 (N_11051,N_10337,N_9857);
nor U11052 (N_11052,N_10321,N_10053);
nor U11053 (N_11053,N_9866,N_10494);
nand U11054 (N_11054,N_9784,N_10135);
nand U11055 (N_11055,N_10281,N_10073);
and U11056 (N_11056,N_10266,N_10020);
nand U11057 (N_11057,N_10405,N_10023);
nor U11058 (N_11058,N_10428,N_9880);
xor U11059 (N_11059,N_9755,N_10394);
nand U11060 (N_11060,N_10441,N_9877);
nor U11061 (N_11061,N_10411,N_10068);
and U11062 (N_11062,N_10087,N_10244);
or U11063 (N_11063,N_10099,N_9813);
or U11064 (N_11064,N_10097,N_9989);
nand U11065 (N_11065,N_10273,N_9753);
or U11066 (N_11066,N_9904,N_10247);
and U11067 (N_11067,N_10188,N_9891);
and U11068 (N_11068,N_10135,N_10409);
and U11069 (N_11069,N_10120,N_10379);
xor U11070 (N_11070,N_10292,N_10201);
nand U11071 (N_11071,N_10239,N_9998);
or U11072 (N_11072,N_10119,N_10220);
and U11073 (N_11073,N_9931,N_9881);
nand U11074 (N_11074,N_10166,N_10331);
and U11075 (N_11075,N_10416,N_9907);
nand U11076 (N_11076,N_10276,N_10286);
and U11077 (N_11077,N_10237,N_9813);
or U11078 (N_11078,N_10290,N_9804);
or U11079 (N_11079,N_10154,N_9823);
xor U11080 (N_11080,N_10430,N_10429);
or U11081 (N_11081,N_10345,N_10430);
nor U11082 (N_11082,N_10023,N_10242);
nand U11083 (N_11083,N_10384,N_10334);
nand U11084 (N_11084,N_9971,N_9998);
or U11085 (N_11085,N_10069,N_10004);
or U11086 (N_11086,N_10162,N_9848);
or U11087 (N_11087,N_10483,N_9988);
or U11088 (N_11088,N_10046,N_10266);
xor U11089 (N_11089,N_10224,N_10412);
nor U11090 (N_11090,N_9998,N_9988);
or U11091 (N_11091,N_10378,N_10054);
nand U11092 (N_11092,N_10332,N_9848);
xor U11093 (N_11093,N_10036,N_10232);
xnor U11094 (N_11094,N_10446,N_10246);
xnor U11095 (N_11095,N_10005,N_10278);
and U11096 (N_11096,N_10434,N_9983);
or U11097 (N_11097,N_10112,N_10425);
and U11098 (N_11098,N_10286,N_10311);
nand U11099 (N_11099,N_9809,N_9953);
nor U11100 (N_11100,N_10336,N_9831);
or U11101 (N_11101,N_10169,N_10307);
nand U11102 (N_11102,N_10279,N_10207);
xnor U11103 (N_11103,N_10434,N_10008);
and U11104 (N_11104,N_10210,N_10248);
xor U11105 (N_11105,N_10057,N_10211);
nor U11106 (N_11106,N_10372,N_10396);
and U11107 (N_11107,N_9904,N_10292);
nor U11108 (N_11108,N_10152,N_10313);
xnor U11109 (N_11109,N_9973,N_10023);
xnor U11110 (N_11110,N_10417,N_10338);
and U11111 (N_11111,N_10065,N_10136);
xnor U11112 (N_11112,N_10380,N_9751);
and U11113 (N_11113,N_10285,N_10246);
or U11114 (N_11114,N_9894,N_9875);
or U11115 (N_11115,N_10142,N_10407);
nand U11116 (N_11116,N_9854,N_10161);
and U11117 (N_11117,N_10361,N_9992);
xor U11118 (N_11118,N_9898,N_10468);
xor U11119 (N_11119,N_9918,N_10495);
xnor U11120 (N_11120,N_10178,N_10404);
nor U11121 (N_11121,N_10028,N_10097);
nand U11122 (N_11122,N_10492,N_10266);
and U11123 (N_11123,N_10172,N_9851);
nand U11124 (N_11124,N_10229,N_10242);
and U11125 (N_11125,N_10341,N_10191);
xor U11126 (N_11126,N_10429,N_10242);
nand U11127 (N_11127,N_9909,N_10205);
and U11128 (N_11128,N_9987,N_9998);
nand U11129 (N_11129,N_10147,N_10034);
xnor U11130 (N_11130,N_9902,N_10250);
nand U11131 (N_11131,N_10097,N_9971);
xor U11132 (N_11132,N_10114,N_9948);
xor U11133 (N_11133,N_10292,N_10250);
and U11134 (N_11134,N_10402,N_9809);
and U11135 (N_11135,N_10103,N_10235);
nor U11136 (N_11136,N_10063,N_9814);
nand U11137 (N_11137,N_10230,N_10131);
xor U11138 (N_11138,N_10046,N_10443);
nand U11139 (N_11139,N_10363,N_10185);
nor U11140 (N_11140,N_10204,N_9806);
or U11141 (N_11141,N_10083,N_10086);
xor U11142 (N_11142,N_10417,N_10204);
xnor U11143 (N_11143,N_9992,N_9995);
nand U11144 (N_11144,N_10095,N_9996);
xnor U11145 (N_11145,N_10461,N_10382);
nor U11146 (N_11146,N_9834,N_9867);
or U11147 (N_11147,N_9951,N_10366);
or U11148 (N_11148,N_10359,N_10118);
xor U11149 (N_11149,N_9898,N_10253);
or U11150 (N_11150,N_10169,N_10449);
nor U11151 (N_11151,N_9953,N_9886);
nand U11152 (N_11152,N_10339,N_10165);
nor U11153 (N_11153,N_9958,N_10490);
nor U11154 (N_11154,N_9821,N_10161);
xor U11155 (N_11155,N_10363,N_10380);
or U11156 (N_11156,N_9845,N_10126);
and U11157 (N_11157,N_10367,N_9821);
xor U11158 (N_11158,N_9852,N_9775);
and U11159 (N_11159,N_9828,N_9927);
and U11160 (N_11160,N_9920,N_9834);
nand U11161 (N_11161,N_9852,N_9878);
and U11162 (N_11162,N_10036,N_10090);
or U11163 (N_11163,N_10438,N_10365);
or U11164 (N_11164,N_10272,N_10308);
or U11165 (N_11165,N_10122,N_10270);
and U11166 (N_11166,N_9978,N_10102);
and U11167 (N_11167,N_10183,N_10185);
or U11168 (N_11168,N_10335,N_9918);
and U11169 (N_11169,N_10147,N_9991);
and U11170 (N_11170,N_9962,N_10080);
xor U11171 (N_11171,N_10390,N_9803);
nor U11172 (N_11172,N_9769,N_9899);
and U11173 (N_11173,N_10225,N_9792);
nor U11174 (N_11174,N_9837,N_10031);
or U11175 (N_11175,N_10408,N_9871);
nor U11176 (N_11176,N_10436,N_10457);
nand U11177 (N_11177,N_10117,N_10411);
xnor U11178 (N_11178,N_9868,N_10198);
nor U11179 (N_11179,N_10415,N_9918);
nand U11180 (N_11180,N_10024,N_10102);
nor U11181 (N_11181,N_9867,N_10220);
or U11182 (N_11182,N_10251,N_9853);
nand U11183 (N_11183,N_10268,N_9944);
nand U11184 (N_11184,N_9834,N_9752);
and U11185 (N_11185,N_10133,N_10216);
nor U11186 (N_11186,N_9914,N_9761);
xor U11187 (N_11187,N_10132,N_10275);
nand U11188 (N_11188,N_9803,N_9953);
and U11189 (N_11189,N_10272,N_10349);
nand U11190 (N_11190,N_9806,N_10040);
nor U11191 (N_11191,N_10473,N_10171);
nand U11192 (N_11192,N_10484,N_10217);
nand U11193 (N_11193,N_10393,N_10147);
nand U11194 (N_11194,N_10154,N_10221);
xnor U11195 (N_11195,N_10315,N_10372);
xor U11196 (N_11196,N_9854,N_10480);
nor U11197 (N_11197,N_9941,N_9786);
or U11198 (N_11198,N_10154,N_9904);
xnor U11199 (N_11199,N_9828,N_9904);
nor U11200 (N_11200,N_10420,N_10467);
xnor U11201 (N_11201,N_10479,N_9873);
and U11202 (N_11202,N_10232,N_10109);
and U11203 (N_11203,N_10033,N_10221);
or U11204 (N_11204,N_10493,N_10045);
and U11205 (N_11205,N_10136,N_10006);
nor U11206 (N_11206,N_10051,N_10371);
nand U11207 (N_11207,N_9969,N_10302);
or U11208 (N_11208,N_9844,N_10015);
or U11209 (N_11209,N_10388,N_10107);
and U11210 (N_11210,N_9867,N_10189);
and U11211 (N_11211,N_10373,N_10144);
xnor U11212 (N_11212,N_10111,N_9927);
and U11213 (N_11213,N_9824,N_10205);
nor U11214 (N_11214,N_9962,N_10453);
or U11215 (N_11215,N_10341,N_10152);
nand U11216 (N_11216,N_10110,N_9957);
or U11217 (N_11217,N_9987,N_10058);
xnor U11218 (N_11218,N_10085,N_10141);
and U11219 (N_11219,N_9923,N_9899);
xnor U11220 (N_11220,N_10421,N_10077);
nor U11221 (N_11221,N_10272,N_9964);
nand U11222 (N_11222,N_10492,N_10044);
nor U11223 (N_11223,N_9931,N_10167);
or U11224 (N_11224,N_10001,N_10005);
xor U11225 (N_11225,N_9780,N_9986);
nand U11226 (N_11226,N_10194,N_9860);
or U11227 (N_11227,N_10220,N_10404);
nand U11228 (N_11228,N_9984,N_10224);
and U11229 (N_11229,N_9972,N_10219);
nand U11230 (N_11230,N_10222,N_10389);
xnor U11231 (N_11231,N_10216,N_10283);
xor U11232 (N_11232,N_10138,N_9895);
nor U11233 (N_11233,N_9939,N_9849);
xor U11234 (N_11234,N_10043,N_9823);
xor U11235 (N_11235,N_10370,N_10426);
and U11236 (N_11236,N_10199,N_10098);
nand U11237 (N_11237,N_10208,N_10422);
nor U11238 (N_11238,N_10108,N_9954);
xor U11239 (N_11239,N_9846,N_10132);
nand U11240 (N_11240,N_10034,N_10085);
or U11241 (N_11241,N_10277,N_9821);
or U11242 (N_11242,N_10035,N_9938);
xor U11243 (N_11243,N_10487,N_10183);
or U11244 (N_11244,N_10084,N_9967);
and U11245 (N_11245,N_10380,N_10196);
xnor U11246 (N_11246,N_10368,N_10256);
nor U11247 (N_11247,N_10005,N_9802);
xor U11248 (N_11248,N_10077,N_10168);
xor U11249 (N_11249,N_10169,N_10441);
and U11250 (N_11250,N_10500,N_10974);
nor U11251 (N_11251,N_11119,N_11185);
nor U11252 (N_11252,N_11017,N_10621);
nor U11253 (N_11253,N_10809,N_11087);
and U11254 (N_11254,N_10764,N_10912);
nand U11255 (N_11255,N_11216,N_10588);
nand U11256 (N_11256,N_10850,N_10696);
xor U11257 (N_11257,N_11022,N_10849);
nand U11258 (N_11258,N_10608,N_10758);
nor U11259 (N_11259,N_11238,N_11040);
nor U11260 (N_11260,N_10819,N_10547);
nor U11261 (N_11261,N_11133,N_11114);
and U11262 (N_11262,N_11137,N_10582);
or U11263 (N_11263,N_10871,N_10748);
or U11264 (N_11264,N_11019,N_11071);
nand U11265 (N_11265,N_10839,N_11097);
and U11266 (N_11266,N_10675,N_11234);
and U11267 (N_11267,N_10502,N_10680);
nand U11268 (N_11268,N_10613,N_10730);
xnor U11269 (N_11269,N_10833,N_10860);
and U11270 (N_11270,N_11236,N_10935);
nor U11271 (N_11271,N_10847,N_10549);
or U11272 (N_11272,N_11220,N_10720);
nand U11273 (N_11273,N_10798,N_10727);
nand U11274 (N_11274,N_10583,N_10831);
nand U11275 (N_11275,N_10682,N_10728);
or U11276 (N_11276,N_11230,N_11138);
xor U11277 (N_11277,N_10692,N_10618);
and U11278 (N_11278,N_11165,N_10787);
or U11279 (N_11279,N_11224,N_10842);
nor U11280 (N_11280,N_10548,N_10987);
xnor U11281 (N_11281,N_11247,N_10650);
or U11282 (N_11282,N_11136,N_10633);
xnor U11283 (N_11283,N_11110,N_11099);
xor U11284 (N_11284,N_10814,N_11214);
xnor U11285 (N_11285,N_10725,N_11078);
nand U11286 (N_11286,N_10896,N_10864);
nor U11287 (N_11287,N_11228,N_10830);
xnor U11288 (N_11288,N_10963,N_10979);
nor U11289 (N_11289,N_10607,N_10595);
nor U11290 (N_11290,N_10740,N_10687);
and U11291 (N_11291,N_11015,N_11131);
and U11292 (N_11292,N_10881,N_11160);
or U11293 (N_11293,N_10928,N_10718);
nor U11294 (N_11294,N_10895,N_10704);
and U11295 (N_11295,N_10615,N_10592);
nand U11296 (N_11296,N_10572,N_10706);
nand U11297 (N_11297,N_11079,N_11003);
or U11298 (N_11298,N_11073,N_11018);
nor U11299 (N_11299,N_11227,N_11034);
and U11300 (N_11300,N_10771,N_11070);
nand U11301 (N_11301,N_10872,N_10511);
or U11302 (N_11302,N_10918,N_11237);
and U11303 (N_11303,N_10964,N_10628);
nand U11304 (N_11304,N_11170,N_11181);
nor U11305 (N_11305,N_11067,N_10584);
or U11306 (N_11306,N_10795,N_11207);
or U11307 (N_11307,N_10915,N_10899);
nor U11308 (N_11308,N_10719,N_10676);
and U11309 (N_11309,N_10634,N_10707);
or U11310 (N_11310,N_11244,N_10835);
nor U11311 (N_11311,N_10806,N_10744);
nand U11312 (N_11312,N_10879,N_10555);
and U11313 (N_11313,N_10523,N_11225);
nor U11314 (N_11314,N_10762,N_10664);
xnor U11315 (N_11315,N_10878,N_10884);
and U11316 (N_11316,N_11210,N_10916);
nor U11317 (N_11317,N_11024,N_11113);
nand U11318 (N_11318,N_10891,N_10563);
or U11319 (N_11319,N_10865,N_10942);
nand U11320 (N_11320,N_10559,N_10639);
nor U11321 (N_11321,N_11014,N_10914);
and U11322 (N_11322,N_10827,N_10792);
xnor U11323 (N_11323,N_11130,N_10816);
nand U11324 (N_11324,N_10620,N_10554);
or U11325 (N_11325,N_10610,N_10735);
and U11326 (N_11326,N_10980,N_11032);
nor U11327 (N_11327,N_10505,N_11107);
and U11328 (N_11328,N_10829,N_11001);
nand U11329 (N_11329,N_10514,N_11006);
nor U11330 (N_11330,N_10927,N_10856);
nand U11331 (N_11331,N_10825,N_10875);
and U11332 (N_11332,N_10565,N_10560);
xnor U11333 (N_11333,N_11121,N_11103);
nand U11334 (N_11334,N_10750,N_10978);
nor U11335 (N_11335,N_10997,N_10781);
and U11336 (N_11336,N_11086,N_10524);
and U11337 (N_11337,N_10900,N_11027);
and U11338 (N_11338,N_10773,N_10948);
or U11339 (N_11339,N_10738,N_11231);
nand U11340 (N_11340,N_10810,N_11168);
or U11341 (N_11341,N_10855,N_11148);
nand U11342 (N_11342,N_10820,N_10539);
or U11343 (N_11343,N_10874,N_10695);
nand U11344 (N_11344,N_11115,N_11029);
nand U11345 (N_11345,N_10890,N_10690);
or U11346 (N_11346,N_11028,N_10824);
or U11347 (N_11347,N_10826,N_10800);
and U11348 (N_11348,N_10946,N_10724);
or U11349 (N_11349,N_10779,N_10925);
and U11350 (N_11350,N_10991,N_11164);
nand U11351 (N_11351,N_10546,N_10652);
and U11352 (N_11352,N_10603,N_10536);
xnor U11353 (N_11353,N_10667,N_10538);
nor U11354 (N_11354,N_11104,N_10789);
nand U11355 (N_11355,N_10998,N_10671);
nand U11356 (N_11356,N_10705,N_11140);
nor U11357 (N_11357,N_10954,N_11026);
nand U11358 (N_11358,N_11072,N_11056);
nor U11359 (N_11359,N_10767,N_11043);
and U11360 (N_11360,N_10561,N_11010);
and U11361 (N_11361,N_11201,N_11057);
and U11362 (N_11362,N_11112,N_11052);
nand U11363 (N_11363,N_10863,N_11095);
and U11364 (N_11364,N_10892,N_10817);
or U11365 (N_11365,N_10597,N_11157);
or U11366 (N_11366,N_10852,N_10640);
xor U11367 (N_11367,N_10923,N_10861);
nor U11368 (N_11368,N_11124,N_11005);
and U11369 (N_11369,N_10769,N_11223);
nand U11370 (N_11370,N_10845,N_11091);
or U11371 (N_11371,N_11175,N_11037);
nand U11372 (N_11372,N_10805,N_10977);
nor U11373 (N_11373,N_10818,N_11211);
and U11374 (N_11374,N_11127,N_10732);
nand U11375 (N_11375,N_11069,N_11106);
xnor U11376 (N_11376,N_11186,N_11122);
xor U11377 (N_11377,N_10917,N_11085);
and U11378 (N_11378,N_10813,N_10754);
or U11379 (N_11379,N_10905,N_10777);
nand U11380 (N_11380,N_10670,N_10858);
and U11381 (N_11381,N_10622,N_10699);
or U11382 (N_11382,N_10729,N_10908);
and U11383 (N_11383,N_10868,N_10510);
xnor U11384 (N_11384,N_11241,N_10672);
nor U11385 (N_11385,N_10578,N_10938);
nand U11386 (N_11386,N_11066,N_11033);
and U11387 (N_11387,N_10663,N_10958);
nor U11388 (N_11388,N_10883,N_10721);
xnor U11389 (N_11389,N_10602,N_10904);
or U11390 (N_11390,N_10902,N_10649);
nor U11391 (N_11391,N_11209,N_10552);
nor U11392 (N_11392,N_11042,N_11154);
nand U11393 (N_11393,N_11146,N_11174);
nand U11394 (N_11394,N_10635,N_11023);
and U11395 (N_11395,N_10619,N_10623);
xnor U11396 (N_11396,N_11199,N_11150);
xnor U11397 (N_11397,N_10533,N_10641);
nand U11398 (N_11398,N_10960,N_10526);
nand U11399 (N_11399,N_10741,N_10697);
or U11400 (N_11400,N_11200,N_10966);
or U11401 (N_11401,N_11152,N_11187);
or U11402 (N_11402,N_10975,N_11156);
nor U11403 (N_11403,N_11059,N_10823);
and U11404 (N_11404,N_11083,N_11031);
nor U11405 (N_11405,N_11117,N_10776);
or U11406 (N_11406,N_10971,N_11172);
xnor U11407 (N_11407,N_11147,N_10924);
nand U11408 (N_11408,N_10556,N_10678);
or U11409 (N_11409,N_10828,N_10553);
and U11410 (N_11410,N_10605,N_10886);
nand U11411 (N_11411,N_10543,N_11126);
or U11412 (N_11412,N_10586,N_10617);
nor U11413 (N_11413,N_10537,N_10940);
or U11414 (N_11414,N_11162,N_10911);
and U11415 (N_11415,N_10965,N_11149);
nor U11416 (N_11416,N_10677,N_11101);
or U11417 (N_11417,N_10765,N_11055);
or U11418 (N_11418,N_10519,N_10714);
xor U11419 (N_11419,N_10612,N_10688);
xnor U11420 (N_11420,N_10989,N_10585);
nor U11421 (N_11421,N_11222,N_11190);
and U11422 (N_11422,N_10962,N_11044);
and U11423 (N_11423,N_10929,N_10836);
or U11424 (N_11424,N_10518,N_11098);
xor U11425 (N_11425,N_10821,N_11111);
or U11426 (N_11426,N_11158,N_10742);
xnor U11427 (N_11427,N_11249,N_10631);
or U11428 (N_11428,N_10532,N_11173);
xnor U11429 (N_11429,N_11243,N_10711);
or U11430 (N_11430,N_10712,N_10756);
or U11431 (N_11431,N_10848,N_10801);
or U11432 (N_11432,N_10803,N_10772);
or U11433 (N_11433,N_10564,N_10939);
and U11434 (N_11434,N_11060,N_11178);
and U11435 (N_11435,N_10796,N_11206);
or U11436 (N_11436,N_11159,N_10981);
nor U11437 (N_11437,N_11065,N_10604);
and U11438 (N_11438,N_10843,N_10508);
nor U11439 (N_11439,N_10636,N_10791);
nand U11440 (N_11440,N_10530,N_11096);
nor U11441 (N_11441,N_10609,N_10757);
and U11442 (N_11442,N_10644,N_10625);
nor U11443 (N_11443,N_10713,N_10507);
xnor U11444 (N_11444,N_10674,N_10626);
nor U11445 (N_11445,N_10786,N_10804);
nand U11446 (N_11446,N_10734,N_10837);
xnor U11447 (N_11447,N_11198,N_11179);
xnor U11448 (N_11448,N_11193,N_10726);
nand U11449 (N_11449,N_10600,N_11062);
xor U11450 (N_11450,N_10647,N_11232);
or U11451 (N_11451,N_10577,N_11092);
and U11452 (N_11452,N_10957,N_10802);
or U11453 (N_11453,N_11053,N_10658);
nand U11454 (N_11454,N_10956,N_10751);
and U11455 (N_11455,N_11248,N_10793);
xnor U11456 (N_11456,N_10961,N_10783);
nand U11457 (N_11457,N_10766,N_10969);
nand U11458 (N_11458,N_11221,N_11089);
nand U11459 (N_11459,N_10749,N_11049);
and U11460 (N_11460,N_11202,N_10984);
xnor U11461 (N_11461,N_10606,N_10504);
xor U11462 (N_11462,N_10598,N_10542);
and U11463 (N_11463,N_11082,N_10708);
nor U11464 (N_11464,N_11048,N_10601);
xor U11465 (N_11465,N_11000,N_10659);
or U11466 (N_11466,N_11233,N_10943);
nor U11467 (N_11467,N_10573,N_10703);
and U11468 (N_11468,N_10694,N_10521);
xor U11469 (N_11469,N_11176,N_10876);
nand U11470 (N_11470,N_10866,N_10515);
xnor U11471 (N_11471,N_10580,N_10568);
and U11472 (N_11472,N_11189,N_11008);
or U11473 (N_11473,N_11144,N_10574);
or U11474 (N_11474,N_10562,N_11041);
and U11475 (N_11475,N_10934,N_10873);
nor U11476 (N_11476,N_11075,N_10882);
nand U11477 (N_11477,N_10867,N_10550);
nand U11478 (N_11478,N_11125,N_10522);
nor U11479 (N_11479,N_11004,N_10716);
xnor U11480 (N_11480,N_10887,N_11246);
nor U11481 (N_11481,N_10662,N_10541);
or U11482 (N_11482,N_10941,N_10691);
nand U11483 (N_11483,N_10944,N_11108);
nor U11484 (N_11484,N_10576,N_10838);
nor U11485 (N_11485,N_10759,N_10755);
nor U11486 (N_11486,N_10557,N_11074);
or U11487 (N_11487,N_10651,N_11245);
nand U11488 (N_11488,N_10910,N_11134);
xor U11489 (N_11489,N_11182,N_11204);
and U11490 (N_11490,N_10698,N_10527);
or U11491 (N_11491,N_11215,N_10648);
xnor U11492 (N_11492,N_10534,N_10747);
and U11493 (N_11493,N_10993,N_10591);
and U11494 (N_11494,N_10949,N_11128);
xor U11495 (N_11495,N_10587,N_11039);
nor U11496 (N_11496,N_10907,N_11171);
or U11497 (N_11497,N_10513,N_10945);
xnor U11498 (N_11498,N_10893,N_10785);
and U11499 (N_11499,N_10794,N_10669);
nor U11500 (N_11500,N_10637,N_10529);
or U11501 (N_11501,N_10594,N_11007);
and U11502 (N_11502,N_10709,N_10788);
nand U11503 (N_11503,N_10665,N_10947);
or U11504 (N_11504,N_10501,N_11197);
nand U11505 (N_11505,N_10629,N_10857);
nand U11506 (N_11506,N_11123,N_10930);
or U11507 (N_11507,N_10760,N_11013);
or U11508 (N_11508,N_11217,N_10973);
nor U11509 (N_11509,N_11046,N_10683);
nor U11510 (N_11510,N_10937,N_11102);
nand U11511 (N_11511,N_10784,N_10913);
nor U11512 (N_11512,N_10517,N_10976);
nand U11513 (N_11513,N_11239,N_10885);
or U11514 (N_11514,N_10880,N_11021);
xnor U11515 (N_11515,N_10888,N_10516);
xnor U11516 (N_11516,N_10571,N_11132);
nand U11517 (N_11517,N_11045,N_11012);
nand U11518 (N_11518,N_11169,N_11076);
xnor U11519 (N_11519,N_10983,N_10655);
and U11520 (N_11520,N_10717,N_10632);
and U11521 (N_11521,N_10723,N_10822);
nor U11522 (N_11522,N_10614,N_10870);
nor U11523 (N_11523,N_10968,N_11050);
and U11524 (N_11524,N_10710,N_11155);
xnor U11525 (N_11525,N_10684,N_10862);
nor U11526 (N_11526,N_10811,N_11145);
and U11527 (N_11527,N_11167,N_10972);
or U11528 (N_11528,N_10596,N_10763);
and U11529 (N_11529,N_10528,N_10558);
xnor U11530 (N_11530,N_10778,N_11194);
nor U11531 (N_11531,N_10761,N_10745);
and U11532 (N_11532,N_11009,N_10666);
nor U11533 (N_11533,N_10921,N_11077);
and U11534 (N_11534,N_10679,N_10654);
nor U11535 (N_11535,N_10545,N_10689);
nor U11536 (N_11536,N_10731,N_10869);
or U11537 (N_11537,N_10898,N_10599);
and U11538 (N_11538,N_10986,N_11016);
nor U11539 (N_11539,N_11161,N_11177);
nor U11540 (N_11540,N_11143,N_10660);
or U11541 (N_11541,N_10990,N_10753);
nand U11542 (N_11542,N_11002,N_10952);
xnor U11543 (N_11543,N_11038,N_11142);
or U11544 (N_11544,N_10922,N_10780);
and U11545 (N_11545,N_10686,N_10722);
nand U11546 (N_11546,N_10936,N_10733);
and U11547 (N_11547,N_10700,N_10859);
or U11548 (N_11548,N_10544,N_10701);
xnor U11549 (N_11549,N_10645,N_10509);
or U11550 (N_11550,N_10931,N_11035);
or U11551 (N_11551,N_10953,N_10920);
nand U11552 (N_11552,N_11100,N_10877);
and U11553 (N_11553,N_10782,N_11183);
and U11554 (N_11554,N_11061,N_10775);
and U11555 (N_11555,N_10579,N_11020);
xnor U11556 (N_11556,N_10590,N_10630);
and U11557 (N_11557,N_10919,N_10593);
xor U11558 (N_11558,N_11205,N_11229);
xnor U11559 (N_11559,N_11192,N_10569);
or U11560 (N_11560,N_10808,N_10681);
xor U11561 (N_11561,N_10797,N_10959);
nand U11562 (N_11562,N_11105,N_11196);
nor U11563 (N_11563,N_10840,N_10967);
xor U11564 (N_11564,N_10851,N_10616);
xor U11565 (N_11565,N_10985,N_11242);
nor U11566 (N_11566,N_10581,N_10531);
or U11567 (N_11567,N_11191,N_10894);
nand U11568 (N_11568,N_10807,N_11080);
xnor U11569 (N_11569,N_10846,N_10525);
or U11570 (N_11570,N_11203,N_10812);
nor U11571 (N_11571,N_10506,N_11090);
nor U11572 (N_11572,N_10832,N_11081);
and U11573 (N_11573,N_10570,N_10932);
nor U11574 (N_11574,N_11063,N_11240);
nand U11575 (N_11575,N_10853,N_10535);
nor U11576 (N_11576,N_10624,N_11120);
or U11577 (N_11577,N_10512,N_10657);
nor U11578 (N_11578,N_10627,N_11188);
or U11579 (N_11579,N_10567,N_11139);
or U11580 (N_11580,N_10743,N_10889);
or U11581 (N_11581,N_11212,N_10951);
or U11582 (N_11582,N_10673,N_10909);
nor U11583 (N_11583,N_10643,N_11163);
nor U11584 (N_11584,N_10841,N_11068);
xor U11585 (N_11585,N_10992,N_11208);
nor U11586 (N_11586,N_10950,N_11058);
nor U11587 (N_11587,N_11153,N_11088);
and U11588 (N_11588,N_10611,N_10897);
nor U11589 (N_11589,N_10988,N_10768);
and U11590 (N_11590,N_10702,N_10520);
nand U11591 (N_11591,N_10854,N_11213);
and U11592 (N_11592,N_10955,N_10815);
nor U11593 (N_11593,N_11011,N_10994);
or U11594 (N_11594,N_10551,N_11135);
or U11595 (N_11595,N_10903,N_10999);
or U11596 (N_11596,N_10503,N_11226);
nand U11597 (N_11597,N_10996,N_10774);
xnor U11598 (N_11598,N_10737,N_11184);
or U11599 (N_11599,N_10844,N_11166);
nand U11600 (N_11600,N_10566,N_11054);
xnor U11601 (N_11601,N_11118,N_10638);
xnor U11602 (N_11602,N_11093,N_10901);
nor U11603 (N_11603,N_11047,N_11141);
nand U11604 (N_11604,N_10715,N_10790);
and U11605 (N_11605,N_11195,N_11218);
and U11606 (N_11606,N_11151,N_10656);
nor U11607 (N_11607,N_11036,N_10685);
and U11608 (N_11608,N_10739,N_10540);
and U11609 (N_11609,N_10995,N_10736);
nand U11610 (N_11610,N_10668,N_11025);
xnor U11611 (N_11611,N_10589,N_11116);
xnor U11612 (N_11612,N_11235,N_10746);
nor U11613 (N_11613,N_10693,N_10926);
or U11614 (N_11614,N_10834,N_10653);
and U11615 (N_11615,N_10752,N_11129);
and U11616 (N_11616,N_10799,N_11180);
xnor U11617 (N_11617,N_10575,N_11064);
or U11618 (N_11618,N_10970,N_11094);
and U11619 (N_11619,N_11109,N_10982);
nand U11620 (N_11620,N_11030,N_10646);
or U11621 (N_11621,N_10906,N_10661);
and U11622 (N_11622,N_10933,N_10642);
nor U11623 (N_11623,N_11219,N_11051);
nand U11624 (N_11624,N_10770,N_11084);
nand U11625 (N_11625,N_10717,N_11056);
nor U11626 (N_11626,N_10970,N_11144);
and U11627 (N_11627,N_10705,N_10704);
or U11628 (N_11628,N_11058,N_10570);
or U11629 (N_11629,N_10937,N_10507);
xor U11630 (N_11630,N_11075,N_11124);
nand U11631 (N_11631,N_10840,N_11062);
nor U11632 (N_11632,N_10798,N_10739);
nor U11633 (N_11633,N_10786,N_10622);
and U11634 (N_11634,N_11178,N_10521);
nand U11635 (N_11635,N_10649,N_10748);
nand U11636 (N_11636,N_10675,N_10515);
xnor U11637 (N_11637,N_10598,N_10619);
nor U11638 (N_11638,N_11016,N_10764);
or U11639 (N_11639,N_11108,N_10710);
and U11640 (N_11640,N_10616,N_11095);
nand U11641 (N_11641,N_11098,N_10891);
nand U11642 (N_11642,N_11093,N_10893);
nor U11643 (N_11643,N_11061,N_10912);
nor U11644 (N_11644,N_10794,N_10584);
xor U11645 (N_11645,N_10597,N_10610);
or U11646 (N_11646,N_10500,N_10574);
nor U11647 (N_11647,N_10848,N_11211);
nor U11648 (N_11648,N_11205,N_10871);
or U11649 (N_11649,N_11124,N_10532);
nor U11650 (N_11650,N_10590,N_11247);
nor U11651 (N_11651,N_10715,N_10744);
nand U11652 (N_11652,N_10667,N_10844);
nor U11653 (N_11653,N_10924,N_10964);
and U11654 (N_11654,N_11029,N_10660);
nor U11655 (N_11655,N_10953,N_10976);
and U11656 (N_11656,N_10565,N_10820);
nor U11657 (N_11657,N_10847,N_10984);
or U11658 (N_11658,N_10965,N_10654);
or U11659 (N_11659,N_10812,N_10915);
nand U11660 (N_11660,N_10528,N_11221);
nand U11661 (N_11661,N_10757,N_11099);
nor U11662 (N_11662,N_10567,N_10919);
xor U11663 (N_11663,N_10557,N_10558);
and U11664 (N_11664,N_11121,N_10975);
nor U11665 (N_11665,N_11149,N_11226);
nand U11666 (N_11666,N_10993,N_11036);
and U11667 (N_11667,N_10526,N_10764);
nand U11668 (N_11668,N_11017,N_11231);
nor U11669 (N_11669,N_10709,N_10911);
nand U11670 (N_11670,N_10682,N_11227);
or U11671 (N_11671,N_10914,N_10817);
and U11672 (N_11672,N_10601,N_10825);
nand U11673 (N_11673,N_10608,N_10786);
nor U11674 (N_11674,N_11186,N_11229);
and U11675 (N_11675,N_10664,N_10795);
nand U11676 (N_11676,N_10653,N_11122);
and U11677 (N_11677,N_11079,N_10836);
and U11678 (N_11678,N_11248,N_11060);
nand U11679 (N_11679,N_11060,N_10546);
and U11680 (N_11680,N_11068,N_10774);
nand U11681 (N_11681,N_10860,N_10736);
xnor U11682 (N_11682,N_10689,N_11165);
and U11683 (N_11683,N_10758,N_10562);
nand U11684 (N_11684,N_10862,N_11194);
nand U11685 (N_11685,N_11248,N_11101);
nor U11686 (N_11686,N_10501,N_10895);
xor U11687 (N_11687,N_10887,N_11206);
nand U11688 (N_11688,N_10805,N_10660);
nand U11689 (N_11689,N_11189,N_10693);
or U11690 (N_11690,N_10615,N_10714);
and U11691 (N_11691,N_10662,N_10556);
and U11692 (N_11692,N_10736,N_10953);
or U11693 (N_11693,N_10590,N_10563);
nand U11694 (N_11694,N_10596,N_10542);
nor U11695 (N_11695,N_11039,N_11092);
xnor U11696 (N_11696,N_10547,N_11140);
nand U11697 (N_11697,N_10958,N_10881);
nor U11698 (N_11698,N_10966,N_10808);
xor U11699 (N_11699,N_10559,N_11038);
nor U11700 (N_11700,N_10933,N_10982);
or U11701 (N_11701,N_10549,N_11100);
nand U11702 (N_11702,N_10619,N_10671);
xor U11703 (N_11703,N_11030,N_10997);
and U11704 (N_11704,N_11002,N_10891);
and U11705 (N_11705,N_10825,N_10853);
nand U11706 (N_11706,N_10788,N_10994);
and U11707 (N_11707,N_10929,N_11226);
nand U11708 (N_11708,N_10924,N_10759);
nor U11709 (N_11709,N_10762,N_10624);
nand U11710 (N_11710,N_10945,N_10624);
or U11711 (N_11711,N_10914,N_10963);
nor U11712 (N_11712,N_10784,N_10682);
xor U11713 (N_11713,N_10553,N_10810);
and U11714 (N_11714,N_10843,N_11052);
or U11715 (N_11715,N_10557,N_11008);
and U11716 (N_11716,N_10976,N_10679);
nor U11717 (N_11717,N_11143,N_11184);
nor U11718 (N_11718,N_11135,N_10563);
xnor U11719 (N_11719,N_10609,N_11049);
nand U11720 (N_11720,N_10997,N_11024);
or U11721 (N_11721,N_10756,N_10772);
xnor U11722 (N_11722,N_10507,N_11217);
nand U11723 (N_11723,N_11222,N_10579);
nand U11724 (N_11724,N_10724,N_11239);
xor U11725 (N_11725,N_11074,N_10577);
xnor U11726 (N_11726,N_11243,N_11022);
and U11727 (N_11727,N_11096,N_10748);
nand U11728 (N_11728,N_10919,N_11152);
xor U11729 (N_11729,N_10800,N_11137);
xnor U11730 (N_11730,N_10923,N_10933);
and U11731 (N_11731,N_10606,N_10814);
nand U11732 (N_11732,N_10903,N_10786);
xor U11733 (N_11733,N_11053,N_10503);
nor U11734 (N_11734,N_10773,N_10658);
or U11735 (N_11735,N_10836,N_11031);
xnor U11736 (N_11736,N_10930,N_10561);
xor U11737 (N_11737,N_10530,N_11122);
nor U11738 (N_11738,N_11114,N_11247);
and U11739 (N_11739,N_10751,N_10925);
nand U11740 (N_11740,N_11219,N_10561);
or U11741 (N_11741,N_10697,N_10993);
xor U11742 (N_11742,N_10595,N_10688);
or U11743 (N_11743,N_10947,N_10841);
or U11744 (N_11744,N_11002,N_10684);
xor U11745 (N_11745,N_10789,N_10620);
or U11746 (N_11746,N_11164,N_10636);
or U11747 (N_11747,N_11235,N_10967);
nor U11748 (N_11748,N_10872,N_10608);
or U11749 (N_11749,N_11059,N_11053);
or U11750 (N_11750,N_10898,N_10732);
xnor U11751 (N_11751,N_10881,N_10506);
xor U11752 (N_11752,N_11156,N_10795);
and U11753 (N_11753,N_10764,N_11117);
nand U11754 (N_11754,N_11231,N_10762);
nor U11755 (N_11755,N_10747,N_11163);
or U11756 (N_11756,N_10681,N_10719);
nor U11757 (N_11757,N_10775,N_10618);
or U11758 (N_11758,N_10596,N_10753);
or U11759 (N_11759,N_11061,N_10962);
nor U11760 (N_11760,N_10871,N_10540);
nand U11761 (N_11761,N_11039,N_10594);
or U11762 (N_11762,N_10861,N_10583);
nor U11763 (N_11763,N_10736,N_10839);
and U11764 (N_11764,N_10963,N_11004);
and U11765 (N_11765,N_10892,N_10984);
or U11766 (N_11766,N_10510,N_11233);
nand U11767 (N_11767,N_11087,N_10838);
nor U11768 (N_11768,N_10741,N_10648);
or U11769 (N_11769,N_10623,N_10979);
nor U11770 (N_11770,N_11068,N_10546);
nand U11771 (N_11771,N_11075,N_10873);
and U11772 (N_11772,N_10541,N_10798);
nor U11773 (N_11773,N_10851,N_11202);
nor U11774 (N_11774,N_10767,N_11039);
nand U11775 (N_11775,N_11186,N_10753);
and U11776 (N_11776,N_11170,N_10505);
and U11777 (N_11777,N_11097,N_10947);
nor U11778 (N_11778,N_10541,N_10789);
nand U11779 (N_11779,N_11090,N_10738);
or U11780 (N_11780,N_10741,N_10843);
or U11781 (N_11781,N_11207,N_10643);
nand U11782 (N_11782,N_10613,N_11135);
and U11783 (N_11783,N_11249,N_10985);
and U11784 (N_11784,N_10507,N_11228);
xor U11785 (N_11785,N_10994,N_10940);
xor U11786 (N_11786,N_10674,N_11242);
nor U11787 (N_11787,N_10956,N_10516);
nor U11788 (N_11788,N_10705,N_10726);
nor U11789 (N_11789,N_11089,N_11128);
xor U11790 (N_11790,N_11015,N_11079);
nor U11791 (N_11791,N_10695,N_10620);
xor U11792 (N_11792,N_10883,N_11055);
and U11793 (N_11793,N_11194,N_10569);
or U11794 (N_11794,N_11147,N_10545);
or U11795 (N_11795,N_10604,N_11153);
and U11796 (N_11796,N_11046,N_11120);
xnor U11797 (N_11797,N_10999,N_10564);
nor U11798 (N_11798,N_10798,N_10889);
or U11799 (N_11799,N_10872,N_10916);
xnor U11800 (N_11800,N_10969,N_10569);
nand U11801 (N_11801,N_10879,N_11069);
nor U11802 (N_11802,N_10537,N_11178);
nor U11803 (N_11803,N_10930,N_11138);
nand U11804 (N_11804,N_10806,N_11199);
nor U11805 (N_11805,N_10981,N_10644);
xor U11806 (N_11806,N_10511,N_10675);
or U11807 (N_11807,N_10562,N_10785);
or U11808 (N_11808,N_10506,N_10691);
or U11809 (N_11809,N_11245,N_10516);
nor U11810 (N_11810,N_10776,N_10624);
or U11811 (N_11811,N_10693,N_10939);
nor U11812 (N_11812,N_11045,N_10787);
xnor U11813 (N_11813,N_11099,N_11080);
nand U11814 (N_11814,N_11201,N_11095);
or U11815 (N_11815,N_10672,N_10794);
xor U11816 (N_11816,N_11029,N_10608);
xnor U11817 (N_11817,N_10992,N_10907);
and U11818 (N_11818,N_10819,N_10972);
xnor U11819 (N_11819,N_11089,N_11028);
and U11820 (N_11820,N_11212,N_11034);
nand U11821 (N_11821,N_10593,N_10508);
and U11822 (N_11822,N_11215,N_11110);
nand U11823 (N_11823,N_10540,N_11017);
nor U11824 (N_11824,N_10866,N_10897);
nand U11825 (N_11825,N_10793,N_10876);
nand U11826 (N_11826,N_10899,N_10640);
nor U11827 (N_11827,N_11044,N_11174);
nand U11828 (N_11828,N_10946,N_10592);
xor U11829 (N_11829,N_10858,N_10925);
xnor U11830 (N_11830,N_11149,N_10881);
nand U11831 (N_11831,N_10937,N_10649);
nor U11832 (N_11832,N_10566,N_11120);
and U11833 (N_11833,N_10689,N_10702);
or U11834 (N_11834,N_10665,N_11079);
nor U11835 (N_11835,N_11090,N_10790);
nor U11836 (N_11836,N_10509,N_10527);
nor U11837 (N_11837,N_10675,N_10713);
nand U11838 (N_11838,N_10862,N_10705);
xor U11839 (N_11839,N_11118,N_11078);
and U11840 (N_11840,N_10882,N_10937);
nor U11841 (N_11841,N_11188,N_11119);
and U11842 (N_11842,N_10630,N_10608);
nand U11843 (N_11843,N_10572,N_10755);
nor U11844 (N_11844,N_11174,N_10509);
nor U11845 (N_11845,N_10579,N_11121);
nor U11846 (N_11846,N_11183,N_11104);
nor U11847 (N_11847,N_10744,N_11002);
and U11848 (N_11848,N_10878,N_10752);
or U11849 (N_11849,N_10668,N_10853);
xnor U11850 (N_11850,N_10517,N_10732);
xnor U11851 (N_11851,N_10585,N_11171);
xor U11852 (N_11852,N_10992,N_10948);
or U11853 (N_11853,N_10783,N_11050);
and U11854 (N_11854,N_10836,N_10977);
nand U11855 (N_11855,N_11107,N_10949);
nand U11856 (N_11856,N_11083,N_11229);
and U11857 (N_11857,N_11051,N_10784);
nor U11858 (N_11858,N_11076,N_11068);
or U11859 (N_11859,N_10919,N_11033);
xor U11860 (N_11860,N_10757,N_11168);
xnor U11861 (N_11861,N_10580,N_10920);
nand U11862 (N_11862,N_10971,N_10641);
nor U11863 (N_11863,N_10982,N_11073);
or U11864 (N_11864,N_11209,N_11034);
and U11865 (N_11865,N_10658,N_10768);
nor U11866 (N_11866,N_10960,N_10604);
nand U11867 (N_11867,N_10789,N_10937);
and U11868 (N_11868,N_10882,N_10974);
and U11869 (N_11869,N_11178,N_10753);
nor U11870 (N_11870,N_10807,N_11032);
or U11871 (N_11871,N_11000,N_11159);
xor U11872 (N_11872,N_10790,N_10545);
nand U11873 (N_11873,N_11006,N_11225);
xor U11874 (N_11874,N_10963,N_10739);
and U11875 (N_11875,N_10614,N_10779);
or U11876 (N_11876,N_10807,N_10737);
nor U11877 (N_11877,N_10614,N_11214);
or U11878 (N_11878,N_11209,N_10670);
nor U11879 (N_11879,N_11184,N_10828);
xor U11880 (N_11880,N_10859,N_11007);
or U11881 (N_11881,N_10648,N_10582);
xor U11882 (N_11882,N_10543,N_10619);
xor U11883 (N_11883,N_10878,N_11121);
and U11884 (N_11884,N_10756,N_11144);
or U11885 (N_11885,N_10939,N_11103);
nand U11886 (N_11886,N_11136,N_10724);
or U11887 (N_11887,N_10679,N_10557);
or U11888 (N_11888,N_10854,N_11169);
xnor U11889 (N_11889,N_10760,N_10662);
nor U11890 (N_11890,N_10788,N_11132);
xnor U11891 (N_11891,N_10807,N_10931);
and U11892 (N_11892,N_10978,N_10983);
or U11893 (N_11893,N_11202,N_11007);
or U11894 (N_11894,N_10808,N_11125);
nand U11895 (N_11895,N_10789,N_11122);
or U11896 (N_11896,N_10981,N_11231);
nor U11897 (N_11897,N_11014,N_10562);
and U11898 (N_11898,N_10720,N_10824);
nor U11899 (N_11899,N_10661,N_10653);
nor U11900 (N_11900,N_11125,N_10826);
xor U11901 (N_11901,N_10561,N_10898);
and U11902 (N_11902,N_10817,N_11000);
nand U11903 (N_11903,N_10729,N_10626);
or U11904 (N_11904,N_11219,N_11188);
nand U11905 (N_11905,N_10676,N_11015);
and U11906 (N_11906,N_10854,N_10652);
xor U11907 (N_11907,N_10930,N_10716);
nand U11908 (N_11908,N_10618,N_11128);
nor U11909 (N_11909,N_10818,N_10647);
or U11910 (N_11910,N_10817,N_10580);
nand U11911 (N_11911,N_10541,N_10871);
and U11912 (N_11912,N_11008,N_10933);
nand U11913 (N_11913,N_10890,N_11037);
nand U11914 (N_11914,N_11192,N_10974);
xnor U11915 (N_11915,N_10772,N_11228);
nand U11916 (N_11916,N_10728,N_10667);
nor U11917 (N_11917,N_11109,N_10898);
and U11918 (N_11918,N_11188,N_11090);
nand U11919 (N_11919,N_10894,N_10721);
nor U11920 (N_11920,N_10980,N_10792);
or U11921 (N_11921,N_10746,N_10849);
nand U11922 (N_11922,N_10946,N_10824);
nor U11923 (N_11923,N_10815,N_10685);
or U11924 (N_11924,N_11216,N_10897);
nand U11925 (N_11925,N_10756,N_10608);
xnor U11926 (N_11926,N_11214,N_10964);
and U11927 (N_11927,N_10940,N_10645);
or U11928 (N_11928,N_10992,N_10822);
xor U11929 (N_11929,N_10928,N_11019);
xor U11930 (N_11930,N_11236,N_10634);
nand U11931 (N_11931,N_10836,N_10589);
xnor U11932 (N_11932,N_10692,N_10771);
nor U11933 (N_11933,N_10579,N_10615);
xnor U11934 (N_11934,N_10808,N_11133);
nor U11935 (N_11935,N_11134,N_10835);
nand U11936 (N_11936,N_10616,N_10885);
or U11937 (N_11937,N_10635,N_11088);
xor U11938 (N_11938,N_10908,N_10535);
nor U11939 (N_11939,N_11247,N_11063);
nand U11940 (N_11940,N_10977,N_10681);
and U11941 (N_11941,N_10566,N_10861);
nand U11942 (N_11942,N_10703,N_11148);
or U11943 (N_11943,N_10884,N_10628);
nand U11944 (N_11944,N_11134,N_11025);
nand U11945 (N_11945,N_11134,N_10920);
nand U11946 (N_11946,N_10671,N_11083);
xor U11947 (N_11947,N_10589,N_10530);
or U11948 (N_11948,N_11029,N_10766);
or U11949 (N_11949,N_10776,N_11190);
xor U11950 (N_11950,N_11237,N_10661);
and U11951 (N_11951,N_10893,N_10534);
xor U11952 (N_11952,N_11050,N_11248);
and U11953 (N_11953,N_10899,N_11200);
nand U11954 (N_11954,N_10826,N_11178);
or U11955 (N_11955,N_10932,N_10658);
or U11956 (N_11956,N_10859,N_10796);
nand U11957 (N_11957,N_11165,N_10790);
nor U11958 (N_11958,N_10724,N_10803);
nand U11959 (N_11959,N_11205,N_10624);
nor U11960 (N_11960,N_10898,N_11134);
and U11961 (N_11961,N_10940,N_10815);
or U11962 (N_11962,N_10864,N_10581);
or U11963 (N_11963,N_11166,N_10504);
nor U11964 (N_11964,N_11193,N_10908);
xor U11965 (N_11965,N_10990,N_10786);
xor U11966 (N_11966,N_10633,N_10732);
nand U11967 (N_11967,N_10797,N_10721);
nor U11968 (N_11968,N_10971,N_10714);
nor U11969 (N_11969,N_11077,N_10947);
nand U11970 (N_11970,N_10648,N_10934);
nand U11971 (N_11971,N_10831,N_10672);
nor U11972 (N_11972,N_10987,N_10645);
nand U11973 (N_11973,N_10795,N_10923);
xnor U11974 (N_11974,N_11198,N_10986);
or U11975 (N_11975,N_11136,N_10688);
xnor U11976 (N_11976,N_11229,N_10532);
nor U11977 (N_11977,N_11247,N_10944);
or U11978 (N_11978,N_11099,N_11200);
or U11979 (N_11979,N_10849,N_10540);
and U11980 (N_11980,N_10754,N_10805);
xor U11981 (N_11981,N_10745,N_10684);
nor U11982 (N_11982,N_10569,N_10845);
and U11983 (N_11983,N_10690,N_11179);
nand U11984 (N_11984,N_10802,N_10690);
or U11985 (N_11985,N_10908,N_10603);
nand U11986 (N_11986,N_10769,N_10658);
and U11987 (N_11987,N_11150,N_10707);
xnor U11988 (N_11988,N_10854,N_10722);
nand U11989 (N_11989,N_10541,N_10673);
nand U11990 (N_11990,N_10822,N_10827);
nand U11991 (N_11991,N_11204,N_11219);
xnor U11992 (N_11992,N_10965,N_10608);
nand U11993 (N_11993,N_10504,N_10796);
nand U11994 (N_11994,N_10805,N_11114);
nand U11995 (N_11995,N_10899,N_10989);
xnor U11996 (N_11996,N_10614,N_11089);
or U11997 (N_11997,N_10886,N_10814);
nand U11998 (N_11998,N_11189,N_10813);
nor U11999 (N_11999,N_10585,N_11097);
or U12000 (N_12000,N_11665,N_11624);
nor U12001 (N_12001,N_11931,N_11304);
and U12002 (N_12002,N_11942,N_11656);
nand U12003 (N_12003,N_11367,N_11677);
or U12004 (N_12004,N_11684,N_11464);
nor U12005 (N_12005,N_11643,N_11469);
or U12006 (N_12006,N_11660,N_11833);
xnor U12007 (N_12007,N_11793,N_11352);
or U12008 (N_12008,N_11622,N_11542);
nor U12009 (N_12009,N_11824,N_11891);
or U12010 (N_12010,N_11341,N_11477);
nand U12011 (N_12011,N_11313,N_11435);
xor U12012 (N_12012,N_11338,N_11438);
or U12013 (N_12013,N_11798,N_11609);
nor U12014 (N_12014,N_11727,N_11849);
xnor U12015 (N_12015,N_11443,N_11962);
and U12016 (N_12016,N_11810,N_11707);
or U12017 (N_12017,N_11493,N_11776);
and U12018 (N_12018,N_11799,N_11552);
nor U12019 (N_12019,N_11281,N_11723);
xnor U12020 (N_12020,N_11548,N_11441);
nand U12021 (N_12021,N_11759,N_11844);
nor U12022 (N_12022,N_11641,N_11371);
or U12023 (N_12023,N_11610,N_11662);
nor U12024 (N_12024,N_11750,N_11454);
or U12025 (N_12025,N_11835,N_11358);
and U12026 (N_12026,N_11733,N_11451);
nand U12027 (N_12027,N_11393,N_11604);
nand U12028 (N_12028,N_11452,N_11459);
xor U12029 (N_12029,N_11502,N_11461);
nor U12030 (N_12030,N_11586,N_11331);
nand U12031 (N_12031,N_11456,N_11715);
xor U12032 (N_12032,N_11334,N_11601);
or U12033 (N_12033,N_11813,N_11420);
and U12034 (N_12034,N_11259,N_11975);
nand U12035 (N_12035,N_11644,N_11611);
nor U12036 (N_12036,N_11623,N_11859);
xor U12037 (N_12037,N_11433,N_11721);
xor U12038 (N_12038,N_11335,N_11319);
or U12039 (N_12039,N_11717,N_11979);
xor U12040 (N_12040,N_11589,N_11786);
or U12041 (N_12041,N_11299,N_11503);
nand U12042 (N_12042,N_11689,N_11893);
and U12043 (N_12043,N_11928,N_11366);
xor U12044 (N_12044,N_11995,N_11694);
or U12045 (N_12045,N_11364,N_11935);
xnor U12046 (N_12046,N_11588,N_11817);
or U12047 (N_12047,N_11445,N_11587);
nor U12048 (N_12048,N_11582,N_11905);
or U12049 (N_12049,N_11574,N_11908);
and U12050 (N_12050,N_11386,N_11402);
or U12051 (N_12051,N_11379,N_11323);
or U12052 (N_12052,N_11682,N_11470);
xor U12053 (N_12053,N_11255,N_11939);
nand U12054 (N_12054,N_11360,N_11567);
nand U12055 (N_12055,N_11388,N_11541);
nor U12056 (N_12056,N_11779,N_11834);
or U12057 (N_12057,N_11520,N_11639);
nor U12058 (N_12058,N_11573,N_11632);
xor U12059 (N_12059,N_11855,N_11982);
xnor U12060 (N_12060,N_11326,N_11288);
nor U12061 (N_12061,N_11809,N_11581);
and U12062 (N_12062,N_11620,N_11322);
and U12063 (N_12063,N_11400,N_11612);
nor U12064 (N_12064,N_11349,N_11501);
nor U12065 (N_12065,N_11256,N_11564);
and U12066 (N_12066,N_11683,N_11792);
xnor U12067 (N_12067,N_11621,N_11351);
nor U12068 (N_12068,N_11330,N_11828);
nor U12069 (N_12069,N_11712,N_11411);
or U12070 (N_12070,N_11932,N_11987);
xor U12071 (N_12071,N_11709,N_11312);
nor U12072 (N_12072,N_11457,N_11812);
and U12073 (N_12073,N_11640,N_11679);
and U12074 (N_12074,N_11480,N_11743);
or U12075 (N_12075,N_11412,N_11897);
nor U12076 (N_12076,N_11851,N_11636);
and U12077 (N_12077,N_11602,N_11909);
nor U12078 (N_12078,N_11568,N_11549);
and U12079 (N_12079,N_11430,N_11691);
nand U12080 (N_12080,N_11698,N_11442);
and U12081 (N_12081,N_11847,N_11376);
xnor U12082 (N_12082,N_11951,N_11695);
and U12083 (N_12083,N_11910,N_11261);
or U12084 (N_12084,N_11446,N_11283);
nand U12085 (N_12085,N_11332,N_11972);
or U12086 (N_12086,N_11466,N_11497);
nand U12087 (N_12087,N_11463,N_11956);
xor U12088 (N_12088,N_11681,N_11667);
xor U12089 (N_12089,N_11362,N_11553);
nand U12090 (N_12090,N_11565,N_11292);
xor U12091 (N_12091,N_11773,N_11751);
or U12092 (N_12092,N_11781,N_11678);
and U12093 (N_12093,N_11607,N_11954);
or U12094 (N_12094,N_11543,N_11378);
xnor U12095 (N_12095,N_11518,N_11722);
and U12096 (N_12096,N_11790,N_11895);
and U12097 (N_12097,N_11274,N_11713);
or U12098 (N_12098,N_11558,N_11576);
or U12099 (N_12099,N_11846,N_11980);
and U12100 (N_12100,N_11287,N_11339);
nand U12101 (N_12101,N_11468,N_11890);
or U12102 (N_12102,N_11926,N_11737);
nand U12103 (N_12103,N_11585,N_11372);
nor U12104 (N_12104,N_11989,N_11422);
and U12105 (N_12105,N_11762,N_11566);
xor U12106 (N_12106,N_11509,N_11746);
and U12107 (N_12107,N_11559,N_11324);
nand U12108 (N_12108,N_11788,N_11535);
nor U12109 (N_12109,N_11580,N_11266);
nand U12110 (N_12110,N_11860,N_11447);
and U12111 (N_12111,N_11342,N_11986);
and U12112 (N_12112,N_11250,N_11419);
xnor U12113 (N_12113,N_11439,N_11265);
nor U12114 (N_12114,N_11894,N_11489);
nand U12115 (N_12115,N_11853,N_11827);
nor U12116 (N_12116,N_11595,N_11763);
nor U12117 (N_12117,N_11770,N_11384);
or U12118 (N_12118,N_11596,N_11729);
or U12119 (N_12119,N_11654,N_11383);
nor U12120 (N_12120,N_11804,N_11510);
xor U12121 (N_12121,N_11831,N_11485);
nand U12122 (N_12122,N_11760,N_11768);
nand U12123 (N_12123,N_11949,N_11732);
and U12124 (N_12124,N_11742,N_11373);
or U12125 (N_12125,N_11301,N_11767);
and U12126 (N_12126,N_11747,N_11839);
nor U12127 (N_12127,N_11592,N_11772);
and U12128 (N_12128,N_11655,N_11803);
or U12129 (N_12129,N_11391,N_11785);
nand U12130 (N_12130,N_11782,N_11883);
and U12131 (N_12131,N_11608,N_11830);
xor U12132 (N_12132,N_11865,N_11325);
nand U12133 (N_12133,N_11857,N_11481);
xnor U12134 (N_12134,N_11886,N_11448);
or U12135 (N_12135,N_11739,N_11514);
xor U12136 (N_12136,N_11885,N_11688);
or U12137 (N_12137,N_11755,N_11692);
xor U12138 (N_12138,N_11554,N_11561);
xnor U12139 (N_12139,N_11506,N_11523);
and U12140 (N_12140,N_11504,N_11437);
nand U12141 (N_12141,N_11850,N_11825);
and U12142 (N_12142,N_11328,N_11368);
nor U12143 (N_12143,N_11981,N_11431);
and U12144 (N_12144,N_11529,N_11795);
nand U12145 (N_12145,N_11693,N_11780);
and U12146 (N_12146,N_11416,N_11344);
nor U12147 (N_12147,N_11436,N_11944);
nand U12148 (N_12148,N_11873,N_11471);
nand U12149 (N_12149,N_11512,N_11591);
and U12150 (N_12150,N_11871,N_11498);
xor U12151 (N_12151,N_11474,N_11957);
nor U12152 (N_12152,N_11359,N_11794);
nor U12153 (N_12153,N_11560,N_11872);
nor U12154 (N_12154,N_11634,N_11590);
nand U12155 (N_12155,N_11937,N_11700);
xnor U12156 (N_12156,N_11413,N_11973);
nand U12157 (N_12157,N_11526,N_11630);
xnor U12158 (N_12158,N_11519,N_11365);
and U12159 (N_12159,N_11736,N_11960);
and U12160 (N_12160,N_11818,N_11916);
nand U12161 (N_12161,N_11947,N_11347);
xnor U12162 (N_12162,N_11361,N_11686);
nand U12163 (N_12163,N_11740,N_11966);
nor U12164 (N_12164,N_11569,N_11533);
nor U12165 (N_12165,N_11728,N_11866);
nand U12166 (N_12166,N_11346,N_11613);
nor U12167 (N_12167,N_11718,N_11598);
nor U12168 (N_12168,N_11556,N_11867);
and U12169 (N_12169,N_11575,N_11414);
nor U12170 (N_12170,N_11906,N_11670);
xnor U12171 (N_12171,N_11531,N_11614);
xnor U12172 (N_12172,N_11653,N_11583);
nor U12173 (N_12173,N_11912,N_11923);
nand U12174 (N_12174,N_11748,N_11964);
xnor U12175 (N_12175,N_11842,N_11726);
nand U12176 (N_12176,N_11837,N_11486);
and U12177 (N_12177,N_11492,N_11298);
and U12178 (N_12178,N_11625,N_11303);
xnor U12179 (N_12179,N_11756,N_11778);
nor U12180 (N_12180,N_11952,N_11711);
and U12181 (N_12181,N_11637,N_11253);
xor U12182 (N_12182,N_11530,N_11652);
and U12183 (N_12183,N_11968,N_11924);
nand U12184 (N_12184,N_11690,N_11421);
and U12185 (N_12185,N_11638,N_11826);
nand U12186 (N_12186,N_11532,N_11955);
xnor U12187 (N_12187,N_11998,N_11343);
nand U12188 (N_12188,N_11807,N_11337);
nor U12189 (N_12189,N_11271,N_11647);
and U12190 (N_12190,N_11467,N_11275);
nand U12191 (N_12191,N_11348,N_11888);
nand U12192 (N_12192,N_11482,N_11946);
and U12193 (N_12193,N_11902,N_11270);
nor U12194 (N_12194,N_11434,N_11615);
xnor U12195 (N_12195,N_11852,N_11879);
and U12196 (N_12196,N_11950,N_11725);
xnor U12197 (N_12197,N_11970,N_11808);
or U12198 (N_12198,N_11544,N_11426);
nand U12199 (N_12199,N_11599,N_11407);
and U12200 (N_12200,N_11864,N_11996);
or U12201 (N_12201,N_11450,N_11490);
or U12202 (N_12202,N_11741,N_11516);
nand U12203 (N_12203,N_11706,N_11405);
xor U12204 (N_12204,N_11282,N_11293);
nor U12205 (N_12205,N_11505,N_11524);
and U12206 (N_12206,N_11843,N_11878);
nor U12207 (N_12207,N_11563,N_11577);
or U12208 (N_12208,N_11633,N_11269);
and U12209 (N_12209,N_11537,N_11976);
or U12210 (N_12210,N_11821,N_11983);
nor U12211 (N_12211,N_11738,N_11994);
and U12212 (N_12212,N_11649,N_11258);
xor U12213 (N_12213,N_11992,N_11687);
xnor U12214 (N_12214,N_11917,N_11385);
or U12215 (N_12215,N_11491,N_11432);
or U12216 (N_12216,N_11765,N_11820);
and U12217 (N_12217,N_11455,N_11401);
nand U12218 (N_12218,N_11494,N_11495);
nand U12219 (N_12219,N_11473,N_11317);
xnor U12220 (N_12220,N_11648,N_11295);
nand U12221 (N_12221,N_11953,N_11327);
nand U12222 (N_12222,N_11761,N_11941);
or U12223 (N_12223,N_11404,N_11657);
nor U12224 (N_12224,N_11701,N_11676);
or U12225 (N_12225,N_11929,N_11398);
xor U12226 (N_12226,N_11919,N_11369);
and U12227 (N_12227,N_11836,N_11719);
nand U12228 (N_12228,N_11579,N_11316);
nand U12229 (N_12229,N_11540,N_11936);
or U12230 (N_12230,N_11899,N_11380);
and U12231 (N_12231,N_11527,N_11300);
xor U12232 (N_12232,N_11796,N_11965);
xnor U12233 (N_12233,N_11744,N_11771);
xor U12234 (N_12234,N_11854,N_11922);
and U12235 (N_12235,N_11285,N_11720);
xnor U12236 (N_12236,N_11315,N_11584);
nor U12237 (N_12237,N_11546,N_11410);
xor U12238 (N_12238,N_11555,N_11479);
and U12239 (N_12239,N_11472,N_11444);
nand U12240 (N_12240,N_11605,N_11958);
or U12241 (N_12241,N_11777,N_11882);
or U12242 (N_12242,N_11704,N_11967);
or U12243 (N_12243,N_11749,N_11805);
and U12244 (N_12244,N_11507,N_11600);
or U12245 (N_12245,N_11874,N_11353);
and U12246 (N_12246,N_11458,N_11307);
xor U12247 (N_12247,N_11626,N_11832);
nand U12248 (N_12248,N_11517,N_11267);
xnor U12249 (N_12249,N_11862,N_11714);
and U12250 (N_12250,N_11496,N_11508);
or U12251 (N_12251,N_11815,N_11791);
xnor U12252 (N_12252,N_11664,N_11534);
nor U12253 (N_12253,N_11515,N_11789);
or U12254 (N_12254,N_11783,N_11408);
nor U12255 (N_12255,N_11417,N_11903);
nand U12256 (N_12256,N_11429,N_11696);
and U12257 (N_12257,N_11674,N_11397);
xor U12258 (N_12258,N_11889,N_11900);
nand U12259 (N_12259,N_11863,N_11550);
and U12260 (N_12260,N_11990,N_11884);
or U12261 (N_12261,N_11356,N_11774);
and U12262 (N_12262,N_11276,N_11845);
or U12263 (N_12263,N_11381,N_11666);
and U12264 (N_12264,N_11672,N_11395);
nand U12265 (N_12265,N_11310,N_11449);
nand U12266 (N_12266,N_11877,N_11263);
xor U12267 (N_12267,N_11974,N_11675);
or U12268 (N_12268,N_11658,N_11930);
or U12269 (N_12269,N_11753,N_11333);
and U12270 (N_12270,N_11671,N_11345);
or U12271 (N_12271,N_11279,N_11428);
nand U12272 (N_12272,N_11856,N_11940);
xnor U12273 (N_12273,N_11769,N_11716);
nor U12274 (N_12274,N_11784,N_11943);
nor U12275 (N_12275,N_11921,N_11927);
xnor U12276 (N_12276,N_11374,N_11984);
nand U12277 (N_12277,N_11881,N_11651);
nor U12278 (N_12278,N_11961,N_11802);
or U12279 (N_12279,N_11308,N_11702);
or U12280 (N_12280,N_11619,N_11819);
or U12281 (N_12281,N_11354,N_11387);
xor U12282 (N_12282,N_11571,N_11465);
or U12283 (N_12283,N_11286,N_11336);
nor U12284 (N_12284,N_11475,N_11500);
xnor U12285 (N_12285,N_11617,N_11396);
or U12286 (N_12286,N_11499,N_11389);
xor U12287 (N_12287,N_11991,N_11306);
nand U12288 (N_12288,N_11551,N_11284);
nand U12289 (N_12289,N_11264,N_11969);
xnor U12290 (N_12290,N_11277,N_11309);
or U12291 (N_12291,N_11616,N_11294);
nand U12292 (N_12292,N_11415,N_11999);
nor U12293 (N_12293,N_11731,N_11280);
xnor U12294 (N_12294,N_11476,N_11948);
nor U12295 (N_12295,N_11659,N_11668);
or U12296 (N_12296,N_11370,N_11513);
xnor U12297 (N_12297,N_11823,N_11735);
and U12298 (N_12298,N_11511,N_11822);
nand U12299 (N_12299,N_11829,N_11650);
and U12300 (N_12300,N_11997,N_11764);
xor U12301 (N_12301,N_11816,N_11363);
and U12302 (N_12302,N_11959,N_11904);
nand U12303 (N_12303,N_11594,N_11403);
nor U12304 (N_12304,N_11705,N_11673);
nand U12305 (N_12305,N_11766,N_11278);
and U12306 (N_12306,N_11730,N_11484);
and U12307 (N_12307,N_11382,N_11314);
and U12308 (N_12308,N_11806,N_11800);
nor U12309 (N_12309,N_11557,N_11710);
nand U12310 (N_12310,N_11251,N_11289);
or U12311 (N_12311,N_11635,N_11978);
nand U12312 (N_12312,N_11272,N_11869);
xnor U12313 (N_12313,N_11907,N_11409);
and U12314 (N_12314,N_11562,N_11290);
nor U12315 (N_12315,N_11318,N_11911);
and U12316 (N_12316,N_11925,N_11811);
nor U12317 (N_12317,N_11302,N_11724);
or U12318 (N_12318,N_11801,N_11977);
and U12319 (N_12319,N_11787,N_11525);
xnor U12320 (N_12320,N_11685,N_11971);
nor U12321 (N_12321,N_11320,N_11870);
xor U12322 (N_12322,N_11483,N_11661);
xnor U12323 (N_12323,N_11528,N_11861);
or U12324 (N_12324,N_11392,N_11311);
xor U12325 (N_12325,N_11868,N_11642);
nor U12326 (N_12326,N_11752,N_11262);
or U12327 (N_12327,N_11321,N_11521);
nor U12328 (N_12328,N_11896,N_11252);
xor U12329 (N_12329,N_11291,N_11775);
nand U12330 (N_12330,N_11570,N_11572);
xor U12331 (N_12331,N_11918,N_11377);
or U12332 (N_12332,N_11993,N_11478);
nor U12333 (N_12333,N_11629,N_11669);
xnor U12334 (N_12334,N_11933,N_11260);
and U12335 (N_12335,N_11536,N_11522);
and U12336 (N_12336,N_11758,N_11938);
or U12337 (N_12337,N_11838,N_11547);
nor U12338 (N_12338,N_11757,N_11627);
nand U12339 (N_12339,N_11915,N_11296);
or U12340 (N_12340,N_11754,N_11708);
nor U12341 (N_12341,N_11423,N_11394);
nor U12342 (N_12342,N_11988,N_11539);
xnor U12343 (N_12343,N_11603,N_11538);
nor U12344 (N_12344,N_11985,N_11273);
nor U12345 (N_12345,N_11390,N_11418);
or U12346 (N_12346,N_11257,N_11887);
and U12347 (N_12347,N_11578,N_11399);
nand U12348 (N_12348,N_11628,N_11329);
nand U12349 (N_12349,N_11680,N_11697);
and U12350 (N_12350,N_11357,N_11424);
and U12351 (N_12351,N_11898,N_11945);
and U12352 (N_12352,N_11453,N_11268);
xor U12353 (N_12353,N_11462,N_11914);
xor U12354 (N_12354,N_11963,N_11875);
nor U12355 (N_12355,N_11848,N_11920);
and U12356 (N_12356,N_11858,N_11841);
nand U12357 (N_12357,N_11460,N_11814);
or U12358 (N_12358,N_11876,N_11425);
or U12359 (N_12359,N_11297,N_11340);
nor U12360 (N_12360,N_11375,N_11254);
or U12361 (N_12361,N_11593,N_11645);
xor U12362 (N_12362,N_11597,N_11797);
or U12363 (N_12363,N_11440,N_11663);
and U12364 (N_12364,N_11901,N_11703);
or U12365 (N_12365,N_11618,N_11545);
nand U12366 (N_12366,N_11406,N_11892);
and U12367 (N_12367,N_11350,N_11913);
xnor U12368 (N_12368,N_11487,N_11880);
or U12369 (N_12369,N_11488,N_11745);
xnor U12370 (N_12370,N_11646,N_11840);
and U12371 (N_12371,N_11734,N_11427);
nor U12372 (N_12372,N_11606,N_11699);
nor U12373 (N_12373,N_11305,N_11355);
nor U12374 (N_12374,N_11934,N_11631);
and U12375 (N_12375,N_11375,N_11291);
xor U12376 (N_12376,N_11774,N_11826);
nor U12377 (N_12377,N_11468,N_11396);
or U12378 (N_12378,N_11417,N_11716);
nand U12379 (N_12379,N_11426,N_11826);
or U12380 (N_12380,N_11637,N_11491);
nand U12381 (N_12381,N_11340,N_11626);
nor U12382 (N_12382,N_11953,N_11363);
nand U12383 (N_12383,N_11281,N_11340);
xnor U12384 (N_12384,N_11894,N_11258);
nor U12385 (N_12385,N_11785,N_11412);
and U12386 (N_12386,N_11387,N_11961);
or U12387 (N_12387,N_11568,N_11435);
xor U12388 (N_12388,N_11562,N_11687);
nand U12389 (N_12389,N_11635,N_11453);
nand U12390 (N_12390,N_11705,N_11919);
xor U12391 (N_12391,N_11603,N_11518);
xor U12392 (N_12392,N_11795,N_11655);
and U12393 (N_12393,N_11674,N_11809);
and U12394 (N_12394,N_11499,N_11825);
and U12395 (N_12395,N_11736,N_11306);
nor U12396 (N_12396,N_11563,N_11990);
or U12397 (N_12397,N_11470,N_11573);
and U12398 (N_12398,N_11842,N_11839);
xor U12399 (N_12399,N_11373,N_11273);
xnor U12400 (N_12400,N_11690,N_11882);
nand U12401 (N_12401,N_11322,N_11458);
nand U12402 (N_12402,N_11667,N_11829);
xnor U12403 (N_12403,N_11774,N_11276);
and U12404 (N_12404,N_11507,N_11327);
nor U12405 (N_12405,N_11750,N_11596);
xor U12406 (N_12406,N_11547,N_11777);
nand U12407 (N_12407,N_11255,N_11377);
xor U12408 (N_12408,N_11687,N_11733);
nor U12409 (N_12409,N_11696,N_11295);
nor U12410 (N_12410,N_11872,N_11589);
nor U12411 (N_12411,N_11675,N_11673);
nand U12412 (N_12412,N_11959,N_11584);
xor U12413 (N_12413,N_11827,N_11584);
nor U12414 (N_12414,N_11391,N_11283);
or U12415 (N_12415,N_11439,N_11451);
xnor U12416 (N_12416,N_11669,N_11757);
and U12417 (N_12417,N_11714,N_11882);
nand U12418 (N_12418,N_11301,N_11875);
nor U12419 (N_12419,N_11645,N_11903);
xor U12420 (N_12420,N_11812,N_11533);
nor U12421 (N_12421,N_11451,N_11514);
or U12422 (N_12422,N_11999,N_11356);
nand U12423 (N_12423,N_11862,N_11926);
and U12424 (N_12424,N_11898,N_11723);
and U12425 (N_12425,N_11409,N_11782);
xnor U12426 (N_12426,N_11764,N_11964);
nor U12427 (N_12427,N_11419,N_11714);
nor U12428 (N_12428,N_11943,N_11764);
or U12429 (N_12429,N_11739,N_11633);
nand U12430 (N_12430,N_11333,N_11673);
xor U12431 (N_12431,N_11437,N_11292);
or U12432 (N_12432,N_11783,N_11413);
nand U12433 (N_12433,N_11559,N_11333);
or U12434 (N_12434,N_11779,N_11560);
xnor U12435 (N_12435,N_11571,N_11334);
or U12436 (N_12436,N_11766,N_11575);
nand U12437 (N_12437,N_11976,N_11969);
or U12438 (N_12438,N_11517,N_11401);
nor U12439 (N_12439,N_11685,N_11955);
xor U12440 (N_12440,N_11744,N_11945);
nor U12441 (N_12441,N_11420,N_11649);
nor U12442 (N_12442,N_11687,N_11296);
xnor U12443 (N_12443,N_11623,N_11669);
and U12444 (N_12444,N_11766,N_11659);
and U12445 (N_12445,N_11876,N_11862);
nand U12446 (N_12446,N_11654,N_11901);
nand U12447 (N_12447,N_11812,N_11585);
or U12448 (N_12448,N_11721,N_11738);
xnor U12449 (N_12449,N_11661,N_11927);
nand U12450 (N_12450,N_11341,N_11784);
xnor U12451 (N_12451,N_11785,N_11924);
nand U12452 (N_12452,N_11894,N_11370);
or U12453 (N_12453,N_11657,N_11884);
or U12454 (N_12454,N_11773,N_11464);
and U12455 (N_12455,N_11855,N_11495);
nand U12456 (N_12456,N_11458,N_11959);
nor U12457 (N_12457,N_11923,N_11346);
xor U12458 (N_12458,N_11702,N_11721);
nand U12459 (N_12459,N_11451,N_11472);
nand U12460 (N_12460,N_11279,N_11335);
nand U12461 (N_12461,N_11871,N_11889);
or U12462 (N_12462,N_11801,N_11272);
or U12463 (N_12463,N_11943,N_11767);
and U12464 (N_12464,N_11609,N_11965);
or U12465 (N_12465,N_11519,N_11264);
xor U12466 (N_12466,N_11625,N_11735);
and U12467 (N_12467,N_11754,N_11680);
and U12468 (N_12468,N_11781,N_11881);
xor U12469 (N_12469,N_11668,N_11414);
or U12470 (N_12470,N_11673,N_11913);
and U12471 (N_12471,N_11420,N_11602);
or U12472 (N_12472,N_11531,N_11638);
nand U12473 (N_12473,N_11436,N_11322);
nor U12474 (N_12474,N_11779,N_11633);
or U12475 (N_12475,N_11367,N_11709);
nor U12476 (N_12476,N_11763,N_11506);
xnor U12477 (N_12477,N_11934,N_11923);
or U12478 (N_12478,N_11317,N_11832);
xor U12479 (N_12479,N_11773,N_11994);
and U12480 (N_12480,N_11273,N_11342);
and U12481 (N_12481,N_11760,N_11398);
or U12482 (N_12482,N_11382,N_11390);
nor U12483 (N_12483,N_11329,N_11841);
nor U12484 (N_12484,N_11837,N_11976);
and U12485 (N_12485,N_11505,N_11791);
nand U12486 (N_12486,N_11346,N_11764);
and U12487 (N_12487,N_11795,N_11695);
and U12488 (N_12488,N_11782,N_11945);
or U12489 (N_12489,N_11990,N_11777);
nor U12490 (N_12490,N_11644,N_11714);
nor U12491 (N_12491,N_11609,N_11384);
nand U12492 (N_12492,N_11928,N_11970);
nand U12493 (N_12493,N_11430,N_11562);
and U12494 (N_12494,N_11748,N_11468);
nand U12495 (N_12495,N_11348,N_11765);
xnor U12496 (N_12496,N_11383,N_11442);
or U12497 (N_12497,N_11752,N_11974);
nor U12498 (N_12498,N_11314,N_11746);
nand U12499 (N_12499,N_11799,N_11807);
or U12500 (N_12500,N_11487,N_11997);
or U12501 (N_12501,N_11931,N_11637);
nand U12502 (N_12502,N_11923,N_11309);
and U12503 (N_12503,N_11440,N_11629);
and U12504 (N_12504,N_11390,N_11716);
and U12505 (N_12505,N_11465,N_11776);
or U12506 (N_12506,N_11711,N_11357);
nand U12507 (N_12507,N_11781,N_11978);
xnor U12508 (N_12508,N_11362,N_11817);
xnor U12509 (N_12509,N_11505,N_11605);
or U12510 (N_12510,N_11598,N_11773);
or U12511 (N_12511,N_11587,N_11720);
nand U12512 (N_12512,N_11413,N_11970);
xor U12513 (N_12513,N_11844,N_11792);
or U12514 (N_12514,N_11625,N_11347);
nor U12515 (N_12515,N_11706,N_11853);
xor U12516 (N_12516,N_11872,N_11815);
nor U12517 (N_12517,N_11532,N_11669);
nor U12518 (N_12518,N_11810,N_11939);
nor U12519 (N_12519,N_11930,N_11306);
nand U12520 (N_12520,N_11893,N_11493);
nand U12521 (N_12521,N_11419,N_11284);
and U12522 (N_12522,N_11476,N_11722);
and U12523 (N_12523,N_11723,N_11856);
or U12524 (N_12524,N_11858,N_11458);
and U12525 (N_12525,N_11992,N_11295);
and U12526 (N_12526,N_11942,N_11799);
and U12527 (N_12527,N_11386,N_11459);
and U12528 (N_12528,N_11568,N_11355);
xor U12529 (N_12529,N_11917,N_11921);
and U12530 (N_12530,N_11379,N_11566);
nor U12531 (N_12531,N_11322,N_11531);
and U12532 (N_12532,N_11946,N_11368);
and U12533 (N_12533,N_11462,N_11736);
nand U12534 (N_12534,N_11401,N_11425);
nand U12535 (N_12535,N_11603,N_11893);
or U12536 (N_12536,N_11564,N_11425);
xor U12537 (N_12537,N_11969,N_11578);
or U12538 (N_12538,N_11282,N_11951);
or U12539 (N_12539,N_11676,N_11308);
xnor U12540 (N_12540,N_11451,N_11709);
xnor U12541 (N_12541,N_11274,N_11449);
nand U12542 (N_12542,N_11276,N_11599);
xor U12543 (N_12543,N_11415,N_11421);
and U12544 (N_12544,N_11625,N_11794);
or U12545 (N_12545,N_11706,N_11377);
nor U12546 (N_12546,N_11301,N_11493);
or U12547 (N_12547,N_11998,N_11458);
nor U12548 (N_12548,N_11698,N_11711);
nor U12549 (N_12549,N_11619,N_11813);
nor U12550 (N_12550,N_11698,N_11890);
xor U12551 (N_12551,N_11362,N_11824);
nor U12552 (N_12552,N_11324,N_11832);
or U12553 (N_12553,N_11412,N_11924);
xor U12554 (N_12554,N_11505,N_11322);
or U12555 (N_12555,N_11488,N_11497);
or U12556 (N_12556,N_11477,N_11319);
nor U12557 (N_12557,N_11824,N_11898);
and U12558 (N_12558,N_11715,N_11367);
or U12559 (N_12559,N_11997,N_11744);
nor U12560 (N_12560,N_11551,N_11542);
and U12561 (N_12561,N_11764,N_11967);
or U12562 (N_12562,N_11420,N_11767);
and U12563 (N_12563,N_11614,N_11857);
or U12564 (N_12564,N_11283,N_11451);
xnor U12565 (N_12565,N_11986,N_11338);
nor U12566 (N_12566,N_11799,N_11904);
nor U12567 (N_12567,N_11541,N_11933);
xor U12568 (N_12568,N_11362,N_11506);
nor U12569 (N_12569,N_11351,N_11513);
xnor U12570 (N_12570,N_11868,N_11421);
nand U12571 (N_12571,N_11725,N_11886);
or U12572 (N_12572,N_11997,N_11675);
and U12573 (N_12573,N_11276,N_11994);
xor U12574 (N_12574,N_11508,N_11837);
or U12575 (N_12575,N_11362,N_11302);
or U12576 (N_12576,N_11353,N_11627);
or U12577 (N_12577,N_11318,N_11489);
nor U12578 (N_12578,N_11707,N_11948);
xnor U12579 (N_12579,N_11793,N_11856);
or U12580 (N_12580,N_11623,N_11832);
or U12581 (N_12581,N_11352,N_11620);
xor U12582 (N_12582,N_11431,N_11255);
nand U12583 (N_12583,N_11832,N_11738);
nor U12584 (N_12584,N_11530,N_11734);
nand U12585 (N_12585,N_11950,N_11812);
nor U12586 (N_12586,N_11879,N_11353);
or U12587 (N_12587,N_11884,N_11264);
nand U12588 (N_12588,N_11394,N_11602);
nand U12589 (N_12589,N_11751,N_11340);
nand U12590 (N_12590,N_11829,N_11627);
and U12591 (N_12591,N_11838,N_11408);
or U12592 (N_12592,N_11695,N_11899);
or U12593 (N_12593,N_11907,N_11503);
nor U12594 (N_12594,N_11811,N_11393);
nand U12595 (N_12595,N_11763,N_11758);
xnor U12596 (N_12596,N_11543,N_11843);
nand U12597 (N_12597,N_11420,N_11372);
or U12598 (N_12598,N_11405,N_11275);
nor U12599 (N_12599,N_11400,N_11443);
nor U12600 (N_12600,N_11297,N_11760);
nand U12601 (N_12601,N_11273,N_11414);
or U12602 (N_12602,N_11996,N_11859);
xnor U12603 (N_12603,N_11990,N_11421);
or U12604 (N_12604,N_11390,N_11955);
nand U12605 (N_12605,N_11556,N_11668);
and U12606 (N_12606,N_11905,N_11693);
and U12607 (N_12607,N_11301,N_11798);
or U12608 (N_12608,N_11291,N_11342);
nor U12609 (N_12609,N_11711,N_11967);
or U12610 (N_12610,N_11384,N_11307);
xor U12611 (N_12611,N_11454,N_11254);
and U12612 (N_12612,N_11906,N_11338);
and U12613 (N_12613,N_11250,N_11694);
or U12614 (N_12614,N_11704,N_11560);
and U12615 (N_12615,N_11669,N_11737);
or U12616 (N_12616,N_11392,N_11515);
or U12617 (N_12617,N_11362,N_11496);
or U12618 (N_12618,N_11625,N_11995);
and U12619 (N_12619,N_11740,N_11528);
nor U12620 (N_12620,N_11645,N_11503);
xnor U12621 (N_12621,N_11971,N_11782);
and U12622 (N_12622,N_11284,N_11899);
nand U12623 (N_12623,N_11888,N_11760);
or U12624 (N_12624,N_11424,N_11836);
nor U12625 (N_12625,N_11938,N_11731);
xor U12626 (N_12626,N_11391,N_11478);
xnor U12627 (N_12627,N_11298,N_11572);
and U12628 (N_12628,N_11276,N_11642);
nor U12629 (N_12629,N_11618,N_11971);
and U12630 (N_12630,N_11927,N_11942);
nor U12631 (N_12631,N_11296,N_11662);
and U12632 (N_12632,N_11577,N_11649);
and U12633 (N_12633,N_11293,N_11928);
or U12634 (N_12634,N_11869,N_11813);
or U12635 (N_12635,N_11725,N_11409);
nand U12636 (N_12636,N_11491,N_11594);
and U12637 (N_12637,N_11390,N_11642);
nand U12638 (N_12638,N_11636,N_11849);
and U12639 (N_12639,N_11378,N_11779);
nand U12640 (N_12640,N_11888,N_11648);
or U12641 (N_12641,N_11792,N_11350);
nand U12642 (N_12642,N_11722,N_11338);
nand U12643 (N_12643,N_11612,N_11415);
xnor U12644 (N_12644,N_11344,N_11564);
or U12645 (N_12645,N_11620,N_11845);
nand U12646 (N_12646,N_11802,N_11737);
or U12647 (N_12647,N_11818,N_11938);
xnor U12648 (N_12648,N_11873,N_11543);
nand U12649 (N_12649,N_11516,N_11801);
nor U12650 (N_12650,N_11609,N_11516);
nor U12651 (N_12651,N_11561,N_11949);
nand U12652 (N_12652,N_11669,N_11626);
and U12653 (N_12653,N_11526,N_11857);
xor U12654 (N_12654,N_11770,N_11600);
or U12655 (N_12655,N_11260,N_11877);
nor U12656 (N_12656,N_11292,N_11407);
xnor U12657 (N_12657,N_11345,N_11290);
nor U12658 (N_12658,N_11957,N_11682);
or U12659 (N_12659,N_11403,N_11802);
nor U12660 (N_12660,N_11889,N_11346);
xnor U12661 (N_12661,N_11695,N_11863);
nand U12662 (N_12662,N_11349,N_11859);
nand U12663 (N_12663,N_11852,N_11596);
nand U12664 (N_12664,N_11792,N_11400);
xor U12665 (N_12665,N_11412,N_11515);
or U12666 (N_12666,N_11305,N_11414);
xnor U12667 (N_12667,N_11977,N_11405);
nor U12668 (N_12668,N_11879,N_11341);
nor U12669 (N_12669,N_11586,N_11513);
or U12670 (N_12670,N_11515,N_11807);
nand U12671 (N_12671,N_11257,N_11309);
xnor U12672 (N_12672,N_11466,N_11324);
or U12673 (N_12673,N_11722,N_11988);
and U12674 (N_12674,N_11966,N_11496);
or U12675 (N_12675,N_11660,N_11484);
nor U12676 (N_12676,N_11725,N_11629);
nor U12677 (N_12677,N_11263,N_11557);
or U12678 (N_12678,N_11711,N_11258);
or U12679 (N_12679,N_11278,N_11495);
nand U12680 (N_12680,N_11913,N_11440);
and U12681 (N_12681,N_11391,N_11544);
nand U12682 (N_12682,N_11811,N_11449);
xnor U12683 (N_12683,N_11953,N_11583);
or U12684 (N_12684,N_11800,N_11642);
nand U12685 (N_12685,N_11485,N_11777);
xnor U12686 (N_12686,N_11767,N_11531);
or U12687 (N_12687,N_11739,N_11759);
nand U12688 (N_12688,N_11363,N_11779);
nand U12689 (N_12689,N_11717,N_11721);
and U12690 (N_12690,N_11460,N_11910);
nor U12691 (N_12691,N_11991,N_11740);
xnor U12692 (N_12692,N_11690,N_11643);
nor U12693 (N_12693,N_11791,N_11393);
xnor U12694 (N_12694,N_11859,N_11279);
or U12695 (N_12695,N_11607,N_11848);
and U12696 (N_12696,N_11854,N_11253);
xnor U12697 (N_12697,N_11686,N_11634);
nor U12698 (N_12698,N_11760,N_11379);
nand U12699 (N_12699,N_11997,N_11350);
or U12700 (N_12700,N_11870,N_11604);
nor U12701 (N_12701,N_11465,N_11995);
nand U12702 (N_12702,N_11901,N_11612);
or U12703 (N_12703,N_11399,N_11374);
xnor U12704 (N_12704,N_11854,N_11609);
nand U12705 (N_12705,N_11455,N_11453);
nor U12706 (N_12706,N_11879,N_11504);
or U12707 (N_12707,N_11738,N_11768);
nand U12708 (N_12708,N_11666,N_11279);
or U12709 (N_12709,N_11867,N_11474);
nor U12710 (N_12710,N_11652,N_11886);
or U12711 (N_12711,N_11254,N_11290);
nor U12712 (N_12712,N_11657,N_11914);
and U12713 (N_12713,N_11940,N_11758);
or U12714 (N_12714,N_11285,N_11412);
xor U12715 (N_12715,N_11688,N_11536);
nand U12716 (N_12716,N_11752,N_11876);
or U12717 (N_12717,N_11607,N_11498);
nor U12718 (N_12718,N_11891,N_11814);
or U12719 (N_12719,N_11476,N_11305);
nand U12720 (N_12720,N_11855,N_11404);
or U12721 (N_12721,N_11389,N_11948);
nand U12722 (N_12722,N_11378,N_11588);
nand U12723 (N_12723,N_11408,N_11463);
nor U12724 (N_12724,N_11362,N_11788);
xor U12725 (N_12725,N_11584,N_11772);
or U12726 (N_12726,N_11493,N_11835);
and U12727 (N_12727,N_11483,N_11503);
or U12728 (N_12728,N_11812,N_11911);
and U12729 (N_12729,N_11926,N_11653);
or U12730 (N_12730,N_11294,N_11580);
nand U12731 (N_12731,N_11462,N_11945);
and U12732 (N_12732,N_11857,N_11423);
and U12733 (N_12733,N_11554,N_11262);
xor U12734 (N_12734,N_11621,N_11825);
xnor U12735 (N_12735,N_11980,N_11361);
nor U12736 (N_12736,N_11319,N_11737);
xor U12737 (N_12737,N_11837,N_11321);
nor U12738 (N_12738,N_11932,N_11608);
nor U12739 (N_12739,N_11906,N_11735);
or U12740 (N_12740,N_11687,N_11633);
xor U12741 (N_12741,N_11532,N_11638);
or U12742 (N_12742,N_11445,N_11653);
and U12743 (N_12743,N_11858,N_11601);
nor U12744 (N_12744,N_11879,N_11258);
and U12745 (N_12745,N_11894,N_11828);
nand U12746 (N_12746,N_11531,N_11824);
nor U12747 (N_12747,N_11878,N_11416);
nand U12748 (N_12748,N_11682,N_11708);
and U12749 (N_12749,N_11436,N_11274);
and U12750 (N_12750,N_12735,N_12390);
xor U12751 (N_12751,N_12335,N_12315);
nand U12752 (N_12752,N_12068,N_12040);
xor U12753 (N_12753,N_12495,N_12314);
nand U12754 (N_12754,N_12233,N_12131);
nand U12755 (N_12755,N_12083,N_12457);
or U12756 (N_12756,N_12599,N_12052);
nor U12757 (N_12757,N_12522,N_12331);
nor U12758 (N_12758,N_12603,N_12373);
nand U12759 (N_12759,N_12125,N_12737);
and U12760 (N_12760,N_12254,N_12088);
xnor U12761 (N_12761,N_12329,N_12313);
or U12762 (N_12762,N_12643,N_12382);
xor U12763 (N_12763,N_12047,N_12702);
nor U12764 (N_12764,N_12187,N_12160);
and U12765 (N_12765,N_12654,N_12394);
or U12766 (N_12766,N_12053,N_12202);
and U12767 (N_12767,N_12708,N_12017);
or U12768 (N_12768,N_12296,N_12147);
nand U12769 (N_12769,N_12110,N_12176);
or U12770 (N_12770,N_12118,N_12551);
nand U12771 (N_12771,N_12220,N_12617);
and U12772 (N_12772,N_12606,N_12071);
or U12773 (N_12773,N_12289,N_12016);
or U12774 (N_12774,N_12662,N_12561);
nor U12775 (N_12775,N_12264,N_12489);
or U12776 (N_12776,N_12509,N_12531);
and U12777 (N_12777,N_12683,N_12007);
nand U12778 (N_12778,N_12598,N_12135);
nor U12779 (N_12779,N_12694,N_12341);
nor U12780 (N_12780,N_12615,N_12396);
nand U12781 (N_12781,N_12574,N_12405);
xor U12782 (N_12782,N_12387,N_12165);
nand U12783 (N_12783,N_12241,N_12723);
xor U12784 (N_12784,N_12043,N_12480);
and U12785 (N_12785,N_12089,N_12580);
nand U12786 (N_12786,N_12031,N_12228);
nor U12787 (N_12787,N_12065,N_12247);
nand U12788 (N_12788,N_12630,N_12577);
and U12789 (N_12789,N_12720,N_12347);
xnor U12790 (N_12790,N_12510,N_12297);
xnor U12791 (N_12791,N_12098,N_12651);
nand U12792 (N_12792,N_12116,N_12557);
nor U12793 (N_12793,N_12338,N_12463);
xnor U12794 (N_12794,N_12409,N_12403);
nand U12795 (N_12795,N_12020,N_12234);
nor U12796 (N_12796,N_12648,N_12140);
and U12797 (N_12797,N_12478,N_12177);
or U12798 (N_12798,N_12022,N_12719);
xnor U12799 (N_12799,N_12427,N_12129);
xor U12800 (N_12800,N_12466,N_12298);
nand U12801 (N_12801,N_12608,N_12721);
nand U12802 (N_12802,N_12182,N_12502);
nand U12803 (N_12803,N_12590,N_12079);
nor U12804 (N_12804,N_12487,N_12078);
xor U12805 (N_12805,N_12303,N_12733);
nand U12806 (N_12806,N_12404,N_12601);
xnor U12807 (N_12807,N_12265,N_12594);
or U12808 (N_12808,N_12475,N_12285);
nand U12809 (N_12809,N_12372,N_12205);
nand U12810 (N_12810,N_12467,N_12619);
xor U12811 (N_12811,N_12039,N_12240);
xor U12812 (N_12812,N_12092,N_12173);
xnor U12813 (N_12813,N_12628,N_12521);
nand U12814 (N_12814,N_12633,N_12159);
nor U12815 (N_12815,N_12326,N_12674);
nand U12816 (N_12816,N_12362,N_12414);
or U12817 (N_12817,N_12620,N_12048);
and U12818 (N_12818,N_12491,N_12639);
nor U12819 (N_12819,N_12516,N_12271);
and U12820 (N_12820,N_12622,N_12355);
xnor U12821 (N_12821,N_12056,N_12381);
or U12822 (N_12822,N_12525,N_12210);
or U12823 (N_12823,N_12357,N_12099);
and U12824 (N_12824,N_12520,N_12174);
and U12825 (N_12825,N_12268,N_12636);
nand U12826 (N_12826,N_12144,N_12400);
xnor U12827 (N_12827,N_12343,N_12380);
nor U12828 (N_12828,N_12003,N_12658);
or U12829 (N_12829,N_12739,N_12378);
nand U12830 (N_12830,N_12352,N_12600);
and U12831 (N_12831,N_12217,N_12232);
nand U12832 (N_12832,N_12703,N_12196);
or U12833 (N_12833,N_12740,N_12275);
and U12834 (N_12834,N_12449,N_12299);
xnor U12835 (N_12835,N_12340,N_12493);
and U12836 (N_12836,N_12519,N_12700);
or U12837 (N_12837,N_12255,N_12158);
and U12838 (N_12838,N_12416,N_12586);
xnor U12839 (N_12839,N_12153,N_12348);
and U12840 (N_12840,N_12459,N_12469);
and U12841 (N_12841,N_12245,N_12665);
nor U12842 (N_12842,N_12527,N_12582);
nor U12843 (N_12843,N_12269,N_12395);
nor U12844 (N_12844,N_12432,N_12709);
or U12845 (N_12845,N_12413,N_12670);
or U12846 (N_12846,N_12066,N_12446);
xnor U12847 (N_12847,N_12250,N_12011);
and U12848 (N_12848,N_12434,N_12441);
and U12849 (N_12849,N_12183,N_12034);
xor U12850 (N_12850,N_12682,N_12000);
or U12851 (N_12851,N_12081,N_12325);
or U12852 (N_12852,N_12455,N_12496);
nand U12853 (N_12853,N_12663,N_12744);
nor U12854 (N_12854,N_12545,N_12049);
or U12855 (N_12855,N_12345,N_12546);
or U12856 (N_12856,N_12472,N_12100);
nor U12857 (N_12857,N_12675,N_12587);
xnor U12858 (N_12858,N_12386,N_12536);
nand U12859 (N_12859,N_12625,N_12199);
or U12860 (N_12860,N_12529,N_12745);
nor U12861 (N_12861,N_12732,N_12393);
xnor U12862 (N_12862,N_12030,N_12517);
or U12863 (N_12863,N_12544,N_12318);
and U12864 (N_12864,N_12316,N_12481);
or U12865 (N_12865,N_12259,N_12293);
xnor U12866 (N_12866,N_12033,N_12181);
nand U12867 (N_12867,N_12686,N_12253);
xor U12868 (N_12868,N_12067,N_12164);
and U12869 (N_12869,N_12419,N_12283);
nor U12870 (N_12870,N_12638,N_12548);
or U12871 (N_12871,N_12488,N_12337);
nor U12872 (N_12872,N_12402,N_12330);
xnor U12873 (N_12873,N_12252,N_12659);
nand U12874 (N_12874,N_12503,N_12595);
xnor U12875 (N_12875,N_12554,N_12451);
nor U12876 (N_12876,N_12514,N_12621);
nor U12877 (N_12877,N_12421,N_12713);
or U12878 (N_12878,N_12399,N_12175);
and U12879 (N_12879,N_12374,N_12607);
xnor U12880 (N_12880,N_12422,N_12148);
xnor U12881 (N_12881,N_12440,N_12443);
nand U12882 (N_12882,N_12260,N_12353);
xnor U12883 (N_12883,N_12748,N_12311);
and U12884 (N_12884,N_12504,N_12149);
or U12885 (N_12885,N_12714,N_12684);
nor U12886 (N_12886,N_12500,N_12038);
nand U12887 (N_12887,N_12555,N_12257);
nand U12888 (N_12888,N_12547,N_12631);
and U12889 (N_12889,N_12146,N_12698);
xor U12890 (N_12890,N_12712,N_12741);
nand U12891 (N_12891,N_12192,N_12671);
nor U12892 (N_12892,N_12368,N_12470);
nor U12893 (N_12893,N_12024,N_12279);
nor U12894 (N_12894,N_12308,N_12219);
nand U12895 (N_12895,N_12157,N_12094);
nand U12896 (N_12896,N_12435,N_12108);
or U12897 (N_12897,N_12729,N_12431);
and U12898 (N_12898,N_12082,N_12305);
nand U12899 (N_12899,N_12239,N_12609);
or U12900 (N_12900,N_12201,N_12156);
xnor U12901 (N_12901,N_12602,N_12333);
nor U12902 (N_12902,N_12746,N_12074);
nor U12903 (N_12903,N_12623,N_12163);
xor U12904 (N_12904,N_12208,N_12019);
nor U12905 (N_12905,N_12666,N_12567);
nor U12906 (N_12906,N_12307,N_12121);
and U12907 (N_12907,N_12673,N_12013);
nand U12908 (N_12908,N_12236,N_12640);
nand U12909 (N_12909,N_12185,N_12650);
or U12910 (N_12910,N_12575,N_12632);
nor U12911 (N_12911,N_12055,N_12262);
nor U12912 (N_12912,N_12320,N_12282);
and U12913 (N_12913,N_12454,N_12653);
nor U12914 (N_12914,N_12730,N_12170);
xnor U12915 (N_12915,N_12218,N_12734);
nand U12916 (N_12916,N_12014,N_12501);
xnor U12917 (N_12917,N_12462,N_12354);
xor U12918 (N_12918,N_12699,N_12676);
or U12919 (N_12919,N_12072,N_12132);
or U12920 (N_12920,N_12476,N_12572);
nor U12921 (N_12921,N_12188,N_12407);
nand U12922 (N_12922,N_12090,N_12077);
nor U12923 (N_12923,N_12591,N_12154);
nand U12924 (N_12924,N_12562,N_12565);
xor U12925 (N_12925,N_12351,N_12678);
or U12926 (N_12926,N_12479,N_12634);
and U12927 (N_12927,N_12095,N_12592);
xnor U12928 (N_12928,N_12711,N_12581);
and U12929 (N_12929,N_12243,N_12292);
xnor U12930 (N_12930,N_12637,N_12012);
xnor U12931 (N_12931,N_12656,N_12226);
nand U12932 (N_12932,N_12359,N_12535);
or U12933 (N_12933,N_12685,N_12627);
or U12934 (N_12934,N_12191,N_12468);
and U12935 (N_12935,N_12109,N_12036);
xor U12936 (N_12936,N_12291,N_12687);
xor U12937 (N_12937,N_12123,N_12087);
and U12938 (N_12938,N_12589,N_12091);
nor U12939 (N_12939,N_12190,N_12346);
nor U12940 (N_12940,N_12689,N_12563);
or U12941 (N_12941,N_12126,N_12168);
nor U12942 (N_12942,N_12614,N_12041);
xnor U12943 (N_12943,N_12169,N_12725);
or U12944 (N_12944,N_12556,N_12178);
nand U12945 (N_12945,N_12101,N_12063);
nand U12946 (N_12946,N_12037,N_12568);
nor U12947 (N_12947,N_12626,N_12360);
xor U12948 (N_12948,N_12425,N_12447);
xnor U12949 (N_12949,N_12668,N_12417);
nor U12950 (N_12950,N_12552,N_12406);
xnor U12951 (N_12951,N_12366,N_12138);
and U12952 (N_12952,N_12695,N_12193);
nand U12953 (N_12953,N_12206,N_12515);
xnor U12954 (N_12954,N_12295,N_12005);
xor U12955 (N_12955,N_12198,N_12410);
and U12956 (N_12956,N_12073,N_12104);
nor U12957 (N_12957,N_12057,N_12223);
xor U12958 (N_12958,N_12322,N_12273);
nor U12959 (N_12959,N_12302,N_12278);
nand U12960 (N_12960,N_12549,N_12559);
or U12961 (N_12961,N_12161,N_12195);
nor U12962 (N_12962,N_12415,N_12106);
nand U12963 (N_12963,N_12513,N_12137);
and U12964 (N_12964,N_12306,N_12301);
or U12965 (N_12965,N_12122,N_12680);
xnor U12966 (N_12966,N_12616,N_12008);
and U12967 (N_12967,N_12566,N_12722);
nor U12968 (N_12968,N_12120,N_12604);
or U12969 (N_12969,N_12605,N_12576);
or U12970 (N_12970,N_12391,N_12113);
and U12971 (N_12971,N_12242,N_12032);
and U12972 (N_12972,N_12497,N_12704);
xnor U12973 (N_12973,N_12624,N_12726);
xor U12974 (N_12974,N_12076,N_12426);
and U12975 (N_12975,N_12213,N_12142);
nand U12976 (N_12976,N_12738,N_12485);
nor U12977 (N_12977,N_12436,N_12508);
nor U12978 (N_12978,N_12023,N_12115);
and U12979 (N_12979,N_12511,N_12060);
nor U12980 (N_12980,N_12618,N_12267);
xnor U12981 (N_12981,N_12444,N_12133);
nor U12982 (N_12982,N_12731,N_12539);
and U12983 (N_12983,N_12460,N_12166);
nor U12984 (N_12984,N_12474,N_12477);
or U12985 (N_12985,N_12482,N_12526);
or U12986 (N_12986,N_12179,N_12541);
or U12987 (N_12987,N_12494,N_12376);
xor U12988 (N_12988,N_12323,N_12681);
xor U12989 (N_12989,N_12224,N_12361);
nor U12990 (N_12990,N_12070,N_12385);
and U12991 (N_12991,N_12398,N_12742);
and U12992 (N_12992,N_12001,N_12246);
or U12993 (N_12993,N_12693,N_12180);
or U12994 (N_12994,N_12309,N_12710);
nor U12995 (N_12995,N_12507,N_12570);
and U12996 (N_12996,N_12184,N_12009);
nor U12997 (N_12997,N_12281,N_12028);
nor U12998 (N_12998,N_12097,N_12377);
and U12999 (N_12999,N_12050,N_12484);
or U13000 (N_13000,N_12613,N_12207);
nand U13001 (N_13001,N_12388,N_12743);
nand U13002 (N_13002,N_12237,N_12238);
nand U13003 (N_13003,N_12018,N_12445);
and U13004 (N_13004,N_12518,N_12270);
xor U13005 (N_13005,N_12736,N_12197);
and U13006 (N_13006,N_12465,N_12389);
and U13007 (N_13007,N_12543,N_12214);
nor U13008 (N_13008,N_12629,N_12061);
nor U13009 (N_13009,N_12652,N_12379);
or U13010 (N_13010,N_12528,N_12583);
nand U13011 (N_13011,N_12367,N_12274);
or U13012 (N_13012,N_12051,N_12369);
and U13013 (N_13013,N_12573,N_12134);
nor U13014 (N_13014,N_12408,N_12690);
xnor U13015 (N_13015,N_12046,N_12537);
nor U13016 (N_13016,N_12027,N_12375);
nand U13017 (N_13017,N_12006,N_12287);
or U13018 (N_13018,N_12571,N_12453);
nand U13019 (N_13019,N_12452,N_12429);
or U13020 (N_13020,N_12584,N_12433);
nand U13021 (N_13021,N_12215,N_12284);
and U13022 (N_13022,N_12141,N_12471);
nand U13023 (N_13023,N_12334,N_12171);
xnor U13024 (N_13024,N_12286,N_12204);
xor U13025 (N_13025,N_12715,N_12266);
or U13026 (N_13026,N_12450,N_12512);
and U13027 (N_13027,N_12080,N_12015);
xnor U13028 (N_13028,N_12718,N_12701);
nor U13029 (N_13029,N_12664,N_12438);
xor U13030 (N_13030,N_12263,N_12358);
xnor U13031 (N_13031,N_12442,N_12075);
xor U13032 (N_13032,N_12111,N_12747);
xor U13033 (N_13033,N_12096,N_12697);
nor U13034 (N_13034,N_12059,N_12064);
xnor U13035 (N_13035,N_12045,N_12578);
nand U13036 (N_13036,N_12212,N_12127);
nor U13037 (N_13037,N_12499,N_12716);
and U13038 (N_13038,N_12342,N_12216);
nor U13039 (N_13039,N_12130,N_12294);
nor U13040 (N_13040,N_12418,N_12054);
nor U13041 (N_13041,N_12401,N_12672);
nand U13042 (N_13042,N_12456,N_12117);
xor U13043 (N_13043,N_12200,N_12300);
nor U13044 (N_13044,N_12222,N_12610);
xor U13045 (N_13045,N_12107,N_12069);
nor U13046 (N_13046,N_12203,N_12588);
nand U13047 (N_13047,N_12114,N_12310);
and U13048 (N_13048,N_12439,N_12211);
xor U13049 (N_13049,N_12167,N_12277);
nand U13050 (N_13050,N_12724,N_12085);
and U13051 (N_13051,N_12327,N_12103);
and U13052 (N_13052,N_12251,N_12002);
xor U13053 (N_13053,N_12667,N_12538);
nor U13054 (N_13054,N_12370,N_12564);
nand U13055 (N_13055,N_12646,N_12363);
nand U13056 (N_13056,N_12423,N_12249);
nor U13057 (N_13057,N_12458,N_12151);
nand U13058 (N_13058,N_12428,N_12558);
or U13059 (N_13059,N_12026,N_12705);
nor U13060 (N_13060,N_12483,N_12533);
nor U13061 (N_13061,N_12044,N_12642);
nor U13062 (N_13062,N_12194,N_12657);
and U13063 (N_13063,N_12397,N_12498);
xnor U13064 (N_13064,N_12550,N_12280);
xor U13065 (N_13065,N_12448,N_12229);
nor U13066 (N_13066,N_12350,N_12145);
nand U13067 (N_13067,N_12492,N_12035);
nand U13068 (N_13068,N_12086,N_12688);
xnor U13069 (N_13069,N_12102,N_12025);
nand U13070 (N_13070,N_12231,N_12597);
xor U13071 (N_13071,N_12534,N_12655);
nand U13072 (N_13072,N_12542,N_12392);
and U13073 (N_13073,N_12505,N_12707);
nor U13074 (N_13074,N_12042,N_12244);
or U13075 (N_13075,N_12506,N_12084);
and U13076 (N_13076,N_12553,N_12230);
xnor U13077 (N_13077,N_12172,N_12349);
and U13078 (N_13078,N_12383,N_12649);
xor U13079 (N_13079,N_12706,N_12155);
nand U13080 (N_13080,N_12364,N_12124);
or U13081 (N_13081,N_12540,N_12532);
or U13082 (N_13082,N_12696,N_12225);
xor U13083 (N_13083,N_12611,N_12486);
nand U13084 (N_13084,N_12332,N_12569);
or U13085 (N_13085,N_12430,N_12585);
xor U13086 (N_13086,N_12344,N_12058);
and U13087 (N_13087,N_12523,N_12319);
xnor U13088 (N_13088,N_12660,N_12119);
or U13089 (N_13089,N_12143,N_12304);
nand U13090 (N_13090,N_12412,N_12136);
and U13091 (N_13091,N_12227,N_12596);
nand U13092 (N_13092,N_12221,N_12328);
nand U13093 (N_13093,N_12010,N_12692);
and U13094 (N_13094,N_12647,N_12644);
and U13095 (N_13095,N_12384,N_12717);
and U13096 (N_13096,N_12324,N_12464);
nor U13097 (N_13097,N_12029,N_12105);
or U13098 (N_13098,N_12560,N_12272);
nand U13099 (N_13099,N_12635,N_12162);
nor U13100 (N_13100,N_12579,N_12336);
xor U13101 (N_13101,N_12524,N_12727);
xor U13102 (N_13102,N_12290,N_12248);
or U13103 (N_13103,N_12186,N_12661);
and U13104 (N_13104,N_12490,N_12150);
nand U13105 (N_13105,N_12593,N_12139);
and U13106 (N_13106,N_12371,N_12189);
xnor U13107 (N_13107,N_12728,N_12093);
nor U13108 (N_13108,N_12112,N_12641);
xor U13109 (N_13109,N_12437,N_12004);
xnor U13110 (N_13110,N_12749,N_12021);
nor U13111 (N_13111,N_12062,N_12530);
or U13112 (N_13112,N_12256,N_12261);
nand U13113 (N_13113,N_12312,N_12677);
nand U13114 (N_13114,N_12235,N_12645);
nor U13115 (N_13115,N_12152,N_12258);
or U13116 (N_13116,N_12317,N_12321);
nand U13117 (N_13117,N_12209,N_12411);
xor U13118 (N_13118,N_12424,N_12365);
and U13119 (N_13119,N_12473,N_12679);
or U13120 (N_13120,N_12288,N_12128);
nor U13121 (N_13121,N_12691,N_12420);
and U13122 (N_13122,N_12461,N_12276);
and U13123 (N_13123,N_12339,N_12669);
or U13124 (N_13124,N_12356,N_12612);
or U13125 (N_13125,N_12531,N_12258);
xor U13126 (N_13126,N_12169,N_12437);
nand U13127 (N_13127,N_12233,N_12151);
and U13128 (N_13128,N_12221,N_12583);
and U13129 (N_13129,N_12481,N_12018);
nand U13130 (N_13130,N_12556,N_12442);
xnor U13131 (N_13131,N_12532,N_12677);
xor U13132 (N_13132,N_12589,N_12517);
and U13133 (N_13133,N_12480,N_12048);
nor U13134 (N_13134,N_12560,N_12161);
nor U13135 (N_13135,N_12230,N_12253);
or U13136 (N_13136,N_12224,N_12700);
nor U13137 (N_13137,N_12020,N_12007);
xnor U13138 (N_13138,N_12110,N_12724);
and U13139 (N_13139,N_12618,N_12071);
nand U13140 (N_13140,N_12059,N_12422);
nor U13141 (N_13141,N_12296,N_12308);
and U13142 (N_13142,N_12256,N_12711);
and U13143 (N_13143,N_12680,N_12219);
nand U13144 (N_13144,N_12639,N_12286);
and U13145 (N_13145,N_12633,N_12238);
xnor U13146 (N_13146,N_12443,N_12343);
and U13147 (N_13147,N_12622,N_12749);
nor U13148 (N_13148,N_12398,N_12190);
nor U13149 (N_13149,N_12002,N_12436);
xor U13150 (N_13150,N_12164,N_12112);
nor U13151 (N_13151,N_12165,N_12496);
nor U13152 (N_13152,N_12416,N_12025);
xnor U13153 (N_13153,N_12142,N_12541);
and U13154 (N_13154,N_12010,N_12165);
xor U13155 (N_13155,N_12456,N_12412);
and U13156 (N_13156,N_12301,N_12181);
and U13157 (N_13157,N_12496,N_12472);
xor U13158 (N_13158,N_12468,N_12523);
nor U13159 (N_13159,N_12296,N_12060);
nor U13160 (N_13160,N_12701,N_12498);
or U13161 (N_13161,N_12566,N_12218);
nor U13162 (N_13162,N_12646,N_12628);
or U13163 (N_13163,N_12487,N_12245);
and U13164 (N_13164,N_12713,N_12735);
nand U13165 (N_13165,N_12067,N_12210);
xnor U13166 (N_13166,N_12609,N_12071);
or U13167 (N_13167,N_12113,N_12233);
and U13168 (N_13168,N_12178,N_12706);
and U13169 (N_13169,N_12526,N_12748);
nand U13170 (N_13170,N_12634,N_12559);
or U13171 (N_13171,N_12068,N_12570);
xor U13172 (N_13172,N_12521,N_12207);
and U13173 (N_13173,N_12569,N_12289);
or U13174 (N_13174,N_12484,N_12677);
nand U13175 (N_13175,N_12631,N_12519);
nor U13176 (N_13176,N_12099,N_12029);
nor U13177 (N_13177,N_12352,N_12642);
xor U13178 (N_13178,N_12408,N_12185);
and U13179 (N_13179,N_12477,N_12687);
and U13180 (N_13180,N_12363,N_12694);
and U13181 (N_13181,N_12181,N_12195);
nor U13182 (N_13182,N_12101,N_12078);
or U13183 (N_13183,N_12435,N_12380);
or U13184 (N_13184,N_12577,N_12332);
or U13185 (N_13185,N_12186,N_12479);
xor U13186 (N_13186,N_12111,N_12358);
nor U13187 (N_13187,N_12055,N_12182);
nand U13188 (N_13188,N_12400,N_12695);
xor U13189 (N_13189,N_12731,N_12412);
xnor U13190 (N_13190,N_12240,N_12321);
xor U13191 (N_13191,N_12505,N_12419);
xor U13192 (N_13192,N_12564,N_12315);
and U13193 (N_13193,N_12018,N_12040);
xor U13194 (N_13194,N_12192,N_12640);
or U13195 (N_13195,N_12146,N_12438);
nand U13196 (N_13196,N_12719,N_12622);
and U13197 (N_13197,N_12167,N_12063);
and U13198 (N_13198,N_12502,N_12407);
xnor U13199 (N_13199,N_12449,N_12417);
xor U13200 (N_13200,N_12381,N_12022);
and U13201 (N_13201,N_12118,N_12629);
nand U13202 (N_13202,N_12350,N_12672);
nor U13203 (N_13203,N_12192,N_12647);
nor U13204 (N_13204,N_12738,N_12652);
nor U13205 (N_13205,N_12497,N_12073);
xor U13206 (N_13206,N_12676,N_12376);
nand U13207 (N_13207,N_12532,N_12577);
xnor U13208 (N_13208,N_12152,N_12581);
or U13209 (N_13209,N_12128,N_12247);
xor U13210 (N_13210,N_12719,N_12643);
nand U13211 (N_13211,N_12524,N_12169);
nand U13212 (N_13212,N_12060,N_12237);
nor U13213 (N_13213,N_12162,N_12579);
and U13214 (N_13214,N_12092,N_12059);
nor U13215 (N_13215,N_12704,N_12029);
xor U13216 (N_13216,N_12604,N_12067);
nand U13217 (N_13217,N_12232,N_12745);
xor U13218 (N_13218,N_12465,N_12093);
nand U13219 (N_13219,N_12406,N_12206);
nor U13220 (N_13220,N_12434,N_12175);
nand U13221 (N_13221,N_12033,N_12266);
or U13222 (N_13222,N_12387,N_12208);
xor U13223 (N_13223,N_12018,N_12267);
nand U13224 (N_13224,N_12139,N_12698);
nand U13225 (N_13225,N_12584,N_12409);
and U13226 (N_13226,N_12162,N_12308);
nor U13227 (N_13227,N_12749,N_12266);
and U13228 (N_13228,N_12667,N_12557);
or U13229 (N_13229,N_12429,N_12013);
or U13230 (N_13230,N_12399,N_12405);
and U13231 (N_13231,N_12301,N_12408);
nor U13232 (N_13232,N_12336,N_12240);
xnor U13233 (N_13233,N_12015,N_12329);
xnor U13234 (N_13234,N_12004,N_12055);
or U13235 (N_13235,N_12229,N_12228);
and U13236 (N_13236,N_12583,N_12508);
nand U13237 (N_13237,N_12520,N_12312);
xor U13238 (N_13238,N_12397,N_12585);
or U13239 (N_13239,N_12145,N_12160);
xor U13240 (N_13240,N_12494,N_12226);
or U13241 (N_13241,N_12309,N_12370);
or U13242 (N_13242,N_12268,N_12723);
and U13243 (N_13243,N_12238,N_12288);
xnor U13244 (N_13244,N_12070,N_12538);
and U13245 (N_13245,N_12196,N_12709);
and U13246 (N_13246,N_12197,N_12631);
nand U13247 (N_13247,N_12176,N_12538);
and U13248 (N_13248,N_12418,N_12740);
or U13249 (N_13249,N_12166,N_12375);
nand U13250 (N_13250,N_12350,N_12607);
nor U13251 (N_13251,N_12707,N_12628);
or U13252 (N_13252,N_12174,N_12279);
xor U13253 (N_13253,N_12060,N_12323);
xnor U13254 (N_13254,N_12311,N_12422);
or U13255 (N_13255,N_12020,N_12514);
nand U13256 (N_13256,N_12421,N_12130);
nor U13257 (N_13257,N_12000,N_12027);
or U13258 (N_13258,N_12495,N_12088);
and U13259 (N_13259,N_12267,N_12181);
or U13260 (N_13260,N_12129,N_12190);
or U13261 (N_13261,N_12008,N_12466);
or U13262 (N_13262,N_12165,N_12018);
xor U13263 (N_13263,N_12092,N_12354);
or U13264 (N_13264,N_12573,N_12007);
nor U13265 (N_13265,N_12281,N_12608);
or U13266 (N_13266,N_12427,N_12036);
nand U13267 (N_13267,N_12298,N_12136);
nor U13268 (N_13268,N_12112,N_12695);
or U13269 (N_13269,N_12277,N_12726);
nand U13270 (N_13270,N_12496,N_12152);
xor U13271 (N_13271,N_12456,N_12697);
nor U13272 (N_13272,N_12478,N_12129);
xor U13273 (N_13273,N_12539,N_12339);
and U13274 (N_13274,N_12679,N_12566);
and U13275 (N_13275,N_12224,N_12271);
xnor U13276 (N_13276,N_12011,N_12679);
xnor U13277 (N_13277,N_12187,N_12064);
and U13278 (N_13278,N_12681,N_12142);
and U13279 (N_13279,N_12444,N_12027);
or U13280 (N_13280,N_12642,N_12742);
nor U13281 (N_13281,N_12163,N_12512);
nand U13282 (N_13282,N_12067,N_12660);
nor U13283 (N_13283,N_12339,N_12481);
or U13284 (N_13284,N_12650,N_12245);
or U13285 (N_13285,N_12409,N_12443);
nand U13286 (N_13286,N_12187,N_12611);
and U13287 (N_13287,N_12439,N_12033);
and U13288 (N_13288,N_12434,N_12559);
or U13289 (N_13289,N_12595,N_12633);
and U13290 (N_13290,N_12522,N_12625);
or U13291 (N_13291,N_12513,N_12404);
or U13292 (N_13292,N_12023,N_12616);
xor U13293 (N_13293,N_12348,N_12063);
nand U13294 (N_13294,N_12553,N_12547);
nand U13295 (N_13295,N_12018,N_12100);
nor U13296 (N_13296,N_12327,N_12569);
nor U13297 (N_13297,N_12718,N_12216);
xnor U13298 (N_13298,N_12003,N_12416);
nand U13299 (N_13299,N_12579,N_12349);
nor U13300 (N_13300,N_12705,N_12652);
xor U13301 (N_13301,N_12056,N_12365);
or U13302 (N_13302,N_12242,N_12441);
xor U13303 (N_13303,N_12512,N_12197);
nand U13304 (N_13304,N_12498,N_12632);
or U13305 (N_13305,N_12590,N_12198);
nand U13306 (N_13306,N_12042,N_12248);
xor U13307 (N_13307,N_12256,N_12344);
or U13308 (N_13308,N_12536,N_12737);
xor U13309 (N_13309,N_12673,N_12550);
and U13310 (N_13310,N_12669,N_12039);
nand U13311 (N_13311,N_12162,N_12615);
nand U13312 (N_13312,N_12441,N_12413);
or U13313 (N_13313,N_12375,N_12570);
and U13314 (N_13314,N_12580,N_12013);
or U13315 (N_13315,N_12655,N_12356);
xnor U13316 (N_13316,N_12367,N_12193);
nor U13317 (N_13317,N_12613,N_12707);
or U13318 (N_13318,N_12665,N_12438);
nand U13319 (N_13319,N_12688,N_12060);
nor U13320 (N_13320,N_12009,N_12289);
and U13321 (N_13321,N_12178,N_12016);
nand U13322 (N_13322,N_12351,N_12698);
and U13323 (N_13323,N_12718,N_12406);
or U13324 (N_13324,N_12527,N_12738);
and U13325 (N_13325,N_12690,N_12630);
or U13326 (N_13326,N_12407,N_12199);
nand U13327 (N_13327,N_12694,N_12548);
nand U13328 (N_13328,N_12571,N_12056);
xnor U13329 (N_13329,N_12404,N_12139);
and U13330 (N_13330,N_12659,N_12314);
nor U13331 (N_13331,N_12042,N_12213);
nand U13332 (N_13332,N_12259,N_12341);
nor U13333 (N_13333,N_12197,N_12089);
and U13334 (N_13334,N_12463,N_12340);
and U13335 (N_13335,N_12654,N_12466);
xnor U13336 (N_13336,N_12743,N_12284);
or U13337 (N_13337,N_12290,N_12117);
nor U13338 (N_13338,N_12286,N_12292);
and U13339 (N_13339,N_12366,N_12214);
xor U13340 (N_13340,N_12436,N_12191);
and U13341 (N_13341,N_12260,N_12192);
or U13342 (N_13342,N_12020,N_12208);
or U13343 (N_13343,N_12655,N_12170);
xnor U13344 (N_13344,N_12227,N_12024);
xnor U13345 (N_13345,N_12116,N_12542);
and U13346 (N_13346,N_12083,N_12311);
and U13347 (N_13347,N_12045,N_12066);
xnor U13348 (N_13348,N_12120,N_12699);
or U13349 (N_13349,N_12110,N_12344);
nand U13350 (N_13350,N_12635,N_12308);
and U13351 (N_13351,N_12451,N_12475);
nor U13352 (N_13352,N_12552,N_12094);
nand U13353 (N_13353,N_12570,N_12034);
xnor U13354 (N_13354,N_12034,N_12188);
or U13355 (N_13355,N_12575,N_12433);
or U13356 (N_13356,N_12393,N_12033);
and U13357 (N_13357,N_12682,N_12418);
nand U13358 (N_13358,N_12315,N_12401);
nor U13359 (N_13359,N_12589,N_12685);
xor U13360 (N_13360,N_12629,N_12008);
xnor U13361 (N_13361,N_12333,N_12379);
nor U13362 (N_13362,N_12293,N_12294);
xnor U13363 (N_13363,N_12086,N_12238);
and U13364 (N_13364,N_12344,N_12029);
or U13365 (N_13365,N_12563,N_12389);
and U13366 (N_13366,N_12176,N_12626);
and U13367 (N_13367,N_12063,N_12226);
xor U13368 (N_13368,N_12255,N_12373);
and U13369 (N_13369,N_12123,N_12580);
nand U13370 (N_13370,N_12061,N_12319);
and U13371 (N_13371,N_12320,N_12281);
and U13372 (N_13372,N_12330,N_12294);
xnor U13373 (N_13373,N_12426,N_12683);
and U13374 (N_13374,N_12036,N_12372);
xnor U13375 (N_13375,N_12310,N_12013);
and U13376 (N_13376,N_12307,N_12041);
xnor U13377 (N_13377,N_12413,N_12738);
xnor U13378 (N_13378,N_12028,N_12342);
and U13379 (N_13379,N_12225,N_12128);
or U13380 (N_13380,N_12318,N_12588);
nand U13381 (N_13381,N_12685,N_12141);
xor U13382 (N_13382,N_12516,N_12596);
and U13383 (N_13383,N_12014,N_12241);
xnor U13384 (N_13384,N_12224,N_12525);
and U13385 (N_13385,N_12007,N_12146);
nor U13386 (N_13386,N_12150,N_12669);
nor U13387 (N_13387,N_12230,N_12032);
and U13388 (N_13388,N_12399,N_12543);
or U13389 (N_13389,N_12494,N_12566);
xor U13390 (N_13390,N_12434,N_12006);
nor U13391 (N_13391,N_12540,N_12669);
and U13392 (N_13392,N_12617,N_12479);
xor U13393 (N_13393,N_12066,N_12330);
nand U13394 (N_13394,N_12155,N_12144);
or U13395 (N_13395,N_12072,N_12146);
nor U13396 (N_13396,N_12490,N_12260);
xnor U13397 (N_13397,N_12035,N_12078);
and U13398 (N_13398,N_12399,N_12126);
nor U13399 (N_13399,N_12387,N_12705);
or U13400 (N_13400,N_12411,N_12627);
nand U13401 (N_13401,N_12242,N_12526);
xor U13402 (N_13402,N_12219,N_12611);
or U13403 (N_13403,N_12294,N_12512);
or U13404 (N_13404,N_12570,N_12581);
and U13405 (N_13405,N_12550,N_12336);
nor U13406 (N_13406,N_12015,N_12076);
and U13407 (N_13407,N_12738,N_12683);
xor U13408 (N_13408,N_12246,N_12710);
xnor U13409 (N_13409,N_12731,N_12510);
and U13410 (N_13410,N_12081,N_12296);
nand U13411 (N_13411,N_12071,N_12443);
and U13412 (N_13412,N_12352,N_12720);
and U13413 (N_13413,N_12416,N_12009);
nand U13414 (N_13414,N_12524,N_12454);
nor U13415 (N_13415,N_12205,N_12253);
nand U13416 (N_13416,N_12310,N_12351);
or U13417 (N_13417,N_12385,N_12482);
nor U13418 (N_13418,N_12069,N_12032);
xor U13419 (N_13419,N_12388,N_12010);
and U13420 (N_13420,N_12357,N_12196);
nand U13421 (N_13421,N_12528,N_12232);
or U13422 (N_13422,N_12156,N_12293);
nand U13423 (N_13423,N_12328,N_12214);
xor U13424 (N_13424,N_12439,N_12665);
nand U13425 (N_13425,N_12617,N_12449);
xor U13426 (N_13426,N_12589,N_12532);
nor U13427 (N_13427,N_12601,N_12364);
xor U13428 (N_13428,N_12312,N_12371);
or U13429 (N_13429,N_12536,N_12599);
nand U13430 (N_13430,N_12170,N_12628);
nor U13431 (N_13431,N_12077,N_12517);
nand U13432 (N_13432,N_12393,N_12320);
nor U13433 (N_13433,N_12629,N_12273);
nor U13434 (N_13434,N_12681,N_12476);
nor U13435 (N_13435,N_12705,N_12500);
xnor U13436 (N_13436,N_12543,N_12018);
or U13437 (N_13437,N_12174,N_12482);
and U13438 (N_13438,N_12287,N_12223);
and U13439 (N_13439,N_12102,N_12596);
and U13440 (N_13440,N_12455,N_12695);
and U13441 (N_13441,N_12412,N_12658);
nor U13442 (N_13442,N_12256,N_12376);
nor U13443 (N_13443,N_12684,N_12185);
nor U13444 (N_13444,N_12006,N_12162);
nand U13445 (N_13445,N_12309,N_12207);
and U13446 (N_13446,N_12519,N_12737);
nor U13447 (N_13447,N_12059,N_12463);
nor U13448 (N_13448,N_12326,N_12314);
or U13449 (N_13449,N_12610,N_12676);
or U13450 (N_13450,N_12117,N_12349);
nor U13451 (N_13451,N_12305,N_12239);
xnor U13452 (N_13452,N_12579,N_12603);
nand U13453 (N_13453,N_12248,N_12258);
or U13454 (N_13454,N_12638,N_12276);
nand U13455 (N_13455,N_12638,N_12337);
or U13456 (N_13456,N_12746,N_12288);
and U13457 (N_13457,N_12416,N_12510);
nor U13458 (N_13458,N_12680,N_12188);
or U13459 (N_13459,N_12482,N_12152);
and U13460 (N_13460,N_12303,N_12678);
xnor U13461 (N_13461,N_12131,N_12051);
and U13462 (N_13462,N_12264,N_12455);
nor U13463 (N_13463,N_12661,N_12402);
or U13464 (N_13464,N_12307,N_12172);
nor U13465 (N_13465,N_12494,N_12329);
or U13466 (N_13466,N_12151,N_12350);
nand U13467 (N_13467,N_12440,N_12516);
nand U13468 (N_13468,N_12231,N_12432);
and U13469 (N_13469,N_12249,N_12335);
nand U13470 (N_13470,N_12464,N_12674);
and U13471 (N_13471,N_12341,N_12640);
and U13472 (N_13472,N_12397,N_12614);
nor U13473 (N_13473,N_12076,N_12095);
or U13474 (N_13474,N_12012,N_12730);
xor U13475 (N_13475,N_12363,N_12136);
nand U13476 (N_13476,N_12623,N_12305);
nand U13477 (N_13477,N_12026,N_12423);
and U13478 (N_13478,N_12395,N_12643);
and U13479 (N_13479,N_12361,N_12450);
nand U13480 (N_13480,N_12035,N_12215);
xnor U13481 (N_13481,N_12020,N_12442);
xnor U13482 (N_13482,N_12431,N_12365);
or U13483 (N_13483,N_12096,N_12547);
xnor U13484 (N_13484,N_12718,N_12011);
nand U13485 (N_13485,N_12126,N_12224);
xor U13486 (N_13486,N_12269,N_12543);
xor U13487 (N_13487,N_12087,N_12453);
nor U13488 (N_13488,N_12657,N_12083);
xnor U13489 (N_13489,N_12237,N_12003);
nor U13490 (N_13490,N_12168,N_12252);
nor U13491 (N_13491,N_12258,N_12182);
xnor U13492 (N_13492,N_12682,N_12396);
or U13493 (N_13493,N_12661,N_12054);
nand U13494 (N_13494,N_12160,N_12143);
xor U13495 (N_13495,N_12287,N_12268);
nand U13496 (N_13496,N_12551,N_12464);
and U13497 (N_13497,N_12097,N_12020);
xnor U13498 (N_13498,N_12545,N_12087);
and U13499 (N_13499,N_12615,N_12029);
xor U13500 (N_13500,N_12998,N_12796);
nor U13501 (N_13501,N_13214,N_13139);
nor U13502 (N_13502,N_12783,N_13099);
and U13503 (N_13503,N_13351,N_12894);
or U13504 (N_13504,N_13280,N_12884);
nand U13505 (N_13505,N_13040,N_13465);
nor U13506 (N_13506,N_13007,N_13011);
and U13507 (N_13507,N_12814,N_13039);
and U13508 (N_13508,N_13388,N_12849);
or U13509 (N_13509,N_13485,N_13020);
and U13510 (N_13510,N_12953,N_13321);
nor U13511 (N_13511,N_13364,N_13279);
xor U13512 (N_13512,N_13329,N_12770);
or U13513 (N_13513,N_13356,N_13082);
or U13514 (N_13514,N_13486,N_13073);
nand U13515 (N_13515,N_13110,N_13259);
and U13516 (N_13516,N_13245,N_13322);
nor U13517 (N_13517,N_13103,N_13312);
nand U13518 (N_13518,N_13347,N_13059);
or U13519 (N_13519,N_12799,N_13105);
nand U13520 (N_13520,N_13025,N_13126);
nor U13521 (N_13521,N_13090,N_13019);
xor U13522 (N_13522,N_13392,N_13491);
nor U13523 (N_13523,N_13022,N_13004);
or U13524 (N_13524,N_13077,N_13436);
and U13525 (N_13525,N_13204,N_13151);
xnor U13526 (N_13526,N_13157,N_12981);
nand U13527 (N_13527,N_13201,N_13064);
nand U13528 (N_13528,N_13096,N_13104);
nor U13529 (N_13529,N_13313,N_13093);
nor U13530 (N_13530,N_13240,N_12776);
and U13531 (N_13531,N_13418,N_13235);
xnor U13532 (N_13532,N_13135,N_13424);
xnor U13533 (N_13533,N_12914,N_13206);
nand U13534 (N_13534,N_13297,N_13179);
or U13535 (N_13535,N_13137,N_12948);
and U13536 (N_13536,N_12844,N_13127);
nand U13537 (N_13537,N_13468,N_13480);
nand U13538 (N_13538,N_13397,N_13097);
xor U13539 (N_13539,N_13370,N_12790);
and U13540 (N_13540,N_13407,N_13042);
nor U13541 (N_13541,N_13063,N_13456);
xnor U13542 (N_13542,N_12838,N_13426);
xnor U13543 (N_13543,N_12843,N_13402);
and U13544 (N_13544,N_13215,N_12797);
or U13545 (N_13545,N_12867,N_13242);
xnor U13546 (N_13546,N_12836,N_12754);
nor U13547 (N_13547,N_13287,N_13267);
nand U13548 (N_13548,N_13053,N_13116);
or U13549 (N_13549,N_12777,N_12779);
or U13550 (N_13550,N_12831,N_13270);
or U13551 (N_13551,N_13335,N_13254);
or U13552 (N_13552,N_13078,N_13274);
and U13553 (N_13553,N_12958,N_13412);
nand U13554 (N_13554,N_12971,N_13476);
or U13555 (N_13555,N_13405,N_13479);
and U13556 (N_13556,N_13396,N_13293);
and U13557 (N_13557,N_12815,N_12966);
or U13558 (N_13558,N_12890,N_12988);
nor U13559 (N_13559,N_13380,N_12905);
or U13560 (N_13560,N_12899,N_12828);
or U13561 (N_13561,N_12871,N_13339);
nand U13562 (N_13562,N_13155,N_13271);
nand U13563 (N_13563,N_12888,N_12909);
or U13564 (N_13564,N_13145,N_13186);
xor U13565 (N_13565,N_13140,N_12829);
or U13566 (N_13566,N_13216,N_13406);
and U13567 (N_13567,N_13469,N_13441);
nor U13568 (N_13568,N_12937,N_12985);
xor U13569 (N_13569,N_13049,N_12850);
nor U13570 (N_13570,N_12907,N_13081);
nand U13571 (N_13571,N_12978,N_13260);
xor U13572 (N_13572,N_13171,N_12835);
or U13573 (N_13573,N_13269,N_12932);
nor U13574 (N_13574,N_12913,N_12979);
nand U13575 (N_13575,N_13141,N_12855);
xor U13576 (N_13576,N_12812,N_12986);
or U13577 (N_13577,N_12859,N_13289);
or U13578 (N_13578,N_12788,N_13316);
nand U13579 (N_13579,N_13354,N_13144);
and U13580 (N_13580,N_12769,N_12969);
nor U13581 (N_13581,N_12804,N_12865);
nand U13582 (N_13582,N_13168,N_13383);
or U13583 (N_13583,N_12918,N_13319);
or U13584 (N_13584,N_12980,N_13332);
nor U13585 (N_13585,N_13102,N_13336);
nand U13586 (N_13586,N_12870,N_13047);
and U13587 (N_13587,N_12886,N_13180);
nand U13588 (N_13588,N_13275,N_13299);
or U13589 (N_13589,N_13266,N_13068);
or U13590 (N_13590,N_13146,N_13000);
nor U13591 (N_13591,N_13061,N_13188);
and U13592 (N_13592,N_13443,N_13067);
nand U13593 (N_13593,N_13372,N_13331);
nand U13594 (N_13594,N_12892,N_13130);
xnor U13595 (N_13595,N_12816,N_12781);
nand U13596 (N_13596,N_12996,N_13300);
nor U13597 (N_13597,N_13492,N_13163);
and U13598 (N_13598,N_13337,N_12873);
nor U13599 (N_13599,N_13328,N_13379);
nor U13600 (N_13600,N_13375,N_12938);
nor U13601 (N_13601,N_13109,N_12990);
or U13602 (N_13602,N_13374,N_13400);
and U13603 (N_13603,N_12847,N_13410);
nand U13604 (N_13604,N_13419,N_13481);
xnor U13605 (N_13605,N_13341,N_13199);
and U13606 (N_13606,N_12837,N_12992);
xor U13607 (N_13607,N_13236,N_12911);
nand U13608 (N_13608,N_13449,N_12910);
nand U13609 (N_13609,N_13248,N_13220);
or U13610 (N_13610,N_13307,N_13015);
or U13611 (N_13611,N_12868,N_13045);
xnor U13612 (N_13612,N_12832,N_13393);
and U13613 (N_13613,N_12919,N_13390);
nor U13614 (N_13614,N_13094,N_12750);
nand U13615 (N_13615,N_12775,N_12945);
or U13616 (N_13616,N_13303,N_13273);
xnor U13617 (N_13617,N_12771,N_12951);
xor U13618 (N_13618,N_13205,N_13376);
or U13619 (N_13619,N_13177,N_13498);
xor U13620 (N_13620,N_12944,N_13320);
xnor U13621 (N_13621,N_13120,N_13043);
nand U13622 (N_13622,N_12830,N_13461);
nand U13623 (N_13623,N_13255,N_13253);
and U13624 (N_13624,N_13474,N_12752);
nor U13625 (N_13625,N_13311,N_13262);
and U13626 (N_13626,N_12921,N_12813);
nor U13627 (N_13627,N_12784,N_13089);
or U13628 (N_13628,N_13355,N_13080);
xor U13629 (N_13629,N_12763,N_13198);
nor U13630 (N_13630,N_12874,N_13478);
xnor U13631 (N_13631,N_13249,N_13119);
nand U13632 (N_13632,N_12927,N_12853);
xor U13633 (N_13633,N_12760,N_13176);
or U13634 (N_13634,N_13203,N_13340);
or U13635 (N_13635,N_12798,N_13452);
or U13636 (N_13636,N_13472,N_13010);
nand U13637 (N_13637,N_13184,N_13238);
nand U13638 (N_13638,N_13359,N_13243);
nand U13639 (N_13639,N_13079,N_13463);
or U13640 (N_13640,N_13378,N_13401);
and U13641 (N_13641,N_12972,N_12876);
nor U13642 (N_13642,N_13453,N_13489);
xor U13643 (N_13643,N_13363,N_13098);
nand U13644 (N_13644,N_13034,N_13024);
nor U13645 (N_13645,N_13288,N_13108);
or U13646 (N_13646,N_13228,N_12900);
xnor U13647 (N_13647,N_13369,N_13175);
xor U13648 (N_13648,N_12935,N_13387);
or U13649 (N_13649,N_13128,N_12964);
nand U13650 (N_13650,N_13055,N_12960);
or U13651 (N_13651,N_13324,N_13434);
or U13652 (N_13652,N_12807,N_13196);
xnor U13653 (N_13653,N_13241,N_13033);
or U13654 (N_13654,N_12977,N_13191);
and U13655 (N_13655,N_13227,N_13437);
and U13656 (N_13656,N_12802,N_13352);
xnor U13657 (N_13657,N_12933,N_13057);
or U13658 (N_13658,N_13246,N_13430);
xor U13659 (N_13659,N_13484,N_13030);
and U13660 (N_13660,N_12925,N_13185);
xor U13661 (N_13661,N_13031,N_13281);
or U13662 (N_13662,N_13394,N_13423);
nand U13663 (N_13663,N_12878,N_12952);
xor U13664 (N_13664,N_13237,N_13302);
xnor U13665 (N_13665,N_12756,N_13391);
nor U13666 (N_13666,N_13048,N_12778);
nor U13667 (N_13667,N_12869,N_12872);
and U13668 (N_13668,N_13173,N_13226);
or U13669 (N_13669,N_13131,N_13368);
nand U13670 (N_13670,N_13360,N_13425);
xor U13671 (N_13671,N_13165,N_12846);
and U13672 (N_13672,N_13017,N_13195);
nor U13673 (N_13673,N_12936,N_13471);
and U13674 (N_13674,N_13252,N_13085);
nand U13675 (N_13675,N_13134,N_13366);
or U13676 (N_13676,N_12864,N_13385);
nor U13677 (N_13677,N_13207,N_13159);
xor U13678 (N_13678,N_12800,N_13003);
and U13679 (N_13679,N_13219,N_13052);
nor U13680 (N_13680,N_13037,N_13314);
nand U13681 (N_13681,N_12801,N_12924);
and U13682 (N_13682,N_12811,N_13482);
and U13683 (N_13683,N_13349,N_13218);
xnor U13684 (N_13684,N_13161,N_13247);
or U13685 (N_13685,N_12955,N_13125);
nor U13686 (N_13686,N_13038,N_13149);
or U13687 (N_13687,N_13428,N_13286);
nand U13688 (N_13688,N_12857,N_13106);
nor U13689 (N_13689,N_13263,N_13118);
or U13690 (N_13690,N_13028,N_13202);
and U13691 (N_13691,N_12904,N_13451);
xor U13692 (N_13692,N_12787,N_13101);
nand U13693 (N_13693,N_13092,N_12947);
and U13694 (N_13694,N_12842,N_12789);
nand U13695 (N_13695,N_12968,N_12758);
xor U13696 (N_13696,N_13362,N_13413);
xnor U13697 (N_13697,N_13470,N_13348);
and U13698 (N_13698,N_12908,N_12889);
nand U13699 (N_13699,N_12875,N_13225);
xnor U13700 (N_13700,N_12755,N_13233);
or U13701 (N_13701,N_12896,N_13071);
nor U13702 (N_13702,N_13495,N_13261);
and U13703 (N_13703,N_12768,N_13301);
xor U13704 (N_13704,N_13256,N_12922);
nand U13705 (N_13705,N_12792,N_12950);
nor U13706 (N_13706,N_13292,N_13147);
or U13707 (N_13707,N_13295,N_13018);
and U13708 (N_13708,N_13072,N_13084);
nand U13709 (N_13709,N_13200,N_13066);
nand U13710 (N_13710,N_13386,N_13095);
and U13711 (N_13711,N_13291,N_13210);
nand U13712 (N_13712,N_13221,N_13111);
nor U13713 (N_13713,N_13395,N_13076);
nor U13714 (N_13714,N_13169,N_13258);
and U13715 (N_13715,N_13150,N_12824);
nand U13716 (N_13716,N_13239,N_13283);
nand U13717 (N_13717,N_13193,N_13234);
and U13718 (N_13718,N_12963,N_13070);
nor U13719 (N_13719,N_13431,N_13464);
xnor U13720 (N_13720,N_12965,N_13488);
nand U13721 (N_13721,N_12994,N_13083);
or U13722 (N_13722,N_13467,N_13427);
or U13723 (N_13723,N_13277,N_13035);
nor U13724 (N_13724,N_13009,N_12803);
and U13725 (N_13725,N_12791,N_12767);
and U13726 (N_13726,N_13317,N_13309);
and U13727 (N_13727,N_12840,N_12785);
nor U13728 (N_13728,N_13115,N_12795);
nor U13729 (N_13729,N_13075,N_13244);
and U13730 (N_13730,N_13276,N_13044);
and U13731 (N_13731,N_13357,N_13432);
or U13732 (N_13732,N_13058,N_13483);
or U13733 (N_13733,N_12780,N_13497);
xnor U13734 (N_13734,N_12833,N_12772);
and U13735 (N_13735,N_13284,N_12821);
nand U13736 (N_13736,N_13222,N_13230);
and U13737 (N_13737,N_13123,N_13384);
xnor U13738 (N_13738,N_13152,N_13326);
and U13739 (N_13739,N_13499,N_13250);
nand U13740 (N_13740,N_13416,N_12881);
or U13741 (N_13741,N_13409,N_12962);
or U13742 (N_13742,N_13315,N_13477);
nor U13743 (N_13743,N_13433,N_12982);
xor U13744 (N_13744,N_13178,N_13345);
xnor U13745 (N_13745,N_12826,N_13208);
nor U13746 (N_13746,N_13087,N_13389);
or U13747 (N_13747,N_12995,N_12851);
or U13748 (N_13748,N_12860,N_13414);
xnor U13749 (N_13749,N_13408,N_13023);
and U13750 (N_13750,N_12926,N_13358);
nor U13751 (N_13751,N_12946,N_12761);
nor U13752 (N_13752,N_13466,N_12957);
nand U13753 (N_13753,N_12764,N_13310);
and U13754 (N_13754,N_12753,N_13422);
nor U13755 (N_13755,N_13367,N_12757);
nand U13756 (N_13756,N_13455,N_12806);
or U13757 (N_13757,N_12928,N_13181);
nand U13758 (N_13758,N_12929,N_13026);
xnor U13759 (N_13759,N_13458,N_13330);
nand U13760 (N_13760,N_12923,N_13382);
and U13761 (N_13761,N_12970,N_12765);
and U13762 (N_13762,N_13197,N_12939);
and U13763 (N_13763,N_12861,N_13121);
and U13764 (N_13764,N_12759,N_13448);
xnor U13765 (N_13765,N_12931,N_13027);
and U13766 (N_13766,N_13088,N_13100);
or U13767 (N_13767,N_12906,N_13403);
nand U13768 (N_13768,N_12997,N_12819);
nor U13769 (N_13769,N_12794,N_13074);
nand U13770 (N_13770,N_13166,N_13264);
xnor U13771 (N_13771,N_12920,N_13129);
xor U13772 (N_13772,N_12984,N_12858);
xnor U13773 (N_13773,N_13398,N_13122);
and U13774 (N_13774,N_13132,N_12827);
and U13775 (N_13775,N_13056,N_13444);
nand U13776 (N_13776,N_12974,N_13306);
and U13777 (N_13777,N_13373,N_13346);
nand U13778 (N_13778,N_13232,N_13170);
xor U13779 (N_13779,N_13381,N_13183);
or U13780 (N_13780,N_13429,N_13016);
or U13781 (N_13781,N_13142,N_13174);
xnor U13782 (N_13782,N_12885,N_13377);
nand U13783 (N_13783,N_13029,N_13411);
or U13784 (N_13784,N_12893,N_12852);
xnor U13785 (N_13785,N_12882,N_12810);
xnor U13786 (N_13786,N_13327,N_13005);
nor U13787 (N_13787,N_12967,N_13445);
and U13788 (N_13788,N_13278,N_13365);
nand U13789 (N_13789,N_13399,N_12941);
nor U13790 (N_13790,N_13194,N_12897);
xor U13791 (N_13791,N_13117,N_12880);
xnor U13792 (N_13792,N_13323,N_13060);
nand U13793 (N_13793,N_13334,N_12902);
and U13794 (N_13794,N_12895,N_12866);
or U13795 (N_13795,N_13006,N_12999);
or U13796 (N_13796,N_12766,N_13211);
or U13797 (N_13797,N_12993,N_13344);
or U13798 (N_13798,N_13107,N_12973);
nor U13799 (N_13799,N_12976,N_13493);
nor U13800 (N_13800,N_12903,N_12863);
or U13801 (N_13801,N_13002,N_13473);
nand U13802 (N_13802,N_12773,N_12959);
xor U13803 (N_13803,N_12949,N_12912);
nand U13804 (N_13804,N_13156,N_13308);
xor U13805 (N_13805,N_12877,N_13350);
xnor U13806 (N_13806,N_12883,N_13272);
nand U13807 (N_13807,N_13475,N_12916);
and U13808 (N_13808,N_13187,N_13054);
nor U13809 (N_13809,N_13172,N_12845);
nand U13810 (N_13810,N_12887,N_12901);
nand U13811 (N_13811,N_12879,N_13138);
nor U13812 (N_13812,N_13217,N_13167);
or U13813 (N_13813,N_13012,N_12841);
xnor U13814 (N_13814,N_13421,N_13086);
nand U13815 (N_13815,N_13298,N_13143);
and U13816 (N_13816,N_13268,N_12956);
xor U13817 (N_13817,N_12762,N_13153);
and U13818 (N_13818,N_13459,N_12954);
nor U13819 (N_13819,N_13442,N_13189);
and U13820 (N_13820,N_13457,N_13305);
or U13821 (N_13821,N_12917,N_13133);
nor U13822 (N_13822,N_13154,N_13282);
or U13823 (N_13823,N_13257,N_13001);
xnor U13824 (N_13824,N_13136,N_13251);
and U13825 (N_13825,N_12915,N_13371);
xor U13826 (N_13826,N_13091,N_13190);
and U13827 (N_13827,N_13342,N_13041);
or U13828 (N_13828,N_12822,N_13450);
or U13829 (N_13829,N_13062,N_12751);
xor U13830 (N_13830,N_13318,N_13008);
or U13831 (N_13831,N_12991,N_13046);
or U13832 (N_13832,N_12786,N_12862);
xor U13833 (N_13833,N_13294,N_12823);
nand U13834 (N_13834,N_13021,N_13229);
nor U13835 (N_13835,N_12808,N_13494);
nor U13836 (N_13836,N_13487,N_12820);
xnor U13837 (N_13837,N_13265,N_12898);
or U13838 (N_13838,N_12934,N_13446);
or U13839 (N_13839,N_13404,N_13013);
nor U13840 (N_13840,N_12825,N_13112);
or U13841 (N_13841,N_13113,N_13438);
nor U13842 (N_13842,N_12983,N_12817);
nand U13843 (N_13843,N_12854,N_13209);
or U13844 (N_13844,N_13338,N_13182);
or U13845 (N_13845,N_12793,N_13420);
nand U13846 (N_13846,N_12930,N_12774);
and U13847 (N_13847,N_13032,N_13343);
or U13848 (N_13848,N_13454,N_13148);
nand U13849 (N_13849,N_13417,N_13164);
nor U13850 (N_13850,N_13069,N_12942);
and U13851 (N_13851,N_13440,N_13415);
nand U13852 (N_13852,N_13231,N_12891);
or U13853 (N_13853,N_13462,N_13158);
nand U13854 (N_13854,N_13285,N_12856);
and U13855 (N_13855,N_12782,N_12809);
xnor U13856 (N_13856,N_13304,N_13162);
nor U13857 (N_13857,N_13460,N_12943);
and U13858 (N_13858,N_13361,N_13224);
xnor U13859 (N_13859,N_12834,N_13333);
or U13860 (N_13860,N_13050,N_13160);
xor U13861 (N_13861,N_13435,N_13439);
and U13862 (N_13862,N_13212,N_13490);
nor U13863 (N_13863,N_13325,N_12805);
xor U13864 (N_13864,N_12961,N_13192);
and U13865 (N_13865,N_13353,N_12987);
or U13866 (N_13866,N_13223,N_12839);
nand U13867 (N_13867,N_13065,N_13036);
or U13868 (N_13868,N_12989,N_13051);
xor U13869 (N_13869,N_12818,N_12848);
xor U13870 (N_13870,N_13124,N_13114);
and U13871 (N_13871,N_13296,N_13290);
xor U13872 (N_13872,N_12940,N_13014);
nor U13873 (N_13873,N_13496,N_12975);
nor U13874 (N_13874,N_13447,N_13213);
or U13875 (N_13875,N_13419,N_12873);
nor U13876 (N_13876,N_13141,N_13359);
xnor U13877 (N_13877,N_12933,N_13396);
nor U13878 (N_13878,N_13000,N_13394);
or U13879 (N_13879,N_13499,N_13358);
nand U13880 (N_13880,N_13030,N_13365);
and U13881 (N_13881,N_13070,N_13452);
nand U13882 (N_13882,N_13074,N_13324);
and U13883 (N_13883,N_13272,N_13301);
nand U13884 (N_13884,N_12993,N_13464);
and U13885 (N_13885,N_13294,N_13458);
nor U13886 (N_13886,N_13354,N_12986);
and U13887 (N_13887,N_13242,N_12980);
xor U13888 (N_13888,N_12906,N_13340);
or U13889 (N_13889,N_13356,N_13478);
nor U13890 (N_13890,N_13450,N_12995);
or U13891 (N_13891,N_12777,N_13101);
and U13892 (N_13892,N_13439,N_12996);
xnor U13893 (N_13893,N_12833,N_13112);
nor U13894 (N_13894,N_12938,N_13320);
nor U13895 (N_13895,N_13236,N_12902);
or U13896 (N_13896,N_13295,N_12753);
nand U13897 (N_13897,N_13322,N_12840);
nand U13898 (N_13898,N_12975,N_12838);
xor U13899 (N_13899,N_12904,N_13297);
and U13900 (N_13900,N_13354,N_13214);
and U13901 (N_13901,N_13384,N_13031);
nand U13902 (N_13902,N_13309,N_12766);
or U13903 (N_13903,N_13181,N_12969);
nor U13904 (N_13904,N_13043,N_12833);
or U13905 (N_13905,N_13123,N_13099);
nand U13906 (N_13906,N_13400,N_13464);
and U13907 (N_13907,N_12770,N_13405);
nor U13908 (N_13908,N_13405,N_13252);
nor U13909 (N_13909,N_12949,N_13321);
nand U13910 (N_13910,N_13096,N_13039);
nor U13911 (N_13911,N_12766,N_12900);
nor U13912 (N_13912,N_13185,N_12858);
or U13913 (N_13913,N_13464,N_13339);
nor U13914 (N_13914,N_12857,N_13007);
nor U13915 (N_13915,N_13183,N_13239);
xnor U13916 (N_13916,N_12755,N_12919);
and U13917 (N_13917,N_12817,N_13043);
and U13918 (N_13918,N_13092,N_13355);
nand U13919 (N_13919,N_13091,N_13117);
xor U13920 (N_13920,N_13081,N_12857);
or U13921 (N_13921,N_13245,N_13135);
xor U13922 (N_13922,N_13441,N_13428);
nor U13923 (N_13923,N_13083,N_12860);
xor U13924 (N_13924,N_13432,N_12857);
and U13925 (N_13925,N_12852,N_12949);
or U13926 (N_13926,N_13189,N_13401);
nor U13927 (N_13927,N_13025,N_13466);
and U13928 (N_13928,N_12753,N_13133);
xor U13929 (N_13929,N_13370,N_12955);
nor U13930 (N_13930,N_13203,N_13044);
xnor U13931 (N_13931,N_13112,N_13012);
and U13932 (N_13932,N_13299,N_12765);
or U13933 (N_13933,N_12963,N_13289);
and U13934 (N_13934,N_12809,N_12986);
and U13935 (N_13935,N_13459,N_13011);
nand U13936 (N_13936,N_12902,N_12912);
nor U13937 (N_13937,N_12912,N_12768);
xnor U13938 (N_13938,N_13438,N_13323);
or U13939 (N_13939,N_12941,N_13486);
nor U13940 (N_13940,N_13472,N_13471);
nand U13941 (N_13941,N_13375,N_13409);
or U13942 (N_13942,N_13157,N_13028);
nor U13943 (N_13943,N_12782,N_13241);
and U13944 (N_13944,N_13376,N_12831);
and U13945 (N_13945,N_13300,N_13433);
or U13946 (N_13946,N_13373,N_13084);
or U13947 (N_13947,N_12899,N_12950);
xnor U13948 (N_13948,N_12812,N_13094);
or U13949 (N_13949,N_13260,N_12884);
xor U13950 (N_13950,N_13172,N_12834);
nand U13951 (N_13951,N_12865,N_13014);
xnor U13952 (N_13952,N_13221,N_12953);
nor U13953 (N_13953,N_12949,N_13168);
and U13954 (N_13954,N_13181,N_12923);
or U13955 (N_13955,N_13279,N_13233);
xor U13956 (N_13956,N_12920,N_13155);
nor U13957 (N_13957,N_13465,N_13048);
xor U13958 (N_13958,N_12803,N_13094);
and U13959 (N_13959,N_13370,N_13171);
nand U13960 (N_13960,N_13339,N_12980);
nand U13961 (N_13961,N_13466,N_13171);
nand U13962 (N_13962,N_12797,N_13150);
or U13963 (N_13963,N_12799,N_12828);
nor U13964 (N_13964,N_12856,N_12974);
or U13965 (N_13965,N_13110,N_12974);
and U13966 (N_13966,N_13076,N_13457);
nor U13967 (N_13967,N_13277,N_13354);
nor U13968 (N_13968,N_12774,N_13411);
nor U13969 (N_13969,N_13315,N_13388);
nor U13970 (N_13970,N_13366,N_13349);
nand U13971 (N_13971,N_13429,N_12906);
nor U13972 (N_13972,N_13009,N_13116);
nand U13973 (N_13973,N_13051,N_13121);
nand U13974 (N_13974,N_12807,N_13183);
nand U13975 (N_13975,N_13200,N_13402);
xor U13976 (N_13976,N_12783,N_12807);
nand U13977 (N_13977,N_13187,N_13355);
nand U13978 (N_13978,N_12794,N_13090);
nand U13979 (N_13979,N_12821,N_12870);
nand U13980 (N_13980,N_13300,N_12890);
and U13981 (N_13981,N_13448,N_12933);
nand U13982 (N_13982,N_12882,N_13394);
xor U13983 (N_13983,N_12873,N_12982);
nor U13984 (N_13984,N_13252,N_12759);
xnor U13985 (N_13985,N_13052,N_13308);
nand U13986 (N_13986,N_13190,N_13150);
nor U13987 (N_13987,N_13085,N_12958);
or U13988 (N_13988,N_12942,N_12897);
xnor U13989 (N_13989,N_12960,N_12846);
and U13990 (N_13990,N_13095,N_13033);
xor U13991 (N_13991,N_12949,N_13410);
or U13992 (N_13992,N_12985,N_12785);
nor U13993 (N_13993,N_13412,N_12954);
nand U13994 (N_13994,N_13184,N_12930);
nor U13995 (N_13995,N_13121,N_13377);
and U13996 (N_13996,N_13085,N_13262);
nor U13997 (N_13997,N_12910,N_13468);
xor U13998 (N_13998,N_13258,N_12863);
nor U13999 (N_13999,N_13421,N_12802);
nor U14000 (N_14000,N_12894,N_13479);
nand U14001 (N_14001,N_12821,N_12879);
or U14002 (N_14002,N_12765,N_12865);
or U14003 (N_14003,N_13246,N_12945);
nor U14004 (N_14004,N_12840,N_12911);
nand U14005 (N_14005,N_13290,N_12834);
nand U14006 (N_14006,N_12994,N_13024);
nand U14007 (N_14007,N_12989,N_13384);
xor U14008 (N_14008,N_12958,N_13267);
nor U14009 (N_14009,N_13082,N_13114);
xnor U14010 (N_14010,N_13225,N_13320);
xnor U14011 (N_14011,N_13211,N_13087);
nand U14012 (N_14012,N_13070,N_13114);
nor U14013 (N_14013,N_13244,N_13360);
xor U14014 (N_14014,N_13266,N_12806);
nor U14015 (N_14015,N_12827,N_13087);
or U14016 (N_14016,N_13103,N_13346);
nand U14017 (N_14017,N_13192,N_12833);
and U14018 (N_14018,N_13022,N_13393);
xor U14019 (N_14019,N_12790,N_12927);
and U14020 (N_14020,N_12932,N_12785);
or U14021 (N_14021,N_12789,N_13111);
nor U14022 (N_14022,N_13078,N_13395);
or U14023 (N_14023,N_13188,N_12945);
and U14024 (N_14024,N_12998,N_13394);
xnor U14025 (N_14025,N_13218,N_13261);
nor U14026 (N_14026,N_13379,N_12848);
nand U14027 (N_14027,N_13119,N_12856);
xnor U14028 (N_14028,N_12773,N_13015);
and U14029 (N_14029,N_13249,N_12951);
or U14030 (N_14030,N_13453,N_13413);
nor U14031 (N_14031,N_13041,N_13126);
and U14032 (N_14032,N_13261,N_13289);
and U14033 (N_14033,N_13283,N_13231);
or U14034 (N_14034,N_12841,N_13017);
nand U14035 (N_14035,N_13038,N_13432);
nor U14036 (N_14036,N_12875,N_12934);
or U14037 (N_14037,N_12800,N_12985);
or U14038 (N_14038,N_13132,N_12950);
or U14039 (N_14039,N_13370,N_13404);
or U14040 (N_14040,N_12982,N_12923);
or U14041 (N_14041,N_13340,N_12941);
and U14042 (N_14042,N_13141,N_13085);
and U14043 (N_14043,N_13421,N_13379);
nor U14044 (N_14044,N_13381,N_13214);
nand U14045 (N_14045,N_13051,N_13392);
nand U14046 (N_14046,N_13346,N_12768);
nor U14047 (N_14047,N_12953,N_13102);
xnor U14048 (N_14048,N_13295,N_13250);
or U14049 (N_14049,N_12755,N_13476);
and U14050 (N_14050,N_13029,N_12851);
nor U14051 (N_14051,N_13103,N_12855);
and U14052 (N_14052,N_13025,N_13243);
xnor U14053 (N_14053,N_13127,N_13279);
nor U14054 (N_14054,N_12904,N_13446);
and U14055 (N_14055,N_13357,N_13248);
nor U14056 (N_14056,N_13391,N_13247);
or U14057 (N_14057,N_12979,N_13135);
nor U14058 (N_14058,N_12780,N_13482);
nor U14059 (N_14059,N_13267,N_12979);
and U14060 (N_14060,N_13116,N_13253);
nand U14061 (N_14061,N_13154,N_12856);
xnor U14062 (N_14062,N_13372,N_12919);
and U14063 (N_14063,N_12867,N_13191);
and U14064 (N_14064,N_13472,N_13242);
xnor U14065 (N_14065,N_13065,N_13029);
xnor U14066 (N_14066,N_13360,N_13037);
xor U14067 (N_14067,N_12759,N_13413);
or U14068 (N_14068,N_13212,N_13258);
nand U14069 (N_14069,N_13308,N_12973);
nand U14070 (N_14070,N_13264,N_12855);
nor U14071 (N_14071,N_13483,N_13469);
or U14072 (N_14072,N_13424,N_13449);
and U14073 (N_14073,N_12762,N_13498);
or U14074 (N_14074,N_13145,N_12898);
xor U14075 (N_14075,N_12955,N_13196);
or U14076 (N_14076,N_13170,N_12937);
nor U14077 (N_14077,N_13220,N_13381);
and U14078 (N_14078,N_13386,N_13412);
and U14079 (N_14079,N_13113,N_12778);
nand U14080 (N_14080,N_12981,N_13046);
or U14081 (N_14081,N_13420,N_13242);
and U14082 (N_14082,N_12926,N_13367);
xnor U14083 (N_14083,N_13435,N_13243);
and U14084 (N_14084,N_13082,N_13171);
nor U14085 (N_14085,N_12943,N_13245);
and U14086 (N_14086,N_13310,N_13240);
xor U14087 (N_14087,N_12776,N_12867);
nor U14088 (N_14088,N_13445,N_13285);
or U14089 (N_14089,N_13031,N_13378);
xor U14090 (N_14090,N_12995,N_13003);
xor U14091 (N_14091,N_13143,N_13103);
or U14092 (N_14092,N_12841,N_12923);
nor U14093 (N_14093,N_13358,N_12779);
xnor U14094 (N_14094,N_13410,N_13049);
or U14095 (N_14095,N_13209,N_12898);
or U14096 (N_14096,N_13483,N_13366);
nor U14097 (N_14097,N_12827,N_13041);
xnor U14098 (N_14098,N_13142,N_13372);
nor U14099 (N_14099,N_12984,N_13122);
xor U14100 (N_14100,N_13051,N_13341);
or U14101 (N_14101,N_12931,N_13293);
xnor U14102 (N_14102,N_12939,N_13203);
nand U14103 (N_14103,N_13171,N_13186);
nor U14104 (N_14104,N_13009,N_13019);
xor U14105 (N_14105,N_13432,N_12982);
nand U14106 (N_14106,N_13111,N_12986);
nand U14107 (N_14107,N_12950,N_13345);
nor U14108 (N_14108,N_13336,N_13137);
nand U14109 (N_14109,N_12932,N_12919);
nand U14110 (N_14110,N_13033,N_13207);
nand U14111 (N_14111,N_12882,N_13366);
and U14112 (N_14112,N_12922,N_13080);
nor U14113 (N_14113,N_13367,N_12964);
xnor U14114 (N_14114,N_13313,N_12945);
nor U14115 (N_14115,N_13023,N_13252);
xor U14116 (N_14116,N_12951,N_12784);
or U14117 (N_14117,N_13304,N_12998);
nand U14118 (N_14118,N_12967,N_13371);
nand U14119 (N_14119,N_13023,N_13297);
or U14120 (N_14120,N_13171,N_12878);
nor U14121 (N_14121,N_13366,N_12941);
xor U14122 (N_14122,N_13284,N_13468);
and U14123 (N_14123,N_12853,N_13119);
xnor U14124 (N_14124,N_13407,N_12962);
xnor U14125 (N_14125,N_13082,N_12973);
and U14126 (N_14126,N_13121,N_13228);
or U14127 (N_14127,N_13204,N_13369);
xnor U14128 (N_14128,N_13132,N_13453);
nand U14129 (N_14129,N_13316,N_13389);
nand U14130 (N_14130,N_13028,N_13132);
and U14131 (N_14131,N_13256,N_12813);
or U14132 (N_14132,N_13074,N_13434);
and U14133 (N_14133,N_13156,N_13246);
nor U14134 (N_14134,N_13150,N_13015);
and U14135 (N_14135,N_13318,N_13236);
or U14136 (N_14136,N_13138,N_12750);
nor U14137 (N_14137,N_13193,N_13458);
nor U14138 (N_14138,N_13388,N_13407);
and U14139 (N_14139,N_13023,N_13184);
or U14140 (N_14140,N_13265,N_12882);
xnor U14141 (N_14141,N_12789,N_12937);
nor U14142 (N_14142,N_13439,N_13041);
or U14143 (N_14143,N_13210,N_13179);
or U14144 (N_14144,N_13409,N_13461);
nand U14145 (N_14145,N_13392,N_13189);
and U14146 (N_14146,N_13326,N_13441);
nor U14147 (N_14147,N_13098,N_13420);
nand U14148 (N_14148,N_12897,N_13220);
nor U14149 (N_14149,N_12932,N_13409);
and U14150 (N_14150,N_13351,N_12785);
nor U14151 (N_14151,N_13119,N_13480);
nor U14152 (N_14152,N_13138,N_12831);
or U14153 (N_14153,N_13236,N_13385);
nand U14154 (N_14154,N_13165,N_12988);
nor U14155 (N_14155,N_13194,N_12766);
or U14156 (N_14156,N_13411,N_12809);
nand U14157 (N_14157,N_12912,N_13056);
nor U14158 (N_14158,N_13262,N_13442);
xnor U14159 (N_14159,N_12846,N_12836);
and U14160 (N_14160,N_13239,N_13199);
nor U14161 (N_14161,N_12845,N_13413);
nor U14162 (N_14162,N_13044,N_13181);
xor U14163 (N_14163,N_13167,N_13156);
nand U14164 (N_14164,N_13053,N_12792);
nand U14165 (N_14165,N_13134,N_13444);
and U14166 (N_14166,N_13063,N_13012);
xnor U14167 (N_14167,N_12958,N_13171);
and U14168 (N_14168,N_13024,N_13438);
or U14169 (N_14169,N_13136,N_12946);
nand U14170 (N_14170,N_13099,N_13461);
nand U14171 (N_14171,N_13440,N_13113);
xnor U14172 (N_14172,N_13390,N_13017);
and U14173 (N_14173,N_12983,N_13001);
nor U14174 (N_14174,N_13463,N_13256);
xnor U14175 (N_14175,N_13478,N_13298);
or U14176 (N_14176,N_13237,N_13269);
nor U14177 (N_14177,N_13276,N_13151);
and U14178 (N_14178,N_13069,N_13358);
or U14179 (N_14179,N_13299,N_13108);
or U14180 (N_14180,N_13392,N_12811);
nor U14181 (N_14181,N_12852,N_13444);
and U14182 (N_14182,N_13213,N_13249);
or U14183 (N_14183,N_13327,N_12774);
nor U14184 (N_14184,N_13499,N_12936);
nand U14185 (N_14185,N_12992,N_13047);
xnor U14186 (N_14186,N_12805,N_12796);
or U14187 (N_14187,N_13123,N_13277);
or U14188 (N_14188,N_13379,N_13455);
nand U14189 (N_14189,N_12960,N_13154);
xnor U14190 (N_14190,N_13226,N_13354);
and U14191 (N_14191,N_13264,N_13080);
xnor U14192 (N_14192,N_13388,N_12754);
or U14193 (N_14193,N_13372,N_12975);
or U14194 (N_14194,N_13340,N_12821);
nor U14195 (N_14195,N_12919,N_13479);
xor U14196 (N_14196,N_13288,N_13050);
nor U14197 (N_14197,N_13489,N_12914);
and U14198 (N_14198,N_13182,N_12985);
and U14199 (N_14199,N_13430,N_12987);
or U14200 (N_14200,N_12852,N_12992);
or U14201 (N_14201,N_13110,N_12983);
or U14202 (N_14202,N_12995,N_13414);
nor U14203 (N_14203,N_13471,N_13173);
nand U14204 (N_14204,N_13273,N_12906);
or U14205 (N_14205,N_13099,N_12927);
or U14206 (N_14206,N_13369,N_13005);
xor U14207 (N_14207,N_13271,N_13047);
nor U14208 (N_14208,N_13149,N_13109);
and U14209 (N_14209,N_13125,N_12937);
nor U14210 (N_14210,N_13005,N_13477);
and U14211 (N_14211,N_13004,N_13165);
nand U14212 (N_14212,N_12773,N_13250);
xnor U14213 (N_14213,N_13418,N_13283);
xnor U14214 (N_14214,N_13339,N_12836);
and U14215 (N_14215,N_13205,N_13055);
or U14216 (N_14216,N_13025,N_13338);
xnor U14217 (N_14217,N_13248,N_13155);
or U14218 (N_14218,N_12844,N_13397);
or U14219 (N_14219,N_13080,N_13132);
or U14220 (N_14220,N_13381,N_13421);
nand U14221 (N_14221,N_12821,N_12965);
nor U14222 (N_14222,N_12994,N_13282);
nor U14223 (N_14223,N_13410,N_13472);
xnor U14224 (N_14224,N_13465,N_13227);
or U14225 (N_14225,N_13342,N_12849);
nor U14226 (N_14226,N_13190,N_13329);
and U14227 (N_14227,N_13265,N_12951);
nand U14228 (N_14228,N_13394,N_12849);
nor U14229 (N_14229,N_12893,N_13265);
and U14230 (N_14230,N_12881,N_13033);
or U14231 (N_14231,N_13158,N_13114);
and U14232 (N_14232,N_13442,N_12771);
and U14233 (N_14233,N_13065,N_13035);
and U14234 (N_14234,N_13330,N_13495);
nor U14235 (N_14235,N_12767,N_13061);
nor U14236 (N_14236,N_13376,N_13239);
nor U14237 (N_14237,N_13126,N_13477);
xor U14238 (N_14238,N_12786,N_13042);
nand U14239 (N_14239,N_13403,N_13470);
nand U14240 (N_14240,N_13108,N_13324);
and U14241 (N_14241,N_13140,N_12992);
or U14242 (N_14242,N_13470,N_12889);
and U14243 (N_14243,N_13267,N_13307);
nor U14244 (N_14244,N_13232,N_13247);
and U14245 (N_14245,N_13491,N_13196);
nand U14246 (N_14246,N_13349,N_13284);
nor U14247 (N_14247,N_13368,N_13111);
or U14248 (N_14248,N_13407,N_13367);
nand U14249 (N_14249,N_13486,N_13417);
nand U14250 (N_14250,N_13589,N_13556);
and U14251 (N_14251,N_13529,N_13853);
nor U14252 (N_14252,N_14249,N_14053);
nor U14253 (N_14253,N_13593,N_13646);
or U14254 (N_14254,N_14165,N_13630);
or U14255 (N_14255,N_13877,N_13546);
nor U14256 (N_14256,N_13648,N_14120);
or U14257 (N_14257,N_13692,N_13739);
and U14258 (N_14258,N_13947,N_14154);
nand U14259 (N_14259,N_13520,N_13805);
xnor U14260 (N_14260,N_13974,N_13615);
xor U14261 (N_14261,N_14141,N_13668);
xnor U14262 (N_14262,N_13838,N_13652);
nor U14263 (N_14263,N_13685,N_14086);
or U14264 (N_14264,N_13937,N_13940);
nand U14265 (N_14265,N_13954,N_13898);
or U14266 (N_14266,N_13763,N_13935);
nor U14267 (N_14267,N_13633,N_13899);
or U14268 (N_14268,N_13773,N_14044);
or U14269 (N_14269,N_13582,N_14244);
xnor U14270 (N_14270,N_14189,N_14176);
or U14271 (N_14271,N_13711,N_14240);
nand U14272 (N_14272,N_13799,N_13905);
or U14273 (N_14273,N_13746,N_13665);
xnor U14274 (N_14274,N_13712,N_13851);
nand U14275 (N_14275,N_13531,N_13992);
xor U14276 (N_14276,N_13756,N_13651);
and U14277 (N_14277,N_14020,N_13822);
nand U14278 (N_14278,N_13787,N_13588);
nand U14279 (N_14279,N_13816,N_13536);
nor U14280 (N_14280,N_13620,N_13986);
or U14281 (N_14281,N_13783,N_14047);
or U14282 (N_14282,N_13982,N_13994);
nor U14283 (N_14283,N_14080,N_14190);
or U14284 (N_14284,N_13618,N_13761);
and U14285 (N_14285,N_14200,N_13549);
xnor U14286 (N_14286,N_14220,N_13781);
xnor U14287 (N_14287,N_13628,N_14009);
xor U14288 (N_14288,N_14221,N_13691);
nor U14289 (N_14289,N_14218,N_14081);
and U14290 (N_14290,N_13563,N_13968);
or U14291 (N_14291,N_13721,N_13501);
or U14292 (N_14292,N_13839,N_13797);
and U14293 (N_14293,N_13706,N_14144);
xor U14294 (N_14294,N_14071,N_14056);
or U14295 (N_14295,N_13817,N_14238);
nand U14296 (N_14296,N_13724,N_13865);
nor U14297 (N_14297,N_13580,N_14247);
nand U14298 (N_14298,N_13917,N_14157);
xor U14299 (N_14299,N_13726,N_13671);
or U14300 (N_14300,N_13629,N_13979);
nand U14301 (N_14301,N_13842,N_13846);
nor U14302 (N_14302,N_14094,N_13950);
or U14303 (N_14303,N_13945,N_13507);
or U14304 (N_14304,N_13737,N_14037);
xnor U14305 (N_14305,N_13907,N_13925);
nor U14306 (N_14306,N_14117,N_14112);
and U14307 (N_14307,N_14018,N_13793);
xnor U14308 (N_14308,N_13962,N_14090);
nor U14309 (N_14309,N_14195,N_14214);
nor U14310 (N_14310,N_13570,N_13878);
and U14311 (N_14311,N_13812,N_13991);
or U14312 (N_14312,N_14145,N_14088);
nand U14313 (N_14313,N_14160,N_13894);
or U14314 (N_14314,N_13896,N_14133);
or U14315 (N_14315,N_13682,N_14045);
or U14316 (N_14316,N_13654,N_13697);
nor U14317 (N_14317,N_13873,N_13779);
nor U14318 (N_14318,N_13604,N_13740);
xor U14319 (N_14319,N_14198,N_13802);
nand U14320 (N_14320,N_14215,N_13662);
nand U14321 (N_14321,N_13694,N_13828);
and U14322 (N_14322,N_14073,N_13539);
and U14323 (N_14323,N_13855,N_13999);
xor U14324 (N_14324,N_14107,N_13951);
xor U14325 (N_14325,N_13884,N_13608);
and U14326 (N_14326,N_13576,N_13791);
xor U14327 (N_14327,N_13521,N_13893);
or U14328 (N_14328,N_13619,N_13678);
and U14329 (N_14329,N_14089,N_14017);
xor U14330 (N_14330,N_13681,N_14148);
xnor U14331 (N_14331,N_13923,N_13964);
xor U14332 (N_14332,N_13545,N_14095);
and U14333 (N_14333,N_13577,N_13977);
and U14334 (N_14334,N_13603,N_13769);
or U14335 (N_14335,N_13866,N_14027);
xnor U14336 (N_14336,N_14206,N_13639);
xnor U14337 (N_14337,N_14032,N_14132);
nor U14338 (N_14338,N_14201,N_13742);
nor U14339 (N_14339,N_14004,N_14106);
or U14340 (N_14340,N_14226,N_13760);
xor U14341 (N_14341,N_14139,N_13541);
nand U14342 (N_14342,N_13931,N_13599);
nor U14343 (N_14343,N_14038,N_14219);
or U14344 (N_14344,N_14109,N_14197);
nand U14345 (N_14345,N_13830,N_13581);
xor U14346 (N_14346,N_14022,N_13833);
xor U14347 (N_14347,N_14002,N_13586);
and U14348 (N_14348,N_13774,N_14061);
and U14349 (N_14349,N_13910,N_13792);
and U14350 (N_14350,N_14161,N_14152);
xnor U14351 (N_14351,N_14233,N_13552);
and U14352 (N_14352,N_13789,N_13554);
and U14353 (N_14353,N_13659,N_13672);
nor U14354 (N_14354,N_13882,N_13638);
or U14355 (N_14355,N_14231,N_14057);
and U14356 (N_14356,N_13785,N_13566);
xnor U14357 (N_14357,N_13904,N_13664);
and U14358 (N_14358,N_13673,N_13834);
and U14359 (N_14359,N_13690,N_14102);
nand U14360 (N_14360,N_13730,N_14118);
nor U14361 (N_14361,N_13996,N_13649);
xnor U14362 (N_14362,N_13674,N_14166);
and U14363 (N_14363,N_14125,N_13775);
nor U14364 (N_14364,N_14208,N_14087);
xor U14365 (N_14365,N_13583,N_14051);
nor U14366 (N_14366,N_13868,N_13707);
nor U14367 (N_14367,N_13538,N_13920);
xnor U14368 (N_14368,N_13565,N_13643);
xor U14369 (N_14369,N_13709,N_14043);
nand U14370 (N_14370,N_14021,N_13930);
nor U14371 (N_14371,N_14092,N_13843);
nor U14372 (N_14372,N_14013,N_13891);
nor U14373 (N_14373,N_13537,N_13644);
nor U14374 (N_14374,N_14085,N_14069);
nor U14375 (N_14375,N_13919,N_14025);
xnor U14376 (N_14376,N_13750,N_13729);
and U14377 (N_14377,N_13976,N_13860);
nand U14378 (N_14378,N_13906,N_13625);
xor U14379 (N_14379,N_13605,N_13995);
nor U14380 (N_14380,N_13849,N_13924);
nand U14381 (N_14381,N_13611,N_13575);
nor U14382 (N_14382,N_13578,N_14181);
xor U14383 (N_14383,N_14105,N_13794);
xnor U14384 (N_14384,N_13534,N_14127);
nor U14385 (N_14385,N_13858,N_14093);
and U14386 (N_14386,N_14054,N_13667);
nand U14387 (N_14387,N_13969,N_13523);
nand U14388 (N_14388,N_13510,N_13568);
nand U14389 (N_14389,N_13714,N_14222);
xor U14390 (N_14390,N_13637,N_14033);
and U14391 (N_14391,N_14156,N_13952);
and U14392 (N_14392,N_13768,N_13632);
nand U14393 (N_14393,N_14172,N_14103);
nand U14394 (N_14394,N_13826,N_13998);
nor U14395 (N_14395,N_13759,N_13511);
and U14396 (N_14396,N_13591,N_13861);
nand U14397 (N_14397,N_13824,N_14029);
nor U14398 (N_14398,N_13874,N_13770);
and U14399 (N_14399,N_13972,N_13680);
xnor U14400 (N_14400,N_14178,N_13880);
nor U14401 (N_14401,N_13796,N_13832);
and U14402 (N_14402,N_14224,N_14097);
and U14403 (N_14403,N_13879,N_14163);
or U14404 (N_14404,N_13616,N_13515);
or U14405 (N_14405,N_13686,N_13738);
and U14406 (N_14406,N_13888,N_13548);
or U14407 (N_14407,N_13687,N_14241);
nor U14408 (N_14408,N_14007,N_13550);
nand U14409 (N_14409,N_13985,N_14173);
and U14410 (N_14410,N_13666,N_13889);
nor U14411 (N_14411,N_13704,N_13916);
or U14412 (N_14412,N_13718,N_13745);
nand U14413 (N_14413,N_13530,N_13696);
or U14414 (N_14414,N_14217,N_13850);
nor U14415 (N_14415,N_14041,N_13755);
nand U14416 (N_14416,N_14040,N_14203);
nor U14417 (N_14417,N_14171,N_14065);
nand U14418 (N_14418,N_14075,N_14100);
and U14419 (N_14419,N_14146,N_13614);
and U14420 (N_14420,N_13825,N_13914);
or U14421 (N_14421,N_14034,N_13913);
xor U14422 (N_14422,N_13725,N_13810);
and U14423 (N_14423,N_14049,N_14168);
xor U14424 (N_14424,N_14019,N_13699);
xnor U14425 (N_14425,N_13973,N_13765);
xor U14426 (N_14426,N_13883,N_14121);
nor U14427 (N_14427,N_13512,N_14137);
xor U14428 (N_14428,N_13795,N_14211);
xor U14429 (N_14429,N_13518,N_13572);
nand U14430 (N_14430,N_13934,N_13771);
and U14431 (N_14431,N_13957,N_14234);
nand U14432 (N_14432,N_13663,N_14023);
or U14433 (N_14433,N_14162,N_13587);
and U14434 (N_14434,N_13936,N_13635);
or U14435 (N_14435,N_13598,N_14175);
nand U14436 (N_14436,N_14114,N_13870);
and U14437 (N_14437,N_13609,N_14182);
nor U14438 (N_14438,N_13650,N_13975);
nand U14439 (N_14439,N_13744,N_14243);
xor U14440 (N_14440,N_13553,N_14210);
and U14441 (N_14441,N_13814,N_14016);
nand U14442 (N_14442,N_13528,N_14024);
and U14443 (N_14443,N_13908,N_13821);
nor U14444 (N_14444,N_14153,N_13532);
xor U14445 (N_14445,N_14188,N_13677);
and U14446 (N_14446,N_14180,N_14110);
and U14447 (N_14447,N_13958,N_14111);
or U14448 (N_14448,N_13728,N_13988);
or U14449 (N_14449,N_13540,N_13856);
or U14450 (N_14450,N_13978,N_13844);
or U14451 (N_14451,N_14028,N_14248);
and U14452 (N_14452,N_13815,N_13758);
xnor U14453 (N_14453,N_13655,N_13684);
and U14454 (N_14454,N_13818,N_13869);
xor U14455 (N_14455,N_13875,N_13607);
nand U14456 (N_14456,N_13669,N_13984);
nor U14457 (N_14457,N_14072,N_13987);
xnor U14458 (N_14458,N_13503,N_13679);
or U14459 (N_14459,N_13720,N_13641);
nand U14460 (N_14460,N_14184,N_13804);
xor U14461 (N_14461,N_14213,N_14204);
xor U14462 (N_14462,N_14077,N_14070);
nand U14463 (N_14463,N_14035,N_14209);
nand U14464 (N_14464,N_13803,N_13871);
or U14465 (N_14465,N_13820,N_14128);
and U14466 (N_14466,N_13980,N_13872);
nor U14467 (N_14467,N_14216,N_13636);
and U14468 (N_14468,N_13733,N_13970);
or U14469 (N_14469,N_14067,N_13622);
nor U14470 (N_14470,N_13612,N_14091);
nor U14471 (N_14471,N_13933,N_14048);
or U14472 (N_14472,N_13788,N_14096);
nand U14473 (N_14473,N_14230,N_13848);
nand U14474 (N_14474,N_13993,N_14062);
nor U14475 (N_14475,N_13959,N_13764);
and U14476 (N_14476,N_13956,N_13653);
nor U14477 (N_14477,N_14229,N_13741);
xor U14478 (N_14478,N_13772,N_14126);
xnor U14479 (N_14479,N_14159,N_13514);
and U14480 (N_14480,N_14079,N_14122);
nor U14481 (N_14481,N_14063,N_14113);
and U14482 (N_14482,N_13784,N_13786);
nor U14483 (N_14483,N_13543,N_14151);
xnor U14484 (N_14484,N_13876,N_13617);
nor U14485 (N_14485,N_14140,N_13723);
xnor U14486 (N_14486,N_14012,N_13573);
or U14487 (N_14487,N_13594,N_13701);
or U14488 (N_14488,N_13961,N_13693);
and U14489 (N_14489,N_13929,N_13960);
or U14490 (N_14490,N_13661,N_13544);
or U14491 (N_14491,N_13863,N_13557);
and U14492 (N_14492,N_13912,N_13927);
nand U14493 (N_14493,N_13955,N_13841);
nand U14494 (N_14494,N_13736,N_14169);
xnor U14495 (N_14495,N_14185,N_14119);
nor U14496 (N_14496,N_14036,N_14099);
nor U14497 (N_14497,N_13525,N_13642);
xnor U14498 (N_14498,N_13519,N_13592);
or U14499 (N_14499,N_13658,N_13504);
xnor U14500 (N_14500,N_14135,N_13660);
and U14501 (N_14501,N_13944,N_13997);
or U14502 (N_14502,N_13790,N_13719);
xnor U14503 (N_14503,N_13634,N_14147);
or U14504 (N_14504,N_13555,N_13513);
and U14505 (N_14505,N_13702,N_13941);
xor U14506 (N_14506,N_14246,N_14052);
or U14507 (N_14507,N_13734,N_14026);
nor U14508 (N_14508,N_14031,N_13807);
or U14509 (N_14509,N_14242,N_14078);
and U14510 (N_14510,N_13840,N_14143);
nand U14511 (N_14511,N_14194,N_13610);
xor U14512 (N_14512,N_14011,N_13915);
and U14513 (N_14513,N_13780,N_13502);
xnor U14514 (N_14514,N_13547,N_13752);
or U14515 (N_14515,N_13670,N_14134);
nand U14516 (N_14516,N_13508,N_14101);
and U14517 (N_14517,N_14136,N_14149);
or U14518 (N_14518,N_14177,N_14039);
nor U14519 (N_14519,N_14084,N_14223);
and U14520 (N_14520,N_14138,N_13683);
xor U14521 (N_14521,N_13657,N_13526);
xnor U14522 (N_14522,N_13727,N_13809);
nand U14523 (N_14523,N_14005,N_13762);
nand U14524 (N_14524,N_13800,N_14150);
nand U14525 (N_14525,N_13942,N_14014);
nand U14526 (N_14526,N_14207,N_14164);
nor U14527 (N_14527,N_14142,N_13777);
or U14528 (N_14528,N_13857,N_13946);
nor U14529 (N_14529,N_13798,N_13749);
and U14530 (N_14530,N_13689,N_14124);
xnor U14531 (N_14531,N_13627,N_13886);
nor U14532 (N_14532,N_13903,N_14098);
or U14533 (N_14533,N_13564,N_13897);
xnor U14534 (N_14534,N_13939,N_13808);
and U14535 (N_14535,N_14030,N_13811);
xnor U14536 (N_14536,N_13895,N_13757);
nor U14537 (N_14537,N_13558,N_13722);
and U14538 (N_14538,N_14104,N_13700);
xnor U14539 (N_14539,N_13517,N_13813);
xor U14540 (N_14540,N_13782,N_14170);
or U14541 (N_14541,N_13579,N_14158);
and U14542 (N_14542,N_13778,N_13695);
and U14543 (N_14543,N_14187,N_13922);
and U14544 (N_14544,N_13731,N_14183);
nand U14545 (N_14545,N_13585,N_14193);
nor U14546 (N_14546,N_13836,N_13852);
or U14547 (N_14547,N_13715,N_13989);
and U14548 (N_14548,N_13831,N_13747);
xor U14549 (N_14549,N_13631,N_14155);
or U14550 (N_14550,N_13735,N_13932);
nand U14551 (N_14551,N_13524,N_13595);
xnor U14552 (N_14552,N_14115,N_13823);
or U14553 (N_14553,N_14167,N_14123);
and U14554 (N_14554,N_13854,N_13560);
or U14555 (N_14555,N_13559,N_13901);
nand U14556 (N_14556,N_14227,N_13713);
nand U14557 (N_14557,N_14131,N_13703);
or U14558 (N_14558,N_13569,N_13656);
or U14559 (N_14559,N_13574,N_13881);
nor U14560 (N_14560,N_13647,N_14129);
xor U14561 (N_14561,N_14205,N_14232);
or U14562 (N_14562,N_13835,N_13621);
and U14563 (N_14563,N_13590,N_14074);
nand U14564 (N_14564,N_13767,N_13613);
or U14565 (N_14565,N_14058,N_13890);
or U14566 (N_14566,N_13902,N_14225);
xor U14567 (N_14567,N_13600,N_14108);
and U14568 (N_14568,N_14082,N_13717);
nor U14569 (N_14569,N_13827,N_14006);
xnor U14570 (N_14570,N_13981,N_13748);
xor U14571 (N_14571,N_14059,N_13698);
xor U14572 (N_14572,N_13601,N_13943);
xor U14573 (N_14573,N_13743,N_13516);
nand U14574 (N_14574,N_13626,N_14060);
nor U14575 (N_14575,N_14130,N_13990);
or U14576 (N_14576,N_13710,N_13965);
nand U14577 (N_14577,N_13776,N_14237);
and U14578 (N_14578,N_14003,N_14000);
or U14579 (N_14579,N_13928,N_14046);
nor U14580 (N_14580,N_13819,N_13509);
or U14581 (N_14581,N_13551,N_13754);
nand U14582 (N_14582,N_13926,N_13949);
or U14583 (N_14583,N_13885,N_13829);
and U14584 (N_14584,N_13971,N_14228);
or U14585 (N_14585,N_13602,N_13909);
xnor U14586 (N_14586,N_13561,N_14010);
xor U14587 (N_14587,N_13864,N_13966);
nand U14588 (N_14588,N_13753,N_14015);
or U14589 (N_14589,N_13506,N_13921);
nand U14590 (N_14590,N_14055,N_13751);
xnor U14591 (N_14591,N_13623,N_13953);
and U14592 (N_14592,N_13948,N_14008);
or U14593 (N_14593,N_14236,N_14239);
nor U14594 (N_14594,N_14179,N_13688);
and U14595 (N_14595,N_13967,N_13887);
or U14596 (N_14596,N_13522,N_13535);
xnor U14597 (N_14597,N_14191,N_14196);
nand U14598 (N_14598,N_14076,N_13542);
nand U14599 (N_14599,N_13606,N_13892);
nor U14600 (N_14600,N_14199,N_14116);
nand U14601 (N_14601,N_14083,N_13845);
nand U14602 (N_14602,N_13624,N_13801);
nor U14603 (N_14603,N_14174,N_13918);
xor U14604 (N_14604,N_13640,N_14064);
xnor U14605 (N_14605,N_14186,N_13571);
nor U14606 (N_14606,N_13806,N_13847);
xnor U14607 (N_14607,N_13983,N_13567);
nand U14608 (N_14608,N_13859,N_13963);
or U14609 (N_14609,N_13716,N_13911);
nand U14610 (N_14610,N_14042,N_13732);
xnor U14611 (N_14611,N_13862,N_13584);
and U14612 (N_14612,N_13596,N_13505);
xor U14613 (N_14613,N_13645,N_13837);
xor U14614 (N_14614,N_14245,N_13867);
or U14615 (N_14615,N_13597,N_14066);
or U14616 (N_14616,N_14192,N_13708);
nand U14617 (N_14617,N_14202,N_13527);
and U14618 (N_14618,N_14235,N_13675);
nor U14619 (N_14619,N_13900,N_14212);
nand U14620 (N_14620,N_13533,N_13938);
nand U14621 (N_14621,N_14068,N_13676);
nand U14622 (N_14622,N_14050,N_13562);
nor U14623 (N_14623,N_13705,N_13766);
nand U14624 (N_14624,N_14001,N_13500);
and U14625 (N_14625,N_14151,N_13813);
nand U14626 (N_14626,N_13663,N_13656);
nand U14627 (N_14627,N_13589,N_13967);
nor U14628 (N_14628,N_13550,N_13945);
nand U14629 (N_14629,N_13699,N_14106);
and U14630 (N_14630,N_13520,N_14038);
and U14631 (N_14631,N_14211,N_13757);
nand U14632 (N_14632,N_13800,N_14143);
nand U14633 (N_14633,N_14037,N_13717);
nor U14634 (N_14634,N_13670,N_14138);
nor U14635 (N_14635,N_14219,N_14156);
or U14636 (N_14636,N_13894,N_13520);
nor U14637 (N_14637,N_13578,N_13544);
and U14638 (N_14638,N_13876,N_13535);
and U14639 (N_14639,N_13836,N_14200);
or U14640 (N_14640,N_13799,N_13944);
and U14641 (N_14641,N_13544,N_13692);
and U14642 (N_14642,N_13685,N_13701);
or U14643 (N_14643,N_13771,N_13880);
nor U14644 (N_14644,N_13653,N_13679);
or U14645 (N_14645,N_13648,N_13769);
and U14646 (N_14646,N_13930,N_13992);
or U14647 (N_14647,N_13566,N_14197);
xnor U14648 (N_14648,N_13775,N_14154);
xor U14649 (N_14649,N_13895,N_13731);
or U14650 (N_14650,N_13859,N_13984);
and U14651 (N_14651,N_13805,N_13730);
and U14652 (N_14652,N_13676,N_13773);
nand U14653 (N_14653,N_13562,N_13742);
and U14654 (N_14654,N_14123,N_13807);
or U14655 (N_14655,N_13525,N_13640);
nor U14656 (N_14656,N_14241,N_13534);
nor U14657 (N_14657,N_13909,N_13598);
xnor U14658 (N_14658,N_14081,N_13846);
nand U14659 (N_14659,N_13786,N_14090);
nand U14660 (N_14660,N_13631,N_14247);
and U14661 (N_14661,N_13998,N_13987);
or U14662 (N_14662,N_14092,N_13732);
xor U14663 (N_14663,N_14059,N_13603);
or U14664 (N_14664,N_13547,N_13598);
nor U14665 (N_14665,N_13883,N_13926);
and U14666 (N_14666,N_13755,N_13768);
xor U14667 (N_14667,N_13641,N_13904);
or U14668 (N_14668,N_13702,N_13906);
and U14669 (N_14669,N_14100,N_14145);
or U14670 (N_14670,N_14080,N_14142);
nor U14671 (N_14671,N_13783,N_13680);
and U14672 (N_14672,N_13775,N_13709);
or U14673 (N_14673,N_14196,N_13583);
nor U14674 (N_14674,N_14186,N_13655);
nand U14675 (N_14675,N_13822,N_13576);
xnor U14676 (N_14676,N_13558,N_13562);
nand U14677 (N_14677,N_14040,N_14181);
xnor U14678 (N_14678,N_14049,N_14057);
xnor U14679 (N_14679,N_13833,N_14132);
nand U14680 (N_14680,N_13824,N_13556);
nor U14681 (N_14681,N_14195,N_13951);
xnor U14682 (N_14682,N_13643,N_13713);
or U14683 (N_14683,N_13853,N_14203);
xnor U14684 (N_14684,N_13747,N_13786);
xnor U14685 (N_14685,N_14167,N_13648);
nand U14686 (N_14686,N_13625,N_14070);
nand U14687 (N_14687,N_14141,N_13575);
and U14688 (N_14688,N_14185,N_13933);
xor U14689 (N_14689,N_13951,N_13831);
or U14690 (N_14690,N_14079,N_13847);
nand U14691 (N_14691,N_14240,N_13810);
xor U14692 (N_14692,N_13783,N_13646);
nand U14693 (N_14693,N_13710,N_13585);
and U14694 (N_14694,N_13876,N_13525);
nor U14695 (N_14695,N_13576,N_13896);
xnor U14696 (N_14696,N_13694,N_13913);
or U14697 (N_14697,N_13618,N_13989);
and U14698 (N_14698,N_13703,N_14152);
nand U14699 (N_14699,N_13514,N_14021);
nor U14700 (N_14700,N_13951,N_13587);
nor U14701 (N_14701,N_13865,N_13830);
or U14702 (N_14702,N_14236,N_13725);
and U14703 (N_14703,N_13997,N_14243);
xor U14704 (N_14704,N_13599,N_14100);
nor U14705 (N_14705,N_13691,N_14228);
nand U14706 (N_14706,N_14010,N_13558);
nand U14707 (N_14707,N_13943,N_13834);
or U14708 (N_14708,N_13844,N_13917);
or U14709 (N_14709,N_13548,N_13663);
xor U14710 (N_14710,N_13569,N_13593);
nand U14711 (N_14711,N_14025,N_13851);
xor U14712 (N_14712,N_13809,N_14065);
or U14713 (N_14713,N_13821,N_13638);
and U14714 (N_14714,N_13750,N_14035);
xnor U14715 (N_14715,N_13750,N_13629);
or U14716 (N_14716,N_14249,N_13919);
and U14717 (N_14717,N_13869,N_14048);
or U14718 (N_14718,N_13781,N_14057);
nor U14719 (N_14719,N_13916,N_14228);
and U14720 (N_14720,N_14081,N_13765);
and U14721 (N_14721,N_13728,N_13967);
nor U14722 (N_14722,N_13787,N_13931);
xor U14723 (N_14723,N_13528,N_13878);
nor U14724 (N_14724,N_13952,N_13740);
and U14725 (N_14725,N_14174,N_13983);
nand U14726 (N_14726,N_13665,N_13726);
and U14727 (N_14727,N_13575,N_13998);
or U14728 (N_14728,N_13987,N_13515);
xor U14729 (N_14729,N_13792,N_13884);
and U14730 (N_14730,N_13904,N_13905);
nor U14731 (N_14731,N_14068,N_13708);
or U14732 (N_14732,N_13868,N_14151);
nor U14733 (N_14733,N_13862,N_13953);
xnor U14734 (N_14734,N_13949,N_13631);
and U14735 (N_14735,N_13581,N_13867);
and U14736 (N_14736,N_13839,N_14121);
and U14737 (N_14737,N_14176,N_14016);
nor U14738 (N_14738,N_13925,N_13944);
nor U14739 (N_14739,N_14108,N_14186);
or U14740 (N_14740,N_13843,N_14025);
or U14741 (N_14741,N_14086,N_13623);
nand U14742 (N_14742,N_14168,N_14023);
xor U14743 (N_14743,N_13681,N_13647);
nand U14744 (N_14744,N_13779,N_13678);
nand U14745 (N_14745,N_14218,N_14133);
nor U14746 (N_14746,N_14176,N_14135);
or U14747 (N_14747,N_13674,N_13559);
nand U14748 (N_14748,N_14223,N_14145);
or U14749 (N_14749,N_13525,N_13893);
and U14750 (N_14750,N_13555,N_13761);
xnor U14751 (N_14751,N_14247,N_13918);
or U14752 (N_14752,N_13766,N_13724);
and U14753 (N_14753,N_13821,N_13997);
nand U14754 (N_14754,N_13860,N_13573);
nor U14755 (N_14755,N_13968,N_14206);
xnor U14756 (N_14756,N_13910,N_14136);
or U14757 (N_14757,N_13671,N_13670);
xnor U14758 (N_14758,N_13520,N_13932);
or U14759 (N_14759,N_13706,N_14022);
or U14760 (N_14760,N_14195,N_14207);
and U14761 (N_14761,N_13515,N_13624);
nor U14762 (N_14762,N_13575,N_13768);
nor U14763 (N_14763,N_13991,N_13716);
nor U14764 (N_14764,N_13596,N_14131);
nor U14765 (N_14765,N_13692,N_14058);
or U14766 (N_14766,N_14222,N_13645);
and U14767 (N_14767,N_13805,N_13600);
and U14768 (N_14768,N_13931,N_13679);
xor U14769 (N_14769,N_13859,N_14075);
xor U14770 (N_14770,N_13668,N_14236);
xor U14771 (N_14771,N_13740,N_14049);
nand U14772 (N_14772,N_13754,N_14190);
and U14773 (N_14773,N_13547,N_13729);
nor U14774 (N_14774,N_13745,N_13764);
and U14775 (N_14775,N_14186,N_13863);
nor U14776 (N_14776,N_13661,N_13872);
nand U14777 (N_14777,N_14004,N_13842);
nor U14778 (N_14778,N_13550,N_13764);
xnor U14779 (N_14779,N_13651,N_13677);
xor U14780 (N_14780,N_13548,N_13752);
nand U14781 (N_14781,N_13909,N_13860);
and U14782 (N_14782,N_14096,N_14224);
xnor U14783 (N_14783,N_14095,N_13658);
nand U14784 (N_14784,N_14239,N_14174);
or U14785 (N_14785,N_13749,N_13672);
xor U14786 (N_14786,N_13960,N_13890);
and U14787 (N_14787,N_13567,N_13669);
nand U14788 (N_14788,N_13809,N_13673);
nor U14789 (N_14789,N_13743,N_14055);
or U14790 (N_14790,N_14125,N_13545);
and U14791 (N_14791,N_13869,N_13734);
and U14792 (N_14792,N_13891,N_14042);
and U14793 (N_14793,N_13788,N_13615);
or U14794 (N_14794,N_14007,N_14207);
nor U14795 (N_14795,N_13515,N_13775);
nand U14796 (N_14796,N_14043,N_14208);
nor U14797 (N_14797,N_13902,N_13864);
or U14798 (N_14798,N_13650,N_14161);
nor U14799 (N_14799,N_14163,N_14094);
xor U14800 (N_14800,N_13667,N_13615);
xnor U14801 (N_14801,N_13900,N_13707);
nor U14802 (N_14802,N_13920,N_14051);
and U14803 (N_14803,N_14162,N_14175);
nand U14804 (N_14804,N_14083,N_13851);
nand U14805 (N_14805,N_13557,N_13693);
xor U14806 (N_14806,N_14211,N_13614);
xnor U14807 (N_14807,N_13959,N_14215);
nand U14808 (N_14808,N_14014,N_13614);
xnor U14809 (N_14809,N_14186,N_13951);
nor U14810 (N_14810,N_14213,N_13722);
nor U14811 (N_14811,N_13564,N_14124);
nand U14812 (N_14812,N_14042,N_14166);
or U14813 (N_14813,N_13962,N_13868);
nand U14814 (N_14814,N_13821,N_14063);
xnor U14815 (N_14815,N_13525,N_13715);
nand U14816 (N_14816,N_13755,N_13546);
nand U14817 (N_14817,N_13883,N_13837);
and U14818 (N_14818,N_13811,N_14198);
and U14819 (N_14819,N_14169,N_13650);
nand U14820 (N_14820,N_13548,N_14102);
and U14821 (N_14821,N_13724,N_13984);
or U14822 (N_14822,N_14162,N_13734);
and U14823 (N_14823,N_13701,N_14034);
and U14824 (N_14824,N_14049,N_13968);
nor U14825 (N_14825,N_14021,N_14010);
xnor U14826 (N_14826,N_13863,N_13601);
nand U14827 (N_14827,N_13619,N_13524);
xnor U14828 (N_14828,N_13659,N_13588);
and U14829 (N_14829,N_14173,N_13741);
or U14830 (N_14830,N_13692,N_13600);
and U14831 (N_14831,N_13950,N_13777);
nand U14832 (N_14832,N_13535,N_13527);
or U14833 (N_14833,N_13692,N_13837);
and U14834 (N_14834,N_14247,N_13827);
nor U14835 (N_14835,N_13683,N_13743);
and U14836 (N_14836,N_13538,N_14096);
nand U14837 (N_14837,N_13933,N_14098);
or U14838 (N_14838,N_14148,N_13685);
nor U14839 (N_14839,N_14154,N_13716);
or U14840 (N_14840,N_14086,N_14136);
or U14841 (N_14841,N_13611,N_14071);
nand U14842 (N_14842,N_13899,N_13536);
xnor U14843 (N_14843,N_14126,N_13598);
and U14844 (N_14844,N_14034,N_13580);
or U14845 (N_14845,N_13518,N_13530);
and U14846 (N_14846,N_14082,N_13757);
and U14847 (N_14847,N_13708,N_14036);
and U14848 (N_14848,N_14203,N_14194);
and U14849 (N_14849,N_13756,N_14137);
and U14850 (N_14850,N_13723,N_13933);
and U14851 (N_14851,N_14090,N_13903);
xor U14852 (N_14852,N_14029,N_13599);
nor U14853 (N_14853,N_13897,N_13905);
nor U14854 (N_14854,N_13635,N_13549);
nand U14855 (N_14855,N_13734,N_13669);
and U14856 (N_14856,N_13719,N_13835);
xnor U14857 (N_14857,N_13552,N_13622);
xor U14858 (N_14858,N_13514,N_14033);
or U14859 (N_14859,N_13900,N_13771);
nor U14860 (N_14860,N_13849,N_14138);
xor U14861 (N_14861,N_13640,N_13710);
nand U14862 (N_14862,N_14170,N_13608);
xnor U14863 (N_14863,N_14224,N_14028);
and U14864 (N_14864,N_13847,N_13752);
nor U14865 (N_14865,N_14222,N_14062);
xor U14866 (N_14866,N_14241,N_14225);
xor U14867 (N_14867,N_13820,N_13525);
nor U14868 (N_14868,N_13500,N_13716);
or U14869 (N_14869,N_13871,N_13737);
nor U14870 (N_14870,N_13929,N_14215);
nor U14871 (N_14871,N_14012,N_13571);
and U14872 (N_14872,N_13791,N_13897);
xnor U14873 (N_14873,N_14202,N_14136);
or U14874 (N_14874,N_13946,N_13959);
or U14875 (N_14875,N_13692,N_14077);
xnor U14876 (N_14876,N_13616,N_13760);
xnor U14877 (N_14877,N_14029,N_13820);
and U14878 (N_14878,N_14212,N_13628);
and U14879 (N_14879,N_13945,N_13525);
nor U14880 (N_14880,N_13668,N_13925);
nor U14881 (N_14881,N_13840,N_13666);
or U14882 (N_14882,N_13691,N_13647);
or U14883 (N_14883,N_13552,N_13937);
nor U14884 (N_14884,N_13920,N_14209);
nand U14885 (N_14885,N_13718,N_13638);
and U14886 (N_14886,N_14161,N_14147);
and U14887 (N_14887,N_13717,N_13925);
xor U14888 (N_14888,N_13503,N_13804);
nand U14889 (N_14889,N_13737,N_13907);
nor U14890 (N_14890,N_13627,N_13588);
and U14891 (N_14891,N_14064,N_13945);
and U14892 (N_14892,N_14007,N_13690);
and U14893 (N_14893,N_13953,N_13636);
nand U14894 (N_14894,N_13885,N_13699);
or U14895 (N_14895,N_13628,N_14176);
nor U14896 (N_14896,N_13701,N_13606);
and U14897 (N_14897,N_13789,N_13607);
nor U14898 (N_14898,N_14064,N_13705);
nor U14899 (N_14899,N_13628,N_14069);
nand U14900 (N_14900,N_14137,N_13762);
nand U14901 (N_14901,N_14146,N_13754);
and U14902 (N_14902,N_13861,N_13659);
nand U14903 (N_14903,N_14229,N_13929);
nand U14904 (N_14904,N_14055,N_13807);
nand U14905 (N_14905,N_13819,N_13935);
xor U14906 (N_14906,N_14007,N_14147);
and U14907 (N_14907,N_14189,N_13784);
or U14908 (N_14908,N_13993,N_14020);
xnor U14909 (N_14909,N_13878,N_13573);
nand U14910 (N_14910,N_14080,N_13681);
or U14911 (N_14911,N_14101,N_14044);
nand U14912 (N_14912,N_13639,N_13673);
nor U14913 (N_14913,N_13707,N_14201);
xnor U14914 (N_14914,N_14068,N_14232);
nand U14915 (N_14915,N_13746,N_13541);
or U14916 (N_14916,N_14025,N_14249);
or U14917 (N_14917,N_13588,N_14139);
nor U14918 (N_14918,N_13779,N_13925);
nand U14919 (N_14919,N_13600,N_14048);
xnor U14920 (N_14920,N_14127,N_13895);
xor U14921 (N_14921,N_13575,N_13779);
xnor U14922 (N_14922,N_14018,N_13900);
xor U14923 (N_14923,N_13870,N_13999);
nor U14924 (N_14924,N_14167,N_14113);
or U14925 (N_14925,N_13977,N_14060);
xor U14926 (N_14926,N_14037,N_13643);
or U14927 (N_14927,N_13526,N_13858);
nand U14928 (N_14928,N_13856,N_13957);
nand U14929 (N_14929,N_13658,N_14164);
xnor U14930 (N_14930,N_14095,N_13829);
or U14931 (N_14931,N_13996,N_14067);
nand U14932 (N_14932,N_13583,N_13503);
nor U14933 (N_14933,N_13539,N_13646);
and U14934 (N_14934,N_14003,N_13670);
nor U14935 (N_14935,N_13720,N_14154);
nand U14936 (N_14936,N_13771,N_13857);
xor U14937 (N_14937,N_13898,N_13644);
nor U14938 (N_14938,N_14015,N_13594);
xor U14939 (N_14939,N_13587,N_14164);
and U14940 (N_14940,N_13521,N_13908);
xnor U14941 (N_14941,N_13920,N_13759);
xnor U14942 (N_14942,N_14079,N_13946);
nand U14943 (N_14943,N_13989,N_13949);
and U14944 (N_14944,N_14082,N_13820);
nor U14945 (N_14945,N_13857,N_13671);
nor U14946 (N_14946,N_14160,N_13556);
and U14947 (N_14947,N_14240,N_13671);
or U14948 (N_14948,N_14002,N_13511);
or U14949 (N_14949,N_14096,N_13938);
nor U14950 (N_14950,N_14212,N_14149);
nand U14951 (N_14951,N_13688,N_13834);
and U14952 (N_14952,N_14098,N_14050);
and U14953 (N_14953,N_14199,N_13765);
or U14954 (N_14954,N_13975,N_14043);
nor U14955 (N_14955,N_13701,N_13714);
nand U14956 (N_14956,N_13724,N_13873);
or U14957 (N_14957,N_14159,N_13507);
xnor U14958 (N_14958,N_14010,N_14209);
xnor U14959 (N_14959,N_13740,N_13798);
nand U14960 (N_14960,N_13859,N_13784);
xor U14961 (N_14961,N_13519,N_13522);
xnor U14962 (N_14962,N_13948,N_13823);
nor U14963 (N_14963,N_13529,N_13632);
and U14964 (N_14964,N_13831,N_14097);
or U14965 (N_14965,N_13856,N_13672);
nand U14966 (N_14966,N_13793,N_14083);
and U14967 (N_14967,N_13706,N_13558);
and U14968 (N_14968,N_14087,N_14038);
or U14969 (N_14969,N_13712,N_14018);
or U14970 (N_14970,N_13887,N_14206);
xor U14971 (N_14971,N_13672,N_13836);
nor U14972 (N_14972,N_13636,N_14077);
nor U14973 (N_14973,N_14218,N_13621);
xnor U14974 (N_14974,N_14099,N_13511);
nor U14975 (N_14975,N_13628,N_13583);
xor U14976 (N_14976,N_13980,N_14203);
nor U14977 (N_14977,N_13790,N_14008);
nor U14978 (N_14978,N_13641,N_13737);
xnor U14979 (N_14979,N_14041,N_14023);
xor U14980 (N_14980,N_14150,N_13539);
nand U14981 (N_14981,N_14151,N_13619);
and U14982 (N_14982,N_13721,N_13682);
and U14983 (N_14983,N_13519,N_13591);
nor U14984 (N_14984,N_13970,N_13832);
or U14985 (N_14985,N_13833,N_13742);
nor U14986 (N_14986,N_13638,N_14043);
xor U14987 (N_14987,N_14167,N_13825);
nor U14988 (N_14988,N_14108,N_14147);
nand U14989 (N_14989,N_13744,N_13659);
nor U14990 (N_14990,N_14128,N_13847);
or U14991 (N_14991,N_14241,N_13785);
nor U14992 (N_14992,N_14180,N_13615);
nor U14993 (N_14993,N_13887,N_13635);
xor U14994 (N_14994,N_14239,N_14074);
xor U14995 (N_14995,N_13516,N_13916);
xor U14996 (N_14996,N_13778,N_13682);
nor U14997 (N_14997,N_14144,N_14074);
nor U14998 (N_14998,N_14074,N_13761);
xor U14999 (N_14999,N_13592,N_13531);
nor UO_0 (O_0,N_14279,N_14564);
or UO_1 (O_1,N_14401,N_14324);
nand UO_2 (O_2,N_14256,N_14616);
xor UO_3 (O_3,N_14838,N_14635);
nor UO_4 (O_4,N_14299,N_14847);
nor UO_5 (O_5,N_14553,N_14826);
or UO_6 (O_6,N_14339,N_14284);
or UO_7 (O_7,N_14948,N_14760);
or UO_8 (O_8,N_14493,N_14746);
and UO_9 (O_9,N_14983,N_14541);
nor UO_10 (O_10,N_14506,N_14957);
nor UO_11 (O_11,N_14766,N_14531);
xor UO_12 (O_12,N_14570,N_14621);
and UO_13 (O_13,N_14503,N_14919);
nor UO_14 (O_14,N_14835,N_14703);
nand UO_15 (O_15,N_14912,N_14998);
xnor UO_16 (O_16,N_14972,N_14750);
nand UO_17 (O_17,N_14426,N_14909);
and UO_18 (O_18,N_14813,N_14894);
xor UO_19 (O_19,N_14716,N_14945);
xor UO_20 (O_20,N_14803,N_14368);
xor UO_21 (O_21,N_14706,N_14617);
nor UO_22 (O_22,N_14574,N_14890);
nand UO_23 (O_23,N_14868,N_14512);
nand UO_24 (O_24,N_14968,N_14694);
and UO_25 (O_25,N_14923,N_14304);
and UO_26 (O_26,N_14888,N_14851);
and UO_27 (O_27,N_14350,N_14821);
or UO_28 (O_28,N_14772,N_14395);
nand UO_29 (O_29,N_14657,N_14548);
xnor UO_30 (O_30,N_14474,N_14642);
and UO_31 (O_31,N_14610,N_14402);
or UO_32 (O_32,N_14454,N_14818);
or UO_33 (O_33,N_14475,N_14761);
and UO_34 (O_34,N_14799,N_14332);
nor UO_35 (O_35,N_14549,N_14556);
nor UO_36 (O_36,N_14509,N_14544);
or UO_37 (O_37,N_14595,N_14592);
nand UO_38 (O_38,N_14916,N_14640);
and UO_39 (O_39,N_14251,N_14295);
nand UO_40 (O_40,N_14480,N_14960);
nand UO_41 (O_41,N_14568,N_14529);
nor UO_42 (O_42,N_14313,N_14423);
or UO_43 (O_43,N_14398,N_14977);
nand UO_44 (O_44,N_14921,N_14864);
nor UO_45 (O_45,N_14685,N_14687);
nor UO_46 (O_46,N_14523,N_14354);
nand UO_47 (O_47,N_14320,N_14507);
and UO_48 (O_48,N_14975,N_14442);
nand UO_49 (O_49,N_14405,N_14889);
or UO_50 (O_50,N_14290,N_14824);
xnor UO_51 (O_51,N_14499,N_14725);
nor UO_52 (O_52,N_14976,N_14798);
xnor UO_53 (O_53,N_14433,N_14335);
or UO_54 (O_54,N_14802,N_14591);
xnor UO_55 (O_55,N_14770,N_14298);
xor UO_56 (O_56,N_14626,N_14702);
xnor UO_57 (O_57,N_14740,N_14837);
nand UO_58 (O_58,N_14486,N_14554);
xnor UO_59 (O_59,N_14448,N_14947);
or UO_60 (O_60,N_14559,N_14488);
or UO_61 (O_61,N_14361,N_14757);
nor UO_62 (O_62,N_14422,N_14876);
xnor UO_63 (O_63,N_14863,N_14323);
xnor UO_64 (O_64,N_14494,N_14404);
and UO_65 (O_65,N_14632,N_14815);
and UO_66 (O_66,N_14811,N_14849);
or UO_67 (O_67,N_14788,N_14843);
and UO_68 (O_68,N_14628,N_14904);
nor UO_69 (O_69,N_14833,N_14711);
nand UO_70 (O_70,N_14928,N_14668);
and UO_71 (O_71,N_14828,N_14981);
nor UO_72 (O_72,N_14563,N_14428);
or UO_73 (O_73,N_14884,N_14963);
nor UO_74 (O_74,N_14751,N_14259);
nand UO_75 (O_75,N_14705,N_14790);
nand UO_76 (O_76,N_14593,N_14273);
nor UO_77 (O_77,N_14765,N_14333);
nand UO_78 (O_78,N_14520,N_14974);
or UO_79 (O_79,N_14715,N_14425);
nor UO_80 (O_80,N_14390,N_14801);
nor UO_81 (O_81,N_14791,N_14834);
nor UO_82 (O_82,N_14809,N_14779);
or UO_83 (O_83,N_14625,N_14599);
xor UO_84 (O_84,N_14663,N_14911);
xor UO_85 (O_85,N_14275,N_14491);
or UO_86 (O_86,N_14573,N_14728);
nor UO_87 (O_87,N_14622,N_14690);
xnor UO_88 (O_88,N_14858,N_14495);
and UO_89 (O_89,N_14996,N_14662);
xor UO_90 (O_90,N_14631,N_14340);
or UO_91 (O_91,N_14403,N_14346);
xor UO_92 (O_92,N_14437,N_14759);
nand UO_93 (O_93,N_14973,N_14862);
or UO_94 (O_94,N_14464,N_14933);
and UO_95 (O_95,N_14504,N_14534);
xnor UO_96 (O_96,N_14545,N_14487);
nand UO_97 (O_97,N_14387,N_14327);
and UO_98 (O_98,N_14682,N_14731);
nand UO_99 (O_99,N_14345,N_14754);
xnor UO_100 (O_100,N_14508,N_14807);
nor UO_101 (O_101,N_14250,N_14653);
or UO_102 (O_102,N_14878,N_14594);
nand UO_103 (O_103,N_14936,N_14265);
or UO_104 (O_104,N_14887,N_14476);
xnor UO_105 (O_105,N_14907,N_14565);
xnor UO_106 (O_106,N_14608,N_14695);
nand UO_107 (O_107,N_14900,N_14634);
nor UO_108 (O_108,N_14899,N_14949);
or UO_109 (O_109,N_14436,N_14962);
or UO_110 (O_110,N_14872,N_14458);
xor UO_111 (O_111,N_14661,N_14829);
nor UO_112 (O_112,N_14510,N_14885);
nor UO_113 (O_113,N_14710,N_14886);
nor UO_114 (O_114,N_14649,N_14836);
nor UO_115 (O_115,N_14659,N_14850);
and UO_116 (O_116,N_14421,N_14260);
nand UO_117 (O_117,N_14481,N_14932);
or UO_118 (O_118,N_14674,N_14753);
or UO_119 (O_119,N_14411,N_14471);
nand UO_120 (O_120,N_14418,N_14432);
xor UO_121 (O_121,N_14264,N_14364);
and UO_122 (O_122,N_14302,N_14586);
and UO_123 (O_123,N_14334,N_14860);
nand UO_124 (O_124,N_14789,N_14756);
xnor UO_125 (O_125,N_14514,N_14784);
and UO_126 (O_126,N_14924,N_14712);
nor UO_127 (O_127,N_14796,N_14492);
nor UO_128 (O_128,N_14656,N_14462);
nand UO_129 (O_129,N_14280,N_14539);
and UO_130 (O_130,N_14980,N_14739);
and UO_131 (O_131,N_14646,N_14285);
xor UO_132 (O_132,N_14995,N_14413);
nor UO_133 (O_133,N_14999,N_14956);
nand UO_134 (O_134,N_14954,N_14741);
and UO_135 (O_135,N_14365,N_14312);
and UO_136 (O_136,N_14588,N_14777);
and UO_137 (O_137,N_14352,N_14992);
and UO_138 (O_138,N_14579,N_14859);
nor UO_139 (O_139,N_14839,N_14871);
nor UO_140 (O_140,N_14543,N_14420);
and UO_141 (O_141,N_14666,N_14737);
and UO_142 (O_142,N_14607,N_14611);
or UO_143 (O_143,N_14502,N_14764);
or UO_144 (O_144,N_14315,N_14329);
nor UO_145 (O_145,N_14678,N_14827);
xnor UO_146 (O_146,N_14853,N_14966);
and UO_147 (O_147,N_14767,N_14935);
or UO_148 (O_148,N_14252,N_14517);
xnor UO_149 (O_149,N_14465,N_14638);
or UO_150 (O_150,N_14450,N_14726);
nand UO_151 (O_151,N_14736,N_14268);
or UO_152 (O_152,N_14337,N_14931);
nor UO_153 (O_153,N_14381,N_14944);
and UO_154 (O_154,N_14699,N_14449);
nor UO_155 (O_155,N_14673,N_14624);
xnor UO_156 (O_156,N_14958,N_14644);
xor UO_157 (O_157,N_14892,N_14806);
xnor UO_158 (O_158,N_14865,N_14768);
nand UO_159 (O_159,N_14842,N_14709);
xnor UO_160 (O_160,N_14536,N_14555);
or UO_161 (O_161,N_14910,N_14776);
nor UO_162 (O_162,N_14769,N_14330);
nand UO_163 (O_163,N_14717,N_14881);
and UO_164 (O_164,N_14344,N_14456);
and UO_165 (O_165,N_14987,N_14704);
or UO_166 (O_166,N_14620,N_14321);
nor UO_167 (O_167,N_14747,N_14639);
or UO_168 (O_168,N_14578,N_14990);
nor UO_169 (O_169,N_14901,N_14669);
and UO_170 (O_170,N_14670,N_14526);
or UO_171 (O_171,N_14971,N_14469);
xnor UO_172 (O_172,N_14457,N_14915);
xnor UO_173 (O_173,N_14654,N_14979);
nand UO_174 (O_174,N_14558,N_14742);
nor UO_175 (O_175,N_14794,N_14735);
nand UO_176 (O_176,N_14922,N_14431);
nand UO_177 (O_177,N_14351,N_14501);
nand UO_178 (O_178,N_14580,N_14723);
xor UO_179 (O_179,N_14918,N_14920);
nor UO_180 (O_180,N_14688,N_14874);
or UO_181 (O_181,N_14841,N_14267);
or UO_182 (O_182,N_14745,N_14478);
or UO_183 (O_183,N_14326,N_14623);
nand UO_184 (O_184,N_14961,N_14946);
nand UO_185 (O_185,N_14293,N_14263);
and UO_186 (O_186,N_14410,N_14619);
and UO_187 (O_187,N_14696,N_14883);
or UO_188 (O_188,N_14289,N_14810);
nor UO_189 (O_189,N_14793,N_14743);
or UO_190 (O_190,N_14400,N_14902);
xor UO_191 (O_191,N_14366,N_14399);
xor UO_192 (O_192,N_14521,N_14590);
or UO_193 (O_193,N_14939,N_14376);
or UO_194 (O_194,N_14665,N_14445);
nor UO_195 (O_195,N_14693,N_14880);
nor UO_196 (O_196,N_14409,N_14375);
nor UO_197 (O_197,N_14775,N_14819);
nand UO_198 (O_198,N_14540,N_14371);
and UO_199 (O_199,N_14466,N_14749);
and UO_200 (O_200,N_14562,N_14671);
nand UO_201 (O_201,N_14468,N_14278);
nand UO_202 (O_202,N_14359,N_14530);
and UO_203 (O_203,N_14524,N_14407);
nor UO_204 (O_204,N_14396,N_14986);
and UO_205 (O_205,N_14331,N_14356);
xnor UO_206 (O_206,N_14752,N_14385);
nor UO_207 (O_207,N_14598,N_14882);
and UO_208 (O_208,N_14701,N_14451);
nand UO_209 (O_209,N_14367,N_14758);
nor UO_210 (O_210,N_14729,N_14338);
and UO_211 (O_211,N_14780,N_14276);
or UO_212 (O_212,N_14681,N_14831);
nand UO_213 (O_213,N_14783,N_14261);
nor UO_214 (O_214,N_14773,N_14692);
nand UO_215 (O_215,N_14470,N_14732);
nor UO_216 (O_216,N_14734,N_14720);
nor UO_217 (O_217,N_14898,N_14342);
and UO_218 (O_218,N_14341,N_14569);
nand UO_219 (O_219,N_14389,N_14870);
nor UO_220 (O_220,N_14316,N_14282);
and UO_221 (O_221,N_14730,N_14585);
and UO_222 (O_222,N_14257,N_14527);
or UO_223 (O_223,N_14353,N_14377);
or UO_224 (O_224,N_14877,N_14292);
nor UO_225 (O_225,N_14463,N_14676);
nand UO_226 (O_226,N_14613,N_14417);
and UO_227 (O_227,N_14597,N_14605);
xnor UO_228 (O_228,N_14840,N_14797);
nor UO_229 (O_229,N_14270,N_14427);
or UO_230 (O_230,N_14441,N_14606);
xor UO_231 (O_231,N_14484,N_14473);
xnor UO_232 (O_232,N_14472,N_14255);
nand UO_233 (O_233,N_14258,N_14869);
or UO_234 (O_234,N_14373,N_14680);
nor UO_235 (O_235,N_14805,N_14357);
nand UO_236 (O_236,N_14721,N_14844);
or UO_237 (O_237,N_14926,N_14406);
and UO_238 (O_238,N_14288,N_14698);
nor UO_239 (O_239,N_14627,N_14648);
xnor UO_240 (O_240,N_14479,N_14397);
nor UO_241 (O_241,N_14713,N_14652);
xor UO_242 (O_242,N_14482,N_14286);
and UO_243 (O_243,N_14897,N_14609);
or UO_244 (O_244,N_14893,N_14913);
nor UO_245 (O_245,N_14380,N_14347);
nor UO_246 (O_246,N_14601,N_14550);
xnor UO_247 (O_247,N_14719,N_14615);
xnor UO_248 (O_248,N_14414,N_14408);
xnor UO_249 (O_249,N_14424,N_14384);
xor UO_250 (O_250,N_14496,N_14658);
xor UO_251 (O_251,N_14308,N_14305);
nor UO_252 (O_252,N_14991,N_14439);
nand UO_253 (O_253,N_14274,N_14328);
or UO_254 (O_254,N_14301,N_14489);
and UO_255 (O_255,N_14978,N_14643);
and UO_256 (O_256,N_14786,N_14997);
nor UO_257 (O_257,N_14823,N_14895);
or UO_258 (O_258,N_14287,N_14792);
or UO_259 (O_259,N_14440,N_14820);
nor UO_260 (O_260,N_14655,N_14513);
nor UO_261 (O_261,N_14938,N_14867);
or UO_262 (O_262,N_14814,N_14697);
nor UO_263 (O_263,N_14969,N_14435);
and UO_264 (O_264,N_14708,N_14903);
nand UO_265 (O_265,N_14891,N_14300);
nand UO_266 (O_266,N_14383,N_14447);
nor UO_267 (O_267,N_14774,N_14722);
xnor UO_268 (O_268,N_14355,N_14630);
nand UO_269 (O_269,N_14873,N_14965);
and UO_270 (O_270,N_14645,N_14388);
nand UO_271 (O_271,N_14984,N_14429);
nand UO_272 (O_272,N_14576,N_14684);
nand UO_273 (O_273,N_14412,N_14379);
nor UO_274 (O_274,N_14358,N_14664);
xor UO_275 (O_275,N_14677,N_14994);
xor UO_276 (O_276,N_14940,N_14641);
or UO_277 (O_277,N_14636,N_14434);
nor UO_278 (O_278,N_14755,N_14319);
or UO_279 (O_279,N_14277,N_14430);
nor UO_280 (O_280,N_14532,N_14362);
or UO_281 (O_281,N_14557,N_14309);
or UO_282 (O_282,N_14370,N_14392);
nor UO_283 (O_283,N_14498,N_14336);
nor UO_284 (O_284,N_14505,N_14718);
or UO_285 (O_285,N_14941,N_14571);
nor UO_286 (O_286,N_14587,N_14683);
and UO_287 (O_287,N_14518,N_14461);
nor UO_288 (O_288,N_14296,N_14629);
xnor UO_289 (O_289,N_14438,N_14360);
nor UO_290 (O_290,N_14515,N_14855);
nand UO_291 (O_291,N_14959,N_14262);
or UO_292 (O_292,N_14294,N_14575);
nand UO_293 (O_293,N_14929,N_14378);
and UO_294 (O_294,N_14459,N_14857);
and UO_295 (O_295,N_14650,N_14297);
xor UO_296 (O_296,N_14804,N_14700);
or UO_297 (O_297,N_14393,N_14846);
nor UO_298 (O_298,N_14283,N_14455);
or UO_299 (O_299,N_14989,N_14386);
xor UO_300 (O_300,N_14581,N_14953);
or UO_301 (O_301,N_14583,N_14394);
and UO_302 (O_302,N_14970,N_14943);
nand UO_303 (O_303,N_14917,N_14667);
and UO_304 (O_304,N_14795,N_14614);
or UO_305 (O_305,N_14542,N_14374);
or UO_306 (O_306,N_14930,N_14651);
nor UO_307 (O_307,N_14985,N_14785);
nor UO_308 (O_308,N_14446,N_14602);
xnor UO_309 (O_309,N_14689,N_14444);
and UO_310 (O_310,N_14781,N_14546);
nor UO_311 (O_311,N_14925,N_14908);
and UO_312 (O_312,N_14567,N_14763);
and UO_313 (O_313,N_14861,N_14419);
nand UO_314 (O_314,N_14460,N_14577);
and UO_315 (O_315,N_14253,N_14522);
or UO_316 (O_316,N_14618,N_14993);
xnor UO_317 (O_317,N_14483,N_14955);
nand UO_318 (O_318,N_14875,N_14516);
nand UO_319 (O_319,N_14317,N_14830);
nor UO_320 (O_320,N_14937,N_14714);
or UO_321 (O_321,N_14848,N_14727);
or UO_322 (O_322,N_14511,N_14551);
or UO_323 (O_323,N_14906,N_14879);
or UO_324 (O_324,N_14771,N_14660);
xnor UO_325 (O_325,N_14291,N_14538);
nor UO_326 (O_326,N_14733,N_14343);
nand UO_327 (O_327,N_14254,N_14382);
nor UO_328 (O_328,N_14272,N_14325);
nand UO_329 (O_329,N_14866,N_14782);
or UO_330 (O_330,N_14311,N_14778);
nor UO_331 (O_331,N_14391,N_14416);
xor UO_332 (O_332,N_14363,N_14477);
xor UO_333 (O_333,N_14369,N_14500);
nand UO_334 (O_334,N_14533,N_14535);
and UO_335 (O_335,N_14318,N_14675);
and UO_336 (O_336,N_14547,N_14633);
nor UO_337 (O_337,N_14560,N_14415);
nand UO_338 (O_338,N_14552,N_14572);
nand UO_339 (O_339,N_14738,N_14934);
nor UO_340 (O_340,N_14964,N_14988);
or UO_341 (O_341,N_14281,N_14914);
or UO_342 (O_342,N_14647,N_14856);
or UO_343 (O_343,N_14528,N_14561);
or UO_344 (O_344,N_14679,N_14762);
and UO_345 (O_345,N_14744,N_14822);
or UO_346 (O_346,N_14348,N_14748);
nand UO_347 (O_347,N_14942,N_14307);
and UO_348 (O_348,N_14452,N_14467);
xnor UO_349 (O_349,N_14707,N_14525);
xnor UO_350 (O_350,N_14832,N_14372);
or UO_351 (O_351,N_14306,N_14314);
and UO_352 (O_352,N_14443,N_14905);
nand UO_353 (O_353,N_14603,N_14787);
xnor UO_354 (O_354,N_14310,N_14896);
xnor UO_355 (O_355,N_14584,N_14600);
nand UO_356 (O_356,N_14967,N_14612);
or UO_357 (O_357,N_14566,N_14604);
nor UO_358 (O_358,N_14817,N_14485);
nor UO_359 (O_359,N_14845,N_14952);
and UO_360 (O_360,N_14596,N_14582);
and UO_361 (O_361,N_14271,N_14691);
nand UO_362 (O_362,N_14349,N_14982);
or UO_363 (O_363,N_14950,N_14322);
nand UO_364 (O_364,N_14816,N_14266);
nand UO_365 (O_365,N_14303,N_14808);
nor UO_366 (O_366,N_14927,N_14812);
or UO_367 (O_367,N_14852,N_14453);
nand UO_368 (O_368,N_14800,N_14497);
xnor UO_369 (O_369,N_14537,N_14825);
or UO_370 (O_370,N_14519,N_14269);
or UO_371 (O_371,N_14854,N_14672);
nand UO_372 (O_372,N_14637,N_14490);
nor UO_373 (O_373,N_14724,N_14686);
nor UO_374 (O_374,N_14589,N_14951);
and UO_375 (O_375,N_14969,N_14453);
nor UO_376 (O_376,N_14291,N_14665);
xor UO_377 (O_377,N_14257,N_14741);
nand UO_378 (O_378,N_14721,N_14405);
and UO_379 (O_379,N_14847,N_14586);
or UO_380 (O_380,N_14916,N_14360);
and UO_381 (O_381,N_14979,N_14891);
or UO_382 (O_382,N_14916,N_14790);
nor UO_383 (O_383,N_14722,N_14787);
or UO_384 (O_384,N_14879,N_14453);
nor UO_385 (O_385,N_14272,N_14987);
xor UO_386 (O_386,N_14769,N_14395);
nor UO_387 (O_387,N_14267,N_14781);
xnor UO_388 (O_388,N_14707,N_14667);
and UO_389 (O_389,N_14799,N_14683);
nor UO_390 (O_390,N_14496,N_14594);
nand UO_391 (O_391,N_14817,N_14803);
nand UO_392 (O_392,N_14869,N_14884);
and UO_393 (O_393,N_14297,N_14503);
nand UO_394 (O_394,N_14492,N_14878);
nand UO_395 (O_395,N_14559,N_14796);
xor UO_396 (O_396,N_14905,N_14716);
or UO_397 (O_397,N_14311,N_14486);
and UO_398 (O_398,N_14853,N_14373);
or UO_399 (O_399,N_14855,N_14885);
xnor UO_400 (O_400,N_14328,N_14423);
and UO_401 (O_401,N_14932,N_14810);
nor UO_402 (O_402,N_14868,N_14862);
nand UO_403 (O_403,N_14495,N_14932);
or UO_404 (O_404,N_14771,N_14918);
nand UO_405 (O_405,N_14540,N_14253);
xnor UO_406 (O_406,N_14454,N_14696);
nand UO_407 (O_407,N_14981,N_14339);
or UO_408 (O_408,N_14254,N_14639);
nand UO_409 (O_409,N_14311,N_14891);
or UO_410 (O_410,N_14927,N_14639);
or UO_411 (O_411,N_14591,N_14991);
and UO_412 (O_412,N_14267,N_14947);
or UO_413 (O_413,N_14998,N_14783);
and UO_414 (O_414,N_14299,N_14763);
nor UO_415 (O_415,N_14250,N_14773);
nor UO_416 (O_416,N_14406,N_14252);
and UO_417 (O_417,N_14741,N_14361);
xnor UO_418 (O_418,N_14321,N_14754);
xnor UO_419 (O_419,N_14671,N_14986);
and UO_420 (O_420,N_14772,N_14953);
xor UO_421 (O_421,N_14390,N_14693);
nor UO_422 (O_422,N_14840,N_14525);
nor UO_423 (O_423,N_14297,N_14668);
and UO_424 (O_424,N_14409,N_14720);
nor UO_425 (O_425,N_14751,N_14335);
nand UO_426 (O_426,N_14680,N_14478);
xor UO_427 (O_427,N_14362,N_14571);
xnor UO_428 (O_428,N_14539,N_14637);
nor UO_429 (O_429,N_14820,N_14751);
and UO_430 (O_430,N_14908,N_14503);
and UO_431 (O_431,N_14468,N_14735);
or UO_432 (O_432,N_14869,N_14605);
and UO_433 (O_433,N_14989,N_14424);
or UO_434 (O_434,N_14564,N_14945);
and UO_435 (O_435,N_14760,N_14266);
or UO_436 (O_436,N_14510,N_14783);
nand UO_437 (O_437,N_14338,N_14905);
xor UO_438 (O_438,N_14259,N_14632);
nand UO_439 (O_439,N_14609,N_14335);
and UO_440 (O_440,N_14745,N_14569);
xnor UO_441 (O_441,N_14458,N_14583);
and UO_442 (O_442,N_14849,N_14902);
nor UO_443 (O_443,N_14464,N_14968);
nor UO_444 (O_444,N_14917,N_14590);
or UO_445 (O_445,N_14535,N_14637);
and UO_446 (O_446,N_14300,N_14947);
xor UO_447 (O_447,N_14479,N_14556);
nor UO_448 (O_448,N_14328,N_14521);
xor UO_449 (O_449,N_14505,N_14371);
nor UO_450 (O_450,N_14502,N_14970);
nand UO_451 (O_451,N_14424,N_14338);
and UO_452 (O_452,N_14433,N_14523);
nor UO_453 (O_453,N_14995,N_14433);
or UO_454 (O_454,N_14927,N_14780);
and UO_455 (O_455,N_14646,N_14910);
and UO_456 (O_456,N_14263,N_14328);
or UO_457 (O_457,N_14985,N_14309);
nor UO_458 (O_458,N_14556,N_14855);
nor UO_459 (O_459,N_14466,N_14469);
or UO_460 (O_460,N_14280,N_14306);
xor UO_461 (O_461,N_14413,N_14415);
xnor UO_462 (O_462,N_14868,N_14594);
or UO_463 (O_463,N_14379,N_14847);
and UO_464 (O_464,N_14325,N_14919);
and UO_465 (O_465,N_14413,N_14378);
nor UO_466 (O_466,N_14550,N_14881);
and UO_467 (O_467,N_14296,N_14565);
and UO_468 (O_468,N_14316,N_14264);
nand UO_469 (O_469,N_14730,N_14771);
or UO_470 (O_470,N_14571,N_14977);
nor UO_471 (O_471,N_14436,N_14256);
or UO_472 (O_472,N_14678,N_14682);
or UO_473 (O_473,N_14927,N_14834);
xnor UO_474 (O_474,N_14714,N_14749);
nor UO_475 (O_475,N_14890,N_14750);
xor UO_476 (O_476,N_14428,N_14607);
nor UO_477 (O_477,N_14954,N_14524);
nor UO_478 (O_478,N_14934,N_14852);
xor UO_479 (O_479,N_14958,N_14691);
or UO_480 (O_480,N_14306,N_14368);
or UO_481 (O_481,N_14374,N_14282);
or UO_482 (O_482,N_14445,N_14715);
and UO_483 (O_483,N_14419,N_14564);
xnor UO_484 (O_484,N_14450,N_14418);
and UO_485 (O_485,N_14336,N_14767);
nor UO_486 (O_486,N_14867,N_14591);
nor UO_487 (O_487,N_14863,N_14905);
and UO_488 (O_488,N_14354,N_14618);
xor UO_489 (O_489,N_14467,N_14889);
xor UO_490 (O_490,N_14809,N_14479);
xor UO_491 (O_491,N_14880,N_14919);
nand UO_492 (O_492,N_14974,N_14590);
xor UO_493 (O_493,N_14829,N_14863);
xnor UO_494 (O_494,N_14810,N_14400);
nor UO_495 (O_495,N_14678,N_14584);
nor UO_496 (O_496,N_14373,N_14594);
nand UO_497 (O_497,N_14642,N_14255);
nor UO_498 (O_498,N_14342,N_14784);
or UO_499 (O_499,N_14672,N_14270);
or UO_500 (O_500,N_14599,N_14333);
or UO_501 (O_501,N_14623,N_14764);
xnor UO_502 (O_502,N_14522,N_14817);
nand UO_503 (O_503,N_14756,N_14436);
xor UO_504 (O_504,N_14286,N_14690);
xor UO_505 (O_505,N_14603,N_14348);
and UO_506 (O_506,N_14502,N_14726);
xor UO_507 (O_507,N_14464,N_14276);
or UO_508 (O_508,N_14766,N_14949);
nor UO_509 (O_509,N_14826,N_14715);
nor UO_510 (O_510,N_14949,N_14820);
xnor UO_511 (O_511,N_14559,N_14406);
or UO_512 (O_512,N_14853,N_14413);
nor UO_513 (O_513,N_14430,N_14901);
and UO_514 (O_514,N_14647,N_14807);
and UO_515 (O_515,N_14584,N_14763);
xor UO_516 (O_516,N_14607,N_14406);
nor UO_517 (O_517,N_14570,N_14435);
and UO_518 (O_518,N_14654,N_14502);
xor UO_519 (O_519,N_14387,N_14656);
and UO_520 (O_520,N_14629,N_14809);
nand UO_521 (O_521,N_14271,N_14382);
or UO_522 (O_522,N_14796,N_14281);
nand UO_523 (O_523,N_14799,N_14915);
nor UO_524 (O_524,N_14870,N_14950);
nor UO_525 (O_525,N_14749,N_14259);
and UO_526 (O_526,N_14634,N_14440);
and UO_527 (O_527,N_14463,N_14559);
and UO_528 (O_528,N_14629,N_14684);
and UO_529 (O_529,N_14869,N_14451);
xnor UO_530 (O_530,N_14512,N_14754);
and UO_531 (O_531,N_14584,N_14872);
xor UO_532 (O_532,N_14818,N_14858);
nand UO_533 (O_533,N_14590,N_14423);
or UO_534 (O_534,N_14733,N_14724);
xnor UO_535 (O_535,N_14480,N_14936);
and UO_536 (O_536,N_14581,N_14274);
or UO_537 (O_537,N_14917,N_14523);
and UO_538 (O_538,N_14641,N_14373);
or UO_539 (O_539,N_14886,N_14664);
xor UO_540 (O_540,N_14395,N_14341);
xnor UO_541 (O_541,N_14339,N_14520);
or UO_542 (O_542,N_14424,N_14267);
xor UO_543 (O_543,N_14604,N_14658);
nor UO_544 (O_544,N_14605,N_14715);
nand UO_545 (O_545,N_14761,N_14344);
nor UO_546 (O_546,N_14848,N_14924);
or UO_547 (O_547,N_14978,N_14298);
or UO_548 (O_548,N_14435,N_14648);
xnor UO_549 (O_549,N_14260,N_14750);
nor UO_550 (O_550,N_14379,N_14792);
and UO_551 (O_551,N_14908,N_14675);
and UO_552 (O_552,N_14889,N_14656);
nand UO_553 (O_553,N_14463,N_14671);
nand UO_554 (O_554,N_14842,N_14799);
nand UO_555 (O_555,N_14635,N_14680);
and UO_556 (O_556,N_14930,N_14779);
nor UO_557 (O_557,N_14425,N_14320);
and UO_558 (O_558,N_14397,N_14630);
or UO_559 (O_559,N_14477,N_14787);
or UO_560 (O_560,N_14640,N_14493);
nor UO_561 (O_561,N_14817,N_14476);
xor UO_562 (O_562,N_14644,N_14305);
xor UO_563 (O_563,N_14790,N_14412);
nand UO_564 (O_564,N_14520,N_14447);
and UO_565 (O_565,N_14492,N_14455);
or UO_566 (O_566,N_14295,N_14513);
or UO_567 (O_567,N_14688,N_14468);
nor UO_568 (O_568,N_14452,N_14960);
nor UO_569 (O_569,N_14342,N_14887);
xor UO_570 (O_570,N_14733,N_14965);
and UO_571 (O_571,N_14588,N_14684);
and UO_572 (O_572,N_14984,N_14617);
nor UO_573 (O_573,N_14576,N_14719);
xnor UO_574 (O_574,N_14349,N_14763);
and UO_575 (O_575,N_14568,N_14495);
or UO_576 (O_576,N_14447,N_14588);
nand UO_577 (O_577,N_14439,N_14483);
nand UO_578 (O_578,N_14426,N_14573);
nand UO_579 (O_579,N_14770,N_14372);
nand UO_580 (O_580,N_14339,N_14555);
nor UO_581 (O_581,N_14933,N_14486);
nor UO_582 (O_582,N_14473,N_14515);
or UO_583 (O_583,N_14760,N_14404);
nand UO_584 (O_584,N_14337,N_14705);
xor UO_585 (O_585,N_14659,N_14548);
or UO_586 (O_586,N_14433,N_14909);
or UO_587 (O_587,N_14576,N_14864);
and UO_588 (O_588,N_14358,N_14385);
and UO_589 (O_589,N_14821,N_14421);
xor UO_590 (O_590,N_14620,N_14742);
or UO_591 (O_591,N_14460,N_14258);
or UO_592 (O_592,N_14725,N_14958);
or UO_593 (O_593,N_14509,N_14391);
nor UO_594 (O_594,N_14618,N_14845);
or UO_595 (O_595,N_14488,N_14855);
or UO_596 (O_596,N_14832,N_14734);
xor UO_597 (O_597,N_14852,N_14582);
or UO_598 (O_598,N_14618,N_14858);
and UO_599 (O_599,N_14917,N_14970);
and UO_600 (O_600,N_14828,N_14637);
nor UO_601 (O_601,N_14927,N_14273);
nor UO_602 (O_602,N_14789,N_14737);
xnor UO_603 (O_603,N_14514,N_14851);
nor UO_604 (O_604,N_14409,N_14966);
xor UO_605 (O_605,N_14824,N_14858);
xor UO_606 (O_606,N_14531,N_14856);
nor UO_607 (O_607,N_14929,N_14421);
xor UO_608 (O_608,N_14580,N_14464);
or UO_609 (O_609,N_14397,N_14787);
nand UO_610 (O_610,N_14726,N_14339);
nor UO_611 (O_611,N_14525,N_14472);
and UO_612 (O_612,N_14260,N_14296);
nor UO_613 (O_613,N_14422,N_14502);
and UO_614 (O_614,N_14281,N_14508);
and UO_615 (O_615,N_14877,N_14350);
nor UO_616 (O_616,N_14749,N_14846);
xor UO_617 (O_617,N_14340,N_14745);
xor UO_618 (O_618,N_14368,N_14773);
nor UO_619 (O_619,N_14949,N_14749);
nand UO_620 (O_620,N_14752,N_14998);
nand UO_621 (O_621,N_14838,N_14462);
xnor UO_622 (O_622,N_14784,N_14413);
nor UO_623 (O_623,N_14419,N_14280);
xnor UO_624 (O_624,N_14430,N_14565);
nor UO_625 (O_625,N_14984,N_14499);
or UO_626 (O_626,N_14672,N_14892);
or UO_627 (O_627,N_14782,N_14437);
nand UO_628 (O_628,N_14649,N_14925);
xnor UO_629 (O_629,N_14938,N_14713);
xor UO_630 (O_630,N_14515,N_14832);
and UO_631 (O_631,N_14661,N_14826);
and UO_632 (O_632,N_14421,N_14652);
nor UO_633 (O_633,N_14465,N_14367);
and UO_634 (O_634,N_14603,N_14628);
nor UO_635 (O_635,N_14950,N_14339);
or UO_636 (O_636,N_14813,N_14671);
xnor UO_637 (O_637,N_14444,N_14404);
and UO_638 (O_638,N_14767,N_14960);
xnor UO_639 (O_639,N_14814,N_14432);
xnor UO_640 (O_640,N_14810,N_14386);
or UO_641 (O_641,N_14763,N_14993);
and UO_642 (O_642,N_14953,N_14603);
or UO_643 (O_643,N_14874,N_14804);
and UO_644 (O_644,N_14841,N_14643);
and UO_645 (O_645,N_14667,N_14736);
nor UO_646 (O_646,N_14512,N_14615);
nand UO_647 (O_647,N_14806,N_14738);
nand UO_648 (O_648,N_14464,N_14745);
nor UO_649 (O_649,N_14844,N_14464);
and UO_650 (O_650,N_14583,N_14739);
and UO_651 (O_651,N_14257,N_14549);
and UO_652 (O_652,N_14625,N_14429);
nor UO_653 (O_653,N_14376,N_14753);
nor UO_654 (O_654,N_14369,N_14702);
nand UO_655 (O_655,N_14251,N_14472);
and UO_656 (O_656,N_14885,N_14286);
nand UO_657 (O_657,N_14703,N_14794);
xor UO_658 (O_658,N_14378,N_14402);
or UO_659 (O_659,N_14251,N_14810);
nor UO_660 (O_660,N_14519,N_14744);
xnor UO_661 (O_661,N_14923,N_14735);
and UO_662 (O_662,N_14663,N_14778);
and UO_663 (O_663,N_14600,N_14369);
xnor UO_664 (O_664,N_14718,N_14800);
and UO_665 (O_665,N_14286,N_14318);
xnor UO_666 (O_666,N_14816,N_14253);
nand UO_667 (O_667,N_14413,N_14361);
nor UO_668 (O_668,N_14340,N_14640);
nor UO_669 (O_669,N_14792,N_14951);
xor UO_670 (O_670,N_14981,N_14826);
nor UO_671 (O_671,N_14556,N_14973);
and UO_672 (O_672,N_14579,N_14775);
and UO_673 (O_673,N_14637,N_14510);
nand UO_674 (O_674,N_14931,N_14434);
nor UO_675 (O_675,N_14657,N_14525);
or UO_676 (O_676,N_14942,N_14367);
or UO_677 (O_677,N_14382,N_14713);
nand UO_678 (O_678,N_14955,N_14930);
or UO_679 (O_679,N_14461,N_14930);
or UO_680 (O_680,N_14478,N_14360);
nand UO_681 (O_681,N_14576,N_14295);
nor UO_682 (O_682,N_14675,N_14926);
nand UO_683 (O_683,N_14313,N_14337);
nand UO_684 (O_684,N_14335,N_14573);
or UO_685 (O_685,N_14310,N_14366);
nor UO_686 (O_686,N_14924,N_14958);
xor UO_687 (O_687,N_14717,N_14378);
xor UO_688 (O_688,N_14306,N_14376);
nor UO_689 (O_689,N_14827,N_14823);
and UO_690 (O_690,N_14613,N_14855);
xor UO_691 (O_691,N_14672,N_14957);
xnor UO_692 (O_692,N_14342,N_14675);
or UO_693 (O_693,N_14631,N_14836);
or UO_694 (O_694,N_14627,N_14807);
nand UO_695 (O_695,N_14850,N_14675);
nand UO_696 (O_696,N_14903,N_14484);
nor UO_697 (O_697,N_14944,N_14633);
and UO_698 (O_698,N_14618,N_14657);
and UO_699 (O_699,N_14845,N_14788);
or UO_700 (O_700,N_14934,N_14340);
nand UO_701 (O_701,N_14315,N_14345);
nor UO_702 (O_702,N_14638,N_14291);
nor UO_703 (O_703,N_14431,N_14941);
and UO_704 (O_704,N_14544,N_14724);
or UO_705 (O_705,N_14670,N_14673);
nand UO_706 (O_706,N_14815,N_14415);
nand UO_707 (O_707,N_14480,N_14813);
nor UO_708 (O_708,N_14865,N_14401);
and UO_709 (O_709,N_14421,N_14705);
xor UO_710 (O_710,N_14860,N_14730);
xor UO_711 (O_711,N_14334,N_14964);
or UO_712 (O_712,N_14483,N_14725);
nand UO_713 (O_713,N_14769,N_14522);
nand UO_714 (O_714,N_14338,N_14276);
nand UO_715 (O_715,N_14563,N_14928);
or UO_716 (O_716,N_14571,N_14695);
or UO_717 (O_717,N_14881,N_14955);
nor UO_718 (O_718,N_14742,N_14940);
and UO_719 (O_719,N_14921,N_14858);
and UO_720 (O_720,N_14995,N_14856);
nor UO_721 (O_721,N_14654,N_14590);
and UO_722 (O_722,N_14641,N_14808);
nor UO_723 (O_723,N_14348,N_14912);
nor UO_724 (O_724,N_14637,N_14687);
or UO_725 (O_725,N_14480,N_14535);
and UO_726 (O_726,N_14269,N_14529);
nor UO_727 (O_727,N_14860,N_14597);
or UO_728 (O_728,N_14788,N_14437);
nor UO_729 (O_729,N_14958,N_14303);
xor UO_730 (O_730,N_14840,N_14359);
nor UO_731 (O_731,N_14801,N_14701);
and UO_732 (O_732,N_14539,N_14676);
or UO_733 (O_733,N_14566,N_14989);
nand UO_734 (O_734,N_14611,N_14590);
and UO_735 (O_735,N_14482,N_14468);
xor UO_736 (O_736,N_14404,N_14565);
nor UO_737 (O_737,N_14825,N_14612);
nor UO_738 (O_738,N_14641,N_14778);
nand UO_739 (O_739,N_14829,N_14753);
and UO_740 (O_740,N_14910,N_14950);
nor UO_741 (O_741,N_14285,N_14348);
or UO_742 (O_742,N_14641,N_14357);
nor UO_743 (O_743,N_14446,N_14666);
or UO_744 (O_744,N_14998,N_14547);
nand UO_745 (O_745,N_14529,N_14658);
nor UO_746 (O_746,N_14401,N_14384);
or UO_747 (O_747,N_14434,N_14754);
xnor UO_748 (O_748,N_14748,N_14937);
nand UO_749 (O_749,N_14284,N_14640);
and UO_750 (O_750,N_14881,N_14828);
nand UO_751 (O_751,N_14987,N_14600);
xnor UO_752 (O_752,N_14449,N_14683);
nand UO_753 (O_753,N_14713,N_14583);
nor UO_754 (O_754,N_14907,N_14760);
or UO_755 (O_755,N_14587,N_14537);
nor UO_756 (O_756,N_14452,N_14409);
xnor UO_757 (O_757,N_14497,N_14629);
or UO_758 (O_758,N_14705,N_14730);
and UO_759 (O_759,N_14997,N_14738);
nor UO_760 (O_760,N_14466,N_14340);
nand UO_761 (O_761,N_14456,N_14275);
xnor UO_762 (O_762,N_14629,N_14758);
nand UO_763 (O_763,N_14910,N_14890);
and UO_764 (O_764,N_14873,N_14501);
nor UO_765 (O_765,N_14564,N_14703);
nand UO_766 (O_766,N_14930,N_14361);
or UO_767 (O_767,N_14759,N_14597);
nor UO_768 (O_768,N_14496,N_14364);
xnor UO_769 (O_769,N_14531,N_14347);
or UO_770 (O_770,N_14946,N_14835);
or UO_771 (O_771,N_14693,N_14345);
xor UO_772 (O_772,N_14466,N_14500);
and UO_773 (O_773,N_14932,N_14925);
nor UO_774 (O_774,N_14666,N_14288);
nor UO_775 (O_775,N_14646,N_14300);
nor UO_776 (O_776,N_14331,N_14545);
and UO_777 (O_777,N_14914,N_14343);
or UO_778 (O_778,N_14967,N_14879);
or UO_779 (O_779,N_14798,N_14870);
or UO_780 (O_780,N_14389,N_14626);
and UO_781 (O_781,N_14510,N_14944);
xor UO_782 (O_782,N_14974,N_14997);
nor UO_783 (O_783,N_14973,N_14905);
nor UO_784 (O_784,N_14746,N_14783);
and UO_785 (O_785,N_14863,N_14740);
nand UO_786 (O_786,N_14539,N_14449);
nor UO_787 (O_787,N_14497,N_14811);
xor UO_788 (O_788,N_14440,N_14574);
nand UO_789 (O_789,N_14419,N_14727);
or UO_790 (O_790,N_14802,N_14677);
and UO_791 (O_791,N_14635,N_14973);
nor UO_792 (O_792,N_14968,N_14791);
or UO_793 (O_793,N_14911,N_14593);
nand UO_794 (O_794,N_14716,N_14811);
and UO_795 (O_795,N_14341,N_14358);
and UO_796 (O_796,N_14401,N_14819);
xnor UO_797 (O_797,N_14925,N_14471);
or UO_798 (O_798,N_14740,N_14814);
or UO_799 (O_799,N_14515,N_14403);
nand UO_800 (O_800,N_14558,N_14260);
or UO_801 (O_801,N_14902,N_14254);
nor UO_802 (O_802,N_14770,N_14573);
xnor UO_803 (O_803,N_14452,N_14845);
nor UO_804 (O_804,N_14887,N_14392);
xnor UO_805 (O_805,N_14390,N_14475);
xor UO_806 (O_806,N_14444,N_14471);
xnor UO_807 (O_807,N_14440,N_14359);
nor UO_808 (O_808,N_14695,N_14407);
nand UO_809 (O_809,N_14516,N_14258);
or UO_810 (O_810,N_14368,N_14807);
xnor UO_811 (O_811,N_14380,N_14975);
xor UO_812 (O_812,N_14797,N_14491);
and UO_813 (O_813,N_14783,N_14607);
nor UO_814 (O_814,N_14757,N_14285);
and UO_815 (O_815,N_14534,N_14900);
xor UO_816 (O_816,N_14749,N_14686);
or UO_817 (O_817,N_14546,N_14634);
and UO_818 (O_818,N_14729,N_14505);
nand UO_819 (O_819,N_14725,N_14848);
xnor UO_820 (O_820,N_14555,N_14451);
nand UO_821 (O_821,N_14625,N_14740);
nor UO_822 (O_822,N_14554,N_14961);
nand UO_823 (O_823,N_14783,N_14525);
xnor UO_824 (O_824,N_14352,N_14912);
nand UO_825 (O_825,N_14490,N_14703);
nor UO_826 (O_826,N_14890,N_14539);
nor UO_827 (O_827,N_14519,N_14802);
nand UO_828 (O_828,N_14579,N_14313);
or UO_829 (O_829,N_14543,N_14619);
and UO_830 (O_830,N_14474,N_14592);
and UO_831 (O_831,N_14986,N_14599);
xor UO_832 (O_832,N_14473,N_14360);
and UO_833 (O_833,N_14278,N_14883);
nand UO_834 (O_834,N_14988,N_14800);
and UO_835 (O_835,N_14372,N_14562);
nor UO_836 (O_836,N_14610,N_14621);
and UO_837 (O_837,N_14599,N_14796);
nor UO_838 (O_838,N_14492,N_14376);
and UO_839 (O_839,N_14993,N_14988);
xor UO_840 (O_840,N_14822,N_14734);
and UO_841 (O_841,N_14532,N_14462);
nand UO_842 (O_842,N_14915,N_14482);
or UO_843 (O_843,N_14936,N_14533);
nand UO_844 (O_844,N_14476,N_14948);
and UO_845 (O_845,N_14566,N_14485);
or UO_846 (O_846,N_14620,N_14520);
and UO_847 (O_847,N_14508,N_14701);
nand UO_848 (O_848,N_14822,N_14831);
nand UO_849 (O_849,N_14914,N_14315);
nand UO_850 (O_850,N_14282,N_14831);
nor UO_851 (O_851,N_14645,N_14505);
and UO_852 (O_852,N_14596,N_14668);
nor UO_853 (O_853,N_14260,N_14356);
nand UO_854 (O_854,N_14252,N_14642);
xnor UO_855 (O_855,N_14644,N_14691);
and UO_856 (O_856,N_14910,N_14587);
nand UO_857 (O_857,N_14787,N_14771);
or UO_858 (O_858,N_14842,N_14764);
or UO_859 (O_859,N_14362,N_14599);
and UO_860 (O_860,N_14633,N_14478);
xor UO_861 (O_861,N_14595,N_14549);
and UO_862 (O_862,N_14821,N_14759);
and UO_863 (O_863,N_14648,N_14671);
and UO_864 (O_864,N_14545,N_14722);
xor UO_865 (O_865,N_14589,N_14261);
or UO_866 (O_866,N_14820,N_14883);
nand UO_867 (O_867,N_14779,N_14481);
or UO_868 (O_868,N_14526,N_14914);
nor UO_869 (O_869,N_14728,N_14491);
nand UO_870 (O_870,N_14387,N_14585);
nand UO_871 (O_871,N_14545,N_14520);
or UO_872 (O_872,N_14277,N_14670);
nand UO_873 (O_873,N_14943,N_14649);
nor UO_874 (O_874,N_14527,N_14273);
and UO_875 (O_875,N_14276,N_14751);
nand UO_876 (O_876,N_14590,N_14921);
nand UO_877 (O_877,N_14822,N_14684);
nand UO_878 (O_878,N_14590,N_14645);
nand UO_879 (O_879,N_14967,N_14800);
and UO_880 (O_880,N_14819,N_14828);
nand UO_881 (O_881,N_14952,N_14311);
and UO_882 (O_882,N_14329,N_14620);
nor UO_883 (O_883,N_14696,N_14777);
and UO_884 (O_884,N_14494,N_14285);
nand UO_885 (O_885,N_14728,N_14574);
xnor UO_886 (O_886,N_14755,N_14644);
nor UO_887 (O_887,N_14652,N_14462);
xor UO_888 (O_888,N_14627,N_14961);
nor UO_889 (O_889,N_14345,N_14949);
or UO_890 (O_890,N_14477,N_14815);
nor UO_891 (O_891,N_14653,N_14502);
or UO_892 (O_892,N_14610,N_14805);
or UO_893 (O_893,N_14443,N_14474);
and UO_894 (O_894,N_14555,N_14974);
or UO_895 (O_895,N_14759,N_14459);
or UO_896 (O_896,N_14271,N_14891);
and UO_897 (O_897,N_14568,N_14582);
and UO_898 (O_898,N_14722,N_14325);
xnor UO_899 (O_899,N_14402,N_14275);
nor UO_900 (O_900,N_14447,N_14377);
and UO_901 (O_901,N_14659,N_14839);
nor UO_902 (O_902,N_14776,N_14251);
nor UO_903 (O_903,N_14356,N_14297);
xnor UO_904 (O_904,N_14519,N_14464);
or UO_905 (O_905,N_14821,N_14251);
nor UO_906 (O_906,N_14634,N_14987);
nand UO_907 (O_907,N_14665,N_14477);
nor UO_908 (O_908,N_14986,N_14694);
and UO_909 (O_909,N_14861,N_14685);
nand UO_910 (O_910,N_14935,N_14474);
xor UO_911 (O_911,N_14711,N_14463);
nor UO_912 (O_912,N_14897,N_14788);
or UO_913 (O_913,N_14961,N_14359);
nor UO_914 (O_914,N_14738,N_14589);
xnor UO_915 (O_915,N_14785,N_14407);
xor UO_916 (O_916,N_14980,N_14499);
nor UO_917 (O_917,N_14755,N_14932);
xor UO_918 (O_918,N_14702,N_14849);
nand UO_919 (O_919,N_14392,N_14511);
xor UO_920 (O_920,N_14290,N_14256);
and UO_921 (O_921,N_14501,N_14382);
xor UO_922 (O_922,N_14881,N_14912);
or UO_923 (O_923,N_14703,N_14386);
and UO_924 (O_924,N_14257,N_14419);
nand UO_925 (O_925,N_14291,N_14425);
nor UO_926 (O_926,N_14678,N_14644);
xor UO_927 (O_927,N_14401,N_14458);
or UO_928 (O_928,N_14394,N_14831);
xnor UO_929 (O_929,N_14813,N_14547);
nor UO_930 (O_930,N_14480,N_14471);
xnor UO_931 (O_931,N_14400,N_14355);
xnor UO_932 (O_932,N_14859,N_14630);
nand UO_933 (O_933,N_14888,N_14707);
nor UO_934 (O_934,N_14370,N_14777);
and UO_935 (O_935,N_14971,N_14901);
nand UO_936 (O_936,N_14504,N_14482);
nor UO_937 (O_937,N_14748,N_14699);
xnor UO_938 (O_938,N_14289,N_14683);
nor UO_939 (O_939,N_14736,N_14519);
nor UO_940 (O_940,N_14988,N_14508);
nand UO_941 (O_941,N_14835,N_14634);
nand UO_942 (O_942,N_14664,N_14806);
nor UO_943 (O_943,N_14596,N_14614);
or UO_944 (O_944,N_14639,N_14382);
xor UO_945 (O_945,N_14452,N_14423);
or UO_946 (O_946,N_14354,N_14917);
nor UO_947 (O_947,N_14664,N_14958);
nand UO_948 (O_948,N_14460,N_14707);
or UO_949 (O_949,N_14559,N_14522);
and UO_950 (O_950,N_14916,N_14999);
or UO_951 (O_951,N_14565,N_14323);
or UO_952 (O_952,N_14572,N_14702);
xnor UO_953 (O_953,N_14504,N_14777);
or UO_954 (O_954,N_14480,N_14297);
nand UO_955 (O_955,N_14792,N_14873);
and UO_956 (O_956,N_14281,N_14600);
nor UO_957 (O_957,N_14384,N_14353);
and UO_958 (O_958,N_14283,N_14619);
and UO_959 (O_959,N_14536,N_14304);
xnor UO_960 (O_960,N_14361,N_14672);
or UO_961 (O_961,N_14454,N_14942);
xor UO_962 (O_962,N_14307,N_14977);
and UO_963 (O_963,N_14810,N_14785);
and UO_964 (O_964,N_14296,N_14673);
nor UO_965 (O_965,N_14769,N_14363);
and UO_966 (O_966,N_14757,N_14749);
nand UO_967 (O_967,N_14361,N_14779);
nand UO_968 (O_968,N_14301,N_14510);
xor UO_969 (O_969,N_14769,N_14440);
nor UO_970 (O_970,N_14552,N_14295);
or UO_971 (O_971,N_14441,N_14640);
xor UO_972 (O_972,N_14422,N_14452);
or UO_973 (O_973,N_14994,N_14272);
and UO_974 (O_974,N_14603,N_14534);
and UO_975 (O_975,N_14525,N_14339);
or UO_976 (O_976,N_14661,N_14639);
nand UO_977 (O_977,N_14836,N_14959);
and UO_978 (O_978,N_14299,N_14880);
nor UO_979 (O_979,N_14814,N_14534);
nor UO_980 (O_980,N_14644,N_14360);
nand UO_981 (O_981,N_14334,N_14540);
nor UO_982 (O_982,N_14395,N_14869);
xnor UO_983 (O_983,N_14851,N_14991);
xnor UO_984 (O_984,N_14986,N_14603);
xor UO_985 (O_985,N_14615,N_14393);
and UO_986 (O_986,N_14817,N_14949);
nor UO_987 (O_987,N_14315,N_14459);
xor UO_988 (O_988,N_14595,N_14515);
and UO_989 (O_989,N_14257,N_14963);
nand UO_990 (O_990,N_14451,N_14430);
nand UO_991 (O_991,N_14767,N_14902);
and UO_992 (O_992,N_14834,N_14877);
xor UO_993 (O_993,N_14864,N_14422);
nor UO_994 (O_994,N_14521,N_14313);
nand UO_995 (O_995,N_14846,N_14508);
xnor UO_996 (O_996,N_14589,N_14775);
or UO_997 (O_997,N_14949,N_14618);
xnor UO_998 (O_998,N_14932,N_14471);
xor UO_999 (O_999,N_14343,N_14416);
or UO_1000 (O_1000,N_14460,N_14825);
or UO_1001 (O_1001,N_14660,N_14862);
xnor UO_1002 (O_1002,N_14270,N_14457);
or UO_1003 (O_1003,N_14671,N_14765);
nand UO_1004 (O_1004,N_14465,N_14785);
and UO_1005 (O_1005,N_14901,N_14677);
and UO_1006 (O_1006,N_14725,N_14580);
xor UO_1007 (O_1007,N_14931,N_14776);
nor UO_1008 (O_1008,N_14950,N_14425);
or UO_1009 (O_1009,N_14492,N_14953);
nor UO_1010 (O_1010,N_14346,N_14276);
xor UO_1011 (O_1011,N_14464,N_14405);
nor UO_1012 (O_1012,N_14288,N_14902);
xnor UO_1013 (O_1013,N_14662,N_14696);
nor UO_1014 (O_1014,N_14580,N_14572);
or UO_1015 (O_1015,N_14342,N_14472);
xnor UO_1016 (O_1016,N_14979,N_14310);
nand UO_1017 (O_1017,N_14444,N_14483);
nand UO_1018 (O_1018,N_14434,N_14261);
and UO_1019 (O_1019,N_14320,N_14705);
xnor UO_1020 (O_1020,N_14973,N_14917);
nand UO_1021 (O_1021,N_14789,N_14458);
xnor UO_1022 (O_1022,N_14926,N_14993);
or UO_1023 (O_1023,N_14578,N_14319);
nand UO_1024 (O_1024,N_14877,N_14274);
nand UO_1025 (O_1025,N_14881,N_14674);
nor UO_1026 (O_1026,N_14388,N_14372);
or UO_1027 (O_1027,N_14746,N_14880);
and UO_1028 (O_1028,N_14975,N_14472);
or UO_1029 (O_1029,N_14904,N_14368);
nor UO_1030 (O_1030,N_14486,N_14928);
nand UO_1031 (O_1031,N_14571,N_14912);
or UO_1032 (O_1032,N_14469,N_14321);
nand UO_1033 (O_1033,N_14415,N_14372);
nor UO_1034 (O_1034,N_14791,N_14733);
nor UO_1035 (O_1035,N_14742,N_14881);
and UO_1036 (O_1036,N_14473,N_14642);
nand UO_1037 (O_1037,N_14995,N_14636);
or UO_1038 (O_1038,N_14371,N_14798);
or UO_1039 (O_1039,N_14594,N_14677);
or UO_1040 (O_1040,N_14789,N_14817);
nor UO_1041 (O_1041,N_14994,N_14884);
nand UO_1042 (O_1042,N_14706,N_14987);
or UO_1043 (O_1043,N_14593,N_14902);
xnor UO_1044 (O_1044,N_14737,N_14341);
and UO_1045 (O_1045,N_14531,N_14818);
xor UO_1046 (O_1046,N_14484,N_14553);
nand UO_1047 (O_1047,N_14261,N_14927);
xnor UO_1048 (O_1048,N_14322,N_14366);
and UO_1049 (O_1049,N_14465,N_14829);
nor UO_1050 (O_1050,N_14340,N_14663);
nor UO_1051 (O_1051,N_14275,N_14413);
nor UO_1052 (O_1052,N_14986,N_14951);
xor UO_1053 (O_1053,N_14606,N_14463);
or UO_1054 (O_1054,N_14908,N_14376);
or UO_1055 (O_1055,N_14878,N_14884);
nand UO_1056 (O_1056,N_14812,N_14661);
nor UO_1057 (O_1057,N_14310,N_14407);
nor UO_1058 (O_1058,N_14653,N_14925);
or UO_1059 (O_1059,N_14303,N_14420);
or UO_1060 (O_1060,N_14847,N_14901);
nand UO_1061 (O_1061,N_14409,N_14697);
nor UO_1062 (O_1062,N_14289,N_14395);
and UO_1063 (O_1063,N_14451,N_14634);
and UO_1064 (O_1064,N_14288,N_14539);
and UO_1065 (O_1065,N_14840,N_14326);
nand UO_1066 (O_1066,N_14813,N_14887);
nor UO_1067 (O_1067,N_14283,N_14528);
nand UO_1068 (O_1068,N_14562,N_14698);
xnor UO_1069 (O_1069,N_14515,N_14267);
and UO_1070 (O_1070,N_14481,N_14252);
or UO_1071 (O_1071,N_14927,N_14455);
or UO_1072 (O_1072,N_14417,N_14320);
nand UO_1073 (O_1073,N_14814,N_14785);
and UO_1074 (O_1074,N_14841,N_14250);
nor UO_1075 (O_1075,N_14538,N_14702);
and UO_1076 (O_1076,N_14955,N_14459);
xor UO_1077 (O_1077,N_14997,N_14757);
nand UO_1078 (O_1078,N_14266,N_14511);
nand UO_1079 (O_1079,N_14404,N_14435);
or UO_1080 (O_1080,N_14478,N_14402);
nor UO_1081 (O_1081,N_14483,N_14276);
nor UO_1082 (O_1082,N_14906,N_14611);
or UO_1083 (O_1083,N_14864,N_14899);
or UO_1084 (O_1084,N_14635,N_14282);
nor UO_1085 (O_1085,N_14820,N_14695);
xnor UO_1086 (O_1086,N_14601,N_14402);
nand UO_1087 (O_1087,N_14325,N_14937);
nand UO_1088 (O_1088,N_14742,N_14984);
and UO_1089 (O_1089,N_14828,N_14490);
or UO_1090 (O_1090,N_14500,N_14507);
or UO_1091 (O_1091,N_14616,N_14702);
xor UO_1092 (O_1092,N_14332,N_14330);
xor UO_1093 (O_1093,N_14823,N_14772);
xor UO_1094 (O_1094,N_14932,N_14304);
nand UO_1095 (O_1095,N_14978,N_14902);
and UO_1096 (O_1096,N_14533,N_14429);
or UO_1097 (O_1097,N_14654,N_14626);
nor UO_1098 (O_1098,N_14861,N_14892);
nor UO_1099 (O_1099,N_14590,N_14446);
xor UO_1100 (O_1100,N_14848,N_14738);
or UO_1101 (O_1101,N_14573,N_14748);
or UO_1102 (O_1102,N_14899,N_14938);
or UO_1103 (O_1103,N_14492,N_14884);
or UO_1104 (O_1104,N_14724,N_14339);
or UO_1105 (O_1105,N_14479,N_14719);
xor UO_1106 (O_1106,N_14745,N_14813);
xor UO_1107 (O_1107,N_14607,N_14279);
and UO_1108 (O_1108,N_14574,N_14873);
nand UO_1109 (O_1109,N_14696,N_14458);
nor UO_1110 (O_1110,N_14634,N_14751);
nand UO_1111 (O_1111,N_14951,N_14942);
nor UO_1112 (O_1112,N_14798,N_14502);
nor UO_1113 (O_1113,N_14583,N_14879);
and UO_1114 (O_1114,N_14351,N_14400);
nand UO_1115 (O_1115,N_14804,N_14823);
nor UO_1116 (O_1116,N_14802,N_14291);
nand UO_1117 (O_1117,N_14592,N_14822);
or UO_1118 (O_1118,N_14439,N_14669);
nand UO_1119 (O_1119,N_14279,N_14713);
nand UO_1120 (O_1120,N_14534,N_14821);
nor UO_1121 (O_1121,N_14657,N_14818);
xnor UO_1122 (O_1122,N_14501,N_14385);
xor UO_1123 (O_1123,N_14362,N_14743);
xnor UO_1124 (O_1124,N_14692,N_14434);
nand UO_1125 (O_1125,N_14341,N_14974);
xnor UO_1126 (O_1126,N_14813,N_14429);
nor UO_1127 (O_1127,N_14862,N_14372);
or UO_1128 (O_1128,N_14616,N_14445);
nand UO_1129 (O_1129,N_14368,N_14926);
or UO_1130 (O_1130,N_14737,N_14819);
xor UO_1131 (O_1131,N_14555,N_14664);
nand UO_1132 (O_1132,N_14547,N_14291);
or UO_1133 (O_1133,N_14287,N_14762);
or UO_1134 (O_1134,N_14286,N_14679);
and UO_1135 (O_1135,N_14915,N_14488);
nand UO_1136 (O_1136,N_14478,N_14313);
and UO_1137 (O_1137,N_14791,N_14471);
or UO_1138 (O_1138,N_14356,N_14372);
xor UO_1139 (O_1139,N_14836,N_14286);
nand UO_1140 (O_1140,N_14298,N_14342);
and UO_1141 (O_1141,N_14598,N_14618);
or UO_1142 (O_1142,N_14640,N_14884);
and UO_1143 (O_1143,N_14599,N_14612);
or UO_1144 (O_1144,N_14803,N_14789);
xnor UO_1145 (O_1145,N_14996,N_14841);
and UO_1146 (O_1146,N_14295,N_14911);
nand UO_1147 (O_1147,N_14692,N_14328);
and UO_1148 (O_1148,N_14408,N_14656);
nor UO_1149 (O_1149,N_14915,N_14712);
or UO_1150 (O_1150,N_14696,N_14872);
and UO_1151 (O_1151,N_14994,N_14977);
and UO_1152 (O_1152,N_14740,N_14691);
xor UO_1153 (O_1153,N_14439,N_14650);
nor UO_1154 (O_1154,N_14272,N_14503);
or UO_1155 (O_1155,N_14922,N_14425);
nor UO_1156 (O_1156,N_14645,N_14853);
and UO_1157 (O_1157,N_14272,N_14949);
nand UO_1158 (O_1158,N_14736,N_14889);
or UO_1159 (O_1159,N_14929,N_14256);
nand UO_1160 (O_1160,N_14891,N_14538);
and UO_1161 (O_1161,N_14886,N_14576);
nor UO_1162 (O_1162,N_14538,N_14632);
xor UO_1163 (O_1163,N_14755,N_14410);
or UO_1164 (O_1164,N_14432,N_14784);
nand UO_1165 (O_1165,N_14882,N_14969);
nand UO_1166 (O_1166,N_14820,N_14455);
nand UO_1167 (O_1167,N_14562,N_14640);
nor UO_1168 (O_1168,N_14491,N_14768);
nor UO_1169 (O_1169,N_14656,N_14601);
nand UO_1170 (O_1170,N_14814,N_14640);
and UO_1171 (O_1171,N_14830,N_14739);
xor UO_1172 (O_1172,N_14715,N_14694);
and UO_1173 (O_1173,N_14367,N_14495);
xor UO_1174 (O_1174,N_14860,N_14773);
and UO_1175 (O_1175,N_14691,N_14962);
and UO_1176 (O_1176,N_14698,N_14357);
and UO_1177 (O_1177,N_14901,N_14836);
nand UO_1178 (O_1178,N_14252,N_14568);
or UO_1179 (O_1179,N_14952,N_14591);
and UO_1180 (O_1180,N_14402,N_14414);
xnor UO_1181 (O_1181,N_14835,N_14773);
or UO_1182 (O_1182,N_14481,N_14959);
xnor UO_1183 (O_1183,N_14537,N_14670);
nand UO_1184 (O_1184,N_14935,N_14701);
and UO_1185 (O_1185,N_14741,N_14561);
nor UO_1186 (O_1186,N_14674,N_14724);
or UO_1187 (O_1187,N_14808,N_14331);
xor UO_1188 (O_1188,N_14604,N_14645);
or UO_1189 (O_1189,N_14748,N_14343);
or UO_1190 (O_1190,N_14803,N_14987);
or UO_1191 (O_1191,N_14393,N_14557);
nor UO_1192 (O_1192,N_14891,N_14425);
and UO_1193 (O_1193,N_14696,N_14309);
and UO_1194 (O_1194,N_14817,N_14738);
nand UO_1195 (O_1195,N_14457,N_14467);
nand UO_1196 (O_1196,N_14478,N_14552);
xor UO_1197 (O_1197,N_14360,N_14786);
xnor UO_1198 (O_1198,N_14282,N_14871);
nand UO_1199 (O_1199,N_14366,N_14610);
xnor UO_1200 (O_1200,N_14682,N_14522);
and UO_1201 (O_1201,N_14840,N_14730);
xnor UO_1202 (O_1202,N_14567,N_14942);
and UO_1203 (O_1203,N_14513,N_14564);
nor UO_1204 (O_1204,N_14603,N_14277);
nor UO_1205 (O_1205,N_14513,N_14747);
nor UO_1206 (O_1206,N_14498,N_14605);
nand UO_1207 (O_1207,N_14554,N_14434);
nor UO_1208 (O_1208,N_14390,N_14413);
or UO_1209 (O_1209,N_14324,N_14363);
or UO_1210 (O_1210,N_14646,N_14931);
nand UO_1211 (O_1211,N_14532,N_14850);
xnor UO_1212 (O_1212,N_14390,N_14400);
nand UO_1213 (O_1213,N_14668,N_14820);
nor UO_1214 (O_1214,N_14392,N_14683);
or UO_1215 (O_1215,N_14508,N_14881);
nor UO_1216 (O_1216,N_14645,N_14850);
and UO_1217 (O_1217,N_14765,N_14903);
and UO_1218 (O_1218,N_14699,N_14866);
nor UO_1219 (O_1219,N_14711,N_14466);
and UO_1220 (O_1220,N_14478,N_14265);
xnor UO_1221 (O_1221,N_14879,N_14489);
and UO_1222 (O_1222,N_14909,N_14555);
nand UO_1223 (O_1223,N_14532,N_14543);
xor UO_1224 (O_1224,N_14888,N_14821);
xor UO_1225 (O_1225,N_14594,N_14328);
or UO_1226 (O_1226,N_14877,N_14693);
xnor UO_1227 (O_1227,N_14427,N_14465);
xor UO_1228 (O_1228,N_14554,N_14765);
or UO_1229 (O_1229,N_14640,N_14865);
and UO_1230 (O_1230,N_14569,N_14582);
nand UO_1231 (O_1231,N_14643,N_14337);
nand UO_1232 (O_1232,N_14997,N_14520);
xor UO_1233 (O_1233,N_14818,N_14890);
and UO_1234 (O_1234,N_14690,N_14425);
nor UO_1235 (O_1235,N_14796,N_14820);
nand UO_1236 (O_1236,N_14794,N_14560);
nand UO_1237 (O_1237,N_14645,N_14924);
nor UO_1238 (O_1238,N_14636,N_14319);
or UO_1239 (O_1239,N_14264,N_14354);
nand UO_1240 (O_1240,N_14430,N_14997);
xor UO_1241 (O_1241,N_14692,N_14396);
or UO_1242 (O_1242,N_14256,N_14849);
nand UO_1243 (O_1243,N_14374,N_14967);
and UO_1244 (O_1244,N_14681,N_14632);
nand UO_1245 (O_1245,N_14404,N_14682);
nor UO_1246 (O_1246,N_14477,N_14399);
and UO_1247 (O_1247,N_14612,N_14976);
or UO_1248 (O_1248,N_14742,N_14843);
or UO_1249 (O_1249,N_14971,N_14362);
nor UO_1250 (O_1250,N_14308,N_14456);
xnor UO_1251 (O_1251,N_14708,N_14377);
nor UO_1252 (O_1252,N_14448,N_14754);
nand UO_1253 (O_1253,N_14418,N_14407);
xor UO_1254 (O_1254,N_14975,N_14386);
nand UO_1255 (O_1255,N_14866,N_14739);
nor UO_1256 (O_1256,N_14281,N_14918);
or UO_1257 (O_1257,N_14803,N_14757);
and UO_1258 (O_1258,N_14437,N_14972);
nor UO_1259 (O_1259,N_14759,N_14655);
and UO_1260 (O_1260,N_14700,N_14882);
or UO_1261 (O_1261,N_14521,N_14868);
or UO_1262 (O_1262,N_14919,N_14881);
or UO_1263 (O_1263,N_14413,N_14723);
xor UO_1264 (O_1264,N_14822,N_14302);
and UO_1265 (O_1265,N_14816,N_14972);
or UO_1266 (O_1266,N_14485,N_14929);
xor UO_1267 (O_1267,N_14525,N_14788);
xor UO_1268 (O_1268,N_14458,N_14405);
xor UO_1269 (O_1269,N_14703,N_14284);
or UO_1270 (O_1270,N_14616,N_14314);
nand UO_1271 (O_1271,N_14437,N_14389);
xor UO_1272 (O_1272,N_14428,N_14688);
nand UO_1273 (O_1273,N_14929,N_14608);
xor UO_1274 (O_1274,N_14747,N_14366);
or UO_1275 (O_1275,N_14411,N_14307);
nor UO_1276 (O_1276,N_14431,N_14716);
nand UO_1277 (O_1277,N_14871,N_14442);
and UO_1278 (O_1278,N_14698,N_14348);
nand UO_1279 (O_1279,N_14578,N_14445);
nand UO_1280 (O_1280,N_14653,N_14572);
or UO_1281 (O_1281,N_14539,N_14811);
or UO_1282 (O_1282,N_14585,N_14326);
xnor UO_1283 (O_1283,N_14574,N_14917);
nor UO_1284 (O_1284,N_14291,N_14391);
xor UO_1285 (O_1285,N_14316,N_14288);
and UO_1286 (O_1286,N_14559,N_14255);
nand UO_1287 (O_1287,N_14750,N_14418);
and UO_1288 (O_1288,N_14822,N_14978);
nand UO_1289 (O_1289,N_14367,N_14324);
and UO_1290 (O_1290,N_14850,N_14634);
nand UO_1291 (O_1291,N_14471,N_14615);
or UO_1292 (O_1292,N_14510,N_14644);
and UO_1293 (O_1293,N_14625,N_14694);
nor UO_1294 (O_1294,N_14691,N_14712);
and UO_1295 (O_1295,N_14680,N_14817);
nor UO_1296 (O_1296,N_14787,N_14544);
xor UO_1297 (O_1297,N_14801,N_14335);
nor UO_1298 (O_1298,N_14435,N_14605);
nor UO_1299 (O_1299,N_14755,N_14453);
and UO_1300 (O_1300,N_14588,N_14875);
and UO_1301 (O_1301,N_14986,N_14974);
nor UO_1302 (O_1302,N_14926,N_14408);
and UO_1303 (O_1303,N_14355,N_14578);
and UO_1304 (O_1304,N_14653,N_14616);
or UO_1305 (O_1305,N_14336,N_14788);
and UO_1306 (O_1306,N_14312,N_14622);
or UO_1307 (O_1307,N_14680,N_14362);
xor UO_1308 (O_1308,N_14970,N_14775);
xnor UO_1309 (O_1309,N_14465,N_14605);
nor UO_1310 (O_1310,N_14544,N_14679);
and UO_1311 (O_1311,N_14363,N_14934);
and UO_1312 (O_1312,N_14738,N_14987);
and UO_1313 (O_1313,N_14830,N_14761);
xor UO_1314 (O_1314,N_14997,N_14327);
and UO_1315 (O_1315,N_14473,N_14506);
or UO_1316 (O_1316,N_14530,N_14761);
xor UO_1317 (O_1317,N_14972,N_14331);
nor UO_1318 (O_1318,N_14306,N_14466);
or UO_1319 (O_1319,N_14305,N_14502);
and UO_1320 (O_1320,N_14401,N_14573);
nand UO_1321 (O_1321,N_14931,N_14348);
xor UO_1322 (O_1322,N_14522,N_14732);
xor UO_1323 (O_1323,N_14277,N_14553);
xor UO_1324 (O_1324,N_14786,N_14491);
and UO_1325 (O_1325,N_14873,N_14784);
or UO_1326 (O_1326,N_14565,N_14998);
and UO_1327 (O_1327,N_14446,N_14608);
xor UO_1328 (O_1328,N_14652,N_14848);
nand UO_1329 (O_1329,N_14574,N_14898);
and UO_1330 (O_1330,N_14743,N_14968);
and UO_1331 (O_1331,N_14566,N_14700);
nand UO_1332 (O_1332,N_14554,N_14710);
xor UO_1333 (O_1333,N_14956,N_14513);
or UO_1334 (O_1334,N_14975,N_14259);
and UO_1335 (O_1335,N_14523,N_14583);
xnor UO_1336 (O_1336,N_14780,N_14532);
nand UO_1337 (O_1337,N_14829,N_14936);
and UO_1338 (O_1338,N_14741,N_14927);
or UO_1339 (O_1339,N_14902,N_14644);
or UO_1340 (O_1340,N_14921,N_14566);
nor UO_1341 (O_1341,N_14897,N_14747);
nand UO_1342 (O_1342,N_14376,N_14543);
nand UO_1343 (O_1343,N_14714,N_14365);
and UO_1344 (O_1344,N_14678,N_14570);
nor UO_1345 (O_1345,N_14759,N_14620);
nor UO_1346 (O_1346,N_14970,N_14990);
nor UO_1347 (O_1347,N_14755,N_14539);
or UO_1348 (O_1348,N_14308,N_14682);
and UO_1349 (O_1349,N_14806,N_14855);
nand UO_1350 (O_1350,N_14627,N_14572);
or UO_1351 (O_1351,N_14870,N_14623);
xor UO_1352 (O_1352,N_14403,N_14842);
xor UO_1353 (O_1353,N_14740,N_14862);
nand UO_1354 (O_1354,N_14952,N_14931);
and UO_1355 (O_1355,N_14877,N_14329);
nand UO_1356 (O_1356,N_14777,N_14760);
xnor UO_1357 (O_1357,N_14726,N_14328);
and UO_1358 (O_1358,N_14597,N_14595);
or UO_1359 (O_1359,N_14903,N_14932);
xor UO_1360 (O_1360,N_14724,N_14515);
or UO_1361 (O_1361,N_14938,N_14309);
xnor UO_1362 (O_1362,N_14541,N_14520);
nor UO_1363 (O_1363,N_14698,N_14544);
nand UO_1364 (O_1364,N_14464,N_14994);
xnor UO_1365 (O_1365,N_14954,N_14551);
nor UO_1366 (O_1366,N_14708,N_14423);
nor UO_1367 (O_1367,N_14327,N_14475);
and UO_1368 (O_1368,N_14729,N_14566);
nand UO_1369 (O_1369,N_14426,N_14256);
nand UO_1370 (O_1370,N_14333,N_14971);
nand UO_1371 (O_1371,N_14503,N_14548);
nand UO_1372 (O_1372,N_14449,N_14559);
xnor UO_1373 (O_1373,N_14650,N_14901);
or UO_1374 (O_1374,N_14347,N_14477);
or UO_1375 (O_1375,N_14813,N_14754);
or UO_1376 (O_1376,N_14713,N_14421);
xor UO_1377 (O_1377,N_14515,N_14722);
xor UO_1378 (O_1378,N_14259,N_14280);
nand UO_1379 (O_1379,N_14289,N_14878);
and UO_1380 (O_1380,N_14347,N_14488);
xor UO_1381 (O_1381,N_14568,N_14546);
xor UO_1382 (O_1382,N_14286,N_14822);
and UO_1383 (O_1383,N_14373,N_14767);
nand UO_1384 (O_1384,N_14323,N_14621);
or UO_1385 (O_1385,N_14379,N_14492);
and UO_1386 (O_1386,N_14970,N_14518);
xor UO_1387 (O_1387,N_14407,N_14578);
nor UO_1388 (O_1388,N_14733,N_14788);
and UO_1389 (O_1389,N_14623,N_14751);
nor UO_1390 (O_1390,N_14853,N_14349);
xor UO_1391 (O_1391,N_14336,N_14822);
or UO_1392 (O_1392,N_14497,N_14442);
nor UO_1393 (O_1393,N_14859,N_14521);
xnor UO_1394 (O_1394,N_14368,N_14460);
and UO_1395 (O_1395,N_14751,N_14484);
and UO_1396 (O_1396,N_14283,N_14507);
nor UO_1397 (O_1397,N_14378,N_14761);
nand UO_1398 (O_1398,N_14724,N_14383);
nand UO_1399 (O_1399,N_14275,N_14985);
nand UO_1400 (O_1400,N_14269,N_14870);
nor UO_1401 (O_1401,N_14435,N_14925);
xor UO_1402 (O_1402,N_14367,N_14603);
nand UO_1403 (O_1403,N_14735,N_14303);
and UO_1404 (O_1404,N_14361,N_14311);
nor UO_1405 (O_1405,N_14591,N_14600);
or UO_1406 (O_1406,N_14890,N_14378);
xor UO_1407 (O_1407,N_14751,N_14610);
and UO_1408 (O_1408,N_14469,N_14911);
nand UO_1409 (O_1409,N_14690,N_14659);
and UO_1410 (O_1410,N_14348,N_14417);
or UO_1411 (O_1411,N_14287,N_14729);
xnor UO_1412 (O_1412,N_14503,N_14940);
and UO_1413 (O_1413,N_14644,N_14677);
xnor UO_1414 (O_1414,N_14861,N_14827);
and UO_1415 (O_1415,N_14510,N_14973);
or UO_1416 (O_1416,N_14453,N_14384);
and UO_1417 (O_1417,N_14818,N_14311);
nand UO_1418 (O_1418,N_14797,N_14751);
nor UO_1419 (O_1419,N_14878,N_14882);
nor UO_1420 (O_1420,N_14675,N_14862);
nor UO_1421 (O_1421,N_14365,N_14391);
xnor UO_1422 (O_1422,N_14437,N_14800);
and UO_1423 (O_1423,N_14448,N_14741);
and UO_1424 (O_1424,N_14835,N_14674);
xnor UO_1425 (O_1425,N_14534,N_14818);
xnor UO_1426 (O_1426,N_14736,N_14501);
xnor UO_1427 (O_1427,N_14696,N_14631);
or UO_1428 (O_1428,N_14820,N_14526);
nor UO_1429 (O_1429,N_14308,N_14392);
and UO_1430 (O_1430,N_14935,N_14369);
xor UO_1431 (O_1431,N_14998,N_14957);
nand UO_1432 (O_1432,N_14857,N_14517);
xor UO_1433 (O_1433,N_14268,N_14666);
nand UO_1434 (O_1434,N_14676,N_14493);
nor UO_1435 (O_1435,N_14326,N_14734);
xnor UO_1436 (O_1436,N_14301,N_14894);
nor UO_1437 (O_1437,N_14610,N_14576);
and UO_1438 (O_1438,N_14332,N_14814);
nor UO_1439 (O_1439,N_14870,N_14924);
xnor UO_1440 (O_1440,N_14309,N_14386);
xnor UO_1441 (O_1441,N_14735,N_14309);
or UO_1442 (O_1442,N_14926,N_14984);
nor UO_1443 (O_1443,N_14912,N_14675);
and UO_1444 (O_1444,N_14921,N_14549);
and UO_1445 (O_1445,N_14949,N_14547);
and UO_1446 (O_1446,N_14519,N_14817);
xor UO_1447 (O_1447,N_14382,N_14282);
xnor UO_1448 (O_1448,N_14390,N_14393);
or UO_1449 (O_1449,N_14716,N_14698);
nand UO_1450 (O_1450,N_14795,N_14546);
nor UO_1451 (O_1451,N_14928,N_14384);
and UO_1452 (O_1452,N_14353,N_14715);
and UO_1453 (O_1453,N_14711,N_14534);
or UO_1454 (O_1454,N_14618,N_14758);
xor UO_1455 (O_1455,N_14723,N_14566);
nand UO_1456 (O_1456,N_14681,N_14774);
and UO_1457 (O_1457,N_14417,N_14546);
and UO_1458 (O_1458,N_14999,N_14525);
nand UO_1459 (O_1459,N_14496,N_14345);
and UO_1460 (O_1460,N_14492,N_14808);
or UO_1461 (O_1461,N_14695,N_14724);
nor UO_1462 (O_1462,N_14569,N_14319);
xnor UO_1463 (O_1463,N_14448,N_14486);
nand UO_1464 (O_1464,N_14371,N_14923);
nor UO_1465 (O_1465,N_14642,N_14767);
xnor UO_1466 (O_1466,N_14411,N_14973);
and UO_1467 (O_1467,N_14902,N_14529);
nand UO_1468 (O_1468,N_14266,N_14310);
and UO_1469 (O_1469,N_14923,N_14912);
nand UO_1470 (O_1470,N_14856,N_14942);
and UO_1471 (O_1471,N_14982,N_14893);
and UO_1472 (O_1472,N_14650,N_14660);
or UO_1473 (O_1473,N_14721,N_14541);
nand UO_1474 (O_1474,N_14708,N_14981);
and UO_1475 (O_1475,N_14414,N_14595);
xnor UO_1476 (O_1476,N_14554,N_14689);
or UO_1477 (O_1477,N_14557,N_14993);
xnor UO_1478 (O_1478,N_14847,N_14308);
xnor UO_1479 (O_1479,N_14650,N_14489);
xnor UO_1480 (O_1480,N_14504,N_14925);
nor UO_1481 (O_1481,N_14657,N_14567);
nand UO_1482 (O_1482,N_14945,N_14473);
and UO_1483 (O_1483,N_14800,N_14632);
nor UO_1484 (O_1484,N_14826,N_14407);
xnor UO_1485 (O_1485,N_14872,N_14446);
xnor UO_1486 (O_1486,N_14852,N_14931);
nand UO_1487 (O_1487,N_14935,N_14803);
xnor UO_1488 (O_1488,N_14794,N_14784);
xnor UO_1489 (O_1489,N_14945,N_14664);
and UO_1490 (O_1490,N_14640,N_14656);
nand UO_1491 (O_1491,N_14687,N_14491);
xnor UO_1492 (O_1492,N_14585,N_14311);
nand UO_1493 (O_1493,N_14585,N_14829);
nor UO_1494 (O_1494,N_14337,N_14576);
xnor UO_1495 (O_1495,N_14911,N_14976);
nor UO_1496 (O_1496,N_14914,N_14862);
nand UO_1497 (O_1497,N_14375,N_14439);
nor UO_1498 (O_1498,N_14377,N_14572);
or UO_1499 (O_1499,N_14684,N_14339);
and UO_1500 (O_1500,N_14568,N_14423);
nand UO_1501 (O_1501,N_14496,N_14505);
xnor UO_1502 (O_1502,N_14869,N_14837);
or UO_1503 (O_1503,N_14690,N_14958);
nand UO_1504 (O_1504,N_14402,N_14607);
or UO_1505 (O_1505,N_14812,N_14960);
nand UO_1506 (O_1506,N_14805,N_14666);
or UO_1507 (O_1507,N_14321,N_14523);
xor UO_1508 (O_1508,N_14501,N_14396);
or UO_1509 (O_1509,N_14584,N_14388);
or UO_1510 (O_1510,N_14917,N_14992);
and UO_1511 (O_1511,N_14757,N_14845);
nor UO_1512 (O_1512,N_14905,N_14809);
xor UO_1513 (O_1513,N_14752,N_14744);
nor UO_1514 (O_1514,N_14867,N_14618);
nand UO_1515 (O_1515,N_14833,N_14748);
and UO_1516 (O_1516,N_14904,N_14457);
and UO_1517 (O_1517,N_14712,N_14987);
xor UO_1518 (O_1518,N_14981,N_14838);
nand UO_1519 (O_1519,N_14560,N_14954);
or UO_1520 (O_1520,N_14735,N_14442);
xnor UO_1521 (O_1521,N_14686,N_14542);
and UO_1522 (O_1522,N_14830,N_14697);
and UO_1523 (O_1523,N_14353,N_14920);
nand UO_1524 (O_1524,N_14972,N_14445);
nand UO_1525 (O_1525,N_14349,N_14397);
xor UO_1526 (O_1526,N_14860,N_14538);
xnor UO_1527 (O_1527,N_14758,N_14580);
xor UO_1528 (O_1528,N_14537,N_14911);
or UO_1529 (O_1529,N_14903,N_14500);
nor UO_1530 (O_1530,N_14363,N_14261);
nand UO_1531 (O_1531,N_14666,N_14296);
xnor UO_1532 (O_1532,N_14507,N_14285);
or UO_1533 (O_1533,N_14322,N_14259);
nor UO_1534 (O_1534,N_14731,N_14860);
and UO_1535 (O_1535,N_14419,N_14520);
xnor UO_1536 (O_1536,N_14627,N_14481);
xor UO_1537 (O_1537,N_14372,N_14510);
xor UO_1538 (O_1538,N_14681,N_14647);
xor UO_1539 (O_1539,N_14805,N_14714);
xnor UO_1540 (O_1540,N_14737,N_14758);
nand UO_1541 (O_1541,N_14611,N_14820);
nand UO_1542 (O_1542,N_14370,N_14664);
and UO_1543 (O_1543,N_14841,N_14878);
nand UO_1544 (O_1544,N_14752,N_14902);
or UO_1545 (O_1545,N_14279,N_14744);
and UO_1546 (O_1546,N_14500,N_14519);
and UO_1547 (O_1547,N_14867,N_14770);
xor UO_1548 (O_1548,N_14563,N_14566);
or UO_1549 (O_1549,N_14867,N_14601);
and UO_1550 (O_1550,N_14847,N_14938);
or UO_1551 (O_1551,N_14391,N_14515);
xor UO_1552 (O_1552,N_14661,N_14374);
nor UO_1553 (O_1553,N_14486,N_14978);
nor UO_1554 (O_1554,N_14341,N_14781);
or UO_1555 (O_1555,N_14594,N_14886);
and UO_1556 (O_1556,N_14398,N_14999);
nor UO_1557 (O_1557,N_14533,N_14643);
or UO_1558 (O_1558,N_14314,N_14644);
or UO_1559 (O_1559,N_14564,N_14691);
or UO_1560 (O_1560,N_14559,N_14867);
and UO_1561 (O_1561,N_14478,N_14638);
nand UO_1562 (O_1562,N_14375,N_14480);
nor UO_1563 (O_1563,N_14865,N_14740);
or UO_1564 (O_1564,N_14490,N_14830);
nor UO_1565 (O_1565,N_14726,N_14632);
xor UO_1566 (O_1566,N_14282,N_14558);
xnor UO_1567 (O_1567,N_14384,N_14395);
nand UO_1568 (O_1568,N_14677,N_14542);
and UO_1569 (O_1569,N_14453,N_14620);
or UO_1570 (O_1570,N_14437,N_14302);
or UO_1571 (O_1571,N_14386,N_14620);
nor UO_1572 (O_1572,N_14323,N_14854);
and UO_1573 (O_1573,N_14935,N_14382);
and UO_1574 (O_1574,N_14366,N_14351);
or UO_1575 (O_1575,N_14671,N_14890);
or UO_1576 (O_1576,N_14835,N_14358);
nor UO_1577 (O_1577,N_14339,N_14907);
or UO_1578 (O_1578,N_14509,N_14884);
or UO_1579 (O_1579,N_14827,N_14587);
xnor UO_1580 (O_1580,N_14613,N_14865);
or UO_1581 (O_1581,N_14324,N_14518);
or UO_1582 (O_1582,N_14390,N_14264);
and UO_1583 (O_1583,N_14515,N_14730);
nor UO_1584 (O_1584,N_14729,N_14623);
and UO_1585 (O_1585,N_14980,N_14491);
xnor UO_1586 (O_1586,N_14281,N_14435);
nor UO_1587 (O_1587,N_14855,N_14942);
nand UO_1588 (O_1588,N_14305,N_14723);
nand UO_1589 (O_1589,N_14428,N_14442);
nand UO_1590 (O_1590,N_14475,N_14620);
nand UO_1591 (O_1591,N_14718,N_14560);
or UO_1592 (O_1592,N_14716,N_14577);
nand UO_1593 (O_1593,N_14311,N_14729);
nand UO_1594 (O_1594,N_14313,N_14462);
or UO_1595 (O_1595,N_14790,N_14417);
nand UO_1596 (O_1596,N_14842,N_14269);
nand UO_1597 (O_1597,N_14427,N_14499);
xnor UO_1598 (O_1598,N_14454,N_14275);
and UO_1599 (O_1599,N_14885,N_14640);
xor UO_1600 (O_1600,N_14585,N_14297);
nand UO_1601 (O_1601,N_14311,N_14808);
or UO_1602 (O_1602,N_14323,N_14270);
and UO_1603 (O_1603,N_14489,N_14802);
and UO_1604 (O_1604,N_14917,N_14758);
and UO_1605 (O_1605,N_14766,N_14508);
nand UO_1606 (O_1606,N_14494,N_14673);
nor UO_1607 (O_1607,N_14519,N_14640);
nor UO_1608 (O_1608,N_14342,N_14356);
and UO_1609 (O_1609,N_14369,N_14781);
nor UO_1610 (O_1610,N_14379,N_14885);
xnor UO_1611 (O_1611,N_14355,N_14499);
xnor UO_1612 (O_1612,N_14252,N_14670);
nor UO_1613 (O_1613,N_14377,N_14380);
nor UO_1614 (O_1614,N_14428,N_14572);
and UO_1615 (O_1615,N_14890,N_14352);
xnor UO_1616 (O_1616,N_14820,N_14463);
nor UO_1617 (O_1617,N_14731,N_14494);
and UO_1618 (O_1618,N_14436,N_14472);
and UO_1619 (O_1619,N_14810,N_14394);
nor UO_1620 (O_1620,N_14819,N_14334);
nor UO_1621 (O_1621,N_14816,N_14891);
xnor UO_1622 (O_1622,N_14361,N_14760);
and UO_1623 (O_1623,N_14846,N_14873);
nor UO_1624 (O_1624,N_14766,N_14504);
nor UO_1625 (O_1625,N_14942,N_14485);
xor UO_1626 (O_1626,N_14541,N_14377);
xnor UO_1627 (O_1627,N_14513,N_14301);
xnor UO_1628 (O_1628,N_14259,N_14504);
xor UO_1629 (O_1629,N_14752,N_14905);
nand UO_1630 (O_1630,N_14988,N_14867);
xnor UO_1631 (O_1631,N_14890,N_14888);
or UO_1632 (O_1632,N_14842,N_14694);
nor UO_1633 (O_1633,N_14303,N_14308);
and UO_1634 (O_1634,N_14411,N_14959);
nor UO_1635 (O_1635,N_14437,N_14840);
nor UO_1636 (O_1636,N_14969,N_14315);
nand UO_1637 (O_1637,N_14588,N_14494);
or UO_1638 (O_1638,N_14468,N_14792);
and UO_1639 (O_1639,N_14335,N_14726);
and UO_1640 (O_1640,N_14430,N_14927);
and UO_1641 (O_1641,N_14727,N_14680);
and UO_1642 (O_1642,N_14263,N_14702);
nor UO_1643 (O_1643,N_14504,N_14734);
xnor UO_1644 (O_1644,N_14287,N_14968);
nand UO_1645 (O_1645,N_14986,N_14544);
or UO_1646 (O_1646,N_14282,N_14917);
xor UO_1647 (O_1647,N_14731,N_14978);
nor UO_1648 (O_1648,N_14475,N_14819);
nor UO_1649 (O_1649,N_14404,N_14583);
and UO_1650 (O_1650,N_14723,N_14386);
or UO_1651 (O_1651,N_14347,N_14396);
nand UO_1652 (O_1652,N_14406,N_14809);
xnor UO_1653 (O_1653,N_14865,N_14600);
nand UO_1654 (O_1654,N_14719,N_14930);
nand UO_1655 (O_1655,N_14880,N_14501);
xor UO_1656 (O_1656,N_14671,N_14303);
and UO_1657 (O_1657,N_14830,N_14258);
or UO_1658 (O_1658,N_14896,N_14864);
or UO_1659 (O_1659,N_14298,N_14596);
nand UO_1660 (O_1660,N_14628,N_14743);
or UO_1661 (O_1661,N_14566,N_14533);
or UO_1662 (O_1662,N_14578,N_14688);
xnor UO_1663 (O_1663,N_14403,N_14605);
and UO_1664 (O_1664,N_14790,N_14892);
xor UO_1665 (O_1665,N_14349,N_14776);
nor UO_1666 (O_1666,N_14844,N_14911);
or UO_1667 (O_1667,N_14263,N_14844);
nand UO_1668 (O_1668,N_14821,N_14944);
nand UO_1669 (O_1669,N_14350,N_14268);
nor UO_1670 (O_1670,N_14468,N_14571);
xor UO_1671 (O_1671,N_14477,N_14751);
nand UO_1672 (O_1672,N_14345,N_14896);
nand UO_1673 (O_1673,N_14773,N_14927);
nor UO_1674 (O_1674,N_14720,N_14573);
or UO_1675 (O_1675,N_14515,N_14285);
or UO_1676 (O_1676,N_14923,N_14525);
or UO_1677 (O_1677,N_14969,N_14513);
nand UO_1678 (O_1678,N_14906,N_14476);
nand UO_1679 (O_1679,N_14993,N_14695);
nor UO_1680 (O_1680,N_14535,N_14870);
and UO_1681 (O_1681,N_14633,N_14450);
nor UO_1682 (O_1682,N_14781,N_14610);
xor UO_1683 (O_1683,N_14933,N_14297);
and UO_1684 (O_1684,N_14539,N_14674);
nand UO_1685 (O_1685,N_14297,N_14771);
and UO_1686 (O_1686,N_14601,N_14317);
nor UO_1687 (O_1687,N_14821,N_14551);
xor UO_1688 (O_1688,N_14824,N_14817);
xnor UO_1689 (O_1689,N_14837,N_14711);
nor UO_1690 (O_1690,N_14658,N_14279);
or UO_1691 (O_1691,N_14553,N_14258);
nor UO_1692 (O_1692,N_14397,N_14890);
nand UO_1693 (O_1693,N_14305,N_14701);
xor UO_1694 (O_1694,N_14836,N_14639);
or UO_1695 (O_1695,N_14760,N_14260);
or UO_1696 (O_1696,N_14531,N_14279);
or UO_1697 (O_1697,N_14566,N_14406);
and UO_1698 (O_1698,N_14596,N_14978);
or UO_1699 (O_1699,N_14487,N_14552);
and UO_1700 (O_1700,N_14784,N_14711);
nor UO_1701 (O_1701,N_14428,N_14685);
nor UO_1702 (O_1702,N_14498,N_14711);
or UO_1703 (O_1703,N_14587,N_14636);
xor UO_1704 (O_1704,N_14325,N_14433);
xnor UO_1705 (O_1705,N_14870,N_14813);
and UO_1706 (O_1706,N_14650,N_14925);
and UO_1707 (O_1707,N_14330,N_14597);
nor UO_1708 (O_1708,N_14938,N_14550);
or UO_1709 (O_1709,N_14925,N_14597);
and UO_1710 (O_1710,N_14463,N_14811);
or UO_1711 (O_1711,N_14684,N_14580);
nand UO_1712 (O_1712,N_14727,N_14840);
nand UO_1713 (O_1713,N_14277,N_14731);
nor UO_1714 (O_1714,N_14970,N_14303);
and UO_1715 (O_1715,N_14701,N_14656);
nor UO_1716 (O_1716,N_14477,N_14868);
xor UO_1717 (O_1717,N_14767,N_14486);
nor UO_1718 (O_1718,N_14374,N_14496);
nor UO_1719 (O_1719,N_14999,N_14842);
nor UO_1720 (O_1720,N_14641,N_14395);
nor UO_1721 (O_1721,N_14812,N_14515);
or UO_1722 (O_1722,N_14526,N_14835);
nor UO_1723 (O_1723,N_14953,N_14362);
nor UO_1724 (O_1724,N_14751,N_14457);
nor UO_1725 (O_1725,N_14667,N_14346);
nor UO_1726 (O_1726,N_14579,N_14982);
nor UO_1727 (O_1727,N_14781,N_14444);
nor UO_1728 (O_1728,N_14552,N_14705);
nand UO_1729 (O_1729,N_14449,N_14404);
and UO_1730 (O_1730,N_14660,N_14308);
nand UO_1731 (O_1731,N_14336,N_14690);
or UO_1732 (O_1732,N_14700,N_14414);
nor UO_1733 (O_1733,N_14453,N_14687);
or UO_1734 (O_1734,N_14466,N_14893);
nor UO_1735 (O_1735,N_14280,N_14961);
nand UO_1736 (O_1736,N_14931,N_14327);
nand UO_1737 (O_1737,N_14473,N_14482);
or UO_1738 (O_1738,N_14396,N_14784);
xnor UO_1739 (O_1739,N_14705,N_14545);
nor UO_1740 (O_1740,N_14476,N_14520);
and UO_1741 (O_1741,N_14667,N_14940);
nand UO_1742 (O_1742,N_14577,N_14506);
xor UO_1743 (O_1743,N_14613,N_14383);
nand UO_1744 (O_1744,N_14794,N_14845);
nand UO_1745 (O_1745,N_14817,N_14809);
or UO_1746 (O_1746,N_14500,N_14587);
xnor UO_1747 (O_1747,N_14934,N_14286);
or UO_1748 (O_1748,N_14711,N_14401);
or UO_1749 (O_1749,N_14639,N_14398);
nand UO_1750 (O_1750,N_14921,N_14435);
xnor UO_1751 (O_1751,N_14988,N_14982);
and UO_1752 (O_1752,N_14281,N_14769);
nor UO_1753 (O_1753,N_14439,N_14844);
nor UO_1754 (O_1754,N_14816,N_14431);
or UO_1755 (O_1755,N_14873,N_14492);
nand UO_1756 (O_1756,N_14963,N_14806);
xnor UO_1757 (O_1757,N_14285,N_14627);
xnor UO_1758 (O_1758,N_14637,N_14714);
nand UO_1759 (O_1759,N_14467,N_14767);
and UO_1760 (O_1760,N_14569,N_14583);
and UO_1761 (O_1761,N_14861,N_14911);
nand UO_1762 (O_1762,N_14892,N_14924);
or UO_1763 (O_1763,N_14716,N_14272);
nor UO_1764 (O_1764,N_14800,N_14697);
nand UO_1765 (O_1765,N_14599,N_14740);
nand UO_1766 (O_1766,N_14708,N_14621);
xnor UO_1767 (O_1767,N_14728,N_14581);
or UO_1768 (O_1768,N_14594,N_14622);
or UO_1769 (O_1769,N_14895,N_14602);
nor UO_1770 (O_1770,N_14698,N_14739);
xnor UO_1771 (O_1771,N_14670,N_14319);
nor UO_1772 (O_1772,N_14443,N_14954);
nor UO_1773 (O_1773,N_14830,N_14451);
nor UO_1774 (O_1774,N_14722,N_14475);
or UO_1775 (O_1775,N_14620,N_14438);
nand UO_1776 (O_1776,N_14940,N_14530);
nand UO_1777 (O_1777,N_14562,N_14784);
and UO_1778 (O_1778,N_14455,N_14965);
or UO_1779 (O_1779,N_14610,N_14714);
nor UO_1780 (O_1780,N_14566,N_14937);
nor UO_1781 (O_1781,N_14418,N_14796);
xor UO_1782 (O_1782,N_14852,N_14662);
nand UO_1783 (O_1783,N_14625,N_14849);
nor UO_1784 (O_1784,N_14682,N_14485);
or UO_1785 (O_1785,N_14651,N_14902);
xnor UO_1786 (O_1786,N_14630,N_14572);
or UO_1787 (O_1787,N_14358,N_14670);
or UO_1788 (O_1788,N_14285,N_14366);
nand UO_1789 (O_1789,N_14387,N_14922);
or UO_1790 (O_1790,N_14848,N_14474);
xnor UO_1791 (O_1791,N_14753,N_14321);
nand UO_1792 (O_1792,N_14915,N_14928);
nor UO_1793 (O_1793,N_14853,N_14640);
nand UO_1794 (O_1794,N_14774,N_14657);
nor UO_1795 (O_1795,N_14534,N_14680);
or UO_1796 (O_1796,N_14729,N_14397);
nand UO_1797 (O_1797,N_14259,N_14667);
or UO_1798 (O_1798,N_14683,N_14762);
nand UO_1799 (O_1799,N_14729,N_14448);
nor UO_1800 (O_1800,N_14706,N_14460);
and UO_1801 (O_1801,N_14307,N_14910);
or UO_1802 (O_1802,N_14256,N_14689);
and UO_1803 (O_1803,N_14820,N_14937);
xor UO_1804 (O_1804,N_14448,N_14305);
and UO_1805 (O_1805,N_14569,N_14539);
xnor UO_1806 (O_1806,N_14480,N_14526);
nand UO_1807 (O_1807,N_14810,N_14555);
or UO_1808 (O_1808,N_14926,N_14725);
and UO_1809 (O_1809,N_14618,N_14708);
nand UO_1810 (O_1810,N_14394,N_14929);
or UO_1811 (O_1811,N_14472,N_14277);
or UO_1812 (O_1812,N_14401,N_14928);
xnor UO_1813 (O_1813,N_14455,N_14822);
or UO_1814 (O_1814,N_14870,N_14547);
and UO_1815 (O_1815,N_14918,N_14915);
or UO_1816 (O_1816,N_14664,N_14328);
nor UO_1817 (O_1817,N_14433,N_14740);
or UO_1818 (O_1818,N_14403,N_14776);
and UO_1819 (O_1819,N_14373,N_14425);
nand UO_1820 (O_1820,N_14645,N_14345);
and UO_1821 (O_1821,N_14298,N_14506);
nor UO_1822 (O_1822,N_14684,N_14358);
nand UO_1823 (O_1823,N_14422,N_14322);
or UO_1824 (O_1824,N_14925,N_14469);
and UO_1825 (O_1825,N_14511,N_14336);
and UO_1826 (O_1826,N_14320,N_14915);
and UO_1827 (O_1827,N_14551,N_14378);
nand UO_1828 (O_1828,N_14781,N_14992);
nor UO_1829 (O_1829,N_14378,N_14841);
nor UO_1830 (O_1830,N_14511,N_14809);
nand UO_1831 (O_1831,N_14532,N_14412);
xor UO_1832 (O_1832,N_14895,N_14708);
or UO_1833 (O_1833,N_14557,N_14708);
nor UO_1834 (O_1834,N_14775,N_14890);
nand UO_1835 (O_1835,N_14389,N_14697);
nand UO_1836 (O_1836,N_14912,N_14947);
xnor UO_1837 (O_1837,N_14618,N_14903);
nand UO_1838 (O_1838,N_14895,N_14529);
or UO_1839 (O_1839,N_14653,N_14785);
xnor UO_1840 (O_1840,N_14554,N_14854);
and UO_1841 (O_1841,N_14422,N_14537);
nor UO_1842 (O_1842,N_14368,N_14871);
or UO_1843 (O_1843,N_14322,N_14993);
or UO_1844 (O_1844,N_14467,N_14415);
nor UO_1845 (O_1845,N_14474,N_14705);
or UO_1846 (O_1846,N_14944,N_14714);
xor UO_1847 (O_1847,N_14495,N_14387);
or UO_1848 (O_1848,N_14814,N_14938);
xnor UO_1849 (O_1849,N_14349,N_14790);
xor UO_1850 (O_1850,N_14431,N_14674);
and UO_1851 (O_1851,N_14250,N_14857);
and UO_1852 (O_1852,N_14862,N_14806);
or UO_1853 (O_1853,N_14989,N_14975);
nor UO_1854 (O_1854,N_14783,N_14323);
or UO_1855 (O_1855,N_14849,N_14960);
xnor UO_1856 (O_1856,N_14564,N_14660);
xor UO_1857 (O_1857,N_14599,N_14607);
xor UO_1858 (O_1858,N_14915,N_14446);
xnor UO_1859 (O_1859,N_14364,N_14885);
xnor UO_1860 (O_1860,N_14419,N_14989);
nand UO_1861 (O_1861,N_14962,N_14589);
or UO_1862 (O_1862,N_14605,N_14797);
and UO_1863 (O_1863,N_14530,N_14462);
nand UO_1864 (O_1864,N_14592,N_14428);
nand UO_1865 (O_1865,N_14632,N_14674);
or UO_1866 (O_1866,N_14840,N_14702);
or UO_1867 (O_1867,N_14962,N_14894);
nor UO_1868 (O_1868,N_14354,N_14364);
nor UO_1869 (O_1869,N_14254,N_14456);
and UO_1870 (O_1870,N_14321,N_14888);
nand UO_1871 (O_1871,N_14651,N_14502);
nor UO_1872 (O_1872,N_14852,N_14810);
nand UO_1873 (O_1873,N_14316,N_14716);
or UO_1874 (O_1874,N_14278,N_14414);
nand UO_1875 (O_1875,N_14601,N_14629);
xnor UO_1876 (O_1876,N_14809,N_14575);
nand UO_1877 (O_1877,N_14296,N_14355);
and UO_1878 (O_1878,N_14836,N_14454);
nor UO_1879 (O_1879,N_14697,N_14404);
nand UO_1880 (O_1880,N_14665,N_14718);
nand UO_1881 (O_1881,N_14954,N_14970);
xnor UO_1882 (O_1882,N_14266,N_14498);
and UO_1883 (O_1883,N_14818,N_14795);
nand UO_1884 (O_1884,N_14970,N_14516);
xnor UO_1885 (O_1885,N_14758,N_14895);
nor UO_1886 (O_1886,N_14281,N_14523);
xor UO_1887 (O_1887,N_14372,N_14949);
and UO_1888 (O_1888,N_14772,N_14300);
xnor UO_1889 (O_1889,N_14972,N_14302);
and UO_1890 (O_1890,N_14338,N_14805);
and UO_1891 (O_1891,N_14333,N_14799);
nand UO_1892 (O_1892,N_14913,N_14746);
nand UO_1893 (O_1893,N_14688,N_14253);
nand UO_1894 (O_1894,N_14343,N_14942);
xnor UO_1895 (O_1895,N_14610,N_14298);
or UO_1896 (O_1896,N_14401,N_14309);
and UO_1897 (O_1897,N_14324,N_14765);
or UO_1898 (O_1898,N_14764,N_14539);
nor UO_1899 (O_1899,N_14913,N_14370);
xor UO_1900 (O_1900,N_14396,N_14887);
xor UO_1901 (O_1901,N_14793,N_14447);
nor UO_1902 (O_1902,N_14795,N_14389);
nor UO_1903 (O_1903,N_14915,N_14250);
nand UO_1904 (O_1904,N_14885,N_14578);
nor UO_1905 (O_1905,N_14711,N_14578);
nand UO_1906 (O_1906,N_14791,N_14837);
nor UO_1907 (O_1907,N_14739,N_14846);
and UO_1908 (O_1908,N_14472,N_14327);
xor UO_1909 (O_1909,N_14424,N_14790);
or UO_1910 (O_1910,N_14330,N_14253);
and UO_1911 (O_1911,N_14282,N_14414);
xnor UO_1912 (O_1912,N_14909,N_14544);
nand UO_1913 (O_1913,N_14566,N_14609);
nand UO_1914 (O_1914,N_14590,N_14858);
nor UO_1915 (O_1915,N_14611,N_14454);
xnor UO_1916 (O_1916,N_14634,N_14411);
and UO_1917 (O_1917,N_14857,N_14868);
nand UO_1918 (O_1918,N_14505,N_14276);
nand UO_1919 (O_1919,N_14470,N_14983);
and UO_1920 (O_1920,N_14339,N_14936);
and UO_1921 (O_1921,N_14940,N_14427);
nand UO_1922 (O_1922,N_14674,N_14750);
and UO_1923 (O_1923,N_14504,N_14720);
or UO_1924 (O_1924,N_14271,N_14387);
nand UO_1925 (O_1925,N_14338,N_14339);
or UO_1926 (O_1926,N_14908,N_14544);
nand UO_1927 (O_1927,N_14594,N_14465);
nor UO_1928 (O_1928,N_14638,N_14952);
nor UO_1929 (O_1929,N_14675,N_14941);
or UO_1930 (O_1930,N_14479,N_14806);
nor UO_1931 (O_1931,N_14998,N_14396);
and UO_1932 (O_1932,N_14705,N_14960);
and UO_1933 (O_1933,N_14826,N_14749);
nor UO_1934 (O_1934,N_14258,N_14734);
or UO_1935 (O_1935,N_14838,N_14913);
and UO_1936 (O_1936,N_14934,N_14298);
xnor UO_1937 (O_1937,N_14979,N_14937);
and UO_1938 (O_1938,N_14409,N_14837);
nor UO_1939 (O_1939,N_14308,N_14644);
or UO_1940 (O_1940,N_14438,N_14775);
nor UO_1941 (O_1941,N_14260,N_14658);
and UO_1942 (O_1942,N_14676,N_14591);
and UO_1943 (O_1943,N_14815,N_14657);
or UO_1944 (O_1944,N_14441,N_14419);
nand UO_1945 (O_1945,N_14791,N_14257);
xor UO_1946 (O_1946,N_14689,N_14378);
nand UO_1947 (O_1947,N_14955,N_14446);
xor UO_1948 (O_1948,N_14369,N_14372);
or UO_1949 (O_1949,N_14973,N_14626);
nor UO_1950 (O_1950,N_14350,N_14858);
xnor UO_1951 (O_1951,N_14585,N_14902);
or UO_1952 (O_1952,N_14855,N_14388);
or UO_1953 (O_1953,N_14527,N_14497);
or UO_1954 (O_1954,N_14791,N_14454);
nand UO_1955 (O_1955,N_14562,N_14301);
or UO_1956 (O_1956,N_14503,N_14635);
nor UO_1957 (O_1957,N_14744,N_14503);
nor UO_1958 (O_1958,N_14621,N_14335);
and UO_1959 (O_1959,N_14842,N_14572);
or UO_1960 (O_1960,N_14367,N_14648);
nand UO_1961 (O_1961,N_14677,N_14303);
nand UO_1962 (O_1962,N_14411,N_14305);
or UO_1963 (O_1963,N_14356,N_14532);
and UO_1964 (O_1964,N_14838,N_14576);
and UO_1965 (O_1965,N_14971,N_14364);
nor UO_1966 (O_1966,N_14774,N_14387);
nor UO_1967 (O_1967,N_14285,N_14874);
nand UO_1968 (O_1968,N_14598,N_14814);
or UO_1969 (O_1969,N_14641,N_14680);
or UO_1970 (O_1970,N_14763,N_14337);
nand UO_1971 (O_1971,N_14710,N_14499);
nand UO_1972 (O_1972,N_14519,N_14711);
and UO_1973 (O_1973,N_14869,N_14789);
and UO_1974 (O_1974,N_14743,N_14342);
xnor UO_1975 (O_1975,N_14310,N_14820);
or UO_1976 (O_1976,N_14264,N_14718);
xor UO_1977 (O_1977,N_14544,N_14754);
and UO_1978 (O_1978,N_14297,N_14272);
nor UO_1979 (O_1979,N_14296,N_14604);
nand UO_1980 (O_1980,N_14466,N_14551);
nor UO_1981 (O_1981,N_14293,N_14740);
and UO_1982 (O_1982,N_14410,N_14377);
nand UO_1983 (O_1983,N_14691,N_14912);
xor UO_1984 (O_1984,N_14632,N_14712);
xor UO_1985 (O_1985,N_14591,N_14324);
or UO_1986 (O_1986,N_14591,N_14478);
nand UO_1987 (O_1987,N_14702,N_14658);
xor UO_1988 (O_1988,N_14374,N_14943);
xnor UO_1989 (O_1989,N_14851,N_14712);
or UO_1990 (O_1990,N_14413,N_14589);
xor UO_1991 (O_1991,N_14307,N_14950);
and UO_1992 (O_1992,N_14288,N_14516);
xor UO_1993 (O_1993,N_14736,N_14445);
nand UO_1994 (O_1994,N_14417,N_14676);
and UO_1995 (O_1995,N_14624,N_14999);
and UO_1996 (O_1996,N_14642,N_14625);
xor UO_1997 (O_1997,N_14564,N_14373);
nor UO_1998 (O_1998,N_14599,N_14928);
xnor UO_1999 (O_1999,N_14701,N_14499);
endmodule