module basic_500_3000_500_5_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_241,In_15);
nor U1 (N_1,In_291,In_26);
nand U2 (N_2,In_168,In_94);
nor U3 (N_3,In_471,In_452);
nor U4 (N_4,In_32,In_275);
and U5 (N_5,In_423,In_104);
or U6 (N_6,In_135,In_404);
or U7 (N_7,In_432,In_157);
xnor U8 (N_8,In_303,In_105);
and U9 (N_9,In_220,In_391);
or U10 (N_10,In_162,In_92);
or U11 (N_11,In_328,In_193);
or U12 (N_12,In_8,In_444);
nand U13 (N_13,In_289,In_447);
nor U14 (N_14,In_224,In_167);
and U15 (N_15,In_232,In_258);
nand U16 (N_16,In_468,In_302);
or U17 (N_17,In_3,In_312);
and U18 (N_18,In_424,In_440);
or U19 (N_19,In_309,In_201);
nand U20 (N_20,In_495,In_427);
or U21 (N_21,In_407,In_112);
and U22 (N_22,In_142,In_208);
nor U23 (N_23,In_465,In_421);
and U24 (N_24,In_487,In_307);
nor U25 (N_25,In_172,In_60);
nand U26 (N_26,In_82,In_405);
or U27 (N_27,In_90,In_344);
and U28 (N_28,In_39,In_20);
nand U29 (N_29,In_207,In_107);
and U30 (N_30,In_229,In_349);
and U31 (N_31,In_66,In_70);
and U32 (N_32,In_326,In_223);
and U33 (N_33,In_446,In_370);
nor U34 (N_34,In_438,In_246);
nor U35 (N_35,In_261,In_273);
nand U36 (N_36,In_81,In_377);
or U37 (N_37,In_422,In_170);
nor U38 (N_38,In_247,In_33);
and U39 (N_39,In_319,In_325);
or U40 (N_40,In_433,In_79);
nor U41 (N_41,In_151,In_88);
nand U42 (N_42,In_496,In_351);
and U43 (N_43,In_233,In_57);
and U44 (N_44,In_282,In_97);
xnor U45 (N_45,In_491,In_323);
nand U46 (N_46,In_91,In_279);
nand U47 (N_47,In_205,In_346);
nor U48 (N_48,In_359,In_478);
nand U49 (N_49,In_74,In_454);
nand U50 (N_50,In_86,In_479);
and U51 (N_51,In_296,In_362);
or U52 (N_52,In_24,In_47);
nand U53 (N_53,In_357,In_131);
and U54 (N_54,In_249,In_69);
nand U55 (N_55,In_149,In_330);
and U56 (N_56,In_462,In_467);
and U57 (N_57,In_485,In_191);
nand U58 (N_58,In_59,In_31);
nand U59 (N_59,In_222,In_83);
or U60 (N_60,In_281,In_25);
nor U61 (N_61,In_98,In_400);
nor U62 (N_62,In_499,In_40);
or U63 (N_63,In_408,In_434);
nor U64 (N_64,In_458,In_295);
or U65 (N_65,In_160,In_431);
or U66 (N_66,In_173,In_480);
or U67 (N_67,In_276,In_410);
and U68 (N_68,In_129,In_451);
nand U69 (N_69,In_198,In_445);
nand U70 (N_70,In_363,In_403);
and U71 (N_71,In_235,In_228);
or U72 (N_72,In_381,In_277);
or U73 (N_73,In_484,In_498);
nor U74 (N_74,In_383,In_337);
nor U75 (N_75,In_417,In_293);
or U76 (N_76,In_67,In_287);
or U77 (N_77,In_304,In_199);
and U78 (N_78,In_350,In_269);
or U79 (N_79,In_213,In_290);
or U80 (N_80,In_9,In_30);
nand U81 (N_81,In_270,In_76);
nand U82 (N_82,In_230,In_285);
nor U83 (N_83,In_119,In_243);
and U84 (N_84,In_126,In_211);
nand U85 (N_85,In_202,In_414);
nor U86 (N_86,In_14,In_196);
and U87 (N_87,In_415,In_128);
nand U88 (N_88,In_392,In_368);
nand U89 (N_89,In_150,In_192);
and U90 (N_90,In_85,In_159);
and U91 (N_91,In_371,In_45);
or U92 (N_92,In_475,In_113);
nor U93 (N_93,In_103,In_360);
or U94 (N_94,In_41,In_437);
or U95 (N_95,In_19,In_148);
or U96 (N_96,In_55,In_308);
and U97 (N_97,In_358,In_146);
and U98 (N_98,In_65,In_34);
nand U99 (N_99,In_221,In_464);
nor U100 (N_100,In_286,In_143);
nand U101 (N_101,In_42,In_239);
nor U102 (N_102,In_481,In_382);
nand U103 (N_103,In_5,In_38);
or U104 (N_104,In_367,In_189);
and U105 (N_105,In_152,In_0);
nand U106 (N_106,In_372,In_137);
nor U107 (N_107,In_430,In_18);
nor U108 (N_108,In_399,In_395);
nand U109 (N_109,In_118,In_340);
nor U110 (N_110,In_324,In_334);
and U111 (N_111,In_322,In_29);
nand U112 (N_112,In_166,In_35);
or U113 (N_113,In_178,In_457);
nor U114 (N_114,In_343,In_190);
xor U115 (N_115,In_95,In_409);
nor U116 (N_116,In_71,In_316);
and U117 (N_117,In_78,In_387);
or U118 (N_118,In_96,In_390);
nand U119 (N_119,In_268,In_215);
nor U120 (N_120,In_297,In_265);
or U121 (N_121,In_298,In_206);
nand U122 (N_122,In_188,In_393);
or U123 (N_123,In_251,In_255);
nor U124 (N_124,In_183,In_155);
or U125 (N_125,In_317,In_10);
or U126 (N_126,In_280,In_428);
and U127 (N_127,In_182,In_210);
or U128 (N_128,In_436,In_163);
or U129 (N_129,In_102,In_244);
and U130 (N_130,In_347,In_306);
or U131 (N_131,In_419,In_466);
or U132 (N_132,In_16,In_353);
and U133 (N_133,In_176,In_375);
or U134 (N_134,In_1,In_490);
or U135 (N_135,In_448,In_355);
or U136 (N_136,In_51,In_388);
and U137 (N_137,In_154,In_299);
or U138 (N_138,In_420,In_219);
nor U139 (N_139,In_473,In_68);
and U140 (N_140,In_218,In_169);
and U141 (N_141,In_292,In_6);
nor U142 (N_142,In_109,In_234);
nand U143 (N_143,In_122,In_214);
or U144 (N_144,In_185,In_379);
nor U145 (N_145,In_242,In_385);
or U146 (N_146,In_314,In_352);
and U147 (N_147,In_333,In_127);
nor U148 (N_148,In_426,In_58);
nor U149 (N_149,In_124,In_411);
nand U150 (N_150,In_418,In_116);
nor U151 (N_151,In_46,In_470);
or U152 (N_152,In_364,In_175);
and U153 (N_153,In_144,In_141);
or U154 (N_154,In_61,In_469);
nand U155 (N_155,In_378,In_177);
and U156 (N_156,In_413,In_460);
nand U157 (N_157,In_310,In_386);
nor U158 (N_158,In_187,In_216);
nand U159 (N_159,In_402,In_483);
and U160 (N_160,In_398,In_138);
nand U161 (N_161,In_256,In_361);
nor U162 (N_162,In_331,In_301);
or U163 (N_163,In_89,In_4);
or U164 (N_164,In_266,In_194);
and U165 (N_165,In_477,In_227);
and U166 (N_166,In_87,In_27);
and U167 (N_167,In_72,In_133);
and U168 (N_168,In_369,In_7);
and U169 (N_169,In_130,In_373);
nor U170 (N_170,In_260,In_474);
or U171 (N_171,In_153,In_114);
and U172 (N_172,In_264,In_453);
or U173 (N_173,In_75,In_99);
nor U174 (N_174,In_139,In_132);
nand U175 (N_175,In_165,In_376);
or U176 (N_176,In_455,In_401);
nor U177 (N_177,In_184,In_108);
and U178 (N_178,In_121,In_225);
nor U179 (N_179,In_494,In_226);
nand U180 (N_180,In_488,In_125);
nand U181 (N_181,In_311,In_12);
or U182 (N_182,In_44,In_62);
and U183 (N_183,In_472,In_283);
nand U184 (N_184,In_212,In_406);
or U185 (N_185,In_240,In_456);
nor U186 (N_186,In_63,In_238);
nor U187 (N_187,In_52,In_73);
nor U188 (N_188,In_435,In_449);
nor U189 (N_189,In_332,In_267);
and U190 (N_190,In_374,In_80);
or U191 (N_191,In_342,In_272);
or U192 (N_192,In_197,In_93);
or U193 (N_193,In_294,In_259);
nand U194 (N_194,In_22,In_305);
and U195 (N_195,In_134,In_11);
or U196 (N_196,In_237,In_315);
and U197 (N_197,In_443,In_100);
nor U198 (N_198,In_339,In_425);
and U199 (N_199,In_476,In_356);
or U200 (N_200,In_48,In_106);
or U201 (N_201,In_110,In_120);
or U202 (N_202,In_253,In_140);
and U203 (N_203,In_156,In_313);
or U204 (N_204,In_231,In_365);
and U205 (N_205,In_396,In_348);
nor U206 (N_206,In_248,In_145);
and U207 (N_207,In_50,In_461);
and U208 (N_208,In_397,In_257);
and U209 (N_209,In_123,In_200);
nand U210 (N_210,In_380,In_254);
and U211 (N_211,In_56,In_262);
nor U212 (N_212,In_336,In_53);
and U213 (N_213,In_497,In_329);
nor U214 (N_214,In_463,In_174);
or U215 (N_215,In_17,In_493);
nor U216 (N_216,In_389,In_441);
and U217 (N_217,In_49,In_318);
xnor U218 (N_218,In_204,In_450);
nand U219 (N_219,In_136,In_271);
nand U220 (N_220,In_288,In_37);
or U221 (N_221,In_245,In_320);
or U222 (N_222,In_416,In_64);
and U223 (N_223,In_263,In_161);
or U224 (N_224,In_23,In_217);
or U225 (N_225,In_36,In_321);
nand U226 (N_226,In_21,In_345);
nor U227 (N_227,In_338,In_442);
nand U228 (N_228,In_439,In_250);
and U229 (N_229,In_28,In_354);
or U230 (N_230,In_186,In_164);
and U231 (N_231,In_77,In_195);
and U232 (N_232,In_278,In_492);
nand U233 (N_233,In_84,In_274);
or U234 (N_234,In_486,In_327);
nor U235 (N_235,In_341,In_384);
and U236 (N_236,In_180,In_284);
or U237 (N_237,In_489,In_366);
nand U238 (N_238,In_147,In_171);
nor U239 (N_239,In_203,In_300);
and U240 (N_240,In_179,In_2);
nand U241 (N_241,In_54,In_43);
or U242 (N_242,In_459,In_181);
or U243 (N_243,In_101,In_13);
or U244 (N_244,In_236,In_429);
nand U245 (N_245,In_117,In_335);
nor U246 (N_246,In_158,In_394);
nand U247 (N_247,In_209,In_111);
nor U248 (N_248,In_412,In_252);
nor U249 (N_249,In_482,In_115);
or U250 (N_250,In_6,In_210);
nor U251 (N_251,In_16,In_360);
or U252 (N_252,In_371,In_187);
nor U253 (N_253,In_177,In_311);
nor U254 (N_254,In_76,In_445);
and U255 (N_255,In_110,In_480);
and U256 (N_256,In_294,In_141);
nor U257 (N_257,In_203,In_198);
nand U258 (N_258,In_418,In_497);
nand U259 (N_259,In_195,In_67);
and U260 (N_260,In_496,In_366);
or U261 (N_261,In_52,In_172);
and U262 (N_262,In_365,In_100);
and U263 (N_263,In_113,In_317);
and U264 (N_264,In_282,In_23);
nand U265 (N_265,In_64,In_488);
nand U266 (N_266,In_313,In_354);
nand U267 (N_267,In_464,In_219);
or U268 (N_268,In_151,In_166);
nand U269 (N_269,In_448,In_195);
nand U270 (N_270,In_44,In_138);
and U271 (N_271,In_138,In_232);
nand U272 (N_272,In_206,In_212);
nand U273 (N_273,In_228,In_193);
or U274 (N_274,In_33,In_303);
nand U275 (N_275,In_111,In_432);
and U276 (N_276,In_475,In_308);
and U277 (N_277,In_218,In_253);
or U278 (N_278,In_193,In_454);
or U279 (N_279,In_2,In_303);
and U280 (N_280,In_128,In_184);
and U281 (N_281,In_465,In_114);
nand U282 (N_282,In_293,In_236);
nor U283 (N_283,In_17,In_299);
nor U284 (N_284,In_479,In_431);
or U285 (N_285,In_156,In_494);
or U286 (N_286,In_461,In_468);
nor U287 (N_287,In_437,In_60);
or U288 (N_288,In_391,In_288);
and U289 (N_289,In_288,In_3);
nand U290 (N_290,In_219,In_427);
nor U291 (N_291,In_392,In_143);
or U292 (N_292,In_83,In_252);
and U293 (N_293,In_234,In_293);
or U294 (N_294,In_474,In_1);
or U295 (N_295,In_41,In_195);
or U296 (N_296,In_66,In_359);
nand U297 (N_297,In_463,In_76);
nor U298 (N_298,In_198,In_325);
nand U299 (N_299,In_474,In_241);
nand U300 (N_300,In_144,In_24);
nand U301 (N_301,In_63,In_220);
nand U302 (N_302,In_261,In_178);
nand U303 (N_303,In_340,In_484);
or U304 (N_304,In_198,In_183);
nand U305 (N_305,In_297,In_270);
nor U306 (N_306,In_477,In_201);
nor U307 (N_307,In_336,In_152);
and U308 (N_308,In_333,In_420);
nor U309 (N_309,In_111,In_189);
nor U310 (N_310,In_137,In_58);
nor U311 (N_311,In_471,In_494);
nand U312 (N_312,In_292,In_43);
and U313 (N_313,In_274,In_52);
nand U314 (N_314,In_139,In_123);
nand U315 (N_315,In_492,In_462);
and U316 (N_316,In_369,In_402);
nand U317 (N_317,In_137,In_25);
nor U318 (N_318,In_139,In_146);
and U319 (N_319,In_384,In_37);
and U320 (N_320,In_446,In_226);
nand U321 (N_321,In_370,In_196);
or U322 (N_322,In_247,In_213);
nor U323 (N_323,In_358,In_63);
and U324 (N_324,In_114,In_73);
and U325 (N_325,In_265,In_440);
nand U326 (N_326,In_396,In_387);
nor U327 (N_327,In_379,In_439);
nand U328 (N_328,In_459,In_276);
nand U329 (N_329,In_16,In_209);
nand U330 (N_330,In_172,In_294);
and U331 (N_331,In_438,In_19);
nor U332 (N_332,In_328,In_438);
or U333 (N_333,In_54,In_180);
or U334 (N_334,In_290,In_420);
or U335 (N_335,In_189,In_337);
and U336 (N_336,In_186,In_400);
nand U337 (N_337,In_23,In_234);
or U338 (N_338,In_40,In_80);
and U339 (N_339,In_185,In_463);
and U340 (N_340,In_420,In_426);
nand U341 (N_341,In_355,In_99);
and U342 (N_342,In_378,In_195);
nand U343 (N_343,In_302,In_254);
nand U344 (N_344,In_446,In_163);
and U345 (N_345,In_181,In_432);
nor U346 (N_346,In_34,In_446);
and U347 (N_347,In_232,In_349);
nor U348 (N_348,In_334,In_463);
and U349 (N_349,In_396,In_320);
and U350 (N_350,In_218,In_382);
nor U351 (N_351,In_204,In_136);
or U352 (N_352,In_399,In_4);
and U353 (N_353,In_79,In_9);
nor U354 (N_354,In_83,In_394);
and U355 (N_355,In_319,In_226);
nor U356 (N_356,In_237,In_288);
nand U357 (N_357,In_363,In_381);
and U358 (N_358,In_498,In_367);
and U359 (N_359,In_92,In_488);
and U360 (N_360,In_108,In_154);
or U361 (N_361,In_343,In_42);
and U362 (N_362,In_251,In_98);
nor U363 (N_363,In_365,In_275);
or U364 (N_364,In_118,In_105);
nor U365 (N_365,In_120,In_426);
and U366 (N_366,In_121,In_446);
nor U367 (N_367,In_276,In_389);
and U368 (N_368,In_475,In_122);
nor U369 (N_369,In_231,In_300);
and U370 (N_370,In_105,In_264);
or U371 (N_371,In_374,In_393);
and U372 (N_372,In_307,In_54);
nor U373 (N_373,In_140,In_309);
or U374 (N_374,In_438,In_178);
nor U375 (N_375,In_429,In_404);
or U376 (N_376,In_16,In_69);
and U377 (N_377,In_484,In_7);
nor U378 (N_378,In_49,In_119);
or U379 (N_379,In_444,In_255);
or U380 (N_380,In_344,In_446);
and U381 (N_381,In_341,In_151);
nand U382 (N_382,In_340,In_413);
and U383 (N_383,In_56,In_228);
nor U384 (N_384,In_49,In_102);
xnor U385 (N_385,In_249,In_100);
or U386 (N_386,In_498,In_236);
or U387 (N_387,In_98,In_263);
and U388 (N_388,In_98,In_304);
nand U389 (N_389,In_115,In_483);
nand U390 (N_390,In_71,In_394);
and U391 (N_391,In_323,In_133);
and U392 (N_392,In_193,In_198);
and U393 (N_393,In_379,In_328);
nor U394 (N_394,In_198,In_177);
or U395 (N_395,In_52,In_491);
nor U396 (N_396,In_418,In_154);
nand U397 (N_397,In_102,In_458);
or U398 (N_398,In_106,In_304);
or U399 (N_399,In_155,In_195);
nand U400 (N_400,In_158,In_443);
nor U401 (N_401,In_110,In_376);
and U402 (N_402,In_322,In_20);
nand U403 (N_403,In_23,In_433);
or U404 (N_404,In_206,In_401);
nor U405 (N_405,In_357,In_31);
nor U406 (N_406,In_33,In_177);
and U407 (N_407,In_21,In_238);
nand U408 (N_408,In_277,In_251);
nand U409 (N_409,In_100,In_488);
and U410 (N_410,In_392,In_266);
nor U411 (N_411,In_200,In_3);
and U412 (N_412,In_338,In_391);
or U413 (N_413,In_60,In_199);
and U414 (N_414,In_381,In_327);
nand U415 (N_415,In_176,In_302);
or U416 (N_416,In_256,In_9);
and U417 (N_417,In_470,In_251);
nor U418 (N_418,In_311,In_178);
or U419 (N_419,In_170,In_344);
or U420 (N_420,In_221,In_206);
and U421 (N_421,In_260,In_16);
nand U422 (N_422,In_309,In_25);
and U423 (N_423,In_273,In_287);
nor U424 (N_424,In_308,In_237);
nand U425 (N_425,In_75,In_352);
nor U426 (N_426,In_68,In_7);
nor U427 (N_427,In_191,In_480);
nand U428 (N_428,In_261,In_391);
nand U429 (N_429,In_465,In_456);
or U430 (N_430,In_490,In_211);
nor U431 (N_431,In_316,In_286);
and U432 (N_432,In_46,In_237);
and U433 (N_433,In_321,In_467);
nand U434 (N_434,In_418,In_380);
nand U435 (N_435,In_186,In_71);
or U436 (N_436,In_420,In_385);
and U437 (N_437,In_42,In_352);
nor U438 (N_438,In_68,In_35);
and U439 (N_439,In_474,In_434);
nand U440 (N_440,In_340,In_201);
or U441 (N_441,In_7,In_220);
nor U442 (N_442,In_379,In_8);
nor U443 (N_443,In_156,In_322);
nand U444 (N_444,In_343,In_485);
nor U445 (N_445,In_1,In_381);
or U446 (N_446,In_378,In_21);
or U447 (N_447,In_185,In_283);
xor U448 (N_448,In_460,In_296);
nor U449 (N_449,In_449,In_28);
and U450 (N_450,In_152,In_308);
nand U451 (N_451,In_209,In_91);
or U452 (N_452,In_112,In_97);
or U453 (N_453,In_171,In_495);
nor U454 (N_454,In_427,In_392);
nand U455 (N_455,In_324,In_353);
and U456 (N_456,In_250,In_129);
nand U457 (N_457,In_398,In_370);
and U458 (N_458,In_248,In_446);
nor U459 (N_459,In_324,In_4);
nor U460 (N_460,In_13,In_367);
nor U461 (N_461,In_204,In_260);
nor U462 (N_462,In_278,In_355);
nand U463 (N_463,In_445,In_382);
nor U464 (N_464,In_472,In_222);
and U465 (N_465,In_175,In_113);
or U466 (N_466,In_331,In_350);
or U467 (N_467,In_39,In_132);
and U468 (N_468,In_7,In_164);
nor U469 (N_469,In_187,In_421);
and U470 (N_470,In_471,In_365);
nand U471 (N_471,In_320,In_95);
or U472 (N_472,In_358,In_96);
nand U473 (N_473,In_477,In_455);
nor U474 (N_474,In_135,In_465);
and U475 (N_475,In_213,In_437);
or U476 (N_476,In_3,In_366);
nor U477 (N_477,In_143,In_57);
or U478 (N_478,In_406,In_6);
nor U479 (N_479,In_201,In_324);
or U480 (N_480,In_219,In_201);
nand U481 (N_481,In_452,In_225);
nor U482 (N_482,In_317,In_107);
nor U483 (N_483,In_87,In_25);
nand U484 (N_484,In_445,In_136);
or U485 (N_485,In_129,In_458);
and U486 (N_486,In_244,In_110);
or U487 (N_487,In_5,In_308);
nor U488 (N_488,In_439,In_348);
nand U489 (N_489,In_259,In_277);
or U490 (N_490,In_153,In_271);
and U491 (N_491,In_168,In_494);
and U492 (N_492,In_239,In_443);
and U493 (N_493,In_66,In_122);
nor U494 (N_494,In_329,In_420);
nor U495 (N_495,In_463,In_128);
or U496 (N_496,In_131,In_97);
nor U497 (N_497,In_377,In_230);
nor U498 (N_498,In_167,In_168);
or U499 (N_499,In_423,In_214);
nor U500 (N_500,In_43,In_499);
nor U501 (N_501,In_466,In_359);
nor U502 (N_502,In_172,In_410);
and U503 (N_503,In_311,In_114);
nor U504 (N_504,In_2,In_17);
or U505 (N_505,In_175,In_360);
or U506 (N_506,In_274,In_148);
nand U507 (N_507,In_462,In_36);
and U508 (N_508,In_123,In_91);
and U509 (N_509,In_312,In_185);
and U510 (N_510,In_465,In_499);
nand U511 (N_511,In_92,In_220);
and U512 (N_512,In_44,In_473);
nor U513 (N_513,In_97,In_325);
nand U514 (N_514,In_331,In_20);
xor U515 (N_515,In_86,In_124);
or U516 (N_516,In_377,In_425);
and U517 (N_517,In_27,In_190);
nor U518 (N_518,In_407,In_167);
nand U519 (N_519,In_428,In_138);
or U520 (N_520,In_329,In_343);
and U521 (N_521,In_283,In_359);
and U522 (N_522,In_145,In_356);
nand U523 (N_523,In_132,In_329);
and U524 (N_524,In_477,In_281);
and U525 (N_525,In_294,In_430);
nand U526 (N_526,In_64,In_494);
and U527 (N_527,In_50,In_480);
nand U528 (N_528,In_492,In_456);
nand U529 (N_529,In_189,In_159);
nor U530 (N_530,In_294,In_158);
nand U531 (N_531,In_338,In_135);
and U532 (N_532,In_115,In_338);
or U533 (N_533,In_254,In_439);
nor U534 (N_534,In_160,In_248);
xor U535 (N_535,In_469,In_232);
nor U536 (N_536,In_483,In_463);
nand U537 (N_537,In_323,In_467);
nor U538 (N_538,In_323,In_465);
or U539 (N_539,In_439,In_488);
and U540 (N_540,In_463,In_57);
and U541 (N_541,In_96,In_209);
nand U542 (N_542,In_137,In_290);
xnor U543 (N_543,In_207,In_142);
nand U544 (N_544,In_90,In_375);
and U545 (N_545,In_109,In_437);
nor U546 (N_546,In_8,In_351);
or U547 (N_547,In_386,In_266);
and U548 (N_548,In_86,In_4);
or U549 (N_549,In_341,In_95);
or U550 (N_550,In_51,In_486);
or U551 (N_551,In_497,In_415);
nor U552 (N_552,In_471,In_41);
and U553 (N_553,In_86,In_288);
or U554 (N_554,In_478,In_10);
or U555 (N_555,In_295,In_411);
or U556 (N_556,In_265,In_474);
nand U557 (N_557,In_135,In_241);
and U558 (N_558,In_265,In_12);
nor U559 (N_559,In_312,In_130);
and U560 (N_560,In_256,In_486);
nand U561 (N_561,In_305,In_155);
nand U562 (N_562,In_429,In_112);
nand U563 (N_563,In_340,In_422);
or U564 (N_564,In_250,In_301);
or U565 (N_565,In_469,In_171);
nor U566 (N_566,In_476,In_472);
nor U567 (N_567,In_86,In_145);
nand U568 (N_568,In_334,In_428);
or U569 (N_569,In_278,In_360);
nand U570 (N_570,In_183,In_158);
or U571 (N_571,In_233,In_167);
or U572 (N_572,In_79,In_479);
nand U573 (N_573,In_298,In_329);
nor U574 (N_574,In_401,In_166);
nor U575 (N_575,In_422,In_23);
nand U576 (N_576,In_353,In_87);
nor U577 (N_577,In_165,In_307);
nand U578 (N_578,In_55,In_402);
nand U579 (N_579,In_183,In_161);
nor U580 (N_580,In_222,In_164);
nand U581 (N_581,In_223,In_232);
or U582 (N_582,In_80,In_342);
and U583 (N_583,In_250,In_36);
nor U584 (N_584,In_252,In_376);
or U585 (N_585,In_488,In_7);
nor U586 (N_586,In_327,In_417);
and U587 (N_587,In_408,In_420);
or U588 (N_588,In_220,In_202);
nor U589 (N_589,In_131,In_454);
and U590 (N_590,In_116,In_287);
or U591 (N_591,In_412,In_392);
nand U592 (N_592,In_167,In_303);
and U593 (N_593,In_370,In_122);
nor U594 (N_594,In_432,In_241);
and U595 (N_595,In_184,In_426);
and U596 (N_596,In_272,In_430);
and U597 (N_597,In_437,In_230);
and U598 (N_598,In_235,In_418);
nand U599 (N_599,In_198,In_143);
and U600 (N_600,N_280,N_135);
or U601 (N_601,N_564,N_346);
and U602 (N_602,N_490,N_26);
nand U603 (N_603,N_151,N_279);
nand U604 (N_604,N_494,N_202);
nor U605 (N_605,N_464,N_77);
or U606 (N_606,N_304,N_283);
nor U607 (N_607,N_259,N_446);
nand U608 (N_608,N_595,N_542);
nor U609 (N_609,N_502,N_261);
nand U610 (N_610,N_398,N_404);
and U611 (N_611,N_530,N_253);
and U612 (N_612,N_399,N_84);
nand U613 (N_613,N_110,N_289);
or U614 (N_614,N_303,N_332);
and U615 (N_615,N_80,N_563);
nor U616 (N_616,N_256,N_411);
and U617 (N_617,N_277,N_192);
or U618 (N_618,N_162,N_52);
nand U619 (N_619,N_394,N_248);
nand U620 (N_620,N_267,N_87);
nand U621 (N_621,N_72,N_90);
and U622 (N_622,N_217,N_58);
and U623 (N_623,N_353,N_104);
or U624 (N_624,N_526,N_426);
and U625 (N_625,N_462,N_10);
or U626 (N_626,N_455,N_363);
nand U627 (N_627,N_489,N_215);
and U628 (N_628,N_42,N_307);
or U629 (N_629,N_543,N_550);
nor U630 (N_630,N_518,N_492);
and U631 (N_631,N_246,N_323);
and U632 (N_632,N_82,N_234);
or U633 (N_633,N_64,N_22);
and U634 (N_634,N_218,N_481);
or U635 (N_635,N_231,N_458);
nand U636 (N_636,N_30,N_561);
nor U637 (N_637,N_206,N_37);
nand U638 (N_638,N_28,N_385);
xnor U639 (N_639,N_457,N_222);
nor U640 (N_640,N_381,N_228);
nor U641 (N_641,N_498,N_125);
and U642 (N_642,N_448,N_435);
nand U643 (N_643,N_520,N_547);
nand U644 (N_644,N_414,N_252);
or U645 (N_645,N_389,N_97);
nor U646 (N_646,N_198,N_456);
and U647 (N_647,N_161,N_432);
nor U648 (N_648,N_210,N_321);
and U649 (N_649,N_529,N_255);
or U650 (N_650,N_75,N_418);
nor U651 (N_651,N_560,N_453);
or U652 (N_652,N_83,N_515);
and U653 (N_653,N_434,N_141);
nand U654 (N_654,N_355,N_102);
nor U655 (N_655,N_144,N_233);
nand U656 (N_656,N_584,N_430);
and U657 (N_657,N_372,N_528);
and U658 (N_658,N_377,N_205);
or U659 (N_659,N_316,N_582);
nor U660 (N_660,N_326,N_585);
or U661 (N_661,N_554,N_291);
and U662 (N_662,N_366,N_195);
nand U663 (N_663,N_512,N_45);
and U664 (N_664,N_6,N_567);
or U665 (N_665,N_589,N_176);
and U666 (N_666,N_501,N_516);
and U667 (N_667,N_467,N_71);
nor U668 (N_668,N_220,N_136);
nand U669 (N_669,N_118,N_374);
nand U670 (N_670,N_380,N_350);
nand U671 (N_671,N_343,N_287);
nand U672 (N_672,N_440,N_296);
and U673 (N_673,N_211,N_40);
and U674 (N_674,N_491,N_157);
and U675 (N_675,N_495,N_148);
nand U676 (N_676,N_5,N_460);
and U677 (N_677,N_61,N_46);
and U678 (N_678,N_194,N_362);
and U679 (N_679,N_478,N_579);
nor U680 (N_680,N_14,N_238);
nand U681 (N_681,N_245,N_54);
or U682 (N_682,N_269,N_201);
and U683 (N_683,N_570,N_549);
nand U684 (N_684,N_535,N_517);
and U685 (N_685,N_558,N_309);
and U686 (N_686,N_341,N_573);
nand U687 (N_687,N_425,N_576);
and U688 (N_688,N_168,N_587);
nor U689 (N_689,N_532,N_361);
or U690 (N_690,N_171,N_70);
nor U691 (N_691,N_123,N_57);
and U692 (N_692,N_143,N_236);
or U693 (N_693,N_514,N_207);
or U694 (N_694,N_300,N_265);
xor U695 (N_695,N_486,N_13);
nor U696 (N_696,N_281,N_66);
or U697 (N_697,N_50,N_165);
or U698 (N_698,N_271,N_276);
or U699 (N_699,N_342,N_334);
and U700 (N_700,N_451,N_408);
nor U701 (N_701,N_329,N_203);
or U702 (N_702,N_74,N_449);
nor U703 (N_703,N_557,N_384);
nand U704 (N_704,N_559,N_120);
nor U705 (N_705,N_181,N_500);
nand U706 (N_706,N_131,N_47);
or U707 (N_707,N_376,N_349);
or U708 (N_708,N_229,N_436);
nor U709 (N_709,N_63,N_117);
nand U710 (N_710,N_298,N_67);
nor U711 (N_711,N_439,N_590);
or U712 (N_712,N_487,N_292);
nor U713 (N_713,N_392,N_403);
nor U714 (N_714,N_310,N_56);
nand U715 (N_715,N_415,N_428);
or U716 (N_716,N_581,N_427);
nand U717 (N_717,N_393,N_209);
nor U718 (N_718,N_358,N_68);
nor U719 (N_719,N_365,N_484);
and U720 (N_720,N_16,N_119);
nand U721 (N_721,N_60,N_24);
nand U722 (N_722,N_167,N_593);
or U723 (N_723,N_146,N_262);
nor U724 (N_724,N_177,N_196);
or U725 (N_725,N_158,N_179);
or U726 (N_726,N_476,N_367);
or U727 (N_727,N_189,N_396);
nand U728 (N_728,N_422,N_340);
and U729 (N_729,N_32,N_475);
and U730 (N_730,N_525,N_410);
nand U731 (N_731,N_147,N_306);
nor U732 (N_732,N_35,N_356);
nor U733 (N_733,N_139,N_186);
or U734 (N_734,N_536,N_270);
and U735 (N_735,N_17,N_313);
xnor U736 (N_736,N_438,N_224);
nand U737 (N_737,N_364,N_43);
nand U738 (N_738,N_320,N_540);
or U739 (N_739,N_330,N_299);
nand U740 (N_740,N_521,N_184);
or U741 (N_741,N_333,N_134);
and U742 (N_742,N_477,N_409);
and U743 (N_743,N_221,N_553);
nor U744 (N_744,N_391,N_447);
nor U745 (N_745,N_130,N_15);
or U746 (N_746,N_401,N_479);
nor U747 (N_747,N_85,N_556);
and U748 (N_748,N_424,N_96);
nand U749 (N_749,N_473,N_339);
or U750 (N_750,N_124,N_95);
or U751 (N_751,N_347,N_103);
nand U752 (N_752,N_423,N_73);
nor U753 (N_753,N_523,N_368);
nor U754 (N_754,N_472,N_336);
nor U755 (N_755,N_213,N_122);
or U756 (N_756,N_507,N_263);
and U757 (N_757,N_133,N_185);
or U758 (N_758,N_105,N_44);
nor U759 (N_759,N_417,N_565);
or U760 (N_760,N_129,N_174);
or U761 (N_761,N_311,N_578);
nor U762 (N_762,N_397,N_524);
or U763 (N_763,N_140,N_383);
or U764 (N_764,N_496,N_2);
nand U765 (N_765,N_155,N_388);
nand U766 (N_766,N_12,N_216);
or U767 (N_767,N_493,N_1);
and U768 (N_768,N_36,N_183);
and U769 (N_769,N_480,N_294);
nor U770 (N_770,N_577,N_327);
and U771 (N_771,N_328,N_509);
and U772 (N_772,N_284,N_508);
nor U773 (N_773,N_324,N_7);
nand U774 (N_774,N_178,N_226);
nor U775 (N_775,N_375,N_232);
and U776 (N_776,N_308,N_266);
nor U777 (N_777,N_597,N_27);
nor U778 (N_778,N_588,N_527);
and U779 (N_779,N_9,N_152);
xor U780 (N_780,N_314,N_562);
nor U781 (N_781,N_370,N_8);
or U782 (N_782,N_240,N_33);
nor U783 (N_783,N_369,N_208);
nor U784 (N_784,N_379,N_575);
or U785 (N_785,N_128,N_441);
and U786 (N_786,N_499,N_170);
nor U787 (N_787,N_78,N_373);
or U788 (N_788,N_285,N_537);
nor U789 (N_789,N_574,N_318);
or U790 (N_790,N_182,N_503);
nor U791 (N_791,N_533,N_506);
and U792 (N_792,N_249,N_337);
or U793 (N_793,N_568,N_325);
nand U794 (N_794,N_443,N_94);
and U795 (N_795,N_386,N_160);
and U796 (N_796,N_445,N_88);
nand U797 (N_797,N_112,N_461);
nand U798 (N_798,N_19,N_235);
and U799 (N_799,N_180,N_126);
nor U800 (N_800,N_172,N_345);
and U801 (N_801,N_154,N_264);
or U802 (N_802,N_286,N_538);
or U803 (N_803,N_400,N_59);
or U804 (N_804,N_421,N_53);
nand U805 (N_805,N_257,N_250);
and U806 (N_806,N_190,N_437);
nand U807 (N_807,N_348,N_452);
or U808 (N_808,N_544,N_38);
or U809 (N_809,N_251,N_92);
nand U810 (N_810,N_199,N_219);
and U811 (N_811,N_429,N_359);
or U812 (N_812,N_223,N_511);
or U813 (N_813,N_48,N_91);
nand U814 (N_814,N_89,N_471);
nor U815 (N_815,N_145,N_101);
nor U816 (N_816,N_301,N_539);
nor U817 (N_817,N_107,N_18);
nor U818 (N_818,N_302,N_485);
and U819 (N_819,N_295,N_566);
nor U820 (N_820,N_86,N_450);
nor U821 (N_821,N_106,N_413);
or U822 (N_822,N_488,N_29);
nand U823 (N_823,N_187,N_156);
nor U824 (N_824,N_244,N_100);
and U825 (N_825,N_49,N_382);
and U826 (N_826,N_371,N_297);
nand U827 (N_827,N_108,N_191);
nand U828 (N_828,N_132,N_354);
nand U829 (N_829,N_583,N_3);
nand U830 (N_830,N_331,N_21);
nand U831 (N_831,N_387,N_204);
and U832 (N_832,N_351,N_142);
nand U833 (N_833,N_474,N_278);
xor U834 (N_834,N_483,N_197);
nor U835 (N_835,N_510,N_531);
and U836 (N_836,N_571,N_166);
nor U837 (N_837,N_20,N_545);
nand U838 (N_838,N_431,N_111);
xnor U839 (N_839,N_282,N_482);
or U840 (N_840,N_230,N_594);
nand U841 (N_841,N_260,N_406);
or U842 (N_842,N_164,N_344);
and U843 (N_843,N_247,N_360);
nand U844 (N_844,N_193,N_137);
xor U845 (N_845,N_555,N_153);
nor U846 (N_846,N_11,N_288);
nand U847 (N_847,N_513,N_39);
nor U848 (N_848,N_34,N_51);
xor U849 (N_849,N_569,N_596);
nor U850 (N_850,N_357,N_212);
and U851 (N_851,N_237,N_99);
and U852 (N_852,N_534,N_81);
and U853 (N_853,N_227,N_116);
and U854 (N_854,N_315,N_420);
and U855 (N_855,N_274,N_551);
and U856 (N_856,N_522,N_62);
and U857 (N_857,N_159,N_395);
or U858 (N_858,N_113,N_390);
or U859 (N_859,N_469,N_31);
nand U860 (N_860,N_466,N_552);
or U861 (N_861,N_548,N_243);
nand U862 (N_862,N_275,N_317);
nand U863 (N_863,N_79,N_305);
and U864 (N_864,N_290,N_454);
or U865 (N_865,N_598,N_242);
or U866 (N_866,N_115,N_65);
nand U867 (N_867,N_572,N_93);
and U868 (N_868,N_505,N_378);
or U869 (N_869,N_402,N_225);
and U870 (N_870,N_0,N_322);
and U871 (N_871,N_405,N_149);
or U872 (N_872,N_312,N_239);
nand U873 (N_873,N_293,N_127);
nor U874 (N_874,N_121,N_41);
and U875 (N_875,N_268,N_258);
and U876 (N_876,N_98,N_433);
nor U877 (N_877,N_419,N_55);
or U878 (N_878,N_163,N_76);
nand U879 (N_879,N_504,N_200);
or U880 (N_880,N_416,N_497);
nor U881 (N_881,N_519,N_319);
nor U882 (N_882,N_109,N_541);
nor U883 (N_883,N_465,N_352);
and U884 (N_884,N_138,N_25);
and U885 (N_885,N_273,N_338);
and U886 (N_886,N_470,N_335);
or U887 (N_887,N_69,N_169);
nor U888 (N_888,N_150,N_23);
nor U889 (N_889,N_586,N_580);
nand U890 (N_890,N_592,N_254);
nor U891 (N_891,N_214,N_241);
nand U892 (N_892,N_459,N_407);
or U893 (N_893,N_442,N_412);
nor U894 (N_894,N_188,N_444);
nand U895 (N_895,N_4,N_463);
or U896 (N_896,N_468,N_114);
or U897 (N_897,N_599,N_173);
and U898 (N_898,N_591,N_175);
nor U899 (N_899,N_546,N_272);
and U900 (N_900,N_371,N_441);
or U901 (N_901,N_96,N_422);
nand U902 (N_902,N_590,N_560);
nor U903 (N_903,N_552,N_72);
and U904 (N_904,N_488,N_444);
and U905 (N_905,N_348,N_219);
nand U906 (N_906,N_361,N_204);
nor U907 (N_907,N_114,N_500);
nand U908 (N_908,N_118,N_547);
nor U909 (N_909,N_96,N_430);
nor U910 (N_910,N_312,N_160);
nand U911 (N_911,N_42,N_229);
nor U912 (N_912,N_459,N_23);
or U913 (N_913,N_578,N_552);
or U914 (N_914,N_381,N_417);
nor U915 (N_915,N_408,N_205);
nand U916 (N_916,N_135,N_19);
nand U917 (N_917,N_553,N_540);
nand U918 (N_918,N_79,N_56);
or U919 (N_919,N_466,N_64);
nor U920 (N_920,N_486,N_92);
or U921 (N_921,N_113,N_115);
and U922 (N_922,N_58,N_158);
or U923 (N_923,N_45,N_58);
and U924 (N_924,N_263,N_16);
nor U925 (N_925,N_168,N_402);
nand U926 (N_926,N_160,N_198);
or U927 (N_927,N_294,N_36);
nor U928 (N_928,N_56,N_87);
nor U929 (N_929,N_167,N_401);
or U930 (N_930,N_237,N_299);
nor U931 (N_931,N_291,N_493);
xor U932 (N_932,N_355,N_393);
and U933 (N_933,N_433,N_379);
nand U934 (N_934,N_405,N_35);
nor U935 (N_935,N_39,N_396);
nor U936 (N_936,N_174,N_34);
or U937 (N_937,N_473,N_90);
and U938 (N_938,N_240,N_331);
or U939 (N_939,N_519,N_594);
and U940 (N_940,N_185,N_324);
nand U941 (N_941,N_567,N_132);
and U942 (N_942,N_462,N_84);
or U943 (N_943,N_414,N_503);
nand U944 (N_944,N_480,N_260);
or U945 (N_945,N_459,N_525);
nor U946 (N_946,N_559,N_230);
nand U947 (N_947,N_536,N_164);
nor U948 (N_948,N_403,N_218);
nor U949 (N_949,N_124,N_178);
nor U950 (N_950,N_266,N_224);
nand U951 (N_951,N_570,N_89);
nand U952 (N_952,N_192,N_545);
nor U953 (N_953,N_23,N_446);
nand U954 (N_954,N_389,N_413);
nand U955 (N_955,N_71,N_394);
or U956 (N_956,N_583,N_138);
and U957 (N_957,N_122,N_509);
and U958 (N_958,N_427,N_194);
or U959 (N_959,N_416,N_77);
nand U960 (N_960,N_169,N_519);
nor U961 (N_961,N_212,N_139);
nand U962 (N_962,N_389,N_377);
nand U963 (N_963,N_228,N_276);
nand U964 (N_964,N_142,N_112);
nand U965 (N_965,N_382,N_581);
nor U966 (N_966,N_579,N_466);
or U967 (N_967,N_164,N_534);
nor U968 (N_968,N_402,N_182);
and U969 (N_969,N_331,N_414);
nor U970 (N_970,N_588,N_302);
nor U971 (N_971,N_267,N_469);
nand U972 (N_972,N_43,N_429);
nor U973 (N_973,N_544,N_105);
nor U974 (N_974,N_457,N_50);
nand U975 (N_975,N_394,N_302);
or U976 (N_976,N_34,N_263);
nand U977 (N_977,N_527,N_535);
and U978 (N_978,N_383,N_449);
nor U979 (N_979,N_163,N_560);
and U980 (N_980,N_469,N_161);
nor U981 (N_981,N_94,N_364);
nor U982 (N_982,N_588,N_406);
or U983 (N_983,N_221,N_411);
and U984 (N_984,N_99,N_408);
or U985 (N_985,N_209,N_409);
nor U986 (N_986,N_453,N_427);
nor U987 (N_987,N_361,N_495);
nand U988 (N_988,N_108,N_269);
nand U989 (N_989,N_357,N_340);
and U990 (N_990,N_585,N_455);
nor U991 (N_991,N_434,N_314);
and U992 (N_992,N_478,N_337);
and U993 (N_993,N_196,N_200);
nor U994 (N_994,N_575,N_506);
nand U995 (N_995,N_237,N_380);
or U996 (N_996,N_469,N_576);
and U997 (N_997,N_278,N_563);
or U998 (N_998,N_428,N_520);
nand U999 (N_999,N_365,N_31);
nor U1000 (N_1000,N_278,N_78);
nand U1001 (N_1001,N_550,N_373);
nand U1002 (N_1002,N_345,N_288);
nor U1003 (N_1003,N_539,N_499);
nand U1004 (N_1004,N_347,N_453);
nand U1005 (N_1005,N_361,N_166);
and U1006 (N_1006,N_579,N_197);
and U1007 (N_1007,N_117,N_332);
or U1008 (N_1008,N_305,N_191);
nand U1009 (N_1009,N_504,N_308);
nor U1010 (N_1010,N_312,N_130);
nor U1011 (N_1011,N_109,N_451);
nand U1012 (N_1012,N_6,N_374);
and U1013 (N_1013,N_560,N_227);
and U1014 (N_1014,N_331,N_517);
and U1015 (N_1015,N_589,N_92);
and U1016 (N_1016,N_59,N_197);
nand U1017 (N_1017,N_15,N_29);
nor U1018 (N_1018,N_395,N_108);
nand U1019 (N_1019,N_11,N_523);
and U1020 (N_1020,N_155,N_599);
or U1021 (N_1021,N_374,N_12);
nor U1022 (N_1022,N_428,N_99);
and U1023 (N_1023,N_454,N_247);
or U1024 (N_1024,N_366,N_38);
and U1025 (N_1025,N_123,N_135);
nor U1026 (N_1026,N_127,N_96);
and U1027 (N_1027,N_142,N_380);
and U1028 (N_1028,N_290,N_23);
nand U1029 (N_1029,N_590,N_200);
or U1030 (N_1030,N_234,N_415);
or U1031 (N_1031,N_474,N_551);
nor U1032 (N_1032,N_209,N_153);
or U1033 (N_1033,N_347,N_133);
nor U1034 (N_1034,N_65,N_222);
nand U1035 (N_1035,N_290,N_596);
nand U1036 (N_1036,N_237,N_252);
and U1037 (N_1037,N_373,N_342);
or U1038 (N_1038,N_377,N_118);
nor U1039 (N_1039,N_578,N_350);
nand U1040 (N_1040,N_184,N_96);
nand U1041 (N_1041,N_476,N_498);
or U1042 (N_1042,N_87,N_314);
nor U1043 (N_1043,N_116,N_514);
nor U1044 (N_1044,N_449,N_506);
and U1045 (N_1045,N_300,N_452);
nand U1046 (N_1046,N_350,N_493);
nand U1047 (N_1047,N_170,N_557);
and U1048 (N_1048,N_15,N_245);
nor U1049 (N_1049,N_189,N_151);
nand U1050 (N_1050,N_222,N_157);
nor U1051 (N_1051,N_227,N_13);
and U1052 (N_1052,N_267,N_62);
or U1053 (N_1053,N_313,N_336);
nor U1054 (N_1054,N_478,N_112);
nor U1055 (N_1055,N_495,N_164);
nand U1056 (N_1056,N_128,N_97);
nand U1057 (N_1057,N_401,N_598);
nand U1058 (N_1058,N_320,N_75);
nor U1059 (N_1059,N_466,N_480);
nand U1060 (N_1060,N_361,N_210);
nor U1061 (N_1061,N_203,N_590);
or U1062 (N_1062,N_268,N_77);
nor U1063 (N_1063,N_314,N_466);
nor U1064 (N_1064,N_474,N_105);
nand U1065 (N_1065,N_452,N_197);
and U1066 (N_1066,N_459,N_79);
nand U1067 (N_1067,N_365,N_106);
and U1068 (N_1068,N_362,N_452);
and U1069 (N_1069,N_40,N_375);
and U1070 (N_1070,N_12,N_575);
xor U1071 (N_1071,N_4,N_43);
and U1072 (N_1072,N_577,N_496);
or U1073 (N_1073,N_267,N_312);
and U1074 (N_1074,N_377,N_441);
or U1075 (N_1075,N_336,N_195);
nand U1076 (N_1076,N_18,N_336);
nor U1077 (N_1077,N_496,N_173);
nor U1078 (N_1078,N_347,N_191);
nand U1079 (N_1079,N_452,N_211);
nand U1080 (N_1080,N_528,N_159);
nand U1081 (N_1081,N_173,N_149);
and U1082 (N_1082,N_16,N_150);
nand U1083 (N_1083,N_588,N_332);
nor U1084 (N_1084,N_39,N_177);
nor U1085 (N_1085,N_433,N_187);
nand U1086 (N_1086,N_109,N_403);
nand U1087 (N_1087,N_438,N_314);
or U1088 (N_1088,N_474,N_125);
or U1089 (N_1089,N_455,N_354);
nand U1090 (N_1090,N_542,N_306);
nand U1091 (N_1091,N_448,N_499);
nand U1092 (N_1092,N_580,N_275);
and U1093 (N_1093,N_532,N_220);
or U1094 (N_1094,N_478,N_157);
and U1095 (N_1095,N_209,N_496);
nor U1096 (N_1096,N_34,N_410);
and U1097 (N_1097,N_337,N_96);
or U1098 (N_1098,N_37,N_264);
nand U1099 (N_1099,N_22,N_163);
nor U1100 (N_1100,N_337,N_508);
and U1101 (N_1101,N_200,N_46);
nor U1102 (N_1102,N_554,N_240);
nand U1103 (N_1103,N_315,N_88);
nand U1104 (N_1104,N_461,N_491);
or U1105 (N_1105,N_82,N_161);
and U1106 (N_1106,N_540,N_161);
and U1107 (N_1107,N_399,N_463);
or U1108 (N_1108,N_129,N_265);
and U1109 (N_1109,N_541,N_241);
nor U1110 (N_1110,N_266,N_195);
or U1111 (N_1111,N_79,N_113);
nor U1112 (N_1112,N_297,N_51);
nor U1113 (N_1113,N_41,N_31);
nand U1114 (N_1114,N_558,N_81);
nand U1115 (N_1115,N_598,N_297);
and U1116 (N_1116,N_456,N_68);
or U1117 (N_1117,N_578,N_438);
nand U1118 (N_1118,N_534,N_6);
nor U1119 (N_1119,N_236,N_138);
nand U1120 (N_1120,N_390,N_161);
nand U1121 (N_1121,N_127,N_590);
xor U1122 (N_1122,N_585,N_444);
nand U1123 (N_1123,N_156,N_384);
or U1124 (N_1124,N_260,N_279);
nand U1125 (N_1125,N_69,N_317);
nand U1126 (N_1126,N_348,N_120);
nor U1127 (N_1127,N_111,N_95);
nand U1128 (N_1128,N_13,N_586);
nor U1129 (N_1129,N_70,N_262);
and U1130 (N_1130,N_398,N_172);
or U1131 (N_1131,N_101,N_413);
and U1132 (N_1132,N_147,N_296);
and U1133 (N_1133,N_156,N_426);
nor U1134 (N_1134,N_235,N_256);
and U1135 (N_1135,N_522,N_537);
and U1136 (N_1136,N_558,N_412);
nor U1137 (N_1137,N_19,N_151);
and U1138 (N_1138,N_349,N_377);
nand U1139 (N_1139,N_348,N_195);
and U1140 (N_1140,N_404,N_148);
nand U1141 (N_1141,N_375,N_345);
nand U1142 (N_1142,N_471,N_168);
nor U1143 (N_1143,N_566,N_21);
or U1144 (N_1144,N_588,N_228);
nand U1145 (N_1145,N_312,N_425);
nor U1146 (N_1146,N_582,N_531);
nand U1147 (N_1147,N_159,N_38);
nand U1148 (N_1148,N_63,N_486);
or U1149 (N_1149,N_220,N_364);
nor U1150 (N_1150,N_364,N_202);
nand U1151 (N_1151,N_365,N_268);
or U1152 (N_1152,N_78,N_505);
nor U1153 (N_1153,N_185,N_146);
or U1154 (N_1154,N_563,N_195);
nor U1155 (N_1155,N_409,N_421);
nor U1156 (N_1156,N_574,N_8);
or U1157 (N_1157,N_62,N_295);
nand U1158 (N_1158,N_176,N_435);
nor U1159 (N_1159,N_4,N_184);
nand U1160 (N_1160,N_324,N_444);
nor U1161 (N_1161,N_273,N_94);
nor U1162 (N_1162,N_68,N_170);
nand U1163 (N_1163,N_468,N_405);
xnor U1164 (N_1164,N_359,N_524);
nor U1165 (N_1165,N_427,N_17);
nand U1166 (N_1166,N_571,N_392);
nand U1167 (N_1167,N_81,N_580);
or U1168 (N_1168,N_488,N_580);
nand U1169 (N_1169,N_396,N_252);
and U1170 (N_1170,N_582,N_377);
or U1171 (N_1171,N_93,N_243);
nand U1172 (N_1172,N_196,N_204);
and U1173 (N_1173,N_360,N_388);
and U1174 (N_1174,N_46,N_515);
or U1175 (N_1175,N_516,N_562);
or U1176 (N_1176,N_145,N_399);
nand U1177 (N_1177,N_441,N_82);
and U1178 (N_1178,N_334,N_595);
or U1179 (N_1179,N_517,N_582);
or U1180 (N_1180,N_517,N_148);
nor U1181 (N_1181,N_263,N_95);
nor U1182 (N_1182,N_240,N_97);
and U1183 (N_1183,N_292,N_154);
or U1184 (N_1184,N_253,N_349);
and U1185 (N_1185,N_75,N_347);
nand U1186 (N_1186,N_403,N_590);
nor U1187 (N_1187,N_569,N_450);
nand U1188 (N_1188,N_107,N_423);
or U1189 (N_1189,N_548,N_446);
and U1190 (N_1190,N_345,N_155);
xor U1191 (N_1191,N_130,N_570);
or U1192 (N_1192,N_313,N_409);
or U1193 (N_1193,N_80,N_504);
or U1194 (N_1194,N_276,N_328);
nor U1195 (N_1195,N_320,N_502);
and U1196 (N_1196,N_502,N_4);
nor U1197 (N_1197,N_401,N_121);
nor U1198 (N_1198,N_444,N_556);
nand U1199 (N_1199,N_58,N_430);
nand U1200 (N_1200,N_875,N_1016);
and U1201 (N_1201,N_828,N_1110);
nand U1202 (N_1202,N_720,N_985);
nor U1203 (N_1203,N_1081,N_682);
nand U1204 (N_1204,N_1126,N_939);
nor U1205 (N_1205,N_1164,N_908);
nor U1206 (N_1206,N_987,N_1027);
or U1207 (N_1207,N_696,N_704);
nor U1208 (N_1208,N_920,N_1043);
or U1209 (N_1209,N_817,N_1074);
or U1210 (N_1210,N_813,N_856);
xor U1211 (N_1211,N_902,N_650);
or U1212 (N_1212,N_623,N_659);
nand U1213 (N_1213,N_724,N_969);
and U1214 (N_1214,N_938,N_1096);
and U1215 (N_1215,N_1083,N_1188);
and U1216 (N_1216,N_714,N_1029);
and U1217 (N_1217,N_1009,N_1093);
or U1218 (N_1218,N_654,N_864);
nor U1219 (N_1219,N_721,N_1069);
or U1220 (N_1220,N_1003,N_841);
or U1221 (N_1221,N_753,N_824);
nor U1222 (N_1222,N_889,N_1176);
or U1223 (N_1223,N_797,N_1089);
nand U1224 (N_1224,N_1025,N_625);
and U1225 (N_1225,N_1041,N_1028);
nor U1226 (N_1226,N_899,N_612);
or U1227 (N_1227,N_983,N_781);
nor U1228 (N_1228,N_733,N_626);
or U1229 (N_1229,N_765,N_709);
or U1230 (N_1230,N_883,N_1147);
nand U1231 (N_1231,N_1080,N_636);
nor U1232 (N_1232,N_1156,N_1199);
nand U1233 (N_1233,N_727,N_853);
nand U1234 (N_1234,N_638,N_862);
nor U1235 (N_1235,N_995,N_1082);
nand U1236 (N_1236,N_627,N_992);
and U1237 (N_1237,N_955,N_988);
nor U1238 (N_1238,N_904,N_768);
nand U1239 (N_1239,N_1157,N_1075);
or U1240 (N_1240,N_1113,N_695);
or U1241 (N_1241,N_924,N_646);
and U1242 (N_1242,N_1150,N_741);
and U1243 (N_1243,N_1123,N_644);
nand U1244 (N_1244,N_1024,N_993);
and U1245 (N_1245,N_1065,N_870);
or U1246 (N_1246,N_1149,N_900);
or U1247 (N_1247,N_1192,N_831);
or U1248 (N_1248,N_1159,N_830);
nor U1249 (N_1249,N_705,N_1165);
and U1250 (N_1250,N_686,N_848);
nor U1251 (N_1251,N_749,N_867);
nor U1252 (N_1252,N_1131,N_736);
or U1253 (N_1253,N_1022,N_1152);
nand U1254 (N_1254,N_731,N_799);
nor U1255 (N_1255,N_1148,N_1106);
and U1256 (N_1256,N_754,N_671);
or U1257 (N_1257,N_1034,N_1181);
nor U1258 (N_1258,N_1114,N_897);
nand U1259 (N_1259,N_877,N_1142);
nor U1260 (N_1260,N_732,N_961);
nand U1261 (N_1261,N_673,N_688);
and U1262 (N_1262,N_681,N_666);
or U1263 (N_1263,N_930,N_1153);
nor U1264 (N_1264,N_871,N_665);
nand U1265 (N_1265,N_1044,N_725);
or U1266 (N_1266,N_986,N_868);
or U1267 (N_1267,N_611,N_726);
or U1268 (N_1268,N_1120,N_1112);
nand U1269 (N_1269,N_1039,N_743);
or U1270 (N_1270,N_818,N_850);
or U1271 (N_1271,N_1088,N_963);
and U1272 (N_1272,N_887,N_808);
or U1273 (N_1273,N_834,N_640);
and U1274 (N_1274,N_910,N_635);
nand U1275 (N_1275,N_1072,N_953);
nor U1276 (N_1276,N_1122,N_1099);
nand U1277 (N_1277,N_723,N_1138);
or U1278 (N_1278,N_748,N_1076);
nand U1279 (N_1279,N_1042,N_1079);
nand U1280 (N_1280,N_888,N_835);
nand U1281 (N_1281,N_735,N_717);
nand U1282 (N_1282,N_691,N_1007);
and U1283 (N_1283,N_1001,N_1014);
nor U1284 (N_1284,N_702,N_829);
nand U1285 (N_1285,N_1021,N_861);
nor U1286 (N_1286,N_970,N_1071);
nor U1287 (N_1287,N_648,N_913);
or U1288 (N_1288,N_1167,N_839);
nand U1289 (N_1289,N_901,N_943);
nor U1290 (N_1290,N_1118,N_798);
and U1291 (N_1291,N_892,N_1018);
nand U1292 (N_1292,N_621,N_619);
and U1293 (N_1293,N_1166,N_645);
nor U1294 (N_1294,N_872,N_1063);
or U1295 (N_1295,N_785,N_613);
xnor U1296 (N_1296,N_1066,N_707);
and U1297 (N_1297,N_787,N_819);
nand U1298 (N_1298,N_1023,N_926);
or U1299 (N_1299,N_775,N_1011);
nor U1300 (N_1300,N_715,N_1100);
nor U1301 (N_1301,N_1013,N_911);
or U1302 (N_1302,N_1070,N_620);
and U1303 (N_1303,N_974,N_639);
nand U1304 (N_1304,N_1160,N_914);
nand U1305 (N_1305,N_1109,N_1179);
and U1306 (N_1306,N_773,N_1172);
and U1307 (N_1307,N_1017,N_791);
and U1308 (N_1308,N_701,N_942);
or U1309 (N_1309,N_784,N_652);
or U1310 (N_1310,N_771,N_616);
nand U1311 (N_1311,N_958,N_710);
or U1312 (N_1312,N_617,N_832);
or U1313 (N_1313,N_764,N_869);
nor U1314 (N_1314,N_1101,N_1154);
or U1315 (N_1315,N_1115,N_601);
or U1316 (N_1316,N_972,N_1078);
nand U1317 (N_1317,N_615,N_886);
or U1318 (N_1318,N_751,N_1091);
and U1319 (N_1319,N_814,N_789);
nor U1320 (N_1320,N_905,N_1056);
nand U1321 (N_1321,N_1004,N_1174);
and U1322 (N_1322,N_921,N_1026);
and U1323 (N_1323,N_804,N_1186);
nand U1324 (N_1324,N_1162,N_821);
nand U1325 (N_1325,N_761,N_1092);
nand U1326 (N_1326,N_922,N_1040);
and U1327 (N_1327,N_622,N_999);
or U1328 (N_1328,N_989,N_647);
or U1329 (N_1329,N_1141,N_1094);
and U1330 (N_1330,N_783,N_600);
and U1331 (N_1331,N_738,N_1006);
or U1332 (N_1332,N_941,N_952);
nor U1333 (N_1333,N_827,N_602);
nand U1334 (N_1334,N_1008,N_1111);
nor U1335 (N_1335,N_757,N_854);
and U1336 (N_1336,N_894,N_1020);
nor U1337 (N_1337,N_766,N_697);
or U1338 (N_1338,N_909,N_1032);
or U1339 (N_1339,N_959,N_676);
and U1340 (N_1340,N_729,N_801);
nor U1341 (N_1341,N_1133,N_708);
nor U1342 (N_1342,N_712,N_843);
or U1343 (N_1343,N_758,N_1151);
nor U1344 (N_1344,N_632,N_1053);
or U1345 (N_1345,N_672,N_846);
or U1346 (N_1346,N_965,N_763);
nor U1347 (N_1347,N_893,N_1128);
and U1348 (N_1348,N_994,N_896);
and U1349 (N_1349,N_1119,N_1098);
nand U1350 (N_1350,N_982,N_1005);
nor U1351 (N_1351,N_700,N_865);
or U1352 (N_1352,N_614,N_770);
or U1353 (N_1353,N_945,N_1035);
nand U1354 (N_1354,N_1054,N_1077);
nand U1355 (N_1355,N_1135,N_1140);
and U1356 (N_1356,N_742,N_1068);
and U1357 (N_1357,N_649,N_778);
nand U1358 (N_1358,N_825,N_933);
nor U1359 (N_1359,N_928,N_1171);
and U1360 (N_1360,N_651,N_1173);
nor U1361 (N_1361,N_971,N_807);
nand U1362 (N_1362,N_1124,N_793);
or U1363 (N_1363,N_669,N_876);
nor U1364 (N_1364,N_1051,N_1050);
nor U1365 (N_1365,N_934,N_826);
or U1366 (N_1366,N_603,N_802);
or U1367 (N_1367,N_1169,N_859);
nand U1368 (N_1368,N_806,N_1177);
nor U1369 (N_1369,N_948,N_956);
and U1370 (N_1370,N_842,N_1030);
nand U1371 (N_1371,N_805,N_932);
nand U1372 (N_1372,N_1183,N_847);
nor U1373 (N_1373,N_1125,N_745);
nor U1374 (N_1374,N_604,N_929);
nand U1375 (N_1375,N_1175,N_852);
and U1376 (N_1376,N_838,N_884);
nor U1377 (N_1377,N_923,N_1158);
nand U1378 (N_1378,N_874,N_873);
nand U1379 (N_1379,N_949,N_734);
or U1380 (N_1380,N_816,N_947);
nand U1381 (N_1381,N_678,N_1198);
nor U1382 (N_1382,N_858,N_1073);
or U1383 (N_1383,N_1161,N_1060);
nand U1384 (N_1384,N_674,N_752);
nand U1385 (N_1385,N_1190,N_634);
or U1386 (N_1386,N_1178,N_1121);
and U1387 (N_1387,N_1102,N_1058);
nor U1388 (N_1388,N_1031,N_1194);
and U1389 (N_1389,N_1045,N_1136);
or U1390 (N_1390,N_1000,N_1116);
or U1391 (N_1391,N_1134,N_1097);
nand U1392 (N_1392,N_1055,N_719);
and U1393 (N_1393,N_1002,N_1057);
or U1394 (N_1394,N_1197,N_975);
and U1395 (N_1395,N_1037,N_747);
or U1396 (N_1396,N_629,N_642);
and U1397 (N_1397,N_1104,N_1095);
and U1398 (N_1398,N_912,N_916);
nor U1399 (N_1399,N_1143,N_739);
nand U1400 (N_1400,N_1015,N_879);
nor U1401 (N_1401,N_815,N_1196);
or U1402 (N_1402,N_1146,N_722);
or U1403 (N_1403,N_657,N_984);
and U1404 (N_1404,N_962,N_946);
or U1405 (N_1405,N_1191,N_906);
and U1406 (N_1406,N_667,N_1087);
or U1407 (N_1407,N_796,N_692);
and U1408 (N_1408,N_931,N_810);
and U1409 (N_1409,N_607,N_919);
nand U1410 (N_1410,N_936,N_756);
nor U1411 (N_1411,N_610,N_1117);
nor U1412 (N_1412,N_680,N_795);
or U1413 (N_1413,N_631,N_1052);
nand U1414 (N_1414,N_849,N_837);
nand U1415 (N_1415,N_890,N_836);
or U1416 (N_1416,N_718,N_746);
nand U1417 (N_1417,N_755,N_658);
or U1418 (N_1418,N_954,N_1127);
and U1419 (N_1419,N_917,N_991);
or U1420 (N_1420,N_728,N_1130);
or U1421 (N_1421,N_762,N_786);
nor U1422 (N_1422,N_779,N_737);
nand U1423 (N_1423,N_630,N_689);
nor U1424 (N_1424,N_608,N_968);
xor U1425 (N_1425,N_1062,N_918);
or U1426 (N_1426,N_744,N_643);
and U1427 (N_1427,N_973,N_690);
nor U1428 (N_1428,N_1036,N_809);
nor U1429 (N_1429,N_845,N_792);
nand U1430 (N_1430,N_951,N_857);
nor U1431 (N_1431,N_698,N_606);
nand U1432 (N_1432,N_656,N_776);
nor U1433 (N_1433,N_1168,N_1046);
nor U1434 (N_1434,N_618,N_664);
nor U1435 (N_1435,N_1137,N_800);
and U1436 (N_1436,N_1038,N_1103);
or U1437 (N_1437,N_977,N_1019);
nand U1438 (N_1438,N_895,N_1064);
or U1439 (N_1439,N_609,N_1107);
nand U1440 (N_1440,N_1108,N_767);
nand U1441 (N_1441,N_885,N_937);
nor U1442 (N_1442,N_851,N_782);
nor U1443 (N_1443,N_1180,N_706);
nand U1444 (N_1444,N_660,N_1195);
nand U1445 (N_1445,N_1047,N_1048);
or U1446 (N_1446,N_624,N_679);
or U1447 (N_1447,N_967,N_730);
nand U1448 (N_1448,N_935,N_605);
nand U1449 (N_1449,N_957,N_1049);
and U1450 (N_1450,N_1033,N_1185);
nor U1451 (N_1451,N_711,N_978);
nand U1452 (N_1452,N_1129,N_655);
nand U1453 (N_1453,N_683,N_1132);
or U1454 (N_1454,N_907,N_663);
nor U1455 (N_1455,N_1145,N_820);
and U1456 (N_1456,N_759,N_833);
or U1457 (N_1457,N_633,N_1184);
nor U1458 (N_1458,N_990,N_866);
nor U1459 (N_1459,N_860,N_966);
nor U1460 (N_1460,N_1189,N_1144);
or U1461 (N_1461,N_1086,N_637);
or U1462 (N_1462,N_794,N_878);
nor U1463 (N_1463,N_944,N_823);
and U1464 (N_1464,N_1139,N_662);
nor U1465 (N_1465,N_1193,N_1059);
and U1466 (N_1466,N_903,N_675);
and U1467 (N_1467,N_772,N_1010);
and U1468 (N_1468,N_811,N_880);
and U1469 (N_1469,N_1163,N_693);
nand U1470 (N_1470,N_694,N_780);
or U1471 (N_1471,N_1012,N_915);
and U1472 (N_1472,N_998,N_716);
and U1473 (N_1473,N_1105,N_891);
nor U1474 (N_1474,N_882,N_979);
or U1475 (N_1475,N_788,N_881);
nand U1476 (N_1476,N_844,N_777);
nor U1477 (N_1477,N_670,N_980);
or U1478 (N_1478,N_628,N_687);
nor U1479 (N_1479,N_898,N_964);
or U1480 (N_1480,N_760,N_981);
nor U1481 (N_1481,N_1084,N_927);
and U1482 (N_1482,N_997,N_653);
or U1483 (N_1483,N_822,N_1155);
nand U1484 (N_1484,N_790,N_1182);
nor U1485 (N_1485,N_699,N_1170);
and U1486 (N_1486,N_1061,N_668);
and U1487 (N_1487,N_641,N_1090);
and U1488 (N_1488,N_769,N_803);
and U1489 (N_1489,N_925,N_740);
or U1490 (N_1490,N_1187,N_996);
nand U1491 (N_1491,N_684,N_855);
or U1492 (N_1492,N_960,N_976);
nand U1493 (N_1493,N_703,N_950);
and U1494 (N_1494,N_774,N_940);
nand U1495 (N_1495,N_750,N_863);
or U1496 (N_1496,N_812,N_713);
nand U1497 (N_1497,N_661,N_677);
or U1498 (N_1498,N_1067,N_840);
or U1499 (N_1499,N_1085,N_685);
or U1500 (N_1500,N_947,N_925);
or U1501 (N_1501,N_607,N_902);
or U1502 (N_1502,N_1006,N_915);
and U1503 (N_1503,N_779,N_849);
and U1504 (N_1504,N_1141,N_746);
or U1505 (N_1505,N_624,N_1008);
nand U1506 (N_1506,N_614,N_725);
or U1507 (N_1507,N_759,N_841);
nand U1508 (N_1508,N_1113,N_620);
or U1509 (N_1509,N_896,N_695);
and U1510 (N_1510,N_728,N_754);
or U1511 (N_1511,N_1187,N_1125);
nor U1512 (N_1512,N_736,N_1164);
and U1513 (N_1513,N_606,N_763);
or U1514 (N_1514,N_1146,N_962);
nand U1515 (N_1515,N_860,N_1157);
or U1516 (N_1516,N_1115,N_742);
and U1517 (N_1517,N_966,N_1095);
nand U1518 (N_1518,N_944,N_1152);
or U1519 (N_1519,N_697,N_858);
or U1520 (N_1520,N_1192,N_809);
and U1521 (N_1521,N_633,N_1023);
nor U1522 (N_1522,N_1012,N_1035);
nand U1523 (N_1523,N_690,N_619);
and U1524 (N_1524,N_889,N_1040);
nor U1525 (N_1525,N_1167,N_691);
nor U1526 (N_1526,N_824,N_1106);
and U1527 (N_1527,N_954,N_838);
nor U1528 (N_1528,N_953,N_1097);
and U1529 (N_1529,N_781,N_938);
and U1530 (N_1530,N_803,N_721);
nand U1531 (N_1531,N_780,N_957);
nand U1532 (N_1532,N_842,N_905);
nor U1533 (N_1533,N_696,N_827);
or U1534 (N_1534,N_1043,N_678);
nand U1535 (N_1535,N_884,N_858);
nand U1536 (N_1536,N_1160,N_799);
nand U1537 (N_1537,N_832,N_1195);
or U1538 (N_1538,N_1162,N_980);
nand U1539 (N_1539,N_1014,N_735);
nor U1540 (N_1540,N_774,N_996);
xnor U1541 (N_1541,N_1156,N_999);
xor U1542 (N_1542,N_1168,N_1145);
nand U1543 (N_1543,N_1187,N_803);
nor U1544 (N_1544,N_1148,N_1072);
and U1545 (N_1545,N_840,N_1096);
and U1546 (N_1546,N_1078,N_948);
or U1547 (N_1547,N_961,N_1163);
and U1548 (N_1548,N_985,N_650);
and U1549 (N_1549,N_720,N_737);
nor U1550 (N_1550,N_600,N_1060);
and U1551 (N_1551,N_769,N_1099);
nor U1552 (N_1552,N_1022,N_751);
nor U1553 (N_1553,N_644,N_716);
nand U1554 (N_1554,N_716,N_704);
and U1555 (N_1555,N_895,N_613);
nand U1556 (N_1556,N_676,N_708);
nor U1557 (N_1557,N_1196,N_900);
nand U1558 (N_1558,N_632,N_1036);
or U1559 (N_1559,N_618,N_761);
nand U1560 (N_1560,N_886,N_1090);
nor U1561 (N_1561,N_641,N_1102);
nand U1562 (N_1562,N_1108,N_733);
nand U1563 (N_1563,N_1097,N_783);
nor U1564 (N_1564,N_610,N_1058);
nand U1565 (N_1565,N_1111,N_1044);
and U1566 (N_1566,N_808,N_965);
or U1567 (N_1567,N_805,N_846);
or U1568 (N_1568,N_754,N_717);
or U1569 (N_1569,N_778,N_639);
or U1570 (N_1570,N_919,N_708);
nand U1571 (N_1571,N_1018,N_965);
or U1572 (N_1572,N_820,N_975);
nand U1573 (N_1573,N_1158,N_610);
nand U1574 (N_1574,N_993,N_905);
or U1575 (N_1575,N_660,N_814);
or U1576 (N_1576,N_622,N_851);
nand U1577 (N_1577,N_707,N_651);
or U1578 (N_1578,N_1026,N_812);
nor U1579 (N_1579,N_655,N_755);
or U1580 (N_1580,N_1132,N_944);
or U1581 (N_1581,N_1057,N_1153);
and U1582 (N_1582,N_981,N_961);
and U1583 (N_1583,N_723,N_1068);
nor U1584 (N_1584,N_841,N_638);
or U1585 (N_1585,N_728,N_902);
or U1586 (N_1586,N_1177,N_957);
nand U1587 (N_1587,N_854,N_750);
nand U1588 (N_1588,N_826,N_1073);
or U1589 (N_1589,N_898,N_868);
and U1590 (N_1590,N_627,N_916);
nand U1591 (N_1591,N_1064,N_723);
nand U1592 (N_1592,N_780,N_756);
and U1593 (N_1593,N_1089,N_843);
and U1594 (N_1594,N_878,N_964);
nor U1595 (N_1595,N_978,N_1031);
and U1596 (N_1596,N_821,N_1010);
nand U1597 (N_1597,N_858,N_767);
or U1598 (N_1598,N_1073,N_692);
or U1599 (N_1599,N_636,N_689);
nor U1600 (N_1600,N_962,N_683);
nor U1601 (N_1601,N_1006,N_1136);
nand U1602 (N_1602,N_1196,N_953);
nand U1603 (N_1603,N_906,N_829);
and U1604 (N_1604,N_833,N_1074);
or U1605 (N_1605,N_613,N_1089);
nand U1606 (N_1606,N_684,N_643);
nand U1607 (N_1607,N_851,N_637);
or U1608 (N_1608,N_1130,N_1052);
nand U1609 (N_1609,N_984,N_656);
nand U1610 (N_1610,N_785,N_712);
nor U1611 (N_1611,N_985,N_605);
and U1612 (N_1612,N_1199,N_919);
or U1613 (N_1613,N_975,N_642);
nand U1614 (N_1614,N_698,N_930);
or U1615 (N_1615,N_1126,N_1187);
and U1616 (N_1616,N_845,N_825);
nand U1617 (N_1617,N_982,N_912);
or U1618 (N_1618,N_650,N_1090);
or U1619 (N_1619,N_794,N_1125);
nor U1620 (N_1620,N_823,N_810);
nand U1621 (N_1621,N_907,N_759);
or U1622 (N_1622,N_989,N_894);
and U1623 (N_1623,N_885,N_610);
nor U1624 (N_1624,N_773,N_1090);
nand U1625 (N_1625,N_967,N_893);
nor U1626 (N_1626,N_782,N_744);
or U1627 (N_1627,N_957,N_1196);
nor U1628 (N_1628,N_1131,N_1174);
and U1629 (N_1629,N_742,N_801);
nand U1630 (N_1630,N_628,N_825);
nor U1631 (N_1631,N_659,N_652);
nor U1632 (N_1632,N_1198,N_763);
or U1633 (N_1633,N_920,N_867);
nor U1634 (N_1634,N_793,N_1100);
nand U1635 (N_1635,N_600,N_1070);
nor U1636 (N_1636,N_1139,N_643);
and U1637 (N_1637,N_957,N_1118);
nand U1638 (N_1638,N_1052,N_1119);
nand U1639 (N_1639,N_915,N_680);
or U1640 (N_1640,N_786,N_829);
nand U1641 (N_1641,N_978,N_913);
or U1642 (N_1642,N_629,N_857);
nand U1643 (N_1643,N_780,N_1031);
nor U1644 (N_1644,N_857,N_1070);
or U1645 (N_1645,N_764,N_858);
and U1646 (N_1646,N_666,N_866);
nand U1647 (N_1647,N_600,N_644);
nand U1648 (N_1648,N_785,N_975);
nor U1649 (N_1649,N_818,N_809);
nor U1650 (N_1650,N_923,N_1142);
nor U1651 (N_1651,N_964,N_998);
nand U1652 (N_1652,N_1070,N_924);
and U1653 (N_1653,N_645,N_817);
nor U1654 (N_1654,N_1197,N_795);
and U1655 (N_1655,N_949,N_695);
or U1656 (N_1656,N_684,N_833);
nor U1657 (N_1657,N_932,N_734);
nand U1658 (N_1658,N_1041,N_888);
nand U1659 (N_1659,N_927,N_684);
nor U1660 (N_1660,N_1122,N_1136);
or U1661 (N_1661,N_1021,N_688);
nand U1662 (N_1662,N_1048,N_960);
and U1663 (N_1663,N_656,N_860);
or U1664 (N_1664,N_1035,N_620);
or U1665 (N_1665,N_989,N_765);
nor U1666 (N_1666,N_1042,N_853);
nor U1667 (N_1667,N_1174,N_1044);
nand U1668 (N_1668,N_692,N_984);
or U1669 (N_1669,N_1070,N_1089);
or U1670 (N_1670,N_716,N_887);
and U1671 (N_1671,N_1126,N_878);
and U1672 (N_1672,N_853,N_1075);
or U1673 (N_1673,N_1107,N_740);
or U1674 (N_1674,N_627,N_950);
or U1675 (N_1675,N_971,N_678);
or U1676 (N_1676,N_893,N_827);
or U1677 (N_1677,N_964,N_958);
or U1678 (N_1678,N_1083,N_1101);
or U1679 (N_1679,N_1064,N_1196);
or U1680 (N_1680,N_744,N_711);
nor U1681 (N_1681,N_1169,N_999);
nand U1682 (N_1682,N_755,N_743);
and U1683 (N_1683,N_917,N_680);
nand U1684 (N_1684,N_888,N_1132);
nand U1685 (N_1685,N_1060,N_1027);
nand U1686 (N_1686,N_743,N_624);
or U1687 (N_1687,N_620,N_614);
or U1688 (N_1688,N_733,N_676);
nor U1689 (N_1689,N_624,N_722);
and U1690 (N_1690,N_829,N_683);
and U1691 (N_1691,N_608,N_1099);
nor U1692 (N_1692,N_1192,N_956);
nand U1693 (N_1693,N_1132,N_1137);
nor U1694 (N_1694,N_1118,N_793);
or U1695 (N_1695,N_808,N_1150);
nor U1696 (N_1696,N_1072,N_850);
or U1697 (N_1697,N_925,N_1108);
or U1698 (N_1698,N_707,N_1168);
or U1699 (N_1699,N_653,N_1146);
nor U1700 (N_1700,N_879,N_891);
nor U1701 (N_1701,N_779,N_615);
nand U1702 (N_1702,N_801,N_863);
or U1703 (N_1703,N_632,N_625);
and U1704 (N_1704,N_932,N_1073);
nor U1705 (N_1705,N_718,N_698);
nor U1706 (N_1706,N_1169,N_800);
nor U1707 (N_1707,N_1096,N_1198);
or U1708 (N_1708,N_857,N_632);
and U1709 (N_1709,N_892,N_815);
or U1710 (N_1710,N_796,N_816);
xor U1711 (N_1711,N_1140,N_960);
or U1712 (N_1712,N_1040,N_907);
or U1713 (N_1713,N_780,N_930);
and U1714 (N_1714,N_835,N_837);
nand U1715 (N_1715,N_709,N_706);
or U1716 (N_1716,N_801,N_822);
nor U1717 (N_1717,N_1096,N_691);
and U1718 (N_1718,N_950,N_880);
nand U1719 (N_1719,N_1018,N_756);
nand U1720 (N_1720,N_783,N_1005);
nor U1721 (N_1721,N_669,N_882);
nand U1722 (N_1722,N_848,N_1001);
or U1723 (N_1723,N_991,N_783);
nand U1724 (N_1724,N_1026,N_1156);
nor U1725 (N_1725,N_956,N_774);
or U1726 (N_1726,N_1043,N_843);
or U1727 (N_1727,N_999,N_1035);
and U1728 (N_1728,N_1084,N_962);
or U1729 (N_1729,N_703,N_721);
nor U1730 (N_1730,N_625,N_839);
nand U1731 (N_1731,N_987,N_853);
nand U1732 (N_1732,N_949,N_609);
nor U1733 (N_1733,N_1078,N_1068);
nor U1734 (N_1734,N_819,N_852);
and U1735 (N_1735,N_1079,N_866);
and U1736 (N_1736,N_688,N_1011);
and U1737 (N_1737,N_1140,N_835);
nor U1738 (N_1738,N_1037,N_815);
xor U1739 (N_1739,N_603,N_1139);
and U1740 (N_1740,N_999,N_1002);
and U1741 (N_1741,N_1126,N_936);
nand U1742 (N_1742,N_938,N_1174);
nand U1743 (N_1743,N_1065,N_1177);
or U1744 (N_1744,N_1009,N_909);
nand U1745 (N_1745,N_1170,N_1192);
and U1746 (N_1746,N_607,N_670);
or U1747 (N_1747,N_779,N_1011);
and U1748 (N_1748,N_604,N_873);
or U1749 (N_1749,N_913,N_1151);
or U1750 (N_1750,N_789,N_1146);
nor U1751 (N_1751,N_1102,N_1178);
nand U1752 (N_1752,N_943,N_1034);
or U1753 (N_1753,N_943,N_1083);
or U1754 (N_1754,N_734,N_1001);
nand U1755 (N_1755,N_684,N_1034);
and U1756 (N_1756,N_1012,N_843);
nand U1757 (N_1757,N_886,N_990);
nand U1758 (N_1758,N_806,N_834);
or U1759 (N_1759,N_1186,N_1021);
nor U1760 (N_1760,N_947,N_997);
and U1761 (N_1761,N_1113,N_770);
xnor U1762 (N_1762,N_808,N_1148);
and U1763 (N_1763,N_818,N_616);
nand U1764 (N_1764,N_1001,N_600);
nor U1765 (N_1765,N_923,N_984);
or U1766 (N_1766,N_667,N_976);
nor U1767 (N_1767,N_668,N_1011);
nor U1768 (N_1768,N_1194,N_930);
and U1769 (N_1769,N_819,N_1127);
nand U1770 (N_1770,N_611,N_1014);
nand U1771 (N_1771,N_605,N_1058);
and U1772 (N_1772,N_1111,N_1197);
nor U1773 (N_1773,N_1156,N_1057);
or U1774 (N_1774,N_1121,N_736);
or U1775 (N_1775,N_842,N_639);
and U1776 (N_1776,N_612,N_944);
nand U1777 (N_1777,N_1052,N_673);
and U1778 (N_1778,N_877,N_807);
and U1779 (N_1779,N_764,N_1142);
nand U1780 (N_1780,N_1161,N_1000);
nor U1781 (N_1781,N_836,N_602);
nand U1782 (N_1782,N_933,N_613);
nand U1783 (N_1783,N_1127,N_619);
nor U1784 (N_1784,N_646,N_747);
nand U1785 (N_1785,N_786,N_904);
and U1786 (N_1786,N_876,N_786);
nor U1787 (N_1787,N_792,N_1053);
and U1788 (N_1788,N_874,N_1161);
and U1789 (N_1789,N_648,N_858);
and U1790 (N_1790,N_833,N_1035);
nand U1791 (N_1791,N_1108,N_823);
or U1792 (N_1792,N_1163,N_1115);
nor U1793 (N_1793,N_1158,N_854);
nand U1794 (N_1794,N_778,N_821);
nand U1795 (N_1795,N_783,N_1163);
or U1796 (N_1796,N_877,N_961);
nand U1797 (N_1797,N_1126,N_608);
nand U1798 (N_1798,N_1087,N_630);
and U1799 (N_1799,N_634,N_870);
or U1800 (N_1800,N_1208,N_1664);
and U1801 (N_1801,N_1259,N_1312);
nand U1802 (N_1802,N_1645,N_1723);
nor U1803 (N_1803,N_1622,N_1660);
nor U1804 (N_1804,N_1762,N_1548);
and U1805 (N_1805,N_1559,N_1528);
nand U1806 (N_1806,N_1397,N_1783);
nand U1807 (N_1807,N_1641,N_1751);
nand U1808 (N_1808,N_1368,N_1781);
nand U1809 (N_1809,N_1687,N_1296);
and U1810 (N_1810,N_1514,N_1434);
nand U1811 (N_1811,N_1663,N_1530);
nor U1812 (N_1812,N_1387,N_1728);
xnor U1813 (N_1813,N_1484,N_1444);
and U1814 (N_1814,N_1381,N_1202);
and U1815 (N_1815,N_1411,N_1347);
nor U1816 (N_1816,N_1759,N_1386);
or U1817 (N_1817,N_1705,N_1709);
and U1818 (N_1818,N_1704,N_1694);
and U1819 (N_1819,N_1509,N_1336);
nor U1820 (N_1820,N_1582,N_1589);
or U1821 (N_1821,N_1313,N_1266);
nand U1822 (N_1822,N_1287,N_1451);
nand U1823 (N_1823,N_1238,N_1719);
nor U1824 (N_1824,N_1334,N_1211);
or U1825 (N_1825,N_1649,N_1419);
and U1826 (N_1826,N_1575,N_1608);
nand U1827 (N_1827,N_1477,N_1407);
or U1828 (N_1828,N_1669,N_1489);
or U1829 (N_1829,N_1526,N_1349);
xnor U1830 (N_1830,N_1683,N_1460);
or U1831 (N_1831,N_1416,N_1706);
and U1832 (N_1832,N_1616,N_1634);
nor U1833 (N_1833,N_1466,N_1539);
nand U1834 (N_1834,N_1772,N_1670);
nand U1835 (N_1835,N_1724,N_1638);
and U1836 (N_1836,N_1281,N_1495);
nand U1837 (N_1837,N_1506,N_1674);
and U1838 (N_1838,N_1666,N_1456);
nor U1839 (N_1839,N_1417,N_1682);
or U1840 (N_1840,N_1439,N_1250);
and U1841 (N_1841,N_1760,N_1251);
or U1842 (N_1842,N_1301,N_1327);
and U1843 (N_1843,N_1345,N_1586);
or U1844 (N_1844,N_1615,N_1343);
and U1845 (N_1845,N_1453,N_1237);
nor U1846 (N_1846,N_1303,N_1512);
or U1847 (N_1847,N_1621,N_1295);
or U1848 (N_1848,N_1525,N_1227);
or U1849 (N_1849,N_1423,N_1502);
or U1850 (N_1850,N_1756,N_1225);
or U1851 (N_1851,N_1628,N_1277);
or U1852 (N_1852,N_1410,N_1798);
or U1853 (N_1853,N_1403,N_1642);
and U1854 (N_1854,N_1556,N_1306);
or U1855 (N_1855,N_1372,N_1401);
nand U1856 (N_1856,N_1521,N_1684);
nor U1857 (N_1857,N_1209,N_1631);
or U1858 (N_1858,N_1604,N_1662);
nor U1859 (N_1859,N_1445,N_1602);
nor U1860 (N_1860,N_1424,N_1440);
nand U1861 (N_1861,N_1206,N_1763);
nor U1862 (N_1862,N_1464,N_1665);
or U1863 (N_1863,N_1790,N_1226);
nand U1864 (N_1864,N_1718,N_1532);
and U1865 (N_1865,N_1203,N_1777);
nor U1866 (N_1866,N_1335,N_1243);
and U1867 (N_1867,N_1292,N_1776);
or U1868 (N_1868,N_1467,N_1293);
and U1869 (N_1869,N_1324,N_1560);
nor U1870 (N_1870,N_1613,N_1761);
nand U1871 (N_1871,N_1657,N_1519);
and U1872 (N_1872,N_1508,N_1536);
and U1873 (N_1873,N_1627,N_1275);
nand U1874 (N_1874,N_1764,N_1435);
nand U1875 (N_1875,N_1352,N_1216);
nor U1876 (N_1876,N_1429,N_1461);
nand U1877 (N_1877,N_1624,N_1780);
nor U1878 (N_1878,N_1448,N_1637);
and U1879 (N_1879,N_1591,N_1733);
and U1880 (N_1880,N_1233,N_1430);
nor U1881 (N_1881,N_1205,N_1747);
nand U1882 (N_1882,N_1558,N_1650);
nand U1883 (N_1883,N_1374,N_1223);
nand U1884 (N_1884,N_1779,N_1738);
nand U1885 (N_1885,N_1305,N_1737);
and U1886 (N_1886,N_1260,N_1778);
and U1887 (N_1887,N_1354,N_1362);
nand U1888 (N_1888,N_1715,N_1702);
nand U1889 (N_1889,N_1332,N_1241);
nand U1890 (N_1890,N_1302,N_1325);
or U1891 (N_1891,N_1446,N_1735);
and U1892 (N_1892,N_1271,N_1428);
or U1893 (N_1893,N_1252,N_1585);
and U1894 (N_1894,N_1623,N_1597);
nand U1895 (N_1895,N_1677,N_1462);
and U1896 (N_1896,N_1393,N_1283);
nor U1897 (N_1897,N_1341,N_1771);
nand U1898 (N_1898,N_1552,N_1520);
and U1899 (N_1899,N_1257,N_1413);
and U1900 (N_1900,N_1708,N_1543);
nor U1901 (N_1901,N_1745,N_1443);
nor U1902 (N_1902,N_1554,N_1563);
nand U1903 (N_1903,N_1425,N_1373);
nor U1904 (N_1904,N_1310,N_1245);
and U1905 (N_1905,N_1395,N_1505);
and U1906 (N_1906,N_1782,N_1319);
nor U1907 (N_1907,N_1307,N_1794);
nand U1908 (N_1908,N_1311,N_1688);
nor U1909 (N_1909,N_1655,N_1398);
and U1910 (N_1910,N_1567,N_1450);
and U1911 (N_1911,N_1330,N_1344);
and U1912 (N_1912,N_1339,N_1584);
nor U1913 (N_1913,N_1775,N_1490);
nor U1914 (N_1914,N_1691,N_1480);
and U1915 (N_1915,N_1361,N_1437);
nand U1916 (N_1916,N_1699,N_1300);
and U1917 (N_1917,N_1698,N_1230);
nor U1918 (N_1918,N_1679,N_1545);
nor U1919 (N_1919,N_1647,N_1493);
nor U1920 (N_1920,N_1384,N_1507);
and U1921 (N_1921,N_1577,N_1531);
xor U1922 (N_1922,N_1676,N_1400);
or U1923 (N_1923,N_1355,N_1269);
and U1924 (N_1924,N_1219,N_1406);
nand U1925 (N_1925,N_1766,N_1522);
nor U1926 (N_1926,N_1309,N_1418);
nand U1927 (N_1927,N_1727,N_1713);
nor U1928 (N_1928,N_1431,N_1267);
or U1929 (N_1929,N_1314,N_1712);
and U1930 (N_1930,N_1726,N_1753);
nand U1931 (N_1931,N_1675,N_1394);
or U1932 (N_1932,N_1652,N_1498);
and U1933 (N_1933,N_1298,N_1569);
and U1934 (N_1934,N_1632,N_1633);
nor U1935 (N_1935,N_1286,N_1572);
nor U1936 (N_1936,N_1366,N_1482);
and U1937 (N_1937,N_1204,N_1468);
and U1938 (N_1938,N_1686,N_1768);
and U1939 (N_1939,N_1785,N_1457);
nand U1940 (N_1940,N_1658,N_1239);
or U1941 (N_1941,N_1426,N_1646);
and U1942 (N_1942,N_1290,N_1562);
nand U1943 (N_1943,N_1576,N_1262);
and U1944 (N_1944,N_1741,N_1360);
nor U1945 (N_1945,N_1744,N_1578);
and U1946 (N_1946,N_1371,N_1568);
and U1947 (N_1947,N_1470,N_1308);
or U1948 (N_1948,N_1249,N_1500);
and U1949 (N_1949,N_1255,N_1784);
nand U1950 (N_1950,N_1217,N_1438);
nand U1951 (N_1951,N_1581,N_1542);
nand U1952 (N_1952,N_1769,N_1382);
nor U1953 (N_1953,N_1357,N_1452);
nor U1954 (N_1954,N_1210,N_1421);
nor U1955 (N_1955,N_1590,N_1654);
nor U1956 (N_1956,N_1504,N_1236);
nor U1957 (N_1957,N_1304,N_1717);
nor U1958 (N_1958,N_1510,N_1617);
nand U1959 (N_1959,N_1587,N_1524);
or U1960 (N_1960,N_1285,N_1232);
and U1961 (N_1961,N_1333,N_1626);
nand U1962 (N_1962,N_1496,N_1573);
nor U1963 (N_1963,N_1329,N_1714);
or U1964 (N_1964,N_1291,N_1318);
nor U1965 (N_1965,N_1538,N_1566);
or U1966 (N_1966,N_1475,N_1680);
and U1967 (N_1967,N_1580,N_1774);
or U1968 (N_1968,N_1793,N_1516);
and U1969 (N_1969,N_1494,N_1253);
nand U1970 (N_1970,N_1734,N_1415);
or U1971 (N_1971,N_1246,N_1600);
and U1972 (N_1972,N_1212,N_1732);
nand U1973 (N_1973,N_1746,N_1549);
nand U1974 (N_1974,N_1661,N_1513);
nand U1975 (N_1975,N_1263,N_1337);
nor U1976 (N_1976,N_1517,N_1297);
or U1977 (N_1977,N_1265,N_1659);
or U1978 (N_1978,N_1240,N_1380);
nor U1979 (N_1979,N_1553,N_1598);
and U1980 (N_1980,N_1791,N_1376);
and U1981 (N_1981,N_1388,N_1218);
and U1982 (N_1982,N_1635,N_1449);
and U1983 (N_1983,N_1221,N_1593);
or U1984 (N_1984,N_1511,N_1757);
or U1985 (N_1985,N_1765,N_1579);
nor U1986 (N_1986,N_1340,N_1409);
nand U1987 (N_1987,N_1748,N_1213);
nor U1988 (N_1988,N_1640,N_1673);
nand U1989 (N_1989,N_1685,N_1595);
or U1990 (N_1990,N_1322,N_1476);
nor U1991 (N_1991,N_1359,N_1279);
nor U1992 (N_1992,N_1328,N_1799);
xnor U1993 (N_1993,N_1541,N_1721);
nand U1994 (N_1994,N_1527,N_1299);
or U1995 (N_1995,N_1551,N_1264);
nor U1996 (N_1996,N_1316,N_1703);
or U1997 (N_1997,N_1550,N_1377);
and U1998 (N_1998,N_1228,N_1535);
nand U1999 (N_1999,N_1441,N_1594);
nor U2000 (N_2000,N_1770,N_1612);
nor U2001 (N_2001,N_1648,N_1326);
and U2002 (N_2002,N_1391,N_1605);
and U2003 (N_2003,N_1485,N_1606);
nand U2004 (N_2004,N_1792,N_1363);
and U2005 (N_2005,N_1651,N_1729);
nand U2006 (N_2006,N_1672,N_1789);
and U2007 (N_2007,N_1378,N_1557);
or U2008 (N_2008,N_1348,N_1404);
and U2009 (N_2009,N_1294,N_1282);
or U2010 (N_2010,N_1220,N_1201);
or U2011 (N_2011,N_1358,N_1465);
nor U2012 (N_2012,N_1620,N_1454);
and U2013 (N_2013,N_1639,N_1596);
or U2014 (N_2014,N_1501,N_1546);
or U2015 (N_2015,N_1408,N_1323);
and U2016 (N_2016,N_1716,N_1214);
xor U2017 (N_2017,N_1571,N_1280);
nand U2018 (N_2018,N_1272,N_1405);
or U2019 (N_2019,N_1678,N_1614);
or U2020 (N_2020,N_1518,N_1739);
nand U2021 (N_2021,N_1697,N_1399);
and U2022 (N_2022,N_1367,N_1534);
nand U2023 (N_2023,N_1643,N_1711);
nor U2024 (N_2024,N_1479,N_1742);
nor U2025 (N_2025,N_1433,N_1787);
nand U2026 (N_2026,N_1599,N_1365);
and U2027 (N_2027,N_1379,N_1420);
or U2028 (N_2028,N_1603,N_1317);
nor U2029 (N_2029,N_1222,N_1390);
nand U2030 (N_2030,N_1544,N_1385);
or U2031 (N_2031,N_1472,N_1258);
nand U2032 (N_2032,N_1389,N_1402);
and U2033 (N_2033,N_1321,N_1481);
nor U2034 (N_2034,N_1488,N_1592);
and U2035 (N_2035,N_1707,N_1610);
or U2036 (N_2036,N_1273,N_1276);
nand U2037 (N_2037,N_1555,N_1619);
xor U2038 (N_2038,N_1289,N_1644);
nor U2039 (N_2039,N_1436,N_1795);
nand U2040 (N_2040,N_1215,N_1547);
and U2041 (N_2041,N_1474,N_1200);
nor U2042 (N_2042,N_1392,N_1254);
nand U2043 (N_2043,N_1268,N_1564);
or U2044 (N_2044,N_1740,N_1749);
nand U2045 (N_2045,N_1629,N_1455);
and U2046 (N_2046,N_1736,N_1693);
and U2047 (N_2047,N_1414,N_1483);
nand U2048 (N_2048,N_1375,N_1229);
nand U2049 (N_2049,N_1618,N_1731);
or U2050 (N_2050,N_1695,N_1459);
nand U2051 (N_2051,N_1491,N_1320);
or U2052 (N_2052,N_1346,N_1447);
nand U2053 (N_2053,N_1611,N_1247);
nand U2054 (N_2054,N_1533,N_1523);
nand U2055 (N_2055,N_1463,N_1537);
xor U2056 (N_2056,N_1607,N_1667);
or U2057 (N_2057,N_1730,N_1725);
nor U2058 (N_2058,N_1499,N_1471);
and U2059 (N_2059,N_1656,N_1540);
nor U2060 (N_2060,N_1231,N_1284);
and U2061 (N_2061,N_1242,N_1492);
nor U2062 (N_2062,N_1369,N_1248);
nor U2063 (N_2063,N_1353,N_1689);
or U2064 (N_2064,N_1256,N_1356);
nor U2065 (N_2065,N_1754,N_1574);
nand U2066 (N_2066,N_1288,N_1364);
nor U2067 (N_2067,N_1692,N_1351);
nand U2068 (N_2068,N_1690,N_1235);
nand U2069 (N_2069,N_1503,N_1486);
nor U2070 (N_2070,N_1427,N_1473);
or U2071 (N_2071,N_1788,N_1758);
nand U2072 (N_2072,N_1331,N_1696);
nand U2073 (N_2073,N_1350,N_1261);
and U2074 (N_2074,N_1750,N_1422);
and U2075 (N_2075,N_1700,N_1570);
nand U2076 (N_2076,N_1342,N_1478);
nand U2077 (N_2077,N_1755,N_1458);
and U2078 (N_2078,N_1412,N_1383);
nor U2079 (N_2079,N_1207,N_1668);
and U2080 (N_2080,N_1224,N_1671);
nand U2081 (N_2081,N_1244,N_1487);
nand U2082 (N_2082,N_1722,N_1625);
and U2083 (N_2083,N_1630,N_1601);
nand U2084 (N_2084,N_1278,N_1442);
or U2085 (N_2085,N_1681,N_1773);
and U2086 (N_2086,N_1338,N_1767);
nor U2087 (N_2087,N_1796,N_1797);
and U2088 (N_2088,N_1497,N_1432);
or U2089 (N_2089,N_1561,N_1469);
and U2090 (N_2090,N_1270,N_1710);
or U2091 (N_2091,N_1720,N_1583);
nor U2092 (N_2092,N_1396,N_1701);
and U2093 (N_2093,N_1315,N_1274);
or U2094 (N_2094,N_1786,N_1370);
nor U2095 (N_2095,N_1609,N_1588);
nor U2096 (N_2096,N_1515,N_1234);
and U2097 (N_2097,N_1743,N_1653);
or U2098 (N_2098,N_1529,N_1636);
nand U2099 (N_2099,N_1752,N_1565);
or U2100 (N_2100,N_1413,N_1728);
or U2101 (N_2101,N_1224,N_1738);
nand U2102 (N_2102,N_1402,N_1420);
and U2103 (N_2103,N_1719,N_1307);
nor U2104 (N_2104,N_1275,N_1655);
nor U2105 (N_2105,N_1563,N_1435);
nor U2106 (N_2106,N_1785,N_1657);
or U2107 (N_2107,N_1328,N_1468);
nor U2108 (N_2108,N_1396,N_1441);
nand U2109 (N_2109,N_1332,N_1579);
and U2110 (N_2110,N_1738,N_1663);
or U2111 (N_2111,N_1516,N_1219);
and U2112 (N_2112,N_1635,N_1536);
and U2113 (N_2113,N_1303,N_1773);
nor U2114 (N_2114,N_1735,N_1554);
nand U2115 (N_2115,N_1789,N_1700);
or U2116 (N_2116,N_1751,N_1406);
nor U2117 (N_2117,N_1797,N_1229);
nand U2118 (N_2118,N_1334,N_1577);
and U2119 (N_2119,N_1366,N_1281);
or U2120 (N_2120,N_1357,N_1265);
or U2121 (N_2121,N_1392,N_1631);
nor U2122 (N_2122,N_1399,N_1694);
and U2123 (N_2123,N_1532,N_1382);
nand U2124 (N_2124,N_1495,N_1541);
nand U2125 (N_2125,N_1598,N_1246);
nor U2126 (N_2126,N_1355,N_1614);
and U2127 (N_2127,N_1714,N_1785);
or U2128 (N_2128,N_1619,N_1355);
and U2129 (N_2129,N_1223,N_1636);
nand U2130 (N_2130,N_1405,N_1243);
and U2131 (N_2131,N_1759,N_1306);
nor U2132 (N_2132,N_1340,N_1572);
nor U2133 (N_2133,N_1448,N_1720);
or U2134 (N_2134,N_1450,N_1215);
nand U2135 (N_2135,N_1466,N_1256);
nand U2136 (N_2136,N_1410,N_1567);
or U2137 (N_2137,N_1201,N_1464);
nor U2138 (N_2138,N_1434,N_1567);
nor U2139 (N_2139,N_1687,N_1404);
or U2140 (N_2140,N_1296,N_1558);
nand U2141 (N_2141,N_1214,N_1548);
nand U2142 (N_2142,N_1448,N_1430);
nor U2143 (N_2143,N_1661,N_1754);
nand U2144 (N_2144,N_1557,N_1453);
nor U2145 (N_2145,N_1571,N_1793);
nand U2146 (N_2146,N_1548,N_1464);
or U2147 (N_2147,N_1534,N_1315);
nand U2148 (N_2148,N_1585,N_1202);
and U2149 (N_2149,N_1721,N_1442);
and U2150 (N_2150,N_1475,N_1226);
nand U2151 (N_2151,N_1667,N_1656);
or U2152 (N_2152,N_1278,N_1628);
nand U2153 (N_2153,N_1643,N_1665);
nand U2154 (N_2154,N_1768,N_1780);
nor U2155 (N_2155,N_1446,N_1613);
xor U2156 (N_2156,N_1263,N_1399);
or U2157 (N_2157,N_1501,N_1556);
and U2158 (N_2158,N_1557,N_1675);
nand U2159 (N_2159,N_1692,N_1232);
nand U2160 (N_2160,N_1586,N_1374);
nand U2161 (N_2161,N_1493,N_1353);
or U2162 (N_2162,N_1277,N_1509);
or U2163 (N_2163,N_1371,N_1522);
nor U2164 (N_2164,N_1248,N_1226);
nand U2165 (N_2165,N_1528,N_1453);
or U2166 (N_2166,N_1542,N_1566);
nand U2167 (N_2167,N_1259,N_1621);
nor U2168 (N_2168,N_1614,N_1727);
or U2169 (N_2169,N_1370,N_1764);
nand U2170 (N_2170,N_1461,N_1259);
nor U2171 (N_2171,N_1275,N_1707);
nand U2172 (N_2172,N_1728,N_1509);
nor U2173 (N_2173,N_1524,N_1476);
nand U2174 (N_2174,N_1239,N_1243);
and U2175 (N_2175,N_1308,N_1500);
or U2176 (N_2176,N_1605,N_1504);
nor U2177 (N_2177,N_1302,N_1469);
nand U2178 (N_2178,N_1336,N_1334);
nor U2179 (N_2179,N_1320,N_1777);
or U2180 (N_2180,N_1475,N_1730);
or U2181 (N_2181,N_1556,N_1591);
nand U2182 (N_2182,N_1751,N_1341);
nor U2183 (N_2183,N_1726,N_1602);
nor U2184 (N_2184,N_1544,N_1653);
and U2185 (N_2185,N_1424,N_1547);
nand U2186 (N_2186,N_1221,N_1566);
nor U2187 (N_2187,N_1594,N_1462);
or U2188 (N_2188,N_1347,N_1746);
and U2189 (N_2189,N_1603,N_1256);
nor U2190 (N_2190,N_1234,N_1629);
and U2191 (N_2191,N_1642,N_1661);
nor U2192 (N_2192,N_1507,N_1537);
and U2193 (N_2193,N_1436,N_1628);
and U2194 (N_2194,N_1250,N_1398);
or U2195 (N_2195,N_1689,N_1775);
or U2196 (N_2196,N_1303,N_1638);
or U2197 (N_2197,N_1201,N_1519);
nor U2198 (N_2198,N_1354,N_1649);
and U2199 (N_2199,N_1695,N_1691);
and U2200 (N_2200,N_1545,N_1416);
and U2201 (N_2201,N_1790,N_1287);
and U2202 (N_2202,N_1493,N_1329);
nand U2203 (N_2203,N_1333,N_1741);
nand U2204 (N_2204,N_1275,N_1527);
or U2205 (N_2205,N_1334,N_1644);
or U2206 (N_2206,N_1326,N_1638);
and U2207 (N_2207,N_1358,N_1760);
and U2208 (N_2208,N_1536,N_1564);
nor U2209 (N_2209,N_1217,N_1710);
nand U2210 (N_2210,N_1773,N_1554);
nand U2211 (N_2211,N_1747,N_1506);
or U2212 (N_2212,N_1503,N_1294);
or U2213 (N_2213,N_1705,N_1647);
nand U2214 (N_2214,N_1233,N_1761);
nor U2215 (N_2215,N_1506,N_1209);
nor U2216 (N_2216,N_1572,N_1484);
nand U2217 (N_2217,N_1329,N_1713);
and U2218 (N_2218,N_1521,N_1449);
and U2219 (N_2219,N_1248,N_1471);
or U2220 (N_2220,N_1461,N_1716);
and U2221 (N_2221,N_1215,N_1432);
nand U2222 (N_2222,N_1437,N_1501);
or U2223 (N_2223,N_1398,N_1436);
and U2224 (N_2224,N_1430,N_1557);
nand U2225 (N_2225,N_1358,N_1214);
nand U2226 (N_2226,N_1275,N_1337);
or U2227 (N_2227,N_1375,N_1790);
nor U2228 (N_2228,N_1444,N_1458);
or U2229 (N_2229,N_1376,N_1632);
nor U2230 (N_2230,N_1385,N_1396);
or U2231 (N_2231,N_1545,N_1445);
and U2232 (N_2232,N_1766,N_1748);
and U2233 (N_2233,N_1472,N_1719);
nand U2234 (N_2234,N_1343,N_1625);
nand U2235 (N_2235,N_1351,N_1693);
nand U2236 (N_2236,N_1550,N_1563);
nand U2237 (N_2237,N_1421,N_1695);
and U2238 (N_2238,N_1392,N_1691);
nor U2239 (N_2239,N_1366,N_1227);
and U2240 (N_2240,N_1750,N_1773);
and U2241 (N_2241,N_1375,N_1525);
nor U2242 (N_2242,N_1502,N_1751);
and U2243 (N_2243,N_1400,N_1234);
nor U2244 (N_2244,N_1669,N_1363);
nor U2245 (N_2245,N_1275,N_1768);
nand U2246 (N_2246,N_1485,N_1379);
or U2247 (N_2247,N_1603,N_1628);
and U2248 (N_2248,N_1210,N_1721);
nand U2249 (N_2249,N_1281,N_1665);
and U2250 (N_2250,N_1728,N_1211);
and U2251 (N_2251,N_1523,N_1245);
xor U2252 (N_2252,N_1695,N_1209);
nand U2253 (N_2253,N_1205,N_1721);
nor U2254 (N_2254,N_1641,N_1382);
nand U2255 (N_2255,N_1431,N_1527);
and U2256 (N_2256,N_1299,N_1470);
nor U2257 (N_2257,N_1742,N_1674);
and U2258 (N_2258,N_1433,N_1518);
nor U2259 (N_2259,N_1263,N_1327);
and U2260 (N_2260,N_1207,N_1525);
and U2261 (N_2261,N_1521,N_1761);
or U2262 (N_2262,N_1202,N_1729);
nand U2263 (N_2263,N_1695,N_1625);
or U2264 (N_2264,N_1265,N_1534);
or U2265 (N_2265,N_1408,N_1566);
nor U2266 (N_2266,N_1542,N_1750);
and U2267 (N_2267,N_1579,N_1385);
nor U2268 (N_2268,N_1307,N_1328);
nand U2269 (N_2269,N_1222,N_1301);
and U2270 (N_2270,N_1578,N_1326);
or U2271 (N_2271,N_1273,N_1698);
and U2272 (N_2272,N_1447,N_1595);
nand U2273 (N_2273,N_1524,N_1321);
nor U2274 (N_2274,N_1264,N_1319);
and U2275 (N_2275,N_1492,N_1307);
and U2276 (N_2276,N_1466,N_1443);
or U2277 (N_2277,N_1527,N_1495);
nand U2278 (N_2278,N_1286,N_1624);
nor U2279 (N_2279,N_1313,N_1570);
nor U2280 (N_2280,N_1388,N_1649);
nor U2281 (N_2281,N_1625,N_1423);
nand U2282 (N_2282,N_1378,N_1738);
or U2283 (N_2283,N_1552,N_1793);
nand U2284 (N_2284,N_1288,N_1373);
nand U2285 (N_2285,N_1259,N_1469);
nand U2286 (N_2286,N_1693,N_1619);
nand U2287 (N_2287,N_1661,N_1550);
and U2288 (N_2288,N_1660,N_1507);
nand U2289 (N_2289,N_1416,N_1581);
and U2290 (N_2290,N_1738,N_1692);
and U2291 (N_2291,N_1275,N_1658);
nand U2292 (N_2292,N_1781,N_1631);
nor U2293 (N_2293,N_1541,N_1408);
or U2294 (N_2294,N_1666,N_1460);
or U2295 (N_2295,N_1416,N_1661);
and U2296 (N_2296,N_1718,N_1536);
nand U2297 (N_2297,N_1543,N_1262);
or U2298 (N_2298,N_1708,N_1733);
nand U2299 (N_2299,N_1764,N_1224);
nor U2300 (N_2300,N_1291,N_1360);
or U2301 (N_2301,N_1397,N_1729);
or U2302 (N_2302,N_1707,N_1651);
nor U2303 (N_2303,N_1469,N_1794);
or U2304 (N_2304,N_1531,N_1774);
nor U2305 (N_2305,N_1229,N_1463);
xor U2306 (N_2306,N_1382,N_1566);
nand U2307 (N_2307,N_1300,N_1710);
or U2308 (N_2308,N_1397,N_1646);
nor U2309 (N_2309,N_1320,N_1769);
nor U2310 (N_2310,N_1454,N_1682);
nand U2311 (N_2311,N_1562,N_1542);
or U2312 (N_2312,N_1559,N_1717);
or U2313 (N_2313,N_1421,N_1376);
nand U2314 (N_2314,N_1287,N_1420);
or U2315 (N_2315,N_1317,N_1781);
and U2316 (N_2316,N_1692,N_1261);
or U2317 (N_2317,N_1216,N_1550);
or U2318 (N_2318,N_1532,N_1272);
and U2319 (N_2319,N_1325,N_1639);
nor U2320 (N_2320,N_1319,N_1342);
and U2321 (N_2321,N_1280,N_1523);
nor U2322 (N_2322,N_1289,N_1358);
nor U2323 (N_2323,N_1215,N_1373);
nand U2324 (N_2324,N_1673,N_1477);
and U2325 (N_2325,N_1326,N_1621);
nand U2326 (N_2326,N_1219,N_1571);
and U2327 (N_2327,N_1693,N_1416);
nand U2328 (N_2328,N_1656,N_1356);
or U2329 (N_2329,N_1313,N_1293);
or U2330 (N_2330,N_1574,N_1200);
and U2331 (N_2331,N_1559,N_1361);
nor U2332 (N_2332,N_1700,N_1320);
nor U2333 (N_2333,N_1613,N_1370);
nand U2334 (N_2334,N_1554,N_1422);
nand U2335 (N_2335,N_1314,N_1671);
and U2336 (N_2336,N_1648,N_1523);
nand U2337 (N_2337,N_1732,N_1218);
and U2338 (N_2338,N_1647,N_1307);
nor U2339 (N_2339,N_1365,N_1376);
nor U2340 (N_2340,N_1636,N_1270);
or U2341 (N_2341,N_1586,N_1377);
or U2342 (N_2342,N_1429,N_1589);
and U2343 (N_2343,N_1317,N_1441);
nand U2344 (N_2344,N_1775,N_1553);
nand U2345 (N_2345,N_1235,N_1395);
or U2346 (N_2346,N_1773,N_1406);
nand U2347 (N_2347,N_1234,N_1353);
and U2348 (N_2348,N_1736,N_1647);
or U2349 (N_2349,N_1479,N_1758);
or U2350 (N_2350,N_1545,N_1309);
nand U2351 (N_2351,N_1425,N_1749);
or U2352 (N_2352,N_1645,N_1253);
nand U2353 (N_2353,N_1528,N_1344);
nand U2354 (N_2354,N_1258,N_1544);
or U2355 (N_2355,N_1486,N_1727);
and U2356 (N_2356,N_1531,N_1683);
or U2357 (N_2357,N_1279,N_1521);
and U2358 (N_2358,N_1390,N_1647);
nand U2359 (N_2359,N_1504,N_1674);
nor U2360 (N_2360,N_1426,N_1469);
nor U2361 (N_2361,N_1481,N_1581);
nor U2362 (N_2362,N_1573,N_1226);
or U2363 (N_2363,N_1722,N_1533);
nand U2364 (N_2364,N_1759,N_1583);
nand U2365 (N_2365,N_1486,N_1775);
or U2366 (N_2366,N_1679,N_1699);
nand U2367 (N_2367,N_1201,N_1505);
nand U2368 (N_2368,N_1543,N_1757);
nor U2369 (N_2369,N_1659,N_1686);
or U2370 (N_2370,N_1572,N_1559);
and U2371 (N_2371,N_1631,N_1468);
xor U2372 (N_2372,N_1702,N_1414);
and U2373 (N_2373,N_1632,N_1623);
nor U2374 (N_2374,N_1423,N_1406);
or U2375 (N_2375,N_1612,N_1347);
nor U2376 (N_2376,N_1668,N_1694);
or U2377 (N_2377,N_1569,N_1415);
nor U2378 (N_2378,N_1526,N_1248);
nand U2379 (N_2379,N_1234,N_1491);
xnor U2380 (N_2380,N_1636,N_1368);
nor U2381 (N_2381,N_1363,N_1378);
or U2382 (N_2382,N_1510,N_1480);
nand U2383 (N_2383,N_1480,N_1773);
nand U2384 (N_2384,N_1455,N_1321);
or U2385 (N_2385,N_1739,N_1775);
or U2386 (N_2386,N_1726,N_1368);
and U2387 (N_2387,N_1285,N_1501);
or U2388 (N_2388,N_1475,N_1374);
nand U2389 (N_2389,N_1705,N_1330);
and U2390 (N_2390,N_1244,N_1605);
or U2391 (N_2391,N_1650,N_1495);
nand U2392 (N_2392,N_1639,N_1267);
and U2393 (N_2393,N_1692,N_1451);
or U2394 (N_2394,N_1250,N_1207);
or U2395 (N_2395,N_1482,N_1466);
or U2396 (N_2396,N_1577,N_1309);
xor U2397 (N_2397,N_1231,N_1404);
and U2398 (N_2398,N_1763,N_1440);
nor U2399 (N_2399,N_1662,N_1549);
and U2400 (N_2400,N_2078,N_2112);
and U2401 (N_2401,N_2229,N_1960);
or U2402 (N_2402,N_2309,N_1913);
nor U2403 (N_2403,N_1869,N_2194);
or U2404 (N_2404,N_1995,N_1966);
nand U2405 (N_2405,N_2014,N_1837);
nor U2406 (N_2406,N_2137,N_2086);
or U2407 (N_2407,N_2385,N_2381);
nor U2408 (N_2408,N_1959,N_1862);
and U2409 (N_2409,N_1917,N_2280);
nand U2410 (N_2410,N_2089,N_2173);
nand U2411 (N_2411,N_2267,N_2313);
nor U2412 (N_2412,N_1934,N_2247);
or U2413 (N_2413,N_2343,N_1908);
nand U2414 (N_2414,N_2205,N_2043);
and U2415 (N_2415,N_2350,N_2285);
nand U2416 (N_2416,N_2379,N_2045);
or U2417 (N_2417,N_1870,N_1859);
nand U2418 (N_2418,N_2129,N_2212);
and U2419 (N_2419,N_2095,N_2273);
and U2420 (N_2420,N_2087,N_2241);
or U2421 (N_2421,N_1809,N_2115);
nor U2422 (N_2422,N_2314,N_2103);
nor U2423 (N_2423,N_1979,N_2189);
nor U2424 (N_2424,N_2344,N_2026);
xor U2425 (N_2425,N_2196,N_2307);
or U2426 (N_2426,N_2108,N_2353);
nor U2427 (N_2427,N_2066,N_2370);
and U2428 (N_2428,N_1834,N_2117);
and U2429 (N_2429,N_2050,N_2101);
or U2430 (N_2430,N_1986,N_2223);
nor U2431 (N_2431,N_2290,N_1932);
nand U2432 (N_2432,N_2039,N_2292);
or U2433 (N_2433,N_2357,N_1806);
or U2434 (N_2434,N_2220,N_2358);
nor U2435 (N_2435,N_2080,N_2021);
nor U2436 (N_2436,N_1852,N_2148);
and U2437 (N_2437,N_2378,N_1849);
and U2438 (N_2438,N_1897,N_2305);
xor U2439 (N_2439,N_2393,N_1952);
and U2440 (N_2440,N_1984,N_2107);
nor U2441 (N_2441,N_2396,N_1957);
nand U2442 (N_2442,N_1896,N_2061);
or U2443 (N_2443,N_2372,N_2152);
nor U2444 (N_2444,N_2252,N_2369);
and U2445 (N_2445,N_2338,N_2232);
and U2446 (N_2446,N_2085,N_2142);
and U2447 (N_2447,N_2111,N_2371);
nand U2448 (N_2448,N_2074,N_1976);
nor U2449 (N_2449,N_1983,N_2394);
nor U2450 (N_2450,N_1882,N_2254);
and U2451 (N_2451,N_1999,N_2041);
nand U2452 (N_2452,N_1991,N_1839);
nand U2453 (N_2453,N_2166,N_1945);
or U2454 (N_2454,N_1969,N_1821);
nand U2455 (N_2455,N_2055,N_1866);
nand U2456 (N_2456,N_1864,N_1878);
nor U2457 (N_2457,N_2183,N_2013);
nor U2458 (N_2458,N_1916,N_2335);
nand U2459 (N_2459,N_2174,N_2002);
or U2460 (N_2460,N_2195,N_2236);
xor U2461 (N_2461,N_1985,N_1840);
nand U2462 (N_2462,N_2118,N_2160);
nor U2463 (N_2463,N_2368,N_2054);
and U2464 (N_2464,N_2058,N_1954);
and U2465 (N_2465,N_2263,N_1965);
nor U2466 (N_2466,N_1915,N_2298);
nand U2467 (N_2467,N_1838,N_1816);
nor U2468 (N_2468,N_1938,N_2068);
nor U2469 (N_2469,N_1876,N_2375);
or U2470 (N_2470,N_1935,N_2181);
nand U2471 (N_2471,N_2168,N_2059);
nor U2472 (N_2472,N_2145,N_2144);
or U2473 (N_2473,N_2178,N_2186);
nand U2474 (N_2474,N_2215,N_2354);
nor U2475 (N_2475,N_2076,N_2140);
nor U2476 (N_2476,N_2128,N_1970);
or U2477 (N_2477,N_2270,N_2139);
or U2478 (N_2478,N_1899,N_2034);
nand U2479 (N_2479,N_2345,N_1804);
or U2480 (N_2480,N_2098,N_2193);
nor U2481 (N_2481,N_2218,N_2106);
and U2482 (N_2482,N_1843,N_2114);
and U2483 (N_2483,N_1922,N_1868);
nand U2484 (N_2484,N_2207,N_2213);
and U2485 (N_2485,N_2015,N_1937);
and U2486 (N_2486,N_2093,N_2006);
or U2487 (N_2487,N_1972,N_2356);
or U2488 (N_2488,N_1883,N_2238);
or U2489 (N_2489,N_2274,N_2003);
or U2490 (N_2490,N_2242,N_2102);
or U2491 (N_2491,N_1822,N_2262);
and U2492 (N_2492,N_2303,N_2047);
nand U2493 (N_2493,N_1875,N_1841);
and U2494 (N_2494,N_2395,N_2032);
nor U2495 (N_2495,N_1955,N_1818);
nand U2496 (N_2496,N_2294,N_2233);
or U2497 (N_2497,N_1953,N_2293);
or U2498 (N_2498,N_1973,N_2031);
nand U2499 (N_2499,N_2105,N_2022);
or U2500 (N_2500,N_1902,N_2188);
nand U2501 (N_2501,N_1963,N_2020);
or U2502 (N_2502,N_1924,N_2190);
nand U2503 (N_2503,N_1831,N_1828);
and U2504 (N_2504,N_2033,N_2306);
and U2505 (N_2505,N_2200,N_2230);
xnor U2506 (N_2506,N_1989,N_2038);
nor U2507 (N_2507,N_2301,N_2170);
nor U2508 (N_2508,N_1962,N_2341);
nand U2509 (N_2509,N_1826,N_1964);
and U2510 (N_2510,N_2390,N_2235);
nor U2511 (N_2511,N_1860,N_1884);
nor U2512 (N_2512,N_1853,N_2197);
or U2513 (N_2513,N_2199,N_1880);
nand U2514 (N_2514,N_2126,N_1961);
nor U2515 (N_2515,N_2081,N_1944);
nand U2516 (N_2516,N_2127,N_2042);
nor U2517 (N_2517,N_2175,N_1858);
or U2518 (N_2518,N_1927,N_2284);
or U2519 (N_2519,N_2090,N_2261);
nor U2520 (N_2520,N_2179,N_2062);
xnor U2521 (N_2521,N_2184,N_1855);
and U2522 (N_2522,N_1997,N_2219);
or U2523 (N_2523,N_2163,N_2147);
nor U2524 (N_2524,N_2304,N_2167);
nand U2525 (N_2525,N_2332,N_1846);
or U2526 (N_2526,N_2100,N_1836);
nor U2527 (N_2527,N_2388,N_2326);
or U2528 (N_2528,N_2330,N_2329);
nand U2529 (N_2529,N_2282,N_2323);
or U2530 (N_2530,N_2311,N_2331);
nor U2531 (N_2531,N_2281,N_2151);
or U2532 (N_2532,N_2214,N_2094);
and U2533 (N_2533,N_2365,N_2347);
and U2534 (N_2534,N_1856,N_1819);
nor U2535 (N_2535,N_2071,N_2243);
and U2536 (N_2536,N_1851,N_2245);
and U2537 (N_2537,N_1981,N_1912);
nand U2538 (N_2538,N_2134,N_2130);
nand U2539 (N_2539,N_1811,N_1921);
nor U2540 (N_2540,N_2237,N_1803);
nor U2541 (N_2541,N_2008,N_2052);
and U2542 (N_2542,N_2367,N_2053);
nand U2543 (N_2543,N_2383,N_2122);
and U2544 (N_2544,N_2096,N_2072);
nand U2545 (N_2545,N_2192,N_2120);
nand U2546 (N_2546,N_2024,N_2209);
nand U2547 (N_2547,N_1971,N_2362);
nand U2548 (N_2548,N_2239,N_2234);
and U2549 (N_2549,N_2377,N_2222);
or U2550 (N_2550,N_2269,N_2333);
nor U2551 (N_2551,N_1874,N_2392);
or U2552 (N_2552,N_2016,N_2202);
nor U2553 (N_2553,N_2224,N_1990);
and U2554 (N_2554,N_1808,N_1926);
nor U2555 (N_2555,N_2391,N_2386);
nor U2556 (N_2556,N_2155,N_2321);
and U2557 (N_2557,N_2320,N_1911);
nand U2558 (N_2558,N_1936,N_2005);
nand U2559 (N_2559,N_1919,N_2275);
or U2560 (N_2560,N_2176,N_2000);
and U2561 (N_2561,N_2069,N_2044);
nand U2562 (N_2562,N_2240,N_2012);
nand U2563 (N_2563,N_2374,N_1861);
or U2564 (N_2564,N_1890,N_2171);
nor U2565 (N_2565,N_2056,N_1877);
nand U2566 (N_2566,N_2387,N_1928);
and U2567 (N_2567,N_1873,N_2327);
nand U2568 (N_2568,N_1891,N_2091);
nor U2569 (N_2569,N_1980,N_2116);
and U2570 (N_2570,N_2060,N_2373);
nor U2571 (N_2571,N_2035,N_1823);
nor U2572 (N_2572,N_2177,N_1865);
and U2573 (N_2573,N_2077,N_2048);
and U2574 (N_2574,N_1845,N_2255);
nor U2575 (N_2575,N_2113,N_1904);
and U2576 (N_2576,N_1894,N_2159);
nor U2577 (N_2577,N_1923,N_1886);
nor U2578 (N_2578,N_2266,N_2040);
and U2579 (N_2579,N_2380,N_1910);
and U2580 (N_2580,N_2007,N_1847);
nand U2581 (N_2581,N_2110,N_2182);
or U2582 (N_2582,N_1881,N_1832);
or U2583 (N_2583,N_2231,N_1988);
nor U2584 (N_2584,N_2153,N_2083);
nor U2585 (N_2585,N_2337,N_2019);
nand U2586 (N_2586,N_2185,N_1950);
nor U2587 (N_2587,N_2297,N_1898);
or U2588 (N_2588,N_1968,N_1978);
or U2589 (N_2589,N_1802,N_2289);
nand U2590 (N_2590,N_2271,N_2011);
nand U2591 (N_2591,N_2010,N_2366);
nor U2592 (N_2592,N_2121,N_2030);
nand U2593 (N_2593,N_2322,N_1998);
and U2594 (N_2594,N_2180,N_1824);
nor U2595 (N_2595,N_1889,N_1958);
or U2596 (N_2596,N_2064,N_2328);
nor U2597 (N_2597,N_1887,N_2300);
nor U2598 (N_2598,N_2316,N_1967);
nand U2599 (N_2599,N_2154,N_2291);
and U2600 (N_2600,N_1920,N_1918);
and U2601 (N_2601,N_1830,N_1949);
and U2602 (N_2602,N_1951,N_2135);
nor U2603 (N_2603,N_1933,N_2250);
nor U2604 (N_2604,N_1879,N_2248);
nor U2605 (N_2605,N_1807,N_2027);
nand U2606 (N_2606,N_2260,N_1892);
nand U2607 (N_2607,N_1929,N_1871);
and U2608 (N_2608,N_1942,N_1931);
nor U2609 (N_2609,N_2187,N_2227);
nand U2610 (N_2610,N_1827,N_2226);
or U2611 (N_2611,N_2208,N_2302);
nor U2612 (N_2612,N_2063,N_1941);
nor U2613 (N_2613,N_2123,N_2259);
nor U2614 (N_2614,N_1914,N_1854);
nand U2615 (N_2615,N_2288,N_1940);
nand U2616 (N_2616,N_2004,N_2143);
or U2617 (N_2617,N_2399,N_2308);
nor U2618 (N_2618,N_1895,N_2310);
or U2619 (N_2619,N_1906,N_2299);
and U2620 (N_2620,N_2109,N_1948);
nand U2621 (N_2621,N_1813,N_2075);
and U2622 (N_2622,N_2169,N_2049);
nand U2623 (N_2623,N_2162,N_2324);
and U2624 (N_2624,N_2018,N_2277);
nand U2625 (N_2625,N_1850,N_2295);
nor U2626 (N_2626,N_1817,N_1842);
nor U2627 (N_2627,N_2336,N_1974);
or U2628 (N_2628,N_1800,N_2256);
nand U2629 (N_2629,N_1982,N_2206);
and U2630 (N_2630,N_2272,N_2073);
nor U2631 (N_2631,N_1867,N_1872);
nor U2632 (N_2632,N_1975,N_2037);
nor U2633 (N_2633,N_2001,N_1801);
or U2634 (N_2634,N_2092,N_2246);
or U2635 (N_2635,N_2104,N_2172);
or U2636 (N_2636,N_2191,N_2161);
and U2637 (N_2637,N_2067,N_2346);
nor U2638 (N_2638,N_2351,N_1925);
or U2639 (N_2639,N_2257,N_2070);
nand U2640 (N_2640,N_2082,N_2398);
or U2641 (N_2641,N_1812,N_2009);
nor U2642 (N_2642,N_2216,N_2023);
and U2643 (N_2643,N_1900,N_2244);
or U2644 (N_2644,N_2349,N_2164);
or U2645 (N_2645,N_2251,N_2132);
nand U2646 (N_2646,N_2057,N_2340);
or U2647 (N_2647,N_2228,N_2384);
nor U2648 (N_2648,N_2287,N_2217);
or U2649 (N_2649,N_2258,N_2141);
or U2650 (N_2650,N_2025,N_2296);
or U2651 (N_2651,N_2119,N_2125);
nand U2652 (N_2652,N_2158,N_2286);
or U2653 (N_2653,N_1901,N_2278);
and U2654 (N_2654,N_2150,N_1888);
and U2655 (N_2655,N_2312,N_1810);
and U2656 (N_2656,N_1947,N_2319);
or U2657 (N_2657,N_1829,N_2265);
or U2658 (N_2658,N_2097,N_1893);
nand U2659 (N_2659,N_2211,N_2317);
and U2660 (N_2660,N_2382,N_1930);
or U2661 (N_2661,N_1820,N_2325);
nand U2662 (N_2662,N_1835,N_1909);
or U2663 (N_2663,N_2028,N_1833);
nor U2664 (N_2664,N_1848,N_2363);
or U2665 (N_2665,N_2157,N_2279);
or U2666 (N_2666,N_2389,N_2355);
and U2667 (N_2667,N_2029,N_1939);
nor U2668 (N_2668,N_1805,N_2221);
and U2669 (N_2669,N_2315,N_2051);
nand U2670 (N_2670,N_2133,N_1993);
nand U2671 (N_2671,N_2201,N_1946);
nor U2672 (N_2672,N_2165,N_2360);
nor U2673 (N_2673,N_2036,N_2334);
or U2674 (N_2674,N_2079,N_2376);
nand U2675 (N_2675,N_1814,N_2364);
and U2676 (N_2676,N_1943,N_2198);
nand U2677 (N_2677,N_1857,N_2352);
and U2678 (N_2678,N_2397,N_2088);
nor U2679 (N_2679,N_2318,N_2268);
nor U2680 (N_2680,N_2348,N_1885);
and U2681 (N_2681,N_2099,N_2225);
nand U2682 (N_2682,N_2264,N_2017);
nand U2683 (N_2683,N_2136,N_1977);
or U2684 (N_2684,N_2065,N_2210);
nand U2685 (N_2685,N_1907,N_1815);
nor U2686 (N_2686,N_2283,N_2149);
and U2687 (N_2687,N_2359,N_2249);
and U2688 (N_2688,N_2276,N_2156);
and U2689 (N_2689,N_1996,N_2138);
nor U2690 (N_2690,N_2253,N_2203);
nand U2691 (N_2691,N_2204,N_2084);
and U2692 (N_2692,N_1994,N_1987);
nand U2693 (N_2693,N_1956,N_2361);
nand U2694 (N_2694,N_2342,N_1903);
nor U2695 (N_2695,N_1844,N_1992);
nor U2696 (N_2696,N_1905,N_2146);
or U2697 (N_2697,N_2339,N_1863);
nand U2698 (N_2698,N_2046,N_2131);
or U2699 (N_2699,N_1825,N_2124);
or U2700 (N_2700,N_2121,N_2380);
nor U2701 (N_2701,N_1870,N_2345);
and U2702 (N_2702,N_2238,N_1823);
nor U2703 (N_2703,N_2276,N_2143);
or U2704 (N_2704,N_2006,N_2132);
nor U2705 (N_2705,N_2012,N_2382);
nand U2706 (N_2706,N_1803,N_2279);
nand U2707 (N_2707,N_2155,N_2306);
nor U2708 (N_2708,N_1852,N_2128);
and U2709 (N_2709,N_2359,N_2319);
or U2710 (N_2710,N_2199,N_2284);
or U2711 (N_2711,N_2250,N_2091);
nand U2712 (N_2712,N_1964,N_2288);
nand U2713 (N_2713,N_1818,N_2026);
or U2714 (N_2714,N_1861,N_2349);
or U2715 (N_2715,N_1824,N_2042);
nor U2716 (N_2716,N_2153,N_2036);
nand U2717 (N_2717,N_1816,N_1991);
and U2718 (N_2718,N_2284,N_1805);
or U2719 (N_2719,N_2020,N_2190);
or U2720 (N_2720,N_1897,N_2028);
nand U2721 (N_2721,N_2375,N_1957);
nand U2722 (N_2722,N_2152,N_2350);
nor U2723 (N_2723,N_2272,N_1916);
and U2724 (N_2724,N_1878,N_1939);
or U2725 (N_2725,N_1916,N_1932);
nand U2726 (N_2726,N_2090,N_2213);
or U2727 (N_2727,N_1844,N_2085);
or U2728 (N_2728,N_1932,N_2344);
nand U2729 (N_2729,N_1951,N_1887);
nand U2730 (N_2730,N_2095,N_1936);
and U2731 (N_2731,N_1808,N_2186);
and U2732 (N_2732,N_2267,N_1855);
nor U2733 (N_2733,N_2291,N_2359);
nor U2734 (N_2734,N_2373,N_2005);
nand U2735 (N_2735,N_2345,N_2343);
and U2736 (N_2736,N_2264,N_2071);
nor U2737 (N_2737,N_1800,N_2330);
or U2738 (N_2738,N_1812,N_1900);
nand U2739 (N_2739,N_2048,N_2313);
nor U2740 (N_2740,N_2133,N_2364);
nor U2741 (N_2741,N_1902,N_2382);
nand U2742 (N_2742,N_2066,N_2337);
nand U2743 (N_2743,N_2254,N_2047);
or U2744 (N_2744,N_2006,N_2294);
nor U2745 (N_2745,N_1925,N_2014);
nor U2746 (N_2746,N_2282,N_2329);
nor U2747 (N_2747,N_1853,N_2211);
and U2748 (N_2748,N_2088,N_1880);
or U2749 (N_2749,N_1878,N_2108);
or U2750 (N_2750,N_1857,N_2377);
and U2751 (N_2751,N_1946,N_2357);
and U2752 (N_2752,N_2317,N_1915);
nor U2753 (N_2753,N_1901,N_2199);
and U2754 (N_2754,N_2154,N_1910);
nand U2755 (N_2755,N_2188,N_2361);
nor U2756 (N_2756,N_2101,N_2296);
and U2757 (N_2757,N_2253,N_2063);
or U2758 (N_2758,N_2163,N_2214);
nand U2759 (N_2759,N_2213,N_2264);
and U2760 (N_2760,N_2192,N_2056);
and U2761 (N_2761,N_1817,N_2352);
and U2762 (N_2762,N_2102,N_1854);
or U2763 (N_2763,N_1847,N_2325);
and U2764 (N_2764,N_1850,N_1905);
or U2765 (N_2765,N_1923,N_2179);
nand U2766 (N_2766,N_2098,N_2077);
nand U2767 (N_2767,N_2136,N_2297);
nand U2768 (N_2768,N_2209,N_2053);
or U2769 (N_2769,N_2376,N_2048);
and U2770 (N_2770,N_2275,N_1960);
and U2771 (N_2771,N_1919,N_2318);
nor U2772 (N_2772,N_2294,N_2164);
and U2773 (N_2773,N_2185,N_2078);
and U2774 (N_2774,N_2222,N_2056);
or U2775 (N_2775,N_2120,N_2063);
nand U2776 (N_2776,N_1838,N_2076);
nand U2777 (N_2777,N_2177,N_1900);
and U2778 (N_2778,N_2023,N_2210);
and U2779 (N_2779,N_1894,N_2380);
or U2780 (N_2780,N_1809,N_2194);
or U2781 (N_2781,N_2281,N_2172);
xor U2782 (N_2782,N_2170,N_1878);
and U2783 (N_2783,N_2365,N_2396);
or U2784 (N_2784,N_1945,N_2129);
or U2785 (N_2785,N_1872,N_1804);
nor U2786 (N_2786,N_1952,N_2309);
nor U2787 (N_2787,N_1870,N_1961);
and U2788 (N_2788,N_1949,N_1828);
and U2789 (N_2789,N_1845,N_2246);
and U2790 (N_2790,N_2346,N_2052);
and U2791 (N_2791,N_2235,N_1930);
nor U2792 (N_2792,N_1915,N_2158);
xnor U2793 (N_2793,N_2122,N_1986);
nand U2794 (N_2794,N_2359,N_2041);
or U2795 (N_2795,N_2319,N_2382);
nor U2796 (N_2796,N_2255,N_2296);
nor U2797 (N_2797,N_2204,N_2232);
or U2798 (N_2798,N_1921,N_2171);
nand U2799 (N_2799,N_1976,N_2352);
nor U2800 (N_2800,N_1914,N_1951);
or U2801 (N_2801,N_2275,N_2149);
nor U2802 (N_2802,N_1995,N_1879);
nor U2803 (N_2803,N_2260,N_2152);
or U2804 (N_2804,N_2315,N_2381);
nand U2805 (N_2805,N_2316,N_2217);
or U2806 (N_2806,N_2393,N_2394);
nor U2807 (N_2807,N_2160,N_2297);
nand U2808 (N_2808,N_1962,N_2372);
nand U2809 (N_2809,N_2249,N_1809);
or U2810 (N_2810,N_2316,N_1824);
and U2811 (N_2811,N_1965,N_2186);
or U2812 (N_2812,N_2211,N_1892);
nor U2813 (N_2813,N_2189,N_1857);
or U2814 (N_2814,N_2069,N_2065);
or U2815 (N_2815,N_1868,N_2188);
nand U2816 (N_2816,N_1936,N_2047);
nor U2817 (N_2817,N_2089,N_1889);
nand U2818 (N_2818,N_2325,N_1875);
or U2819 (N_2819,N_1995,N_2344);
nand U2820 (N_2820,N_1838,N_1810);
nor U2821 (N_2821,N_2239,N_2284);
nor U2822 (N_2822,N_2262,N_2396);
and U2823 (N_2823,N_2306,N_2066);
and U2824 (N_2824,N_2003,N_1860);
nand U2825 (N_2825,N_2272,N_2006);
or U2826 (N_2826,N_2355,N_2371);
nand U2827 (N_2827,N_1846,N_1823);
and U2828 (N_2828,N_2185,N_2260);
or U2829 (N_2829,N_2204,N_2202);
nor U2830 (N_2830,N_2046,N_2389);
and U2831 (N_2831,N_2249,N_2227);
nor U2832 (N_2832,N_2301,N_1842);
xnor U2833 (N_2833,N_2267,N_1840);
and U2834 (N_2834,N_2312,N_2068);
nor U2835 (N_2835,N_2351,N_2089);
or U2836 (N_2836,N_1903,N_2105);
nor U2837 (N_2837,N_1946,N_2270);
or U2838 (N_2838,N_2361,N_1824);
and U2839 (N_2839,N_2103,N_2362);
nor U2840 (N_2840,N_1920,N_1914);
or U2841 (N_2841,N_2005,N_1865);
or U2842 (N_2842,N_2116,N_2069);
and U2843 (N_2843,N_1810,N_1828);
or U2844 (N_2844,N_2270,N_2227);
nor U2845 (N_2845,N_2256,N_2129);
and U2846 (N_2846,N_2024,N_1973);
or U2847 (N_2847,N_2387,N_2354);
nand U2848 (N_2848,N_1890,N_2117);
or U2849 (N_2849,N_2151,N_1816);
or U2850 (N_2850,N_2122,N_2177);
nor U2851 (N_2851,N_2192,N_1896);
nor U2852 (N_2852,N_2364,N_2181);
nand U2853 (N_2853,N_1849,N_2298);
and U2854 (N_2854,N_1887,N_2034);
nand U2855 (N_2855,N_2109,N_1810);
nor U2856 (N_2856,N_2301,N_2050);
and U2857 (N_2857,N_1907,N_1915);
or U2858 (N_2858,N_2322,N_2111);
nor U2859 (N_2859,N_2235,N_2004);
nor U2860 (N_2860,N_2384,N_2337);
and U2861 (N_2861,N_2279,N_2212);
nand U2862 (N_2862,N_2101,N_2383);
nand U2863 (N_2863,N_1959,N_1961);
nand U2864 (N_2864,N_2184,N_2081);
nand U2865 (N_2865,N_2249,N_2391);
nand U2866 (N_2866,N_1816,N_2170);
and U2867 (N_2867,N_2199,N_2304);
or U2868 (N_2868,N_1903,N_2077);
and U2869 (N_2869,N_2350,N_1939);
or U2870 (N_2870,N_2054,N_1948);
nand U2871 (N_2871,N_1873,N_2137);
and U2872 (N_2872,N_2028,N_1896);
nand U2873 (N_2873,N_1965,N_2044);
nor U2874 (N_2874,N_1953,N_2196);
nand U2875 (N_2875,N_2072,N_1872);
nand U2876 (N_2876,N_2186,N_2086);
nand U2877 (N_2877,N_2348,N_2059);
or U2878 (N_2878,N_1998,N_2373);
nor U2879 (N_2879,N_1905,N_1809);
xor U2880 (N_2880,N_2123,N_1942);
nand U2881 (N_2881,N_1910,N_2302);
nor U2882 (N_2882,N_1824,N_1907);
nor U2883 (N_2883,N_1997,N_1873);
and U2884 (N_2884,N_1944,N_2214);
and U2885 (N_2885,N_2190,N_2086);
nor U2886 (N_2886,N_2365,N_2318);
nand U2887 (N_2887,N_1885,N_2263);
nand U2888 (N_2888,N_1956,N_2225);
nor U2889 (N_2889,N_1917,N_1874);
and U2890 (N_2890,N_2369,N_2280);
and U2891 (N_2891,N_2250,N_1998);
nor U2892 (N_2892,N_1856,N_2344);
nor U2893 (N_2893,N_2376,N_2360);
and U2894 (N_2894,N_2093,N_2129);
and U2895 (N_2895,N_1864,N_1976);
nand U2896 (N_2896,N_2130,N_2381);
nand U2897 (N_2897,N_1942,N_2098);
or U2898 (N_2898,N_1970,N_1865);
or U2899 (N_2899,N_2207,N_2198);
nor U2900 (N_2900,N_2253,N_1838);
or U2901 (N_2901,N_2032,N_2180);
or U2902 (N_2902,N_1838,N_2046);
nand U2903 (N_2903,N_1921,N_2364);
or U2904 (N_2904,N_1812,N_2240);
nand U2905 (N_2905,N_2367,N_1978);
nor U2906 (N_2906,N_2042,N_2116);
nand U2907 (N_2907,N_1903,N_2208);
nand U2908 (N_2908,N_2305,N_2131);
and U2909 (N_2909,N_2150,N_2117);
nor U2910 (N_2910,N_2316,N_2081);
nand U2911 (N_2911,N_1992,N_2053);
nand U2912 (N_2912,N_2326,N_1969);
and U2913 (N_2913,N_1819,N_1820);
or U2914 (N_2914,N_1917,N_2115);
nand U2915 (N_2915,N_2176,N_2170);
nand U2916 (N_2916,N_1994,N_2222);
nor U2917 (N_2917,N_2313,N_1841);
and U2918 (N_2918,N_2335,N_2314);
or U2919 (N_2919,N_2226,N_1974);
nor U2920 (N_2920,N_2164,N_2360);
nor U2921 (N_2921,N_1947,N_2253);
nor U2922 (N_2922,N_2294,N_2305);
or U2923 (N_2923,N_2166,N_2225);
and U2924 (N_2924,N_2390,N_1890);
nand U2925 (N_2925,N_1971,N_2167);
nand U2926 (N_2926,N_1885,N_2346);
nand U2927 (N_2927,N_2071,N_2387);
nor U2928 (N_2928,N_1995,N_1864);
or U2929 (N_2929,N_2055,N_1952);
and U2930 (N_2930,N_1852,N_1868);
or U2931 (N_2931,N_1973,N_2387);
and U2932 (N_2932,N_2206,N_2319);
and U2933 (N_2933,N_2207,N_2197);
and U2934 (N_2934,N_1907,N_2342);
and U2935 (N_2935,N_2229,N_1830);
and U2936 (N_2936,N_2149,N_2056);
nand U2937 (N_2937,N_1891,N_1968);
nand U2938 (N_2938,N_1884,N_1922);
nand U2939 (N_2939,N_2293,N_1830);
and U2940 (N_2940,N_2132,N_1951);
nand U2941 (N_2941,N_1922,N_2044);
nor U2942 (N_2942,N_1991,N_1892);
nor U2943 (N_2943,N_2164,N_1959);
nand U2944 (N_2944,N_2105,N_1987);
nand U2945 (N_2945,N_2103,N_2347);
or U2946 (N_2946,N_2242,N_2031);
and U2947 (N_2947,N_1803,N_1839);
nor U2948 (N_2948,N_2081,N_2377);
nand U2949 (N_2949,N_1936,N_2239);
or U2950 (N_2950,N_2335,N_2065);
nor U2951 (N_2951,N_1833,N_1872);
and U2952 (N_2952,N_1935,N_2270);
or U2953 (N_2953,N_2143,N_1998);
and U2954 (N_2954,N_2124,N_2174);
or U2955 (N_2955,N_2132,N_1804);
nor U2956 (N_2956,N_1832,N_2190);
or U2957 (N_2957,N_2289,N_2154);
nand U2958 (N_2958,N_2282,N_2053);
or U2959 (N_2959,N_2080,N_2317);
nand U2960 (N_2960,N_1977,N_1969);
or U2961 (N_2961,N_2159,N_2297);
xor U2962 (N_2962,N_2293,N_2209);
or U2963 (N_2963,N_2345,N_2089);
nand U2964 (N_2964,N_2168,N_2099);
nor U2965 (N_2965,N_2329,N_2291);
and U2966 (N_2966,N_1869,N_2209);
nand U2967 (N_2967,N_2054,N_1870);
nor U2968 (N_2968,N_2163,N_1965);
nand U2969 (N_2969,N_1909,N_2221);
or U2970 (N_2970,N_2022,N_2306);
nand U2971 (N_2971,N_2391,N_2257);
xnor U2972 (N_2972,N_2314,N_2101);
or U2973 (N_2973,N_2391,N_1997);
nor U2974 (N_2974,N_1875,N_2032);
or U2975 (N_2975,N_1826,N_2263);
nand U2976 (N_2976,N_1806,N_1812);
nor U2977 (N_2977,N_1811,N_2333);
nand U2978 (N_2978,N_2017,N_2326);
or U2979 (N_2979,N_2009,N_2346);
and U2980 (N_2980,N_1826,N_2295);
or U2981 (N_2981,N_2339,N_2103);
or U2982 (N_2982,N_1829,N_2269);
and U2983 (N_2983,N_2373,N_2296);
nand U2984 (N_2984,N_2065,N_2044);
nand U2985 (N_2985,N_1821,N_1900);
and U2986 (N_2986,N_2222,N_2025);
or U2987 (N_2987,N_2035,N_2066);
or U2988 (N_2988,N_2110,N_1945);
and U2989 (N_2989,N_2318,N_2078);
or U2990 (N_2990,N_2037,N_2141);
nand U2991 (N_2991,N_2201,N_2015);
nor U2992 (N_2992,N_2392,N_2188);
and U2993 (N_2993,N_2212,N_2197);
nand U2994 (N_2994,N_1942,N_2208);
or U2995 (N_2995,N_2020,N_2316);
nand U2996 (N_2996,N_2166,N_2172);
and U2997 (N_2997,N_2057,N_2122);
and U2998 (N_2998,N_2327,N_2025);
nor U2999 (N_2999,N_2065,N_2348);
or UO_0 (O_0,N_2626,N_2559);
or UO_1 (O_1,N_2711,N_2655);
or UO_2 (O_2,N_2945,N_2955);
nor UO_3 (O_3,N_2685,N_2533);
nor UO_4 (O_4,N_2650,N_2770);
and UO_5 (O_5,N_2731,N_2769);
nor UO_6 (O_6,N_2557,N_2712);
nand UO_7 (O_7,N_2700,N_2708);
nor UO_8 (O_8,N_2473,N_2490);
or UO_9 (O_9,N_2461,N_2483);
nor UO_10 (O_10,N_2824,N_2995);
nor UO_11 (O_11,N_2682,N_2753);
and UO_12 (O_12,N_2836,N_2807);
nand UO_13 (O_13,N_2965,N_2773);
nand UO_14 (O_14,N_2625,N_2605);
nand UO_15 (O_15,N_2998,N_2725);
or UO_16 (O_16,N_2783,N_2428);
xnor UO_17 (O_17,N_2762,N_2893);
or UO_18 (O_18,N_2832,N_2950);
and UO_19 (O_19,N_2932,N_2814);
or UO_20 (O_20,N_2687,N_2829);
and UO_21 (O_21,N_2432,N_2589);
and UO_22 (O_22,N_2787,N_2583);
or UO_23 (O_23,N_2610,N_2582);
and UO_24 (O_24,N_2604,N_2899);
xnor UO_25 (O_25,N_2948,N_2684);
and UO_26 (O_26,N_2830,N_2699);
and UO_27 (O_27,N_2532,N_2407);
nand UO_28 (O_28,N_2840,N_2431);
and UO_29 (O_29,N_2617,N_2594);
and UO_30 (O_30,N_2569,N_2596);
and UO_31 (O_31,N_2906,N_2908);
nand UO_32 (O_32,N_2846,N_2881);
or UO_33 (O_33,N_2624,N_2941);
or UO_34 (O_34,N_2933,N_2651);
nor UO_35 (O_35,N_2668,N_2622);
nand UO_36 (O_36,N_2534,N_2877);
nor UO_37 (O_37,N_2737,N_2630);
or UO_38 (O_38,N_2554,N_2518);
or UO_39 (O_39,N_2789,N_2522);
nor UO_40 (O_40,N_2648,N_2584);
and UO_41 (O_41,N_2992,N_2747);
or UO_42 (O_42,N_2957,N_2450);
and UO_43 (O_43,N_2987,N_2419);
and UO_44 (O_44,N_2646,N_2619);
nor UO_45 (O_45,N_2511,N_2784);
or UO_46 (O_46,N_2776,N_2879);
nand UO_47 (O_47,N_2601,N_2459);
and UO_48 (O_48,N_2714,N_2756);
or UO_49 (O_49,N_2615,N_2577);
nor UO_50 (O_50,N_2822,N_2867);
nor UO_51 (O_51,N_2971,N_2930);
or UO_52 (O_52,N_2695,N_2482);
and UO_53 (O_53,N_2856,N_2400);
and UO_54 (O_54,N_2420,N_2425);
nor UO_55 (O_55,N_2692,N_2732);
and UO_56 (O_56,N_2905,N_2471);
nand UO_57 (O_57,N_2705,N_2723);
and UO_58 (O_58,N_2664,N_2813);
nor UO_59 (O_59,N_2942,N_2408);
or UO_60 (O_60,N_2728,N_2478);
or UO_61 (O_61,N_2984,N_2456);
and UO_62 (O_62,N_2865,N_2764);
and UO_63 (O_63,N_2854,N_2567);
or UO_64 (O_64,N_2669,N_2496);
nor UO_65 (O_65,N_2959,N_2652);
nand UO_66 (O_66,N_2703,N_2544);
or UO_67 (O_67,N_2542,N_2477);
and UO_68 (O_68,N_2620,N_2936);
nor UO_69 (O_69,N_2973,N_2526);
and UO_70 (O_70,N_2489,N_2458);
nor UO_71 (O_71,N_2633,N_2454);
nor UO_72 (O_72,N_2676,N_2778);
and UO_73 (O_73,N_2882,N_2863);
or UO_74 (O_74,N_2686,N_2562);
or UO_75 (O_75,N_2427,N_2581);
or UO_76 (O_76,N_2476,N_2535);
nor UO_77 (O_77,N_2979,N_2525);
nand UO_78 (O_78,N_2497,N_2403);
and UO_79 (O_79,N_2913,N_2969);
nand UO_80 (O_80,N_2749,N_2663);
or UO_81 (O_81,N_2976,N_2873);
nand UO_82 (O_82,N_2411,N_2565);
nor UO_83 (O_83,N_2637,N_2818);
nor UO_84 (O_84,N_2444,N_2972);
nor UO_85 (O_85,N_2896,N_2795);
nor UO_86 (O_86,N_2548,N_2733);
and UO_87 (O_87,N_2883,N_2493);
nand UO_88 (O_88,N_2429,N_2516);
nor UO_89 (O_89,N_2927,N_2947);
nand UO_90 (O_90,N_2597,N_2667);
and UO_91 (O_91,N_2592,N_2697);
nand UO_92 (O_92,N_2709,N_2885);
nand UO_93 (O_93,N_2740,N_2726);
and UO_94 (O_94,N_2887,N_2587);
nor UO_95 (O_95,N_2819,N_2853);
nand UO_96 (O_96,N_2735,N_2794);
or UO_97 (O_97,N_2745,N_2455);
or UO_98 (O_98,N_2401,N_2501);
or UO_99 (O_99,N_2674,N_2670);
nand UO_100 (O_100,N_2999,N_2568);
and UO_101 (O_101,N_2938,N_2467);
nor UO_102 (O_102,N_2701,N_2926);
nor UO_103 (O_103,N_2835,N_2977);
and UO_104 (O_104,N_2975,N_2734);
nor UO_105 (O_105,N_2507,N_2848);
nand UO_106 (O_106,N_2717,N_2917);
nor UO_107 (O_107,N_2851,N_2842);
nor UO_108 (O_108,N_2491,N_2484);
and UO_109 (O_109,N_2470,N_2884);
nand UO_110 (O_110,N_2962,N_2791);
nor UO_111 (O_111,N_2614,N_2549);
or UO_112 (O_112,N_2989,N_2993);
xnor UO_113 (O_113,N_2693,N_2481);
nand UO_114 (O_114,N_2445,N_2754);
or UO_115 (O_115,N_2460,N_2801);
and UO_116 (O_116,N_2447,N_2591);
nor UO_117 (O_117,N_2677,N_2869);
or UO_118 (O_118,N_2698,N_2657);
and UO_119 (O_119,N_2994,N_2763);
nand UO_120 (O_120,N_2876,N_2616);
or UO_121 (O_121,N_2436,N_2742);
or UO_122 (O_122,N_2985,N_2416);
nor UO_123 (O_123,N_2804,N_2574);
nor UO_124 (O_124,N_2662,N_2585);
nor UO_125 (O_125,N_2864,N_2815);
and UO_126 (O_126,N_2966,N_2744);
or UO_127 (O_127,N_2833,N_2766);
and UO_128 (O_128,N_2440,N_2452);
nor UO_129 (O_129,N_2739,N_2555);
and UO_130 (O_130,N_2462,N_2943);
and UO_131 (O_131,N_2844,N_2406);
nor UO_132 (O_132,N_2914,N_2506);
nand UO_133 (O_133,N_2817,N_2426);
and UO_134 (O_134,N_2576,N_2857);
or UO_135 (O_135,N_2860,N_2551);
or UO_136 (O_136,N_2607,N_2593);
or UO_137 (O_137,N_2472,N_2826);
or UO_138 (O_138,N_2422,N_2777);
or UO_139 (O_139,N_2654,N_2465);
or UO_140 (O_140,N_2681,N_2874);
nand UO_141 (O_141,N_2892,N_2730);
or UO_142 (O_142,N_2797,N_2839);
nor UO_143 (O_143,N_2485,N_2451);
nor UO_144 (O_144,N_2515,N_2897);
or UO_145 (O_145,N_2768,N_2528);
nand UO_146 (O_146,N_2858,N_2508);
nand UO_147 (O_147,N_2788,N_2982);
nor UO_148 (O_148,N_2751,N_2954);
or UO_149 (O_149,N_2771,N_2598);
or UO_150 (O_150,N_2931,N_2752);
or UO_151 (O_151,N_2631,N_2678);
or UO_152 (O_152,N_2722,N_2871);
nand UO_153 (O_153,N_2602,N_2890);
nand UO_154 (O_154,N_2643,N_2635);
nor UO_155 (O_155,N_2675,N_2916);
or UO_156 (O_156,N_2823,N_2718);
or UO_157 (O_157,N_2634,N_2628);
nor UO_158 (O_158,N_2924,N_2870);
or UO_159 (O_159,N_2793,N_2514);
xnor UO_160 (O_160,N_2872,N_2702);
and UO_161 (O_161,N_2691,N_2792);
and UO_162 (O_162,N_2939,N_2561);
nor UO_163 (O_163,N_2658,N_2688);
or UO_164 (O_164,N_2967,N_2573);
nor UO_165 (O_165,N_2828,N_2530);
or UO_166 (O_166,N_2547,N_2413);
nor UO_167 (O_167,N_2757,N_2843);
nor UO_168 (O_168,N_2782,N_2618);
and UO_169 (O_169,N_2434,N_2433);
and UO_170 (O_170,N_2921,N_2812);
nor UO_171 (O_171,N_2475,N_2850);
nand UO_172 (O_172,N_2940,N_2510);
nor UO_173 (O_173,N_2636,N_2901);
nand UO_174 (O_174,N_2755,N_2517);
xnor UO_175 (O_175,N_2531,N_2759);
nand UO_176 (O_176,N_2661,N_2767);
and UO_177 (O_177,N_2743,N_2430);
or UO_178 (O_178,N_2609,N_2861);
nor UO_179 (O_179,N_2494,N_2642);
nor UO_180 (O_180,N_2834,N_2539);
and UO_181 (O_181,N_2512,N_2588);
or UO_182 (O_182,N_2612,N_2919);
and UO_183 (O_183,N_2796,N_2781);
nor UO_184 (O_184,N_2603,N_2779);
nor UO_185 (O_185,N_2802,N_2423);
nor UO_186 (O_186,N_2640,N_2521);
and UO_187 (O_187,N_2509,N_2847);
xor UO_188 (O_188,N_2719,N_2556);
or UO_189 (O_189,N_2785,N_2627);
or UO_190 (O_190,N_2920,N_2715);
or UO_191 (O_191,N_2629,N_2412);
or UO_192 (O_192,N_2894,N_2438);
nor UO_193 (O_193,N_2727,N_2964);
nand UO_194 (O_194,N_2448,N_2953);
nand UO_195 (O_195,N_2404,N_2666);
nand UO_196 (O_196,N_2520,N_2566);
and UO_197 (O_197,N_2457,N_2845);
nor UO_198 (O_198,N_2922,N_2799);
or UO_199 (O_199,N_2586,N_2523);
and UO_200 (O_200,N_2418,N_2513);
nand UO_201 (O_201,N_2750,N_2621);
and UO_202 (O_202,N_2632,N_2495);
nor UO_203 (O_203,N_2469,N_2487);
nor UO_204 (O_204,N_2645,N_2679);
or UO_205 (O_205,N_2623,N_2519);
nor UO_206 (O_206,N_2935,N_2696);
nor UO_207 (O_207,N_2409,N_2421);
nor UO_208 (O_208,N_2827,N_2417);
nor UO_209 (O_209,N_2990,N_2553);
or UO_210 (O_210,N_2649,N_2564);
nand UO_211 (O_211,N_2820,N_2500);
nand UO_212 (O_212,N_2590,N_2852);
or UO_213 (O_213,N_2552,N_2704);
and UO_214 (O_214,N_2720,N_2660);
nand UO_215 (O_215,N_2886,N_2758);
or UO_216 (O_216,N_2595,N_2925);
and UO_217 (O_217,N_2572,N_2952);
nor UO_218 (O_218,N_2672,N_2505);
and UO_219 (O_219,N_2798,N_2504);
nor UO_220 (O_220,N_2963,N_2446);
and UO_221 (O_221,N_2915,N_2806);
and UO_222 (O_222,N_2659,N_2683);
or UO_223 (O_223,N_2541,N_2875);
or UO_224 (O_224,N_2831,N_2912);
nand UO_225 (O_225,N_2443,N_2849);
or UO_226 (O_226,N_2499,N_2644);
and UO_227 (O_227,N_2599,N_2880);
and UO_228 (O_228,N_2414,N_2479);
nand UO_229 (O_229,N_2790,N_2974);
nor UO_230 (O_230,N_2464,N_2761);
nand UO_231 (O_231,N_2997,N_2575);
nor UO_232 (O_232,N_2956,N_2838);
nand UO_233 (O_233,N_2944,N_2558);
or UO_234 (O_234,N_2606,N_2641);
nor UO_235 (O_235,N_2811,N_2608);
and UO_236 (O_236,N_2748,N_2862);
or UO_237 (O_237,N_2825,N_2690);
or UO_238 (O_238,N_2980,N_2809);
nor UO_239 (O_239,N_2611,N_2673);
and UO_240 (O_240,N_2405,N_2498);
or UO_241 (O_241,N_2441,N_2437);
nor UO_242 (O_242,N_2909,N_2888);
nand UO_243 (O_243,N_2978,N_2529);
or UO_244 (O_244,N_2653,N_2415);
and UO_245 (O_245,N_2468,N_2868);
or UO_246 (O_246,N_2803,N_2929);
nand UO_247 (O_247,N_2424,N_2579);
nor UO_248 (O_248,N_2895,N_2902);
nand UO_249 (O_249,N_2524,N_2600);
nor UO_250 (O_250,N_2918,N_2527);
or UO_251 (O_251,N_2910,N_2639);
or UO_252 (O_252,N_2951,N_2536);
nand UO_253 (O_253,N_2904,N_2808);
nand UO_254 (O_254,N_2563,N_2503);
nand UO_255 (O_255,N_2671,N_2866);
nand UO_256 (O_256,N_2746,N_2638);
nor UO_257 (O_257,N_2923,N_2435);
and UO_258 (O_258,N_2800,N_2410);
nand UO_259 (O_259,N_2837,N_2760);
nand UO_260 (O_260,N_2466,N_2738);
and UO_261 (O_261,N_2694,N_2492);
and UO_262 (O_262,N_2928,N_2889);
and UO_263 (O_263,N_2996,N_2713);
nand UO_264 (O_264,N_2772,N_2724);
nand UO_265 (O_265,N_2934,N_2786);
nor UO_266 (O_266,N_2970,N_2710);
or UO_267 (O_267,N_2937,N_2545);
nor UO_268 (O_268,N_2480,N_2946);
nor UO_269 (O_269,N_2729,N_2463);
nor UO_270 (O_270,N_2960,N_2780);
or UO_271 (O_271,N_2775,N_2988);
nand UO_272 (O_272,N_2841,N_2449);
and UO_273 (O_273,N_2736,N_2859);
nand UO_274 (O_274,N_2765,N_2816);
nand UO_275 (O_275,N_2810,N_2550);
and UO_276 (O_276,N_2898,N_2907);
or UO_277 (O_277,N_2706,N_2647);
or UO_278 (O_278,N_2900,N_2486);
and UO_279 (O_279,N_2453,N_2891);
nor UO_280 (O_280,N_2689,N_2991);
nor UO_281 (O_281,N_2774,N_2981);
or UO_282 (O_282,N_2903,N_2571);
nand UO_283 (O_283,N_2958,N_2968);
nor UO_284 (O_284,N_2741,N_2721);
or UO_285 (O_285,N_2474,N_2540);
or UO_286 (O_286,N_2911,N_2656);
nor UO_287 (O_287,N_2613,N_2560);
and UO_288 (O_288,N_2546,N_2502);
nand UO_289 (O_289,N_2442,N_2961);
or UO_290 (O_290,N_2949,N_2986);
and UO_291 (O_291,N_2878,N_2439);
nor UO_292 (O_292,N_2543,N_2680);
or UO_293 (O_293,N_2707,N_2578);
nand UO_294 (O_294,N_2570,N_2537);
nand UO_295 (O_295,N_2983,N_2805);
or UO_296 (O_296,N_2665,N_2402);
nor UO_297 (O_297,N_2821,N_2538);
and UO_298 (O_298,N_2716,N_2855);
or UO_299 (O_299,N_2488,N_2580);
nor UO_300 (O_300,N_2751,N_2784);
and UO_301 (O_301,N_2638,N_2612);
or UO_302 (O_302,N_2806,N_2637);
and UO_303 (O_303,N_2473,N_2591);
or UO_304 (O_304,N_2573,N_2953);
nand UO_305 (O_305,N_2778,N_2449);
nand UO_306 (O_306,N_2457,N_2501);
nand UO_307 (O_307,N_2793,N_2559);
or UO_308 (O_308,N_2709,N_2418);
nor UO_309 (O_309,N_2886,N_2899);
nor UO_310 (O_310,N_2441,N_2719);
nor UO_311 (O_311,N_2568,N_2818);
nor UO_312 (O_312,N_2719,N_2579);
nor UO_313 (O_313,N_2858,N_2995);
or UO_314 (O_314,N_2896,N_2742);
or UO_315 (O_315,N_2519,N_2647);
and UO_316 (O_316,N_2906,N_2728);
or UO_317 (O_317,N_2732,N_2538);
and UO_318 (O_318,N_2872,N_2723);
and UO_319 (O_319,N_2788,N_2821);
and UO_320 (O_320,N_2754,N_2400);
nor UO_321 (O_321,N_2406,N_2420);
or UO_322 (O_322,N_2409,N_2762);
nand UO_323 (O_323,N_2494,N_2540);
and UO_324 (O_324,N_2992,N_2986);
and UO_325 (O_325,N_2423,N_2892);
or UO_326 (O_326,N_2701,N_2633);
or UO_327 (O_327,N_2697,N_2510);
nor UO_328 (O_328,N_2516,N_2657);
nand UO_329 (O_329,N_2948,N_2765);
nor UO_330 (O_330,N_2798,N_2873);
nor UO_331 (O_331,N_2570,N_2978);
nand UO_332 (O_332,N_2933,N_2697);
nor UO_333 (O_333,N_2771,N_2745);
and UO_334 (O_334,N_2732,N_2669);
or UO_335 (O_335,N_2658,N_2689);
and UO_336 (O_336,N_2492,N_2610);
nand UO_337 (O_337,N_2926,N_2449);
and UO_338 (O_338,N_2753,N_2843);
or UO_339 (O_339,N_2617,N_2752);
nand UO_340 (O_340,N_2504,N_2529);
or UO_341 (O_341,N_2730,N_2415);
nand UO_342 (O_342,N_2500,N_2599);
nor UO_343 (O_343,N_2691,N_2719);
or UO_344 (O_344,N_2816,N_2587);
nand UO_345 (O_345,N_2840,N_2438);
or UO_346 (O_346,N_2461,N_2567);
nand UO_347 (O_347,N_2976,N_2923);
and UO_348 (O_348,N_2746,N_2577);
nor UO_349 (O_349,N_2791,N_2724);
or UO_350 (O_350,N_2920,N_2682);
nand UO_351 (O_351,N_2983,N_2890);
nor UO_352 (O_352,N_2489,N_2940);
or UO_353 (O_353,N_2469,N_2523);
nand UO_354 (O_354,N_2591,N_2874);
nor UO_355 (O_355,N_2993,N_2413);
and UO_356 (O_356,N_2624,N_2499);
nor UO_357 (O_357,N_2931,N_2814);
or UO_358 (O_358,N_2856,N_2629);
and UO_359 (O_359,N_2636,N_2742);
nand UO_360 (O_360,N_2845,N_2754);
nand UO_361 (O_361,N_2974,N_2892);
and UO_362 (O_362,N_2785,N_2461);
nand UO_363 (O_363,N_2880,N_2598);
nand UO_364 (O_364,N_2621,N_2966);
nor UO_365 (O_365,N_2892,N_2445);
or UO_366 (O_366,N_2801,N_2453);
nand UO_367 (O_367,N_2565,N_2513);
and UO_368 (O_368,N_2794,N_2725);
or UO_369 (O_369,N_2451,N_2943);
or UO_370 (O_370,N_2425,N_2414);
or UO_371 (O_371,N_2742,N_2778);
and UO_372 (O_372,N_2527,N_2827);
and UO_373 (O_373,N_2990,N_2816);
or UO_374 (O_374,N_2729,N_2652);
or UO_375 (O_375,N_2435,N_2780);
nand UO_376 (O_376,N_2968,N_2536);
nand UO_377 (O_377,N_2449,N_2500);
and UO_378 (O_378,N_2797,N_2822);
nor UO_379 (O_379,N_2910,N_2983);
nand UO_380 (O_380,N_2492,N_2449);
or UO_381 (O_381,N_2456,N_2963);
nand UO_382 (O_382,N_2695,N_2736);
or UO_383 (O_383,N_2949,N_2862);
nand UO_384 (O_384,N_2837,N_2973);
or UO_385 (O_385,N_2555,N_2993);
nand UO_386 (O_386,N_2658,N_2615);
nor UO_387 (O_387,N_2508,N_2807);
nor UO_388 (O_388,N_2995,N_2770);
and UO_389 (O_389,N_2486,N_2557);
and UO_390 (O_390,N_2428,N_2676);
or UO_391 (O_391,N_2838,N_2518);
nand UO_392 (O_392,N_2632,N_2928);
nand UO_393 (O_393,N_2581,N_2446);
nor UO_394 (O_394,N_2921,N_2668);
or UO_395 (O_395,N_2523,N_2815);
nor UO_396 (O_396,N_2511,N_2547);
nand UO_397 (O_397,N_2877,N_2505);
nor UO_398 (O_398,N_2505,N_2736);
nor UO_399 (O_399,N_2684,N_2818);
or UO_400 (O_400,N_2846,N_2835);
or UO_401 (O_401,N_2409,N_2674);
nand UO_402 (O_402,N_2610,N_2457);
and UO_403 (O_403,N_2780,N_2948);
xor UO_404 (O_404,N_2885,N_2748);
and UO_405 (O_405,N_2665,N_2534);
nand UO_406 (O_406,N_2511,N_2839);
and UO_407 (O_407,N_2768,N_2929);
and UO_408 (O_408,N_2951,N_2420);
or UO_409 (O_409,N_2405,N_2419);
and UO_410 (O_410,N_2480,N_2938);
nand UO_411 (O_411,N_2814,N_2641);
nor UO_412 (O_412,N_2937,N_2980);
nor UO_413 (O_413,N_2467,N_2844);
or UO_414 (O_414,N_2700,N_2677);
nand UO_415 (O_415,N_2951,N_2878);
or UO_416 (O_416,N_2877,N_2783);
and UO_417 (O_417,N_2796,N_2477);
nand UO_418 (O_418,N_2913,N_2884);
or UO_419 (O_419,N_2637,N_2657);
nor UO_420 (O_420,N_2935,N_2679);
and UO_421 (O_421,N_2678,N_2912);
nand UO_422 (O_422,N_2545,N_2732);
or UO_423 (O_423,N_2946,N_2526);
and UO_424 (O_424,N_2874,N_2764);
xnor UO_425 (O_425,N_2472,N_2425);
and UO_426 (O_426,N_2871,N_2864);
and UO_427 (O_427,N_2881,N_2442);
or UO_428 (O_428,N_2594,N_2472);
nand UO_429 (O_429,N_2812,N_2920);
nor UO_430 (O_430,N_2651,N_2928);
or UO_431 (O_431,N_2628,N_2846);
nand UO_432 (O_432,N_2733,N_2757);
and UO_433 (O_433,N_2972,N_2936);
or UO_434 (O_434,N_2649,N_2422);
nor UO_435 (O_435,N_2512,N_2805);
nand UO_436 (O_436,N_2700,N_2647);
or UO_437 (O_437,N_2675,N_2776);
or UO_438 (O_438,N_2666,N_2454);
and UO_439 (O_439,N_2560,N_2734);
or UO_440 (O_440,N_2464,N_2946);
nand UO_441 (O_441,N_2930,N_2571);
or UO_442 (O_442,N_2453,N_2938);
and UO_443 (O_443,N_2623,N_2995);
or UO_444 (O_444,N_2415,N_2686);
nand UO_445 (O_445,N_2819,N_2471);
nor UO_446 (O_446,N_2699,N_2931);
nand UO_447 (O_447,N_2921,N_2560);
nor UO_448 (O_448,N_2807,N_2933);
or UO_449 (O_449,N_2715,N_2623);
and UO_450 (O_450,N_2755,N_2461);
or UO_451 (O_451,N_2627,N_2554);
nor UO_452 (O_452,N_2985,N_2710);
or UO_453 (O_453,N_2453,N_2570);
nor UO_454 (O_454,N_2961,N_2714);
or UO_455 (O_455,N_2955,N_2929);
nor UO_456 (O_456,N_2442,N_2536);
or UO_457 (O_457,N_2825,N_2785);
nand UO_458 (O_458,N_2642,N_2976);
nor UO_459 (O_459,N_2759,N_2895);
nand UO_460 (O_460,N_2748,N_2402);
and UO_461 (O_461,N_2689,N_2820);
nand UO_462 (O_462,N_2627,N_2620);
or UO_463 (O_463,N_2600,N_2658);
and UO_464 (O_464,N_2686,N_2708);
nor UO_465 (O_465,N_2995,N_2639);
nand UO_466 (O_466,N_2510,N_2840);
nor UO_467 (O_467,N_2667,N_2699);
nor UO_468 (O_468,N_2879,N_2796);
nor UO_469 (O_469,N_2425,N_2906);
nor UO_470 (O_470,N_2450,N_2833);
nor UO_471 (O_471,N_2895,N_2472);
nor UO_472 (O_472,N_2700,N_2535);
or UO_473 (O_473,N_2544,N_2453);
or UO_474 (O_474,N_2958,N_2818);
nand UO_475 (O_475,N_2768,N_2976);
nand UO_476 (O_476,N_2591,N_2822);
and UO_477 (O_477,N_2826,N_2873);
nand UO_478 (O_478,N_2768,N_2444);
and UO_479 (O_479,N_2866,N_2812);
and UO_480 (O_480,N_2718,N_2998);
nor UO_481 (O_481,N_2806,N_2722);
and UO_482 (O_482,N_2796,N_2583);
and UO_483 (O_483,N_2740,N_2978);
and UO_484 (O_484,N_2902,N_2736);
or UO_485 (O_485,N_2510,N_2516);
nor UO_486 (O_486,N_2891,N_2696);
and UO_487 (O_487,N_2441,N_2447);
nor UO_488 (O_488,N_2965,N_2967);
or UO_489 (O_489,N_2918,N_2494);
or UO_490 (O_490,N_2856,N_2476);
nor UO_491 (O_491,N_2790,N_2628);
and UO_492 (O_492,N_2494,N_2948);
and UO_493 (O_493,N_2847,N_2973);
and UO_494 (O_494,N_2518,N_2768);
or UO_495 (O_495,N_2490,N_2914);
nor UO_496 (O_496,N_2757,N_2675);
and UO_497 (O_497,N_2722,N_2528);
and UO_498 (O_498,N_2484,N_2983);
or UO_499 (O_499,N_2979,N_2575);
endmodule