module basic_500_3000_500_4_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xor U0 (N_0,In_146,In_479);
or U1 (N_1,In_444,In_30);
nand U2 (N_2,In_74,In_142);
nand U3 (N_3,In_9,In_160);
and U4 (N_4,In_254,In_398);
xor U5 (N_5,In_393,In_497);
nor U6 (N_6,In_239,In_166);
and U7 (N_7,In_240,In_199);
xnor U8 (N_8,In_456,In_144);
nand U9 (N_9,In_169,In_449);
nor U10 (N_10,In_349,In_491);
or U11 (N_11,In_457,In_27);
xor U12 (N_12,In_106,In_492);
xnor U13 (N_13,In_45,In_185);
nand U14 (N_14,In_280,In_462);
nor U15 (N_15,In_277,In_348);
or U16 (N_16,In_435,In_136);
nor U17 (N_17,In_147,In_253);
nand U18 (N_18,In_149,In_412);
xor U19 (N_19,In_214,In_172);
xor U20 (N_20,In_145,In_422);
or U21 (N_21,In_250,In_126);
nand U22 (N_22,In_18,In_208);
or U23 (N_23,In_51,In_347);
nand U24 (N_24,In_446,In_68);
xnor U25 (N_25,In_490,In_419);
nor U26 (N_26,In_105,In_235);
and U27 (N_27,In_252,In_210);
and U28 (N_28,In_247,In_223);
and U29 (N_29,In_372,In_191);
nor U30 (N_30,In_82,In_120);
nor U31 (N_31,In_148,In_287);
or U32 (N_32,In_324,In_282);
xor U33 (N_33,In_284,In_478);
nor U34 (N_34,In_440,In_111);
nor U35 (N_35,In_487,In_383);
and U36 (N_36,In_98,In_171);
and U37 (N_37,In_63,In_392);
nand U38 (N_38,In_156,In_413);
or U39 (N_39,In_218,In_415);
nand U40 (N_40,In_410,In_110);
and U41 (N_41,In_202,In_139);
nand U42 (N_42,In_228,In_87);
nor U43 (N_43,In_367,In_450);
and U44 (N_44,In_49,In_436);
nand U45 (N_45,In_134,In_445);
and U46 (N_46,In_396,In_453);
and U47 (N_47,In_22,In_288);
or U48 (N_48,In_438,In_267);
nand U49 (N_49,In_231,In_67);
nor U50 (N_50,In_353,In_431);
nor U51 (N_51,In_154,In_269);
or U52 (N_52,In_59,In_115);
xor U53 (N_53,In_471,In_296);
nand U54 (N_54,In_245,In_265);
xor U55 (N_55,In_97,In_314);
and U56 (N_56,In_81,In_366);
xnor U57 (N_57,In_326,In_317);
or U58 (N_58,In_60,In_163);
or U59 (N_59,In_137,In_88);
nor U60 (N_60,In_211,In_132);
or U61 (N_61,In_236,In_325);
and U62 (N_62,In_200,In_42);
nor U63 (N_63,In_331,In_403);
and U64 (N_64,In_109,In_258);
nor U65 (N_65,In_44,In_174);
or U66 (N_66,In_429,In_365);
or U67 (N_67,In_151,In_266);
xor U68 (N_68,In_433,In_370);
xor U69 (N_69,In_345,In_143);
and U70 (N_70,In_322,In_53);
xor U71 (N_71,In_489,In_48);
or U72 (N_72,In_119,In_128);
xor U73 (N_73,In_307,In_448);
and U74 (N_74,In_346,In_56);
and U75 (N_75,In_337,In_298);
and U76 (N_76,In_104,In_170);
xor U77 (N_77,In_424,In_55);
xnor U78 (N_78,In_188,In_304);
nand U79 (N_79,In_246,In_83);
nor U80 (N_80,In_310,In_274);
or U81 (N_81,In_472,In_73);
or U82 (N_82,In_182,In_350);
and U83 (N_83,In_31,In_230);
or U84 (N_84,In_96,In_224);
nand U85 (N_85,In_173,In_375);
nor U86 (N_86,In_447,In_164);
xor U87 (N_87,In_434,In_452);
nor U88 (N_88,In_90,In_72);
nand U89 (N_89,In_293,In_432);
and U90 (N_90,In_339,In_305);
and U91 (N_91,In_464,In_0);
and U92 (N_92,In_256,In_77);
and U93 (N_93,In_10,In_28);
nor U94 (N_94,In_481,In_54);
nor U95 (N_95,In_232,In_391);
or U96 (N_96,In_292,In_11);
or U97 (N_97,In_175,In_99);
and U98 (N_98,In_333,In_43);
nor U99 (N_99,In_37,In_207);
nand U100 (N_100,In_385,In_6);
xor U101 (N_101,In_152,In_36);
xnor U102 (N_102,In_319,In_332);
xor U103 (N_103,In_338,In_386);
and U104 (N_104,In_13,In_276);
xnor U105 (N_105,In_342,In_183);
and U106 (N_106,In_47,In_114);
or U107 (N_107,In_430,In_219);
or U108 (N_108,In_356,In_21);
or U109 (N_109,In_470,In_93);
nor U110 (N_110,In_113,In_485);
or U111 (N_111,In_401,In_2);
nand U112 (N_112,In_255,In_368);
nand U113 (N_113,In_417,In_29);
xnor U114 (N_114,In_272,In_124);
nand U115 (N_115,In_177,In_389);
nand U116 (N_116,In_343,In_468);
or U117 (N_117,In_474,In_290);
and U118 (N_118,In_150,In_25);
and U119 (N_119,In_493,In_397);
nor U120 (N_120,In_420,In_108);
nor U121 (N_121,In_461,In_50);
nand U122 (N_122,In_388,In_390);
and U123 (N_123,In_34,In_380);
or U124 (N_124,In_123,In_103);
xnor U125 (N_125,In_416,In_369);
nand U126 (N_126,In_117,In_414);
xor U127 (N_127,In_19,In_165);
xnor U128 (N_128,In_190,In_138);
xor U129 (N_129,In_264,In_498);
nand U130 (N_130,In_130,In_141);
or U131 (N_131,In_459,In_285);
nand U132 (N_132,In_61,In_455);
nor U133 (N_133,In_294,In_358);
or U134 (N_134,In_312,In_14);
xnor U135 (N_135,In_38,In_91);
or U136 (N_136,In_354,In_283);
or U137 (N_137,In_32,In_313);
or U138 (N_138,In_352,In_162);
xnor U139 (N_139,In_494,In_168);
and U140 (N_140,In_249,In_155);
nor U141 (N_141,In_355,In_281);
xor U142 (N_142,In_220,In_39);
nor U143 (N_143,In_480,In_122);
or U144 (N_144,In_242,In_483);
nand U145 (N_145,In_241,In_351);
nand U146 (N_146,In_308,In_127);
xor U147 (N_147,In_167,In_159);
or U148 (N_148,In_306,In_24);
or U149 (N_149,In_65,In_300);
or U150 (N_150,In_262,In_7);
and U151 (N_151,In_411,In_437);
nand U152 (N_152,In_309,In_179);
and U153 (N_153,In_5,In_484);
or U154 (N_154,In_248,In_35);
and U155 (N_155,In_94,In_395);
nand U156 (N_156,In_263,In_71);
or U157 (N_157,In_216,In_328);
nor U158 (N_158,In_79,In_102);
xor U159 (N_159,In_64,In_374);
and U160 (N_160,In_463,In_244);
nor U161 (N_161,In_311,In_299);
and U162 (N_162,In_344,In_291);
or U163 (N_163,In_460,In_466);
xnor U164 (N_164,In_95,In_261);
and U165 (N_165,In_157,In_204);
xnor U166 (N_166,In_381,In_251);
nor U167 (N_167,In_499,In_180);
xnor U168 (N_168,In_441,In_186);
xor U169 (N_169,In_423,In_271);
and U170 (N_170,In_407,In_315);
nor U171 (N_171,In_62,In_4);
xnor U172 (N_172,In_221,In_476);
or U173 (N_173,In_229,In_327);
nand U174 (N_174,In_486,In_357);
nor U175 (N_175,In_70,In_107);
xor U176 (N_176,In_330,In_329);
xnor U177 (N_177,In_86,In_406);
nand U178 (N_178,In_451,In_217);
or U179 (N_179,In_268,In_206);
nor U180 (N_180,In_212,In_57);
or U181 (N_181,In_213,In_33);
nor U182 (N_182,In_379,In_259);
xor U183 (N_183,In_289,In_238);
nand U184 (N_184,In_84,In_16);
nand U185 (N_185,In_477,In_243);
nor U186 (N_186,In_376,In_408);
nor U187 (N_187,In_402,In_442);
nand U188 (N_188,In_153,In_428);
and U189 (N_189,In_40,In_469);
nand U190 (N_190,In_184,In_360);
xor U191 (N_191,In_302,In_76);
and U192 (N_192,In_359,In_394);
and U193 (N_193,In_125,In_335);
nor U194 (N_194,In_400,In_270);
nand U195 (N_195,In_197,In_80);
and U196 (N_196,In_205,In_334);
nor U197 (N_197,In_189,In_278);
and U198 (N_198,In_58,In_286);
xor U199 (N_199,In_439,In_473);
nor U200 (N_200,In_46,In_66);
nor U201 (N_201,In_467,In_233);
nor U202 (N_202,In_297,In_321);
and U203 (N_203,In_52,In_362);
xor U204 (N_204,In_373,In_260);
or U205 (N_205,In_303,In_192);
and U206 (N_206,In_195,In_273);
xnor U207 (N_207,In_418,In_496);
xor U208 (N_208,In_133,In_215);
nand U209 (N_209,In_101,In_404);
and U210 (N_210,In_1,In_301);
and U211 (N_211,In_237,In_194);
nor U212 (N_212,In_458,In_140);
nand U213 (N_213,In_198,In_118);
or U214 (N_214,In_340,In_279);
and U215 (N_215,In_409,In_378);
and U216 (N_216,In_361,In_12);
or U217 (N_217,In_475,In_26);
or U218 (N_218,In_129,In_465);
xnor U219 (N_219,In_116,In_161);
or U220 (N_220,In_69,In_295);
nor U221 (N_221,In_181,In_193);
nor U222 (N_222,In_158,In_92);
nor U223 (N_223,In_425,In_427);
and U224 (N_224,In_178,In_41);
xnor U225 (N_225,In_454,In_363);
xor U226 (N_226,In_488,In_341);
and U227 (N_227,In_8,In_364);
nor U228 (N_228,In_275,In_17);
xor U229 (N_229,In_482,In_382);
nor U230 (N_230,In_196,In_85);
nand U231 (N_231,In_426,In_227);
nand U232 (N_232,In_226,In_135);
nand U233 (N_233,In_15,In_100);
xor U234 (N_234,In_3,In_203);
or U235 (N_235,In_20,In_23);
nand U236 (N_236,In_320,In_443);
and U237 (N_237,In_222,In_377);
xnor U238 (N_238,In_75,In_318);
nor U239 (N_239,In_405,In_176);
xor U240 (N_240,In_316,In_336);
or U241 (N_241,In_209,In_225);
and U242 (N_242,In_257,In_495);
xnor U243 (N_243,In_234,In_187);
xnor U244 (N_244,In_131,In_371);
xnor U245 (N_245,In_201,In_121);
xor U246 (N_246,In_421,In_323);
nand U247 (N_247,In_78,In_387);
xnor U248 (N_248,In_384,In_112);
or U249 (N_249,In_89,In_399);
and U250 (N_250,In_488,In_151);
and U251 (N_251,In_386,In_333);
and U252 (N_252,In_360,In_320);
nor U253 (N_253,In_404,In_281);
and U254 (N_254,In_359,In_269);
xnor U255 (N_255,In_270,In_357);
nor U256 (N_256,In_327,In_79);
and U257 (N_257,In_31,In_120);
nor U258 (N_258,In_407,In_144);
nor U259 (N_259,In_450,In_79);
and U260 (N_260,In_266,In_70);
and U261 (N_261,In_199,In_89);
and U262 (N_262,In_441,In_412);
nand U263 (N_263,In_172,In_6);
and U264 (N_264,In_242,In_310);
nor U265 (N_265,In_302,In_443);
nor U266 (N_266,In_480,In_149);
nand U267 (N_267,In_408,In_33);
xnor U268 (N_268,In_166,In_200);
or U269 (N_269,In_178,In_285);
xnor U270 (N_270,In_459,In_181);
nand U271 (N_271,In_168,In_170);
or U272 (N_272,In_422,In_485);
nand U273 (N_273,In_350,In_247);
nor U274 (N_274,In_72,In_492);
or U275 (N_275,In_121,In_79);
or U276 (N_276,In_24,In_105);
xor U277 (N_277,In_197,In_199);
or U278 (N_278,In_242,In_225);
and U279 (N_279,In_389,In_211);
xor U280 (N_280,In_112,In_175);
or U281 (N_281,In_419,In_308);
and U282 (N_282,In_459,In_224);
and U283 (N_283,In_141,In_152);
or U284 (N_284,In_275,In_141);
and U285 (N_285,In_412,In_203);
and U286 (N_286,In_484,In_485);
xnor U287 (N_287,In_444,In_224);
xnor U288 (N_288,In_208,In_260);
xnor U289 (N_289,In_86,In_11);
and U290 (N_290,In_265,In_424);
and U291 (N_291,In_440,In_315);
and U292 (N_292,In_145,In_418);
nor U293 (N_293,In_319,In_375);
and U294 (N_294,In_310,In_312);
nand U295 (N_295,In_246,In_19);
xor U296 (N_296,In_270,In_332);
or U297 (N_297,In_80,In_417);
nand U298 (N_298,In_183,In_442);
nand U299 (N_299,In_294,In_161);
nand U300 (N_300,In_42,In_225);
or U301 (N_301,In_373,In_43);
xnor U302 (N_302,In_396,In_114);
or U303 (N_303,In_51,In_498);
and U304 (N_304,In_24,In_466);
and U305 (N_305,In_368,In_309);
or U306 (N_306,In_458,In_150);
or U307 (N_307,In_367,In_382);
xnor U308 (N_308,In_88,In_232);
and U309 (N_309,In_219,In_122);
nand U310 (N_310,In_306,In_2);
nand U311 (N_311,In_357,In_412);
nor U312 (N_312,In_196,In_327);
xor U313 (N_313,In_488,In_86);
and U314 (N_314,In_156,In_47);
nor U315 (N_315,In_400,In_402);
and U316 (N_316,In_125,In_162);
or U317 (N_317,In_69,In_196);
or U318 (N_318,In_25,In_16);
nor U319 (N_319,In_448,In_15);
or U320 (N_320,In_404,In_240);
and U321 (N_321,In_151,In_466);
or U322 (N_322,In_51,In_283);
and U323 (N_323,In_239,In_296);
nor U324 (N_324,In_361,In_294);
or U325 (N_325,In_71,In_185);
nor U326 (N_326,In_377,In_40);
or U327 (N_327,In_133,In_38);
nand U328 (N_328,In_81,In_272);
nand U329 (N_329,In_111,In_184);
nand U330 (N_330,In_73,In_230);
nand U331 (N_331,In_214,In_355);
nand U332 (N_332,In_55,In_269);
nor U333 (N_333,In_252,In_396);
or U334 (N_334,In_247,In_406);
and U335 (N_335,In_105,In_118);
xnor U336 (N_336,In_27,In_46);
nand U337 (N_337,In_183,In_340);
or U338 (N_338,In_62,In_168);
and U339 (N_339,In_84,In_173);
nand U340 (N_340,In_477,In_151);
nor U341 (N_341,In_433,In_314);
xor U342 (N_342,In_438,In_365);
nor U343 (N_343,In_383,In_249);
and U344 (N_344,In_75,In_176);
xnor U345 (N_345,In_389,In_411);
or U346 (N_346,In_94,In_217);
and U347 (N_347,In_1,In_181);
nor U348 (N_348,In_451,In_464);
nand U349 (N_349,In_498,In_64);
nor U350 (N_350,In_99,In_338);
xnor U351 (N_351,In_464,In_244);
nor U352 (N_352,In_202,In_484);
nand U353 (N_353,In_285,In_30);
and U354 (N_354,In_156,In_424);
nand U355 (N_355,In_67,In_265);
nand U356 (N_356,In_96,In_215);
nor U357 (N_357,In_448,In_355);
or U358 (N_358,In_407,In_319);
xor U359 (N_359,In_221,In_495);
or U360 (N_360,In_83,In_133);
and U361 (N_361,In_454,In_291);
nand U362 (N_362,In_245,In_258);
nand U363 (N_363,In_397,In_20);
xnor U364 (N_364,In_236,In_470);
nand U365 (N_365,In_152,In_111);
or U366 (N_366,In_449,In_413);
xor U367 (N_367,In_338,In_300);
or U368 (N_368,In_122,In_470);
and U369 (N_369,In_107,In_398);
xnor U370 (N_370,In_498,In_494);
nand U371 (N_371,In_271,In_399);
nor U372 (N_372,In_394,In_49);
xnor U373 (N_373,In_95,In_284);
or U374 (N_374,In_367,In_240);
nand U375 (N_375,In_344,In_72);
or U376 (N_376,In_81,In_227);
xnor U377 (N_377,In_199,In_40);
and U378 (N_378,In_465,In_220);
and U379 (N_379,In_125,In_203);
nor U380 (N_380,In_427,In_370);
nand U381 (N_381,In_399,In_416);
or U382 (N_382,In_240,In_254);
nand U383 (N_383,In_417,In_33);
and U384 (N_384,In_135,In_278);
and U385 (N_385,In_467,In_336);
and U386 (N_386,In_400,In_242);
and U387 (N_387,In_397,In_245);
nand U388 (N_388,In_224,In_355);
nand U389 (N_389,In_99,In_465);
nor U390 (N_390,In_488,In_259);
xnor U391 (N_391,In_328,In_279);
and U392 (N_392,In_50,In_275);
or U393 (N_393,In_141,In_211);
and U394 (N_394,In_489,In_446);
or U395 (N_395,In_447,In_321);
or U396 (N_396,In_83,In_400);
or U397 (N_397,In_315,In_240);
or U398 (N_398,In_486,In_120);
xnor U399 (N_399,In_98,In_380);
nor U400 (N_400,In_113,In_496);
xor U401 (N_401,In_247,In_215);
or U402 (N_402,In_361,In_49);
xnor U403 (N_403,In_456,In_77);
nand U404 (N_404,In_239,In_190);
nand U405 (N_405,In_317,In_65);
nand U406 (N_406,In_482,In_415);
or U407 (N_407,In_101,In_132);
or U408 (N_408,In_208,In_296);
and U409 (N_409,In_171,In_111);
nor U410 (N_410,In_65,In_55);
xnor U411 (N_411,In_261,In_320);
and U412 (N_412,In_33,In_272);
nor U413 (N_413,In_423,In_133);
nor U414 (N_414,In_299,In_437);
and U415 (N_415,In_90,In_443);
and U416 (N_416,In_467,In_279);
and U417 (N_417,In_156,In_295);
nor U418 (N_418,In_39,In_113);
nor U419 (N_419,In_195,In_427);
xnor U420 (N_420,In_271,In_71);
nand U421 (N_421,In_494,In_26);
xor U422 (N_422,In_136,In_89);
and U423 (N_423,In_142,In_254);
nand U424 (N_424,In_88,In_398);
xor U425 (N_425,In_342,In_142);
nand U426 (N_426,In_155,In_367);
and U427 (N_427,In_147,In_226);
xor U428 (N_428,In_337,In_354);
xor U429 (N_429,In_363,In_42);
or U430 (N_430,In_417,In_155);
or U431 (N_431,In_311,In_81);
and U432 (N_432,In_379,In_395);
nand U433 (N_433,In_247,In_487);
nor U434 (N_434,In_343,In_375);
nand U435 (N_435,In_227,In_378);
xnor U436 (N_436,In_395,In_479);
or U437 (N_437,In_79,In_27);
and U438 (N_438,In_203,In_378);
nor U439 (N_439,In_375,In_271);
xor U440 (N_440,In_37,In_370);
and U441 (N_441,In_325,In_481);
or U442 (N_442,In_365,In_238);
or U443 (N_443,In_49,In_232);
xnor U444 (N_444,In_26,In_84);
or U445 (N_445,In_441,In_399);
nand U446 (N_446,In_244,In_84);
xor U447 (N_447,In_495,In_435);
or U448 (N_448,In_359,In_232);
xor U449 (N_449,In_390,In_410);
and U450 (N_450,In_396,In_432);
nand U451 (N_451,In_50,In_264);
nand U452 (N_452,In_208,In_455);
or U453 (N_453,In_415,In_154);
and U454 (N_454,In_60,In_461);
and U455 (N_455,In_186,In_499);
and U456 (N_456,In_10,In_422);
and U457 (N_457,In_399,In_365);
nand U458 (N_458,In_260,In_465);
or U459 (N_459,In_216,In_335);
and U460 (N_460,In_53,In_14);
nor U461 (N_461,In_378,In_349);
xor U462 (N_462,In_54,In_115);
xnor U463 (N_463,In_422,In_169);
and U464 (N_464,In_495,In_465);
and U465 (N_465,In_375,In_51);
and U466 (N_466,In_454,In_436);
nand U467 (N_467,In_44,In_417);
or U468 (N_468,In_303,In_258);
or U469 (N_469,In_294,In_455);
and U470 (N_470,In_312,In_146);
xnor U471 (N_471,In_266,In_475);
nor U472 (N_472,In_45,In_39);
xnor U473 (N_473,In_37,In_2);
nor U474 (N_474,In_62,In_20);
or U475 (N_475,In_421,In_190);
nor U476 (N_476,In_253,In_333);
nand U477 (N_477,In_96,In_188);
and U478 (N_478,In_122,In_316);
and U479 (N_479,In_410,In_405);
nand U480 (N_480,In_396,In_454);
nand U481 (N_481,In_227,In_36);
xor U482 (N_482,In_213,In_186);
nand U483 (N_483,In_408,In_19);
and U484 (N_484,In_18,In_152);
and U485 (N_485,In_5,In_421);
or U486 (N_486,In_287,In_58);
nor U487 (N_487,In_70,In_186);
nor U488 (N_488,In_1,In_473);
xor U489 (N_489,In_463,In_297);
and U490 (N_490,In_325,In_7);
nand U491 (N_491,In_1,In_56);
or U492 (N_492,In_421,In_202);
nor U493 (N_493,In_383,In_12);
or U494 (N_494,In_496,In_179);
or U495 (N_495,In_137,In_198);
and U496 (N_496,In_104,In_478);
and U497 (N_497,In_285,In_130);
xor U498 (N_498,In_289,In_12);
or U499 (N_499,In_187,In_401);
xor U500 (N_500,In_54,In_240);
and U501 (N_501,In_345,In_420);
nand U502 (N_502,In_236,In_294);
and U503 (N_503,In_304,In_62);
nand U504 (N_504,In_20,In_368);
xor U505 (N_505,In_125,In_65);
xnor U506 (N_506,In_138,In_294);
nor U507 (N_507,In_202,In_315);
xnor U508 (N_508,In_9,In_244);
nor U509 (N_509,In_409,In_13);
xor U510 (N_510,In_11,In_131);
or U511 (N_511,In_199,In_173);
and U512 (N_512,In_160,In_478);
or U513 (N_513,In_240,In_301);
nor U514 (N_514,In_117,In_57);
and U515 (N_515,In_167,In_126);
and U516 (N_516,In_277,In_211);
and U517 (N_517,In_73,In_20);
nor U518 (N_518,In_97,In_251);
nand U519 (N_519,In_44,In_369);
or U520 (N_520,In_116,In_55);
or U521 (N_521,In_346,In_29);
nor U522 (N_522,In_488,In_220);
nand U523 (N_523,In_300,In_362);
nand U524 (N_524,In_293,In_365);
or U525 (N_525,In_402,In_42);
or U526 (N_526,In_427,In_283);
and U527 (N_527,In_405,In_345);
and U528 (N_528,In_438,In_240);
xor U529 (N_529,In_174,In_163);
nor U530 (N_530,In_65,In_472);
nor U531 (N_531,In_382,In_98);
nand U532 (N_532,In_185,In_89);
or U533 (N_533,In_408,In_10);
xnor U534 (N_534,In_446,In_391);
nand U535 (N_535,In_71,In_23);
nand U536 (N_536,In_418,In_173);
xnor U537 (N_537,In_255,In_31);
and U538 (N_538,In_313,In_315);
or U539 (N_539,In_133,In_184);
and U540 (N_540,In_282,In_164);
or U541 (N_541,In_322,In_443);
nor U542 (N_542,In_457,In_425);
xor U543 (N_543,In_147,In_306);
nand U544 (N_544,In_471,In_261);
nand U545 (N_545,In_472,In_475);
nand U546 (N_546,In_224,In_123);
xnor U547 (N_547,In_69,In_66);
nand U548 (N_548,In_271,In_72);
and U549 (N_549,In_376,In_368);
and U550 (N_550,In_173,In_124);
and U551 (N_551,In_346,In_219);
xor U552 (N_552,In_410,In_201);
xnor U553 (N_553,In_72,In_63);
and U554 (N_554,In_48,In_56);
nand U555 (N_555,In_70,In_419);
nor U556 (N_556,In_301,In_69);
nand U557 (N_557,In_418,In_200);
nand U558 (N_558,In_314,In_360);
nor U559 (N_559,In_497,In_143);
xor U560 (N_560,In_306,In_77);
nor U561 (N_561,In_70,In_295);
or U562 (N_562,In_198,In_394);
nand U563 (N_563,In_96,In_328);
or U564 (N_564,In_36,In_218);
xnor U565 (N_565,In_65,In_398);
or U566 (N_566,In_33,In_118);
nor U567 (N_567,In_499,In_147);
and U568 (N_568,In_60,In_339);
nor U569 (N_569,In_298,In_324);
nand U570 (N_570,In_314,In_126);
xor U571 (N_571,In_440,In_303);
xnor U572 (N_572,In_271,In_482);
nand U573 (N_573,In_140,In_485);
nor U574 (N_574,In_297,In_384);
xnor U575 (N_575,In_113,In_452);
and U576 (N_576,In_161,In_302);
xnor U577 (N_577,In_267,In_377);
nor U578 (N_578,In_33,In_423);
xnor U579 (N_579,In_305,In_392);
and U580 (N_580,In_43,In_326);
nand U581 (N_581,In_141,In_171);
and U582 (N_582,In_356,In_423);
and U583 (N_583,In_480,In_12);
nand U584 (N_584,In_166,In_280);
and U585 (N_585,In_95,In_210);
nand U586 (N_586,In_426,In_137);
nand U587 (N_587,In_392,In_429);
nor U588 (N_588,In_192,In_422);
or U589 (N_589,In_70,In_420);
nand U590 (N_590,In_217,In_84);
xnor U591 (N_591,In_171,In_448);
xor U592 (N_592,In_61,In_281);
xor U593 (N_593,In_97,In_79);
nor U594 (N_594,In_247,In_225);
or U595 (N_595,In_381,In_403);
nand U596 (N_596,In_177,In_450);
and U597 (N_597,In_327,In_80);
nand U598 (N_598,In_189,In_288);
or U599 (N_599,In_154,In_174);
and U600 (N_600,In_366,In_407);
nand U601 (N_601,In_417,In_205);
or U602 (N_602,In_235,In_54);
and U603 (N_603,In_423,In_340);
or U604 (N_604,In_126,In_84);
and U605 (N_605,In_153,In_50);
xnor U606 (N_606,In_12,In_7);
nand U607 (N_607,In_251,In_255);
xor U608 (N_608,In_0,In_15);
nand U609 (N_609,In_487,In_401);
and U610 (N_610,In_169,In_145);
or U611 (N_611,In_436,In_426);
and U612 (N_612,In_101,In_432);
or U613 (N_613,In_321,In_481);
or U614 (N_614,In_157,In_420);
or U615 (N_615,In_119,In_54);
nor U616 (N_616,In_413,In_421);
xnor U617 (N_617,In_252,In_48);
nand U618 (N_618,In_54,In_16);
nand U619 (N_619,In_427,In_397);
nor U620 (N_620,In_413,In_215);
or U621 (N_621,In_466,In_153);
nand U622 (N_622,In_357,In_477);
xnor U623 (N_623,In_361,In_57);
nand U624 (N_624,In_269,In_176);
xnor U625 (N_625,In_309,In_425);
nand U626 (N_626,In_482,In_410);
nor U627 (N_627,In_206,In_150);
or U628 (N_628,In_416,In_340);
or U629 (N_629,In_447,In_180);
xnor U630 (N_630,In_408,In_295);
xor U631 (N_631,In_146,In_156);
nand U632 (N_632,In_31,In_195);
nand U633 (N_633,In_89,In_382);
xor U634 (N_634,In_63,In_343);
or U635 (N_635,In_466,In_2);
and U636 (N_636,In_133,In_421);
nand U637 (N_637,In_445,In_491);
or U638 (N_638,In_393,In_216);
nor U639 (N_639,In_67,In_443);
or U640 (N_640,In_180,In_185);
nor U641 (N_641,In_107,In_289);
nor U642 (N_642,In_364,In_325);
nand U643 (N_643,In_303,In_89);
nand U644 (N_644,In_477,In_8);
or U645 (N_645,In_435,In_359);
and U646 (N_646,In_369,In_400);
nand U647 (N_647,In_137,In_119);
nand U648 (N_648,In_441,In_144);
nand U649 (N_649,In_432,In_374);
or U650 (N_650,In_143,In_193);
nor U651 (N_651,In_286,In_299);
xnor U652 (N_652,In_123,In_442);
nand U653 (N_653,In_456,In_251);
nand U654 (N_654,In_272,In_45);
nand U655 (N_655,In_405,In_239);
or U656 (N_656,In_73,In_310);
and U657 (N_657,In_422,In_242);
xor U658 (N_658,In_349,In_32);
and U659 (N_659,In_246,In_251);
or U660 (N_660,In_278,In_118);
and U661 (N_661,In_358,In_106);
nand U662 (N_662,In_140,In_419);
nor U663 (N_663,In_400,In_5);
nand U664 (N_664,In_342,In_274);
xor U665 (N_665,In_287,In_222);
xor U666 (N_666,In_334,In_130);
xnor U667 (N_667,In_158,In_347);
or U668 (N_668,In_347,In_461);
xor U669 (N_669,In_333,In_97);
or U670 (N_670,In_302,In_277);
or U671 (N_671,In_278,In_40);
and U672 (N_672,In_266,In_203);
xnor U673 (N_673,In_86,In_37);
or U674 (N_674,In_282,In_48);
xnor U675 (N_675,In_483,In_285);
nor U676 (N_676,In_74,In_371);
nor U677 (N_677,In_399,In_296);
xor U678 (N_678,In_105,In_176);
xnor U679 (N_679,In_76,In_458);
nor U680 (N_680,In_129,In_322);
nand U681 (N_681,In_117,In_268);
nand U682 (N_682,In_445,In_171);
or U683 (N_683,In_456,In_313);
or U684 (N_684,In_355,In_159);
nor U685 (N_685,In_239,In_71);
nand U686 (N_686,In_91,In_0);
nor U687 (N_687,In_287,In_201);
nand U688 (N_688,In_249,In_428);
nor U689 (N_689,In_494,In_40);
xor U690 (N_690,In_206,In_478);
nand U691 (N_691,In_194,In_393);
or U692 (N_692,In_436,In_62);
and U693 (N_693,In_162,In_276);
nand U694 (N_694,In_78,In_98);
and U695 (N_695,In_219,In_317);
nand U696 (N_696,In_56,In_259);
nor U697 (N_697,In_448,In_89);
and U698 (N_698,In_306,In_426);
nand U699 (N_699,In_258,In_190);
nand U700 (N_700,In_383,In_170);
or U701 (N_701,In_103,In_422);
xnor U702 (N_702,In_488,In_281);
xnor U703 (N_703,In_404,In_330);
xor U704 (N_704,In_206,In_156);
and U705 (N_705,In_108,In_251);
nand U706 (N_706,In_296,In_437);
or U707 (N_707,In_183,In_253);
and U708 (N_708,In_197,In_201);
or U709 (N_709,In_466,In_346);
xnor U710 (N_710,In_265,In_209);
or U711 (N_711,In_32,In_121);
nand U712 (N_712,In_486,In_459);
nand U713 (N_713,In_497,In_458);
and U714 (N_714,In_202,In_250);
nand U715 (N_715,In_135,In_145);
or U716 (N_716,In_402,In_204);
and U717 (N_717,In_315,In_361);
nand U718 (N_718,In_383,In_281);
xnor U719 (N_719,In_296,In_153);
xnor U720 (N_720,In_165,In_24);
xnor U721 (N_721,In_134,In_248);
nand U722 (N_722,In_406,In_38);
nor U723 (N_723,In_275,In_105);
xor U724 (N_724,In_241,In_207);
nand U725 (N_725,In_59,In_182);
nand U726 (N_726,In_280,In_3);
nand U727 (N_727,In_58,In_297);
nand U728 (N_728,In_12,In_254);
or U729 (N_729,In_415,In_374);
nand U730 (N_730,In_35,In_44);
xnor U731 (N_731,In_251,In_430);
nor U732 (N_732,In_451,In_452);
nor U733 (N_733,In_446,In_31);
and U734 (N_734,In_324,In_150);
nor U735 (N_735,In_363,In_399);
or U736 (N_736,In_71,In_476);
nand U737 (N_737,In_143,In_394);
xor U738 (N_738,In_175,In_329);
nor U739 (N_739,In_474,In_220);
nor U740 (N_740,In_236,In_335);
nor U741 (N_741,In_213,In_440);
or U742 (N_742,In_281,In_356);
nor U743 (N_743,In_333,In_331);
or U744 (N_744,In_207,In_476);
nor U745 (N_745,In_70,In_275);
nor U746 (N_746,In_486,In_457);
xor U747 (N_747,In_457,In_54);
xor U748 (N_748,In_199,In_289);
xnor U749 (N_749,In_193,In_374);
or U750 (N_750,N_176,N_481);
xnor U751 (N_751,N_547,N_265);
xnor U752 (N_752,N_624,N_68);
or U753 (N_753,N_454,N_324);
or U754 (N_754,N_46,N_183);
and U755 (N_755,N_720,N_269);
nor U756 (N_756,N_107,N_270);
nor U757 (N_757,N_552,N_337);
and U758 (N_758,N_210,N_313);
or U759 (N_759,N_19,N_274);
and U760 (N_760,N_302,N_30);
nand U761 (N_761,N_564,N_241);
or U762 (N_762,N_296,N_194);
nor U763 (N_763,N_96,N_698);
and U764 (N_764,N_204,N_66);
xor U765 (N_765,N_655,N_600);
xor U766 (N_766,N_128,N_171);
and U767 (N_767,N_160,N_81);
xnor U768 (N_768,N_432,N_705);
and U769 (N_769,N_189,N_669);
and U770 (N_770,N_122,N_315);
and U771 (N_771,N_246,N_277);
and U772 (N_772,N_629,N_214);
or U773 (N_773,N_403,N_587);
or U774 (N_774,N_548,N_649);
or U775 (N_775,N_380,N_222);
xnor U776 (N_776,N_163,N_557);
xor U777 (N_777,N_240,N_43);
or U778 (N_778,N_563,N_331);
xor U779 (N_779,N_44,N_436);
or U780 (N_780,N_47,N_111);
and U781 (N_781,N_259,N_482);
nor U782 (N_782,N_650,N_4);
nand U783 (N_783,N_80,N_499);
xnor U784 (N_784,N_585,N_492);
nand U785 (N_785,N_400,N_618);
or U786 (N_786,N_441,N_479);
nand U787 (N_787,N_673,N_369);
nor U788 (N_788,N_622,N_376);
and U789 (N_789,N_472,N_565);
and U790 (N_790,N_249,N_219);
nand U791 (N_791,N_465,N_216);
or U792 (N_792,N_459,N_395);
and U793 (N_793,N_474,N_155);
xnor U794 (N_794,N_97,N_736);
and U795 (N_795,N_225,N_575);
nor U796 (N_796,N_693,N_642);
xor U797 (N_797,N_312,N_31);
and U798 (N_798,N_527,N_363);
and U799 (N_799,N_560,N_182);
or U800 (N_800,N_540,N_298);
xnor U801 (N_801,N_62,N_3);
and U802 (N_802,N_491,N_330);
xor U803 (N_803,N_130,N_581);
and U804 (N_804,N_285,N_672);
and U805 (N_805,N_319,N_228);
nand U806 (N_806,N_251,N_407);
nor U807 (N_807,N_687,N_351);
xnor U808 (N_808,N_510,N_2);
or U809 (N_809,N_706,N_52);
and U810 (N_810,N_341,N_645);
or U811 (N_811,N_725,N_694);
xnor U812 (N_812,N_686,N_635);
xor U813 (N_813,N_5,N_9);
nand U814 (N_814,N_316,N_367);
xor U815 (N_815,N_539,N_93);
xor U816 (N_816,N_192,N_737);
or U817 (N_817,N_731,N_524);
and U818 (N_818,N_48,N_431);
nand U819 (N_819,N_411,N_28);
or U820 (N_820,N_250,N_89);
or U821 (N_821,N_385,N_551);
and U822 (N_822,N_329,N_21);
nand U823 (N_823,N_724,N_484);
nor U824 (N_824,N_289,N_100);
and U825 (N_825,N_701,N_72);
or U826 (N_826,N_366,N_397);
nor U827 (N_827,N_136,N_476);
xnor U828 (N_828,N_461,N_384);
and U829 (N_829,N_180,N_446);
nand U830 (N_830,N_166,N_118);
and U831 (N_831,N_55,N_8);
nor U832 (N_832,N_526,N_729);
nand U833 (N_833,N_20,N_27);
nand U834 (N_834,N_389,N_239);
nor U835 (N_835,N_158,N_511);
xnor U836 (N_836,N_417,N_595);
nand U837 (N_837,N_414,N_447);
and U838 (N_838,N_311,N_606);
and U839 (N_839,N_625,N_735);
or U840 (N_840,N_50,N_456);
or U841 (N_841,N_279,N_549);
and U842 (N_842,N_79,N_742);
and U843 (N_843,N_119,N_36);
xnor U844 (N_844,N_611,N_231);
nor U845 (N_845,N_323,N_267);
xnor U846 (N_846,N_147,N_434);
or U847 (N_847,N_37,N_377);
or U848 (N_848,N_309,N_238);
nor U849 (N_849,N_576,N_232);
nor U850 (N_850,N_318,N_18);
or U851 (N_851,N_556,N_151);
nand U852 (N_852,N_691,N_747);
nand U853 (N_853,N_139,N_22);
and U854 (N_854,N_467,N_378);
nor U855 (N_855,N_442,N_105);
or U856 (N_856,N_390,N_42);
nor U857 (N_857,N_102,N_51);
and U858 (N_858,N_17,N_708);
or U859 (N_859,N_45,N_373);
and U860 (N_860,N_498,N_525);
xor U861 (N_861,N_264,N_266);
xnor U862 (N_862,N_577,N_541);
or U863 (N_863,N_658,N_529);
or U864 (N_864,N_272,N_418);
nand U865 (N_865,N_327,N_26);
nand U866 (N_866,N_332,N_416);
nand U867 (N_867,N_697,N_356);
xor U868 (N_868,N_590,N_170);
xnor U869 (N_869,N_670,N_457);
and U870 (N_870,N_471,N_174);
xnor U871 (N_871,N_287,N_288);
and U872 (N_872,N_678,N_15);
nand U873 (N_873,N_480,N_294);
or U874 (N_874,N_199,N_184);
xor U875 (N_875,N_344,N_514);
nand U876 (N_876,N_388,N_534);
nor U877 (N_877,N_743,N_383);
and U878 (N_878,N_634,N_382);
and U879 (N_879,N_544,N_610);
and U880 (N_880,N_71,N_92);
nor U881 (N_881,N_515,N_602);
xnor U882 (N_882,N_715,N_64);
nor U883 (N_883,N_433,N_6);
and U884 (N_884,N_229,N_252);
xor U885 (N_885,N_520,N_109);
nand U886 (N_886,N_710,N_223);
nor U887 (N_887,N_404,N_422);
nand U888 (N_888,N_116,N_579);
nor U889 (N_889,N_732,N_340);
and U890 (N_890,N_489,N_127);
nor U891 (N_891,N_640,N_509);
xnor U892 (N_892,N_464,N_500);
nor U893 (N_893,N_521,N_545);
nand U894 (N_894,N_322,N_550);
and U895 (N_895,N_745,N_167);
nor U896 (N_896,N_603,N_343);
nor U897 (N_897,N_33,N_11);
nor U898 (N_898,N_614,N_198);
and U899 (N_899,N_609,N_7);
nand U900 (N_900,N_106,N_643);
or U901 (N_901,N_748,N_202);
xnor U902 (N_902,N_501,N_25);
and U903 (N_903,N_676,N_409);
and U904 (N_904,N_588,N_387);
xnor U905 (N_905,N_451,N_439);
nand U906 (N_906,N_230,N_601);
and U907 (N_907,N_712,N_38);
nor U908 (N_908,N_94,N_468);
nor U909 (N_909,N_16,N_365);
nor U910 (N_910,N_435,N_700);
xnor U911 (N_911,N_300,N_161);
xnor U912 (N_912,N_740,N_131);
or U913 (N_913,N_148,N_342);
and U914 (N_914,N_40,N_217);
nor U915 (N_915,N_469,N_352);
nor U916 (N_916,N_683,N_34);
nor U917 (N_917,N_145,N_211);
nand U918 (N_918,N_473,N_716);
xor U919 (N_919,N_412,N_584);
nand U920 (N_920,N_739,N_195);
xnor U921 (N_921,N_371,N_205);
xnor U922 (N_922,N_206,N_651);
nand U923 (N_923,N_320,N_159);
or U924 (N_924,N_664,N_717);
or U925 (N_925,N_67,N_727);
or U926 (N_926,N_426,N_535);
nand U927 (N_927,N_310,N_76);
or U928 (N_928,N_644,N_162);
and U929 (N_929,N_70,N_359);
or U930 (N_930,N_522,N_637);
or U931 (N_931,N_227,N_314);
or U932 (N_932,N_255,N_621);
xor U933 (N_933,N_408,N_69);
nand U934 (N_934,N_680,N_262);
and U935 (N_935,N_734,N_589);
xor U936 (N_936,N_391,N_140);
or U937 (N_937,N_630,N_592);
nor U938 (N_938,N_84,N_104);
or U939 (N_939,N_536,N_428);
and U940 (N_940,N_455,N_623);
and U941 (N_941,N_172,N_233);
and U942 (N_942,N_684,N_349);
nand U943 (N_943,N_675,N_627);
nand U944 (N_944,N_236,N_306);
nor U945 (N_945,N_628,N_90);
and U946 (N_946,N_78,N_574);
xor U947 (N_947,N_150,N_244);
nand U948 (N_948,N_487,N_242);
nor U949 (N_949,N_125,N_113);
nand U950 (N_950,N_23,N_87);
and U951 (N_951,N_396,N_690);
nor U952 (N_952,N_243,N_512);
xnor U953 (N_953,N_613,N_596);
nand U954 (N_954,N_594,N_413);
nor U955 (N_955,N_452,N_98);
and U956 (N_956,N_646,N_695);
and U957 (N_957,N_478,N_129);
and U958 (N_958,N_215,N_709);
nand U959 (N_959,N_304,N_667);
nand U960 (N_960,N_141,N_677);
nor U961 (N_961,N_401,N_164);
xnor U962 (N_962,N_201,N_308);
xnor U963 (N_963,N_507,N_247);
nor U964 (N_964,N_604,N_714);
nor U965 (N_965,N_718,N_399);
xor U966 (N_966,N_293,N_0);
and U967 (N_967,N_704,N_533);
or U968 (N_968,N_746,N_490);
or U969 (N_969,N_286,N_420);
xor U970 (N_970,N_57,N_144);
nor U971 (N_971,N_336,N_271);
and U972 (N_972,N_448,N_453);
and U973 (N_973,N_460,N_493);
nor U974 (N_974,N_538,N_537);
or U975 (N_975,N_32,N_186);
nand U976 (N_976,N_95,N_555);
nand U977 (N_977,N_398,N_633);
nand U978 (N_978,N_276,N_405);
nand U979 (N_979,N_652,N_462);
nand U980 (N_980,N_13,N_504);
or U981 (N_981,N_273,N_593);
or U982 (N_982,N_438,N_368);
xnor U983 (N_983,N_466,N_364);
and U984 (N_984,N_82,N_513);
nor U985 (N_985,N_234,N_347);
or U986 (N_986,N_553,N_370);
or U987 (N_987,N_648,N_245);
and U988 (N_988,N_165,N_185);
nor U989 (N_989,N_253,N_599);
xnor U990 (N_990,N_280,N_357);
xnor U991 (N_991,N_696,N_662);
nor U992 (N_992,N_179,N_354);
and U993 (N_993,N_224,N_458);
xnor U994 (N_994,N_138,N_61);
nor U995 (N_995,N_738,N_361);
and U996 (N_996,N_263,N_711);
nor U997 (N_997,N_719,N_730);
nor U998 (N_998,N_260,N_543);
and U999 (N_999,N_10,N_620);
nand U1000 (N_1000,N_406,N_668);
nor U1001 (N_1001,N_49,N_12);
xor U1002 (N_1002,N_117,N_218);
nand U1003 (N_1003,N_374,N_674);
nor U1004 (N_1004,N_749,N_134);
xnor U1005 (N_1005,N_567,N_608);
nor U1006 (N_1006,N_722,N_74);
nand U1007 (N_1007,N_578,N_566);
xor U1008 (N_1008,N_108,N_187);
xor U1009 (N_1009,N_591,N_77);
nand U1010 (N_1010,N_58,N_124);
and U1011 (N_1011,N_605,N_339);
nor U1012 (N_1012,N_149,N_350);
or U1013 (N_1013,N_157,N_641);
nand U1014 (N_1014,N_723,N_483);
and U1015 (N_1015,N_317,N_132);
nand U1016 (N_1016,N_326,N_572);
or U1017 (N_1017,N_415,N_427);
xor U1018 (N_1018,N_477,N_307);
or U1019 (N_1019,N_123,N_671);
nand U1020 (N_1020,N_688,N_60);
or U1021 (N_1021,N_99,N_394);
xnor U1022 (N_1022,N_35,N_598);
nor U1023 (N_1023,N_168,N_190);
or U1024 (N_1024,N_505,N_278);
or U1025 (N_1025,N_65,N_663);
nor U1026 (N_1026,N_713,N_386);
xor U1027 (N_1027,N_657,N_532);
or U1028 (N_1028,N_39,N_362);
nand U1029 (N_1029,N_647,N_121);
or U1030 (N_1030,N_86,N_689);
or U1031 (N_1031,N_188,N_665);
nor U1032 (N_1032,N_419,N_424);
nor U1033 (N_1033,N_741,N_290);
nand U1034 (N_1034,N_1,N_226);
or U1035 (N_1035,N_299,N_173);
xor U1036 (N_1036,N_213,N_733);
nor U1037 (N_1037,N_379,N_177);
nand U1038 (N_1038,N_305,N_303);
nand U1039 (N_1039,N_56,N_392);
xnor U1040 (N_1040,N_626,N_91);
xnor U1041 (N_1041,N_220,N_702);
nor U1042 (N_1042,N_568,N_450);
xnor U1043 (N_1043,N_338,N_83);
nand U1044 (N_1044,N_519,N_346);
nor U1045 (N_1045,N_653,N_181);
nand U1046 (N_1046,N_496,N_421);
or U1047 (N_1047,N_393,N_485);
nor U1048 (N_1048,N_410,N_582);
and U1049 (N_1049,N_203,N_169);
or U1050 (N_1050,N_353,N_143);
xnor U1051 (N_1051,N_685,N_573);
and U1052 (N_1052,N_41,N_328);
nor U1053 (N_1053,N_281,N_197);
nand U1054 (N_1054,N_488,N_546);
nor U1055 (N_1055,N_531,N_268);
and U1056 (N_1056,N_728,N_495);
nor U1057 (N_1057,N_444,N_73);
and U1058 (N_1058,N_571,N_191);
or U1059 (N_1059,N_120,N_707);
nand U1060 (N_1060,N_617,N_430);
and U1061 (N_1061,N_517,N_235);
nand U1062 (N_1062,N_744,N_597);
xnor U1063 (N_1063,N_494,N_193);
xor U1064 (N_1064,N_360,N_443);
xor U1065 (N_1065,N_59,N_292);
nand U1066 (N_1066,N_638,N_297);
and U1067 (N_1067,N_348,N_475);
or U1068 (N_1068,N_256,N_660);
and U1069 (N_1069,N_14,N_518);
and U1070 (N_1070,N_196,N_75);
or U1071 (N_1071,N_178,N_153);
nand U1072 (N_1072,N_445,N_24);
nor U1073 (N_1073,N_508,N_569);
nand U1074 (N_1074,N_703,N_135);
and U1075 (N_1075,N_284,N_63);
or U1076 (N_1076,N_321,N_248);
nand U1077 (N_1077,N_142,N_470);
or U1078 (N_1078,N_639,N_679);
and U1079 (N_1079,N_207,N_530);
and U1080 (N_1080,N_152,N_372);
nor U1081 (N_1081,N_291,N_636);
or U1082 (N_1082,N_607,N_523);
xnor U1083 (N_1083,N_682,N_486);
nand U1084 (N_1084,N_381,N_554);
nand U1085 (N_1085,N_133,N_208);
nand U1086 (N_1086,N_275,N_402);
and U1087 (N_1087,N_666,N_542);
xnor U1088 (N_1088,N_502,N_85);
nand U1089 (N_1089,N_692,N_355);
xor U1090 (N_1090,N_112,N_497);
nor U1091 (N_1091,N_570,N_283);
xor U1092 (N_1092,N_257,N_295);
or U1093 (N_1093,N_175,N_333);
nor U1094 (N_1094,N_681,N_154);
nand U1095 (N_1095,N_659,N_146);
xor U1096 (N_1096,N_29,N_423);
nand U1097 (N_1097,N_282,N_221);
and U1098 (N_1098,N_88,N_661);
nand U1099 (N_1099,N_425,N_53);
nand U1100 (N_1100,N_580,N_559);
nor U1101 (N_1101,N_503,N_506);
or U1102 (N_1102,N_516,N_619);
nor U1103 (N_1103,N_632,N_429);
or U1104 (N_1104,N_558,N_654);
nor U1105 (N_1105,N_110,N_334);
and U1106 (N_1106,N_631,N_358);
nor U1107 (N_1107,N_115,N_212);
or U1108 (N_1108,N_726,N_437);
nor U1109 (N_1109,N_615,N_258);
xnor U1110 (N_1110,N_583,N_586);
nand U1111 (N_1111,N_528,N_375);
nand U1112 (N_1112,N_440,N_562);
or U1113 (N_1113,N_103,N_200);
nand U1114 (N_1114,N_54,N_209);
and U1115 (N_1115,N_156,N_301);
nor U1116 (N_1116,N_254,N_463);
nand U1117 (N_1117,N_561,N_126);
nand U1118 (N_1118,N_616,N_101);
xor U1119 (N_1119,N_137,N_612);
xnor U1120 (N_1120,N_325,N_721);
and U1121 (N_1121,N_114,N_345);
nand U1122 (N_1122,N_656,N_261);
xnor U1123 (N_1123,N_335,N_449);
xor U1124 (N_1124,N_699,N_237);
nand U1125 (N_1125,N_520,N_605);
xor U1126 (N_1126,N_11,N_543);
nand U1127 (N_1127,N_580,N_5);
and U1128 (N_1128,N_5,N_192);
nor U1129 (N_1129,N_24,N_507);
or U1130 (N_1130,N_742,N_321);
or U1131 (N_1131,N_556,N_587);
nor U1132 (N_1132,N_245,N_177);
xor U1133 (N_1133,N_301,N_539);
nand U1134 (N_1134,N_68,N_279);
and U1135 (N_1135,N_95,N_624);
nor U1136 (N_1136,N_273,N_397);
xnor U1137 (N_1137,N_199,N_59);
xor U1138 (N_1138,N_109,N_483);
xor U1139 (N_1139,N_571,N_583);
and U1140 (N_1140,N_502,N_716);
xnor U1141 (N_1141,N_494,N_459);
nand U1142 (N_1142,N_633,N_632);
and U1143 (N_1143,N_208,N_381);
nand U1144 (N_1144,N_217,N_747);
nor U1145 (N_1145,N_685,N_590);
or U1146 (N_1146,N_538,N_101);
nor U1147 (N_1147,N_588,N_313);
or U1148 (N_1148,N_585,N_16);
xor U1149 (N_1149,N_543,N_307);
xnor U1150 (N_1150,N_205,N_670);
or U1151 (N_1151,N_81,N_456);
nand U1152 (N_1152,N_243,N_382);
nor U1153 (N_1153,N_356,N_562);
or U1154 (N_1154,N_662,N_250);
and U1155 (N_1155,N_508,N_446);
nor U1156 (N_1156,N_717,N_6);
or U1157 (N_1157,N_209,N_230);
and U1158 (N_1158,N_344,N_106);
or U1159 (N_1159,N_410,N_244);
xor U1160 (N_1160,N_346,N_168);
nor U1161 (N_1161,N_148,N_644);
or U1162 (N_1162,N_371,N_598);
and U1163 (N_1163,N_300,N_588);
xor U1164 (N_1164,N_286,N_739);
nor U1165 (N_1165,N_210,N_335);
nand U1166 (N_1166,N_212,N_40);
xnor U1167 (N_1167,N_198,N_223);
xnor U1168 (N_1168,N_163,N_304);
and U1169 (N_1169,N_617,N_168);
nor U1170 (N_1170,N_57,N_707);
xnor U1171 (N_1171,N_158,N_233);
xor U1172 (N_1172,N_260,N_280);
xor U1173 (N_1173,N_83,N_667);
nand U1174 (N_1174,N_573,N_333);
and U1175 (N_1175,N_540,N_437);
or U1176 (N_1176,N_93,N_550);
or U1177 (N_1177,N_634,N_125);
nor U1178 (N_1178,N_437,N_391);
xnor U1179 (N_1179,N_38,N_158);
nand U1180 (N_1180,N_440,N_682);
and U1181 (N_1181,N_482,N_520);
xor U1182 (N_1182,N_557,N_108);
nand U1183 (N_1183,N_532,N_319);
nand U1184 (N_1184,N_246,N_622);
or U1185 (N_1185,N_275,N_641);
nand U1186 (N_1186,N_322,N_679);
and U1187 (N_1187,N_366,N_441);
nand U1188 (N_1188,N_404,N_609);
nor U1189 (N_1189,N_278,N_415);
nand U1190 (N_1190,N_169,N_661);
and U1191 (N_1191,N_485,N_392);
xnor U1192 (N_1192,N_358,N_41);
xnor U1193 (N_1193,N_405,N_469);
nand U1194 (N_1194,N_747,N_652);
and U1195 (N_1195,N_622,N_89);
or U1196 (N_1196,N_711,N_524);
nor U1197 (N_1197,N_580,N_308);
nand U1198 (N_1198,N_747,N_138);
nor U1199 (N_1199,N_35,N_68);
xnor U1200 (N_1200,N_731,N_349);
nand U1201 (N_1201,N_595,N_114);
and U1202 (N_1202,N_630,N_41);
and U1203 (N_1203,N_183,N_108);
or U1204 (N_1204,N_213,N_514);
xor U1205 (N_1205,N_259,N_128);
or U1206 (N_1206,N_568,N_432);
and U1207 (N_1207,N_710,N_47);
nand U1208 (N_1208,N_375,N_62);
and U1209 (N_1209,N_441,N_142);
xnor U1210 (N_1210,N_586,N_426);
xor U1211 (N_1211,N_434,N_486);
and U1212 (N_1212,N_590,N_177);
xor U1213 (N_1213,N_237,N_564);
xnor U1214 (N_1214,N_418,N_39);
nand U1215 (N_1215,N_720,N_743);
and U1216 (N_1216,N_676,N_522);
nand U1217 (N_1217,N_114,N_407);
or U1218 (N_1218,N_0,N_450);
or U1219 (N_1219,N_744,N_100);
nor U1220 (N_1220,N_63,N_622);
or U1221 (N_1221,N_527,N_723);
or U1222 (N_1222,N_99,N_668);
xnor U1223 (N_1223,N_500,N_545);
or U1224 (N_1224,N_462,N_70);
or U1225 (N_1225,N_98,N_336);
nor U1226 (N_1226,N_643,N_12);
or U1227 (N_1227,N_92,N_127);
nand U1228 (N_1228,N_259,N_286);
xor U1229 (N_1229,N_458,N_618);
and U1230 (N_1230,N_21,N_342);
xor U1231 (N_1231,N_107,N_702);
and U1232 (N_1232,N_654,N_286);
nand U1233 (N_1233,N_475,N_405);
nor U1234 (N_1234,N_43,N_640);
nand U1235 (N_1235,N_184,N_354);
nand U1236 (N_1236,N_82,N_268);
nor U1237 (N_1237,N_546,N_1);
and U1238 (N_1238,N_368,N_457);
nand U1239 (N_1239,N_690,N_86);
nor U1240 (N_1240,N_689,N_675);
nand U1241 (N_1241,N_428,N_710);
or U1242 (N_1242,N_265,N_116);
nor U1243 (N_1243,N_206,N_641);
and U1244 (N_1244,N_638,N_334);
xnor U1245 (N_1245,N_90,N_594);
nand U1246 (N_1246,N_296,N_375);
nand U1247 (N_1247,N_31,N_647);
xor U1248 (N_1248,N_157,N_470);
nor U1249 (N_1249,N_307,N_490);
xnor U1250 (N_1250,N_191,N_421);
xor U1251 (N_1251,N_228,N_144);
nand U1252 (N_1252,N_106,N_736);
nor U1253 (N_1253,N_222,N_445);
xnor U1254 (N_1254,N_203,N_740);
and U1255 (N_1255,N_524,N_366);
nand U1256 (N_1256,N_741,N_642);
xnor U1257 (N_1257,N_480,N_575);
or U1258 (N_1258,N_251,N_542);
or U1259 (N_1259,N_449,N_142);
xor U1260 (N_1260,N_245,N_11);
or U1261 (N_1261,N_50,N_711);
or U1262 (N_1262,N_525,N_161);
or U1263 (N_1263,N_605,N_439);
nor U1264 (N_1264,N_623,N_421);
and U1265 (N_1265,N_622,N_175);
nor U1266 (N_1266,N_55,N_704);
or U1267 (N_1267,N_421,N_346);
nand U1268 (N_1268,N_442,N_643);
xnor U1269 (N_1269,N_502,N_615);
or U1270 (N_1270,N_371,N_545);
or U1271 (N_1271,N_31,N_86);
or U1272 (N_1272,N_228,N_612);
nor U1273 (N_1273,N_653,N_739);
or U1274 (N_1274,N_274,N_71);
and U1275 (N_1275,N_132,N_288);
xor U1276 (N_1276,N_646,N_371);
or U1277 (N_1277,N_235,N_307);
nor U1278 (N_1278,N_282,N_243);
nand U1279 (N_1279,N_422,N_9);
or U1280 (N_1280,N_476,N_14);
nand U1281 (N_1281,N_538,N_355);
nor U1282 (N_1282,N_705,N_126);
nand U1283 (N_1283,N_588,N_529);
xnor U1284 (N_1284,N_326,N_589);
nand U1285 (N_1285,N_580,N_156);
or U1286 (N_1286,N_476,N_480);
and U1287 (N_1287,N_79,N_184);
or U1288 (N_1288,N_576,N_438);
xor U1289 (N_1289,N_120,N_111);
nor U1290 (N_1290,N_452,N_470);
nor U1291 (N_1291,N_439,N_334);
xnor U1292 (N_1292,N_601,N_627);
or U1293 (N_1293,N_312,N_536);
xnor U1294 (N_1294,N_26,N_605);
xor U1295 (N_1295,N_327,N_270);
or U1296 (N_1296,N_345,N_590);
xor U1297 (N_1297,N_101,N_13);
or U1298 (N_1298,N_95,N_199);
xor U1299 (N_1299,N_299,N_636);
nor U1300 (N_1300,N_589,N_66);
or U1301 (N_1301,N_580,N_491);
or U1302 (N_1302,N_33,N_23);
and U1303 (N_1303,N_1,N_22);
xnor U1304 (N_1304,N_637,N_423);
nor U1305 (N_1305,N_249,N_308);
or U1306 (N_1306,N_604,N_724);
nand U1307 (N_1307,N_533,N_85);
and U1308 (N_1308,N_575,N_384);
nor U1309 (N_1309,N_696,N_619);
and U1310 (N_1310,N_508,N_171);
or U1311 (N_1311,N_292,N_506);
and U1312 (N_1312,N_371,N_449);
or U1313 (N_1313,N_362,N_723);
nor U1314 (N_1314,N_551,N_242);
nand U1315 (N_1315,N_183,N_390);
or U1316 (N_1316,N_218,N_466);
and U1317 (N_1317,N_384,N_244);
xor U1318 (N_1318,N_706,N_169);
and U1319 (N_1319,N_441,N_452);
nor U1320 (N_1320,N_734,N_666);
nor U1321 (N_1321,N_122,N_497);
nand U1322 (N_1322,N_457,N_648);
xnor U1323 (N_1323,N_541,N_360);
xnor U1324 (N_1324,N_142,N_393);
and U1325 (N_1325,N_416,N_454);
xor U1326 (N_1326,N_313,N_329);
or U1327 (N_1327,N_238,N_18);
nor U1328 (N_1328,N_286,N_550);
or U1329 (N_1329,N_220,N_637);
or U1330 (N_1330,N_724,N_590);
and U1331 (N_1331,N_170,N_74);
nand U1332 (N_1332,N_311,N_428);
nor U1333 (N_1333,N_656,N_499);
xor U1334 (N_1334,N_127,N_116);
nand U1335 (N_1335,N_158,N_459);
or U1336 (N_1336,N_35,N_275);
xnor U1337 (N_1337,N_325,N_240);
nor U1338 (N_1338,N_548,N_271);
and U1339 (N_1339,N_184,N_120);
or U1340 (N_1340,N_674,N_596);
or U1341 (N_1341,N_654,N_98);
or U1342 (N_1342,N_293,N_182);
nor U1343 (N_1343,N_183,N_510);
and U1344 (N_1344,N_401,N_382);
and U1345 (N_1345,N_327,N_500);
xor U1346 (N_1346,N_724,N_721);
nand U1347 (N_1347,N_718,N_639);
nor U1348 (N_1348,N_433,N_412);
nand U1349 (N_1349,N_67,N_662);
xnor U1350 (N_1350,N_531,N_264);
nand U1351 (N_1351,N_75,N_399);
or U1352 (N_1352,N_202,N_568);
or U1353 (N_1353,N_677,N_389);
nand U1354 (N_1354,N_487,N_444);
xor U1355 (N_1355,N_612,N_232);
or U1356 (N_1356,N_239,N_549);
and U1357 (N_1357,N_488,N_183);
nand U1358 (N_1358,N_725,N_22);
xnor U1359 (N_1359,N_100,N_422);
and U1360 (N_1360,N_629,N_243);
xnor U1361 (N_1361,N_293,N_699);
or U1362 (N_1362,N_206,N_356);
nand U1363 (N_1363,N_75,N_361);
nand U1364 (N_1364,N_147,N_406);
nor U1365 (N_1365,N_151,N_227);
nand U1366 (N_1366,N_308,N_545);
nand U1367 (N_1367,N_470,N_609);
nand U1368 (N_1368,N_229,N_543);
nor U1369 (N_1369,N_415,N_600);
nand U1370 (N_1370,N_387,N_570);
xor U1371 (N_1371,N_421,N_201);
nand U1372 (N_1372,N_441,N_644);
xor U1373 (N_1373,N_469,N_421);
or U1374 (N_1374,N_560,N_340);
nor U1375 (N_1375,N_549,N_624);
nand U1376 (N_1376,N_540,N_43);
nand U1377 (N_1377,N_210,N_660);
and U1378 (N_1378,N_239,N_457);
nand U1379 (N_1379,N_62,N_261);
nor U1380 (N_1380,N_70,N_41);
or U1381 (N_1381,N_473,N_443);
nor U1382 (N_1382,N_330,N_420);
nand U1383 (N_1383,N_18,N_192);
nor U1384 (N_1384,N_284,N_303);
nand U1385 (N_1385,N_215,N_107);
nor U1386 (N_1386,N_583,N_446);
or U1387 (N_1387,N_206,N_366);
xnor U1388 (N_1388,N_354,N_34);
xnor U1389 (N_1389,N_452,N_68);
xor U1390 (N_1390,N_73,N_507);
nor U1391 (N_1391,N_354,N_112);
nand U1392 (N_1392,N_641,N_307);
nor U1393 (N_1393,N_274,N_338);
or U1394 (N_1394,N_63,N_305);
or U1395 (N_1395,N_449,N_625);
nor U1396 (N_1396,N_610,N_218);
or U1397 (N_1397,N_176,N_233);
nor U1398 (N_1398,N_284,N_296);
nor U1399 (N_1399,N_508,N_325);
xnor U1400 (N_1400,N_476,N_679);
or U1401 (N_1401,N_136,N_43);
and U1402 (N_1402,N_9,N_625);
and U1403 (N_1403,N_331,N_99);
xnor U1404 (N_1404,N_48,N_410);
xnor U1405 (N_1405,N_222,N_612);
or U1406 (N_1406,N_209,N_139);
nand U1407 (N_1407,N_1,N_457);
or U1408 (N_1408,N_576,N_746);
nor U1409 (N_1409,N_671,N_536);
and U1410 (N_1410,N_102,N_346);
and U1411 (N_1411,N_277,N_257);
nor U1412 (N_1412,N_14,N_178);
nor U1413 (N_1413,N_318,N_13);
or U1414 (N_1414,N_479,N_393);
xnor U1415 (N_1415,N_15,N_706);
or U1416 (N_1416,N_652,N_73);
xnor U1417 (N_1417,N_274,N_396);
nor U1418 (N_1418,N_313,N_246);
nor U1419 (N_1419,N_612,N_433);
and U1420 (N_1420,N_399,N_364);
and U1421 (N_1421,N_206,N_673);
and U1422 (N_1422,N_512,N_529);
xor U1423 (N_1423,N_390,N_154);
or U1424 (N_1424,N_64,N_437);
xnor U1425 (N_1425,N_434,N_77);
and U1426 (N_1426,N_566,N_255);
or U1427 (N_1427,N_66,N_166);
xnor U1428 (N_1428,N_213,N_371);
nor U1429 (N_1429,N_599,N_694);
xnor U1430 (N_1430,N_22,N_154);
and U1431 (N_1431,N_665,N_493);
xor U1432 (N_1432,N_481,N_471);
nand U1433 (N_1433,N_607,N_241);
xnor U1434 (N_1434,N_615,N_68);
nand U1435 (N_1435,N_129,N_214);
nand U1436 (N_1436,N_25,N_586);
and U1437 (N_1437,N_567,N_467);
xnor U1438 (N_1438,N_627,N_282);
and U1439 (N_1439,N_116,N_682);
xnor U1440 (N_1440,N_276,N_413);
nor U1441 (N_1441,N_231,N_187);
xnor U1442 (N_1442,N_673,N_457);
and U1443 (N_1443,N_214,N_134);
nand U1444 (N_1444,N_180,N_322);
or U1445 (N_1445,N_199,N_56);
nand U1446 (N_1446,N_146,N_307);
nand U1447 (N_1447,N_245,N_5);
or U1448 (N_1448,N_79,N_740);
and U1449 (N_1449,N_257,N_586);
and U1450 (N_1450,N_360,N_742);
nor U1451 (N_1451,N_292,N_661);
nor U1452 (N_1452,N_343,N_520);
nand U1453 (N_1453,N_401,N_631);
nor U1454 (N_1454,N_704,N_247);
xor U1455 (N_1455,N_446,N_473);
and U1456 (N_1456,N_46,N_474);
nand U1457 (N_1457,N_354,N_11);
xor U1458 (N_1458,N_600,N_565);
and U1459 (N_1459,N_355,N_105);
or U1460 (N_1460,N_336,N_196);
or U1461 (N_1461,N_142,N_491);
or U1462 (N_1462,N_294,N_98);
nand U1463 (N_1463,N_9,N_269);
or U1464 (N_1464,N_653,N_649);
and U1465 (N_1465,N_670,N_185);
or U1466 (N_1466,N_317,N_393);
or U1467 (N_1467,N_515,N_60);
nor U1468 (N_1468,N_118,N_661);
xnor U1469 (N_1469,N_297,N_254);
or U1470 (N_1470,N_509,N_678);
and U1471 (N_1471,N_287,N_238);
nand U1472 (N_1472,N_632,N_64);
xor U1473 (N_1473,N_367,N_579);
or U1474 (N_1474,N_38,N_346);
and U1475 (N_1475,N_719,N_238);
xor U1476 (N_1476,N_381,N_303);
nor U1477 (N_1477,N_473,N_592);
xor U1478 (N_1478,N_517,N_413);
nand U1479 (N_1479,N_542,N_712);
nand U1480 (N_1480,N_84,N_222);
and U1481 (N_1481,N_275,N_78);
or U1482 (N_1482,N_605,N_554);
nand U1483 (N_1483,N_324,N_4);
nand U1484 (N_1484,N_108,N_588);
or U1485 (N_1485,N_624,N_656);
or U1486 (N_1486,N_652,N_408);
xnor U1487 (N_1487,N_31,N_411);
nand U1488 (N_1488,N_264,N_653);
and U1489 (N_1489,N_287,N_527);
and U1490 (N_1490,N_296,N_653);
nand U1491 (N_1491,N_68,N_300);
and U1492 (N_1492,N_251,N_551);
nand U1493 (N_1493,N_18,N_661);
or U1494 (N_1494,N_484,N_514);
or U1495 (N_1495,N_373,N_380);
and U1496 (N_1496,N_228,N_87);
and U1497 (N_1497,N_513,N_404);
or U1498 (N_1498,N_404,N_643);
or U1499 (N_1499,N_235,N_690);
nor U1500 (N_1500,N_1418,N_855);
and U1501 (N_1501,N_1444,N_1295);
xor U1502 (N_1502,N_1394,N_1145);
and U1503 (N_1503,N_1364,N_1196);
xnor U1504 (N_1504,N_1079,N_1319);
xor U1505 (N_1505,N_1450,N_1238);
nor U1506 (N_1506,N_1329,N_1449);
and U1507 (N_1507,N_1351,N_1222);
and U1508 (N_1508,N_994,N_1333);
xor U1509 (N_1509,N_1380,N_999);
or U1510 (N_1510,N_1470,N_926);
or U1511 (N_1511,N_821,N_1378);
nand U1512 (N_1512,N_1382,N_1401);
nand U1513 (N_1513,N_1226,N_856);
or U1514 (N_1514,N_922,N_1147);
xor U1515 (N_1515,N_1135,N_980);
nor U1516 (N_1516,N_844,N_1117);
and U1517 (N_1517,N_1101,N_1198);
nor U1518 (N_1518,N_1395,N_882);
nor U1519 (N_1519,N_1109,N_830);
xnor U1520 (N_1520,N_801,N_1456);
xor U1521 (N_1521,N_1362,N_1331);
nand U1522 (N_1522,N_923,N_1451);
xor U1523 (N_1523,N_967,N_783);
and U1524 (N_1524,N_819,N_1170);
or U1525 (N_1525,N_1471,N_1130);
and U1526 (N_1526,N_1050,N_1320);
and U1527 (N_1527,N_1365,N_1197);
and U1528 (N_1528,N_1439,N_1258);
nand U1529 (N_1529,N_1400,N_1497);
nor U1530 (N_1530,N_1288,N_773);
or U1531 (N_1531,N_917,N_1052);
xnor U1532 (N_1532,N_1324,N_1070);
xor U1533 (N_1533,N_1411,N_786);
nand U1534 (N_1534,N_939,N_1459);
nand U1535 (N_1535,N_787,N_1491);
nand U1536 (N_1536,N_941,N_1097);
nor U1537 (N_1537,N_808,N_832);
nand U1538 (N_1538,N_1321,N_1116);
and U1539 (N_1539,N_1408,N_1367);
xor U1540 (N_1540,N_776,N_1013);
nand U1541 (N_1541,N_1022,N_1448);
nand U1542 (N_1542,N_1091,N_1064);
nor U1543 (N_1543,N_1312,N_1384);
nand U1544 (N_1544,N_1115,N_992);
nand U1545 (N_1545,N_796,N_1330);
nor U1546 (N_1546,N_1006,N_1100);
or U1547 (N_1547,N_1025,N_1252);
nor U1548 (N_1548,N_913,N_777);
or U1549 (N_1549,N_1307,N_1402);
xnor U1550 (N_1550,N_995,N_1447);
nor U1551 (N_1551,N_1202,N_1271);
nand U1552 (N_1552,N_934,N_867);
or U1553 (N_1553,N_909,N_1191);
or U1554 (N_1554,N_1148,N_1298);
nand U1555 (N_1555,N_1166,N_788);
xor U1556 (N_1556,N_1179,N_1088);
xor U1557 (N_1557,N_1421,N_1019);
and U1558 (N_1558,N_1335,N_1363);
xor U1559 (N_1559,N_1140,N_841);
nand U1560 (N_1560,N_842,N_802);
xnor U1561 (N_1561,N_1063,N_766);
nand U1562 (N_1562,N_961,N_816);
nor U1563 (N_1563,N_1205,N_1280);
nand U1564 (N_1564,N_929,N_1247);
nor U1565 (N_1565,N_988,N_814);
xor U1566 (N_1566,N_1262,N_1061);
nor U1567 (N_1567,N_1326,N_858);
xor U1568 (N_1568,N_1424,N_931);
xor U1569 (N_1569,N_1499,N_1003);
and U1570 (N_1570,N_1397,N_1286);
or U1571 (N_1571,N_1094,N_791);
xor U1572 (N_1572,N_803,N_1308);
or U1573 (N_1573,N_1077,N_1478);
and U1574 (N_1574,N_1152,N_1156);
or U1575 (N_1575,N_1095,N_789);
nand U1576 (N_1576,N_1124,N_897);
and U1577 (N_1577,N_1386,N_772);
nand U1578 (N_1578,N_784,N_1347);
xnor U1579 (N_1579,N_1192,N_1492);
xnor U1580 (N_1580,N_893,N_1015);
nand U1581 (N_1581,N_1203,N_1315);
and U1582 (N_1582,N_1241,N_1138);
or U1583 (N_1583,N_1260,N_1187);
nand U1584 (N_1584,N_1043,N_1432);
xor U1585 (N_1585,N_1493,N_1028);
xor U1586 (N_1586,N_1002,N_872);
or U1587 (N_1587,N_1181,N_868);
nor U1588 (N_1588,N_970,N_1127);
nand U1589 (N_1589,N_1428,N_911);
and U1590 (N_1590,N_1165,N_1248);
nand U1591 (N_1591,N_1169,N_1090);
xnor U1592 (N_1592,N_997,N_1009);
nand U1593 (N_1593,N_1318,N_1339);
nor U1594 (N_1594,N_1472,N_876);
nor U1595 (N_1595,N_1162,N_973);
xnor U1596 (N_1596,N_870,N_1008);
and U1597 (N_1597,N_1429,N_1132);
xor U1598 (N_1598,N_1161,N_1361);
xor U1599 (N_1599,N_840,N_906);
nor U1600 (N_1600,N_1246,N_883);
xor U1601 (N_1601,N_1416,N_874);
or U1602 (N_1602,N_958,N_1484);
nor U1603 (N_1603,N_1026,N_985);
or U1604 (N_1604,N_938,N_1149);
nand U1605 (N_1605,N_1306,N_930);
nand U1606 (N_1606,N_1270,N_1186);
nand U1607 (N_1607,N_1084,N_1105);
or U1608 (N_1608,N_1235,N_831);
or U1609 (N_1609,N_1476,N_1427);
or U1610 (N_1610,N_1322,N_1216);
nand U1611 (N_1611,N_850,N_1311);
nor U1612 (N_1612,N_864,N_863);
or U1613 (N_1613,N_1058,N_881);
nand U1614 (N_1614,N_1184,N_822);
nand U1615 (N_1615,N_1004,N_1081);
or U1616 (N_1616,N_891,N_943);
and U1617 (N_1617,N_974,N_779);
and U1618 (N_1618,N_903,N_1431);
nand U1619 (N_1619,N_1388,N_1485);
or U1620 (N_1620,N_1207,N_915);
nand U1621 (N_1621,N_820,N_888);
or U1622 (N_1622,N_1422,N_1236);
xor U1623 (N_1623,N_920,N_1358);
xnor U1624 (N_1624,N_1325,N_957);
xor U1625 (N_1625,N_1349,N_949);
or U1626 (N_1626,N_932,N_1245);
xnor U1627 (N_1627,N_877,N_1419);
or U1628 (N_1628,N_1481,N_990);
nand U1629 (N_1629,N_1264,N_968);
nand U1630 (N_1630,N_1039,N_998);
nand U1631 (N_1631,N_951,N_1218);
xor U1632 (N_1632,N_1167,N_1399);
and U1633 (N_1633,N_1446,N_1385);
or U1634 (N_1634,N_1296,N_948);
and U1635 (N_1635,N_1237,N_1368);
nor U1636 (N_1636,N_817,N_1049);
and U1637 (N_1637,N_1204,N_1305);
and U1638 (N_1638,N_824,N_1182);
nor U1639 (N_1639,N_1338,N_966);
xnor U1640 (N_1640,N_982,N_1060);
xor U1641 (N_1641,N_1377,N_1021);
and U1642 (N_1642,N_1120,N_940);
or U1643 (N_1643,N_1276,N_1030);
nor U1644 (N_1644,N_845,N_1096);
xor U1645 (N_1645,N_1348,N_1461);
and U1646 (N_1646,N_1299,N_795);
nor U1647 (N_1647,N_1035,N_1215);
and U1648 (N_1648,N_1302,N_910);
xor U1649 (N_1649,N_1045,N_1494);
nand U1650 (N_1650,N_1495,N_1406);
nand U1651 (N_1651,N_871,N_828);
and U1652 (N_1652,N_1176,N_1220);
nand U1653 (N_1653,N_1044,N_1265);
nand U1654 (N_1654,N_1212,N_1083);
nor U1655 (N_1655,N_1396,N_1037);
xor U1656 (N_1656,N_1048,N_1137);
xor U1657 (N_1657,N_1445,N_1154);
or U1658 (N_1658,N_759,N_1417);
nor U1659 (N_1659,N_1355,N_1342);
xnor U1660 (N_1660,N_875,N_1407);
nand U1661 (N_1661,N_1332,N_942);
nor U1662 (N_1662,N_1233,N_1200);
and U1663 (N_1663,N_1387,N_1496);
and U1664 (N_1664,N_813,N_849);
and U1665 (N_1665,N_1261,N_1000);
and U1666 (N_1666,N_1389,N_835);
nor U1667 (N_1667,N_1099,N_879);
xnor U1668 (N_1668,N_1125,N_1457);
nand U1669 (N_1669,N_818,N_764);
and U1670 (N_1670,N_1243,N_1278);
nor U1671 (N_1671,N_904,N_972);
xnor U1672 (N_1672,N_1460,N_887);
nand U1673 (N_1673,N_1468,N_1066);
nor U1674 (N_1674,N_1413,N_1151);
and U1675 (N_1675,N_1051,N_1228);
xnor U1676 (N_1676,N_1054,N_1310);
xnor U1677 (N_1677,N_1194,N_860);
nand U1678 (N_1678,N_1438,N_991);
or U1679 (N_1679,N_1269,N_1078);
and U1680 (N_1680,N_977,N_1111);
or U1681 (N_1681,N_1024,N_1435);
xnor U1682 (N_1682,N_878,N_794);
and U1683 (N_1683,N_1005,N_771);
nor U1684 (N_1684,N_1328,N_1313);
and U1685 (N_1685,N_1087,N_918);
and U1686 (N_1686,N_1434,N_1180);
xnor U1687 (N_1687,N_785,N_854);
nand U1688 (N_1688,N_1023,N_798);
xor U1689 (N_1689,N_1211,N_847);
nand U1690 (N_1690,N_1464,N_1327);
xor U1691 (N_1691,N_1304,N_1455);
and U1692 (N_1692,N_1359,N_1150);
and U1693 (N_1693,N_1110,N_950);
and U1694 (N_1694,N_851,N_1221);
nand U1695 (N_1695,N_1136,N_760);
xor U1696 (N_1696,N_1282,N_935);
xor U1697 (N_1697,N_862,N_1443);
nand U1698 (N_1698,N_1010,N_1113);
xor U1699 (N_1699,N_1174,N_1163);
nand U1700 (N_1700,N_1201,N_838);
xnor U1701 (N_1701,N_754,N_1069);
nand U1702 (N_1702,N_763,N_1404);
nand U1703 (N_1703,N_1185,N_1251);
and U1704 (N_1704,N_1480,N_1412);
nor U1705 (N_1705,N_1268,N_1350);
nor U1706 (N_1706,N_1036,N_1142);
or U1707 (N_1707,N_956,N_1383);
nand U1708 (N_1708,N_964,N_898);
nor U1709 (N_1709,N_1014,N_833);
or U1710 (N_1710,N_1244,N_1272);
xor U1711 (N_1711,N_986,N_1267);
and U1712 (N_1712,N_921,N_843);
nand U1713 (N_1713,N_1229,N_1230);
xnor U1714 (N_1714,N_1287,N_1466);
nand U1715 (N_1715,N_1055,N_1454);
or U1716 (N_1716,N_1467,N_1441);
and U1717 (N_1717,N_1131,N_1209);
nand U1718 (N_1718,N_1178,N_1415);
and U1719 (N_1719,N_1346,N_1092);
nor U1720 (N_1720,N_1223,N_1283);
nor U1721 (N_1721,N_775,N_1277);
xor U1722 (N_1722,N_1477,N_1393);
nand U1723 (N_1723,N_836,N_1102);
nor U1724 (N_1724,N_1195,N_965);
and U1725 (N_1725,N_1391,N_1316);
nor U1726 (N_1726,N_1452,N_1224);
or U1727 (N_1727,N_928,N_1007);
or U1728 (N_1728,N_751,N_1498);
nand U1729 (N_1729,N_1104,N_1336);
or U1730 (N_1730,N_770,N_750);
and U1731 (N_1731,N_1234,N_1309);
xnor U1732 (N_1732,N_936,N_1217);
or U1733 (N_1733,N_812,N_1232);
xor U1734 (N_1734,N_782,N_1371);
xnor U1735 (N_1735,N_1255,N_1020);
nand U1736 (N_1736,N_1250,N_1381);
and U1737 (N_1737,N_780,N_1038);
xnor U1738 (N_1738,N_1121,N_946);
xor U1739 (N_1739,N_1240,N_1158);
nand U1740 (N_1740,N_1403,N_1289);
nand U1741 (N_1741,N_1076,N_1073);
nor U1742 (N_1742,N_1107,N_1345);
or U1743 (N_1743,N_1344,N_981);
or U1744 (N_1744,N_1360,N_1175);
xnor U1745 (N_1745,N_861,N_1190);
and U1746 (N_1746,N_885,N_1453);
and U1747 (N_1747,N_778,N_955);
xor U1748 (N_1748,N_1171,N_1089);
or U1749 (N_1749,N_1119,N_1337);
nor U1750 (N_1750,N_1442,N_1486);
nor U1751 (N_1751,N_774,N_1249);
and U1752 (N_1752,N_971,N_1071);
and U1753 (N_1753,N_848,N_1275);
or U1754 (N_1754,N_1159,N_1294);
and U1755 (N_1755,N_962,N_1098);
nand U1756 (N_1756,N_1108,N_1193);
and U1757 (N_1757,N_1279,N_1259);
nand U1758 (N_1758,N_1093,N_809);
xor U1759 (N_1759,N_1256,N_1062);
nor U1760 (N_1760,N_880,N_960);
nor U1761 (N_1761,N_1293,N_1475);
nand U1762 (N_1762,N_1239,N_1012);
or U1763 (N_1763,N_1353,N_799);
nor U1764 (N_1764,N_869,N_1057);
xor U1765 (N_1765,N_975,N_959);
nand U1766 (N_1766,N_866,N_1018);
xor U1767 (N_1767,N_1059,N_927);
xor U1768 (N_1768,N_1080,N_1177);
xnor U1769 (N_1769,N_873,N_1366);
and U1770 (N_1770,N_815,N_1016);
and U1771 (N_1771,N_1273,N_1266);
nand U1772 (N_1772,N_1046,N_810);
or U1773 (N_1773,N_823,N_1189);
nand U1774 (N_1774,N_1047,N_1290);
nor U1775 (N_1775,N_837,N_1085);
and U1776 (N_1776,N_1164,N_1129);
nor U1777 (N_1777,N_1040,N_1254);
or U1778 (N_1778,N_1291,N_1430);
xnor U1779 (N_1779,N_1488,N_1056);
nor U1780 (N_1780,N_1065,N_1033);
and U1781 (N_1781,N_1074,N_1420);
nand U1782 (N_1782,N_1357,N_1409);
nand U1783 (N_1783,N_1426,N_894);
xnor U1784 (N_1784,N_1374,N_752);
or U1785 (N_1785,N_1398,N_1490);
or U1786 (N_1786,N_1144,N_1213);
xor U1787 (N_1787,N_1160,N_853);
nor U1788 (N_1788,N_1340,N_1031);
nor U1789 (N_1789,N_1122,N_1133);
nand U1790 (N_1790,N_916,N_1214);
and U1791 (N_1791,N_781,N_944);
nand U1792 (N_1792,N_792,N_993);
xnor U1793 (N_1793,N_1334,N_1375);
xnor U1794 (N_1794,N_865,N_1106);
or U1795 (N_1795,N_1208,N_1086);
or U1796 (N_1796,N_989,N_1487);
and U1797 (N_1797,N_963,N_933);
or U1798 (N_1798,N_1231,N_1118);
nor U1799 (N_1799,N_952,N_1284);
or U1800 (N_1800,N_902,N_1323);
or U1801 (N_1801,N_954,N_826);
xnor U1802 (N_1802,N_805,N_755);
nor U1803 (N_1803,N_1303,N_1227);
and U1804 (N_1804,N_1053,N_1352);
nand U1805 (N_1805,N_1001,N_768);
or U1806 (N_1806,N_757,N_908);
xnor U1807 (N_1807,N_900,N_1082);
or U1808 (N_1808,N_825,N_1463);
nand U1809 (N_1809,N_1172,N_1465);
nand U1810 (N_1810,N_1314,N_976);
nor U1811 (N_1811,N_919,N_892);
xor U1812 (N_1812,N_987,N_1301);
nor U1813 (N_1813,N_983,N_852);
nand U1814 (N_1814,N_1317,N_1300);
and U1815 (N_1815,N_1274,N_804);
xor U1816 (N_1816,N_886,N_984);
xnor U1817 (N_1817,N_924,N_1479);
or U1818 (N_1818,N_793,N_1114);
nor U1819 (N_1819,N_1134,N_769);
or U1820 (N_1820,N_1103,N_1141);
or U1821 (N_1821,N_953,N_1292);
or U1822 (N_1822,N_1469,N_1146);
nor U1823 (N_1823,N_806,N_800);
and U1824 (N_1824,N_1075,N_945);
and U1825 (N_1825,N_1032,N_1199);
nor U1826 (N_1826,N_758,N_1153);
or U1827 (N_1827,N_1297,N_979);
xnor U1828 (N_1828,N_884,N_1112);
nand U1829 (N_1829,N_890,N_905);
or U1830 (N_1830,N_899,N_1372);
and U1831 (N_1831,N_1433,N_1155);
nand U1832 (N_1832,N_846,N_857);
and U1833 (N_1833,N_1370,N_834);
nor U1834 (N_1834,N_914,N_1458);
nor U1835 (N_1835,N_1425,N_912);
or U1836 (N_1836,N_1157,N_807);
or U1837 (N_1837,N_827,N_1225);
and U1838 (N_1838,N_1436,N_1011);
xor U1839 (N_1839,N_1072,N_1263);
nand U1840 (N_1840,N_839,N_1414);
or U1841 (N_1841,N_1462,N_1029);
xnor U1842 (N_1842,N_1410,N_1183);
and U1843 (N_1843,N_1067,N_1042);
nand U1844 (N_1844,N_1440,N_756);
nor U1845 (N_1845,N_1343,N_1041);
and U1846 (N_1846,N_1242,N_907);
xor U1847 (N_1847,N_765,N_761);
nand U1848 (N_1848,N_753,N_1253);
and U1849 (N_1849,N_1126,N_925);
xor U1850 (N_1850,N_1482,N_1356);
nand U1851 (N_1851,N_1437,N_1392);
nand U1852 (N_1852,N_1128,N_762);
nor U1853 (N_1853,N_1219,N_1373);
xnor U1854 (N_1854,N_901,N_1473);
nand U1855 (N_1855,N_1257,N_1285);
nand U1856 (N_1856,N_889,N_1390);
and U1857 (N_1857,N_895,N_896);
nor U1858 (N_1858,N_1341,N_1405);
xor U1859 (N_1859,N_1068,N_1489);
nand U1860 (N_1860,N_947,N_767);
xor U1861 (N_1861,N_1376,N_1354);
or U1862 (N_1862,N_1281,N_969);
nor U1863 (N_1863,N_859,N_1173);
nand U1864 (N_1864,N_1168,N_829);
nand U1865 (N_1865,N_790,N_996);
nor U1866 (N_1866,N_797,N_1379);
or U1867 (N_1867,N_1483,N_1017);
and U1868 (N_1868,N_1143,N_1188);
or U1869 (N_1869,N_1123,N_1139);
and U1870 (N_1870,N_1369,N_1474);
or U1871 (N_1871,N_811,N_937);
xnor U1872 (N_1872,N_978,N_1034);
nand U1873 (N_1873,N_1210,N_1027);
xor U1874 (N_1874,N_1423,N_1206);
nand U1875 (N_1875,N_1070,N_1010);
or U1876 (N_1876,N_986,N_851);
and U1877 (N_1877,N_1253,N_1349);
xnor U1878 (N_1878,N_1061,N_1476);
and U1879 (N_1879,N_934,N_769);
or U1880 (N_1880,N_1194,N_1285);
or U1881 (N_1881,N_779,N_1270);
nand U1882 (N_1882,N_795,N_1303);
nor U1883 (N_1883,N_800,N_1344);
and U1884 (N_1884,N_1056,N_1220);
nand U1885 (N_1885,N_1140,N_870);
or U1886 (N_1886,N_1316,N_1064);
xnor U1887 (N_1887,N_916,N_843);
xnor U1888 (N_1888,N_781,N_766);
and U1889 (N_1889,N_1081,N_948);
xnor U1890 (N_1890,N_847,N_1349);
and U1891 (N_1891,N_961,N_1206);
nand U1892 (N_1892,N_1442,N_1006);
and U1893 (N_1893,N_980,N_1049);
nand U1894 (N_1894,N_754,N_955);
xnor U1895 (N_1895,N_1355,N_821);
or U1896 (N_1896,N_1152,N_843);
xnor U1897 (N_1897,N_1106,N_1277);
nor U1898 (N_1898,N_936,N_766);
nor U1899 (N_1899,N_1433,N_1005);
nor U1900 (N_1900,N_1460,N_1374);
and U1901 (N_1901,N_854,N_1337);
and U1902 (N_1902,N_969,N_1238);
nand U1903 (N_1903,N_1045,N_1307);
or U1904 (N_1904,N_838,N_1206);
or U1905 (N_1905,N_771,N_1377);
nor U1906 (N_1906,N_855,N_1189);
xor U1907 (N_1907,N_1485,N_1109);
nor U1908 (N_1908,N_851,N_1424);
nor U1909 (N_1909,N_1342,N_989);
nor U1910 (N_1910,N_866,N_1318);
nor U1911 (N_1911,N_1468,N_1373);
and U1912 (N_1912,N_781,N_979);
xnor U1913 (N_1913,N_939,N_1446);
or U1914 (N_1914,N_1133,N_1156);
or U1915 (N_1915,N_953,N_1394);
nand U1916 (N_1916,N_930,N_1017);
xor U1917 (N_1917,N_1097,N_914);
xnor U1918 (N_1918,N_1084,N_976);
nor U1919 (N_1919,N_869,N_1321);
nand U1920 (N_1920,N_1218,N_1487);
and U1921 (N_1921,N_1487,N_946);
nand U1922 (N_1922,N_760,N_848);
and U1923 (N_1923,N_916,N_1434);
nand U1924 (N_1924,N_1264,N_1358);
nand U1925 (N_1925,N_783,N_1220);
and U1926 (N_1926,N_1484,N_821);
or U1927 (N_1927,N_1224,N_1051);
or U1928 (N_1928,N_801,N_816);
and U1929 (N_1929,N_1302,N_1477);
nand U1930 (N_1930,N_1275,N_922);
nor U1931 (N_1931,N_1412,N_813);
nor U1932 (N_1932,N_1044,N_1360);
nand U1933 (N_1933,N_859,N_804);
and U1934 (N_1934,N_1168,N_1258);
xnor U1935 (N_1935,N_1211,N_817);
nor U1936 (N_1936,N_1407,N_831);
nand U1937 (N_1937,N_751,N_818);
and U1938 (N_1938,N_985,N_931);
nand U1939 (N_1939,N_1405,N_907);
and U1940 (N_1940,N_1169,N_897);
nor U1941 (N_1941,N_1140,N_1169);
or U1942 (N_1942,N_1286,N_1291);
nand U1943 (N_1943,N_861,N_1270);
xnor U1944 (N_1944,N_770,N_1401);
and U1945 (N_1945,N_1097,N_943);
xor U1946 (N_1946,N_1229,N_1143);
xor U1947 (N_1947,N_787,N_882);
nand U1948 (N_1948,N_1473,N_1187);
and U1949 (N_1949,N_848,N_1313);
or U1950 (N_1950,N_1231,N_927);
xnor U1951 (N_1951,N_1026,N_945);
or U1952 (N_1952,N_1260,N_1170);
and U1953 (N_1953,N_1033,N_1045);
xor U1954 (N_1954,N_1320,N_1195);
xnor U1955 (N_1955,N_1095,N_823);
nor U1956 (N_1956,N_1083,N_888);
and U1957 (N_1957,N_1053,N_961);
nand U1958 (N_1958,N_846,N_1474);
xnor U1959 (N_1959,N_1207,N_1051);
nor U1960 (N_1960,N_1390,N_1275);
nor U1961 (N_1961,N_794,N_1097);
xnor U1962 (N_1962,N_1301,N_1165);
and U1963 (N_1963,N_1307,N_1295);
nand U1964 (N_1964,N_1030,N_822);
nand U1965 (N_1965,N_1416,N_1126);
nand U1966 (N_1966,N_863,N_1262);
nor U1967 (N_1967,N_1488,N_1137);
or U1968 (N_1968,N_1180,N_1179);
nand U1969 (N_1969,N_1060,N_1365);
xnor U1970 (N_1970,N_932,N_858);
nand U1971 (N_1971,N_1206,N_928);
and U1972 (N_1972,N_1269,N_822);
nor U1973 (N_1973,N_1341,N_1186);
or U1974 (N_1974,N_812,N_1220);
nand U1975 (N_1975,N_1072,N_846);
or U1976 (N_1976,N_977,N_860);
xnor U1977 (N_1977,N_796,N_790);
and U1978 (N_1978,N_1230,N_1316);
nor U1979 (N_1979,N_1347,N_775);
xnor U1980 (N_1980,N_931,N_1247);
and U1981 (N_1981,N_1081,N_1370);
nand U1982 (N_1982,N_792,N_1492);
nor U1983 (N_1983,N_1133,N_867);
nand U1984 (N_1984,N_1361,N_1143);
nand U1985 (N_1985,N_1017,N_1488);
and U1986 (N_1986,N_774,N_1335);
and U1987 (N_1987,N_863,N_955);
xnor U1988 (N_1988,N_1447,N_1485);
nand U1989 (N_1989,N_1316,N_1485);
and U1990 (N_1990,N_1189,N_1066);
xor U1991 (N_1991,N_1133,N_1429);
nor U1992 (N_1992,N_870,N_1317);
nand U1993 (N_1993,N_998,N_978);
nor U1994 (N_1994,N_1151,N_886);
nor U1995 (N_1995,N_1398,N_802);
nand U1996 (N_1996,N_1009,N_1486);
xor U1997 (N_1997,N_1140,N_1101);
and U1998 (N_1998,N_1392,N_1110);
nor U1999 (N_1999,N_1330,N_1322);
nand U2000 (N_2000,N_1338,N_1047);
nand U2001 (N_2001,N_1037,N_1389);
nand U2002 (N_2002,N_797,N_1106);
and U2003 (N_2003,N_1046,N_999);
or U2004 (N_2004,N_1446,N_1106);
nor U2005 (N_2005,N_1358,N_1349);
nor U2006 (N_2006,N_1114,N_1302);
nor U2007 (N_2007,N_1310,N_787);
nand U2008 (N_2008,N_1228,N_1329);
xnor U2009 (N_2009,N_871,N_1368);
and U2010 (N_2010,N_821,N_1166);
xnor U2011 (N_2011,N_1027,N_810);
or U2012 (N_2012,N_1105,N_1392);
and U2013 (N_2013,N_1497,N_1070);
or U2014 (N_2014,N_828,N_1154);
nand U2015 (N_2015,N_1460,N_1084);
xnor U2016 (N_2016,N_1137,N_1293);
and U2017 (N_2017,N_938,N_1211);
nor U2018 (N_2018,N_1307,N_1217);
and U2019 (N_2019,N_963,N_1268);
nand U2020 (N_2020,N_1349,N_962);
or U2021 (N_2021,N_1131,N_909);
nor U2022 (N_2022,N_1444,N_1356);
nor U2023 (N_2023,N_775,N_1247);
nor U2024 (N_2024,N_1027,N_1236);
and U2025 (N_2025,N_785,N_923);
and U2026 (N_2026,N_808,N_903);
and U2027 (N_2027,N_1311,N_1449);
nand U2028 (N_2028,N_1348,N_983);
or U2029 (N_2029,N_1473,N_1076);
xnor U2030 (N_2030,N_1305,N_1282);
nand U2031 (N_2031,N_1444,N_1230);
xnor U2032 (N_2032,N_1146,N_1007);
nand U2033 (N_2033,N_815,N_796);
nand U2034 (N_2034,N_951,N_878);
xnor U2035 (N_2035,N_1193,N_885);
nand U2036 (N_2036,N_1119,N_1085);
nand U2037 (N_2037,N_1406,N_958);
xnor U2038 (N_2038,N_1221,N_1039);
nand U2039 (N_2039,N_1432,N_1062);
xnor U2040 (N_2040,N_1413,N_1068);
or U2041 (N_2041,N_1325,N_1369);
nor U2042 (N_2042,N_1441,N_1376);
xor U2043 (N_2043,N_1012,N_1351);
or U2044 (N_2044,N_1374,N_1434);
nand U2045 (N_2045,N_1341,N_1134);
and U2046 (N_2046,N_1423,N_1394);
or U2047 (N_2047,N_815,N_892);
and U2048 (N_2048,N_1478,N_1107);
and U2049 (N_2049,N_1024,N_1238);
and U2050 (N_2050,N_1157,N_767);
or U2051 (N_2051,N_1120,N_942);
xnor U2052 (N_2052,N_813,N_1406);
nor U2053 (N_2053,N_997,N_1439);
nand U2054 (N_2054,N_842,N_1474);
nand U2055 (N_2055,N_1308,N_1077);
or U2056 (N_2056,N_1068,N_982);
or U2057 (N_2057,N_1283,N_1472);
nor U2058 (N_2058,N_1387,N_1461);
and U2059 (N_2059,N_1304,N_837);
nor U2060 (N_2060,N_971,N_1132);
and U2061 (N_2061,N_1438,N_959);
nor U2062 (N_2062,N_1162,N_1434);
or U2063 (N_2063,N_1267,N_1181);
nor U2064 (N_2064,N_878,N_1179);
xor U2065 (N_2065,N_1165,N_752);
and U2066 (N_2066,N_1307,N_1123);
nor U2067 (N_2067,N_1253,N_1055);
nor U2068 (N_2068,N_1133,N_945);
nor U2069 (N_2069,N_1084,N_1076);
or U2070 (N_2070,N_1470,N_755);
nand U2071 (N_2071,N_1134,N_1392);
nor U2072 (N_2072,N_840,N_1389);
xor U2073 (N_2073,N_1163,N_1104);
nand U2074 (N_2074,N_1305,N_1067);
or U2075 (N_2075,N_1072,N_857);
nand U2076 (N_2076,N_1198,N_759);
and U2077 (N_2077,N_1423,N_1108);
nand U2078 (N_2078,N_1225,N_1098);
or U2079 (N_2079,N_1412,N_803);
nand U2080 (N_2080,N_1202,N_971);
or U2081 (N_2081,N_751,N_1113);
and U2082 (N_2082,N_949,N_951);
nor U2083 (N_2083,N_866,N_1329);
nand U2084 (N_2084,N_1106,N_1035);
nor U2085 (N_2085,N_783,N_1184);
or U2086 (N_2086,N_1157,N_780);
nor U2087 (N_2087,N_758,N_1038);
xor U2088 (N_2088,N_1050,N_925);
or U2089 (N_2089,N_1486,N_1220);
or U2090 (N_2090,N_1446,N_1033);
xnor U2091 (N_2091,N_1038,N_1369);
xnor U2092 (N_2092,N_1214,N_798);
or U2093 (N_2093,N_1437,N_1262);
and U2094 (N_2094,N_1209,N_1135);
nand U2095 (N_2095,N_1198,N_1263);
nand U2096 (N_2096,N_1195,N_1156);
nor U2097 (N_2097,N_1332,N_1349);
nand U2098 (N_2098,N_1380,N_791);
nor U2099 (N_2099,N_752,N_893);
xnor U2100 (N_2100,N_767,N_1429);
nor U2101 (N_2101,N_1314,N_1301);
nor U2102 (N_2102,N_964,N_845);
nand U2103 (N_2103,N_810,N_1471);
or U2104 (N_2104,N_762,N_819);
nor U2105 (N_2105,N_1022,N_1390);
nand U2106 (N_2106,N_1124,N_933);
xor U2107 (N_2107,N_1297,N_1291);
and U2108 (N_2108,N_1131,N_1290);
nor U2109 (N_2109,N_920,N_795);
xor U2110 (N_2110,N_1432,N_855);
nand U2111 (N_2111,N_766,N_1182);
nand U2112 (N_2112,N_1161,N_1311);
and U2113 (N_2113,N_1371,N_1498);
or U2114 (N_2114,N_817,N_1031);
or U2115 (N_2115,N_1170,N_1060);
or U2116 (N_2116,N_1340,N_1235);
nand U2117 (N_2117,N_1164,N_990);
nor U2118 (N_2118,N_1003,N_1353);
nor U2119 (N_2119,N_1438,N_940);
xnor U2120 (N_2120,N_1068,N_1234);
nor U2121 (N_2121,N_983,N_797);
or U2122 (N_2122,N_809,N_1406);
nor U2123 (N_2123,N_1311,N_1159);
or U2124 (N_2124,N_1409,N_958);
and U2125 (N_2125,N_897,N_1036);
xor U2126 (N_2126,N_1027,N_1479);
nand U2127 (N_2127,N_910,N_864);
and U2128 (N_2128,N_927,N_774);
xnor U2129 (N_2129,N_847,N_1161);
and U2130 (N_2130,N_795,N_986);
or U2131 (N_2131,N_960,N_799);
nor U2132 (N_2132,N_1342,N_1349);
or U2133 (N_2133,N_1276,N_1192);
or U2134 (N_2134,N_925,N_1363);
nor U2135 (N_2135,N_813,N_830);
nor U2136 (N_2136,N_1363,N_1268);
nor U2137 (N_2137,N_1452,N_1004);
nand U2138 (N_2138,N_758,N_1341);
or U2139 (N_2139,N_807,N_1103);
nand U2140 (N_2140,N_1253,N_1233);
or U2141 (N_2141,N_1035,N_982);
nor U2142 (N_2142,N_1343,N_868);
and U2143 (N_2143,N_981,N_1030);
xor U2144 (N_2144,N_869,N_1488);
nor U2145 (N_2145,N_1370,N_932);
nor U2146 (N_2146,N_992,N_1453);
nand U2147 (N_2147,N_936,N_1347);
and U2148 (N_2148,N_1021,N_1153);
xor U2149 (N_2149,N_844,N_971);
nand U2150 (N_2150,N_1158,N_894);
xnor U2151 (N_2151,N_1052,N_1458);
xor U2152 (N_2152,N_1206,N_1485);
xor U2153 (N_2153,N_1449,N_1370);
nand U2154 (N_2154,N_1454,N_886);
or U2155 (N_2155,N_1178,N_955);
or U2156 (N_2156,N_1057,N_1134);
or U2157 (N_2157,N_875,N_1140);
and U2158 (N_2158,N_1131,N_1154);
or U2159 (N_2159,N_837,N_1321);
nand U2160 (N_2160,N_984,N_1370);
and U2161 (N_2161,N_1096,N_1265);
nand U2162 (N_2162,N_1461,N_1122);
xnor U2163 (N_2163,N_916,N_866);
xnor U2164 (N_2164,N_850,N_1314);
and U2165 (N_2165,N_1230,N_1349);
and U2166 (N_2166,N_983,N_1276);
nor U2167 (N_2167,N_790,N_875);
nor U2168 (N_2168,N_857,N_913);
xnor U2169 (N_2169,N_1149,N_1346);
nor U2170 (N_2170,N_764,N_850);
nand U2171 (N_2171,N_1111,N_1023);
and U2172 (N_2172,N_1376,N_1124);
xnor U2173 (N_2173,N_852,N_764);
and U2174 (N_2174,N_1378,N_962);
nand U2175 (N_2175,N_1351,N_778);
or U2176 (N_2176,N_923,N_1442);
nor U2177 (N_2177,N_909,N_1166);
or U2178 (N_2178,N_804,N_1440);
and U2179 (N_2179,N_1377,N_1425);
and U2180 (N_2180,N_1292,N_965);
nand U2181 (N_2181,N_1155,N_1086);
and U2182 (N_2182,N_791,N_1170);
xnor U2183 (N_2183,N_1497,N_1313);
xnor U2184 (N_2184,N_825,N_1356);
nor U2185 (N_2185,N_1135,N_981);
or U2186 (N_2186,N_1162,N_1350);
xor U2187 (N_2187,N_1213,N_914);
or U2188 (N_2188,N_793,N_1117);
or U2189 (N_2189,N_1465,N_1203);
nand U2190 (N_2190,N_841,N_1499);
nor U2191 (N_2191,N_921,N_845);
nand U2192 (N_2192,N_866,N_1350);
nor U2193 (N_2193,N_1010,N_898);
xor U2194 (N_2194,N_1410,N_968);
or U2195 (N_2195,N_1116,N_922);
nand U2196 (N_2196,N_927,N_1293);
and U2197 (N_2197,N_968,N_1338);
nand U2198 (N_2198,N_1267,N_1240);
nor U2199 (N_2199,N_1034,N_1239);
nor U2200 (N_2200,N_965,N_794);
nor U2201 (N_2201,N_809,N_1058);
nor U2202 (N_2202,N_777,N_1227);
or U2203 (N_2203,N_798,N_1126);
and U2204 (N_2204,N_1367,N_858);
or U2205 (N_2205,N_955,N_1279);
nor U2206 (N_2206,N_1277,N_1394);
nor U2207 (N_2207,N_1076,N_819);
xor U2208 (N_2208,N_1148,N_1450);
nor U2209 (N_2209,N_1076,N_1269);
and U2210 (N_2210,N_1062,N_1153);
nor U2211 (N_2211,N_1152,N_960);
and U2212 (N_2212,N_883,N_844);
xor U2213 (N_2213,N_1361,N_1319);
nand U2214 (N_2214,N_1406,N_1409);
or U2215 (N_2215,N_949,N_1362);
nand U2216 (N_2216,N_1313,N_1374);
xor U2217 (N_2217,N_761,N_992);
and U2218 (N_2218,N_974,N_1305);
or U2219 (N_2219,N_920,N_1247);
or U2220 (N_2220,N_1102,N_1359);
xor U2221 (N_2221,N_993,N_1008);
nor U2222 (N_2222,N_1165,N_1357);
and U2223 (N_2223,N_949,N_1389);
nand U2224 (N_2224,N_932,N_1459);
xnor U2225 (N_2225,N_1029,N_1219);
nor U2226 (N_2226,N_943,N_1115);
or U2227 (N_2227,N_1406,N_934);
nor U2228 (N_2228,N_840,N_883);
nor U2229 (N_2229,N_771,N_1268);
and U2230 (N_2230,N_1216,N_777);
xor U2231 (N_2231,N_1068,N_1078);
nor U2232 (N_2232,N_1089,N_1418);
nand U2233 (N_2233,N_844,N_764);
and U2234 (N_2234,N_881,N_1356);
xor U2235 (N_2235,N_1102,N_1188);
and U2236 (N_2236,N_866,N_836);
nand U2237 (N_2237,N_839,N_932);
nor U2238 (N_2238,N_1255,N_997);
nor U2239 (N_2239,N_1055,N_1184);
or U2240 (N_2240,N_929,N_1471);
xor U2241 (N_2241,N_1476,N_1021);
xor U2242 (N_2242,N_797,N_1225);
or U2243 (N_2243,N_1440,N_1439);
nand U2244 (N_2244,N_1466,N_840);
xor U2245 (N_2245,N_1048,N_912);
or U2246 (N_2246,N_762,N_1162);
nor U2247 (N_2247,N_967,N_1173);
nand U2248 (N_2248,N_1404,N_1485);
xnor U2249 (N_2249,N_1341,N_1222);
or U2250 (N_2250,N_1577,N_1717);
or U2251 (N_2251,N_1672,N_2136);
or U2252 (N_2252,N_2100,N_1849);
or U2253 (N_2253,N_2220,N_1993);
or U2254 (N_2254,N_1893,N_1847);
nand U2255 (N_2255,N_2204,N_1851);
and U2256 (N_2256,N_1797,N_1733);
and U2257 (N_2257,N_1818,N_1828);
and U2258 (N_2258,N_1613,N_2201);
xor U2259 (N_2259,N_1933,N_1894);
xor U2260 (N_2260,N_1647,N_1583);
nand U2261 (N_2261,N_1830,N_1927);
nor U2262 (N_2262,N_1665,N_2000);
nand U2263 (N_2263,N_1860,N_2181);
nor U2264 (N_2264,N_2027,N_1579);
xor U2265 (N_2265,N_1926,N_1697);
nor U2266 (N_2266,N_1712,N_1671);
nand U2267 (N_2267,N_1663,N_2109);
nand U2268 (N_2268,N_1689,N_1758);
and U2269 (N_2269,N_2089,N_1941);
and U2270 (N_2270,N_1527,N_2036);
or U2271 (N_2271,N_1965,N_1901);
and U2272 (N_2272,N_1952,N_2126);
and U2273 (N_2273,N_2221,N_2055);
nor U2274 (N_2274,N_1884,N_1994);
nor U2275 (N_2275,N_1881,N_1617);
nand U2276 (N_2276,N_2169,N_1564);
xnor U2277 (N_2277,N_1516,N_2164);
xor U2278 (N_2278,N_1547,N_2131);
xor U2279 (N_2279,N_2014,N_2125);
or U2280 (N_2280,N_2080,N_1554);
nand U2281 (N_2281,N_2038,N_1968);
and U2282 (N_2282,N_2149,N_1509);
nor U2283 (N_2283,N_1925,N_1869);
or U2284 (N_2284,N_2033,N_2034);
nand U2285 (N_2285,N_2167,N_2042);
nor U2286 (N_2286,N_1838,N_1676);
or U2287 (N_2287,N_2016,N_1747);
and U2288 (N_2288,N_2240,N_1951);
xnor U2289 (N_2289,N_1619,N_1740);
nor U2290 (N_2290,N_1690,N_2105);
nand U2291 (N_2291,N_1726,N_1662);
nor U2292 (N_2292,N_1687,N_1789);
xor U2293 (N_2293,N_1624,N_2088);
nand U2294 (N_2294,N_1948,N_2123);
or U2295 (N_2295,N_2052,N_1693);
and U2296 (N_2296,N_2056,N_2077);
nand U2297 (N_2297,N_1678,N_2004);
and U2298 (N_2298,N_2205,N_1634);
nand U2299 (N_2299,N_1594,N_1856);
nand U2300 (N_2300,N_1908,N_1803);
xor U2301 (N_2301,N_1521,N_2176);
nand U2302 (N_2302,N_1599,N_1807);
nor U2303 (N_2303,N_1708,N_1783);
xnor U2304 (N_2304,N_2041,N_1653);
and U2305 (N_2305,N_1855,N_2020);
nor U2306 (N_2306,N_1819,N_1660);
nand U2307 (N_2307,N_2121,N_2009);
nand U2308 (N_2308,N_1916,N_1754);
or U2309 (N_2309,N_1764,N_2120);
and U2310 (N_2310,N_1798,N_1742);
nor U2311 (N_2311,N_2186,N_2231);
or U2312 (N_2312,N_1762,N_1722);
xor U2313 (N_2313,N_1749,N_2032);
and U2314 (N_2314,N_1787,N_1848);
and U2315 (N_2315,N_2170,N_2189);
or U2316 (N_2316,N_2141,N_1745);
and U2317 (N_2317,N_1863,N_2165);
or U2318 (N_2318,N_1767,N_2063);
nand U2319 (N_2319,N_1954,N_2104);
and U2320 (N_2320,N_2198,N_2081);
nand U2321 (N_2321,N_2107,N_2196);
nand U2322 (N_2322,N_1539,N_1889);
xor U2323 (N_2323,N_1610,N_1661);
nand U2324 (N_2324,N_1560,N_1861);
xor U2325 (N_2325,N_1667,N_1545);
xor U2326 (N_2326,N_1604,N_2015);
and U2327 (N_2327,N_1563,N_1729);
nand U2328 (N_2328,N_2192,N_1589);
and U2329 (N_2329,N_1595,N_1652);
or U2330 (N_2330,N_1804,N_2114);
and U2331 (N_2331,N_1942,N_1971);
nor U2332 (N_2332,N_1921,N_1966);
and U2333 (N_2333,N_2024,N_1845);
nand U2334 (N_2334,N_1643,N_1518);
nor U2335 (N_2335,N_1912,N_1780);
xor U2336 (N_2336,N_1898,N_2005);
nand U2337 (N_2337,N_1562,N_1650);
nand U2338 (N_2338,N_1530,N_2103);
and U2339 (N_2339,N_1775,N_2068);
nor U2340 (N_2340,N_1679,N_1826);
nand U2341 (N_2341,N_2151,N_2237);
or U2342 (N_2342,N_1788,N_1909);
xor U2343 (N_2343,N_2083,N_1580);
nor U2344 (N_2344,N_2101,N_1732);
nand U2345 (N_2345,N_2044,N_2249);
nand U2346 (N_2346,N_1628,N_1645);
and U2347 (N_2347,N_1738,N_2243);
or U2348 (N_2348,N_1872,N_1612);
or U2349 (N_2349,N_1769,N_1696);
xor U2350 (N_2350,N_2172,N_1811);
nand U2351 (N_2351,N_1753,N_1825);
and U2352 (N_2352,N_1963,N_1888);
nand U2353 (N_2353,N_2070,N_1873);
nand U2354 (N_2354,N_2146,N_1718);
and U2355 (N_2355,N_1915,N_1936);
nand U2356 (N_2356,N_1844,N_2049);
and U2357 (N_2357,N_1559,N_1770);
nand U2358 (N_2358,N_2145,N_1506);
nor U2359 (N_2359,N_2232,N_1649);
and U2360 (N_2360,N_1984,N_1555);
xnor U2361 (N_2361,N_1957,N_2174);
nor U2362 (N_2362,N_1786,N_2215);
nor U2363 (N_2363,N_1627,N_2021);
nand U2364 (N_2364,N_1953,N_2245);
nand U2365 (N_2365,N_1695,N_2122);
nand U2366 (N_2366,N_1836,N_1785);
or U2367 (N_2367,N_2029,N_1846);
nand U2368 (N_2368,N_2212,N_1685);
nand U2369 (N_2369,N_2244,N_1566);
and U2370 (N_2370,N_2072,N_1698);
nor U2371 (N_2371,N_1841,N_1934);
or U2372 (N_2372,N_1985,N_1501);
nand U2373 (N_2373,N_2013,N_1657);
xnor U2374 (N_2374,N_1977,N_1618);
nor U2375 (N_2375,N_1962,N_1939);
nor U2376 (N_2376,N_2143,N_1978);
nor U2377 (N_2377,N_1902,N_1537);
nor U2378 (N_2378,N_1937,N_1871);
nor U2379 (N_2379,N_2069,N_2202);
or U2380 (N_2380,N_1983,N_1546);
xnor U2381 (N_2381,N_1990,N_2085);
and U2382 (N_2382,N_2133,N_1969);
nand U2383 (N_2383,N_2054,N_1883);
nor U2384 (N_2384,N_1996,N_1731);
xnor U2385 (N_2385,N_1633,N_1588);
nand U2386 (N_2386,N_1741,N_2028);
xnor U2387 (N_2387,N_1887,N_1774);
nand U2388 (N_2388,N_1648,N_2175);
or U2389 (N_2389,N_2248,N_1569);
nor U2390 (N_2390,N_2045,N_2211);
xnor U2391 (N_2391,N_2019,N_1593);
and U2392 (N_2392,N_2190,N_2116);
nor U2393 (N_2393,N_1616,N_1552);
xor U2394 (N_2394,N_1701,N_1611);
or U2395 (N_2395,N_1799,N_1532);
nand U2396 (N_2396,N_1905,N_2193);
nand U2397 (N_2397,N_1814,N_1550);
xnor U2398 (N_2398,N_1958,N_2071);
nor U2399 (N_2399,N_1620,N_1556);
and U2400 (N_2400,N_1704,N_1714);
and U2401 (N_2401,N_2002,N_1919);
nand U2402 (N_2402,N_2227,N_2112);
nor U2403 (N_2403,N_1528,N_1680);
nor U2404 (N_2404,N_2007,N_1568);
nor U2405 (N_2405,N_1991,N_2037);
nand U2406 (N_2406,N_1922,N_1558);
or U2407 (N_2407,N_1561,N_1864);
xor U2408 (N_2408,N_1866,N_1614);
nand U2409 (N_2409,N_1531,N_2162);
nand U2410 (N_2410,N_1513,N_1763);
xnor U2411 (N_2411,N_2159,N_2209);
xnor U2412 (N_2412,N_2062,N_2207);
nor U2413 (N_2413,N_1734,N_2030);
and U2414 (N_2414,N_1791,N_1533);
nor U2415 (N_2415,N_1813,N_1808);
or U2416 (N_2416,N_2048,N_1673);
and U2417 (N_2417,N_2157,N_2006);
nor U2418 (N_2418,N_1706,N_1526);
xor U2419 (N_2419,N_1795,N_1536);
nand U2420 (N_2420,N_1756,N_2058);
and U2421 (N_2421,N_1820,N_1641);
nand U2422 (N_2422,N_1998,N_2241);
or U2423 (N_2423,N_2188,N_1903);
or U2424 (N_2424,N_2155,N_1683);
xnor U2425 (N_2425,N_2210,N_2066);
nor U2426 (N_2426,N_1575,N_1542);
nand U2427 (N_2427,N_1582,N_1636);
nand U2428 (N_2428,N_2091,N_2096);
nor U2429 (N_2429,N_1730,N_2092);
or U2430 (N_2430,N_1600,N_1668);
xor U2431 (N_2431,N_1572,N_1892);
or U2432 (N_2432,N_2082,N_2067);
nand U2433 (N_2433,N_1891,N_1674);
or U2434 (N_2434,N_2135,N_1739);
and U2435 (N_2435,N_1987,N_1615);
or U2436 (N_2436,N_1867,N_1874);
and U2437 (N_2437,N_1793,N_1543);
xnor U2438 (N_2438,N_1810,N_1534);
and U2439 (N_2439,N_1736,N_2074);
xnor U2440 (N_2440,N_2187,N_1629);
and U2441 (N_2441,N_1525,N_2213);
nor U2442 (N_2442,N_1659,N_1557);
nand U2443 (N_2443,N_1829,N_1761);
xor U2444 (N_2444,N_1549,N_2086);
nor U2445 (N_2445,N_1809,N_2173);
and U2446 (N_2446,N_1623,N_1517);
nor U2447 (N_2447,N_1602,N_2168);
or U2448 (N_2448,N_2191,N_2144);
or U2449 (N_2449,N_1920,N_2129);
xor U2450 (N_2450,N_2093,N_1520);
xor U2451 (N_2451,N_1802,N_2098);
xnor U2452 (N_2452,N_2226,N_1924);
nand U2453 (N_2453,N_1502,N_1637);
and U2454 (N_2454,N_1862,N_1827);
xor U2455 (N_2455,N_1776,N_2117);
and U2456 (N_2456,N_2017,N_1705);
or U2457 (N_2457,N_1551,N_2097);
and U2458 (N_2458,N_1938,N_1587);
and U2459 (N_2459,N_1821,N_1976);
and U2460 (N_2460,N_2147,N_1904);
or U2461 (N_2461,N_1682,N_1630);
xnor U2462 (N_2462,N_1765,N_2118);
nand U2463 (N_2463,N_1837,N_2040);
nor U2464 (N_2464,N_1956,N_1806);
nor U2465 (N_2465,N_2235,N_1694);
or U2466 (N_2466,N_1656,N_1932);
xnor U2467 (N_2467,N_1707,N_1515);
nor U2468 (N_2468,N_1720,N_1635);
nand U2469 (N_2469,N_1870,N_1975);
and U2470 (N_2470,N_1505,N_1815);
or U2471 (N_2471,N_1716,N_1523);
nor U2472 (N_2472,N_2043,N_1843);
xor U2473 (N_2473,N_1750,N_1522);
and U2474 (N_2474,N_1603,N_1607);
xor U2475 (N_2475,N_2156,N_2222);
or U2476 (N_2476,N_2184,N_2023);
nor U2477 (N_2477,N_2022,N_1597);
and U2478 (N_2478,N_1596,N_1725);
or U2479 (N_2479,N_1960,N_1746);
xnor U2480 (N_2480,N_1955,N_1824);
nand U2481 (N_2481,N_2199,N_1681);
and U2482 (N_2482,N_2078,N_2154);
xor U2483 (N_2483,N_2214,N_2064);
and U2484 (N_2484,N_1868,N_1833);
nand U2485 (N_2485,N_1743,N_1529);
xnor U2486 (N_2486,N_1713,N_1727);
nor U2487 (N_2487,N_1947,N_2229);
or U2488 (N_2488,N_1642,N_1839);
or U2489 (N_2489,N_1875,N_1688);
or U2490 (N_2490,N_1510,N_1974);
nor U2491 (N_2491,N_2084,N_1675);
xnor U2492 (N_2492,N_1606,N_1608);
xor U2493 (N_2493,N_2182,N_2206);
nor U2494 (N_2494,N_2179,N_1570);
xor U2495 (N_2495,N_2113,N_2150);
xnor U2496 (N_2496,N_1897,N_1748);
xor U2497 (N_2497,N_2242,N_1508);
nor U2498 (N_2498,N_1519,N_1778);
xor U2499 (N_2499,N_1914,N_2035);
xnor U2500 (N_2500,N_1900,N_1686);
nand U2501 (N_2501,N_1885,N_1930);
xor U2502 (N_2502,N_1639,N_1999);
nand U2503 (N_2503,N_1858,N_1541);
or U2504 (N_2504,N_2203,N_1711);
nor U2505 (N_2505,N_1638,N_1782);
nand U2506 (N_2506,N_1752,N_1598);
nor U2507 (N_2507,N_1514,N_1944);
and U2508 (N_2508,N_2180,N_1840);
nand U2509 (N_2509,N_2060,N_1800);
nand U2510 (N_2510,N_1805,N_1548);
nor U2511 (N_2511,N_1857,N_1771);
nand U2512 (N_2512,N_2010,N_1700);
or U2513 (N_2513,N_1970,N_1982);
xnor U2514 (N_2514,N_2234,N_1507);
or U2515 (N_2515,N_1773,N_2177);
xor U2516 (N_2516,N_1997,N_1512);
and U2517 (N_2517,N_1524,N_1801);
nand U2518 (N_2518,N_1654,N_2166);
nand U2519 (N_2519,N_1859,N_1832);
nor U2520 (N_2520,N_2178,N_1972);
and U2521 (N_2521,N_1876,N_1853);
nor U2522 (N_2522,N_2185,N_1565);
and U2523 (N_2523,N_2115,N_1699);
nand U2524 (N_2524,N_1735,N_1950);
nor U2525 (N_2525,N_2223,N_1586);
nand U2526 (N_2526,N_2090,N_1766);
xor U2527 (N_2527,N_1581,N_2246);
nor U2528 (N_2528,N_1906,N_2026);
xnor U2529 (N_2529,N_1590,N_2110);
and U2530 (N_2530,N_1723,N_1895);
nor U2531 (N_2531,N_2224,N_2219);
and U2532 (N_2532,N_2108,N_2160);
or U2533 (N_2533,N_2047,N_1834);
or U2534 (N_2534,N_2152,N_1923);
nor U2535 (N_2535,N_2200,N_1724);
nor U2536 (N_2536,N_1911,N_1751);
nand U2537 (N_2537,N_1842,N_1877);
nor U2538 (N_2538,N_1728,N_2217);
nand U2539 (N_2539,N_2142,N_1703);
nor U2540 (N_2540,N_1719,N_2132);
xnor U2541 (N_2541,N_2095,N_2171);
or U2542 (N_2542,N_2228,N_1677);
and U2543 (N_2543,N_1755,N_1979);
or U2544 (N_2544,N_2050,N_1910);
or U2545 (N_2545,N_1772,N_2138);
and U2546 (N_2546,N_1658,N_1784);
or U2547 (N_2547,N_2039,N_1980);
nor U2548 (N_2548,N_1666,N_1768);
nand U2549 (N_2549,N_1626,N_1640);
nand U2550 (N_2550,N_2161,N_2127);
or U2551 (N_2551,N_2025,N_1621);
nand U2552 (N_2552,N_1757,N_2008);
xor U2553 (N_2553,N_1812,N_2247);
xor U2554 (N_2554,N_2094,N_1721);
or U2555 (N_2555,N_2239,N_1831);
and U2556 (N_2556,N_2075,N_1651);
and U2557 (N_2557,N_1779,N_2111);
or U2558 (N_2558,N_2031,N_2183);
xor U2559 (N_2559,N_1571,N_2130);
nand U2560 (N_2560,N_1882,N_1794);
or U2561 (N_2561,N_1880,N_2225);
or U2562 (N_2562,N_1967,N_1670);
or U2563 (N_2563,N_2195,N_1777);
xor U2564 (N_2564,N_1973,N_1544);
nor U2565 (N_2565,N_2139,N_1578);
or U2566 (N_2566,N_1709,N_2046);
nor U2567 (N_2567,N_1609,N_1959);
and U2568 (N_2568,N_1929,N_1540);
and U2569 (N_2569,N_2087,N_1760);
nand U2570 (N_2570,N_2124,N_2140);
and U2571 (N_2571,N_2119,N_1865);
nor U2572 (N_2572,N_1790,N_1796);
xor U2573 (N_2573,N_1913,N_1822);
and U2574 (N_2574,N_1943,N_1792);
nand U2575 (N_2575,N_1744,N_2194);
or U2576 (N_2576,N_1928,N_1655);
or U2577 (N_2577,N_1935,N_2061);
nor U2578 (N_2578,N_1946,N_1759);
or U2579 (N_2579,N_2148,N_1945);
nor U2580 (N_2580,N_2153,N_2208);
or U2581 (N_2581,N_1574,N_1644);
nand U2582 (N_2582,N_2099,N_1500);
and U2583 (N_2583,N_2057,N_1878);
xor U2584 (N_2584,N_1622,N_1890);
and U2585 (N_2585,N_1992,N_1737);
or U2586 (N_2586,N_2233,N_1835);
nand U2587 (N_2587,N_2158,N_2079);
and U2588 (N_2588,N_1692,N_2053);
nand U2589 (N_2589,N_1646,N_1504);
nor U2590 (N_2590,N_1605,N_1918);
nand U2591 (N_2591,N_1879,N_2065);
or U2592 (N_2592,N_1632,N_1989);
or U2593 (N_2593,N_1669,N_1535);
xor U2594 (N_2594,N_1823,N_2128);
or U2595 (N_2595,N_1592,N_1931);
nor U2596 (N_2596,N_1852,N_2001);
nor U2597 (N_2597,N_2137,N_1511);
and U2598 (N_2598,N_2230,N_1567);
nand U2599 (N_2599,N_2218,N_1986);
and U2600 (N_2600,N_1684,N_1917);
nor U2601 (N_2601,N_1854,N_2011);
nor U2602 (N_2602,N_2197,N_1601);
xor U2603 (N_2603,N_2216,N_1995);
nand U2604 (N_2604,N_1584,N_1816);
nand U2605 (N_2605,N_1538,N_2102);
nor U2606 (N_2606,N_1702,N_2059);
and U2607 (N_2607,N_2051,N_1886);
nand U2608 (N_2608,N_1691,N_1907);
nor U2609 (N_2609,N_1591,N_1817);
or U2610 (N_2610,N_2018,N_1553);
nand U2611 (N_2611,N_1631,N_2134);
nor U2612 (N_2612,N_1981,N_1503);
nand U2613 (N_2613,N_1664,N_1710);
nor U2614 (N_2614,N_1949,N_1585);
xor U2615 (N_2615,N_1988,N_2003);
or U2616 (N_2616,N_1940,N_1961);
or U2617 (N_2617,N_2106,N_1715);
and U2618 (N_2618,N_2076,N_1576);
nor U2619 (N_2619,N_1850,N_1896);
nand U2620 (N_2620,N_2238,N_1964);
nor U2621 (N_2621,N_1573,N_2073);
nor U2622 (N_2622,N_2236,N_2012);
or U2623 (N_2623,N_1781,N_1625);
nand U2624 (N_2624,N_2163,N_1899);
or U2625 (N_2625,N_1715,N_2185);
nand U2626 (N_2626,N_1866,N_1961);
and U2627 (N_2627,N_2112,N_1721);
or U2628 (N_2628,N_1545,N_1994);
nor U2629 (N_2629,N_1557,N_1578);
nand U2630 (N_2630,N_1850,N_1842);
xnor U2631 (N_2631,N_2069,N_1725);
nand U2632 (N_2632,N_2200,N_2215);
or U2633 (N_2633,N_1749,N_1907);
or U2634 (N_2634,N_2152,N_1506);
nand U2635 (N_2635,N_1957,N_1931);
nand U2636 (N_2636,N_1955,N_2189);
xor U2637 (N_2637,N_2073,N_2126);
or U2638 (N_2638,N_1633,N_2068);
xnor U2639 (N_2639,N_2069,N_1930);
or U2640 (N_2640,N_1947,N_1728);
xor U2641 (N_2641,N_1893,N_1786);
nor U2642 (N_2642,N_1807,N_2038);
or U2643 (N_2643,N_1864,N_2222);
nand U2644 (N_2644,N_2023,N_1860);
and U2645 (N_2645,N_2181,N_1660);
nand U2646 (N_2646,N_1783,N_1897);
or U2647 (N_2647,N_1851,N_1980);
or U2648 (N_2648,N_1556,N_1937);
and U2649 (N_2649,N_1873,N_1759);
nand U2650 (N_2650,N_1512,N_2147);
xor U2651 (N_2651,N_1679,N_1756);
or U2652 (N_2652,N_1746,N_2054);
and U2653 (N_2653,N_1818,N_1829);
nor U2654 (N_2654,N_2202,N_1508);
or U2655 (N_2655,N_2110,N_1876);
nand U2656 (N_2656,N_1541,N_1667);
nor U2657 (N_2657,N_2157,N_2083);
and U2658 (N_2658,N_2245,N_2206);
nand U2659 (N_2659,N_2065,N_2246);
nand U2660 (N_2660,N_1702,N_1705);
nand U2661 (N_2661,N_1533,N_1749);
nor U2662 (N_2662,N_1521,N_1624);
xnor U2663 (N_2663,N_2117,N_1681);
and U2664 (N_2664,N_2167,N_2016);
and U2665 (N_2665,N_2061,N_2230);
xnor U2666 (N_2666,N_2161,N_2131);
nor U2667 (N_2667,N_1551,N_2036);
nor U2668 (N_2668,N_1620,N_1588);
xnor U2669 (N_2669,N_2245,N_2110);
and U2670 (N_2670,N_2231,N_1618);
nor U2671 (N_2671,N_1577,N_2138);
nor U2672 (N_2672,N_2226,N_1899);
xor U2673 (N_2673,N_1902,N_1662);
nor U2674 (N_2674,N_2040,N_1523);
xnor U2675 (N_2675,N_1560,N_1733);
xor U2676 (N_2676,N_1648,N_2075);
xor U2677 (N_2677,N_2110,N_1920);
nand U2678 (N_2678,N_1852,N_2102);
and U2679 (N_2679,N_1579,N_1598);
xor U2680 (N_2680,N_1711,N_1576);
nand U2681 (N_2681,N_1856,N_2202);
xnor U2682 (N_2682,N_2062,N_2053);
xor U2683 (N_2683,N_1531,N_1737);
or U2684 (N_2684,N_1559,N_1551);
nor U2685 (N_2685,N_2187,N_1569);
nor U2686 (N_2686,N_2089,N_1990);
nor U2687 (N_2687,N_2232,N_2211);
nor U2688 (N_2688,N_1519,N_2175);
xnor U2689 (N_2689,N_1516,N_1841);
or U2690 (N_2690,N_1763,N_2038);
or U2691 (N_2691,N_1659,N_2112);
xor U2692 (N_2692,N_1500,N_2112);
nand U2693 (N_2693,N_1853,N_2179);
and U2694 (N_2694,N_1806,N_2166);
nor U2695 (N_2695,N_1952,N_1663);
nand U2696 (N_2696,N_1985,N_1597);
or U2697 (N_2697,N_2002,N_2229);
or U2698 (N_2698,N_1593,N_1863);
nand U2699 (N_2699,N_1930,N_1840);
nand U2700 (N_2700,N_1967,N_2109);
nand U2701 (N_2701,N_1839,N_1771);
nor U2702 (N_2702,N_1582,N_1771);
xor U2703 (N_2703,N_2021,N_2221);
xnor U2704 (N_2704,N_2069,N_1516);
xnor U2705 (N_2705,N_1592,N_1824);
nor U2706 (N_2706,N_2080,N_2088);
nand U2707 (N_2707,N_1779,N_1589);
nor U2708 (N_2708,N_1856,N_2101);
or U2709 (N_2709,N_1914,N_1798);
or U2710 (N_2710,N_1844,N_1744);
or U2711 (N_2711,N_1842,N_1635);
or U2712 (N_2712,N_2069,N_1783);
or U2713 (N_2713,N_1542,N_1768);
and U2714 (N_2714,N_1788,N_2118);
nor U2715 (N_2715,N_2144,N_1813);
or U2716 (N_2716,N_1802,N_2099);
xnor U2717 (N_2717,N_1541,N_2053);
xor U2718 (N_2718,N_1866,N_2047);
or U2719 (N_2719,N_2237,N_1863);
xnor U2720 (N_2720,N_2075,N_2088);
or U2721 (N_2721,N_2249,N_2222);
or U2722 (N_2722,N_2242,N_2248);
or U2723 (N_2723,N_1865,N_1799);
and U2724 (N_2724,N_1752,N_1764);
and U2725 (N_2725,N_2249,N_1523);
xnor U2726 (N_2726,N_2124,N_1691);
or U2727 (N_2727,N_1808,N_1912);
nor U2728 (N_2728,N_2210,N_1837);
or U2729 (N_2729,N_1699,N_2197);
or U2730 (N_2730,N_1561,N_1511);
or U2731 (N_2731,N_2089,N_2046);
nand U2732 (N_2732,N_1778,N_1958);
nand U2733 (N_2733,N_2023,N_1689);
nor U2734 (N_2734,N_2148,N_2061);
and U2735 (N_2735,N_1907,N_1710);
or U2736 (N_2736,N_1579,N_2144);
xnor U2737 (N_2737,N_1919,N_1855);
and U2738 (N_2738,N_2234,N_2149);
xnor U2739 (N_2739,N_2171,N_2118);
or U2740 (N_2740,N_1864,N_2243);
nor U2741 (N_2741,N_2091,N_1616);
or U2742 (N_2742,N_1752,N_1820);
xnor U2743 (N_2743,N_2196,N_1932);
and U2744 (N_2744,N_1822,N_1582);
nor U2745 (N_2745,N_1812,N_1935);
or U2746 (N_2746,N_1963,N_1921);
and U2747 (N_2747,N_1850,N_1653);
or U2748 (N_2748,N_1685,N_1697);
nor U2749 (N_2749,N_1560,N_2056);
and U2750 (N_2750,N_2199,N_2158);
xor U2751 (N_2751,N_1509,N_1539);
or U2752 (N_2752,N_2015,N_1944);
and U2753 (N_2753,N_1723,N_2074);
nor U2754 (N_2754,N_2097,N_2080);
nor U2755 (N_2755,N_2184,N_1788);
or U2756 (N_2756,N_1943,N_1996);
nand U2757 (N_2757,N_1591,N_1548);
nor U2758 (N_2758,N_2000,N_2021);
nand U2759 (N_2759,N_2103,N_2191);
and U2760 (N_2760,N_1551,N_1754);
and U2761 (N_2761,N_1950,N_1990);
and U2762 (N_2762,N_1732,N_1538);
nor U2763 (N_2763,N_2130,N_1878);
nor U2764 (N_2764,N_1528,N_2184);
nor U2765 (N_2765,N_1701,N_2079);
xor U2766 (N_2766,N_2119,N_2087);
and U2767 (N_2767,N_1777,N_1519);
or U2768 (N_2768,N_2186,N_2046);
nor U2769 (N_2769,N_1854,N_1936);
xnor U2770 (N_2770,N_1733,N_2221);
nor U2771 (N_2771,N_2004,N_2084);
nand U2772 (N_2772,N_1752,N_1934);
nor U2773 (N_2773,N_2046,N_1956);
and U2774 (N_2774,N_2138,N_1515);
nor U2775 (N_2775,N_2147,N_2246);
xor U2776 (N_2776,N_2132,N_1912);
and U2777 (N_2777,N_1619,N_2028);
and U2778 (N_2778,N_1507,N_2137);
nor U2779 (N_2779,N_1992,N_1958);
nor U2780 (N_2780,N_1860,N_1735);
xnor U2781 (N_2781,N_1985,N_1837);
xor U2782 (N_2782,N_1966,N_1865);
nand U2783 (N_2783,N_1919,N_2100);
xor U2784 (N_2784,N_1643,N_1578);
nor U2785 (N_2785,N_1663,N_1706);
and U2786 (N_2786,N_1634,N_1667);
nor U2787 (N_2787,N_1622,N_1742);
nand U2788 (N_2788,N_1943,N_1604);
xnor U2789 (N_2789,N_1515,N_2234);
xnor U2790 (N_2790,N_1564,N_1561);
nand U2791 (N_2791,N_1844,N_1680);
and U2792 (N_2792,N_1554,N_1890);
nor U2793 (N_2793,N_2157,N_2123);
nor U2794 (N_2794,N_2032,N_2000);
nor U2795 (N_2795,N_1968,N_2129);
nand U2796 (N_2796,N_1779,N_1612);
xnor U2797 (N_2797,N_1836,N_1755);
nor U2798 (N_2798,N_1611,N_1503);
nor U2799 (N_2799,N_1652,N_2168);
nand U2800 (N_2800,N_1695,N_2064);
xor U2801 (N_2801,N_1989,N_2127);
and U2802 (N_2802,N_2180,N_1751);
xor U2803 (N_2803,N_2162,N_1948);
nand U2804 (N_2804,N_1791,N_1870);
and U2805 (N_2805,N_1527,N_1855);
xnor U2806 (N_2806,N_1783,N_1540);
xor U2807 (N_2807,N_2030,N_1716);
nand U2808 (N_2808,N_1517,N_1896);
xnor U2809 (N_2809,N_2183,N_2243);
and U2810 (N_2810,N_2085,N_2073);
and U2811 (N_2811,N_1500,N_1832);
nor U2812 (N_2812,N_1764,N_1584);
nor U2813 (N_2813,N_1515,N_1834);
nand U2814 (N_2814,N_1503,N_1523);
nand U2815 (N_2815,N_1932,N_2079);
or U2816 (N_2816,N_1506,N_2130);
nor U2817 (N_2817,N_1923,N_1507);
or U2818 (N_2818,N_1671,N_1888);
nand U2819 (N_2819,N_2031,N_1601);
nor U2820 (N_2820,N_1766,N_1820);
and U2821 (N_2821,N_2163,N_2223);
and U2822 (N_2822,N_2223,N_1594);
nand U2823 (N_2823,N_1765,N_1812);
nor U2824 (N_2824,N_1821,N_2051);
xnor U2825 (N_2825,N_1954,N_2087);
and U2826 (N_2826,N_2228,N_2215);
nand U2827 (N_2827,N_1692,N_1922);
xnor U2828 (N_2828,N_1834,N_2179);
or U2829 (N_2829,N_1614,N_2051);
and U2830 (N_2830,N_2204,N_2078);
or U2831 (N_2831,N_1516,N_2009);
xor U2832 (N_2832,N_1951,N_1849);
nor U2833 (N_2833,N_1578,N_1574);
or U2834 (N_2834,N_1824,N_2036);
nand U2835 (N_2835,N_1597,N_1996);
nand U2836 (N_2836,N_1920,N_2050);
nor U2837 (N_2837,N_1651,N_2064);
and U2838 (N_2838,N_1531,N_1635);
nand U2839 (N_2839,N_1792,N_2162);
nand U2840 (N_2840,N_2206,N_2117);
nand U2841 (N_2841,N_1953,N_1899);
and U2842 (N_2842,N_2097,N_1687);
xnor U2843 (N_2843,N_1745,N_2071);
or U2844 (N_2844,N_1988,N_1587);
nand U2845 (N_2845,N_1718,N_1797);
xnor U2846 (N_2846,N_1650,N_1529);
nor U2847 (N_2847,N_1514,N_1528);
nor U2848 (N_2848,N_1697,N_1701);
or U2849 (N_2849,N_2218,N_1808);
or U2850 (N_2850,N_1783,N_1664);
or U2851 (N_2851,N_1510,N_2069);
nor U2852 (N_2852,N_2013,N_1640);
and U2853 (N_2853,N_2100,N_1727);
nor U2854 (N_2854,N_1849,N_2189);
and U2855 (N_2855,N_1824,N_1975);
or U2856 (N_2856,N_1900,N_1575);
nand U2857 (N_2857,N_1599,N_1977);
xor U2858 (N_2858,N_1746,N_1636);
xnor U2859 (N_2859,N_1782,N_1748);
xor U2860 (N_2860,N_1912,N_1821);
nor U2861 (N_2861,N_1627,N_2202);
and U2862 (N_2862,N_2156,N_1906);
xor U2863 (N_2863,N_1883,N_2066);
or U2864 (N_2864,N_1562,N_1987);
nor U2865 (N_2865,N_2213,N_1835);
or U2866 (N_2866,N_2206,N_1593);
xnor U2867 (N_2867,N_1955,N_2239);
nor U2868 (N_2868,N_1969,N_2032);
nand U2869 (N_2869,N_1585,N_1713);
xnor U2870 (N_2870,N_1578,N_1938);
or U2871 (N_2871,N_2172,N_1915);
nand U2872 (N_2872,N_1621,N_1821);
nand U2873 (N_2873,N_1955,N_2120);
xor U2874 (N_2874,N_1629,N_1782);
and U2875 (N_2875,N_2194,N_1951);
nor U2876 (N_2876,N_1665,N_1655);
nand U2877 (N_2877,N_2067,N_2077);
and U2878 (N_2878,N_2146,N_2203);
and U2879 (N_2879,N_2119,N_1544);
or U2880 (N_2880,N_1626,N_2183);
or U2881 (N_2881,N_2059,N_1833);
nor U2882 (N_2882,N_1683,N_2087);
or U2883 (N_2883,N_1680,N_1882);
or U2884 (N_2884,N_2136,N_1898);
or U2885 (N_2885,N_2218,N_1970);
xor U2886 (N_2886,N_1555,N_2078);
nand U2887 (N_2887,N_2220,N_1922);
and U2888 (N_2888,N_2041,N_1659);
xnor U2889 (N_2889,N_2016,N_2147);
nand U2890 (N_2890,N_2223,N_1779);
xor U2891 (N_2891,N_1629,N_1586);
or U2892 (N_2892,N_1546,N_1621);
or U2893 (N_2893,N_1806,N_2096);
and U2894 (N_2894,N_1894,N_2184);
xor U2895 (N_2895,N_2211,N_1993);
or U2896 (N_2896,N_1752,N_1867);
nor U2897 (N_2897,N_2234,N_1504);
nand U2898 (N_2898,N_1935,N_1677);
and U2899 (N_2899,N_1683,N_2226);
and U2900 (N_2900,N_2195,N_1593);
and U2901 (N_2901,N_1936,N_1794);
or U2902 (N_2902,N_2097,N_1509);
nor U2903 (N_2903,N_1923,N_1652);
nand U2904 (N_2904,N_2214,N_1511);
nor U2905 (N_2905,N_2208,N_1947);
nand U2906 (N_2906,N_1612,N_2019);
nor U2907 (N_2907,N_1560,N_1741);
or U2908 (N_2908,N_1539,N_1541);
and U2909 (N_2909,N_1958,N_1776);
and U2910 (N_2910,N_2126,N_2034);
xor U2911 (N_2911,N_1948,N_1783);
or U2912 (N_2912,N_2165,N_1944);
nor U2913 (N_2913,N_2208,N_1625);
or U2914 (N_2914,N_2152,N_2027);
nor U2915 (N_2915,N_2062,N_1564);
nor U2916 (N_2916,N_1923,N_1525);
nand U2917 (N_2917,N_1840,N_2117);
and U2918 (N_2918,N_1963,N_1973);
and U2919 (N_2919,N_1939,N_1977);
nor U2920 (N_2920,N_1552,N_2124);
and U2921 (N_2921,N_1713,N_2110);
and U2922 (N_2922,N_1986,N_1837);
nor U2923 (N_2923,N_2104,N_1623);
nor U2924 (N_2924,N_1896,N_1875);
or U2925 (N_2925,N_2135,N_1975);
nor U2926 (N_2926,N_1949,N_2113);
nand U2927 (N_2927,N_1987,N_1714);
or U2928 (N_2928,N_1711,N_1740);
nand U2929 (N_2929,N_1607,N_1535);
xnor U2930 (N_2930,N_1787,N_1551);
or U2931 (N_2931,N_2163,N_1974);
nor U2932 (N_2932,N_2074,N_1824);
nor U2933 (N_2933,N_2127,N_1688);
and U2934 (N_2934,N_1878,N_2035);
or U2935 (N_2935,N_1990,N_1571);
and U2936 (N_2936,N_2086,N_1885);
nor U2937 (N_2937,N_1979,N_1577);
and U2938 (N_2938,N_1747,N_1992);
nand U2939 (N_2939,N_1767,N_1936);
xor U2940 (N_2940,N_2243,N_1724);
xnor U2941 (N_2941,N_1807,N_2158);
nor U2942 (N_2942,N_2218,N_1950);
xnor U2943 (N_2943,N_1999,N_1857);
or U2944 (N_2944,N_2074,N_2013);
xnor U2945 (N_2945,N_1843,N_1883);
and U2946 (N_2946,N_1869,N_1646);
and U2947 (N_2947,N_2068,N_1845);
xnor U2948 (N_2948,N_1664,N_2195);
xor U2949 (N_2949,N_2004,N_1513);
xnor U2950 (N_2950,N_2196,N_2243);
nand U2951 (N_2951,N_2021,N_2216);
xor U2952 (N_2952,N_2154,N_1717);
nor U2953 (N_2953,N_1684,N_2155);
nand U2954 (N_2954,N_2097,N_2070);
xor U2955 (N_2955,N_1980,N_2036);
or U2956 (N_2956,N_1686,N_1731);
and U2957 (N_2957,N_1627,N_2189);
xor U2958 (N_2958,N_1598,N_2048);
nor U2959 (N_2959,N_1723,N_2131);
or U2960 (N_2960,N_2189,N_1777);
or U2961 (N_2961,N_1993,N_1667);
and U2962 (N_2962,N_1895,N_2224);
nor U2963 (N_2963,N_1591,N_1988);
xnor U2964 (N_2964,N_1673,N_1638);
nand U2965 (N_2965,N_2160,N_1729);
and U2966 (N_2966,N_1571,N_2006);
nor U2967 (N_2967,N_1961,N_1935);
nand U2968 (N_2968,N_1770,N_1531);
nand U2969 (N_2969,N_1785,N_2011);
and U2970 (N_2970,N_1661,N_1564);
and U2971 (N_2971,N_1875,N_2085);
nor U2972 (N_2972,N_1560,N_2176);
nor U2973 (N_2973,N_1570,N_1746);
nand U2974 (N_2974,N_1947,N_1906);
and U2975 (N_2975,N_1801,N_2202);
and U2976 (N_2976,N_1976,N_1550);
nand U2977 (N_2977,N_2029,N_2022);
nor U2978 (N_2978,N_1528,N_2036);
xor U2979 (N_2979,N_2137,N_1803);
xnor U2980 (N_2980,N_1911,N_1864);
nand U2981 (N_2981,N_1500,N_1600);
and U2982 (N_2982,N_1769,N_1580);
nor U2983 (N_2983,N_2113,N_1945);
and U2984 (N_2984,N_1710,N_1866);
or U2985 (N_2985,N_1962,N_2155);
nand U2986 (N_2986,N_1854,N_1728);
nor U2987 (N_2987,N_1687,N_1856);
nor U2988 (N_2988,N_1850,N_2133);
nor U2989 (N_2989,N_1529,N_1623);
or U2990 (N_2990,N_1666,N_1806);
or U2991 (N_2991,N_1951,N_2210);
or U2992 (N_2992,N_2242,N_1610);
nor U2993 (N_2993,N_2144,N_1818);
or U2994 (N_2994,N_1931,N_1842);
or U2995 (N_2995,N_1980,N_1708);
nor U2996 (N_2996,N_1671,N_1709);
and U2997 (N_2997,N_1833,N_2228);
and U2998 (N_2998,N_1980,N_1752);
xnor U2999 (N_2999,N_1908,N_1624);
or UO_0 (O_0,N_2925,N_2488);
and UO_1 (O_1,N_2593,N_2835);
and UO_2 (O_2,N_2923,N_2381);
or UO_3 (O_3,N_2967,N_2714);
nand UO_4 (O_4,N_2599,N_2755);
and UO_5 (O_5,N_2857,N_2694);
and UO_6 (O_6,N_2756,N_2358);
nand UO_7 (O_7,N_2252,N_2870);
and UO_8 (O_8,N_2421,N_2760);
and UO_9 (O_9,N_2422,N_2389);
nor UO_10 (O_10,N_2569,N_2695);
nor UO_11 (O_11,N_2973,N_2785);
xnor UO_12 (O_12,N_2879,N_2312);
or UO_13 (O_13,N_2899,N_2414);
or UO_14 (O_14,N_2662,N_2439);
nand UO_15 (O_15,N_2462,N_2922);
or UO_16 (O_16,N_2814,N_2385);
or UO_17 (O_17,N_2465,N_2473);
nand UO_18 (O_18,N_2393,N_2304);
xnor UO_19 (O_19,N_2992,N_2951);
xor UO_20 (O_20,N_2515,N_2768);
or UO_21 (O_21,N_2797,N_2657);
or UO_22 (O_22,N_2485,N_2608);
and UO_23 (O_23,N_2444,N_2952);
or UO_24 (O_24,N_2826,N_2280);
or UO_25 (O_25,N_2668,N_2748);
nor UO_26 (O_26,N_2821,N_2484);
xor UO_27 (O_27,N_2666,N_2711);
or UO_28 (O_28,N_2977,N_2430);
or UO_29 (O_29,N_2782,N_2710);
or UO_30 (O_30,N_2661,N_2908);
or UO_31 (O_31,N_2638,N_2436);
xor UO_32 (O_32,N_2452,N_2536);
and UO_33 (O_33,N_2830,N_2631);
and UO_34 (O_34,N_2397,N_2704);
nand UO_35 (O_35,N_2734,N_2867);
or UO_36 (O_36,N_2617,N_2621);
nand UO_37 (O_37,N_2596,N_2565);
nor UO_38 (O_38,N_2969,N_2732);
nor UO_39 (O_39,N_2915,N_2772);
and UO_40 (O_40,N_2776,N_2813);
or UO_41 (O_41,N_2490,N_2965);
xnor UO_42 (O_42,N_2623,N_2349);
or UO_43 (O_43,N_2309,N_2635);
nand UO_44 (O_44,N_2298,N_2602);
and UO_45 (O_45,N_2663,N_2636);
or UO_46 (O_46,N_2698,N_2978);
xnor UO_47 (O_47,N_2427,N_2767);
nor UO_48 (O_48,N_2649,N_2726);
or UO_49 (O_49,N_2472,N_2268);
and UO_50 (O_50,N_2700,N_2853);
and UO_51 (O_51,N_2927,N_2983);
or UO_52 (O_52,N_2913,N_2939);
or UO_53 (O_53,N_2722,N_2543);
nand UO_54 (O_54,N_2463,N_2297);
and UO_55 (O_55,N_2750,N_2671);
or UO_56 (O_56,N_2934,N_2262);
and UO_57 (O_57,N_2719,N_2567);
nand UO_58 (O_58,N_2431,N_2530);
nand UO_59 (O_59,N_2633,N_2441);
xor UO_60 (O_60,N_2350,N_2342);
or UO_61 (O_61,N_2932,N_2387);
nand UO_62 (O_62,N_2942,N_2535);
nand UO_63 (O_63,N_2859,N_2693);
and UO_64 (O_64,N_2251,N_2611);
xnor UO_65 (O_65,N_2654,N_2771);
or UO_66 (O_66,N_2401,N_2327);
and UO_67 (O_67,N_2948,N_2866);
and UO_68 (O_68,N_2770,N_2855);
nor UO_69 (O_69,N_2950,N_2678);
nor UO_70 (O_70,N_2261,N_2460);
xnor UO_71 (O_71,N_2820,N_2556);
or UO_72 (O_72,N_2322,N_2676);
and UO_73 (O_73,N_2408,N_2798);
xnor UO_74 (O_74,N_2286,N_2330);
xnor UO_75 (O_75,N_2898,N_2720);
and UO_76 (O_76,N_2699,N_2862);
nand UO_77 (O_77,N_2659,N_2572);
nand UO_78 (O_78,N_2517,N_2291);
xnor UO_79 (O_79,N_2412,N_2434);
and UO_80 (O_80,N_2903,N_2664);
nor UO_81 (O_81,N_2975,N_2725);
or UO_82 (O_82,N_2954,N_2613);
and UO_83 (O_83,N_2630,N_2931);
nor UO_84 (O_84,N_2318,N_2514);
and UO_85 (O_85,N_2889,N_2735);
nand UO_86 (O_86,N_2254,N_2348);
or UO_87 (O_87,N_2592,N_2283);
nor UO_88 (O_88,N_2407,N_2731);
or UO_89 (O_89,N_2791,N_2747);
nand UO_90 (O_90,N_2739,N_2945);
or UO_91 (O_91,N_2609,N_2751);
or UO_92 (O_92,N_2582,N_2980);
xor UO_93 (O_93,N_2993,N_2886);
and UO_94 (O_94,N_2924,N_2428);
nor UO_95 (O_95,N_2683,N_2634);
nor UO_96 (O_96,N_2920,N_2270);
nand UO_97 (O_97,N_2354,N_2483);
or UO_98 (O_98,N_2869,N_2919);
xor UO_99 (O_99,N_2881,N_2542);
nor UO_100 (O_100,N_2406,N_2339);
or UO_101 (O_101,N_2674,N_2794);
or UO_102 (O_102,N_2278,N_2822);
or UO_103 (O_103,N_2705,N_2475);
or UO_104 (O_104,N_2761,N_2544);
or UO_105 (O_105,N_2274,N_2558);
xnor UO_106 (O_106,N_2679,N_2597);
nand UO_107 (O_107,N_2321,N_2590);
nor UO_108 (O_108,N_2885,N_2376);
xor UO_109 (O_109,N_2854,N_2518);
nor UO_110 (O_110,N_2470,N_2757);
nand UO_111 (O_111,N_2876,N_2364);
nand UO_112 (O_112,N_2847,N_2324);
and UO_113 (O_113,N_2926,N_2579);
xnor UO_114 (O_114,N_2627,N_2493);
or UO_115 (O_115,N_2413,N_2928);
or UO_116 (O_116,N_2790,N_2494);
nor UO_117 (O_117,N_2269,N_2691);
nand UO_118 (O_118,N_2644,N_2587);
xnor UO_119 (O_119,N_2758,N_2896);
nor UO_120 (O_120,N_2837,N_2534);
nor UO_121 (O_121,N_2581,N_2733);
and UO_122 (O_122,N_2420,N_2724);
xor UO_123 (O_123,N_2508,N_2645);
xnor UO_124 (O_124,N_2404,N_2585);
nand UO_125 (O_125,N_2545,N_2382);
xor UO_126 (O_126,N_2641,N_2639);
or UO_127 (O_127,N_2386,N_2701);
nand UO_128 (O_128,N_2504,N_2675);
nor UO_129 (O_129,N_2480,N_2914);
nor UO_130 (O_130,N_2571,N_2285);
xnor UO_131 (O_131,N_2833,N_2877);
or UO_132 (O_132,N_2281,N_2652);
nor UO_133 (O_133,N_2712,N_2606);
xor UO_134 (O_134,N_2843,N_2378);
nand UO_135 (O_135,N_2910,N_2686);
and UO_136 (O_136,N_2865,N_2509);
or UO_137 (O_137,N_2537,N_2555);
nand UO_138 (O_138,N_2754,N_2792);
nor UO_139 (O_139,N_2966,N_2972);
or UO_140 (O_140,N_2655,N_2684);
and UO_141 (O_141,N_2702,N_2976);
and UO_142 (O_142,N_2294,N_2445);
nor UO_143 (O_143,N_2839,N_2963);
nor UO_144 (O_144,N_2356,N_2982);
and UO_145 (O_145,N_2667,N_2366);
or UO_146 (O_146,N_2333,N_2805);
nor UO_147 (O_147,N_2259,N_2314);
and UO_148 (O_148,N_2409,N_2374);
nor UO_149 (O_149,N_2672,N_2548);
xnor UO_150 (O_150,N_2738,N_2838);
or UO_151 (O_151,N_2650,N_2812);
nor UO_152 (O_152,N_2315,N_2442);
and UO_153 (O_153,N_2313,N_2955);
nand UO_154 (O_154,N_2818,N_2763);
xor UO_155 (O_155,N_2443,N_2562);
xor UO_156 (O_156,N_2566,N_2689);
nand UO_157 (O_157,N_2799,N_2958);
xnor UO_158 (O_158,N_2784,N_2471);
nand UO_159 (O_159,N_2559,N_2301);
xor UO_160 (O_160,N_2894,N_2303);
or UO_161 (O_161,N_2605,N_2403);
or UO_162 (O_162,N_2933,N_2986);
and UO_163 (O_163,N_2529,N_2351);
and UO_164 (O_164,N_2308,N_2988);
nor UO_165 (O_165,N_2713,N_2815);
nor UO_166 (O_166,N_2753,N_2891);
nor UO_167 (O_167,N_2823,N_2956);
xnor UO_168 (O_168,N_2989,N_2878);
xnor UO_169 (O_169,N_2446,N_2888);
nor UO_170 (O_170,N_2391,N_2468);
nor UO_171 (O_171,N_2840,N_2432);
nor UO_172 (O_172,N_2601,N_2500);
and UO_173 (O_173,N_2410,N_2550);
nand UO_174 (O_174,N_2653,N_2890);
nand UO_175 (O_175,N_2959,N_2907);
and UO_176 (O_176,N_2801,N_2293);
and UO_177 (O_177,N_2568,N_2744);
and UO_178 (O_178,N_2680,N_2651);
nor UO_179 (O_179,N_2519,N_2614);
nor UO_180 (O_180,N_2287,N_2457);
and UO_181 (O_181,N_2525,N_2858);
nand UO_182 (O_182,N_2999,N_2937);
nand UO_183 (O_183,N_2995,N_2829);
xor UO_184 (O_184,N_2574,N_2806);
xor UO_185 (O_185,N_2461,N_2373);
and UO_186 (O_186,N_2265,N_2271);
nor UO_187 (O_187,N_2935,N_2363);
xnor UO_188 (O_188,N_2355,N_2658);
nor UO_189 (O_189,N_2916,N_2466);
nor UO_190 (O_190,N_2594,N_2326);
xnor UO_191 (O_191,N_2807,N_2433);
nand UO_192 (O_192,N_2380,N_2873);
or UO_193 (O_193,N_2390,N_2987);
nand UO_194 (O_194,N_2477,N_2752);
nor UO_195 (O_195,N_2455,N_2576);
nand UO_196 (O_196,N_2991,N_2295);
nor UO_197 (O_197,N_2570,N_2578);
xor UO_198 (O_198,N_2399,N_2632);
nand UO_199 (O_199,N_2554,N_2943);
nor UO_200 (O_200,N_2706,N_2549);
xnor UO_201 (O_201,N_2603,N_2912);
and UO_202 (O_202,N_2783,N_2646);
and UO_203 (O_203,N_2604,N_2272);
and UO_204 (O_204,N_2893,N_2588);
nand UO_205 (O_205,N_2848,N_2502);
and UO_206 (O_206,N_2533,N_2637);
xnor UO_207 (O_207,N_2852,N_2697);
nand UO_208 (O_208,N_2643,N_2253);
xnor UO_209 (O_209,N_2424,N_2629);
nand UO_210 (O_210,N_2727,N_2900);
nor UO_211 (O_211,N_2482,N_2715);
xor UO_212 (O_212,N_2425,N_2622);
and UO_213 (O_213,N_2828,N_2419);
and UO_214 (O_214,N_2803,N_2759);
nand UO_215 (O_215,N_2331,N_2737);
nor UO_216 (O_216,N_2346,N_2372);
nand UO_217 (O_217,N_2334,N_2941);
xnor UO_218 (O_218,N_2789,N_2398);
or UO_219 (O_219,N_2478,N_2400);
and UO_220 (O_220,N_2872,N_2343);
and UO_221 (O_221,N_2552,N_2749);
nand UO_222 (O_222,N_2856,N_2573);
or UO_223 (O_223,N_2394,N_2670);
or UO_224 (O_224,N_2619,N_2560);
xnor UO_225 (O_225,N_2307,N_2474);
or UO_226 (O_226,N_2764,N_2844);
nand UO_227 (O_227,N_2337,N_2357);
nor UO_228 (O_228,N_2338,N_2447);
nand UO_229 (O_229,N_2962,N_2396);
and UO_230 (O_230,N_2620,N_2429);
or UO_231 (O_231,N_2448,N_2551);
nand UO_232 (O_232,N_2263,N_2362);
xor UO_233 (O_233,N_2368,N_2591);
nor UO_234 (O_234,N_2540,N_2769);
nor UO_235 (O_235,N_2902,N_2897);
or UO_236 (O_236,N_2612,N_2709);
or UO_237 (O_237,N_2777,N_2345);
nor UO_238 (O_238,N_2522,N_2938);
xnor UO_239 (O_239,N_2996,N_2600);
xnor UO_240 (O_240,N_2904,N_2788);
and UO_241 (O_241,N_2825,N_2365);
nand UO_242 (O_242,N_2486,N_2846);
nor UO_243 (O_243,N_2766,N_2729);
xnor UO_244 (O_244,N_2796,N_2503);
nor UO_245 (O_245,N_2746,N_2598);
xnor UO_246 (O_246,N_2685,N_2688);
or UO_247 (O_247,N_2526,N_2359);
and UO_248 (O_248,N_2944,N_2467);
or UO_249 (O_249,N_2618,N_2880);
xnor UO_250 (O_250,N_2660,N_2625);
and UO_251 (O_251,N_2267,N_2469);
or UO_252 (O_252,N_2824,N_2964);
nand UO_253 (O_253,N_2516,N_2831);
or UO_254 (O_254,N_2786,N_2994);
and UO_255 (O_255,N_2450,N_2780);
and UO_256 (O_256,N_2415,N_2809);
nand UO_257 (O_257,N_2997,N_2395);
and UO_258 (O_258,N_2960,N_2832);
nand UO_259 (O_259,N_2707,N_2451);
and UO_260 (O_260,N_2723,N_2787);
nand UO_261 (O_261,N_2875,N_2640);
nand UO_262 (O_262,N_2489,N_2520);
xor UO_263 (O_263,N_2860,N_2834);
nor UO_264 (O_264,N_2284,N_2531);
and UO_265 (O_265,N_2377,N_2906);
and UO_266 (O_266,N_2957,N_2459);
xor UO_267 (O_267,N_2528,N_2793);
or UO_268 (O_268,N_2918,N_2464);
xor UO_269 (O_269,N_2656,N_2341);
and UO_270 (O_270,N_2539,N_2388);
and UO_271 (O_271,N_2811,N_2329);
or UO_272 (O_272,N_2527,N_2949);
nor UO_273 (O_273,N_2495,N_2990);
nor UO_274 (O_274,N_2476,N_2541);
or UO_275 (O_275,N_2320,N_2842);
xnor UO_276 (O_276,N_2849,N_2647);
and UO_277 (O_277,N_2781,N_2580);
xor UO_278 (O_278,N_2716,N_2310);
xor UO_279 (O_279,N_2266,N_2256);
nand UO_280 (O_280,N_2871,N_2940);
and UO_281 (O_281,N_2418,N_2317);
or UO_282 (O_282,N_2861,N_2804);
nor UO_283 (O_283,N_2438,N_2810);
nand UO_284 (O_284,N_2492,N_2895);
nor UO_285 (O_285,N_2610,N_2325);
and UO_286 (O_286,N_2743,N_2615);
xor UO_287 (O_287,N_2277,N_2851);
or UO_288 (O_288,N_2402,N_2423);
xnor UO_289 (O_289,N_2507,N_2481);
xor UO_290 (O_290,N_2513,N_2648);
nor UO_291 (O_291,N_2909,N_2375);
or UO_292 (O_292,N_2319,N_2961);
and UO_293 (O_293,N_2458,N_2905);
nor UO_294 (O_294,N_2817,N_2577);
nor UO_295 (O_295,N_2564,N_2728);
xor UO_296 (O_296,N_2718,N_2981);
or UO_297 (O_297,N_2296,N_2984);
and UO_298 (O_298,N_2311,N_2336);
nor UO_299 (O_299,N_2681,N_2583);
xor UO_300 (O_300,N_2487,N_2347);
xnor UO_301 (O_301,N_2742,N_2392);
nor UO_302 (O_302,N_2335,N_2741);
or UO_303 (O_303,N_2850,N_2289);
nand UO_304 (O_304,N_2521,N_2273);
nand UO_305 (O_305,N_2628,N_2250);
nor UO_306 (O_306,N_2546,N_2730);
and UO_307 (O_307,N_2306,N_2884);
or UO_308 (O_308,N_2288,N_2690);
xnor UO_309 (O_309,N_2506,N_2775);
nand UO_310 (O_310,N_2586,N_2779);
nor UO_311 (O_311,N_2276,N_2370);
nand UO_312 (O_312,N_2491,N_2523);
nor UO_313 (O_313,N_2290,N_2498);
and UO_314 (O_314,N_2607,N_2921);
nand UO_315 (O_315,N_2292,N_2553);
nand UO_316 (O_316,N_2383,N_2745);
xnor UO_317 (O_317,N_2736,N_2819);
nor UO_318 (O_318,N_2416,N_2595);
and UO_319 (O_319,N_2947,N_2708);
xor UO_320 (O_320,N_2677,N_2371);
or UO_321 (O_321,N_2340,N_2411);
and UO_322 (O_322,N_2344,N_2305);
xnor UO_323 (O_323,N_2524,N_2682);
nor UO_324 (O_324,N_2721,N_2974);
xnor UO_325 (O_325,N_2816,N_2275);
nor UO_326 (O_326,N_2328,N_2440);
xnor UO_327 (O_327,N_2808,N_2624);
nand UO_328 (O_328,N_2257,N_2449);
xor UO_329 (O_329,N_2557,N_2901);
xnor UO_330 (O_330,N_2841,N_2626);
or UO_331 (O_331,N_2454,N_2538);
or UO_332 (O_332,N_2836,N_2260);
nand UO_333 (O_333,N_2435,N_2953);
nand UO_334 (O_334,N_2532,N_2845);
xnor UO_335 (O_335,N_2936,N_2501);
nand UO_336 (O_336,N_2864,N_2456);
or UO_337 (O_337,N_2547,N_2773);
nand UO_338 (O_338,N_2665,N_2968);
xor UO_339 (O_339,N_2892,N_2642);
nor UO_340 (O_340,N_2971,N_2332);
nand UO_341 (O_341,N_2563,N_2589);
xnor UO_342 (O_342,N_2316,N_2985);
nor UO_343 (O_343,N_2970,N_2917);
xnor UO_344 (O_344,N_2369,N_2384);
nor UO_345 (O_345,N_2795,N_2765);
and UO_346 (O_346,N_2863,N_2827);
and UO_347 (O_347,N_2437,N_2497);
and UO_348 (O_348,N_2360,N_2740);
or UO_349 (O_349,N_2505,N_2979);
nor UO_350 (O_350,N_2499,N_2868);
nand UO_351 (O_351,N_2352,N_2279);
and UO_352 (O_352,N_2703,N_2453);
xor UO_353 (O_353,N_2512,N_2282);
nor UO_354 (O_354,N_2883,N_2673);
or UO_355 (O_355,N_2887,N_2417);
and UO_356 (O_356,N_2774,N_2800);
nor UO_357 (O_357,N_2367,N_2717);
or UO_358 (O_358,N_2575,N_2616);
or UO_359 (O_359,N_2669,N_2510);
nor UO_360 (O_360,N_2361,N_2379);
or UO_361 (O_361,N_2426,N_2692);
xnor UO_362 (O_362,N_2778,N_2479);
or UO_363 (O_363,N_2911,N_2300);
xor UO_364 (O_364,N_2511,N_2258);
nor UO_365 (O_365,N_2946,N_2255);
xnor UO_366 (O_366,N_2405,N_2584);
nor UO_367 (O_367,N_2496,N_2323);
nor UO_368 (O_368,N_2802,N_2299);
or UO_369 (O_369,N_2874,N_2302);
xnor UO_370 (O_370,N_2998,N_2882);
and UO_371 (O_371,N_2561,N_2762);
nor UO_372 (O_372,N_2264,N_2353);
xor UO_373 (O_373,N_2930,N_2929);
and UO_374 (O_374,N_2696,N_2687);
and UO_375 (O_375,N_2701,N_2955);
xor UO_376 (O_376,N_2750,N_2553);
nand UO_377 (O_377,N_2278,N_2645);
and UO_378 (O_378,N_2523,N_2621);
or UO_379 (O_379,N_2397,N_2517);
xnor UO_380 (O_380,N_2429,N_2366);
and UO_381 (O_381,N_2254,N_2567);
nand UO_382 (O_382,N_2814,N_2996);
or UO_383 (O_383,N_2527,N_2366);
nor UO_384 (O_384,N_2763,N_2698);
and UO_385 (O_385,N_2987,N_2862);
nand UO_386 (O_386,N_2530,N_2603);
nor UO_387 (O_387,N_2754,N_2601);
nor UO_388 (O_388,N_2812,N_2673);
nand UO_389 (O_389,N_2316,N_2916);
xor UO_390 (O_390,N_2815,N_2431);
nand UO_391 (O_391,N_2563,N_2930);
nor UO_392 (O_392,N_2413,N_2812);
xor UO_393 (O_393,N_2356,N_2354);
xnor UO_394 (O_394,N_2489,N_2285);
or UO_395 (O_395,N_2393,N_2694);
and UO_396 (O_396,N_2670,N_2705);
or UO_397 (O_397,N_2460,N_2545);
or UO_398 (O_398,N_2830,N_2857);
nand UO_399 (O_399,N_2965,N_2462);
or UO_400 (O_400,N_2554,N_2508);
and UO_401 (O_401,N_2707,N_2461);
nand UO_402 (O_402,N_2984,N_2484);
nand UO_403 (O_403,N_2395,N_2755);
nor UO_404 (O_404,N_2343,N_2741);
nor UO_405 (O_405,N_2349,N_2995);
nand UO_406 (O_406,N_2904,N_2973);
and UO_407 (O_407,N_2498,N_2689);
and UO_408 (O_408,N_2821,N_2267);
and UO_409 (O_409,N_2845,N_2646);
or UO_410 (O_410,N_2805,N_2663);
nand UO_411 (O_411,N_2600,N_2487);
nor UO_412 (O_412,N_2856,N_2310);
xnor UO_413 (O_413,N_2276,N_2831);
xnor UO_414 (O_414,N_2329,N_2291);
nor UO_415 (O_415,N_2609,N_2918);
xor UO_416 (O_416,N_2454,N_2426);
nand UO_417 (O_417,N_2891,N_2411);
nand UO_418 (O_418,N_2716,N_2942);
xnor UO_419 (O_419,N_2862,N_2844);
xnor UO_420 (O_420,N_2302,N_2306);
nand UO_421 (O_421,N_2571,N_2588);
nand UO_422 (O_422,N_2776,N_2323);
and UO_423 (O_423,N_2716,N_2524);
nand UO_424 (O_424,N_2682,N_2695);
or UO_425 (O_425,N_2658,N_2738);
nor UO_426 (O_426,N_2900,N_2372);
nor UO_427 (O_427,N_2389,N_2766);
and UO_428 (O_428,N_2807,N_2317);
or UO_429 (O_429,N_2316,N_2448);
and UO_430 (O_430,N_2265,N_2788);
or UO_431 (O_431,N_2635,N_2557);
nand UO_432 (O_432,N_2321,N_2997);
xor UO_433 (O_433,N_2459,N_2878);
nand UO_434 (O_434,N_2758,N_2867);
or UO_435 (O_435,N_2756,N_2332);
nor UO_436 (O_436,N_2968,N_2786);
and UO_437 (O_437,N_2841,N_2328);
xnor UO_438 (O_438,N_2974,N_2431);
or UO_439 (O_439,N_2824,N_2479);
nand UO_440 (O_440,N_2793,N_2468);
nor UO_441 (O_441,N_2360,N_2719);
or UO_442 (O_442,N_2468,N_2991);
and UO_443 (O_443,N_2377,N_2976);
xnor UO_444 (O_444,N_2514,N_2987);
or UO_445 (O_445,N_2991,N_2738);
nand UO_446 (O_446,N_2362,N_2806);
or UO_447 (O_447,N_2812,N_2325);
nand UO_448 (O_448,N_2296,N_2705);
nor UO_449 (O_449,N_2488,N_2306);
nand UO_450 (O_450,N_2874,N_2415);
or UO_451 (O_451,N_2807,N_2321);
nand UO_452 (O_452,N_2549,N_2520);
nor UO_453 (O_453,N_2808,N_2408);
and UO_454 (O_454,N_2323,N_2897);
nor UO_455 (O_455,N_2928,N_2712);
and UO_456 (O_456,N_2725,N_2359);
and UO_457 (O_457,N_2477,N_2979);
nand UO_458 (O_458,N_2688,N_2388);
and UO_459 (O_459,N_2521,N_2356);
and UO_460 (O_460,N_2485,N_2826);
and UO_461 (O_461,N_2478,N_2302);
and UO_462 (O_462,N_2865,N_2619);
xnor UO_463 (O_463,N_2962,N_2503);
nor UO_464 (O_464,N_2292,N_2566);
or UO_465 (O_465,N_2331,N_2665);
or UO_466 (O_466,N_2895,N_2363);
and UO_467 (O_467,N_2397,N_2546);
and UO_468 (O_468,N_2772,N_2474);
nor UO_469 (O_469,N_2517,N_2826);
nor UO_470 (O_470,N_2562,N_2265);
nand UO_471 (O_471,N_2529,N_2583);
nand UO_472 (O_472,N_2924,N_2754);
or UO_473 (O_473,N_2538,N_2728);
and UO_474 (O_474,N_2308,N_2736);
xor UO_475 (O_475,N_2973,N_2738);
and UO_476 (O_476,N_2830,N_2585);
and UO_477 (O_477,N_2353,N_2356);
or UO_478 (O_478,N_2373,N_2755);
nor UO_479 (O_479,N_2968,N_2787);
nor UO_480 (O_480,N_2711,N_2455);
and UO_481 (O_481,N_2382,N_2368);
xor UO_482 (O_482,N_2853,N_2574);
and UO_483 (O_483,N_2377,N_2300);
nor UO_484 (O_484,N_2401,N_2927);
or UO_485 (O_485,N_2826,N_2981);
and UO_486 (O_486,N_2511,N_2850);
nand UO_487 (O_487,N_2526,N_2550);
or UO_488 (O_488,N_2918,N_2258);
and UO_489 (O_489,N_2706,N_2806);
xnor UO_490 (O_490,N_2981,N_2253);
nor UO_491 (O_491,N_2666,N_2871);
and UO_492 (O_492,N_2735,N_2941);
and UO_493 (O_493,N_2305,N_2493);
or UO_494 (O_494,N_2970,N_2423);
nand UO_495 (O_495,N_2474,N_2508);
nand UO_496 (O_496,N_2367,N_2974);
nor UO_497 (O_497,N_2822,N_2877);
and UO_498 (O_498,N_2684,N_2745);
nand UO_499 (O_499,N_2661,N_2826);
endmodule