module basic_3000_30000_3500_6_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_1756,In_2788);
xnor U1 (N_1,In_871,In_2668);
nor U2 (N_2,In_1414,In_1636);
or U3 (N_3,In_2891,In_978);
nand U4 (N_4,In_2243,In_2986);
or U5 (N_5,In_868,In_854);
nor U6 (N_6,In_533,In_2097);
xnor U7 (N_7,In_1098,In_2978);
nand U8 (N_8,In_1547,In_705);
or U9 (N_9,In_882,In_2774);
xnor U10 (N_10,In_1443,In_1826);
and U11 (N_11,In_2434,In_463);
nor U12 (N_12,In_36,In_1690);
nand U13 (N_13,In_1980,In_1574);
or U14 (N_14,In_1940,In_1191);
nor U15 (N_15,In_1462,In_1758);
nand U16 (N_16,In_1737,In_588);
and U17 (N_17,In_1245,In_3);
xnor U18 (N_18,In_483,In_490);
or U19 (N_19,In_544,In_1288);
nand U20 (N_20,In_373,In_2307);
or U21 (N_21,In_2551,In_2317);
or U22 (N_22,In_770,In_1201);
xor U23 (N_23,In_1426,In_1333);
or U24 (N_24,In_2994,In_1731);
nor U25 (N_25,In_819,In_2290);
xnor U26 (N_26,In_269,In_2867);
xor U27 (N_27,In_2442,In_2359);
xnor U28 (N_28,In_1339,In_2742);
nor U29 (N_29,In_2106,In_1087);
xnor U30 (N_30,In_1799,In_1732);
nand U31 (N_31,In_934,In_2870);
and U32 (N_32,In_2211,In_2068);
or U33 (N_33,In_1870,In_432);
nor U34 (N_34,In_1919,In_948);
nand U35 (N_35,In_2067,In_1229);
xnor U36 (N_36,In_1956,In_1223);
nor U37 (N_37,In_2032,In_2917);
nand U38 (N_38,In_1225,In_1267);
nand U39 (N_39,In_1748,In_1941);
or U40 (N_40,In_733,In_2132);
or U41 (N_41,In_2661,In_701);
and U42 (N_42,In_1865,In_55);
or U43 (N_43,In_636,In_756);
nor U44 (N_44,In_2477,In_844);
or U45 (N_45,In_2529,In_2142);
or U46 (N_46,In_178,In_229);
or U47 (N_47,In_23,In_1469);
nand U48 (N_48,In_1480,In_2125);
nor U49 (N_49,In_384,In_1929);
and U50 (N_50,In_1741,In_1221);
nand U51 (N_51,In_594,In_1879);
and U52 (N_52,In_410,In_2966);
or U53 (N_53,In_2482,In_674);
and U54 (N_54,In_1592,In_680);
or U55 (N_55,In_2822,In_1935);
nand U56 (N_56,In_1358,In_267);
or U57 (N_57,In_2223,In_2023);
xor U58 (N_58,In_1202,In_2943);
xnor U59 (N_59,In_17,In_1280);
nand U60 (N_60,In_1735,In_28);
or U61 (N_61,In_200,In_1257);
xor U62 (N_62,In_1562,In_845);
or U63 (N_63,In_34,In_1241);
nor U64 (N_64,In_572,In_626);
nor U65 (N_65,In_352,In_2942);
nor U66 (N_66,In_369,In_631);
xnor U67 (N_67,In_2376,In_2603);
xor U68 (N_68,In_2162,In_2555);
nor U69 (N_69,In_2892,In_1542);
and U70 (N_70,In_2240,In_1504);
nor U71 (N_71,In_1988,In_2425);
or U72 (N_72,In_379,In_2085);
xnor U73 (N_73,In_2972,In_778);
or U74 (N_74,In_668,In_2458);
or U75 (N_75,In_302,In_2399);
or U76 (N_76,In_853,In_264);
and U77 (N_77,In_514,In_2854);
xnor U78 (N_78,In_1477,In_360);
and U79 (N_79,In_2588,In_396);
and U80 (N_80,In_93,In_2453);
nor U81 (N_81,In_951,In_2221);
nor U82 (N_82,In_163,In_1498);
or U83 (N_83,In_2430,In_1132);
and U84 (N_84,In_811,In_1903);
and U85 (N_85,In_2731,In_940);
nor U86 (N_86,In_995,In_2293);
and U87 (N_87,In_950,In_1891);
and U88 (N_88,In_8,In_1964);
and U89 (N_89,In_80,In_1286);
xor U90 (N_90,In_1308,In_608);
nand U91 (N_91,In_773,In_348);
and U92 (N_92,In_2355,In_419);
and U93 (N_93,In_120,In_2183);
or U94 (N_94,In_2487,In_371);
nand U95 (N_95,In_223,In_158);
or U96 (N_96,In_2370,In_504);
or U97 (N_97,In_2564,In_1598);
or U98 (N_98,In_211,In_2801);
nor U99 (N_99,In_2332,In_515);
xor U100 (N_100,In_1528,In_1113);
or U101 (N_101,In_2200,In_915);
xor U102 (N_102,In_1785,In_1141);
or U103 (N_103,In_428,In_2063);
or U104 (N_104,In_2165,In_2787);
and U105 (N_105,In_2439,In_737);
and U106 (N_106,In_31,In_1921);
or U107 (N_107,In_517,In_776);
or U108 (N_108,In_2356,In_532);
nand U109 (N_109,In_1108,In_1440);
or U110 (N_110,In_1079,In_1300);
xnor U111 (N_111,In_2045,In_1782);
nor U112 (N_112,In_1655,In_872);
nor U113 (N_113,In_2987,In_301);
and U114 (N_114,In_1967,In_1470);
and U115 (N_115,In_1698,In_1775);
xor U116 (N_116,In_385,In_1576);
xnor U117 (N_117,In_1990,In_1439);
and U118 (N_118,In_2506,In_255);
or U119 (N_119,In_1500,In_718);
nand U120 (N_120,In_313,In_1068);
xnor U121 (N_121,In_1003,In_2004);
nand U122 (N_122,In_1049,In_326);
xnor U123 (N_123,In_1148,In_1534);
nor U124 (N_124,In_1111,In_1037);
or U125 (N_125,In_1536,In_2009);
or U126 (N_126,In_305,In_2515);
nand U127 (N_127,In_1882,In_760);
or U128 (N_128,In_1188,In_2331);
nand U129 (N_129,In_165,In_164);
nand U130 (N_130,In_168,In_1482);
xnor U131 (N_131,In_2739,In_2929);
and U132 (N_132,In_1293,In_429);
or U133 (N_133,In_374,In_1898);
and U134 (N_134,In_1423,In_698);
nor U135 (N_135,In_1728,In_2753);
nand U136 (N_136,In_1620,In_2608);
nor U137 (N_137,In_114,In_738);
nor U138 (N_138,In_2465,In_2412);
nand U139 (N_139,In_209,In_244);
nand U140 (N_140,In_445,In_2893);
nor U141 (N_141,In_2248,In_2082);
nor U142 (N_142,In_2910,In_911);
xnor U143 (N_143,In_752,In_92);
nand U144 (N_144,In_2298,In_2746);
nand U145 (N_145,In_1118,In_652);
nand U146 (N_146,In_2034,In_1512);
nor U147 (N_147,In_2898,In_2030);
or U148 (N_148,In_2931,In_565);
nand U149 (N_149,In_709,In_696);
nor U150 (N_150,In_1472,In_2022);
nand U151 (N_151,In_2858,In_1187);
and U152 (N_152,In_1085,In_2813);
and U153 (N_153,In_858,In_2397);
and U154 (N_154,In_1294,In_1053);
xor U155 (N_155,In_2951,In_2680);
nor U156 (N_156,In_415,In_245);
or U157 (N_157,In_1046,In_2033);
nor U158 (N_158,In_386,In_720);
and U159 (N_159,In_1829,In_271);
or U160 (N_160,In_97,In_924);
or U161 (N_161,In_1106,In_1774);
nor U162 (N_162,In_1634,In_291);
or U163 (N_163,In_310,In_2559);
nor U164 (N_164,In_2694,In_1934);
and U165 (N_165,In_932,In_381);
or U166 (N_166,In_927,In_2614);
nor U167 (N_167,In_941,In_383);
and U168 (N_168,In_45,In_2872);
nor U169 (N_169,In_1797,In_1112);
and U170 (N_170,In_1939,In_336);
nor U171 (N_171,In_1601,In_2536);
xnor U172 (N_172,In_119,In_1550);
nor U173 (N_173,In_2340,In_279);
or U174 (N_174,In_1184,In_667);
and U175 (N_175,In_1691,In_1169);
xnor U176 (N_176,In_704,In_592);
nor U177 (N_177,In_1984,In_35);
nand U178 (N_178,In_2610,In_1033);
and U179 (N_179,In_1317,In_2567);
nor U180 (N_180,In_9,In_2500);
nor U181 (N_181,In_160,In_426);
xor U182 (N_182,In_723,In_1559);
xnor U183 (N_183,In_15,In_2091);
nand U184 (N_184,In_1247,In_1813);
xor U185 (N_185,In_1757,In_1677);
nor U186 (N_186,In_2761,In_1349);
nand U187 (N_187,In_2541,In_727);
and U188 (N_188,In_46,In_2887);
nand U189 (N_189,In_2020,In_1772);
and U190 (N_190,In_2617,In_574);
xor U191 (N_191,In_2259,In_2584);
xor U192 (N_192,In_2253,In_949);
or U193 (N_193,In_2964,In_187);
xnor U194 (N_194,In_579,In_382);
or U195 (N_195,In_2843,In_2900);
or U196 (N_196,In_420,In_2795);
xnor U197 (N_197,In_1072,In_1059);
nor U198 (N_198,In_1371,In_1804);
nor U199 (N_199,In_982,In_921);
nor U200 (N_200,In_1994,In_1018);
and U201 (N_201,In_1344,In_2424);
xnor U202 (N_202,In_2653,In_1743);
or U203 (N_203,In_2410,In_2764);
and U204 (N_204,In_2153,In_624);
nor U205 (N_205,In_2785,In_909);
xor U206 (N_206,In_670,In_524);
xnor U207 (N_207,In_5,In_1432);
nor U208 (N_208,In_1837,In_2383);
nand U209 (N_209,In_803,In_913);
xnor U210 (N_210,In_24,In_2285);
nand U211 (N_211,In_1022,In_306);
or U212 (N_212,In_2459,In_141);
nor U213 (N_213,In_830,In_2548);
or U214 (N_214,In_1529,In_802);
and U215 (N_215,In_2226,In_1910);
nand U216 (N_216,In_281,In_2136);
and U217 (N_217,In_1164,In_183);
or U218 (N_218,In_240,In_2542);
xor U219 (N_219,In_991,In_2815);
or U220 (N_220,In_1869,In_99);
or U221 (N_221,In_1082,In_2563);
or U222 (N_222,In_2925,In_1136);
xor U223 (N_223,In_1836,In_2543);
xor U224 (N_224,In_2521,In_242);
nand U225 (N_225,In_965,In_26);
nor U226 (N_226,In_1896,In_1137);
nor U227 (N_227,In_591,In_929);
xnor U228 (N_228,In_1971,In_1382);
and U229 (N_229,In_104,In_2039);
nand U230 (N_230,In_2092,In_2646);
and U231 (N_231,In_525,In_1633);
or U232 (N_232,In_2967,In_265);
nand U233 (N_233,In_1224,In_2440);
and U234 (N_234,In_63,In_1716);
nor U235 (N_235,In_2384,In_1906);
nor U236 (N_236,In_1638,In_2703);
xor U237 (N_237,In_2512,In_2156);
nand U238 (N_238,In_1629,In_2520);
or U239 (N_239,In_1263,In_895);
nor U240 (N_240,In_1560,In_74);
nor U241 (N_241,In_1661,In_2656);
nand U242 (N_242,In_2368,In_2489);
or U243 (N_243,In_1133,In_1884);
xor U244 (N_244,In_2171,In_1208);
nand U245 (N_245,In_1454,In_2962);
nand U246 (N_246,In_1139,In_1166);
nand U247 (N_247,In_1025,In_2985);
or U248 (N_248,In_1230,In_2880);
xnor U249 (N_249,In_421,In_1101);
or U250 (N_250,In_2480,In_536);
nand U251 (N_251,In_816,In_2935);
and U252 (N_252,In_954,In_2590);
nor U253 (N_253,In_649,In_1097);
nand U254 (N_254,In_2401,In_1096);
and U255 (N_255,In_2977,In_708);
xnor U256 (N_256,In_2301,In_1515);
or U257 (N_257,In_2704,In_922);
and U258 (N_258,In_769,In_1181);
xor U259 (N_259,In_331,In_2939);
xnor U260 (N_260,In_2343,In_2652);
nor U261 (N_261,In_361,In_604);
or U262 (N_262,In_637,In_2737);
nor U263 (N_263,In_22,In_405);
nor U264 (N_264,In_2545,In_2876);
and U265 (N_265,In_563,In_799);
or U266 (N_266,In_411,In_2629);
and U267 (N_267,In_1199,In_890);
nor U268 (N_268,In_2000,In_1408);
nor U269 (N_269,In_2375,In_2111);
xnor U270 (N_270,In_2110,In_1131);
and U271 (N_271,In_2072,In_1556);
or U272 (N_272,In_886,In_1911);
and U273 (N_273,In_587,In_1114);
or U274 (N_274,In_1438,In_539);
xor U275 (N_275,In_959,In_340);
or U276 (N_276,In_1681,In_2398);
xor U277 (N_277,In_2005,In_1261);
or U278 (N_278,In_174,In_1736);
nand U279 (N_279,In_182,In_1952);
and U280 (N_280,In_10,In_2575);
or U281 (N_281,In_2681,In_238);
or U282 (N_282,In_2561,In_962);
nand U283 (N_283,In_1733,In_1455);
xnor U284 (N_284,In_2201,In_2088);
or U285 (N_285,In_2770,In_377);
nand U286 (N_286,In_2260,In_1399);
nand U287 (N_287,In_2549,In_1285);
or U288 (N_288,In_1959,In_2616);
nor U289 (N_289,In_1369,In_103);
nor U290 (N_290,In_365,In_724);
nand U291 (N_291,In_2798,In_1676);
nor U292 (N_292,In_1525,In_1127);
nor U293 (N_293,In_139,In_2600);
or U294 (N_294,In_1890,In_2621);
nand U295 (N_295,In_1485,In_547);
xnor U296 (N_296,In_641,In_1902);
nor U297 (N_297,In_2413,In_1777);
or U298 (N_298,In_2847,In_1710);
or U299 (N_299,In_732,In_2449);
nor U300 (N_300,In_1218,In_2921);
nor U301 (N_301,In_2474,In_2249);
nand U302 (N_302,In_2129,In_12);
nand U303 (N_303,In_1771,In_457);
and U304 (N_304,In_98,In_162);
xor U305 (N_305,In_299,In_1787);
xnor U306 (N_306,In_904,In_295);
nand U307 (N_307,In_226,In_2428);
nor U308 (N_308,In_2143,In_1244);
or U309 (N_309,In_741,In_1683);
and U310 (N_310,In_1738,In_131);
nor U311 (N_311,In_1342,In_1305);
xnor U312 (N_312,In_1254,In_2537);
or U313 (N_313,In_276,In_1663);
nor U314 (N_314,In_2041,In_1753);
nand U315 (N_315,In_1965,In_914);
and U316 (N_316,In_1657,In_1255);
nor U317 (N_317,In_952,In_2958);
and U318 (N_318,In_2291,In_208);
or U319 (N_319,In_2391,In_653);
xor U320 (N_320,In_2297,In_1502);
nand U321 (N_321,In_611,In_2006);
or U322 (N_322,In_685,In_312);
nor U323 (N_323,In_2322,In_475);
nand U324 (N_324,In_1064,In_1887);
nand U325 (N_325,In_146,In_263);
nor U326 (N_326,In_1613,In_171);
nor U327 (N_327,In_656,In_699);
and U328 (N_328,In_745,In_353);
xnor U329 (N_329,In_1564,In_2818);
xor U330 (N_330,In_1778,In_2175);
and U331 (N_331,In_1316,In_2485);
nand U332 (N_332,In_2982,In_150);
xor U333 (N_333,In_2155,In_842);
and U334 (N_334,In_235,In_1554);
or U335 (N_335,In_87,In_2507);
nor U336 (N_336,In_2856,In_391);
and U337 (N_337,In_2258,In_2105);
and U338 (N_338,In_2468,In_731);
and U339 (N_339,In_792,In_878);
nor U340 (N_340,In_1400,In_2432);
xor U341 (N_341,In_323,In_1841);
nand U342 (N_342,In_2792,In_2251);
xnor U343 (N_343,In_232,In_607);
xnor U344 (N_344,In_2657,In_2745);
or U345 (N_345,In_944,In_2599);
xnor U346 (N_346,In_2579,In_1706);
and U347 (N_347,In_2015,In_1711);
and U348 (N_348,In_1608,In_1495);
nand U349 (N_349,In_42,In_2911);
xor U350 (N_350,In_956,In_1944);
nor U351 (N_351,In_2268,In_450);
xnor U352 (N_352,In_2984,In_2729);
nand U353 (N_353,In_1395,In_994);
xor U354 (N_354,In_1381,In_2674);
nand U355 (N_355,In_2754,In_60);
nand U356 (N_356,In_2637,In_2271);
nand U357 (N_357,In_444,In_970);
or U358 (N_358,In_783,In_1893);
xor U359 (N_359,In_2367,In_1056);
nor U360 (N_360,In_218,In_273);
xor U361 (N_361,In_988,In_1522);
and U362 (N_362,In_2740,In_2855);
or U363 (N_363,In_1093,In_1042);
and U364 (N_364,In_1780,In_2216);
and U365 (N_365,In_2626,In_2250);
nand U366 (N_366,In_2677,In_791);
and U367 (N_367,In_49,In_1957);
and U368 (N_368,In_1960,In_2148);
xor U369 (N_369,In_1198,In_2237);
nand U370 (N_370,In_857,In_1610);
and U371 (N_371,In_1770,In_580);
nand U372 (N_372,In_1066,In_2812);
or U373 (N_373,In_290,In_37);
nor U374 (N_374,In_275,In_512);
or U375 (N_375,In_744,In_1256);
xnor U376 (N_376,In_2885,In_801);
nor U377 (N_377,In_846,In_2077);
xor U378 (N_378,In_2841,In_2641);
nor U379 (N_379,In_378,In_1461);
nand U380 (N_380,In_300,In_2714);
and U381 (N_381,In_1321,In_2938);
nand U382 (N_382,In_710,In_1332);
nor U383 (N_383,In_1850,In_1034);
or U384 (N_384,In_864,In_1745);
and U385 (N_385,In_2934,In_459);
and U386 (N_386,In_2056,In_1326);
nor U387 (N_387,In_838,In_730);
nand U388 (N_388,In_1631,In_2662);
and U389 (N_389,In_1820,In_133);
nor U390 (N_390,In_1206,In_648);
nor U391 (N_391,In_2471,In_810);
nor U392 (N_392,In_917,In_2825);
and U393 (N_393,In_589,In_1217);
and U394 (N_394,In_2326,In_2918);
and U395 (N_395,In_1784,In_2107);
and U396 (N_396,In_2882,In_422);
and U397 (N_397,In_2286,In_1604);
and U398 (N_398,In_397,In_2347);
nor U399 (N_399,In_751,In_717);
nor U400 (N_400,In_2262,In_2246);
nand U401 (N_401,In_1645,In_1273);
nand U402 (N_402,In_2722,In_25);
nor U403 (N_403,In_347,In_1074);
or U404 (N_404,In_203,In_69);
nor U405 (N_405,In_1212,In_2276);
and U406 (N_406,In_1532,In_394);
nor U407 (N_407,In_1553,In_1912);
and U408 (N_408,In_1015,In_315);
and U409 (N_409,In_1165,In_283);
nand U410 (N_410,In_2344,In_169);
nor U411 (N_411,In_818,In_2065);
nor U412 (N_412,In_1573,In_2360);
and U413 (N_413,In_1005,In_407);
and U414 (N_414,In_1763,In_2470);
and U415 (N_415,In_2491,In_1595);
xnor U416 (N_416,In_2631,In_330);
nand U417 (N_417,In_246,In_1682);
or U418 (N_418,In_1453,In_2669);
xor U419 (N_419,In_111,In_1476);
or U420 (N_420,In_502,In_960);
nor U421 (N_421,In_205,In_2724);
or U422 (N_422,In_1147,In_984);
xor U423 (N_423,In_73,In_317);
xnor U424 (N_424,In_1351,In_1549);
or U425 (N_425,In_1719,In_2752);
xnor U426 (N_426,In_1843,In_6);
or U427 (N_427,In_1411,In_625);
nand U428 (N_428,In_1109,In_2907);
nand U429 (N_429,In_1272,In_2601);
and U430 (N_430,In_1295,In_81);
and U431 (N_431,In_2712,In_1751);
xor U432 (N_432,In_1117,In_1236);
nor U433 (N_433,In_1593,In_1430);
nor U434 (N_434,In_206,In_1897);
and U435 (N_435,In_578,In_1848);
xor U436 (N_436,In_2134,In_2634);
nor U437 (N_437,In_893,In_2509);
xor U438 (N_438,In_1590,In_2896);
xnor U439 (N_439,In_501,In_1999);
nand U440 (N_440,In_477,In_2625);
nor U441 (N_441,In_173,In_322);
or U442 (N_442,In_2450,In_2980);
and U443 (N_443,In_243,In_2647);
nor U444 (N_444,In_774,In_1918);
and U445 (N_445,In_1947,In_474);
nand U446 (N_446,In_2054,In_2596);
xnor U447 (N_447,In_2195,In_543);
nand U448 (N_448,In_387,In_2025);
xor U449 (N_449,In_33,In_815);
nor U450 (N_450,In_393,In_2203);
and U451 (N_451,In_2350,In_481);
nor U452 (N_452,In_1673,In_2803);
or U453 (N_453,In_742,In_86);
nor U454 (N_454,In_2715,In_2008);
or U455 (N_455,In_2152,In_906);
nor U456 (N_456,In_1838,In_1242);
nor U457 (N_457,In_2835,In_77);
and U458 (N_458,In_2619,In_1889);
nand U459 (N_459,In_1614,In_2863);
or U460 (N_460,In_2042,In_754);
or U461 (N_461,In_1986,In_758);
nor U462 (N_462,In_2615,In_2342);
nor U463 (N_463,In_1130,In_2915);
and U464 (N_464,In_2027,In_1185);
nand U465 (N_465,In_2127,In_431);
and U466 (N_466,In_767,In_1311);
nor U467 (N_467,In_1290,In_2264);
xor U468 (N_468,In_1872,In_2313);
nand U469 (N_469,In_0,In_2700);
xor U470 (N_470,In_2577,In_1157);
nand U471 (N_471,In_1177,In_1020);
xnor U472 (N_472,In_2636,In_1805);
or U473 (N_473,In_1142,In_2429);
or U474 (N_474,In_2275,In_850);
or U475 (N_475,In_496,In_2809);
nor U476 (N_476,In_593,In_2169);
or U477 (N_477,In_342,In_2282);
xnor U478 (N_478,In_1880,In_985);
nor U479 (N_479,In_2511,In_561);
or U480 (N_480,In_1266,In_938);
or U481 (N_481,In_1628,In_1240);
and U482 (N_482,In_2963,In_1483);
xor U483 (N_483,In_2050,In_1922);
xor U484 (N_484,In_1159,In_1468);
or U485 (N_485,In_2578,In_1140);
and U486 (N_486,In_1367,In_1600);
nand U487 (N_487,In_1626,In_1781);
or U488 (N_488,In_1589,In_1760);
and U489 (N_489,In_493,In_1943);
xor U490 (N_490,In_2757,In_224);
and U491 (N_491,In_412,In_1403);
or U492 (N_492,In_1588,In_1761);
nand U493 (N_493,In_2877,In_1662);
nand U494 (N_494,In_1834,In_1568);
and U495 (N_495,In_2270,In_1852);
nand U496 (N_496,In_2622,In_1954);
nand U497 (N_497,In_355,In_1209);
or U498 (N_498,In_2035,In_2119);
xnor U499 (N_499,In_2163,In_1660);
xnor U500 (N_500,In_2311,In_2281);
and U501 (N_501,In_1540,In_2922);
and U502 (N_502,In_1161,In_230);
or U503 (N_503,In_1010,In_2678);
nor U504 (N_504,In_2498,In_1647);
xnor U505 (N_505,In_1615,In_1086);
nor U506 (N_506,In_2151,In_1277);
xnor U507 (N_507,In_2396,In_366);
or U508 (N_508,In_1648,In_1656);
and U509 (N_509,In_210,In_2386);
xor U510 (N_510,In_2292,In_1475);
xor U511 (N_511,In_2665,In_1581);
nor U512 (N_512,In_602,In_1653);
xor U513 (N_513,In_1125,In_2036);
nor U514 (N_514,In_1537,In_392);
nand U515 (N_515,In_1584,In_2496);
and U516 (N_516,In_2182,In_1669);
nand U517 (N_517,In_2233,In_1864);
nor U518 (N_518,In_196,In_953);
and U519 (N_519,In_2598,In_2352);
and U520 (N_520,In_1077,In_2274);
nor U521 (N_521,In_750,In_138);
and U522 (N_522,In_356,In_1806);
or U523 (N_523,In_1810,In_601);
nand U524 (N_524,In_254,In_2849);
xnor U525 (N_525,In_2024,In_814);
and U526 (N_526,In_454,In_584);
and U527 (N_527,In_2658,In_2975);
or U528 (N_528,In_390,In_116);
and U529 (N_529,In_2354,In_1039);
and U530 (N_530,In_837,In_1110);
or U531 (N_531,In_1531,In_2905);
nor U532 (N_532,In_2012,In_2941);
or U533 (N_533,In_715,In_2130);
nor U534 (N_534,In_1678,In_1302);
nor U535 (N_535,In_2883,In_1160);
or U536 (N_536,In_2374,In_1855);
nor U537 (N_537,In_1019,In_1035);
xnor U538 (N_538,In_2522,In_370);
and U539 (N_539,In_1231,In_1445);
nor U540 (N_540,In_2433,In_1951);
nor U541 (N_541,In_167,In_1765);
nand U542 (N_542,In_376,In_297);
xnor U543 (N_543,In_1192,In_839);
nor U544 (N_544,In_2123,In_1200);
nor U545 (N_545,In_603,In_38);
or U546 (N_546,In_2423,In_1849);
or U547 (N_547,In_1750,In_1196);
nor U548 (N_548,In_1714,In_2701);
nand U549 (N_549,In_1379,In_1665);
xnor U550 (N_550,In_102,In_1494);
nor U551 (N_551,In_615,In_2090);
xor U552 (N_552,In_796,In_1135);
or U553 (N_553,In_2362,In_1625);
and U554 (N_554,In_1586,In_1004);
nor U555 (N_555,In_296,In_2048);
nor U556 (N_556,In_2139,In_2167);
nand U557 (N_557,In_556,In_1450);
xnor U558 (N_558,In_1276,In_806);
and U559 (N_559,In_2087,In_1828);
xor U560 (N_560,In_2059,In_585);
and U561 (N_561,In_1624,In_1124);
and U562 (N_562,In_1684,In_2895);
nor U563 (N_563,In_761,In_1523);
or U564 (N_564,In_1888,In_740);
and U565 (N_565,In_2516,In_765);
nor U566 (N_566,In_1417,In_1579);
nand U567 (N_567,In_321,In_2190);
and U568 (N_568,In_90,In_623);
and U569 (N_569,In_706,In_2762);
nand U570 (N_570,In_2562,In_916);
nor U571 (N_571,In_1355,In_2288);
nand U572 (N_572,In_1409,In_1023);
and U573 (N_573,In_847,In_1707);
xnor U574 (N_574,In_646,In_942);
or U575 (N_575,In_919,In_1530);
and U576 (N_576,In_2750,In_654);
and U577 (N_577,In_2414,In_1103);
or U578 (N_578,In_1388,In_2114);
xor U579 (N_579,In_1958,In_2231);
xnor U580 (N_580,In_2379,In_1526);
xor U581 (N_581,In_2671,In_2914);
and U582 (N_582,In_566,In_2533);
xor U583 (N_583,In_1116,In_1366);
or U584 (N_584,In_494,In_1812);
or U585 (N_585,In_2767,In_1027);
xnor U586 (N_586,In_2899,In_2613);
nor U587 (N_587,In_2310,In_1178);
xor U588 (N_588,In_1668,In_1174);
or U589 (N_589,In_1754,In_1394);
nor U590 (N_590,In_1269,In_21);
and U591 (N_591,In_1138,In_2888);
nor U592 (N_592,In_1292,In_1908);
nand U593 (N_593,In_2540,In_1687);
and U594 (N_594,In_2644,In_880);
and U595 (N_595,In_57,In_2446);
nor U596 (N_596,In_1817,In_763);
nand U597 (N_597,In_2569,In_655);
and U598 (N_598,In_2273,In_2388);
and U599 (N_599,In_2829,In_2624);
xnor U600 (N_600,In_47,In_2377);
xnor U601 (N_601,In_1343,In_1458);
nand U602 (N_602,In_939,In_1516);
xor U603 (N_603,In_2538,In_339);
xor U604 (N_604,In_827,In_664);
xor U605 (N_605,In_2832,In_1876);
xnor U606 (N_606,In_2011,In_700);
and U607 (N_607,In_1981,In_2560);
xor U608 (N_608,In_1238,In_1220);
nor U609 (N_609,In_1569,In_2417);
nand U610 (N_610,In_256,In_2776);
xor U611 (N_611,In_2859,In_537);
and U612 (N_612,In_1347,In_359);
or U613 (N_613,In_2699,In_2719);
xnor U614 (N_614,In_2490,In_1524);
or U615 (N_615,In_1877,In_143);
and U616 (N_616,In_1128,In_2051);
or U617 (N_617,In_912,In_2821);
nor U618 (N_618,In_2236,In_337);
and U619 (N_619,In_852,In_1617);
nand U620 (N_620,In_1378,In_983);
or U621 (N_621,In_2808,In_1466);
nor U622 (N_622,In_2959,In_2928);
nor U623 (N_623,In_1794,In_2889);
nand U624 (N_624,In_786,In_2070);
and U625 (N_625,In_1099,In_318);
nor U626 (N_626,In_781,In_294);
xnor U627 (N_627,In_1508,In_1216);
xnor U628 (N_628,In_441,In_1839);
or U629 (N_629,In_568,In_2956);
or U630 (N_630,In_2185,In_2353);
and U631 (N_631,In_461,In_748);
and U632 (N_632,In_947,In_307);
or U633 (N_633,In_179,In_2814);
nand U634 (N_634,In_2604,In_1724);
xnor U635 (N_635,In_1377,In_251);
nor U636 (N_636,In_258,In_1410);
nor U637 (N_637,In_425,In_2709);
or U638 (N_638,In_1237,In_2351);
nor U639 (N_639,In_531,In_682);
or U640 (N_640,In_1413,In_1821);
or U641 (N_641,In_851,In_1544);
nor U642 (N_642,In_553,In_1422);
nor U643 (N_643,In_1641,In_634);
or U644 (N_644,In_686,In_1210);
xor U645 (N_645,In_1709,In_1907);
or U646 (N_646,In_480,In_252);
or U647 (N_647,In_2502,In_1071);
nand U648 (N_648,In_1699,In_2472);
or U649 (N_649,In_39,In_2944);
nand U650 (N_650,In_695,In_1689);
nor U651 (N_651,In_1497,In_2057);
nor U652 (N_652,In_1298,In_2495);
xor U653 (N_653,In_1070,In_1666);
nand U654 (N_654,In_1747,In_571);
nand U655 (N_655,In_2689,In_2643);
or U656 (N_656,In_840,In_2003);
and U657 (N_657,In_2,In_1393);
nor U658 (N_658,In_2390,In_2804);
nand U659 (N_659,In_1664,In_647);
nand U660 (N_660,In_1383,In_2860);
nor U661 (N_661,In_747,In_19);
or U662 (N_662,In_2728,In_1885);
and U663 (N_663,In_675,In_961);
nand U664 (N_664,In_1863,In_1658);
nor U665 (N_665,In_2651,In_1211);
nor U666 (N_666,In_1167,In_2756);
nor U667 (N_667,In_1808,In_1370);
xnor U668 (N_668,In_2630,In_354);
and U669 (N_669,In_622,In_257);
nand U670 (N_670,In_2320,In_1441);
or U671 (N_671,In_1704,In_794);
and U672 (N_672,In_1953,In_1356);
nor U673 (N_673,In_2947,In_1433);
xnor U674 (N_674,In_1606,In_1840);
nor U675 (N_675,In_1705,In_2945);
or U676 (N_676,In_1832,In_438);
and U677 (N_677,In_1041,In_1926);
xnor U678 (N_678,In_2639,In_149);
xnor U679 (N_679,In_2089,In_2204);
or U680 (N_680,In_2389,In_805);
and U681 (N_681,In_228,In_2137);
xor U682 (N_682,In_2627,In_2193);
nand U683 (N_683,In_825,In_2079);
or U684 (N_684,In_2664,In_777);
and U685 (N_685,In_1189,In_1444);
nand U686 (N_686,In_2772,In_1402);
xor U687 (N_687,In_1437,In_2912);
or U688 (N_688,In_2328,In_285);
and U689 (N_689,In_2611,In_367);
nand U690 (N_690,In_1992,In_1718);
xnor U691 (N_691,In_2196,In_552);
or U692 (N_692,In_2705,In_2294);
xor U693 (N_693,In_436,In_2261);
or U694 (N_694,In_1779,In_2744);
xnor U695 (N_695,In_107,In_1203);
nand U696 (N_696,In_1640,In_2903);
nor U697 (N_697,In_1875,In_1013);
or U698 (N_698,In_2791,In_888);
and U699 (N_699,In_1451,In_1091);
or U700 (N_700,In_905,In_2830);
or U701 (N_701,In_2407,In_780);
or U702 (N_702,In_2284,In_509);
xnor U703 (N_703,In_1028,In_808);
nand U704 (N_704,In_1977,In_1252);
nand U705 (N_705,In_2846,In_1353);
and U706 (N_706,In_1949,In_651);
nor U707 (N_707,In_1583,In_32);
or U708 (N_708,In_2698,In_1274);
and U709 (N_709,In_2467,In_1802);
and U710 (N_710,In_1197,In_2099);
xnor U711 (N_711,In_1854,In_1501);
or U712 (N_712,In_1162,In_677);
and U713 (N_713,In_1966,In_856);
xnor U714 (N_714,In_1092,In_2706);
or U715 (N_715,In_2265,In_2209);
nand U716 (N_716,In_14,In_2215);
nand U717 (N_717,In_1175,In_2161);
nand U718 (N_718,In_2404,In_212);
nand U719 (N_719,In_1868,In_1492);
or U720 (N_720,In_40,In_687);
xnor U721 (N_721,In_460,In_2325);
nor U722 (N_722,In_1611,In_2278);
and U723 (N_723,In_2186,In_345);
nand U724 (N_724,In_2831,In_2807);
nand U725 (N_725,In_2102,In_2513);
or U726 (N_726,In_2295,In_153);
nand U727 (N_727,In_101,In_1916);
or U728 (N_728,In_1642,In_351);
and U729 (N_729,In_1798,In_1612);
nor U730 (N_730,In_2527,In_1637);
or U731 (N_731,In_1412,In_1734);
nor U732 (N_732,In_2074,In_557);
xor U733 (N_733,In_2989,In_2763);
and U734 (N_734,In_2688,In_753);
or U735 (N_735,In_2749,In_1467);
nand U736 (N_736,In_2920,In_1696);
nand U737 (N_737,In_79,In_2333);
or U738 (N_738,In_2990,In_1519);
xnor U739 (N_739,In_1151,In_2842);
and U740 (N_740,In_1243,In_2805);
nand U741 (N_741,In_1373,In_1713);
nor U742 (N_742,In_2224,In_1183);
nand U743 (N_743,In_2154,In_719);
nor U744 (N_744,In_1350,In_2323);
xor U745 (N_745,In_2418,In_1487);
and U746 (N_746,In_518,In_2363);
xor U747 (N_747,In_2451,In_217);
xnor U748 (N_748,In_2777,In_2881);
or U749 (N_749,In_2837,In_2773);
xnor U750 (N_750,In_2150,In_134);
nor U751 (N_751,In_346,In_2164);
nand U752 (N_752,In_1258,In_2933);
nand U753 (N_753,In_1831,In_1670);
nor U754 (N_754,In_1945,In_1322);
or U755 (N_755,In_2607,In_2239);
xnor U756 (N_756,In_1156,In_2733);
xnor U757 (N_757,In_1715,In_2748);
xnor U758 (N_758,In_1909,In_1180);
nand U759 (N_759,In_892,In_1051);
and U760 (N_760,In_262,In_875);
xnor U761 (N_761,In_2810,In_2147);
xor U762 (N_762,In_722,In_2210);
xor U763 (N_763,In_2334,In_449);
and U764 (N_764,In_2602,In_1712);
or U765 (N_765,In_2387,In_974);
xor U766 (N_766,In_638,In_437);
or U767 (N_767,In_1702,In_1320);
or U768 (N_768,In_274,In_1291);
and U769 (N_769,In_2444,In_1597);
nor U770 (N_770,In_1521,In_124);
or U771 (N_771,In_234,In_2718);
nor U772 (N_772,In_2174,In_1561);
nor U773 (N_773,In_2086,In_225);
and U774 (N_774,In_1851,In_1917);
xor U775 (N_775,In_123,In_976);
or U776 (N_776,In_2635,In_1357);
nand U777 (N_777,In_2071,In_2031);
nor U778 (N_778,In_693,In_800);
nand U779 (N_779,In_889,In_1105);
and U780 (N_780,In_1040,In_1535);
nand U781 (N_781,In_787,In_2369);
xnor U782 (N_782,In_2280,In_2973);
nand U783 (N_783,In_1948,In_729);
nand U784 (N_784,In_1630,In_1009);
xnor U785 (N_785,In_2597,In_1674);
and U786 (N_786,In_891,In_2642);
and U787 (N_787,In_2122,In_2064);
xnor U788 (N_788,In_488,In_2488);
and U789 (N_789,In_835,In_197);
and U790 (N_790,In_848,In_1892);
and U791 (N_791,In_1859,In_734);
nand U792 (N_792,In_2927,In_1284);
or U793 (N_793,In_1920,In_1816);
or U794 (N_794,In_1420,In_817);
or U795 (N_795,In_1759,In_433);
or U796 (N_796,In_314,In_508);
nor U797 (N_797,In_2845,In_1352);
nand U798 (N_798,In_1154,In_2256);
xnor U799 (N_799,In_2727,In_2593);
nor U800 (N_800,In_1328,In_448);
and U801 (N_801,In_408,In_1749);
nand U802 (N_802,In_1260,In_1900);
or U803 (N_803,In_380,In_13);
xnor U804 (N_804,In_467,In_628);
xor U805 (N_805,In_1845,In_94);
or U806 (N_806,In_2075,In_1930);
nand U807 (N_807,In_2539,In_2547);
or U808 (N_808,In_413,In_586);
nor U809 (N_809,In_1102,In_2241);
and U810 (N_810,In_2638,In_2118);
nand U811 (N_811,In_1987,In_665);
and U812 (N_812,In_530,In_2436);
or U813 (N_813,In_430,In_689);
nor U814 (N_814,In_52,In_1324);
or U815 (N_815,In_1163,In_2940);
nor U816 (N_816,In_2871,In_2420);
nand U817 (N_817,In_2371,In_2672);
or U818 (N_818,In_1835,In_2946);
or U819 (N_819,In_227,In_1993);
and U820 (N_820,In_248,In_2851);
nor U821 (N_821,In_1415,In_1858);
or U822 (N_822,In_375,In_755);
or U823 (N_823,In_873,In_1739);
nor U824 (N_824,In_2393,In_2277);
or U825 (N_825,In_2572,In_1686);
or U826 (N_826,In_2208,In_1672);
nor U827 (N_827,In_1222,In_96);
xnor U828 (N_828,In_478,In_1011);
nand U829 (N_829,In_2645,In_928);
nor U830 (N_830,In_2519,In_2014);
or U831 (N_831,In_287,In_268);
and U832 (N_832,In_2811,In_1310);
nand U833 (N_833,In_703,In_2225);
nor U834 (N_834,In_2199,In_121);
and U835 (N_835,In_2178,In_1539);
xnor U836 (N_836,In_1570,In_2349);
nor U837 (N_837,In_1895,In_1693);
xnor U838 (N_838,In_7,In_1464);
xnor U839 (N_839,In_870,In_286);
nor U840 (N_840,In_2995,In_713);
nand U841 (N_841,In_2720,In_2696);
or U842 (N_842,In_1296,In_2850);
and U843 (N_843,In_2784,In_1639);
or U844 (N_844,In_2405,In_2403);
nor U845 (N_845,In_1146,In_1143);
nor U846 (N_846,In_491,In_100);
nand U847 (N_847,In_192,In_2866);
xor U848 (N_848,In_485,In_2969);
nor U849 (N_849,In_1061,In_1271);
and U850 (N_850,In_404,In_2053);
nor U851 (N_851,In_2766,In_881);
xor U852 (N_852,In_798,In_2457);
nor U853 (N_853,In_2052,In_2663);
and U854 (N_854,In_304,In_401);
xor U855 (N_855,In_2769,In_1416);
or U856 (N_856,In_2738,In_2550);
and U857 (N_857,In_2255,In_826);
xor U858 (N_858,In_510,In_797);
and U859 (N_859,In_507,In_2001);
nor U860 (N_860,In_546,In_920);
xor U861 (N_861,In_2484,In_1856);
and U862 (N_862,In_1936,In_456);
nor U863 (N_863,In_298,In_1318);
and U864 (N_864,In_1622,In_1435);
or U865 (N_865,In_1538,In_503);
or U866 (N_866,In_1619,In_1607);
nor U867 (N_867,In_2247,In_2957);
xor U868 (N_868,In_2029,In_1490);
or U869 (N_869,In_2932,In_1717);
nor U870 (N_870,In_902,In_2654);
xor U871 (N_871,In_1818,In_2840);
nor U872 (N_872,In_2628,In_2454);
or U873 (N_873,In_1545,In_129);
and U874 (N_874,In_2552,In_1179);
or U875 (N_875,In_1878,In_2535);
and U876 (N_876,In_2768,In_2267);
nor U877 (N_877,In_529,In_2501);
xnor U878 (N_878,In_599,In_468);
nand U879 (N_879,In_464,In_1995);
and U880 (N_880,In_1488,In_1172);
nor U881 (N_881,In_759,In_1030);
xor U882 (N_882,In_2345,In_2166);
nor U883 (N_883,In_1558,In_202);
nor U884 (N_884,In_91,In_2659);
nor U885 (N_885,In_2466,In_2786);
nor U886 (N_886,In_2104,In_127);
nor U887 (N_887,In_1038,In_813);
xnor U888 (N_888,In_2517,In_2443);
nor U889 (N_889,In_633,In_505);
nor U890 (N_890,In_2864,In_2886);
nand U891 (N_891,In_1251,In_2518);
nor U892 (N_892,In_618,In_1398);
nor U893 (N_893,In_2416,In_2483);
xnor U894 (N_894,In_1924,In_1396);
or U895 (N_895,In_899,In_2721);
xnor U896 (N_896,In_213,In_1431);
and U897 (N_897,In_1048,In_746);
nor U898 (N_898,In_148,In_550);
nand U899 (N_899,In_2976,In_2198);
and U900 (N_900,In_1591,In_358);
nand U901 (N_901,In_1546,In_1679);
nand U902 (N_902,In_2263,In_2212);
xnor U903 (N_903,In_1582,In_1755);
and U904 (N_904,In_2395,In_898);
and U905 (N_905,In_484,In_1227);
nand U906 (N_906,In_2875,In_2794);
nand U907 (N_907,In_2955,In_678);
or U908 (N_908,In_1983,In_155);
and U909 (N_909,In_1474,In_694);
nand U910 (N_910,In_1002,In_1998);
nand U911 (N_911,In_2116,In_1866);
or U912 (N_912,In_1170,In_901);
nand U913 (N_913,In_1384,In_495);
or U914 (N_914,In_1786,In_2452);
and U915 (N_915,In_1844,In_1942);
or U916 (N_916,In_749,In_2026);
or U917 (N_917,In_1587,In_1278);
or U918 (N_918,In_2983,In_2775);
nor U919 (N_919,In_2916,In_2479);
xor U920 (N_920,In_945,In_1297);
and U921 (N_921,In_2133,In_1688);
nand U922 (N_922,In_2269,In_2965);
nor U923 (N_923,In_2826,In_534);
nor U924 (N_924,In_1685,In_53);
nor U925 (N_925,In_1335,In_122);
and U926 (N_926,In_56,In_2609);
nand U927 (N_927,In_2834,In_2016);
nand U928 (N_928,In_2828,In_1193);
or U929 (N_929,In_2289,In_2018);
or U930 (N_930,In_1069,In_1923);
nor U931 (N_931,In_1815,In_2574);
and U932 (N_932,In_2191,In_1792);
nand U933 (N_933,In_2702,In_2108);
or U934 (N_934,In_498,In_2038);
nand U935 (N_935,In_997,In_1289);
and U936 (N_936,In_190,In_2968);
nor U937 (N_937,In_521,In_350);
nor U938 (N_938,In_596,In_112);
and U939 (N_939,In_2385,In_925);
and U940 (N_940,In_2558,In_2974);
and U941 (N_941,In_1052,In_620);
nand U942 (N_942,In_2207,In_2117);
xnor U943 (N_943,In_11,In_417);
and U944 (N_944,In_2257,In_2230);
or U945 (N_945,In_204,In_115);
or U946 (N_946,In_201,In_1505);
and U947 (N_947,In_2338,In_1567);
nand U948 (N_948,In_1123,In_2580);
and U949 (N_949,In_721,In_2179);
or U950 (N_950,In_1652,In_859);
and U951 (N_951,In_1375,In_541);
nand U952 (N_952,In_542,In_272);
nor U953 (N_953,In_1968,In_2514);
and U954 (N_954,In_2667,In_1213);
and U955 (N_955,In_972,In_2675);
or U956 (N_956,In_2463,In_1727);
xnor U957 (N_957,In_1486,In_1788);
or U958 (N_958,In_2146,In_1667);
nand U959 (N_959,In_2227,In_2504);
and U960 (N_960,In_516,In_62);
nand U961 (N_961,In_1575,In_1186);
nand U962 (N_962,In_1833,In_44);
xor U963 (N_963,In_2632,In_1259);
nor U964 (N_964,In_1153,In_883);
xor U965 (N_965,In_1694,In_1449);
and U966 (N_966,In_2321,In_1932);
nor U967 (N_967,In_726,In_1007);
nor U968 (N_968,In_176,In_329);
nor U969 (N_969,In_30,In_2202);
or U970 (N_970,In_519,In_673);
or U971 (N_971,In_1571,In_1618);
and U972 (N_972,In_1963,In_2824);
or U973 (N_973,In_548,In_319);
and U974 (N_974,In_2476,In_2462);
xnor U975 (N_975,In_629,In_2464);
nor U976 (N_976,In_1972,In_918);
or U977 (N_977,In_2017,In_2790);
nor U978 (N_978,In_159,In_1078);
xnor U979 (N_979,In_1058,In_2408);
and U980 (N_980,In_581,In_2741);
or U981 (N_981,In_1790,In_820);
xnor U982 (N_982,In_154,In_2244);
xor U983 (N_983,In_1032,In_650);
and U984 (N_984,In_1905,In_447);
xor U985 (N_985,In_963,In_1385);
nand U986 (N_986,In_1773,In_2758);
xor U987 (N_987,In_2848,In_849);
or U988 (N_988,In_71,In_1860);
and U989 (N_989,In_2080,In_1397);
and U990 (N_990,In_990,In_980);
xor U991 (N_991,In_2013,In_1460);
and U992 (N_992,In_1204,In_943);
nor U993 (N_993,In_126,In_1746);
nand U994 (N_994,In_946,In_2095);
nand U995 (N_995,In_1471,In_1931);
and U996 (N_996,In_399,In_1914);
nor U997 (N_997,In_1447,In_2684);
xnor U998 (N_998,In_1446,In_1329);
or U999 (N_999,In_1533,In_1946);
nor U1000 (N_1000,In_2556,In_1809);
or U1001 (N_1001,In_2582,In_1473);
nand U1002 (N_1002,In_834,In_2305);
xor U1003 (N_1003,In_2531,In_1764);
nor U1004 (N_1004,In_2073,In_1726);
and U1005 (N_1005,In_1119,In_1627);
nor U1006 (N_1006,In_2197,In_527);
xor U1007 (N_1007,In_2228,In_1171);
and U1008 (N_1008,In_423,In_1361);
and U1009 (N_1009,In_1359,In_632);
nor U1010 (N_1010,In_619,In_1006);
xor U1011 (N_1011,In_1605,In_1692);
nor U1012 (N_1012,In_2525,In_2760);
xor U1013 (N_1013,In_2492,In_2234);
xnor U1014 (N_1014,In_2318,In_2981);
or U1015 (N_1015,In_479,In_95);
xnor U1016 (N_1016,In_400,In_2469);
or U1017 (N_1017,In_630,In_979);
or U1018 (N_1018,In_2557,In_2218);
xor U1019 (N_1019,In_237,In_2587);
and U1020 (N_1020,In_1427,In_147);
nand U1021 (N_1021,In_1503,In_964);
nand U1022 (N_1022,In_926,In_2783);
and U1023 (N_1023,In_823,In_635);
and U1024 (N_1024,In_2098,In_2861);
nand U1025 (N_1025,In_545,In_1345);
and U1026 (N_1026,In_1248,In_1150);
xnor U1027 (N_1027,In_247,In_669);
nand U1028 (N_1028,In_2061,In_145);
xor U1029 (N_1029,In_1513,In_1100);
xor U1030 (N_1030,In_1270,In_2112);
or U1031 (N_1031,In_1659,In_1392);
or U1032 (N_1032,In_2586,In_2735);
xor U1033 (N_1033,In_1509,In_231);
nand U1034 (N_1034,In_809,In_128);
nand U1035 (N_1035,In_492,In_427);
nand U1036 (N_1036,In_969,In_471);
or U1037 (N_1037,In_1239,In_1842);
and U1038 (N_1038,In_2019,In_1448);
nor U1039 (N_1039,In_2486,In_1800);
and U1040 (N_1040,In_113,In_1742);
nand U1041 (N_1041,In_993,In_836);
xor U1042 (N_1042,In_325,In_1089);
or U1043 (N_1043,In_117,In_1867);
nor U1044 (N_1044,In_967,In_2904);
nor U1045 (N_1045,In_1299,In_2327);
nand U1046 (N_1046,In_2923,In_2180);
nand U1047 (N_1047,In_1978,In_771);
or U1048 (N_1048,In_975,In_1017);
nor U1049 (N_1049,In_2930,In_616);
nor U1050 (N_1050,In_486,In_1234);
or U1051 (N_1051,In_2300,In_335);
nand U1052 (N_1052,In_923,In_1363);
nand U1053 (N_1053,In_582,In_2508);
xor U1054 (N_1054,In_2544,In_175);
nor U1055 (N_1055,In_2021,In_1783);
nor U1056 (N_1056,In_2205,In_1814);
or U1057 (N_1057,In_2591,In_538);
or U1058 (N_1058,In_1031,In_1283);
and U1059 (N_1059,In_2426,In_707);
or U1060 (N_1060,In_683,In_68);
and U1061 (N_1061,In_2220,In_194);
xor U1062 (N_1062,In_324,In_1264);
xnor U1063 (N_1063,In_215,In_2238);
or U1064 (N_1064,In_1348,In_166);
nand U1065 (N_1065,In_2999,In_1014);
or U1066 (N_1066,In_1045,In_996);
nor U1067 (N_1067,In_2682,In_2666);
nand U1068 (N_1068,In_1047,In_725);
and U1069 (N_1069,In_1158,In_2926);
and U1070 (N_1070,In_293,In_1418);
nor U1071 (N_1071,In_1846,In_2172);
or U1072 (N_1072,In_452,In_84);
xnor U1073 (N_1073,In_1552,In_2949);
and U1074 (N_1074,In_2316,In_2364);
nor U1075 (N_1075,In_1376,In_860);
and U1076 (N_1076,In_1822,In_1811);
nand U1077 (N_1077,In_2394,In_132);
and U1078 (N_1078,In_1518,In_1649);
or U1079 (N_1079,In_338,In_1060);
and U1080 (N_1080,In_659,In_2101);
and U1081 (N_1081,In_2996,In_1306);
nand U1082 (N_1082,In_2252,In_1722);
or U1083 (N_1083,In_1309,In_1680);
or U1084 (N_1084,In_1874,In_2734);
or U1085 (N_1085,In_362,In_1623);
xor U1086 (N_1086,In_289,In_879);
xnor U1087 (N_1087,In_135,In_1572);
or U1088 (N_1088,In_2066,In_1076);
or U1089 (N_1089,In_2692,In_1012);
or U1090 (N_1090,In_1643,In_327);
and U1091 (N_1091,In_41,In_1566);
xor U1092 (N_1092,In_2188,In_1001);
nor U1093 (N_1093,In_2158,In_1173);
xnor U1094 (N_1094,In_2324,In_1428);
xor U1095 (N_1095,In_2109,In_526);
nand U1096 (N_1096,In_897,In_2120);
and U1097 (N_1097,In_554,In_435);
and U1098 (N_1098,In_284,In_195);
nor U1099 (N_1099,In_2103,In_2723);
nor U1100 (N_1100,In_613,In_472);
or U1101 (N_1101,In_2992,In_1090);
nor U1102 (N_1102,In_869,In_1372);
and U1103 (N_1103,In_1725,In_372);
or U1104 (N_1104,In_2747,In_679);
nand U1105 (N_1105,In_2128,In_1789);
xor U1106 (N_1106,In_966,In_2565);
nor U1107 (N_1107,In_59,In_253);
and U1108 (N_1108,In_222,In_2494);
nand U1109 (N_1109,In_414,In_821);
xnor U1110 (N_1110,In_2961,In_768);
nor U1111 (N_1111,In_2380,In_1057);
or U1112 (N_1112,In_1307,In_2184);
and U1113 (N_1113,In_2697,In_1520);
nor U1114 (N_1114,In_595,In_2187);
nor U1115 (N_1115,In_1120,In_2687);
nand U1116 (N_1116,In_2382,In_260);
or U1117 (N_1117,In_470,In_2115);
or U1118 (N_1118,In_930,In_2919);
and U1119 (N_1119,In_1456,In_2640);
and U1120 (N_1120,In_562,In_697);
xor U1121 (N_1121,In_1301,In_1340);
xnor U1122 (N_1122,In_2365,In_2683);
nor U1123 (N_1123,In_2595,In_1499);
xor U1124 (N_1124,In_612,In_1081);
nand U1125 (N_1125,In_1026,In_907);
and U1126 (N_1126,In_528,In_506);
nand U1127 (N_1127,In_987,In_971);
and U1128 (N_1128,In_1479,In_520);
nor U1129 (N_1129,In_1671,In_88);
or U1130 (N_1130,In_2302,In_1527);
xnor U1131 (N_1131,In_2566,In_1857);
or U1132 (N_1132,In_20,In_2028);
and U1133 (N_1133,In_887,In_1122);
xor U1134 (N_1134,In_2144,In_466);
or U1135 (N_1135,In_992,In_2010);
nand U1136 (N_1136,In_2445,In_1088);
and U1137 (N_1137,In_2897,In_1327);
or U1138 (N_1138,In_564,In_2782);
or U1139 (N_1139,In_2793,In_2493);
nor U1140 (N_1140,In_439,In_1489);
and U1141 (N_1141,In_2553,In_692);
and U1142 (N_1142,In_1901,In_779);
nor U1143 (N_1143,In_2695,In_1235);
nor U1144 (N_1144,In_2796,In_1075);
xor U1145 (N_1145,In_931,In_2820);
nor U1146 (N_1146,In_2168,In_1894);
nand U1147 (N_1147,In_2062,In_2378);
or U1148 (N_1148,In_2455,In_343);
nor U1149 (N_1149,In_2232,In_2751);
nor U1150 (N_1150,In_1368,In_1632);
xnor U1151 (N_1151,In_48,In_1644);
or U1152 (N_1152,In_1596,In_789);
nand U1153 (N_1153,In_627,In_1364);
nand U1154 (N_1154,In_403,In_2716);
and U1155 (N_1155,In_643,In_1424);
and U1156 (N_1156,In_1149,In_2100);
nand U1157 (N_1157,In_1769,In_1915);
and U1158 (N_1158,In_2319,In_559);
and U1159 (N_1159,In_161,In_2913);
or U1160 (N_1160,In_2532,In_788);
nor U1161 (N_1161,In_764,In_2366);
nand U1162 (N_1162,In_2113,In_170);
nand U1163 (N_1163,In_1126,In_2581);
nand U1164 (N_1164,In_743,In_2998);
nand U1165 (N_1165,In_712,In_89);
nor U1166 (N_1166,In_2526,In_110);
nor U1167 (N_1167,In_523,In_1955);
and U1168 (N_1168,In_2475,In_1330);
nor U1169 (N_1169,In_1406,In_2283);
or U1170 (N_1170,In_1063,In_16);
nand U1171 (N_1171,In_2711,In_85);
or U1172 (N_1172,In_1827,In_241);
nand U1173 (N_1173,In_136,In_1551);
nor U1174 (N_1174,In_50,In_1312);
or U1175 (N_1175,In_497,In_363);
xor U1176 (N_1176,In_2838,In_78);
and U1177 (N_1177,In_862,In_1913);
and U1178 (N_1178,In_874,In_2655);
xor U1179 (N_1179,In_671,In_1387);
and U1180 (N_1180,In_1541,In_2392);
and U1181 (N_1181,In_989,In_2725);
xnor U1182 (N_1182,In_2908,In_657);
nand U1183 (N_1183,In_1095,In_482);
xor U1184 (N_1184,In_1050,In_2732);
xor U1185 (N_1185,In_1616,In_451);
or U1186 (N_1186,In_2685,In_2419);
and U1187 (N_1187,In_188,In_1281);
and U1188 (N_1188,In_540,In_2309);
or U1189 (N_1189,In_1341,In_2890);
and U1190 (N_1190,In_1730,In_2431);
and U1191 (N_1191,In_1134,In_2341);
or U1192 (N_1192,In_180,In_555);
and U1193 (N_1193,In_1144,In_702);
or U1194 (N_1194,In_2650,In_189);
and U1195 (N_1195,In_535,In_1168);
nand U1196 (N_1196,In_2879,In_644);
nor U1197 (N_1197,In_270,In_303);
nand U1198 (N_1198,In_522,In_1262);
and U1199 (N_1199,In_1723,In_487);
nand U1200 (N_1200,In_2673,In_660);
and U1201 (N_1201,In_332,In_676);
and U1202 (N_1202,In_288,In_2612);
or U1203 (N_1203,In_82,In_357);
and U1204 (N_1204,In_2779,In_2869);
nor U1205 (N_1205,In_832,In_489);
nor U1206 (N_1206,In_2437,In_191);
nor U1207 (N_1207,In_2235,In_1721);
nor U1208 (N_1208,In_109,In_473);
xor U1209 (N_1209,In_446,In_364);
xnor U1210 (N_1210,In_2192,In_309);
or U1211 (N_1211,In_1459,In_2329);
or U1212 (N_1212,In_2789,In_513);
or U1213 (N_1213,In_2676,In_1514);
nor U1214 (N_1214,In_67,In_1084);
xnor U1215 (N_1215,In_1024,In_1970);
and U1216 (N_1216,In_2194,In_2730);
nor U1217 (N_1217,In_1190,In_716);
xnor U1218 (N_1218,In_1465,In_894);
nand U1219 (N_1219,In_2589,In_2971);
or U1220 (N_1220,In_2058,In_2623);
nor U1221 (N_1221,In_1729,In_434);
or U1222 (N_1222,In_2819,In_409);
and U1223 (N_1223,In_1635,In_1510);
or U1224 (N_1224,In_2448,In_193);
xor U1225 (N_1225,In_1452,In_2594);
xor U1226 (N_1226,In_1463,In_2802);
and U1227 (N_1227,In_2346,In_1651);
or U1228 (N_1228,In_1752,In_2726);
xor U1229 (N_1229,In_2780,In_1708);
nor U1230 (N_1230,In_320,In_1928);
nand U1231 (N_1231,In_261,In_1881);
or U1232 (N_1232,In_2081,In_2873);
and U1233 (N_1233,In_2473,In_1493);
nor U1234 (N_1234,In_2229,In_863);
nor U1235 (N_1235,In_877,In_2149);
nor U1236 (N_1236,In_933,In_2040);
xor U1237 (N_1237,In_973,In_476);
nor U1238 (N_1238,In_2083,In_1080);
nand U1239 (N_1239,In_569,In_1253);
nand U1240 (N_1240,In_2076,In_2373);
and U1241 (N_1241,In_684,In_442);
xor U1242 (N_1242,In_1803,In_1933);
or U1243 (N_1243,In_2002,In_2481);
and U1244 (N_1244,In_936,In_1104);
xor U1245 (N_1245,In_2924,In_1314);
or U1246 (N_1246,In_455,In_1338);
or U1247 (N_1247,In_2988,In_1997);
and U1248 (N_1248,In_177,In_130);
nor U1249 (N_1249,In_1152,In_661);
xnor U1250 (N_1250,In_1599,In_1982);
nand U1251 (N_1251,In_2717,In_418);
nand U1252 (N_1252,In_1517,In_1740);
and U1253 (N_1253,In_2060,In_1565);
nand U1254 (N_1254,In_1067,In_2348);
xor U1255 (N_1255,In_2409,In_666);
nor U1256 (N_1256,In_2585,In_1268);
xnor U1257 (N_1257,In_1720,In_2173);
xor U1258 (N_1258,In_2633,In_1609);
nor U1259 (N_1259,In_1401,In_76);
nor U1260 (N_1260,In_968,In_739);
or U1261 (N_1261,In_867,In_2510);
nand U1262 (N_1262,In_65,In_822);
and U1263 (N_1263,In_2497,In_1507);
or U1264 (N_1264,In_1315,In_642);
or U1265 (N_1265,In_424,In_1938);
or U1266 (N_1266,In_1873,In_2400);
xor U1267 (N_1267,In_398,In_2447);
and U1268 (N_1268,In_462,In_590);
xnor U1269 (N_1269,In_214,In_2303);
nand U1270 (N_1270,In_2308,In_2245);
nor U1271 (N_1271,In_1129,In_1481);
or U1272 (N_1272,In_614,In_1585);
xnor U1273 (N_1273,In_2159,In_1434);
nor U1274 (N_1274,In_1603,In_2299);
xor U1275 (N_1275,In_1577,In_2755);
or U1276 (N_1276,In_1226,In_2902);
nand U1277 (N_1277,In_2160,In_2759);
xnor U1278 (N_1278,In_316,In_2936);
nor U1279 (N_1279,In_151,In_1700);
nand U1280 (N_1280,In_2857,In_1801);
xor U1281 (N_1281,In_266,In_577);
nor U1282 (N_1282,In_1323,In_43);
or U1283 (N_1283,In_2503,In_186);
and U1284 (N_1284,In_790,In_2606);
and U1285 (N_1285,In_453,In_1429);
or U1286 (N_1286,In_2330,In_2411);
nand U1287 (N_1287,In_27,In_1937);
nor U1288 (N_1288,In_458,In_1043);
nor U1289 (N_1289,In_1334,In_2007);
nor U1290 (N_1290,In_2272,In_1776);
nand U1291 (N_1291,In_843,In_1044);
and U1292 (N_1292,In_1390,In_4);
nand U1293 (N_1293,In_249,In_1478);
nor U1294 (N_1294,In_1250,In_2312);
xor U1295 (N_1295,In_2381,In_465);
nand U1296 (N_1296,In_334,In_2438);
and U1297 (N_1297,In_1228,In_2874);
nor U1298 (N_1298,In_1578,In_1380);
xnor U1299 (N_1299,In_1389,In_2707);
and U1300 (N_1300,In_1021,In_833);
and U1301 (N_1301,In_221,In_2570);
xnor U1302 (N_1302,In_118,In_691);
and U1303 (N_1303,In_1862,In_2660);
and U1304 (N_1304,In_1796,In_2901);
nand U1305 (N_1305,In_981,In_1975);
xnor U1306 (N_1306,In_2461,In_1362);
xor U1307 (N_1307,In_1650,In_2157);
and U1308 (N_1308,In_125,In_2441);
nor U1309 (N_1309,In_977,In_2817);
or U1310 (N_1310,In_2037,In_2049);
nor U1311 (N_1311,In_1036,In_903);
or U1312 (N_1312,In_236,In_772);
nand U1313 (N_1313,In_2693,In_714);
nand U1314 (N_1314,In_662,In_1029);
nand U1315 (N_1315,In_184,In_551);
and U1316 (N_1316,In_583,In_639);
and U1317 (N_1317,In_999,In_1207);
nor U1318 (N_1318,In_1621,In_2937);
and U1319 (N_1319,In_469,In_1793);
or U1320 (N_1320,In_2816,In_1973);
and U1321 (N_1321,In_29,In_2422);
nand U1322 (N_1322,In_785,In_1094);
nand U1323 (N_1323,In_2649,In_1436);
and U1324 (N_1324,In_1925,In_140);
nor U1325 (N_1325,In_1219,In_1594);
nor U1326 (N_1326,In_1950,In_2771);
and U1327 (N_1327,In_1819,In_2044);
nor U1328 (N_1328,In_500,In_2145);
nand U1329 (N_1329,In_2140,In_681);
or U1330 (N_1330,In_2618,In_1766);
xor U1331 (N_1331,In_2141,In_185);
or U1332 (N_1332,In_575,In_2853);
or U1333 (N_1333,In_1182,In_621);
and U1334 (N_1334,In_137,In_1904);
xnor U1335 (N_1335,In_2336,In_2499);
nand U1336 (N_1336,In_2266,In_2708);
and U1337 (N_1337,In_2361,In_2868);
nand U1338 (N_1338,In_259,In_1215);
xnor U1339 (N_1339,In_829,In_2093);
nor U1340 (N_1340,In_824,In_1303);
or U1341 (N_1341,In_1511,In_1506);
xor U1342 (N_1342,In_2402,In_2839);
nor U1343 (N_1343,In_1407,In_2954);
nor U1344 (N_1344,In_2554,In_2573);
nor U1345 (N_1345,In_1121,In_1176);
or U1346 (N_1346,In_2797,In_280);
or U1347 (N_1347,In_2571,In_1155);
and U1348 (N_1348,In_499,In_606);
or U1349 (N_1349,In_1391,In_1374);
xnor U1350 (N_1350,In_2736,In_1563);
or U1351 (N_1351,In_1265,In_1331);
nor U1352 (N_1352,In_1000,In_1107);
and U1353 (N_1353,In_2181,In_775);
nor U1354 (N_1354,In_311,In_884);
nand U1355 (N_1355,In_2546,In_2435);
nor U1356 (N_1356,In_2827,In_617);
nand U1357 (N_1357,In_1962,In_2806);
and U1358 (N_1358,In_250,In_2862);
and U1359 (N_1359,In_1695,In_757);
nor U1360 (N_1360,In_2884,In_1974);
nand U1361 (N_1361,In_2993,In_986);
nor U1362 (N_1362,In_1703,In_2979);
nor U1363 (N_1363,In_2960,In_2991);
nand U1364 (N_1364,In_957,In_108);
or U1365 (N_1365,In_1795,In_2427);
xor U1366 (N_1366,In_2279,In_2524);
xor U1367 (N_1367,In_885,In_1346);
or U1368 (N_1368,In_277,In_1602);
nor U1369 (N_1369,In_1386,In_416);
xnor U1370 (N_1370,In_1883,In_736);
and U1371 (N_1371,In_2460,In_1491);
and U1372 (N_1372,In_560,In_2950);
and U1373 (N_1373,In_1054,In_1991);
and U1374 (N_1374,In_1304,In_2047);
nor U1375 (N_1375,In_1214,In_663);
or U1376 (N_1376,In_2878,In_2055);
nor U1377 (N_1377,In_18,In_2865);
nor U1378 (N_1378,In_2357,In_1145);
xnor U1379 (N_1379,In_1830,In_828);
nand U1380 (N_1380,In_75,In_2823);
or U1381 (N_1381,In_1861,In_2177);
nor U1382 (N_1382,In_597,In_1419);
and U1383 (N_1383,In_1927,In_1768);
and U1384 (N_1384,In_344,In_1325);
and U1385 (N_1385,In_908,In_64);
nand U1386 (N_1386,In_570,In_2339);
nor U1387 (N_1387,In_2287,In_1791);
nor U1388 (N_1388,In_1996,In_1232);
or U1389 (N_1389,In_2686,In_233);
nand U1390 (N_1390,In_855,In_935);
or U1391 (N_1391,In_937,In_2948);
xnor U1392 (N_1392,In_51,In_1360);
nand U1393 (N_1393,In_1421,In_1762);
xor U1394 (N_1394,In_2456,In_2778);
and U1395 (N_1395,In_292,In_1055);
xor U1396 (N_1396,In_728,In_2213);
nand U1397 (N_1397,In_688,In_640);
nor U1398 (N_1398,In_1249,In_807);
nand U1399 (N_1399,In_333,In_308);
or U1400 (N_1400,In_2315,In_406);
or U1401 (N_1401,In_368,In_645);
xor U1402 (N_1402,In_658,In_2094);
xor U1403 (N_1403,In_609,In_199);
nand U1404 (N_1404,In_2406,In_2800);
or U1405 (N_1405,In_2335,In_1654);
nand U1406 (N_1406,In_2069,In_1233);
nand U1407 (N_1407,In_841,In_2713);
nor U1408 (N_1408,In_2242,In_1337);
nand U1409 (N_1409,In_1313,In_2505);
and U1410 (N_1410,In_1065,In_2799);
and U1411 (N_1411,In_1115,In_955);
or U1412 (N_1412,In_1989,In_1548);
and U1413 (N_1413,In_610,In_1195);
nand U1414 (N_1414,In_998,In_105);
xnor U1415 (N_1415,In_278,In_395);
or U1416 (N_1416,In_866,In_2084);
or U1417 (N_1417,In_784,In_1425);
nand U1418 (N_1418,In_576,In_2131);
and U1419 (N_1419,In_181,In_2691);
nor U1420 (N_1420,In_1557,In_1961);
and U1421 (N_1421,In_672,In_1194);
xor U1422 (N_1422,In_402,In_2337);
nand U1423 (N_1423,In_2176,In_876);
and U1424 (N_1424,In_1744,In_1824);
and U1425 (N_1425,In_72,In_1279);
xnor U1426 (N_1426,In_2530,In_605);
xnor U1427 (N_1427,In_2690,In_2592);
nand U1428 (N_1428,In_1847,In_1985);
and U1429 (N_1429,In_2528,In_2906);
nor U1430 (N_1430,In_83,In_2523);
xnor U1431 (N_1431,In_2314,In_2710);
nand U1432 (N_1432,In_1319,In_58);
nand U1433 (N_1433,In_2583,In_2304);
and U1434 (N_1434,In_1580,In_2534);
and U1435 (N_1435,In_2043,In_511);
xor U1436 (N_1436,In_567,In_2214);
or U1437 (N_1437,In_1246,In_793);
nor U1438 (N_1438,In_2970,In_2296);
nor U1439 (N_1439,In_388,In_2576);
or U1440 (N_1440,In_1496,In_2568);
or U1441 (N_1441,In_782,In_762);
nand U1442 (N_1442,In_207,In_1275);
nand U1443 (N_1443,In_157,In_2679);
xnor U1444 (N_1444,In_2743,In_690);
nand U1445 (N_1445,In_2121,In_2894);
or U1446 (N_1446,In_2765,In_1354);
or U1447 (N_1447,In_804,In_2254);
nor U1448 (N_1448,In_389,In_239);
or U1449 (N_1449,In_795,In_1062);
or U1450 (N_1450,In_1767,In_1701);
nand U1451 (N_1451,In_142,In_152);
and U1452 (N_1452,In_1807,In_900);
nand U1453 (N_1453,In_220,In_2852);
or U1454 (N_1454,In_2126,In_1853);
nand U1455 (N_1455,In_2189,In_61);
xnor U1456 (N_1456,In_1675,In_1365);
nor U1457 (N_1457,In_1205,In_106);
nand U1458 (N_1458,In_958,In_2170);
nand U1459 (N_1459,In_2605,In_349);
or U1460 (N_1460,In_2953,In_1976);
or U1461 (N_1461,In_216,In_861);
xor U1462 (N_1462,In_144,In_219);
nor U1463 (N_1463,In_2478,In_1016);
nand U1464 (N_1464,In_2415,In_831);
or U1465 (N_1465,In_2358,In_2997);
nand U1466 (N_1466,In_2833,In_2952);
nor U1467 (N_1467,In_172,In_66);
nand U1468 (N_1468,In_440,In_1457);
nand U1469 (N_1469,In_1083,In_54);
nand U1470 (N_1470,In_1405,In_2135);
xnor U1471 (N_1471,In_598,In_1697);
xnor U1472 (N_1472,In_198,In_896);
nand U1473 (N_1473,In_2421,In_1886);
nand U1474 (N_1474,In_1336,In_2219);
and U1475 (N_1475,In_2124,In_558);
or U1476 (N_1476,In_2206,In_2222);
and U1477 (N_1477,In_2046,In_70);
nand U1478 (N_1478,In_812,In_156);
xnor U1479 (N_1479,In_443,In_2781);
or U1480 (N_1480,In_2306,In_2648);
nand U1481 (N_1481,In_341,In_1404);
or U1482 (N_1482,In_328,In_2078);
nand U1483 (N_1483,In_1,In_711);
and U1484 (N_1484,In_2138,In_1073);
nand U1485 (N_1485,In_1646,In_573);
nand U1486 (N_1486,In_1543,In_2836);
xor U1487 (N_1487,In_2620,In_910);
nor U1488 (N_1488,In_1823,In_1484);
and U1489 (N_1489,In_1008,In_2909);
nor U1490 (N_1490,In_600,In_865);
or U1491 (N_1491,In_2096,In_1871);
nor U1492 (N_1492,In_2670,In_2844);
nor U1493 (N_1493,In_1899,In_1282);
and U1494 (N_1494,In_1969,In_1555);
nor U1495 (N_1495,In_282,In_2217);
nor U1496 (N_1496,In_549,In_766);
nor U1497 (N_1497,In_1442,In_1287);
xor U1498 (N_1498,In_735,In_1979);
xnor U1499 (N_1499,In_2372,In_1825);
and U1500 (N_1500,In_1469,In_1302);
and U1501 (N_1501,In_1916,In_42);
nor U1502 (N_1502,In_566,In_1599);
or U1503 (N_1503,In_923,In_2979);
and U1504 (N_1504,In_1278,In_2694);
and U1505 (N_1505,In_2580,In_1534);
or U1506 (N_1506,In_1504,In_2612);
or U1507 (N_1507,In_1077,In_819);
or U1508 (N_1508,In_1886,In_1604);
or U1509 (N_1509,In_1309,In_1254);
and U1510 (N_1510,In_2314,In_810);
and U1511 (N_1511,In_2400,In_2904);
and U1512 (N_1512,In_2856,In_2940);
xnor U1513 (N_1513,In_1677,In_1397);
nand U1514 (N_1514,In_569,In_277);
nor U1515 (N_1515,In_584,In_868);
and U1516 (N_1516,In_559,In_671);
or U1517 (N_1517,In_1412,In_1868);
nor U1518 (N_1518,In_636,In_1441);
nor U1519 (N_1519,In_2193,In_192);
nand U1520 (N_1520,In_2848,In_7);
xnor U1521 (N_1521,In_1735,In_2586);
and U1522 (N_1522,In_2937,In_2762);
nor U1523 (N_1523,In_1503,In_2205);
nand U1524 (N_1524,In_2537,In_1962);
nand U1525 (N_1525,In_906,In_1700);
or U1526 (N_1526,In_2160,In_1873);
or U1527 (N_1527,In_2459,In_1928);
nor U1528 (N_1528,In_1667,In_1440);
nand U1529 (N_1529,In_2178,In_2924);
nor U1530 (N_1530,In_1843,In_1317);
xor U1531 (N_1531,In_1546,In_1962);
nor U1532 (N_1532,In_2782,In_2917);
and U1533 (N_1533,In_2530,In_588);
and U1534 (N_1534,In_374,In_2990);
nand U1535 (N_1535,In_1693,In_1569);
and U1536 (N_1536,In_2677,In_657);
and U1537 (N_1537,In_466,In_706);
nor U1538 (N_1538,In_950,In_1596);
xnor U1539 (N_1539,In_298,In_993);
or U1540 (N_1540,In_991,In_1440);
or U1541 (N_1541,In_397,In_1790);
or U1542 (N_1542,In_1358,In_2962);
or U1543 (N_1543,In_671,In_607);
xor U1544 (N_1544,In_106,In_671);
or U1545 (N_1545,In_276,In_2338);
and U1546 (N_1546,In_1032,In_2829);
nor U1547 (N_1547,In_1085,In_2718);
xnor U1548 (N_1548,In_2184,In_977);
or U1549 (N_1549,In_795,In_366);
nand U1550 (N_1550,In_1701,In_1292);
or U1551 (N_1551,In_179,In_2741);
nand U1552 (N_1552,In_2738,In_1827);
and U1553 (N_1553,In_1426,In_1703);
nand U1554 (N_1554,In_241,In_478);
or U1555 (N_1555,In_2190,In_540);
nand U1556 (N_1556,In_523,In_1765);
nand U1557 (N_1557,In_2495,In_916);
and U1558 (N_1558,In_2791,In_2788);
and U1559 (N_1559,In_972,In_327);
xnor U1560 (N_1560,In_338,In_2562);
nor U1561 (N_1561,In_1366,In_2406);
nor U1562 (N_1562,In_1643,In_2068);
xor U1563 (N_1563,In_1452,In_1608);
nand U1564 (N_1564,In_532,In_2059);
or U1565 (N_1565,In_913,In_667);
xor U1566 (N_1566,In_2358,In_2627);
or U1567 (N_1567,In_398,In_1527);
nand U1568 (N_1568,In_686,In_2818);
and U1569 (N_1569,In_367,In_2175);
nor U1570 (N_1570,In_231,In_1039);
nor U1571 (N_1571,In_2020,In_295);
xnor U1572 (N_1572,In_2242,In_1834);
xnor U1573 (N_1573,In_1997,In_2528);
nand U1574 (N_1574,In_244,In_300);
xnor U1575 (N_1575,In_269,In_431);
or U1576 (N_1576,In_947,In_865);
or U1577 (N_1577,In_2846,In_646);
and U1578 (N_1578,In_1942,In_377);
and U1579 (N_1579,In_537,In_1951);
nand U1580 (N_1580,In_1700,In_1708);
nor U1581 (N_1581,In_2209,In_2693);
or U1582 (N_1582,In_1020,In_2941);
or U1583 (N_1583,In_1773,In_746);
nand U1584 (N_1584,In_388,In_85);
xor U1585 (N_1585,In_124,In_185);
or U1586 (N_1586,In_2212,In_82);
xor U1587 (N_1587,In_109,In_1484);
or U1588 (N_1588,In_1856,In_1759);
and U1589 (N_1589,In_1442,In_383);
nor U1590 (N_1590,In_2492,In_783);
nand U1591 (N_1591,In_2944,In_1183);
nor U1592 (N_1592,In_1069,In_2449);
xor U1593 (N_1593,In_2242,In_4);
and U1594 (N_1594,In_43,In_2585);
xor U1595 (N_1595,In_2532,In_1885);
nor U1596 (N_1596,In_1671,In_956);
nor U1597 (N_1597,In_986,In_2889);
and U1598 (N_1598,In_1011,In_207);
nor U1599 (N_1599,In_849,In_2912);
or U1600 (N_1600,In_976,In_2239);
xnor U1601 (N_1601,In_12,In_220);
xor U1602 (N_1602,In_243,In_2949);
nor U1603 (N_1603,In_113,In_1245);
nor U1604 (N_1604,In_245,In_840);
and U1605 (N_1605,In_2845,In_685);
nand U1606 (N_1606,In_1407,In_271);
and U1607 (N_1607,In_2952,In_2724);
and U1608 (N_1608,In_424,In_115);
nand U1609 (N_1609,In_2546,In_46);
and U1610 (N_1610,In_2600,In_2418);
nor U1611 (N_1611,In_76,In_1639);
nor U1612 (N_1612,In_2871,In_1234);
and U1613 (N_1613,In_1163,In_2855);
or U1614 (N_1614,In_1168,In_675);
or U1615 (N_1615,In_135,In_1597);
nand U1616 (N_1616,In_2878,In_1512);
nand U1617 (N_1617,In_866,In_1729);
xor U1618 (N_1618,In_1980,In_2296);
nand U1619 (N_1619,In_307,In_243);
and U1620 (N_1620,In_519,In_896);
and U1621 (N_1621,In_195,In_721);
nand U1622 (N_1622,In_2474,In_1159);
nor U1623 (N_1623,In_929,In_1287);
and U1624 (N_1624,In_2863,In_2349);
or U1625 (N_1625,In_1466,In_2089);
nor U1626 (N_1626,In_2563,In_2229);
and U1627 (N_1627,In_1272,In_1080);
nor U1628 (N_1628,In_686,In_2631);
nor U1629 (N_1629,In_1291,In_53);
nand U1630 (N_1630,In_2026,In_2652);
xor U1631 (N_1631,In_2153,In_760);
nand U1632 (N_1632,In_551,In_761);
nand U1633 (N_1633,In_2178,In_2647);
nor U1634 (N_1634,In_2785,In_0);
or U1635 (N_1635,In_701,In_576);
or U1636 (N_1636,In_1830,In_1936);
xor U1637 (N_1637,In_271,In_2794);
nand U1638 (N_1638,In_508,In_2625);
and U1639 (N_1639,In_2728,In_1675);
xor U1640 (N_1640,In_330,In_819);
nand U1641 (N_1641,In_2562,In_2714);
nor U1642 (N_1642,In_2984,In_2010);
nor U1643 (N_1643,In_2151,In_1807);
or U1644 (N_1644,In_2755,In_2206);
nand U1645 (N_1645,In_1286,In_1812);
and U1646 (N_1646,In_773,In_208);
and U1647 (N_1647,In_638,In_1482);
or U1648 (N_1648,In_1380,In_1249);
and U1649 (N_1649,In_2225,In_2198);
and U1650 (N_1650,In_1317,In_2586);
xor U1651 (N_1651,In_1973,In_2204);
xor U1652 (N_1652,In_177,In_332);
xor U1653 (N_1653,In_2546,In_1490);
or U1654 (N_1654,In_865,In_32);
and U1655 (N_1655,In_2018,In_1020);
nor U1656 (N_1656,In_2994,In_1744);
nor U1657 (N_1657,In_386,In_2684);
xor U1658 (N_1658,In_2784,In_2704);
and U1659 (N_1659,In_408,In_2329);
nor U1660 (N_1660,In_1291,In_2526);
xnor U1661 (N_1661,In_699,In_945);
xor U1662 (N_1662,In_1598,In_2342);
and U1663 (N_1663,In_493,In_2293);
xnor U1664 (N_1664,In_947,In_2060);
nor U1665 (N_1665,In_1742,In_1190);
and U1666 (N_1666,In_1866,In_660);
xnor U1667 (N_1667,In_1720,In_2852);
and U1668 (N_1668,In_1486,In_1209);
nand U1669 (N_1669,In_1440,In_1268);
nor U1670 (N_1670,In_2152,In_856);
nand U1671 (N_1671,In_2537,In_2213);
nor U1672 (N_1672,In_157,In_1027);
and U1673 (N_1673,In_2832,In_2303);
xor U1674 (N_1674,In_722,In_2973);
or U1675 (N_1675,In_398,In_1621);
and U1676 (N_1676,In_1222,In_2206);
nand U1677 (N_1677,In_733,In_2792);
or U1678 (N_1678,In_2952,In_115);
nor U1679 (N_1679,In_1255,In_2315);
and U1680 (N_1680,In_1026,In_1186);
xnor U1681 (N_1681,In_2868,In_685);
nand U1682 (N_1682,In_184,In_2483);
xor U1683 (N_1683,In_2800,In_2844);
xor U1684 (N_1684,In_2622,In_2726);
and U1685 (N_1685,In_1182,In_2617);
or U1686 (N_1686,In_1126,In_587);
or U1687 (N_1687,In_2158,In_2747);
nand U1688 (N_1688,In_2514,In_836);
xnor U1689 (N_1689,In_1411,In_1439);
nor U1690 (N_1690,In_443,In_543);
nor U1691 (N_1691,In_2883,In_1987);
or U1692 (N_1692,In_2264,In_1391);
nor U1693 (N_1693,In_2294,In_1995);
nand U1694 (N_1694,In_632,In_2158);
nor U1695 (N_1695,In_2911,In_1463);
xor U1696 (N_1696,In_2733,In_316);
xor U1697 (N_1697,In_1750,In_1363);
or U1698 (N_1698,In_1771,In_1447);
nand U1699 (N_1699,In_2836,In_2680);
or U1700 (N_1700,In_1691,In_2480);
xnor U1701 (N_1701,In_690,In_341);
and U1702 (N_1702,In_918,In_2990);
xnor U1703 (N_1703,In_913,In_5);
xor U1704 (N_1704,In_1991,In_2584);
xnor U1705 (N_1705,In_1494,In_2018);
nor U1706 (N_1706,In_1734,In_587);
nand U1707 (N_1707,In_2418,In_795);
xnor U1708 (N_1708,In_1588,In_1647);
xor U1709 (N_1709,In_1188,In_2108);
or U1710 (N_1710,In_1477,In_1337);
or U1711 (N_1711,In_778,In_498);
xnor U1712 (N_1712,In_2052,In_1810);
or U1713 (N_1713,In_2534,In_1719);
and U1714 (N_1714,In_1507,In_1717);
or U1715 (N_1715,In_1455,In_2239);
or U1716 (N_1716,In_2405,In_1582);
nand U1717 (N_1717,In_1774,In_2281);
xor U1718 (N_1718,In_1502,In_1067);
nor U1719 (N_1719,In_485,In_325);
nand U1720 (N_1720,In_1956,In_160);
and U1721 (N_1721,In_786,In_422);
nor U1722 (N_1722,In_480,In_1224);
and U1723 (N_1723,In_2388,In_1441);
nand U1724 (N_1724,In_798,In_549);
nand U1725 (N_1725,In_2765,In_1115);
xor U1726 (N_1726,In_766,In_67);
nor U1727 (N_1727,In_1491,In_2565);
xnor U1728 (N_1728,In_135,In_2148);
xnor U1729 (N_1729,In_2091,In_1053);
and U1730 (N_1730,In_1011,In_1925);
nor U1731 (N_1731,In_1211,In_328);
xnor U1732 (N_1732,In_1152,In_1902);
nand U1733 (N_1733,In_2059,In_1848);
or U1734 (N_1734,In_521,In_1786);
or U1735 (N_1735,In_2890,In_1446);
nand U1736 (N_1736,In_1393,In_2154);
nor U1737 (N_1737,In_192,In_1567);
or U1738 (N_1738,In_374,In_19);
nand U1739 (N_1739,In_2879,In_2382);
xnor U1740 (N_1740,In_823,In_2685);
xnor U1741 (N_1741,In_1626,In_2463);
or U1742 (N_1742,In_256,In_1224);
nor U1743 (N_1743,In_284,In_1810);
and U1744 (N_1744,In_188,In_541);
and U1745 (N_1745,In_2478,In_2929);
nand U1746 (N_1746,In_1243,In_2589);
and U1747 (N_1747,In_1064,In_292);
xnor U1748 (N_1748,In_2161,In_310);
xnor U1749 (N_1749,In_1255,In_545);
and U1750 (N_1750,In_1911,In_2746);
nor U1751 (N_1751,In_1043,In_435);
and U1752 (N_1752,In_167,In_1218);
nor U1753 (N_1753,In_2527,In_2880);
or U1754 (N_1754,In_1592,In_444);
nand U1755 (N_1755,In_1146,In_776);
or U1756 (N_1756,In_2991,In_1821);
or U1757 (N_1757,In_665,In_2623);
xnor U1758 (N_1758,In_2670,In_1711);
nand U1759 (N_1759,In_1860,In_493);
nor U1760 (N_1760,In_1124,In_2944);
or U1761 (N_1761,In_1345,In_2140);
nor U1762 (N_1762,In_2858,In_1218);
xnor U1763 (N_1763,In_568,In_2867);
nand U1764 (N_1764,In_149,In_2134);
or U1765 (N_1765,In_2085,In_129);
or U1766 (N_1766,In_1090,In_327);
nor U1767 (N_1767,In_570,In_728);
and U1768 (N_1768,In_1477,In_477);
or U1769 (N_1769,In_1590,In_843);
nand U1770 (N_1770,In_2883,In_2822);
xor U1771 (N_1771,In_1542,In_2413);
and U1772 (N_1772,In_1706,In_587);
and U1773 (N_1773,In_223,In_483);
nor U1774 (N_1774,In_1878,In_2484);
nand U1775 (N_1775,In_2814,In_641);
nand U1776 (N_1776,In_1735,In_1591);
nor U1777 (N_1777,In_552,In_2046);
nand U1778 (N_1778,In_126,In_1469);
and U1779 (N_1779,In_932,In_1892);
or U1780 (N_1780,In_1443,In_1232);
or U1781 (N_1781,In_850,In_1458);
xor U1782 (N_1782,In_664,In_1024);
and U1783 (N_1783,In_376,In_2048);
nor U1784 (N_1784,In_144,In_1564);
nor U1785 (N_1785,In_2996,In_2448);
nand U1786 (N_1786,In_2449,In_432);
nand U1787 (N_1787,In_1606,In_1682);
and U1788 (N_1788,In_2580,In_2815);
nand U1789 (N_1789,In_803,In_2823);
xor U1790 (N_1790,In_2031,In_1767);
or U1791 (N_1791,In_2434,In_1108);
and U1792 (N_1792,In_2948,In_889);
xor U1793 (N_1793,In_961,In_2930);
nand U1794 (N_1794,In_2598,In_2245);
nor U1795 (N_1795,In_731,In_936);
or U1796 (N_1796,In_1421,In_1085);
nand U1797 (N_1797,In_2302,In_2458);
xor U1798 (N_1798,In_27,In_1426);
and U1799 (N_1799,In_1303,In_1251);
or U1800 (N_1800,In_2232,In_862);
or U1801 (N_1801,In_855,In_1576);
or U1802 (N_1802,In_143,In_2397);
xor U1803 (N_1803,In_2162,In_974);
nand U1804 (N_1804,In_2188,In_1081);
or U1805 (N_1805,In_855,In_2838);
nand U1806 (N_1806,In_1288,In_1685);
nor U1807 (N_1807,In_1161,In_584);
nand U1808 (N_1808,In_1743,In_1947);
nand U1809 (N_1809,In_2220,In_1254);
or U1810 (N_1810,In_2452,In_2265);
and U1811 (N_1811,In_1609,In_2871);
nor U1812 (N_1812,In_472,In_2881);
nor U1813 (N_1813,In_1615,In_2967);
or U1814 (N_1814,In_2459,In_424);
xnor U1815 (N_1815,In_290,In_1737);
and U1816 (N_1816,In_2856,In_1025);
or U1817 (N_1817,In_2962,In_1451);
nor U1818 (N_1818,In_596,In_1076);
xnor U1819 (N_1819,In_440,In_1283);
or U1820 (N_1820,In_2082,In_2657);
xnor U1821 (N_1821,In_1415,In_1675);
nor U1822 (N_1822,In_2355,In_2635);
nor U1823 (N_1823,In_2263,In_1100);
or U1824 (N_1824,In_624,In_677);
xor U1825 (N_1825,In_2165,In_1559);
nand U1826 (N_1826,In_276,In_294);
nor U1827 (N_1827,In_2648,In_2579);
nand U1828 (N_1828,In_505,In_133);
or U1829 (N_1829,In_288,In_2703);
nand U1830 (N_1830,In_689,In_2668);
nand U1831 (N_1831,In_2306,In_449);
nor U1832 (N_1832,In_1115,In_2375);
and U1833 (N_1833,In_1353,In_2005);
and U1834 (N_1834,In_220,In_576);
nand U1835 (N_1835,In_2905,In_1832);
nand U1836 (N_1836,In_1930,In_2403);
or U1837 (N_1837,In_1226,In_1180);
xor U1838 (N_1838,In_260,In_1377);
or U1839 (N_1839,In_2475,In_2478);
nor U1840 (N_1840,In_1357,In_2033);
and U1841 (N_1841,In_2014,In_1498);
nand U1842 (N_1842,In_1826,In_2033);
nand U1843 (N_1843,In_2300,In_662);
nand U1844 (N_1844,In_2928,In_2587);
nand U1845 (N_1845,In_2488,In_1034);
and U1846 (N_1846,In_646,In_2110);
or U1847 (N_1847,In_1158,In_466);
xor U1848 (N_1848,In_2275,In_316);
nand U1849 (N_1849,In_2695,In_1237);
xnor U1850 (N_1850,In_2946,In_2533);
or U1851 (N_1851,In_306,In_1015);
nor U1852 (N_1852,In_2064,In_2000);
nand U1853 (N_1853,In_2606,In_2290);
and U1854 (N_1854,In_657,In_2310);
or U1855 (N_1855,In_2213,In_2004);
or U1856 (N_1856,In_1500,In_1705);
and U1857 (N_1857,In_809,In_335);
or U1858 (N_1858,In_1783,In_803);
or U1859 (N_1859,In_342,In_1062);
nand U1860 (N_1860,In_2589,In_151);
nor U1861 (N_1861,In_614,In_1138);
and U1862 (N_1862,In_1003,In_347);
nor U1863 (N_1863,In_111,In_108);
nor U1864 (N_1864,In_1668,In_2699);
and U1865 (N_1865,In_2094,In_1240);
and U1866 (N_1866,In_400,In_2572);
nand U1867 (N_1867,In_36,In_2290);
and U1868 (N_1868,In_2484,In_625);
xor U1869 (N_1869,In_1919,In_2569);
and U1870 (N_1870,In_2901,In_1607);
nor U1871 (N_1871,In_1994,In_840);
nand U1872 (N_1872,In_1737,In_36);
xnor U1873 (N_1873,In_2331,In_2324);
nand U1874 (N_1874,In_2072,In_2661);
or U1875 (N_1875,In_990,In_1497);
nor U1876 (N_1876,In_1947,In_599);
or U1877 (N_1877,In_2052,In_2221);
xor U1878 (N_1878,In_2014,In_2287);
nand U1879 (N_1879,In_1061,In_1423);
nand U1880 (N_1880,In_496,In_2779);
xnor U1881 (N_1881,In_2703,In_667);
or U1882 (N_1882,In_1216,In_2848);
xnor U1883 (N_1883,In_1758,In_2026);
nand U1884 (N_1884,In_2235,In_2286);
or U1885 (N_1885,In_1135,In_532);
or U1886 (N_1886,In_305,In_2027);
or U1887 (N_1887,In_697,In_2104);
and U1888 (N_1888,In_1349,In_2931);
nand U1889 (N_1889,In_2306,In_1273);
and U1890 (N_1890,In_2353,In_1981);
nand U1891 (N_1891,In_466,In_2175);
or U1892 (N_1892,In_2696,In_1621);
nor U1893 (N_1893,In_2964,In_1039);
and U1894 (N_1894,In_908,In_1216);
nand U1895 (N_1895,In_1148,In_269);
nand U1896 (N_1896,In_1098,In_1307);
or U1897 (N_1897,In_1490,In_943);
or U1898 (N_1898,In_501,In_2521);
or U1899 (N_1899,In_2236,In_2148);
xor U1900 (N_1900,In_1318,In_1550);
or U1901 (N_1901,In_2029,In_1979);
or U1902 (N_1902,In_1891,In_2896);
xnor U1903 (N_1903,In_600,In_438);
xnor U1904 (N_1904,In_393,In_1577);
and U1905 (N_1905,In_487,In_1960);
nand U1906 (N_1906,In_1886,In_741);
and U1907 (N_1907,In_1212,In_5);
and U1908 (N_1908,In_836,In_2139);
nand U1909 (N_1909,In_849,In_1200);
or U1910 (N_1910,In_2356,In_41);
xnor U1911 (N_1911,In_518,In_729);
or U1912 (N_1912,In_2236,In_2);
nor U1913 (N_1913,In_2356,In_1113);
or U1914 (N_1914,In_1140,In_980);
nand U1915 (N_1915,In_762,In_1334);
nand U1916 (N_1916,In_2033,In_1467);
nand U1917 (N_1917,In_2092,In_1014);
xnor U1918 (N_1918,In_2216,In_2935);
xor U1919 (N_1919,In_1054,In_965);
xnor U1920 (N_1920,In_1818,In_2208);
xor U1921 (N_1921,In_1228,In_1926);
and U1922 (N_1922,In_1089,In_648);
and U1923 (N_1923,In_2929,In_1674);
and U1924 (N_1924,In_756,In_1689);
and U1925 (N_1925,In_1252,In_2247);
xnor U1926 (N_1926,In_1064,In_1296);
nor U1927 (N_1927,In_2879,In_1024);
nand U1928 (N_1928,In_1066,In_2761);
nand U1929 (N_1929,In_904,In_540);
nand U1930 (N_1930,In_2892,In_565);
nor U1931 (N_1931,In_501,In_1778);
or U1932 (N_1932,In_2512,In_779);
nand U1933 (N_1933,In_1193,In_1340);
or U1934 (N_1934,In_1453,In_2379);
or U1935 (N_1935,In_1332,In_492);
xnor U1936 (N_1936,In_836,In_1214);
nand U1937 (N_1937,In_1962,In_70);
and U1938 (N_1938,In_380,In_2898);
xor U1939 (N_1939,In_732,In_1244);
xor U1940 (N_1940,In_1212,In_2220);
nand U1941 (N_1941,In_1875,In_2116);
xnor U1942 (N_1942,In_966,In_2328);
nor U1943 (N_1943,In_1133,In_1042);
xor U1944 (N_1944,In_1750,In_1786);
nor U1945 (N_1945,In_2902,In_1116);
or U1946 (N_1946,In_823,In_1745);
nor U1947 (N_1947,In_596,In_2573);
nor U1948 (N_1948,In_1999,In_1544);
or U1949 (N_1949,In_2339,In_106);
nand U1950 (N_1950,In_1775,In_2422);
or U1951 (N_1951,In_1399,In_799);
and U1952 (N_1952,In_662,In_1448);
xor U1953 (N_1953,In_759,In_219);
nand U1954 (N_1954,In_592,In_309);
and U1955 (N_1955,In_1786,In_2274);
xnor U1956 (N_1956,In_395,In_2837);
nor U1957 (N_1957,In_2852,In_2677);
nand U1958 (N_1958,In_551,In_1523);
nand U1959 (N_1959,In_1839,In_529);
nor U1960 (N_1960,In_1701,In_157);
nor U1961 (N_1961,In_1514,In_1359);
or U1962 (N_1962,In_2417,In_1184);
xor U1963 (N_1963,In_2129,In_1427);
or U1964 (N_1964,In_314,In_1745);
nor U1965 (N_1965,In_1427,In_8);
xnor U1966 (N_1966,In_2099,In_1345);
nor U1967 (N_1967,In_2608,In_643);
and U1968 (N_1968,In_1276,In_2239);
nor U1969 (N_1969,In_1850,In_1267);
and U1970 (N_1970,In_2941,In_1208);
nand U1971 (N_1971,In_1964,In_2059);
xnor U1972 (N_1972,In_188,In_2450);
nand U1973 (N_1973,In_647,In_1764);
xor U1974 (N_1974,In_314,In_2638);
xnor U1975 (N_1975,In_2257,In_1893);
nand U1976 (N_1976,In_277,In_2793);
or U1977 (N_1977,In_1378,In_2904);
nor U1978 (N_1978,In_242,In_112);
or U1979 (N_1979,In_2747,In_5);
or U1980 (N_1980,In_767,In_2081);
nand U1981 (N_1981,In_2054,In_263);
or U1982 (N_1982,In_1883,In_853);
xnor U1983 (N_1983,In_1561,In_1791);
or U1984 (N_1984,In_797,In_1099);
nor U1985 (N_1985,In_671,In_2370);
xor U1986 (N_1986,In_1023,In_1751);
or U1987 (N_1987,In_751,In_2448);
nor U1988 (N_1988,In_2753,In_1264);
xnor U1989 (N_1989,In_1856,In_1840);
nor U1990 (N_1990,In_2697,In_39);
nor U1991 (N_1991,In_2784,In_400);
nor U1992 (N_1992,In_232,In_970);
nand U1993 (N_1993,In_2592,In_691);
xor U1994 (N_1994,In_1218,In_977);
xor U1995 (N_1995,In_2213,In_1879);
nor U1996 (N_1996,In_2673,In_224);
and U1997 (N_1997,In_2137,In_1301);
nand U1998 (N_1998,In_927,In_755);
and U1999 (N_1999,In_2829,In_1459);
or U2000 (N_2000,In_471,In_2124);
xnor U2001 (N_2001,In_1160,In_2704);
xor U2002 (N_2002,In_1748,In_872);
xor U2003 (N_2003,In_2453,In_801);
nor U2004 (N_2004,In_1945,In_2584);
and U2005 (N_2005,In_1049,In_2827);
and U2006 (N_2006,In_1943,In_1888);
or U2007 (N_2007,In_2967,In_1521);
and U2008 (N_2008,In_736,In_161);
nor U2009 (N_2009,In_646,In_29);
and U2010 (N_2010,In_1538,In_52);
or U2011 (N_2011,In_378,In_1204);
nand U2012 (N_2012,In_449,In_796);
xor U2013 (N_2013,In_678,In_44);
xnor U2014 (N_2014,In_983,In_2660);
nor U2015 (N_2015,In_1466,In_1567);
nand U2016 (N_2016,In_2140,In_958);
and U2017 (N_2017,In_1420,In_820);
nand U2018 (N_2018,In_2921,In_1244);
nand U2019 (N_2019,In_1893,In_2276);
xor U2020 (N_2020,In_2757,In_704);
or U2021 (N_2021,In_2961,In_2255);
nor U2022 (N_2022,In_1680,In_2509);
nand U2023 (N_2023,In_2803,In_2408);
or U2024 (N_2024,In_2663,In_2732);
xor U2025 (N_2025,In_1597,In_2035);
or U2026 (N_2026,In_389,In_2978);
and U2027 (N_2027,In_2418,In_2713);
xnor U2028 (N_2028,In_1426,In_2963);
or U2029 (N_2029,In_1286,In_1700);
nand U2030 (N_2030,In_374,In_89);
nand U2031 (N_2031,In_736,In_1434);
nand U2032 (N_2032,In_107,In_42);
and U2033 (N_2033,In_1713,In_208);
nor U2034 (N_2034,In_1623,In_709);
or U2035 (N_2035,In_1437,In_1318);
and U2036 (N_2036,In_1438,In_609);
xnor U2037 (N_2037,In_1590,In_2861);
or U2038 (N_2038,In_1520,In_1534);
and U2039 (N_2039,In_2035,In_243);
or U2040 (N_2040,In_1142,In_1698);
and U2041 (N_2041,In_1766,In_1504);
or U2042 (N_2042,In_817,In_387);
and U2043 (N_2043,In_1535,In_908);
nand U2044 (N_2044,In_803,In_747);
or U2045 (N_2045,In_1506,In_1923);
xnor U2046 (N_2046,In_939,In_1817);
or U2047 (N_2047,In_824,In_1084);
nand U2048 (N_2048,In_1252,In_2891);
xor U2049 (N_2049,In_2865,In_2642);
nor U2050 (N_2050,In_2433,In_1202);
or U2051 (N_2051,In_2237,In_110);
nand U2052 (N_2052,In_2239,In_1226);
nand U2053 (N_2053,In_2409,In_812);
or U2054 (N_2054,In_981,In_1453);
and U2055 (N_2055,In_1309,In_89);
xnor U2056 (N_2056,In_1070,In_1780);
xnor U2057 (N_2057,In_1895,In_261);
nand U2058 (N_2058,In_2122,In_2778);
nor U2059 (N_2059,In_50,In_2995);
nor U2060 (N_2060,In_662,In_395);
and U2061 (N_2061,In_42,In_2276);
xnor U2062 (N_2062,In_591,In_2297);
xnor U2063 (N_2063,In_153,In_1049);
or U2064 (N_2064,In_1592,In_120);
xnor U2065 (N_2065,In_1058,In_500);
nor U2066 (N_2066,In_2277,In_2993);
nand U2067 (N_2067,In_2215,In_1408);
nor U2068 (N_2068,In_571,In_1695);
nand U2069 (N_2069,In_887,In_2530);
and U2070 (N_2070,In_93,In_2469);
nor U2071 (N_2071,In_960,In_239);
or U2072 (N_2072,In_683,In_1296);
nand U2073 (N_2073,In_2963,In_1881);
xor U2074 (N_2074,In_2180,In_2913);
nor U2075 (N_2075,In_922,In_2245);
or U2076 (N_2076,In_964,In_2684);
and U2077 (N_2077,In_1444,In_481);
nor U2078 (N_2078,In_1877,In_2879);
or U2079 (N_2079,In_1283,In_2050);
or U2080 (N_2080,In_1608,In_2809);
xnor U2081 (N_2081,In_113,In_1473);
and U2082 (N_2082,In_952,In_65);
xor U2083 (N_2083,In_1577,In_2047);
and U2084 (N_2084,In_2746,In_1204);
nor U2085 (N_2085,In_856,In_1550);
xor U2086 (N_2086,In_2896,In_1602);
and U2087 (N_2087,In_1338,In_135);
or U2088 (N_2088,In_1098,In_1377);
xor U2089 (N_2089,In_754,In_2523);
nand U2090 (N_2090,In_2129,In_1574);
xor U2091 (N_2091,In_269,In_2782);
nand U2092 (N_2092,In_2085,In_1723);
or U2093 (N_2093,In_788,In_1);
or U2094 (N_2094,In_283,In_379);
nand U2095 (N_2095,In_2417,In_784);
and U2096 (N_2096,In_2325,In_777);
nand U2097 (N_2097,In_1412,In_1251);
or U2098 (N_2098,In_2986,In_2648);
and U2099 (N_2099,In_382,In_894);
nand U2100 (N_2100,In_607,In_2864);
or U2101 (N_2101,In_2106,In_2101);
and U2102 (N_2102,In_1437,In_901);
or U2103 (N_2103,In_1136,In_2477);
or U2104 (N_2104,In_949,In_2547);
nor U2105 (N_2105,In_796,In_2778);
and U2106 (N_2106,In_1660,In_1467);
and U2107 (N_2107,In_2646,In_1208);
or U2108 (N_2108,In_534,In_1861);
nand U2109 (N_2109,In_77,In_1503);
or U2110 (N_2110,In_2438,In_1260);
nor U2111 (N_2111,In_177,In_1580);
or U2112 (N_2112,In_2280,In_1048);
nor U2113 (N_2113,In_358,In_1570);
nand U2114 (N_2114,In_1376,In_2802);
or U2115 (N_2115,In_1511,In_104);
and U2116 (N_2116,In_1779,In_2267);
and U2117 (N_2117,In_2828,In_1913);
nor U2118 (N_2118,In_2254,In_1985);
and U2119 (N_2119,In_2540,In_2311);
nor U2120 (N_2120,In_2579,In_1466);
nor U2121 (N_2121,In_322,In_2584);
or U2122 (N_2122,In_549,In_838);
nand U2123 (N_2123,In_2967,In_2742);
nor U2124 (N_2124,In_964,In_2968);
or U2125 (N_2125,In_1708,In_366);
nor U2126 (N_2126,In_1556,In_1628);
or U2127 (N_2127,In_2636,In_1172);
xnor U2128 (N_2128,In_310,In_1907);
nand U2129 (N_2129,In_2422,In_476);
or U2130 (N_2130,In_2460,In_1267);
nor U2131 (N_2131,In_35,In_2034);
xnor U2132 (N_2132,In_918,In_1055);
nor U2133 (N_2133,In_1234,In_267);
xnor U2134 (N_2134,In_2505,In_1273);
nor U2135 (N_2135,In_2187,In_1861);
or U2136 (N_2136,In_2110,In_1490);
xor U2137 (N_2137,In_1953,In_63);
nor U2138 (N_2138,In_1971,In_2098);
xor U2139 (N_2139,In_289,In_1183);
xnor U2140 (N_2140,In_1112,In_2158);
nor U2141 (N_2141,In_2192,In_407);
and U2142 (N_2142,In_1969,In_1395);
nor U2143 (N_2143,In_244,In_923);
xor U2144 (N_2144,In_1081,In_2349);
or U2145 (N_2145,In_1954,In_2398);
and U2146 (N_2146,In_2074,In_2218);
and U2147 (N_2147,In_2634,In_46);
and U2148 (N_2148,In_2824,In_1771);
or U2149 (N_2149,In_900,In_977);
nand U2150 (N_2150,In_1290,In_394);
nor U2151 (N_2151,In_2515,In_342);
nand U2152 (N_2152,In_833,In_501);
or U2153 (N_2153,In_2073,In_2458);
or U2154 (N_2154,In_2726,In_2533);
and U2155 (N_2155,In_2193,In_713);
nor U2156 (N_2156,In_1982,In_1050);
xor U2157 (N_2157,In_2947,In_2205);
nand U2158 (N_2158,In_902,In_2622);
xnor U2159 (N_2159,In_2606,In_660);
nand U2160 (N_2160,In_1782,In_436);
nand U2161 (N_2161,In_1283,In_1458);
nand U2162 (N_2162,In_2098,In_380);
nor U2163 (N_2163,In_2983,In_593);
xnor U2164 (N_2164,In_134,In_2704);
nor U2165 (N_2165,In_1608,In_969);
or U2166 (N_2166,In_2195,In_1021);
xor U2167 (N_2167,In_1809,In_154);
nor U2168 (N_2168,In_1587,In_1997);
and U2169 (N_2169,In_1676,In_2254);
or U2170 (N_2170,In_682,In_493);
and U2171 (N_2171,In_27,In_1047);
or U2172 (N_2172,In_1426,In_2603);
or U2173 (N_2173,In_2435,In_547);
xnor U2174 (N_2174,In_2205,In_92);
nand U2175 (N_2175,In_2331,In_1574);
and U2176 (N_2176,In_707,In_391);
and U2177 (N_2177,In_2253,In_1093);
xor U2178 (N_2178,In_2509,In_371);
nor U2179 (N_2179,In_535,In_133);
and U2180 (N_2180,In_2747,In_601);
nand U2181 (N_2181,In_1815,In_364);
or U2182 (N_2182,In_874,In_2324);
xor U2183 (N_2183,In_798,In_1696);
xnor U2184 (N_2184,In_131,In_1854);
xor U2185 (N_2185,In_2487,In_2337);
xnor U2186 (N_2186,In_1548,In_613);
nor U2187 (N_2187,In_2015,In_2411);
nor U2188 (N_2188,In_449,In_313);
nand U2189 (N_2189,In_2347,In_2715);
nor U2190 (N_2190,In_2037,In_630);
nand U2191 (N_2191,In_1496,In_1273);
xnor U2192 (N_2192,In_2263,In_2693);
nand U2193 (N_2193,In_1487,In_701);
and U2194 (N_2194,In_1687,In_2184);
nor U2195 (N_2195,In_632,In_526);
or U2196 (N_2196,In_2037,In_119);
and U2197 (N_2197,In_400,In_1287);
nor U2198 (N_2198,In_412,In_2117);
nor U2199 (N_2199,In_689,In_1182);
or U2200 (N_2200,In_1684,In_850);
xor U2201 (N_2201,In_970,In_80);
and U2202 (N_2202,In_2097,In_268);
and U2203 (N_2203,In_1621,In_1094);
and U2204 (N_2204,In_1333,In_1826);
nor U2205 (N_2205,In_651,In_70);
xnor U2206 (N_2206,In_1935,In_692);
xnor U2207 (N_2207,In_1604,In_1141);
or U2208 (N_2208,In_2821,In_2756);
nand U2209 (N_2209,In_2239,In_1174);
and U2210 (N_2210,In_1158,In_2639);
and U2211 (N_2211,In_1174,In_1625);
nand U2212 (N_2212,In_2499,In_2192);
and U2213 (N_2213,In_1475,In_1735);
and U2214 (N_2214,In_667,In_593);
or U2215 (N_2215,In_1351,In_1021);
xor U2216 (N_2216,In_2465,In_1676);
and U2217 (N_2217,In_116,In_2187);
and U2218 (N_2218,In_1587,In_996);
nor U2219 (N_2219,In_2729,In_1351);
nand U2220 (N_2220,In_1088,In_1037);
nand U2221 (N_2221,In_1280,In_2640);
nand U2222 (N_2222,In_2573,In_2430);
nand U2223 (N_2223,In_594,In_1184);
or U2224 (N_2224,In_2248,In_2126);
or U2225 (N_2225,In_1809,In_1605);
nor U2226 (N_2226,In_972,In_224);
nand U2227 (N_2227,In_883,In_203);
nand U2228 (N_2228,In_428,In_2131);
or U2229 (N_2229,In_1298,In_773);
or U2230 (N_2230,In_2312,In_1675);
nor U2231 (N_2231,In_84,In_2980);
xor U2232 (N_2232,In_2786,In_2970);
or U2233 (N_2233,In_543,In_85);
and U2234 (N_2234,In_1525,In_2603);
xor U2235 (N_2235,In_200,In_1766);
and U2236 (N_2236,In_965,In_1672);
nor U2237 (N_2237,In_2420,In_2780);
xor U2238 (N_2238,In_2571,In_766);
or U2239 (N_2239,In_682,In_604);
xnor U2240 (N_2240,In_1681,In_1662);
or U2241 (N_2241,In_1102,In_1879);
nand U2242 (N_2242,In_1056,In_577);
and U2243 (N_2243,In_2267,In_1185);
nand U2244 (N_2244,In_166,In_1017);
or U2245 (N_2245,In_1818,In_15);
xor U2246 (N_2246,In_1140,In_1981);
nor U2247 (N_2247,In_1297,In_2492);
and U2248 (N_2248,In_2103,In_2816);
nor U2249 (N_2249,In_888,In_1375);
and U2250 (N_2250,In_2545,In_2100);
or U2251 (N_2251,In_950,In_649);
or U2252 (N_2252,In_2128,In_1860);
and U2253 (N_2253,In_263,In_1330);
nor U2254 (N_2254,In_2194,In_1958);
xnor U2255 (N_2255,In_840,In_2674);
or U2256 (N_2256,In_2617,In_1943);
and U2257 (N_2257,In_60,In_2065);
nor U2258 (N_2258,In_2488,In_1000);
xnor U2259 (N_2259,In_2701,In_1305);
nand U2260 (N_2260,In_2157,In_108);
xnor U2261 (N_2261,In_516,In_2671);
nor U2262 (N_2262,In_330,In_1508);
or U2263 (N_2263,In_2441,In_2419);
nor U2264 (N_2264,In_675,In_334);
or U2265 (N_2265,In_315,In_2164);
or U2266 (N_2266,In_1980,In_1347);
or U2267 (N_2267,In_2909,In_2394);
and U2268 (N_2268,In_1340,In_2948);
nand U2269 (N_2269,In_191,In_1315);
nand U2270 (N_2270,In_1334,In_1973);
xnor U2271 (N_2271,In_739,In_1056);
or U2272 (N_2272,In_2317,In_619);
xor U2273 (N_2273,In_1966,In_1279);
or U2274 (N_2274,In_2893,In_1021);
and U2275 (N_2275,In_1757,In_993);
or U2276 (N_2276,In_989,In_1589);
xnor U2277 (N_2277,In_2740,In_1660);
and U2278 (N_2278,In_931,In_1576);
nor U2279 (N_2279,In_1021,In_2344);
nor U2280 (N_2280,In_1518,In_460);
and U2281 (N_2281,In_1707,In_166);
nor U2282 (N_2282,In_2214,In_170);
nor U2283 (N_2283,In_1922,In_2489);
nor U2284 (N_2284,In_2094,In_2793);
and U2285 (N_2285,In_250,In_2062);
nand U2286 (N_2286,In_2398,In_2432);
nor U2287 (N_2287,In_2992,In_1093);
nor U2288 (N_2288,In_303,In_1005);
or U2289 (N_2289,In_1831,In_1546);
xor U2290 (N_2290,In_2336,In_139);
xor U2291 (N_2291,In_330,In_404);
or U2292 (N_2292,In_2296,In_626);
xor U2293 (N_2293,In_1597,In_2606);
or U2294 (N_2294,In_144,In_2699);
nor U2295 (N_2295,In_501,In_1614);
xor U2296 (N_2296,In_293,In_1220);
nor U2297 (N_2297,In_1810,In_892);
and U2298 (N_2298,In_1909,In_1088);
and U2299 (N_2299,In_1489,In_2286);
nand U2300 (N_2300,In_2010,In_1496);
nand U2301 (N_2301,In_738,In_1870);
nand U2302 (N_2302,In_1201,In_2092);
xnor U2303 (N_2303,In_191,In_1436);
xor U2304 (N_2304,In_2031,In_462);
or U2305 (N_2305,In_626,In_642);
nor U2306 (N_2306,In_1508,In_873);
nand U2307 (N_2307,In_2013,In_870);
and U2308 (N_2308,In_2219,In_1109);
or U2309 (N_2309,In_1189,In_1263);
nand U2310 (N_2310,In_1695,In_168);
xor U2311 (N_2311,In_2316,In_1015);
and U2312 (N_2312,In_2862,In_821);
nor U2313 (N_2313,In_2941,In_1416);
or U2314 (N_2314,In_133,In_618);
nor U2315 (N_2315,In_1161,In_536);
and U2316 (N_2316,In_658,In_866);
or U2317 (N_2317,In_669,In_734);
nand U2318 (N_2318,In_1994,In_96);
xnor U2319 (N_2319,In_1187,In_988);
nand U2320 (N_2320,In_2551,In_2750);
xor U2321 (N_2321,In_610,In_802);
and U2322 (N_2322,In_2818,In_264);
or U2323 (N_2323,In_389,In_1778);
nor U2324 (N_2324,In_2158,In_1507);
or U2325 (N_2325,In_1972,In_2015);
nand U2326 (N_2326,In_64,In_802);
xor U2327 (N_2327,In_1906,In_2927);
and U2328 (N_2328,In_1285,In_2090);
and U2329 (N_2329,In_1969,In_750);
or U2330 (N_2330,In_2815,In_2131);
or U2331 (N_2331,In_2479,In_2755);
nand U2332 (N_2332,In_2708,In_2010);
or U2333 (N_2333,In_1577,In_799);
or U2334 (N_2334,In_540,In_2877);
nor U2335 (N_2335,In_246,In_53);
and U2336 (N_2336,In_495,In_2906);
nand U2337 (N_2337,In_292,In_1050);
nor U2338 (N_2338,In_1012,In_1446);
nor U2339 (N_2339,In_1652,In_1404);
nor U2340 (N_2340,In_1137,In_1962);
xnor U2341 (N_2341,In_2083,In_793);
and U2342 (N_2342,In_1725,In_1435);
or U2343 (N_2343,In_2938,In_1013);
nor U2344 (N_2344,In_758,In_367);
nand U2345 (N_2345,In_2341,In_1662);
nand U2346 (N_2346,In_61,In_1421);
nand U2347 (N_2347,In_2681,In_2318);
or U2348 (N_2348,In_1081,In_885);
nor U2349 (N_2349,In_562,In_1468);
nor U2350 (N_2350,In_1125,In_1658);
nand U2351 (N_2351,In_1779,In_320);
or U2352 (N_2352,In_1699,In_1835);
nand U2353 (N_2353,In_790,In_894);
xnor U2354 (N_2354,In_1159,In_506);
and U2355 (N_2355,In_2862,In_1980);
and U2356 (N_2356,In_2485,In_394);
and U2357 (N_2357,In_202,In_2122);
xnor U2358 (N_2358,In_1218,In_2250);
nand U2359 (N_2359,In_1498,In_1593);
nor U2360 (N_2360,In_2771,In_955);
or U2361 (N_2361,In_2874,In_2289);
or U2362 (N_2362,In_1590,In_2507);
or U2363 (N_2363,In_2682,In_1430);
nand U2364 (N_2364,In_1628,In_211);
xnor U2365 (N_2365,In_50,In_567);
and U2366 (N_2366,In_1679,In_2205);
nand U2367 (N_2367,In_2234,In_870);
xor U2368 (N_2368,In_67,In_525);
or U2369 (N_2369,In_770,In_779);
xnor U2370 (N_2370,In_2242,In_1459);
or U2371 (N_2371,In_1669,In_2023);
or U2372 (N_2372,In_754,In_79);
nor U2373 (N_2373,In_1212,In_927);
or U2374 (N_2374,In_438,In_2513);
nor U2375 (N_2375,In_2347,In_7);
and U2376 (N_2376,In_2394,In_944);
xnor U2377 (N_2377,In_1049,In_1018);
or U2378 (N_2378,In_756,In_2102);
nand U2379 (N_2379,In_2133,In_2875);
xor U2380 (N_2380,In_501,In_2509);
nand U2381 (N_2381,In_417,In_1088);
and U2382 (N_2382,In_584,In_1155);
xnor U2383 (N_2383,In_88,In_2764);
nor U2384 (N_2384,In_1024,In_986);
xor U2385 (N_2385,In_1616,In_2445);
and U2386 (N_2386,In_1049,In_149);
nand U2387 (N_2387,In_2829,In_2834);
nor U2388 (N_2388,In_153,In_2627);
xnor U2389 (N_2389,In_1560,In_670);
nand U2390 (N_2390,In_691,In_2541);
or U2391 (N_2391,In_442,In_2833);
and U2392 (N_2392,In_2224,In_2503);
and U2393 (N_2393,In_1523,In_1310);
and U2394 (N_2394,In_2494,In_417);
nand U2395 (N_2395,In_2679,In_2293);
or U2396 (N_2396,In_942,In_1810);
nor U2397 (N_2397,In_2660,In_764);
nand U2398 (N_2398,In_2487,In_2901);
and U2399 (N_2399,In_2563,In_1179);
and U2400 (N_2400,In_1246,In_1405);
and U2401 (N_2401,In_1851,In_811);
or U2402 (N_2402,In_2675,In_2915);
xnor U2403 (N_2403,In_1405,In_912);
and U2404 (N_2404,In_1019,In_1065);
and U2405 (N_2405,In_2954,In_2858);
and U2406 (N_2406,In_200,In_2866);
nor U2407 (N_2407,In_594,In_2209);
and U2408 (N_2408,In_2729,In_979);
nand U2409 (N_2409,In_1474,In_491);
and U2410 (N_2410,In_2215,In_1857);
xnor U2411 (N_2411,In_1683,In_1505);
xnor U2412 (N_2412,In_1495,In_715);
nor U2413 (N_2413,In_2868,In_1285);
xnor U2414 (N_2414,In_658,In_1947);
xnor U2415 (N_2415,In_2429,In_2924);
nand U2416 (N_2416,In_2706,In_1320);
nor U2417 (N_2417,In_1546,In_922);
or U2418 (N_2418,In_460,In_2830);
nand U2419 (N_2419,In_468,In_2987);
or U2420 (N_2420,In_99,In_34);
and U2421 (N_2421,In_2652,In_2033);
nor U2422 (N_2422,In_2879,In_842);
or U2423 (N_2423,In_1285,In_1441);
nand U2424 (N_2424,In_2403,In_792);
or U2425 (N_2425,In_268,In_2873);
nor U2426 (N_2426,In_2594,In_320);
or U2427 (N_2427,In_608,In_621);
and U2428 (N_2428,In_103,In_1338);
xnor U2429 (N_2429,In_901,In_1430);
or U2430 (N_2430,In_514,In_614);
nand U2431 (N_2431,In_1722,In_2062);
nor U2432 (N_2432,In_97,In_960);
nand U2433 (N_2433,In_1243,In_326);
nor U2434 (N_2434,In_1639,In_1199);
nor U2435 (N_2435,In_626,In_25);
xor U2436 (N_2436,In_552,In_953);
xor U2437 (N_2437,In_1850,In_122);
or U2438 (N_2438,In_1831,In_2071);
nor U2439 (N_2439,In_72,In_950);
xor U2440 (N_2440,In_112,In_2174);
or U2441 (N_2441,In_1934,In_1287);
and U2442 (N_2442,In_1610,In_2310);
and U2443 (N_2443,In_1402,In_2092);
xnor U2444 (N_2444,In_2638,In_2789);
nor U2445 (N_2445,In_2718,In_1677);
nor U2446 (N_2446,In_2915,In_2316);
nor U2447 (N_2447,In_2145,In_1594);
nand U2448 (N_2448,In_390,In_1036);
nand U2449 (N_2449,In_76,In_364);
nand U2450 (N_2450,In_163,In_2025);
nor U2451 (N_2451,In_1849,In_648);
nand U2452 (N_2452,In_2850,In_343);
nor U2453 (N_2453,In_2057,In_382);
and U2454 (N_2454,In_2240,In_2679);
or U2455 (N_2455,In_792,In_232);
nor U2456 (N_2456,In_1601,In_2258);
or U2457 (N_2457,In_771,In_1964);
xnor U2458 (N_2458,In_54,In_117);
xnor U2459 (N_2459,In_2489,In_2049);
or U2460 (N_2460,In_315,In_2519);
nand U2461 (N_2461,In_1622,In_1673);
and U2462 (N_2462,In_2687,In_1061);
xor U2463 (N_2463,In_862,In_1943);
nand U2464 (N_2464,In_1724,In_2395);
xor U2465 (N_2465,In_200,In_55);
xnor U2466 (N_2466,In_388,In_766);
or U2467 (N_2467,In_341,In_2434);
and U2468 (N_2468,In_2847,In_408);
or U2469 (N_2469,In_1599,In_1831);
nor U2470 (N_2470,In_1577,In_1797);
nor U2471 (N_2471,In_2574,In_2162);
and U2472 (N_2472,In_1796,In_1987);
nor U2473 (N_2473,In_2359,In_2354);
xor U2474 (N_2474,In_425,In_2138);
nand U2475 (N_2475,In_913,In_1640);
xor U2476 (N_2476,In_2013,In_2651);
xnor U2477 (N_2477,In_381,In_990);
and U2478 (N_2478,In_1109,In_615);
nand U2479 (N_2479,In_2859,In_95);
xnor U2480 (N_2480,In_2908,In_1139);
or U2481 (N_2481,In_2201,In_636);
or U2482 (N_2482,In_2552,In_388);
nor U2483 (N_2483,In_376,In_604);
nor U2484 (N_2484,In_626,In_981);
nand U2485 (N_2485,In_2873,In_1898);
xor U2486 (N_2486,In_2522,In_2583);
and U2487 (N_2487,In_1890,In_2982);
and U2488 (N_2488,In_2157,In_2502);
and U2489 (N_2489,In_2104,In_1057);
nor U2490 (N_2490,In_862,In_841);
xor U2491 (N_2491,In_2706,In_2816);
or U2492 (N_2492,In_2510,In_1308);
nand U2493 (N_2493,In_1607,In_1182);
nand U2494 (N_2494,In_2257,In_2784);
nor U2495 (N_2495,In_255,In_454);
or U2496 (N_2496,In_1856,In_1048);
and U2497 (N_2497,In_2951,In_2946);
nor U2498 (N_2498,In_1111,In_1626);
xor U2499 (N_2499,In_1881,In_1125);
xor U2500 (N_2500,In_2323,In_163);
nand U2501 (N_2501,In_1431,In_117);
xor U2502 (N_2502,In_150,In_1555);
nand U2503 (N_2503,In_1909,In_2326);
or U2504 (N_2504,In_989,In_2694);
and U2505 (N_2505,In_201,In_1410);
xnor U2506 (N_2506,In_2690,In_1601);
and U2507 (N_2507,In_471,In_2350);
and U2508 (N_2508,In_1797,In_2423);
xnor U2509 (N_2509,In_1006,In_893);
xnor U2510 (N_2510,In_912,In_2658);
nand U2511 (N_2511,In_2443,In_543);
nor U2512 (N_2512,In_932,In_2600);
and U2513 (N_2513,In_131,In_4);
xor U2514 (N_2514,In_1800,In_1597);
nand U2515 (N_2515,In_2370,In_1024);
nand U2516 (N_2516,In_356,In_841);
xnor U2517 (N_2517,In_2755,In_2211);
and U2518 (N_2518,In_2118,In_1548);
nor U2519 (N_2519,In_2620,In_375);
xnor U2520 (N_2520,In_2576,In_1903);
xnor U2521 (N_2521,In_642,In_877);
and U2522 (N_2522,In_664,In_1779);
or U2523 (N_2523,In_1568,In_1451);
and U2524 (N_2524,In_1007,In_407);
or U2525 (N_2525,In_1307,In_697);
nor U2526 (N_2526,In_1061,In_2968);
xor U2527 (N_2527,In_871,In_386);
and U2528 (N_2528,In_2215,In_1900);
or U2529 (N_2529,In_658,In_948);
nand U2530 (N_2530,In_1806,In_27);
and U2531 (N_2531,In_2593,In_1327);
nor U2532 (N_2532,In_45,In_1712);
nor U2533 (N_2533,In_2929,In_2330);
xnor U2534 (N_2534,In_762,In_392);
nand U2535 (N_2535,In_1743,In_908);
xnor U2536 (N_2536,In_691,In_326);
nand U2537 (N_2537,In_2607,In_1746);
and U2538 (N_2538,In_179,In_2247);
or U2539 (N_2539,In_595,In_2380);
nor U2540 (N_2540,In_2982,In_2983);
nor U2541 (N_2541,In_95,In_2802);
and U2542 (N_2542,In_2177,In_1031);
or U2543 (N_2543,In_2984,In_2177);
nor U2544 (N_2544,In_2433,In_2597);
nor U2545 (N_2545,In_12,In_2216);
or U2546 (N_2546,In_735,In_791);
nor U2547 (N_2547,In_13,In_1412);
and U2548 (N_2548,In_2516,In_1681);
and U2549 (N_2549,In_1006,In_617);
or U2550 (N_2550,In_666,In_94);
and U2551 (N_2551,In_1757,In_2191);
nor U2552 (N_2552,In_1026,In_2388);
nand U2553 (N_2553,In_1778,In_2917);
and U2554 (N_2554,In_1424,In_123);
and U2555 (N_2555,In_2930,In_839);
or U2556 (N_2556,In_1619,In_2679);
and U2557 (N_2557,In_979,In_2151);
and U2558 (N_2558,In_2715,In_1875);
and U2559 (N_2559,In_1422,In_2087);
xor U2560 (N_2560,In_566,In_2022);
or U2561 (N_2561,In_1638,In_1730);
nand U2562 (N_2562,In_282,In_188);
nand U2563 (N_2563,In_2903,In_2311);
and U2564 (N_2564,In_2729,In_260);
and U2565 (N_2565,In_2198,In_2287);
or U2566 (N_2566,In_607,In_2292);
xnor U2567 (N_2567,In_313,In_1174);
xnor U2568 (N_2568,In_2043,In_2663);
nand U2569 (N_2569,In_785,In_1727);
and U2570 (N_2570,In_2207,In_334);
nand U2571 (N_2571,In_1421,In_1221);
and U2572 (N_2572,In_1984,In_2131);
xnor U2573 (N_2573,In_1466,In_278);
and U2574 (N_2574,In_2391,In_368);
and U2575 (N_2575,In_774,In_1211);
or U2576 (N_2576,In_1254,In_1866);
xor U2577 (N_2577,In_2265,In_2920);
or U2578 (N_2578,In_896,In_2324);
nor U2579 (N_2579,In_2062,In_69);
and U2580 (N_2580,In_2637,In_1282);
xor U2581 (N_2581,In_673,In_1526);
or U2582 (N_2582,In_2535,In_766);
nor U2583 (N_2583,In_1508,In_1455);
or U2584 (N_2584,In_2886,In_240);
and U2585 (N_2585,In_780,In_2382);
nand U2586 (N_2586,In_879,In_2301);
and U2587 (N_2587,In_2601,In_2229);
and U2588 (N_2588,In_2143,In_1933);
xnor U2589 (N_2589,In_527,In_186);
and U2590 (N_2590,In_2632,In_2945);
xnor U2591 (N_2591,In_258,In_1077);
and U2592 (N_2592,In_1258,In_133);
nand U2593 (N_2593,In_104,In_699);
nand U2594 (N_2594,In_2678,In_419);
xnor U2595 (N_2595,In_848,In_2223);
nand U2596 (N_2596,In_1312,In_2099);
and U2597 (N_2597,In_2233,In_128);
and U2598 (N_2598,In_168,In_613);
xnor U2599 (N_2599,In_170,In_2796);
xnor U2600 (N_2600,In_1649,In_2064);
xor U2601 (N_2601,In_1589,In_248);
nor U2602 (N_2602,In_77,In_1044);
xor U2603 (N_2603,In_542,In_2201);
and U2604 (N_2604,In_88,In_2975);
xor U2605 (N_2605,In_239,In_209);
xor U2606 (N_2606,In_2623,In_39);
xor U2607 (N_2607,In_384,In_206);
and U2608 (N_2608,In_937,In_2101);
nand U2609 (N_2609,In_1737,In_2070);
xor U2610 (N_2610,In_2825,In_941);
or U2611 (N_2611,In_2809,In_2472);
xnor U2612 (N_2612,In_917,In_2584);
nand U2613 (N_2613,In_1292,In_1607);
nand U2614 (N_2614,In_1042,In_715);
nor U2615 (N_2615,In_1752,In_45);
and U2616 (N_2616,In_78,In_382);
nand U2617 (N_2617,In_0,In_1511);
or U2618 (N_2618,In_1760,In_1816);
xor U2619 (N_2619,In_1792,In_441);
xnor U2620 (N_2620,In_32,In_1995);
and U2621 (N_2621,In_1262,In_115);
nand U2622 (N_2622,In_1527,In_1565);
or U2623 (N_2623,In_1313,In_2080);
and U2624 (N_2624,In_2801,In_2130);
nand U2625 (N_2625,In_2945,In_407);
xnor U2626 (N_2626,In_865,In_463);
and U2627 (N_2627,In_867,In_883);
nor U2628 (N_2628,In_1574,In_162);
or U2629 (N_2629,In_1896,In_1159);
or U2630 (N_2630,In_2524,In_2793);
and U2631 (N_2631,In_1289,In_732);
or U2632 (N_2632,In_2145,In_488);
or U2633 (N_2633,In_2980,In_1832);
or U2634 (N_2634,In_1752,In_1666);
nor U2635 (N_2635,In_834,In_1816);
or U2636 (N_2636,In_394,In_757);
or U2637 (N_2637,In_2655,In_1987);
nand U2638 (N_2638,In_1344,In_1433);
or U2639 (N_2639,In_544,In_451);
nand U2640 (N_2640,In_620,In_257);
and U2641 (N_2641,In_2207,In_1419);
xnor U2642 (N_2642,In_2290,In_2442);
nor U2643 (N_2643,In_1529,In_2319);
nor U2644 (N_2644,In_2491,In_2236);
nor U2645 (N_2645,In_1554,In_1222);
nand U2646 (N_2646,In_1811,In_576);
nor U2647 (N_2647,In_588,In_5);
nand U2648 (N_2648,In_464,In_1575);
xor U2649 (N_2649,In_1929,In_927);
xnor U2650 (N_2650,In_2887,In_1166);
xnor U2651 (N_2651,In_2088,In_2943);
nor U2652 (N_2652,In_274,In_424);
nand U2653 (N_2653,In_1547,In_2962);
nand U2654 (N_2654,In_1114,In_1910);
xor U2655 (N_2655,In_1281,In_1789);
or U2656 (N_2656,In_1969,In_2023);
or U2657 (N_2657,In_739,In_2782);
and U2658 (N_2658,In_1123,In_1710);
or U2659 (N_2659,In_121,In_2522);
xor U2660 (N_2660,In_2091,In_1999);
or U2661 (N_2661,In_2561,In_2717);
nor U2662 (N_2662,In_721,In_880);
xnor U2663 (N_2663,In_718,In_2688);
xnor U2664 (N_2664,In_1132,In_2016);
and U2665 (N_2665,In_642,In_1224);
nand U2666 (N_2666,In_2798,In_1668);
nand U2667 (N_2667,In_45,In_979);
xor U2668 (N_2668,In_163,In_2669);
nand U2669 (N_2669,In_2510,In_135);
or U2670 (N_2670,In_318,In_1621);
and U2671 (N_2671,In_1043,In_2974);
nand U2672 (N_2672,In_503,In_2136);
or U2673 (N_2673,In_2568,In_2585);
and U2674 (N_2674,In_286,In_1653);
and U2675 (N_2675,In_2371,In_1926);
nor U2676 (N_2676,In_1376,In_886);
xnor U2677 (N_2677,In_1553,In_1397);
or U2678 (N_2678,In_563,In_560);
nand U2679 (N_2679,In_1827,In_1998);
nor U2680 (N_2680,In_529,In_1942);
and U2681 (N_2681,In_563,In_1224);
nand U2682 (N_2682,In_1648,In_1471);
or U2683 (N_2683,In_1209,In_2759);
xnor U2684 (N_2684,In_1099,In_443);
and U2685 (N_2685,In_98,In_476);
and U2686 (N_2686,In_1273,In_1937);
nor U2687 (N_2687,In_2365,In_1795);
nor U2688 (N_2688,In_847,In_2700);
and U2689 (N_2689,In_106,In_368);
and U2690 (N_2690,In_1626,In_577);
nor U2691 (N_2691,In_2111,In_777);
and U2692 (N_2692,In_474,In_169);
or U2693 (N_2693,In_364,In_2500);
and U2694 (N_2694,In_2865,In_446);
or U2695 (N_2695,In_2606,In_2898);
nor U2696 (N_2696,In_808,In_1625);
xor U2697 (N_2697,In_2106,In_583);
xnor U2698 (N_2698,In_2148,In_2130);
xnor U2699 (N_2699,In_779,In_2541);
nor U2700 (N_2700,In_2439,In_697);
and U2701 (N_2701,In_908,In_92);
or U2702 (N_2702,In_1252,In_628);
xnor U2703 (N_2703,In_2983,In_54);
xor U2704 (N_2704,In_1286,In_1814);
nand U2705 (N_2705,In_669,In_621);
nand U2706 (N_2706,In_1016,In_1293);
nand U2707 (N_2707,In_2394,In_1201);
nand U2708 (N_2708,In_1085,In_1253);
nand U2709 (N_2709,In_2378,In_2174);
and U2710 (N_2710,In_207,In_492);
nor U2711 (N_2711,In_2059,In_1085);
xnor U2712 (N_2712,In_1261,In_2535);
xor U2713 (N_2713,In_1037,In_2921);
nor U2714 (N_2714,In_1620,In_817);
and U2715 (N_2715,In_225,In_1394);
xor U2716 (N_2716,In_625,In_1798);
nor U2717 (N_2717,In_1509,In_2669);
and U2718 (N_2718,In_2222,In_2575);
xnor U2719 (N_2719,In_2035,In_309);
nand U2720 (N_2720,In_1495,In_1592);
xnor U2721 (N_2721,In_2507,In_1252);
and U2722 (N_2722,In_2665,In_1024);
xor U2723 (N_2723,In_1912,In_1408);
and U2724 (N_2724,In_825,In_1455);
and U2725 (N_2725,In_641,In_420);
nand U2726 (N_2726,In_2896,In_1804);
and U2727 (N_2727,In_931,In_2960);
and U2728 (N_2728,In_1139,In_1529);
xnor U2729 (N_2729,In_1653,In_2323);
xor U2730 (N_2730,In_1231,In_487);
xnor U2731 (N_2731,In_1783,In_1412);
xor U2732 (N_2732,In_1457,In_251);
and U2733 (N_2733,In_1767,In_1723);
nor U2734 (N_2734,In_870,In_1797);
nand U2735 (N_2735,In_1827,In_985);
and U2736 (N_2736,In_1251,In_1852);
nand U2737 (N_2737,In_2273,In_1069);
xor U2738 (N_2738,In_2618,In_2812);
xnor U2739 (N_2739,In_2033,In_215);
xor U2740 (N_2740,In_1019,In_2407);
nor U2741 (N_2741,In_2843,In_2376);
xnor U2742 (N_2742,In_1626,In_2995);
nand U2743 (N_2743,In_2777,In_889);
nand U2744 (N_2744,In_781,In_839);
and U2745 (N_2745,In_2798,In_982);
nor U2746 (N_2746,In_1319,In_2677);
xnor U2747 (N_2747,In_606,In_30);
nor U2748 (N_2748,In_2344,In_854);
xor U2749 (N_2749,In_1907,In_2177);
nand U2750 (N_2750,In_1251,In_2433);
and U2751 (N_2751,In_1780,In_832);
and U2752 (N_2752,In_1195,In_2503);
xnor U2753 (N_2753,In_1300,In_2102);
xor U2754 (N_2754,In_2709,In_966);
or U2755 (N_2755,In_2543,In_2218);
nand U2756 (N_2756,In_1599,In_130);
nand U2757 (N_2757,In_2324,In_2914);
nor U2758 (N_2758,In_390,In_578);
nor U2759 (N_2759,In_2865,In_2479);
xor U2760 (N_2760,In_1224,In_2767);
xnor U2761 (N_2761,In_591,In_1740);
or U2762 (N_2762,In_614,In_1842);
nor U2763 (N_2763,In_2698,In_1906);
nor U2764 (N_2764,In_61,In_1264);
nand U2765 (N_2765,In_1395,In_2660);
or U2766 (N_2766,In_602,In_973);
and U2767 (N_2767,In_636,In_2279);
nand U2768 (N_2768,In_928,In_993);
and U2769 (N_2769,In_1474,In_2849);
and U2770 (N_2770,In_557,In_1388);
nand U2771 (N_2771,In_677,In_2807);
or U2772 (N_2772,In_2918,In_1827);
xnor U2773 (N_2773,In_250,In_1329);
nor U2774 (N_2774,In_601,In_430);
xnor U2775 (N_2775,In_2839,In_1841);
or U2776 (N_2776,In_2680,In_2611);
nand U2777 (N_2777,In_993,In_2379);
nor U2778 (N_2778,In_1315,In_1675);
and U2779 (N_2779,In_476,In_2174);
nand U2780 (N_2780,In_1588,In_761);
xor U2781 (N_2781,In_2550,In_1634);
xnor U2782 (N_2782,In_1129,In_98);
nor U2783 (N_2783,In_2031,In_605);
nand U2784 (N_2784,In_622,In_1952);
nand U2785 (N_2785,In_2016,In_1102);
or U2786 (N_2786,In_1838,In_1039);
nand U2787 (N_2787,In_28,In_500);
and U2788 (N_2788,In_915,In_1770);
xor U2789 (N_2789,In_2388,In_2305);
nand U2790 (N_2790,In_2418,In_1498);
xnor U2791 (N_2791,In_2531,In_1710);
nor U2792 (N_2792,In_462,In_799);
nor U2793 (N_2793,In_2040,In_1339);
and U2794 (N_2794,In_2485,In_2109);
and U2795 (N_2795,In_405,In_544);
nor U2796 (N_2796,In_524,In_816);
nand U2797 (N_2797,In_640,In_2045);
nor U2798 (N_2798,In_2934,In_1896);
or U2799 (N_2799,In_1297,In_2586);
nand U2800 (N_2800,In_193,In_1911);
and U2801 (N_2801,In_1159,In_1495);
xor U2802 (N_2802,In_2891,In_2290);
nor U2803 (N_2803,In_418,In_1643);
xnor U2804 (N_2804,In_882,In_1541);
nand U2805 (N_2805,In_2973,In_264);
or U2806 (N_2806,In_2393,In_2077);
nand U2807 (N_2807,In_421,In_457);
and U2808 (N_2808,In_2844,In_2543);
and U2809 (N_2809,In_1126,In_1199);
xor U2810 (N_2810,In_2403,In_1886);
or U2811 (N_2811,In_2696,In_559);
xor U2812 (N_2812,In_192,In_470);
nand U2813 (N_2813,In_534,In_471);
nand U2814 (N_2814,In_631,In_2403);
nand U2815 (N_2815,In_1776,In_1604);
or U2816 (N_2816,In_2927,In_1928);
or U2817 (N_2817,In_29,In_1313);
and U2818 (N_2818,In_1233,In_784);
nor U2819 (N_2819,In_2558,In_2927);
nand U2820 (N_2820,In_2125,In_525);
nor U2821 (N_2821,In_1660,In_1146);
xor U2822 (N_2822,In_1604,In_2431);
xnor U2823 (N_2823,In_722,In_962);
and U2824 (N_2824,In_896,In_369);
and U2825 (N_2825,In_2435,In_2866);
nand U2826 (N_2826,In_1417,In_2892);
nor U2827 (N_2827,In_2845,In_913);
nor U2828 (N_2828,In_2455,In_424);
or U2829 (N_2829,In_1638,In_2128);
xnor U2830 (N_2830,In_7,In_2965);
xor U2831 (N_2831,In_1242,In_1252);
xor U2832 (N_2832,In_1609,In_229);
nand U2833 (N_2833,In_200,In_1262);
nor U2834 (N_2834,In_2471,In_901);
nand U2835 (N_2835,In_2086,In_2317);
and U2836 (N_2836,In_483,In_279);
nor U2837 (N_2837,In_1603,In_655);
nor U2838 (N_2838,In_1970,In_729);
and U2839 (N_2839,In_2510,In_465);
nand U2840 (N_2840,In_1787,In_559);
and U2841 (N_2841,In_2739,In_2718);
and U2842 (N_2842,In_996,In_2649);
or U2843 (N_2843,In_2289,In_1523);
or U2844 (N_2844,In_167,In_2693);
nand U2845 (N_2845,In_291,In_2597);
or U2846 (N_2846,In_1080,In_1175);
nor U2847 (N_2847,In_2632,In_680);
nand U2848 (N_2848,In_2123,In_1027);
xnor U2849 (N_2849,In_446,In_2194);
and U2850 (N_2850,In_115,In_242);
or U2851 (N_2851,In_635,In_870);
xor U2852 (N_2852,In_1821,In_83);
nor U2853 (N_2853,In_2749,In_1437);
nor U2854 (N_2854,In_2114,In_241);
and U2855 (N_2855,In_2669,In_1624);
nand U2856 (N_2856,In_2988,In_512);
xnor U2857 (N_2857,In_74,In_1175);
xnor U2858 (N_2858,In_1960,In_366);
nand U2859 (N_2859,In_1856,In_920);
nor U2860 (N_2860,In_1602,In_830);
and U2861 (N_2861,In_2959,In_2775);
and U2862 (N_2862,In_495,In_1101);
nor U2863 (N_2863,In_2293,In_2595);
xnor U2864 (N_2864,In_1324,In_2576);
or U2865 (N_2865,In_2013,In_852);
and U2866 (N_2866,In_1765,In_2030);
xnor U2867 (N_2867,In_2453,In_1817);
and U2868 (N_2868,In_471,In_891);
and U2869 (N_2869,In_724,In_2268);
and U2870 (N_2870,In_2457,In_2183);
nand U2871 (N_2871,In_538,In_58);
or U2872 (N_2872,In_2535,In_571);
nor U2873 (N_2873,In_1233,In_253);
and U2874 (N_2874,In_2803,In_740);
nor U2875 (N_2875,In_1415,In_2702);
and U2876 (N_2876,In_1562,In_1902);
nand U2877 (N_2877,In_2810,In_332);
and U2878 (N_2878,In_1704,In_2839);
nor U2879 (N_2879,In_1659,In_2248);
nand U2880 (N_2880,In_2860,In_1111);
nand U2881 (N_2881,In_1378,In_1265);
nand U2882 (N_2882,In_1150,In_2574);
or U2883 (N_2883,In_2182,In_815);
or U2884 (N_2884,In_2182,In_1558);
or U2885 (N_2885,In_1764,In_2165);
nand U2886 (N_2886,In_1785,In_632);
xnor U2887 (N_2887,In_320,In_55);
xor U2888 (N_2888,In_136,In_1084);
or U2889 (N_2889,In_2796,In_48);
and U2890 (N_2890,In_2476,In_580);
nand U2891 (N_2891,In_1223,In_1328);
xor U2892 (N_2892,In_1544,In_1308);
and U2893 (N_2893,In_2367,In_21);
and U2894 (N_2894,In_2860,In_828);
xnor U2895 (N_2895,In_2325,In_797);
nor U2896 (N_2896,In_719,In_1756);
or U2897 (N_2897,In_412,In_15);
xor U2898 (N_2898,In_1951,In_846);
or U2899 (N_2899,In_2026,In_2565);
nand U2900 (N_2900,In_597,In_708);
and U2901 (N_2901,In_1226,In_1071);
xnor U2902 (N_2902,In_1397,In_420);
and U2903 (N_2903,In_627,In_2303);
nor U2904 (N_2904,In_2913,In_1580);
xor U2905 (N_2905,In_1425,In_1519);
and U2906 (N_2906,In_679,In_2372);
nand U2907 (N_2907,In_2718,In_2695);
nand U2908 (N_2908,In_2952,In_853);
or U2909 (N_2909,In_2165,In_2806);
or U2910 (N_2910,In_305,In_871);
xor U2911 (N_2911,In_2662,In_2621);
and U2912 (N_2912,In_1966,In_1206);
and U2913 (N_2913,In_828,In_99);
and U2914 (N_2914,In_1100,In_650);
or U2915 (N_2915,In_2495,In_890);
or U2916 (N_2916,In_2093,In_2223);
xor U2917 (N_2917,In_1401,In_2338);
xnor U2918 (N_2918,In_1364,In_554);
or U2919 (N_2919,In_1394,In_354);
nand U2920 (N_2920,In_2226,In_179);
xnor U2921 (N_2921,In_484,In_635);
and U2922 (N_2922,In_2575,In_1238);
nor U2923 (N_2923,In_1895,In_2660);
xnor U2924 (N_2924,In_2360,In_607);
nor U2925 (N_2925,In_1009,In_779);
or U2926 (N_2926,In_2638,In_770);
xnor U2927 (N_2927,In_1864,In_1825);
nor U2928 (N_2928,In_1175,In_2555);
or U2929 (N_2929,In_1186,In_231);
nor U2930 (N_2930,In_2996,In_1191);
or U2931 (N_2931,In_815,In_456);
xor U2932 (N_2932,In_2856,In_2471);
xor U2933 (N_2933,In_833,In_1802);
nor U2934 (N_2934,In_2183,In_2083);
nand U2935 (N_2935,In_1326,In_2657);
and U2936 (N_2936,In_1411,In_2826);
or U2937 (N_2937,In_1839,In_1126);
or U2938 (N_2938,In_2020,In_1640);
nand U2939 (N_2939,In_1555,In_2980);
and U2940 (N_2940,In_2861,In_2157);
nor U2941 (N_2941,In_588,In_361);
or U2942 (N_2942,In_2030,In_1771);
or U2943 (N_2943,In_702,In_1337);
nor U2944 (N_2944,In_945,In_826);
nor U2945 (N_2945,In_69,In_1510);
xnor U2946 (N_2946,In_1173,In_2324);
nor U2947 (N_2947,In_653,In_2787);
and U2948 (N_2948,In_242,In_1402);
or U2949 (N_2949,In_2511,In_2944);
nor U2950 (N_2950,In_383,In_1710);
nor U2951 (N_2951,In_271,In_2756);
or U2952 (N_2952,In_894,In_69);
xor U2953 (N_2953,In_1512,In_637);
nor U2954 (N_2954,In_241,In_2857);
and U2955 (N_2955,In_1938,In_369);
or U2956 (N_2956,In_2810,In_1684);
or U2957 (N_2957,In_1613,In_2815);
or U2958 (N_2958,In_2476,In_1473);
nand U2959 (N_2959,In_2076,In_1052);
nand U2960 (N_2960,In_1768,In_1613);
and U2961 (N_2961,In_1339,In_87);
xnor U2962 (N_2962,In_433,In_251);
nor U2963 (N_2963,In_1534,In_1033);
xor U2964 (N_2964,In_18,In_338);
or U2965 (N_2965,In_2371,In_785);
or U2966 (N_2966,In_2837,In_337);
or U2967 (N_2967,In_311,In_2013);
nor U2968 (N_2968,In_35,In_2210);
xnor U2969 (N_2969,In_1604,In_1174);
xnor U2970 (N_2970,In_159,In_2025);
xnor U2971 (N_2971,In_1659,In_1532);
nor U2972 (N_2972,In_1253,In_387);
and U2973 (N_2973,In_772,In_1519);
or U2974 (N_2974,In_2668,In_79);
xnor U2975 (N_2975,In_386,In_946);
nand U2976 (N_2976,In_2640,In_2686);
xnor U2977 (N_2977,In_1942,In_40);
or U2978 (N_2978,In_2278,In_2751);
nand U2979 (N_2979,In_2972,In_1997);
nand U2980 (N_2980,In_437,In_1906);
or U2981 (N_2981,In_66,In_990);
nand U2982 (N_2982,In_654,In_1933);
nor U2983 (N_2983,In_135,In_2709);
or U2984 (N_2984,In_2064,In_2010);
nor U2985 (N_2985,In_1860,In_2251);
xor U2986 (N_2986,In_1814,In_2074);
and U2987 (N_2987,In_1868,In_1317);
and U2988 (N_2988,In_2403,In_681);
nand U2989 (N_2989,In_402,In_2258);
xor U2990 (N_2990,In_1516,In_2053);
xor U2991 (N_2991,In_2204,In_690);
nor U2992 (N_2992,In_510,In_1090);
or U2993 (N_2993,In_2772,In_608);
nor U2994 (N_2994,In_702,In_2356);
nor U2995 (N_2995,In_671,In_2878);
nand U2996 (N_2996,In_1205,In_2316);
xor U2997 (N_2997,In_2519,In_2914);
nand U2998 (N_2998,In_111,In_2828);
nand U2999 (N_2999,In_504,In_916);
nand U3000 (N_3000,In_1609,In_1601);
and U3001 (N_3001,In_2369,In_1390);
and U3002 (N_3002,In_2228,In_1046);
and U3003 (N_3003,In_822,In_266);
xnor U3004 (N_3004,In_1718,In_2736);
nor U3005 (N_3005,In_783,In_453);
nor U3006 (N_3006,In_339,In_2482);
or U3007 (N_3007,In_1301,In_314);
and U3008 (N_3008,In_750,In_2080);
nand U3009 (N_3009,In_81,In_2990);
nand U3010 (N_3010,In_2661,In_649);
and U3011 (N_3011,In_117,In_2729);
nand U3012 (N_3012,In_2168,In_2120);
or U3013 (N_3013,In_1411,In_2395);
or U3014 (N_3014,In_2506,In_381);
nand U3015 (N_3015,In_2817,In_148);
nand U3016 (N_3016,In_1388,In_1644);
nand U3017 (N_3017,In_2131,In_1098);
xnor U3018 (N_3018,In_2619,In_2537);
nand U3019 (N_3019,In_1063,In_1987);
nand U3020 (N_3020,In_2037,In_1610);
nand U3021 (N_3021,In_603,In_1036);
and U3022 (N_3022,In_2036,In_32);
xnor U3023 (N_3023,In_2173,In_2246);
xnor U3024 (N_3024,In_2490,In_211);
nor U3025 (N_3025,In_1541,In_940);
xor U3026 (N_3026,In_418,In_375);
nand U3027 (N_3027,In_1964,In_653);
xnor U3028 (N_3028,In_897,In_2786);
nor U3029 (N_3029,In_2842,In_165);
or U3030 (N_3030,In_2598,In_560);
xnor U3031 (N_3031,In_1221,In_533);
nand U3032 (N_3032,In_219,In_1417);
nor U3033 (N_3033,In_273,In_1445);
xnor U3034 (N_3034,In_1940,In_1865);
nor U3035 (N_3035,In_1061,In_1955);
nor U3036 (N_3036,In_986,In_2307);
nand U3037 (N_3037,In_2833,In_1012);
nand U3038 (N_3038,In_86,In_2218);
xnor U3039 (N_3039,In_385,In_2642);
nor U3040 (N_3040,In_2908,In_2979);
xor U3041 (N_3041,In_1203,In_684);
xor U3042 (N_3042,In_507,In_1964);
nand U3043 (N_3043,In_82,In_2382);
xor U3044 (N_3044,In_1436,In_1613);
nand U3045 (N_3045,In_288,In_1585);
nor U3046 (N_3046,In_615,In_1814);
and U3047 (N_3047,In_2604,In_1885);
nand U3048 (N_3048,In_1744,In_1911);
nor U3049 (N_3049,In_2460,In_1088);
or U3050 (N_3050,In_235,In_421);
xor U3051 (N_3051,In_958,In_289);
or U3052 (N_3052,In_2852,In_971);
nand U3053 (N_3053,In_597,In_746);
xor U3054 (N_3054,In_842,In_214);
nor U3055 (N_3055,In_2727,In_2275);
nor U3056 (N_3056,In_221,In_2882);
and U3057 (N_3057,In_1382,In_755);
nor U3058 (N_3058,In_2757,In_2826);
xor U3059 (N_3059,In_2705,In_586);
nor U3060 (N_3060,In_1022,In_1897);
xor U3061 (N_3061,In_2453,In_2927);
and U3062 (N_3062,In_2134,In_344);
or U3063 (N_3063,In_1288,In_1124);
or U3064 (N_3064,In_1117,In_1556);
nand U3065 (N_3065,In_419,In_5);
nor U3066 (N_3066,In_2411,In_1765);
nand U3067 (N_3067,In_1600,In_1921);
or U3068 (N_3068,In_1991,In_1742);
and U3069 (N_3069,In_10,In_1812);
xor U3070 (N_3070,In_1091,In_2248);
nor U3071 (N_3071,In_2854,In_729);
and U3072 (N_3072,In_1924,In_602);
or U3073 (N_3073,In_1920,In_2763);
nand U3074 (N_3074,In_2637,In_2516);
or U3075 (N_3075,In_75,In_1956);
and U3076 (N_3076,In_659,In_449);
nand U3077 (N_3077,In_523,In_926);
nor U3078 (N_3078,In_2972,In_2954);
or U3079 (N_3079,In_2307,In_2021);
xor U3080 (N_3080,In_1104,In_2630);
and U3081 (N_3081,In_2596,In_873);
nand U3082 (N_3082,In_494,In_1704);
xor U3083 (N_3083,In_1277,In_2167);
nor U3084 (N_3084,In_1073,In_274);
nor U3085 (N_3085,In_2454,In_1489);
nand U3086 (N_3086,In_1483,In_1475);
nor U3087 (N_3087,In_1639,In_376);
xor U3088 (N_3088,In_372,In_1920);
or U3089 (N_3089,In_109,In_2918);
and U3090 (N_3090,In_1282,In_2478);
and U3091 (N_3091,In_1997,In_1165);
nand U3092 (N_3092,In_279,In_1213);
or U3093 (N_3093,In_1855,In_242);
xnor U3094 (N_3094,In_929,In_2564);
nor U3095 (N_3095,In_1804,In_2717);
and U3096 (N_3096,In_817,In_2271);
and U3097 (N_3097,In_2141,In_2999);
and U3098 (N_3098,In_1753,In_2264);
nor U3099 (N_3099,In_2720,In_2824);
and U3100 (N_3100,In_2113,In_2528);
nor U3101 (N_3101,In_161,In_2532);
or U3102 (N_3102,In_2372,In_2149);
and U3103 (N_3103,In_2591,In_889);
or U3104 (N_3104,In_1116,In_8);
or U3105 (N_3105,In_2896,In_2672);
nor U3106 (N_3106,In_2999,In_2081);
nand U3107 (N_3107,In_1655,In_2781);
or U3108 (N_3108,In_1467,In_221);
nor U3109 (N_3109,In_1440,In_2012);
or U3110 (N_3110,In_2699,In_707);
xnor U3111 (N_3111,In_2124,In_411);
and U3112 (N_3112,In_1363,In_743);
and U3113 (N_3113,In_2508,In_784);
nand U3114 (N_3114,In_2079,In_297);
nand U3115 (N_3115,In_1940,In_964);
or U3116 (N_3116,In_2335,In_1859);
xnor U3117 (N_3117,In_1707,In_2248);
xor U3118 (N_3118,In_151,In_689);
xnor U3119 (N_3119,In_2166,In_1079);
and U3120 (N_3120,In_1899,In_2785);
and U3121 (N_3121,In_2089,In_2435);
and U3122 (N_3122,In_1347,In_1946);
or U3123 (N_3123,In_2946,In_708);
xnor U3124 (N_3124,In_1461,In_1112);
nor U3125 (N_3125,In_1980,In_2570);
xnor U3126 (N_3126,In_870,In_2990);
nor U3127 (N_3127,In_2357,In_1983);
nand U3128 (N_3128,In_215,In_1647);
or U3129 (N_3129,In_483,In_2932);
xor U3130 (N_3130,In_2863,In_2436);
and U3131 (N_3131,In_2111,In_2292);
or U3132 (N_3132,In_2182,In_1205);
nor U3133 (N_3133,In_928,In_807);
nor U3134 (N_3134,In_798,In_1714);
nor U3135 (N_3135,In_2990,In_138);
xnor U3136 (N_3136,In_1324,In_2837);
xnor U3137 (N_3137,In_1853,In_2840);
xnor U3138 (N_3138,In_557,In_2821);
nand U3139 (N_3139,In_1890,In_903);
or U3140 (N_3140,In_351,In_2935);
or U3141 (N_3141,In_1803,In_368);
nand U3142 (N_3142,In_2967,In_396);
nor U3143 (N_3143,In_2362,In_1493);
nor U3144 (N_3144,In_2457,In_698);
and U3145 (N_3145,In_640,In_140);
nand U3146 (N_3146,In_857,In_1201);
and U3147 (N_3147,In_2775,In_668);
nor U3148 (N_3148,In_134,In_2685);
or U3149 (N_3149,In_774,In_1386);
nand U3150 (N_3150,In_318,In_2325);
xor U3151 (N_3151,In_2529,In_1185);
nor U3152 (N_3152,In_87,In_2757);
xor U3153 (N_3153,In_1977,In_1497);
xor U3154 (N_3154,In_122,In_334);
or U3155 (N_3155,In_2516,In_1742);
or U3156 (N_3156,In_1537,In_2913);
nor U3157 (N_3157,In_1815,In_1216);
or U3158 (N_3158,In_842,In_377);
nor U3159 (N_3159,In_1138,In_2847);
nand U3160 (N_3160,In_676,In_2625);
or U3161 (N_3161,In_2967,In_2983);
and U3162 (N_3162,In_2134,In_34);
nor U3163 (N_3163,In_2786,In_1728);
xnor U3164 (N_3164,In_2887,In_2181);
nand U3165 (N_3165,In_2485,In_2133);
nor U3166 (N_3166,In_1614,In_2189);
xnor U3167 (N_3167,In_1118,In_2582);
xor U3168 (N_3168,In_2522,In_1365);
or U3169 (N_3169,In_1441,In_2090);
and U3170 (N_3170,In_2265,In_1255);
nand U3171 (N_3171,In_579,In_2513);
xnor U3172 (N_3172,In_1655,In_60);
nor U3173 (N_3173,In_1383,In_311);
nor U3174 (N_3174,In_2009,In_2819);
nor U3175 (N_3175,In_2248,In_2498);
nand U3176 (N_3176,In_132,In_1141);
nand U3177 (N_3177,In_1490,In_1368);
and U3178 (N_3178,In_554,In_1851);
and U3179 (N_3179,In_2326,In_742);
and U3180 (N_3180,In_2815,In_144);
xnor U3181 (N_3181,In_1898,In_2351);
nand U3182 (N_3182,In_1629,In_48);
xnor U3183 (N_3183,In_1099,In_2023);
xor U3184 (N_3184,In_2830,In_455);
nand U3185 (N_3185,In_797,In_628);
and U3186 (N_3186,In_2692,In_110);
or U3187 (N_3187,In_322,In_1406);
xnor U3188 (N_3188,In_430,In_953);
or U3189 (N_3189,In_2912,In_459);
xor U3190 (N_3190,In_60,In_629);
and U3191 (N_3191,In_1477,In_2092);
nor U3192 (N_3192,In_480,In_2555);
or U3193 (N_3193,In_1026,In_1097);
nand U3194 (N_3194,In_568,In_1766);
or U3195 (N_3195,In_2280,In_2216);
nand U3196 (N_3196,In_2377,In_2620);
nand U3197 (N_3197,In_1933,In_1830);
nand U3198 (N_3198,In_1851,In_2584);
nand U3199 (N_3199,In_2142,In_2913);
and U3200 (N_3200,In_2372,In_583);
nand U3201 (N_3201,In_478,In_94);
nand U3202 (N_3202,In_2584,In_388);
nor U3203 (N_3203,In_32,In_641);
or U3204 (N_3204,In_199,In_661);
and U3205 (N_3205,In_2901,In_1504);
and U3206 (N_3206,In_522,In_1176);
nand U3207 (N_3207,In_2768,In_619);
nand U3208 (N_3208,In_1314,In_2708);
xnor U3209 (N_3209,In_2353,In_233);
and U3210 (N_3210,In_2964,In_1168);
and U3211 (N_3211,In_2166,In_2468);
nor U3212 (N_3212,In_38,In_684);
or U3213 (N_3213,In_2493,In_732);
and U3214 (N_3214,In_86,In_23);
and U3215 (N_3215,In_375,In_206);
and U3216 (N_3216,In_2000,In_1632);
or U3217 (N_3217,In_2334,In_854);
and U3218 (N_3218,In_742,In_231);
nand U3219 (N_3219,In_1174,In_1371);
nand U3220 (N_3220,In_2049,In_1993);
xor U3221 (N_3221,In_1019,In_2360);
nor U3222 (N_3222,In_899,In_760);
nor U3223 (N_3223,In_2399,In_667);
or U3224 (N_3224,In_509,In_2716);
or U3225 (N_3225,In_705,In_1608);
nand U3226 (N_3226,In_993,In_2878);
nor U3227 (N_3227,In_2165,In_2854);
nand U3228 (N_3228,In_2093,In_1056);
and U3229 (N_3229,In_1458,In_783);
nand U3230 (N_3230,In_472,In_1575);
nand U3231 (N_3231,In_467,In_379);
or U3232 (N_3232,In_962,In_2815);
or U3233 (N_3233,In_1862,In_813);
or U3234 (N_3234,In_1755,In_2499);
nand U3235 (N_3235,In_2425,In_1242);
and U3236 (N_3236,In_1002,In_2648);
and U3237 (N_3237,In_782,In_1759);
or U3238 (N_3238,In_2062,In_2954);
xor U3239 (N_3239,In_1035,In_1848);
nor U3240 (N_3240,In_837,In_1532);
and U3241 (N_3241,In_2328,In_2053);
nand U3242 (N_3242,In_1578,In_1001);
xor U3243 (N_3243,In_1794,In_2708);
nor U3244 (N_3244,In_1613,In_598);
nor U3245 (N_3245,In_2194,In_11);
or U3246 (N_3246,In_1693,In_1630);
xnor U3247 (N_3247,In_2602,In_1927);
nor U3248 (N_3248,In_2260,In_2039);
xnor U3249 (N_3249,In_347,In_2019);
nor U3250 (N_3250,In_2110,In_805);
xor U3251 (N_3251,In_2099,In_2047);
nand U3252 (N_3252,In_2926,In_2894);
xnor U3253 (N_3253,In_1013,In_1622);
or U3254 (N_3254,In_885,In_507);
and U3255 (N_3255,In_1123,In_759);
nor U3256 (N_3256,In_2613,In_1356);
nand U3257 (N_3257,In_58,In_702);
nor U3258 (N_3258,In_2511,In_1033);
nor U3259 (N_3259,In_1981,In_411);
xnor U3260 (N_3260,In_1447,In_411);
and U3261 (N_3261,In_2121,In_1411);
nand U3262 (N_3262,In_2143,In_463);
and U3263 (N_3263,In_2267,In_170);
nand U3264 (N_3264,In_1867,In_2411);
or U3265 (N_3265,In_654,In_1281);
nor U3266 (N_3266,In_1468,In_2931);
nor U3267 (N_3267,In_1558,In_2801);
nor U3268 (N_3268,In_1960,In_81);
or U3269 (N_3269,In_1954,In_1008);
or U3270 (N_3270,In_99,In_1572);
and U3271 (N_3271,In_842,In_1606);
and U3272 (N_3272,In_2238,In_102);
and U3273 (N_3273,In_268,In_367);
nand U3274 (N_3274,In_1622,In_1818);
and U3275 (N_3275,In_2536,In_497);
nand U3276 (N_3276,In_822,In_2487);
or U3277 (N_3277,In_2447,In_1463);
nand U3278 (N_3278,In_2033,In_189);
nor U3279 (N_3279,In_673,In_1201);
xor U3280 (N_3280,In_2947,In_538);
nand U3281 (N_3281,In_2292,In_1099);
nor U3282 (N_3282,In_1022,In_868);
and U3283 (N_3283,In_910,In_491);
and U3284 (N_3284,In_2304,In_1649);
or U3285 (N_3285,In_801,In_1671);
or U3286 (N_3286,In_1619,In_863);
and U3287 (N_3287,In_980,In_2381);
xnor U3288 (N_3288,In_2944,In_2820);
xor U3289 (N_3289,In_2402,In_1624);
nor U3290 (N_3290,In_1806,In_459);
nor U3291 (N_3291,In_2614,In_710);
or U3292 (N_3292,In_2154,In_1712);
nor U3293 (N_3293,In_1893,In_2200);
and U3294 (N_3294,In_1971,In_2826);
nand U3295 (N_3295,In_789,In_521);
and U3296 (N_3296,In_1528,In_98);
nor U3297 (N_3297,In_655,In_1892);
or U3298 (N_3298,In_1202,In_199);
nor U3299 (N_3299,In_201,In_2668);
xor U3300 (N_3300,In_232,In_2950);
and U3301 (N_3301,In_675,In_186);
xnor U3302 (N_3302,In_1209,In_1882);
xor U3303 (N_3303,In_44,In_1345);
xor U3304 (N_3304,In_1342,In_362);
nor U3305 (N_3305,In_928,In_2053);
or U3306 (N_3306,In_2633,In_1225);
nor U3307 (N_3307,In_1547,In_1381);
nor U3308 (N_3308,In_1508,In_1019);
nor U3309 (N_3309,In_2099,In_2635);
nand U3310 (N_3310,In_924,In_986);
nand U3311 (N_3311,In_1710,In_406);
or U3312 (N_3312,In_777,In_1229);
or U3313 (N_3313,In_163,In_2984);
xnor U3314 (N_3314,In_913,In_2067);
and U3315 (N_3315,In_2593,In_1868);
nand U3316 (N_3316,In_988,In_387);
xor U3317 (N_3317,In_2191,In_670);
xor U3318 (N_3318,In_978,In_2409);
or U3319 (N_3319,In_695,In_1708);
and U3320 (N_3320,In_1801,In_2339);
xor U3321 (N_3321,In_1155,In_466);
nand U3322 (N_3322,In_1272,In_832);
nand U3323 (N_3323,In_1614,In_11);
and U3324 (N_3324,In_2617,In_1146);
and U3325 (N_3325,In_1874,In_2483);
nor U3326 (N_3326,In_1747,In_43);
nand U3327 (N_3327,In_2268,In_518);
xor U3328 (N_3328,In_1826,In_836);
nand U3329 (N_3329,In_613,In_925);
and U3330 (N_3330,In_2515,In_95);
xor U3331 (N_3331,In_1098,In_1962);
and U3332 (N_3332,In_1868,In_884);
xnor U3333 (N_3333,In_1669,In_830);
nor U3334 (N_3334,In_2631,In_1383);
nand U3335 (N_3335,In_297,In_308);
xnor U3336 (N_3336,In_2919,In_1076);
or U3337 (N_3337,In_2229,In_584);
nand U3338 (N_3338,In_1879,In_1754);
and U3339 (N_3339,In_975,In_1659);
nand U3340 (N_3340,In_2643,In_1744);
nor U3341 (N_3341,In_1260,In_1510);
nand U3342 (N_3342,In_2178,In_1980);
nand U3343 (N_3343,In_664,In_2733);
and U3344 (N_3344,In_256,In_998);
nand U3345 (N_3345,In_2547,In_490);
nand U3346 (N_3346,In_992,In_1841);
nor U3347 (N_3347,In_692,In_116);
xor U3348 (N_3348,In_1817,In_507);
and U3349 (N_3349,In_2959,In_1361);
xnor U3350 (N_3350,In_2712,In_2116);
nand U3351 (N_3351,In_1173,In_656);
or U3352 (N_3352,In_687,In_777);
nand U3353 (N_3353,In_2844,In_369);
or U3354 (N_3354,In_911,In_1046);
and U3355 (N_3355,In_2833,In_980);
nor U3356 (N_3356,In_2137,In_1610);
nor U3357 (N_3357,In_2406,In_2649);
or U3358 (N_3358,In_2284,In_825);
or U3359 (N_3359,In_2102,In_35);
and U3360 (N_3360,In_1903,In_1442);
or U3361 (N_3361,In_1526,In_442);
or U3362 (N_3362,In_850,In_582);
nand U3363 (N_3363,In_809,In_2137);
and U3364 (N_3364,In_1770,In_421);
xnor U3365 (N_3365,In_2350,In_611);
nor U3366 (N_3366,In_196,In_293);
nand U3367 (N_3367,In_1650,In_1687);
nand U3368 (N_3368,In_1085,In_502);
and U3369 (N_3369,In_458,In_1369);
or U3370 (N_3370,In_2090,In_1797);
or U3371 (N_3371,In_2633,In_688);
xnor U3372 (N_3372,In_1744,In_860);
nor U3373 (N_3373,In_2615,In_1358);
nor U3374 (N_3374,In_105,In_607);
xor U3375 (N_3375,In_2484,In_1399);
and U3376 (N_3376,In_2484,In_101);
or U3377 (N_3377,In_2754,In_2943);
nor U3378 (N_3378,In_534,In_1270);
and U3379 (N_3379,In_988,In_2390);
and U3380 (N_3380,In_1696,In_2156);
and U3381 (N_3381,In_2491,In_1091);
or U3382 (N_3382,In_2432,In_1911);
or U3383 (N_3383,In_91,In_672);
xor U3384 (N_3384,In_59,In_887);
and U3385 (N_3385,In_82,In_2779);
xor U3386 (N_3386,In_2563,In_1068);
or U3387 (N_3387,In_1770,In_2424);
and U3388 (N_3388,In_720,In_2950);
or U3389 (N_3389,In_1424,In_193);
nand U3390 (N_3390,In_997,In_1660);
or U3391 (N_3391,In_1473,In_737);
xnor U3392 (N_3392,In_2538,In_741);
or U3393 (N_3393,In_2288,In_1204);
and U3394 (N_3394,In_870,In_954);
or U3395 (N_3395,In_815,In_2870);
or U3396 (N_3396,In_1600,In_2929);
nand U3397 (N_3397,In_1934,In_1756);
nand U3398 (N_3398,In_2209,In_2422);
or U3399 (N_3399,In_2572,In_820);
nor U3400 (N_3400,In_202,In_2254);
xnor U3401 (N_3401,In_2365,In_2116);
nor U3402 (N_3402,In_126,In_1935);
nand U3403 (N_3403,In_1969,In_1333);
or U3404 (N_3404,In_1780,In_1410);
or U3405 (N_3405,In_1309,In_1950);
xnor U3406 (N_3406,In_721,In_2413);
xnor U3407 (N_3407,In_2096,In_1649);
and U3408 (N_3408,In_2184,In_734);
and U3409 (N_3409,In_1755,In_2137);
or U3410 (N_3410,In_1257,In_403);
nand U3411 (N_3411,In_2922,In_2696);
nor U3412 (N_3412,In_49,In_2789);
and U3413 (N_3413,In_1195,In_1818);
nor U3414 (N_3414,In_1842,In_2176);
and U3415 (N_3415,In_2257,In_1507);
and U3416 (N_3416,In_1013,In_2902);
or U3417 (N_3417,In_1505,In_216);
nand U3418 (N_3418,In_2778,In_2160);
nand U3419 (N_3419,In_1149,In_2094);
and U3420 (N_3420,In_2315,In_1116);
and U3421 (N_3421,In_359,In_2106);
nor U3422 (N_3422,In_999,In_741);
nor U3423 (N_3423,In_697,In_2680);
nor U3424 (N_3424,In_405,In_1117);
xor U3425 (N_3425,In_1372,In_2639);
or U3426 (N_3426,In_2870,In_2989);
nand U3427 (N_3427,In_548,In_1249);
xnor U3428 (N_3428,In_2952,In_1458);
xor U3429 (N_3429,In_1085,In_2927);
and U3430 (N_3430,In_655,In_2727);
and U3431 (N_3431,In_1447,In_1769);
and U3432 (N_3432,In_2983,In_2280);
nand U3433 (N_3433,In_127,In_131);
and U3434 (N_3434,In_1173,In_200);
xor U3435 (N_3435,In_1020,In_1385);
nand U3436 (N_3436,In_330,In_2099);
nand U3437 (N_3437,In_1969,In_1872);
or U3438 (N_3438,In_1969,In_1768);
nor U3439 (N_3439,In_1940,In_2287);
xor U3440 (N_3440,In_216,In_1767);
xnor U3441 (N_3441,In_2207,In_1505);
nand U3442 (N_3442,In_197,In_623);
xor U3443 (N_3443,In_576,In_692);
nor U3444 (N_3444,In_2186,In_1586);
or U3445 (N_3445,In_938,In_1738);
nor U3446 (N_3446,In_195,In_2906);
and U3447 (N_3447,In_1926,In_1193);
or U3448 (N_3448,In_1058,In_497);
and U3449 (N_3449,In_2909,In_22);
or U3450 (N_3450,In_2931,In_2170);
and U3451 (N_3451,In_1196,In_2141);
nor U3452 (N_3452,In_2487,In_513);
and U3453 (N_3453,In_2013,In_1861);
xor U3454 (N_3454,In_2295,In_1024);
or U3455 (N_3455,In_2837,In_1183);
nor U3456 (N_3456,In_97,In_1949);
nand U3457 (N_3457,In_574,In_182);
nand U3458 (N_3458,In_1623,In_487);
and U3459 (N_3459,In_2012,In_33);
or U3460 (N_3460,In_438,In_2839);
or U3461 (N_3461,In_228,In_689);
and U3462 (N_3462,In_2735,In_1050);
or U3463 (N_3463,In_80,In_1939);
and U3464 (N_3464,In_2784,In_2673);
xnor U3465 (N_3465,In_2048,In_1200);
nand U3466 (N_3466,In_575,In_1863);
nand U3467 (N_3467,In_742,In_794);
nor U3468 (N_3468,In_1557,In_631);
nor U3469 (N_3469,In_338,In_179);
or U3470 (N_3470,In_375,In_1851);
nand U3471 (N_3471,In_1138,In_2058);
xor U3472 (N_3472,In_2867,In_1104);
nand U3473 (N_3473,In_810,In_1474);
xnor U3474 (N_3474,In_1496,In_2418);
xnor U3475 (N_3475,In_1442,In_643);
xnor U3476 (N_3476,In_2497,In_1988);
xor U3477 (N_3477,In_1259,In_2500);
nor U3478 (N_3478,In_2251,In_449);
nor U3479 (N_3479,In_2181,In_1418);
xor U3480 (N_3480,In_659,In_1866);
xnor U3481 (N_3481,In_903,In_1145);
or U3482 (N_3482,In_858,In_2242);
xor U3483 (N_3483,In_2634,In_1672);
nor U3484 (N_3484,In_341,In_2846);
nor U3485 (N_3485,In_1729,In_33);
and U3486 (N_3486,In_575,In_2986);
or U3487 (N_3487,In_556,In_2177);
nand U3488 (N_3488,In_100,In_787);
nand U3489 (N_3489,In_589,In_1604);
and U3490 (N_3490,In_2760,In_2461);
or U3491 (N_3491,In_1911,In_1202);
or U3492 (N_3492,In_1036,In_2330);
nor U3493 (N_3493,In_2415,In_2475);
or U3494 (N_3494,In_203,In_1939);
and U3495 (N_3495,In_106,In_879);
or U3496 (N_3496,In_815,In_2539);
nor U3497 (N_3497,In_1881,In_810);
xnor U3498 (N_3498,In_1900,In_1323);
or U3499 (N_3499,In_1248,In_2591);
and U3500 (N_3500,In_2908,In_1559);
or U3501 (N_3501,In_702,In_2934);
nand U3502 (N_3502,In_218,In_891);
and U3503 (N_3503,In_2138,In_1156);
nor U3504 (N_3504,In_2664,In_2414);
xor U3505 (N_3505,In_1326,In_699);
xnor U3506 (N_3506,In_1149,In_1984);
xor U3507 (N_3507,In_2819,In_682);
nor U3508 (N_3508,In_2574,In_675);
nand U3509 (N_3509,In_32,In_1111);
xor U3510 (N_3510,In_1099,In_86);
or U3511 (N_3511,In_1680,In_2528);
nand U3512 (N_3512,In_1999,In_1510);
nand U3513 (N_3513,In_2316,In_1479);
xnor U3514 (N_3514,In_1505,In_1675);
xor U3515 (N_3515,In_1298,In_2953);
nand U3516 (N_3516,In_382,In_1565);
nand U3517 (N_3517,In_1350,In_2894);
xnor U3518 (N_3518,In_1895,In_291);
nor U3519 (N_3519,In_141,In_1383);
and U3520 (N_3520,In_1820,In_2379);
xor U3521 (N_3521,In_2118,In_963);
or U3522 (N_3522,In_2622,In_1192);
or U3523 (N_3523,In_1857,In_845);
or U3524 (N_3524,In_2726,In_459);
or U3525 (N_3525,In_851,In_1608);
and U3526 (N_3526,In_2529,In_1995);
nand U3527 (N_3527,In_2982,In_2686);
and U3528 (N_3528,In_420,In_2547);
nor U3529 (N_3529,In_740,In_392);
nand U3530 (N_3530,In_2075,In_2409);
and U3531 (N_3531,In_646,In_1666);
nand U3532 (N_3532,In_146,In_2969);
and U3533 (N_3533,In_1148,In_197);
xnor U3534 (N_3534,In_1769,In_809);
nor U3535 (N_3535,In_2047,In_969);
xor U3536 (N_3536,In_2625,In_2709);
or U3537 (N_3537,In_1654,In_120);
nor U3538 (N_3538,In_818,In_886);
nor U3539 (N_3539,In_900,In_2969);
nand U3540 (N_3540,In_1541,In_2248);
and U3541 (N_3541,In_1017,In_360);
nor U3542 (N_3542,In_700,In_475);
nor U3543 (N_3543,In_1474,In_72);
xnor U3544 (N_3544,In_565,In_2119);
or U3545 (N_3545,In_1273,In_848);
nor U3546 (N_3546,In_740,In_2690);
nor U3547 (N_3547,In_1879,In_1755);
xnor U3548 (N_3548,In_805,In_1943);
nor U3549 (N_3549,In_456,In_2761);
or U3550 (N_3550,In_2789,In_1906);
nand U3551 (N_3551,In_2664,In_2291);
xnor U3552 (N_3552,In_2690,In_2639);
nor U3553 (N_3553,In_1879,In_2622);
or U3554 (N_3554,In_2580,In_183);
xor U3555 (N_3555,In_2903,In_1238);
xnor U3556 (N_3556,In_2021,In_471);
and U3557 (N_3557,In_2493,In_2129);
nand U3558 (N_3558,In_873,In_1186);
nand U3559 (N_3559,In_1745,In_685);
nand U3560 (N_3560,In_962,In_455);
or U3561 (N_3561,In_735,In_1502);
or U3562 (N_3562,In_494,In_868);
xor U3563 (N_3563,In_751,In_616);
xnor U3564 (N_3564,In_1749,In_2695);
nand U3565 (N_3565,In_187,In_1616);
nor U3566 (N_3566,In_625,In_2032);
or U3567 (N_3567,In_2301,In_1149);
or U3568 (N_3568,In_2290,In_1946);
or U3569 (N_3569,In_169,In_408);
nor U3570 (N_3570,In_1173,In_1665);
nor U3571 (N_3571,In_236,In_2655);
or U3572 (N_3572,In_4,In_719);
nor U3573 (N_3573,In_1446,In_2168);
and U3574 (N_3574,In_790,In_1574);
nor U3575 (N_3575,In_2967,In_526);
and U3576 (N_3576,In_832,In_174);
or U3577 (N_3577,In_1129,In_41);
nor U3578 (N_3578,In_1918,In_2772);
xnor U3579 (N_3579,In_2809,In_735);
nand U3580 (N_3580,In_2084,In_600);
xor U3581 (N_3581,In_2928,In_226);
and U3582 (N_3582,In_2980,In_473);
or U3583 (N_3583,In_1482,In_56);
or U3584 (N_3584,In_2207,In_1871);
or U3585 (N_3585,In_364,In_1298);
and U3586 (N_3586,In_123,In_2118);
xnor U3587 (N_3587,In_300,In_2254);
or U3588 (N_3588,In_2804,In_2510);
nand U3589 (N_3589,In_1633,In_1996);
or U3590 (N_3590,In_599,In_1640);
or U3591 (N_3591,In_962,In_415);
or U3592 (N_3592,In_1659,In_2523);
xor U3593 (N_3593,In_1495,In_316);
xor U3594 (N_3594,In_627,In_1996);
nand U3595 (N_3595,In_1623,In_258);
and U3596 (N_3596,In_1511,In_326);
nand U3597 (N_3597,In_1857,In_2321);
nand U3598 (N_3598,In_291,In_2880);
and U3599 (N_3599,In_1915,In_2897);
or U3600 (N_3600,In_888,In_1470);
and U3601 (N_3601,In_2204,In_779);
nor U3602 (N_3602,In_146,In_2167);
xor U3603 (N_3603,In_868,In_2764);
nand U3604 (N_3604,In_1298,In_514);
and U3605 (N_3605,In_1165,In_1592);
nand U3606 (N_3606,In_765,In_141);
nand U3607 (N_3607,In_102,In_770);
and U3608 (N_3608,In_2641,In_88);
xor U3609 (N_3609,In_594,In_790);
nand U3610 (N_3610,In_1897,In_775);
nand U3611 (N_3611,In_2421,In_31);
nor U3612 (N_3612,In_1809,In_2625);
nand U3613 (N_3613,In_804,In_2108);
and U3614 (N_3614,In_411,In_2625);
and U3615 (N_3615,In_234,In_758);
xnor U3616 (N_3616,In_1785,In_2694);
or U3617 (N_3617,In_750,In_1331);
or U3618 (N_3618,In_639,In_1486);
nor U3619 (N_3619,In_902,In_2593);
nor U3620 (N_3620,In_1916,In_1198);
xnor U3621 (N_3621,In_43,In_2154);
or U3622 (N_3622,In_2412,In_1702);
nor U3623 (N_3623,In_2045,In_549);
nand U3624 (N_3624,In_2375,In_1366);
xor U3625 (N_3625,In_225,In_2850);
nor U3626 (N_3626,In_2629,In_2067);
nor U3627 (N_3627,In_2042,In_2500);
nand U3628 (N_3628,In_703,In_2347);
nor U3629 (N_3629,In_1272,In_1597);
xor U3630 (N_3630,In_1953,In_1092);
and U3631 (N_3631,In_223,In_2448);
or U3632 (N_3632,In_1222,In_1506);
xor U3633 (N_3633,In_1317,In_2829);
or U3634 (N_3634,In_2448,In_460);
or U3635 (N_3635,In_42,In_2918);
nand U3636 (N_3636,In_2787,In_1921);
or U3637 (N_3637,In_1704,In_2972);
nor U3638 (N_3638,In_1347,In_2069);
xor U3639 (N_3639,In_1385,In_726);
and U3640 (N_3640,In_576,In_1863);
nor U3641 (N_3641,In_2309,In_1600);
xor U3642 (N_3642,In_2849,In_2138);
or U3643 (N_3643,In_1283,In_697);
or U3644 (N_3644,In_2057,In_2002);
nand U3645 (N_3645,In_2677,In_1148);
or U3646 (N_3646,In_2050,In_537);
xor U3647 (N_3647,In_258,In_2052);
nor U3648 (N_3648,In_2724,In_367);
and U3649 (N_3649,In_1048,In_1941);
or U3650 (N_3650,In_2000,In_226);
or U3651 (N_3651,In_328,In_2280);
and U3652 (N_3652,In_658,In_302);
nand U3653 (N_3653,In_1572,In_2830);
and U3654 (N_3654,In_2794,In_968);
nand U3655 (N_3655,In_2095,In_286);
and U3656 (N_3656,In_1552,In_1932);
nand U3657 (N_3657,In_812,In_1281);
or U3658 (N_3658,In_1404,In_2205);
and U3659 (N_3659,In_855,In_259);
and U3660 (N_3660,In_414,In_1726);
nand U3661 (N_3661,In_2508,In_965);
nand U3662 (N_3662,In_2942,In_2840);
and U3663 (N_3663,In_2397,In_2285);
nand U3664 (N_3664,In_317,In_1460);
and U3665 (N_3665,In_1357,In_2794);
nand U3666 (N_3666,In_951,In_641);
xor U3667 (N_3667,In_2741,In_633);
nand U3668 (N_3668,In_2173,In_2262);
nor U3669 (N_3669,In_1912,In_1995);
or U3670 (N_3670,In_1958,In_1240);
xnor U3671 (N_3671,In_986,In_1929);
and U3672 (N_3672,In_240,In_912);
xor U3673 (N_3673,In_408,In_1551);
and U3674 (N_3674,In_133,In_633);
and U3675 (N_3675,In_1219,In_469);
nand U3676 (N_3676,In_2450,In_1001);
nor U3677 (N_3677,In_2333,In_887);
or U3678 (N_3678,In_153,In_1992);
xnor U3679 (N_3679,In_2180,In_1618);
xor U3680 (N_3680,In_2691,In_366);
nand U3681 (N_3681,In_885,In_2630);
xnor U3682 (N_3682,In_1232,In_2108);
xor U3683 (N_3683,In_2501,In_247);
nor U3684 (N_3684,In_242,In_2575);
and U3685 (N_3685,In_1283,In_853);
and U3686 (N_3686,In_218,In_1694);
xnor U3687 (N_3687,In_2374,In_2337);
and U3688 (N_3688,In_2546,In_2798);
nand U3689 (N_3689,In_2229,In_1533);
or U3690 (N_3690,In_1028,In_920);
or U3691 (N_3691,In_1944,In_2699);
or U3692 (N_3692,In_1689,In_1434);
nor U3693 (N_3693,In_428,In_2122);
or U3694 (N_3694,In_1224,In_1900);
nor U3695 (N_3695,In_1426,In_2576);
nand U3696 (N_3696,In_2673,In_717);
and U3697 (N_3697,In_593,In_2349);
nor U3698 (N_3698,In_115,In_1306);
and U3699 (N_3699,In_2833,In_557);
nand U3700 (N_3700,In_1865,In_1339);
xor U3701 (N_3701,In_53,In_344);
xnor U3702 (N_3702,In_1746,In_2138);
nor U3703 (N_3703,In_1674,In_2755);
or U3704 (N_3704,In_2516,In_2336);
xnor U3705 (N_3705,In_2267,In_2671);
nor U3706 (N_3706,In_1610,In_2308);
nor U3707 (N_3707,In_2874,In_1505);
nor U3708 (N_3708,In_2864,In_1086);
xor U3709 (N_3709,In_2132,In_666);
and U3710 (N_3710,In_2766,In_2676);
xor U3711 (N_3711,In_1907,In_865);
or U3712 (N_3712,In_272,In_40);
or U3713 (N_3713,In_721,In_1858);
and U3714 (N_3714,In_37,In_184);
nand U3715 (N_3715,In_2015,In_1724);
or U3716 (N_3716,In_2252,In_1996);
and U3717 (N_3717,In_2207,In_133);
xnor U3718 (N_3718,In_914,In_2164);
or U3719 (N_3719,In_804,In_1864);
or U3720 (N_3720,In_88,In_2008);
xnor U3721 (N_3721,In_503,In_111);
nor U3722 (N_3722,In_507,In_20);
xnor U3723 (N_3723,In_2795,In_1025);
nor U3724 (N_3724,In_2873,In_220);
or U3725 (N_3725,In_2775,In_2543);
and U3726 (N_3726,In_2745,In_784);
or U3727 (N_3727,In_2405,In_906);
nor U3728 (N_3728,In_2854,In_1489);
nor U3729 (N_3729,In_2905,In_487);
and U3730 (N_3730,In_468,In_837);
or U3731 (N_3731,In_214,In_1771);
xor U3732 (N_3732,In_285,In_2396);
and U3733 (N_3733,In_399,In_579);
and U3734 (N_3734,In_886,In_2148);
xor U3735 (N_3735,In_1294,In_1604);
xnor U3736 (N_3736,In_1225,In_258);
xor U3737 (N_3737,In_2720,In_2450);
nor U3738 (N_3738,In_1724,In_1646);
nor U3739 (N_3739,In_1123,In_1232);
nor U3740 (N_3740,In_764,In_140);
and U3741 (N_3741,In_2568,In_1054);
nand U3742 (N_3742,In_360,In_414);
nand U3743 (N_3743,In_1121,In_1344);
and U3744 (N_3744,In_2783,In_2718);
and U3745 (N_3745,In_2156,In_313);
nand U3746 (N_3746,In_2769,In_602);
nand U3747 (N_3747,In_934,In_1234);
nand U3748 (N_3748,In_1211,In_193);
nand U3749 (N_3749,In_124,In_1475);
xor U3750 (N_3750,In_52,In_542);
and U3751 (N_3751,In_886,In_2626);
or U3752 (N_3752,In_2495,In_2022);
or U3753 (N_3753,In_1778,In_790);
or U3754 (N_3754,In_2902,In_333);
and U3755 (N_3755,In_1190,In_840);
nand U3756 (N_3756,In_146,In_2667);
xnor U3757 (N_3757,In_1945,In_470);
nand U3758 (N_3758,In_1077,In_2427);
nand U3759 (N_3759,In_1079,In_2014);
or U3760 (N_3760,In_1778,In_1752);
nand U3761 (N_3761,In_2116,In_2966);
and U3762 (N_3762,In_678,In_2364);
or U3763 (N_3763,In_1842,In_2854);
or U3764 (N_3764,In_2800,In_2373);
xor U3765 (N_3765,In_2177,In_2290);
xnor U3766 (N_3766,In_115,In_2535);
xor U3767 (N_3767,In_737,In_385);
xor U3768 (N_3768,In_720,In_1638);
xor U3769 (N_3769,In_1342,In_1037);
and U3770 (N_3770,In_2090,In_1498);
nand U3771 (N_3771,In_1190,In_1345);
nor U3772 (N_3772,In_2467,In_80);
and U3773 (N_3773,In_1368,In_365);
and U3774 (N_3774,In_95,In_1214);
nor U3775 (N_3775,In_2520,In_499);
xor U3776 (N_3776,In_1680,In_300);
xor U3777 (N_3777,In_1308,In_267);
xor U3778 (N_3778,In_249,In_739);
xnor U3779 (N_3779,In_1829,In_421);
nor U3780 (N_3780,In_2614,In_1636);
or U3781 (N_3781,In_1178,In_165);
nor U3782 (N_3782,In_1902,In_556);
nand U3783 (N_3783,In_1863,In_1344);
nor U3784 (N_3784,In_2947,In_669);
xnor U3785 (N_3785,In_1534,In_2955);
or U3786 (N_3786,In_2303,In_2515);
nand U3787 (N_3787,In_648,In_1771);
nand U3788 (N_3788,In_1674,In_2752);
and U3789 (N_3789,In_1727,In_1403);
nand U3790 (N_3790,In_314,In_308);
nand U3791 (N_3791,In_2514,In_1622);
and U3792 (N_3792,In_807,In_1153);
or U3793 (N_3793,In_2425,In_746);
xor U3794 (N_3794,In_2973,In_520);
and U3795 (N_3795,In_355,In_2788);
nor U3796 (N_3796,In_2726,In_664);
nor U3797 (N_3797,In_1047,In_2454);
nand U3798 (N_3798,In_168,In_1634);
nor U3799 (N_3799,In_2970,In_2388);
xor U3800 (N_3800,In_2215,In_2683);
nand U3801 (N_3801,In_2438,In_2985);
and U3802 (N_3802,In_979,In_1169);
xor U3803 (N_3803,In_2611,In_354);
or U3804 (N_3804,In_838,In_693);
nand U3805 (N_3805,In_2375,In_292);
nor U3806 (N_3806,In_2316,In_1204);
nand U3807 (N_3807,In_650,In_2260);
nor U3808 (N_3808,In_1951,In_2719);
or U3809 (N_3809,In_1576,In_506);
and U3810 (N_3810,In_1008,In_1842);
xor U3811 (N_3811,In_2617,In_568);
and U3812 (N_3812,In_2509,In_2407);
and U3813 (N_3813,In_1890,In_1696);
xor U3814 (N_3814,In_1850,In_224);
and U3815 (N_3815,In_1266,In_1033);
xor U3816 (N_3816,In_2833,In_2233);
xnor U3817 (N_3817,In_759,In_2832);
or U3818 (N_3818,In_1965,In_1592);
nand U3819 (N_3819,In_678,In_176);
xor U3820 (N_3820,In_361,In_2111);
xnor U3821 (N_3821,In_190,In_213);
and U3822 (N_3822,In_2845,In_1215);
xnor U3823 (N_3823,In_580,In_1280);
xnor U3824 (N_3824,In_1506,In_2662);
nand U3825 (N_3825,In_121,In_2877);
xnor U3826 (N_3826,In_2618,In_1063);
xor U3827 (N_3827,In_1472,In_1085);
or U3828 (N_3828,In_1482,In_2651);
nand U3829 (N_3829,In_176,In_1964);
or U3830 (N_3830,In_595,In_2416);
nor U3831 (N_3831,In_2613,In_2017);
or U3832 (N_3832,In_1906,In_217);
xnor U3833 (N_3833,In_2517,In_2706);
and U3834 (N_3834,In_1239,In_2382);
and U3835 (N_3835,In_2689,In_2518);
or U3836 (N_3836,In_2637,In_154);
nor U3837 (N_3837,In_1080,In_2093);
xor U3838 (N_3838,In_2482,In_2714);
or U3839 (N_3839,In_2125,In_1681);
xnor U3840 (N_3840,In_1103,In_1649);
and U3841 (N_3841,In_2493,In_2650);
xor U3842 (N_3842,In_45,In_1137);
or U3843 (N_3843,In_1064,In_2239);
xor U3844 (N_3844,In_1736,In_107);
nor U3845 (N_3845,In_2069,In_373);
nand U3846 (N_3846,In_520,In_840);
xnor U3847 (N_3847,In_2233,In_237);
xnor U3848 (N_3848,In_1372,In_1601);
xor U3849 (N_3849,In_1301,In_273);
and U3850 (N_3850,In_1242,In_1798);
xnor U3851 (N_3851,In_5,In_2790);
nand U3852 (N_3852,In_2006,In_2973);
nor U3853 (N_3853,In_1731,In_212);
xnor U3854 (N_3854,In_816,In_2961);
nor U3855 (N_3855,In_1902,In_697);
nand U3856 (N_3856,In_24,In_32);
and U3857 (N_3857,In_1705,In_657);
nor U3858 (N_3858,In_1313,In_831);
and U3859 (N_3859,In_2606,In_2125);
xor U3860 (N_3860,In_1155,In_1827);
or U3861 (N_3861,In_2599,In_1964);
and U3862 (N_3862,In_229,In_2893);
nor U3863 (N_3863,In_130,In_1096);
nor U3864 (N_3864,In_2136,In_2760);
xnor U3865 (N_3865,In_1453,In_1828);
nand U3866 (N_3866,In_1837,In_1465);
xor U3867 (N_3867,In_615,In_687);
or U3868 (N_3868,In_1078,In_2418);
xnor U3869 (N_3869,In_1610,In_2320);
xnor U3870 (N_3870,In_767,In_521);
nand U3871 (N_3871,In_1702,In_1079);
nor U3872 (N_3872,In_2315,In_2318);
or U3873 (N_3873,In_941,In_1141);
nor U3874 (N_3874,In_2266,In_508);
xor U3875 (N_3875,In_2283,In_2141);
and U3876 (N_3876,In_2300,In_1176);
or U3877 (N_3877,In_2576,In_2727);
nand U3878 (N_3878,In_1377,In_2420);
xor U3879 (N_3879,In_1693,In_1405);
and U3880 (N_3880,In_1260,In_2874);
nand U3881 (N_3881,In_2282,In_1764);
and U3882 (N_3882,In_2079,In_1967);
xnor U3883 (N_3883,In_596,In_1);
xor U3884 (N_3884,In_1643,In_2942);
nand U3885 (N_3885,In_1220,In_1203);
and U3886 (N_3886,In_907,In_2074);
and U3887 (N_3887,In_1099,In_2248);
nand U3888 (N_3888,In_377,In_75);
and U3889 (N_3889,In_1126,In_2936);
xnor U3890 (N_3890,In_2656,In_1379);
xnor U3891 (N_3891,In_2767,In_645);
xnor U3892 (N_3892,In_1911,In_2553);
and U3893 (N_3893,In_1765,In_193);
nor U3894 (N_3894,In_2601,In_165);
nor U3895 (N_3895,In_2157,In_828);
or U3896 (N_3896,In_2432,In_113);
nand U3897 (N_3897,In_834,In_1785);
nand U3898 (N_3898,In_275,In_2934);
or U3899 (N_3899,In_2229,In_146);
and U3900 (N_3900,In_2494,In_2170);
and U3901 (N_3901,In_1098,In_1531);
nor U3902 (N_3902,In_1131,In_1243);
xnor U3903 (N_3903,In_2604,In_976);
or U3904 (N_3904,In_1050,In_84);
xnor U3905 (N_3905,In_1160,In_2500);
nor U3906 (N_3906,In_407,In_2584);
or U3907 (N_3907,In_328,In_2601);
xor U3908 (N_3908,In_863,In_1153);
or U3909 (N_3909,In_24,In_2746);
xor U3910 (N_3910,In_2739,In_2542);
nand U3911 (N_3911,In_1803,In_2123);
xor U3912 (N_3912,In_80,In_2812);
nor U3913 (N_3913,In_2888,In_1806);
nor U3914 (N_3914,In_679,In_716);
or U3915 (N_3915,In_404,In_1684);
xnor U3916 (N_3916,In_1317,In_1286);
xnor U3917 (N_3917,In_633,In_2796);
or U3918 (N_3918,In_946,In_1909);
nor U3919 (N_3919,In_200,In_2944);
and U3920 (N_3920,In_2774,In_1224);
xor U3921 (N_3921,In_740,In_1025);
nand U3922 (N_3922,In_2274,In_104);
or U3923 (N_3923,In_1104,In_1599);
nor U3924 (N_3924,In_495,In_2171);
nand U3925 (N_3925,In_1240,In_2606);
nor U3926 (N_3926,In_2591,In_363);
nand U3927 (N_3927,In_851,In_1687);
xor U3928 (N_3928,In_1202,In_541);
nand U3929 (N_3929,In_603,In_428);
or U3930 (N_3930,In_1362,In_2987);
xnor U3931 (N_3931,In_1308,In_2757);
xor U3932 (N_3932,In_1497,In_166);
nor U3933 (N_3933,In_1855,In_1301);
xor U3934 (N_3934,In_997,In_2436);
and U3935 (N_3935,In_1920,In_2824);
xnor U3936 (N_3936,In_97,In_2517);
nand U3937 (N_3937,In_2870,In_1464);
xor U3938 (N_3938,In_419,In_50);
or U3939 (N_3939,In_432,In_883);
or U3940 (N_3940,In_1960,In_655);
or U3941 (N_3941,In_179,In_2530);
and U3942 (N_3942,In_832,In_2949);
xnor U3943 (N_3943,In_261,In_818);
xor U3944 (N_3944,In_54,In_347);
nand U3945 (N_3945,In_1196,In_1515);
or U3946 (N_3946,In_1274,In_2111);
nand U3947 (N_3947,In_1164,In_378);
nor U3948 (N_3948,In_2938,In_412);
xor U3949 (N_3949,In_728,In_40);
and U3950 (N_3950,In_556,In_199);
and U3951 (N_3951,In_1226,In_231);
nor U3952 (N_3952,In_710,In_2348);
nand U3953 (N_3953,In_2504,In_1988);
xor U3954 (N_3954,In_104,In_2320);
nand U3955 (N_3955,In_62,In_2677);
or U3956 (N_3956,In_194,In_1363);
xor U3957 (N_3957,In_2214,In_975);
nor U3958 (N_3958,In_2105,In_1247);
and U3959 (N_3959,In_1092,In_81);
or U3960 (N_3960,In_2064,In_2569);
xnor U3961 (N_3961,In_1240,In_2313);
nor U3962 (N_3962,In_42,In_1774);
nor U3963 (N_3963,In_2465,In_2977);
nand U3964 (N_3964,In_678,In_822);
and U3965 (N_3965,In_1510,In_1066);
and U3966 (N_3966,In_532,In_2694);
nor U3967 (N_3967,In_2992,In_1679);
or U3968 (N_3968,In_2735,In_2827);
or U3969 (N_3969,In_1253,In_2105);
or U3970 (N_3970,In_2357,In_2232);
nand U3971 (N_3971,In_2656,In_909);
nand U3972 (N_3972,In_1491,In_2314);
nor U3973 (N_3973,In_2776,In_1262);
xor U3974 (N_3974,In_1804,In_903);
and U3975 (N_3975,In_52,In_2476);
and U3976 (N_3976,In_1148,In_1530);
xor U3977 (N_3977,In_52,In_112);
and U3978 (N_3978,In_2425,In_1595);
nand U3979 (N_3979,In_787,In_1951);
and U3980 (N_3980,In_1179,In_816);
and U3981 (N_3981,In_2992,In_666);
nor U3982 (N_3982,In_1067,In_2246);
or U3983 (N_3983,In_148,In_1251);
nand U3984 (N_3984,In_974,In_2473);
nand U3985 (N_3985,In_2465,In_2130);
nor U3986 (N_3986,In_2320,In_2193);
or U3987 (N_3987,In_1941,In_1434);
nand U3988 (N_3988,In_2975,In_1930);
nor U3989 (N_3989,In_1186,In_655);
or U3990 (N_3990,In_428,In_293);
nand U3991 (N_3991,In_1484,In_588);
nor U3992 (N_3992,In_2416,In_987);
and U3993 (N_3993,In_1472,In_2487);
nand U3994 (N_3994,In_2266,In_2405);
nor U3995 (N_3995,In_1383,In_1457);
nand U3996 (N_3996,In_1796,In_2060);
nand U3997 (N_3997,In_277,In_1649);
or U3998 (N_3998,In_247,In_984);
and U3999 (N_3999,In_2555,In_2157);
nand U4000 (N_4000,In_996,In_859);
xor U4001 (N_4001,In_509,In_1441);
xnor U4002 (N_4002,In_1478,In_2254);
nand U4003 (N_4003,In_1328,In_161);
or U4004 (N_4004,In_1028,In_1319);
or U4005 (N_4005,In_2036,In_2266);
and U4006 (N_4006,In_576,In_1673);
or U4007 (N_4007,In_2502,In_695);
nand U4008 (N_4008,In_1412,In_172);
nor U4009 (N_4009,In_1241,In_2627);
or U4010 (N_4010,In_1398,In_2655);
nand U4011 (N_4011,In_1878,In_2987);
nand U4012 (N_4012,In_2634,In_2591);
or U4013 (N_4013,In_1601,In_1864);
or U4014 (N_4014,In_1712,In_2105);
or U4015 (N_4015,In_1009,In_2843);
nor U4016 (N_4016,In_730,In_2405);
nor U4017 (N_4017,In_432,In_1927);
xor U4018 (N_4018,In_180,In_1912);
nor U4019 (N_4019,In_1852,In_2045);
and U4020 (N_4020,In_2606,In_723);
or U4021 (N_4021,In_2451,In_401);
nor U4022 (N_4022,In_2259,In_2215);
nand U4023 (N_4023,In_454,In_287);
xnor U4024 (N_4024,In_2223,In_2180);
nand U4025 (N_4025,In_2170,In_2721);
nor U4026 (N_4026,In_2986,In_328);
nor U4027 (N_4027,In_324,In_1465);
nand U4028 (N_4028,In_151,In_2231);
or U4029 (N_4029,In_2877,In_930);
nor U4030 (N_4030,In_2065,In_1700);
xnor U4031 (N_4031,In_2902,In_819);
and U4032 (N_4032,In_715,In_2461);
nor U4033 (N_4033,In_1437,In_376);
and U4034 (N_4034,In_2384,In_1975);
nor U4035 (N_4035,In_1631,In_2086);
and U4036 (N_4036,In_1170,In_2658);
xnor U4037 (N_4037,In_1933,In_1866);
nor U4038 (N_4038,In_2100,In_2182);
and U4039 (N_4039,In_2692,In_2483);
and U4040 (N_4040,In_1865,In_1101);
nand U4041 (N_4041,In_2488,In_1312);
and U4042 (N_4042,In_836,In_248);
or U4043 (N_4043,In_2498,In_2430);
or U4044 (N_4044,In_1808,In_2174);
and U4045 (N_4045,In_422,In_2990);
or U4046 (N_4046,In_2302,In_2609);
and U4047 (N_4047,In_1749,In_702);
and U4048 (N_4048,In_2876,In_553);
and U4049 (N_4049,In_1978,In_2205);
or U4050 (N_4050,In_1598,In_2020);
nor U4051 (N_4051,In_1305,In_1845);
nor U4052 (N_4052,In_1805,In_1635);
or U4053 (N_4053,In_708,In_2608);
nand U4054 (N_4054,In_2648,In_436);
xnor U4055 (N_4055,In_1938,In_18);
xor U4056 (N_4056,In_2241,In_1499);
and U4057 (N_4057,In_2285,In_756);
nand U4058 (N_4058,In_96,In_1342);
nand U4059 (N_4059,In_1779,In_1418);
xnor U4060 (N_4060,In_1130,In_1720);
nor U4061 (N_4061,In_2458,In_1948);
xnor U4062 (N_4062,In_1741,In_1007);
xnor U4063 (N_4063,In_2192,In_1091);
or U4064 (N_4064,In_323,In_1933);
nor U4065 (N_4065,In_374,In_2252);
nor U4066 (N_4066,In_1860,In_884);
and U4067 (N_4067,In_2584,In_1830);
and U4068 (N_4068,In_2913,In_2277);
xnor U4069 (N_4069,In_1786,In_1695);
nor U4070 (N_4070,In_42,In_1275);
nor U4071 (N_4071,In_976,In_518);
and U4072 (N_4072,In_1618,In_211);
or U4073 (N_4073,In_504,In_2896);
xor U4074 (N_4074,In_2784,In_233);
xnor U4075 (N_4075,In_703,In_1068);
xnor U4076 (N_4076,In_603,In_2594);
or U4077 (N_4077,In_1999,In_2868);
xor U4078 (N_4078,In_1256,In_459);
or U4079 (N_4079,In_518,In_1163);
xor U4080 (N_4080,In_746,In_1454);
nand U4081 (N_4081,In_1558,In_2658);
nor U4082 (N_4082,In_2915,In_404);
nand U4083 (N_4083,In_437,In_1765);
nor U4084 (N_4084,In_182,In_2646);
xnor U4085 (N_4085,In_2761,In_1944);
nand U4086 (N_4086,In_2707,In_121);
nor U4087 (N_4087,In_1915,In_1307);
xor U4088 (N_4088,In_2274,In_440);
or U4089 (N_4089,In_356,In_1168);
nand U4090 (N_4090,In_2954,In_208);
nand U4091 (N_4091,In_2795,In_1191);
nor U4092 (N_4092,In_1286,In_1706);
nand U4093 (N_4093,In_1885,In_344);
nor U4094 (N_4094,In_1163,In_231);
and U4095 (N_4095,In_2111,In_9);
xor U4096 (N_4096,In_94,In_780);
or U4097 (N_4097,In_2583,In_293);
or U4098 (N_4098,In_1698,In_2852);
or U4099 (N_4099,In_1982,In_2870);
and U4100 (N_4100,In_1476,In_485);
and U4101 (N_4101,In_2001,In_1129);
xor U4102 (N_4102,In_2770,In_1780);
or U4103 (N_4103,In_1862,In_1142);
nand U4104 (N_4104,In_394,In_1488);
nand U4105 (N_4105,In_17,In_110);
nor U4106 (N_4106,In_869,In_750);
xnor U4107 (N_4107,In_851,In_2332);
nor U4108 (N_4108,In_659,In_443);
and U4109 (N_4109,In_2984,In_989);
xnor U4110 (N_4110,In_1604,In_2205);
or U4111 (N_4111,In_80,In_448);
nand U4112 (N_4112,In_2371,In_1804);
or U4113 (N_4113,In_1646,In_1403);
nor U4114 (N_4114,In_1366,In_80);
or U4115 (N_4115,In_2018,In_1023);
nand U4116 (N_4116,In_1749,In_1680);
nor U4117 (N_4117,In_510,In_622);
nand U4118 (N_4118,In_2125,In_2978);
and U4119 (N_4119,In_602,In_2747);
nand U4120 (N_4120,In_2729,In_697);
and U4121 (N_4121,In_1149,In_49);
nand U4122 (N_4122,In_989,In_1112);
nor U4123 (N_4123,In_1914,In_2858);
xnor U4124 (N_4124,In_541,In_2230);
and U4125 (N_4125,In_203,In_1367);
nor U4126 (N_4126,In_946,In_1245);
and U4127 (N_4127,In_779,In_72);
and U4128 (N_4128,In_193,In_680);
xor U4129 (N_4129,In_902,In_839);
nor U4130 (N_4130,In_1744,In_1456);
and U4131 (N_4131,In_773,In_622);
nor U4132 (N_4132,In_1814,In_1824);
and U4133 (N_4133,In_631,In_1454);
nand U4134 (N_4134,In_89,In_8);
xnor U4135 (N_4135,In_2466,In_1767);
nand U4136 (N_4136,In_2872,In_1405);
nor U4137 (N_4137,In_1891,In_1156);
nand U4138 (N_4138,In_957,In_1970);
xor U4139 (N_4139,In_350,In_1261);
nor U4140 (N_4140,In_583,In_472);
and U4141 (N_4141,In_719,In_2368);
and U4142 (N_4142,In_940,In_873);
nor U4143 (N_4143,In_246,In_1244);
nor U4144 (N_4144,In_84,In_1107);
xnor U4145 (N_4145,In_2515,In_57);
and U4146 (N_4146,In_2756,In_853);
nand U4147 (N_4147,In_2756,In_865);
or U4148 (N_4148,In_1391,In_2388);
nor U4149 (N_4149,In_448,In_2573);
nor U4150 (N_4150,In_155,In_1136);
or U4151 (N_4151,In_2318,In_1821);
nor U4152 (N_4152,In_1855,In_2307);
or U4153 (N_4153,In_2798,In_2828);
nor U4154 (N_4154,In_2491,In_1609);
nor U4155 (N_4155,In_490,In_402);
xor U4156 (N_4156,In_1008,In_2680);
nand U4157 (N_4157,In_2829,In_652);
nand U4158 (N_4158,In_651,In_927);
and U4159 (N_4159,In_297,In_994);
and U4160 (N_4160,In_2295,In_1655);
or U4161 (N_4161,In_2848,In_2356);
and U4162 (N_4162,In_253,In_2391);
and U4163 (N_4163,In_949,In_2024);
xor U4164 (N_4164,In_688,In_812);
and U4165 (N_4165,In_1576,In_1187);
or U4166 (N_4166,In_1434,In_2506);
nor U4167 (N_4167,In_548,In_811);
and U4168 (N_4168,In_1853,In_2405);
xor U4169 (N_4169,In_1439,In_98);
nand U4170 (N_4170,In_1402,In_1711);
xor U4171 (N_4171,In_1047,In_379);
xnor U4172 (N_4172,In_753,In_2769);
and U4173 (N_4173,In_2257,In_2909);
nor U4174 (N_4174,In_2144,In_2885);
nand U4175 (N_4175,In_1568,In_585);
nor U4176 (N_4176,In_2019,In_1636);
nand U4177 (N_4177,In_1124,In_923);
nand U4178 (N_4178,In_250,In_302);
or U4179 (N_4179,In_252,In_56);
or U4180 (N_4180,In_1168,In_399);
or U4181 (N_4181,In_2458,In_1136);
nor U4182 (N_4182,In_141,In_1655);
nand U4183 (N_4183,In_581,In_1158);
nand U4184 (N_4184,In_437,In_2675);
nor U4185 (N_4185,In_110,In_634);
nand U4186 (N_4186,In_2235,In_359);
or U4187 (N_4187,In_2299,In_2480);
nor U4188 (N_4188,In_1970,In_2008);
nand U4189 (N_4189,In_2469,In_1852);
xor U4190 (N_4190,In_1712,In_2780);
or U4191 (N_4191,In_1855,In_1318);
nor U4192 (N_4192,In_1259,In_1366);
or U4193 (N_4193,In_1858,In_582);
and U4194 (N_4194,In_919,In_1526);
or U4195 (N_4195,In_1527,In_1744);
nand U4196 (N_4196,In_2826,In_726);
and U4197 (N_4197,In_2398,In_2701);
and U4198 (N_4198,In_2804,In_1097);
or U4199 (N_4199,In_2560,In_148);
or U4200 (N_4200,In_775,In_2094);
and U4201 (N_4201,In_1527,In_131);
nor U4202 (N_4202,In_1585,In_417);
and U4203 (N_4203,In_2454,In_1286);
and U4204 (N_4204,In_2518,In_1300);
or U4205 (N_4205,In_2782,In_903);
or U4206 (N_4206,In_52,In_2207);
xnor U4207 (N_4207,In_553,In_2035);
and U4208 (N_4208,In_2706,In_2445);
xor U4209 (N_4209,In_1094,In_2114);
xor U4210 (N_4210,In_2631,In_1671);
or U4211 (N_4211,In_286,In_1038);
or U4212 (N_4212,In_1696,In_2432);
nor U4213 (N_4213,In_603,In_2043);
or U4214 (N_4214,In_16,In_620);
or U4215 (N_4215,In_70,In_906);
or U4216 (N_4216,In_2043,In_648);
or U4217 (N_4217,In_340,In_1016);
xor U4218 (N_4218,In_522,In_960);
nand U4219 (N_4219,In_973,In_38);
and U4220 (N_4220,In_5,In_1630);
nor U4221 (N_4221,In_188,In_92);
or U4222 (N_4222,In_2764,In_2990);
or U4223 (N_4223,In_365,In_981);
nor U4224 (N_4224,In_1517,In_2599);
and U4225 (N_4225,In_2885,In_1459);
nand U4226 (N_4226,In_235,In_36);
and U4227 (N_4227,In_2402,In_2019);
or U4228 (N_4228,In_1527,In_1309);
xor U4229 (N_4229,In_2638,In_2956);
and U4230 (N_4230,In_1656,In_1833);
xnor U4231 (N_4231,In_1927,In_134);
nand U4232 (N_4232,In_2260,In_1380);
and U4233 (N_4233,In_2106,In_1282);
nor U4234 (N_4234,In_1895,In_1104);
and U4235 (N_4235,In_2140,In_1974);
and U4236 (N_4236,In_48,In_1897);
nor U4237 (N_4237,In_2339,In_1883);
xnor U4238 (N_4238,In_2311,In_30);
nor U4239 (N_4239,In_33,In_2888);
and U4240 (N_4240,In_262,In_119);
or U4241 (N_4241,In_2121,In_343);
xnor U4242 (N_4242,In_1149,In_2320);
xor U4243 (N_4243,In_612,In_2711);
nor U4244 (N_4244,In_2879,In_1161);
xnor U4245 (N_4245,In_1552,In_1956);
or U4246 (N_4246,In_2936,In_1449);
xnor U4247 (N_4247,In_2752,In_709);
and U4248 (N_4248,In_706,In_2437);
nand U4249 (N_4249,In_85,In_913);
and U4250 (N_4250,In_2830,In_102);
xnor U4251 (N_4251,In_179,In_1255);
xnor U4252 (N_4252,In_539,In_1754);
and U4253 (N_4253,In_1721,In_2836);
and U4254 (N_4254,In_2952,In_25);
nor U4255 (N_4255,In_1993,In_1564);
nand U4256 (N_4256,In_2551,In_2894);
and U4257 (N_4257,In_2318,In_1136);
xor U4258 (N_4258,In_1644,In_1886);
nor U4259 (N_4259,In_2311,In_2995);
xor U4260 (N_4260,In_1871,In_615);
and U4261 (N_4261,In_1975,In_1720);
and U4262 (N_4262,In_486,In_1711);
nand U4263 (N_4263,In_2198,In_245);
or U4264 (N_4264,In_264,In_785);
and U4265 (N_4265,In_2264,In_2663);
nand U4266 (N_4266,In_721,In_2208);
and U4267 (N_4267,In_2831,In_2461);
and U4268 (N_4268,In_814,In_2897);
nor U4269 (N_4269,In_2853,In_2465);
or U4270 (N_4270,In_2771,In_1635);
nor U4271 (N_4271,In_341,In_858);
nand U4272 (N_4272,In_813,In_1970);
xnor U4273 (N_4273,In_2628,In_1168);
and U4274 (N_4274,In_501,In_1348);
or U4275 (N_4275,In_1482,In_909);
nor U4276 (N_4276,In_552,In_146);
and U4277 (N_4277,In_2236,In_576);
nand U4278 (N_4278,In_2989,In_2907);
nor U4279 (N_4279,In_2295,In_1322);
or U4280 (N_4280,In_703,In_124);
and U4281 (N_4281,In_490,In_418);
nor U4282 (N_4282,In_1993,In_1015);
nand U4283 (N_4283,In_1527,In_113);
xor U4284 (N_4284,In_2077,In_1112);
and U4285 (N_4285,In_787,In_666);
and U4286 (N_4286,In_2800,In_1990);
or U4287 (N_4287,In_2958,In_1173);
xnor U4288 (N_4288,In_1074,In_1111);
nand U4289 (N_4289,In_2857,In_1024);
or U4290 (N_4290,In_2479,In_2625);
nand U4291 (N_4291,In_2131,In_2311);
and U4292 (N_4292,In_2740,In_571);
nand U4293 (N_4293,In_1401,In_738);
or U4294 (N_4294,In_2341,In_682);
nor U4295 (N_4295,In_592,In_2657);
or U4296 (N_4296,In_2662,In_1179);
and U4297 (N_4297,In_1693,In_1702);
and U4298 (N_4298,In_2976,In_212);
nand U4299 (N_4299,In_908,In_740);
and U4300 (N_4300,In_1213,In_44);
or U4301 (N_4301,In_1715,In_1427);
nor U4302 (N_4302,In_945,In_972);
and U4303 (N_4303,In_754,In_1265);
xor U4304 (N_4304,In_1242,In_2401);
or U4305 (N_4305,In_1133,In_515);
and U4306 (N_4306,In_2619,In_2410);
nor U4307 (N_4307,In_2668,In_911);
nor U4308 (N_4308,In_1501,In_2288);
nor U4309 (N_4309,In_850,In_2357);
xor U4310 (N_4310,In_1986,In_1671);
and U4311 (N_4311,In_1483,In_2933);
nor U4312 (N_4312,In_1727,In_2170);
or U4313 (N_4313,In_328,In_1762);
or U4314 (N_4314,In_2544,In_2510);
nand U4315 (N_4315,In_2570,In_1871);
nand U4316 (N_4316,In_1066,In_1769);
nand U4317 (N_4317,In_1310,In_606);
and U4318 (N_4318,In_819,In_1013);
nand U4319 (N_4319,In_2732,In_2996);
or U4320 (N_4320,In_6,In_23);
xor U4321 (N_4321,In_1794,In_902);
or U4322 (N_4322,In_2808,In_2575);
nand U4323 (N_4323,In_1566,In_2596);
xor U4324 (N_4324,In_682,In_288);
nor U4325 (N_4325,In_1106,In_1019);
nand U4326 (N_4326,In_2418,In_796);
nor U4327 (N_4327,In_529,In_851);
nor U4328 (N_4328,In_1672,In_1248);
or U4329 (N_4329,In_1922,In_261);
nor U4330 (N_4330,In_2821,In_1233);
and U4331 (N_4331,In_2980,In_507);
or U4332 (N_4332,In_1842,In_1793);
nor U4333 (N_4333,In_2557,In_2604);
nor U4334 (N_4334,In_1782,In_944);
and U4335 (N_4335,In_312,In_2551);
and U4336 (N_4336,In_1909,In_1938);
nand U4337 (N_4337,In_2447,In_1521);
nor U4338 (N_4338,In_1992,In_877);
xor U4339 (N_4339,In_2906,In_1272);
xor U4340 (N_4340,In_2614,In_1390);
and U4341 (N_4341,In_1139,In_812);
or U4342 (N_4342,In_491,In_892);
and U4343 (N_4343,In_1749,In_2102);
nand U4344 (N_4344,In_754,In_747);
or U4345 (N_4345,In_335,In_808);
or U4346 (N_4346,In_890,In_688);
nand U4347 (N_4347,In_804,In_2673);
nand U4348 (N_4348,In_2700,In_516);
and U4349 (N_4349,In_2473,In_1158);
nor U4350 (N_4350,In_1055,In_1129);
or U4351 (N_4351,In_2084,In_2467);
nor U4352 (N_4352,In_831,In_1788);
and U4353 (N_4353,In_1396,In_6);
nor U4354 (N_4354,In_713,In_400);
xor U4355 (N_4355,In_2044,In_2246);
nand U4356 (N_4356,In_1484,In_1557);
nor U4357 (N_4357,In_1725,In_1574);
nor U4358 (N_4358,In_2230,In_155);
or U4359 (N_4359,In_1095,In_477);
or U4360 (N_4360,In_1196,In_503);
nand U4361 (N_4361,In_882,In_265);
and U4362 (N_4362,In_348,In_1746);
nor U4363 (N_4363,In_631,In_732);
and U4364 (N_4364,In_1983,In_777);
or U4365 (N_4365,In_1565,In_2283);
xor U4366 (N_4366,In_963,In_2886);
and U4367 (N_4367,In_2838,In_1979);
and U4368 (N_4368,In_1148,In_2917);
nor U4369 (N_4369,In_637,In_1232);
xnor U4370 (N_4370,In_26,In_1279);
nand U4371 (N_4371,In_1875,In_1302);
nand U4372 (N_4372,In_312,In_1536);
xor U4373 (N_4373,In_2009,In_335);
and U4374 (N_4374,In_2737,In_2002);
nor U4375 (N_4375,In_1564,In_108);
xor U4376 (N_4376,In_2376,In_795);
xnor U4377 (N_4377,In_999,In_2162);
xor U4378 (N_4378,In_2355,In_1118);
nand U4379 (N_4379,In_262,In_2565);
nand U4380 (N_4380,In_759,In_662);
and U4381 (N_4381,In_2937,In_328);
and U4382 (N_4382,In_217,In_1199);
nand U4383 (N_4383,In_454,In_2890);
nor U4384 (N_4384,In_1425,In_2541);
nand U4385 (N_4385,In_629,In_472);
nand U4386 (N_4386,In_116,In_718);
and U4387 (N_4387,In_2103,In_319);
xor U4388 (N_4388,In_2870,In_218);
nor U4389 (N_4389,In_1865,In_2902);
or U4390 (N_4390,In_669,In_2823);
or U4391 (N_4391,In_2830,In_2368);
nand U4392 (N_4392,In_2516,In_403);
and U4393 (N_4393,In_995,In_2651);
xor U4394 (N_4394,In_2154,In_398);
nor U4395 (N_4395,In_2740,In_469);
xnor U4396 (N_4396,In_907,In_2745);
or U4397 (N_4397,In_959,In_2033);
nand U4398 (N_4398,In_800,In_1192);
nand U4399 (N_4399,In_2675,In_1809);
and U4400 (N_4400,In_281,In_1837);
xor U4401 (N_4401,In_612,In_968);
or U4402 (N_4402,In_947,In_1860);
nor U4403 (N_4403,In_1093,In_2319);
nand U4404 (N_4404,In_1873,In_1557);
and U4405 (N_4405,In_464,In_1856);
nor U4406 (N_4406,In_1522,In_117);
nor U4407 (N_4407,In_1874,In_1246);
xnor U4408 (N_4408,In_2303,In_694);
nand U4409 (N_4409,In_179,In_1669);
nand U4410 (N_4410,In_2199,In_2727);
nand U4411 (N_4411,In_1247,In_1100);
and U4412 (N_4412,In_1185,In_2637);
or U4413 (N_4413,In_1689,In_2724);
or U4414 (N_4414,In_2640,In_2218);
or U4415 (N_4415,In_1561,In_347);
xor U4416 (N_4416,In_488,In_2943);
xnor U4417 (N_4417,In_2573,In_1364);
or U4418 (N_4418,In_1417,In_1971);
and U4419 (N_4419,In_508,In_2183);
xnor U4420 (N_4420,In_2863,In_2384);
nor U4421 (N_4421,In_452,In_1944);
nor U4422 (N_4422,In_674,In_1063);
or U4423 (N_4423,In_1024,In_409);
and U4424 (N_4424,In_2020,In_1937);
and U4425 (N_4425,In_2476,In_1569);
xor U4426 (N_4426,In_2897,In_627);
or U4427 (N_4427,In_1996,In_722);
and U4428 (N_4428,In_2413,In_2209);
nand U4429 (N_4429,In_2712,In_426);
or U4430 (N_4430,In_2972,In_2837);
or U4431 (N_4431,In_2896,In_765);
or U4432 (N_4432,In_1243,In_1818);
nor U4433 (N_4433,In_708,In_2126);
and U4434 (N_4434,In_2273,In_2868);
and U4435 (N_4435,In_459,In_1960);
nand U4436 (N_4436,In_1455,In_83);
nor U4437 (N_4437,In_2092,In_2929);
and U4438 (N_4438,In_632,In_1661);
nor U4439 (N_4439,In_1410,In_1910);
xor U4440 (N_4440,In_925,In_2339);
or U4441 (N_4441,In_556,In_2911);
or U4442 (N_4442,In_710,In_1975);
nor U4443 (N_4443,In_1808,In_1421);
or U4444 (N_4444,In_797,In_2562);
and U4445 (N_4445,In_1412,In_2071);
nand U4446 (N_4446,In_168,In_447);
xnor U4447 (N_4447,In_1386,In_2616);
nor U4448 (N_4448,In_1333,In_2810);
nand U4449 (N_4449,In_2932,In_2734);
nor U4450 (N_4450,In_1918,In_2138);
or U4451 (N_4451,In_1570,In_807);
xor U4452 (N_4452,In_1663,In_2458);
or U4453 (N_4453,In_2883,In_510);
nor U4454 (N_4454,In_628,In_2243);
nor U4455 (N_4455,In_2971,In_1863);
or U4456 (N_4456,In_540,In_85);
xor U4457 (N_4457,In_2918,In_23);
xor U4458 (N_4458,In_2070,In_2748);
nor U4459 (N_4459,In_1982,In_1310);
xnor U4460 (N_4460,In_2945,In_207);
nor U4461 (N_4461,In_2897,In_1829);
xor U4462 (N_4462,In_1751,In_2152);
xor U4463 (N_4463,In_2207,In_1961);
and U4464 (N_4464,In_338,In_2122);
nand U4465 (N_4465,In_1876,In_1639);
xnor U4466 (N_4466,In_2961,In_2026);
and U4467 (N_4467,In_1559,In_2388);
or U4468 (N_4468,In_966,In_1026);
nand U4469 (N_4469,In_1329,In_118);
nand U4470 (N_4470,In_1468,In_2232);
or U4471 (N_4471,In_289,In_781);
and U4472 (N_4472,In_439,In_473);
nand U4473 (N_4473,In_1494,In_2525);
nand U4474 (N_4474,In_526,In_2142);
and U4475 (N_4475,In_2326,In_75);
nor U4476 (N_4476,In_1435,In_2831);
or U4477 (N_4477,In_124,In_497);
and U4478 (N_4478,In_1579,In_633);
nand U4479 (N_4479,In_1807,In_996);
and U4480 (N_4480,In_2676,In_585);
xor U4481 (N_4481,In_2402,In_2061);
and U4482 (N_4482,In_2379,In_1122);
xnor U4483 (N_4483,In_2086,In_426);
xor U4484 (N_4484,In_2028,In_165);
and U4485 (N_4485,In_2292,In_2000);
nand U4486 (N_4486,In_2071,In_2506);
or U4487 (N_4487,In_2718,In_2169);
and U4488 (N_4488,In_1617,In_1201);
xnor U4489 (N_4489,In_2192,In_2149);
and U4490 (N_4490,In_906,In_969);
or U4491 (N_4491,In_609,In_1329);
xor U4492 (N_4492,In_1470,In_717);
nor U4493 (N_4493,In_878,In_230);
xor U4494 (N_4494,In_1598,In_2460);
nand U4495 (N_4495,In_1403,In_2805);
nand U4496 (N_4496,In_933,In_2941);
or U4497 (N_4497,In_219,In_2539);
nand U4498 (N_4498,In_596,In_966);
nor U4499 (N_4499,In_2137,In_2831);
or U4500 (N_4500,In_1118,In_2504);
or U4501 (N_4501,In_2453,In_2923);
and U4502 (N_4502,In_2988,In_1740);
or U4503 (N_4503,In_1918,In_1853);
and U4504 (N_4504,In_907,In_132);
nor U4505 (N_4505,In_225,In_151);
nor U4506 (N_4506,In_1553,In_1801);
and U4507 (N_4507,In_1395,In_1610);
and U4508 (N_4508,In_1846,In_2745);
nand U4509 (N_4509,In_2075,In_1283);
or U4510 (N_4510,In_865,In_2829);
nor U4511 (N_4511,In_1668,In_151);
nor U4512 (N_4512,In_2721,In_1112);
xor U4513 (N_4513,In_1609,In_1935);
xor U4514 (N_4514,In_1134,In_214);
nor U4515 (N_4515,In_1757,In_2006);
and U4516 (N_4516,In_792,In_2118);
nor U4517 (N_4517,In_321,In_2998);
nand U4518 (N_4518,In_2433,In_2009);
nand U4519 (N_4519,In_364,In_2796);
nor U4520 (N_4520,In_343,In_1014);
nand U4521 (N_4521,In_916,In_569);
xnor U4522 (N_4522,In_1770,In_2781);
xnor U4523 (N_4523,In_2747,In_367);
nand U4524 (N_4524,In_565,In_132);
nor U4525 (N_4525,In_440,In_1328);
nor U4526 (N_4526,In_1040,In_991);
or U4527 (N_4527,In_584,In_1426);
or U4528 (N_4528,In_1100,In_1387);
or U4529 (N_4529,In_1992,In_2684);
xor U4530 (N_4530,In_362,In_2478);
and U4531 (N_4531,In_2725,In_2858);
nor U4532 (N_4532,In_1993,In_610);
xnor U4533 (N_4533,In_507,In_655);
nor U4534 (N_4534,In_2494,In_1812);
nand U4535 (N_4535,In_2576,In_1695);
nor U4536 (N_4536,In_2029,In_1677);
or U4537 (N_4537,In_1208,In_638);
nand U4538 (N_4538,In_77,In_517);
and U4539 (N_4539,In_28,In_2574);
or U4540 (N_4540,In_1097,In_2514);
nand U4541 (N_4541,In_1595,In_700);
nor U4542 (N_4542,In_399,In_2288);
or U4543 (N_4543,In_261,In_32);
or U4544 (N_4544,In_1073,In_1369);
nand U4545 (N_4545,In_134,In_1706);
nand U4546 (N_4546,In_1032,In_1256);
nor U4547 (N_4547,In_2073,In_2367);
and U4548 (N_4548,In_1252,In_2451);
or U4549 (N_4549,In_1531,In_1689);
xnor U4550 (N_4550,In_769,In_2838);
or U4551 (N_4551,In_127,In_1100);
xnor U4552 (N_4552,In_114,In_1939);
nand U4553 (N_4553,In_2406,In_1928);
xnor U4554 (N_4554,In_1123,In_1320);
or U4555 (N_4555,In_930,In_712);
or U4556 (N_4556,In_2737,In_2947);
or U4557 (N_4557,In_462,In_1525);
xor U4558 (N_4558,In_870,In_2040);
and U4559 (N_4559,In_2656,In_1333);
and U4560 (N_4560,In_2459,In_2708);
or U4561 (N_4561,In_785,In_1235);
nor U4562 (N_4562,In_306,In_422);
nor U4563 (N_4563,In_1862,In_1048);
or U4564 (N_4564,In_2798,In_2535);
or U4565 (N_4565,In_2101,In_2075);
nor U4566 (N_4566,In_2939,In_447);
or U4567 (N_4567,In_338,In_2376);
xor U4568 (N_4568,In_748,In_2793);
xor U4569 (N_4569,In_253,In_1186);
nor U4570 (N_4570,In_2760,In_992);
nor U4571 (N_4571,In_2636,In_209);
nand U4572 (N_4572,In_97,In_720);
nand U4573 (N_4573,In_2623,In_2463);
xnor U4574 (N_4574,In_2711,In_2163);
or U4575 (N_4575,In_1219,In_1888);
and U4576 (N_4576,In_1245,In_920);
nand U4577 (N_4577,In_2945,In_953);
nor U4578 (N_4578,In_1164,In_1042);
xor U4579 (N_4579,In_2429,In_2404);
or U4580 (N_4580,In_2493,In_759);
nand U4581 (N_4581,In_542,In_2474);
nor U4582 (N_4582,In_617,In_2433);
nor U4583 (N_4583,In_991,In_1589);
or U4584 (N_4584,In_748,In_2584);
xor U4585 (N_4585,In_1837,In_151);
nor U4586 (N_4586,In_2760,In_631);
nand U4587 (N_4587,In_959,In_1682);
xnor U4588 (N_4588,In_542,In_1739);
nor U4589 (N_4589,In_1505,In_1441);
xnor U4590 (N_4590,In_2729,In_1733);
xor U4591 (N_4591,In_1791,In_22);
nor U4592 (N_4592,In_876,In_944);
nand U4593 (N_4593,In_1681,In_237);
xor U4594 (N_4594,In_152,In_2939);
nor U4595 (N_4595,In_1896,In_2111);
and U4596 (N_4596,In_2113,In_893);
nand U4597 (N_4597,In_1447,In_1999);
nor U4598 (N_4598,In_312,In_2096);
nand U4599 (N_4599,In_1868,In_672);
and U4600 (N_4600,In_458,In_1764);
xor U4601 (N_4601,In_1581,In_757);
nand U4602 (N_4602,In_2694,In_1764);
and U4603 (N_4603,In_1028,In_411);
and U4604 (N_4604,In_2679,In_371);
or U4605 (N_4605,In_1773,In_2507);
and U4606 (N_4606,In_149,In_2544);
and U4607 (N_4607,In_380,In_1523);
xnor U4608 (N_4608,In_2991,In_2524);
nor U4609 (N_4609,In_550,In_279);
or U4610 (N_4610,In_607,In_2508);
and U4611 (N_4611,In_2371,In_1549);
xor U4612 (N_4612,In_2624,In_2062);
or U4613 (N_4613,In_1717,In_2596);
and U4614 (N_4614,In_674,In_762);
and U4615 (N_4615,In_1044,In_2853);
xor U4616 (N_4616,In_2550,In_1112);
and U4617 (N_4617,In_234,In_420);
nand U4618 (N_4618,In_359,In_1935);
nand U4619 (N_4619,In_534,In_1875);
xor U4620 (N_4620,In_2212,In_2388);
and U4621 (N_4621,In_2474,In_2282);
xor U4622 (N_4622,In_2439,In_239);
and U4623 (N_4623,In_1250,In_229);
nand U4624 (N_4624,In_522,In_2141);
xnor U4625 (N_4625,In_1479,In_1588);
or U4626 (N_4626,In_1534,In_776);
nand U4627 (N_4627,In_694,In_1509);
nor U4628 (N_4628,In_667,In_26);
or U4629 (N_4629,In_1534,In_1895);
nor U4630 (N_4630,In_483,In_795);
nor U4631 (N_4631,In_1998,In_11);
xor U4632 (N_4632,In_1567,In_2875);
or U4633 (N_4633,In_595,In_1458);
and U4634 (N_4634,In_1823,In_305);
and U4635 (N_4635,In_245,In_2115);
or U4636 (N_4636,In_2587,In_230);
and U4637 (N_4637,In_924,In_1534);
nor U4638 (N_4638,In_2424,In_786);
nand U4639 (N_4639,In_2486,In_1716);
or U4640 (N_4640,In_2412,In_1937);
nor U4641 (N_4641,In_1631,In_714);
or U4642 (N_4642,In_1979,In_2241);
nand U4643 (N_4643,In_1708,In_2002);
xnor U4644 (N_4644,In_847,In_592);
and U4645 (N_4645,In_1458,In_1922);
nand U4646 (N_4646,In_2569,In_1193);
or U4647 (N_4647,In_39,In_760);
xnor U4648 (N_4648,In_532,In_506);
xor U4649 (N_4649,In_407,In_1711);
xor U4650 (N_4650,In_2485,In_1514);
nand U4651 (N_4651,In_544,In_1188);
xnor U4652 (N_4652,In_2379,In_36);
nor U4653 (N_4653,In_1244,In_1380);
xnor U4654 (N_4654,In_1144,In_507);
nand U4655 (N_4655,In_1758,In_167);
nor U4656 (N_4656,In_1239,In_1797);
nor U4657 (N_4657,In_247,In_2009);
nand U4658 (N_4658,In_2562,In_677);
or U4659 (N_4659,In_757,In_1720);
xor U4660 (N_4660,In_607,In_1197);
nor U4661 (N_4661,In_1767,In_63);
and U4662 (N_4662,In_810,In_1585);
nand U4663 (N_4663,In_1170,In_2498);
and U4664 (N_4664,In_1518,In_2305);
xor U4665 (N_4665,In_2525,In_1990);
nor U4666 (N_4666,In_1580,In_1851);
nand U4667 (N_4667,In_806,In_2745);
and U4668 (N_4668,In_2403,In_466);
xnor U4669 (N_4669,In_2936,In_464);
and U4670 (N_4670,In_1953,In_1813);
nand U4671 (N_4671,In_179,In_2851);
and U4672 (N_4672,In_392,In_2128);
nor U4673 (N_4673,In_2484,In_2383);
or U4674 (N_4674,In_983,In_481);
nand U4675 (N_4675,In_2365,In_2579);
nor U4676 (N_4676,In_1767,In_418);
xor U4677 (N_4677,In_1137,In_2341);
xnor U4678 (N_4678,In_2352,In_342);
nor U4679 (N_4679,In_340,In_2187);
nor U4680 (N_4680,In_135,In_2495);
nor U4681 (N_4681,In_1079,In_2523);
nand U4682 (N_4682,In_2093,In_1851);
nor U4683 (N_4683,In_1393,In_469);
nand U4684 (N_4684,In_1580,In_1452);
nand U4685 (N_4685,In_1341,In_32);
xor U4686 (N_4686,In_2577,In_2855);
or U4687 (N_4687,In_2962,In_1533);
nor U4688 (N_4688,In_212,In_252);
or U4689 (N_4689,In_1355,In_411);
and U4690 (N_4690,In_52,In_1140);
and U4691 (N_4691,In_2308,In_1069);
nor U4692 (N_4692,In_2371,In_169);
or U4693 (N_4693,In_295,In_856);
xor U4694 (N_4694,In_1670,In_108);
nor U4695 (N_4695,In_2218,In_813);
and U4696 (N_4696,In_230,In_884);
nor U4697 (N_4697,In_1254,In_1401);
and U4698 (N_4698,In_185,In_1629);
nand U4699 (N_4699,In_322,In_225);
and U4700 (N_4700,In_1069,In_2951);
or U4701 (N_4701,In_2962,In_441);
xnor U4702 (N_4702,In_2101,In_2628);
and U4703 (N_4703,In_891,In_2296);
nor U4704 (N_4704,In_2269,In_2773);
nor U4705 (N_4705,In_2919,In_1346);
xnor U4706 (N_4706,In_1521,In_825);
nor U4707 (N_4707,In_2110,In_426);
xnor U4708 (N_4708,In_1130,In_447);
xnor U4709 (N_4709,In_1544,In_440);
nand U4710 (N_4710,In_2866,In_1540);
or U4711 (N_4711,In_495,In_2904);
or U4712 (N_4712,In_2920,In_1076);
or U4713 (N_4713,In_1938,In_181);
nand U4714 (N_4714,In_2167,In_2631);
and U4715 (N_4715,In_2660,In_2109);
or U4716 (N_4716,In_741,In_68);
and U4717 (N_4717,In_127,In_2952);
nor U4718 (N_4718,In_624,In_466);
nand U4719 (N_4719,In_1144,In_927);
nor U4720 (N_4720,In_760,In_1562);
xor U4721 (N_4721,In_2067,In_703);
nand U4722 (N_4722,In_719,In_2586);
or U4723 (N_4723,In_455,In_437);
and U4724 (N_4724,In_18,In_553);
and U4725 (N_4725,In_2597,In_2120);
nor U4726 (N_4726,In_1481,In_1941);
or U4727 (N_4727,In_1988,In_180);
nor U4728 (N_4728,In_2957,In_293);
nor U4729 (N_4729,In_600,In_392);
nor U4730 (N_4730,In_2341,In_2168);
xnor U4731 (N_4731,In_1863,In_2109);
nand U4732 (N_4732,In_1765,In_875);
nor U4733 (N_4733,In_2639,In_2494);
nand U4734 (N_4734,In_172,In_2369);
xor U4735 (N_4735,In_1096,In_1940);
nor U4736 (N_4736,In_1880,In_2482);
nand U4737 (N_4737,In_1953,In_658);
nor U4738 (N_4738,In_1739,In_2914);
or U4739 (N_4739,In_2968,In_856);
nor U4740 (N_4740,In_1881,In_2701);
or U4741 (N_4741,In_310,In_1511);
nand U4742 (N_4742,In_2107,In_2110);
nor U4743 (N_4743,In_2885,In_1682);
or U4744 (N_4744,In_2607,In_2406);
nand U4745 (N_4745,In_1449,In_1186);
or U4746 (N_4746,In_1239,In_2062);
nor U4747 (N_4747,In_1852,In_2597);
xor U4748 (N_4748,In_2012,In_160);
and U4749 (N_4749,In_1562,In_363);
or U4750 (N_4750,In_602,In_1433);
nand U4751 (N_4751,In_227,In_123);
xor U4752 (N_4752,In_2486,In_1329);
nand U4753 (N_4753,In_188,In_621);
or U4754 (N_4754,In_133,In_1337);
nor U4755 (N_4755,In_1407,In_1305);
xnor U4756 (N_4756,In_2406,In_976);
nor U4757 (N_4757,In_610,In_2198);
nand U4758 (N_4758,In_2252,In_2250);
nand U4759 (N_4759,In_907,In_2893);
nand U4760 (N_4760,In_2233,In_1935);
nor U4761 (N_4761,In_61,In_84);
or U4762 (N_4762,In_711,In_2724);
xnor U4763 (N_4763,In_697,In_2249);
nand U4764 (N_4764,In_2916,In_1624);
xor U4765 (N_4765,In_2971,In_2645);
nor U4766 (N_4766,In_876,In_2860);
nor U4767 (N_4767,In_2332,In_1335);
xnor U4768 (N_4768,In_682,In_1853);
or U4769 (N_4769,In_1306,In_993);
and U4770 (N_4770,In_2500,In_2782);
xor U4771 (N_4771,In_452,In_308);
and U4772 (N_4772,In_2843,In_2005);
or U4773 (N_4773,In_2950,In_745);
nand U4774 (N_4774,In_2069,In_2466);
xnor U4775 (N_4775,In_803,In_916);
nor U4776 (N_4776,In_1032,In_1466);
nand U4777 (N_4777,In_2737,In_890);
and U4778 (N_4778,In_2706,In_2683);
and U4779 (N_4779,In_2888,In_2548);
xnor U4780 (N_4780,In_2638,In_406);
or U4781 (N_4781,In_1187,In_991);
xor U4782 (N_4782,In_2470,In_574);
xor U4783 (N_4783,In_2205,In_1741);
or U4784 (N_4784,In_2264,In_326);
xor U4785 (N_4785,In_2530,In_1391);
nand U4786 (N_4786,In_120,In_2121);
nor U4787 (N_4787,In_1665,In_783);
nor U4788 (N_4788,In_1455,In_259);
or U4789 (N_4789,In_1779,In_2602);
nand U4790 (N_4790,In_1687,In_2419);
nand U4791 (N_4791,In_1272,In_527);
xnor U4792 (N_4792,In_1620,In_1846);
nand U4793 (N_4793,In_2150,In_1517);
and U4794 (N_4794,In_396,In_1573);
nor U4795 (N_4795,In_2344,In_500);
nand U4796 (N_4796,In_550,In_1689);
nand U4797 (N_4797,In_2072,In_2749);
xnor U4798 (N_4798,In_2535,In_2814);
and U4799 (N_4799,In_1679,In_116);
xor U4800 (N_4800,In_941,In_1135);
nor U4801 (N_4801,In_2833,In_706);
and U4802 (N_4802,In_1902,In_268);
nor U4803 (N_4803,In_596,In_2547);
and U4804 (N_4804,In_1179,In_2483);
xor U4805 (N_4805,In_153,In_2111);
or U4806 (N_4806,In_766,In_2579);
nand U4807 (N_4807,In_2020,In_467);
nor U4808 (N_4808,In_1548,In_1564);
and U4809 (N_4809,In_2005,In_1324);
and U4810 (N_4810,In_1171,In_1160);
and U4811 (N_4811,In_2756,In_2291);
nand U4812 (N_4812,In_577,In_1969);
xor U4813 (N_4813,In_2419,In_191);
and U4814 (N_4814,In_2385,In_1574);
nand U4815 (N_4815,In_0,In_1004);
xnor U4816 (N_4816,In_177,In_1385);
or U4817 (N_4817,In_1508,In_1373);
and U4818 (N_4818,In_2742,In_788);
nor U4819 (N_4819,In_2347,In_328);
and U4820 (N_4820,In_133,In_2140);
nor U4821 (N_4821,In_196,In_1716);
or U4822 (N_4822,In_2114,In_1914);
or U4823 (N_4823,In_1676,In_2354);
nor U4824 (N_4824,In_776,In_124);
and U4825 (N_4825,In_844,In_1445);
nand U4826 (N_4826,In_2560,In_633);
xor U4827 (N_4827,In_61,In_342);
nor U4828 (N_4828,In_2372,In_1533);
and U4829 (N_4829,In_899,In_2245);
and U4830 (N_4830,In_2394,In_2534);
nor U4831 (N_4831,In_687,In_2086);
nor U4832 (N_4832,In_2668,In_2989);
and U4833 (N_4833,In_1845,In_2228);
xnor U4834 (N_4834,In_2077,In_800);
nor U4835 (N_4835,In_2082,In_2069);
nor U4836 (N_4836,In_2478,In_1676);
xor U4837 (N_4837,In_838,In_44);
nor U4838 (N_4838,In_1148,In_2878);
xnor U4839 (N_4839,In_1211,In_1924);
nor U4840 (N_4840,In_1736,In_648);
or U4841 (N_4841,In_530,In_1652);
or U4842 (N_4842,In_1664,In_1411);
or U4843 (N_4843,In_1188,In_940);
or U4844 (N_4844,In_1657,In_382);
nand U4845 (N_4845,In_60,In_240);
or U4846 (N_4846,In_316,In_2249);
nor U4847 (N_4847,In_1316,In_1317);
nand U4848 (N_4848,In_2986,In_2860);
nand U4849 (N_4849,In_905,In_1956);
and U4850 (N_4850,In_314,In_680);
nor U4851 (N_4851,In_2609,In_304);
nand U4852 (N_4852,In_2971,In_530);
and U4853 (N_4853,In_375,In_2829);
nand U4854 (N_4854,In_1980,In_2156);
nand U4855 (N_4855,In_1395,In_2423);
nor U4856 (N_4856,In_2729,In_447);
xor U4857 (N_4857,In_1644,In_809);
xnor U4858 (N_4858,In_2796,In_2515);
nor U4859 (N_4859,In_336,In_1176);
xnor U4860 (N_4860,In_1786,In_2082);
nand U4861 (N_4861,In_1406,In_151);
or U4862 (N_4862,In_459,In_1959);
and U4863 (N_4863,In_2178,In_66);
nand U4864 (N_4864,In_343,In_800);
xnor U4865 (N_4865,In_2605,In_273);
or U4866 (N_4866,In_804,In_190);
or U4867 (N_4867,In_2793,In_2634);
or U4868 (N_4868,In_409,In_2403);
xnor U4869 (N_4869,In_1167,In_2066);
or U4870 (N_4870,In_714,In_1135);
xor U4871 (N_4871,In_1781,In_1160);
nor U4872 (N_4872,In_2960,In_2629);
and U4873 (N_4873,In_438,In_1039);
and U4874 (N_4874,In_139,In_786);
nand U4875 (N_4875,In_2598,In_205);
nand U4876 (N_4876,In_233,In_1310);
nor U4877 (N_4877,In_993,In_370);
or U4878 (N_4878,In_1532,In_698);
nand U4879 (N_4879,In_1633,In_2763);
nand U4880 (N_4880,In_2520,In_653);
or U4881 (N_4881,In_598,In_69);
or U4882 (N_4882,In_1774,In_2602);
xor U4883 (N_4883,In_1839,In_1795);
and U4884 (N_4884,In_314,In_918);
nor U4885 (N_4885,In_306,In_1050);
or U4886 (N_4886,In_2202,In_1488);
nand U4887 (N_4887,In_1527,In_2970);
xor U4888 (N_4888,In_20,In_2905);
xor U4889 (N_4889,In_1896,In_2425);
and U4890 (N_4890,In_2909,In_1589);
xor U4891 (N_4891,In_1897,In_1856);
nand U4892 (N_4892,In_1800,In_2972);
xnor U4893 (N_4893,In_1037,In_317);
nand U4894 (N_4894,In_2665,In_30);
or U4895 (N_4895,In_1831,In_2079);
or U4896 (N_4896,In_2587,In_1079);
nand U4897 (N_4897,In_939,In_1751);
xnor U4898 (N_4898,In_1562,In_2197);
nand U4899 (N_4899,In_463,In_459);
and U4900 (N_4900,In_1346,In_660);
or U4901 (N_4901,In_1149,In_1362);
nor U4902 (N_4902,In_2920,In_441);
and U4903 (N_4903,In_2333,In_2389);
nand U4904 (N_4904,In_211,In_1229);
nor U4905 (N_4905,In_2892,In_2145);
nand U4906 (N_4906,In_2820,In_509);
or U4907 (N_4907,In_2442,In_2868);
or U4908 (N_4908,In_711,In_2305);
and U4909 (N_4909,In_2490,In_469);
or U4910 (N_4910,In_1672,In_2747);
nor U4911 (N_4911,In_1514,In_248);
or U4912 (N_4912,In_1338,In_2149);
xnor U4913 (N_4913,In_1968,In_929);
xor U4914 (N_4914,In_883,In_707);
and U4915 (N_4915,In_2727,In_2856);
and U4916 (N_4916,In_1625,In_1365);
and U4917 (N_4917,In_1497,In_1080);
xnor U4918 (N_4918,In_910,In_1127);
nor U4919 (N_4919,In_2298,In_443);
nand U4920 (N_4920,In_2380,In_2009);
nor U4921 (N_4921,In_294,In_1980);
nand U4922 (N_4922,In_619,In_189);
nor U4923 (N_4923,In_1417,In_2915);
nand U4924 (N_4924,In_1847,In_691);
nor U4925 (N_4925,In_1734,In_2864);
or U4926 (N_4926,In_2129,In_317);
and U4927 (N_4927,In_2680,In_39);
and U4928 (N_4928,In_1421,In_1576);
xnor U4929 (N_4929,In_215,In_2624);
nor U4930 (N_4930,In_1841,In_1570);
nor U4931 (N_4931,In_904,In_851);
nor U4932 (N_4932,In_2647,In_791);
nand U4933 (N_4933,In_1206,In_1836);
nand U4934 (N_4934,In_1431,In_1283);
or U4935 (N_4935,In_1475,In_684);
or U4936 (N_4936,In_2936,In_176);
nor U4937 (N_4937,In_1786,In_2076);
and U4938 (N_4938,In_2546,In_1688);
and U4939 (N_4939,In_838,In_2629);
xor U4940 (N_4940,In_478,In_1703);
and U4941 (N_4941,In_2193,In_1514);
or U4942 (N_4942,In_195,In_2663);
xor U4943 (N_4943,In_2907,In_2923);
nand U4944 (N_4944,In_2103,In_1782);
nor U4945 (N_4945,In_460,In_1046);
and U4946 (N_4946,In_368,In_548);
xor U4947 (N_4947,In_2454,In_2893);
nor U4948 (N_4948,In_268,In_884);
nor U4949 (N_4949,In_2350,In_2265);
xor U4950 (N_4950,In_2157,In_2621);
nor U4951 (N_4951,In_2079,In_598);
and U4952 (N_4952,In_498,In_975);
nor U4953 (N_4953,In_2003,In_1484);
nor U4954 (N_4954,In_2003,In_597);
and U4955 (N_4955,In_328,In_2336);
nand U4956 (N_4956,In_380,In_2614);
or U4957 (N_4957,In_1569,In_348);
xor U4958 (N_4958,In_2402,In_668);
nand U4959 (N_4959,In_1359,In_340);
or U4960 (N_4960,In_599,In_560);
nor U4961 (N_4961,In_991,In_1741);
and U4962 (N_4962,In_1464,In_919);
nand U4963 (N_4963,In_937,In_949);
nand U4964 (N_4964,In_1239,In_1428);
or U4965 (N_4965,In_1831,In_2081);
nand U4966 (N_4966,In_2279,In_2844);
nand U4967 (N_4967,In_2297,In_1455);
and U4968 (N_4968,In_1308,In_2103);
xnor U4969 (N_4969,In_2525,In_130);
nor U4970 (N_4970,In_1562,In_2294);
nand U4971 (N_4971,In_1528,In_2605);
or U4972 (N_4972,In_2671,In_1736);
nand U4973 (N_4973,In_1583,In_804);
and U4974 (N_4974,In_45,In_1532);
xor U4975 (N_4975,In_1513,In_2603);
nand U4976 (N_4976,In_1088,In_820);
xor U4977 (N_4977,In_151,In_2988);
xor U4978 (N_4978,In_272,In_2564);
and U4979 (N_4979,In_1407,In_1000);
nand U4980 (N_4980,In_2039,In_2502);
or U4981 (N_4981,In_766,In_1009);
nand U4982 (N_4982,In_1641,In_1373);
nor U4983 (N_4983,In_123,In_1558);
nor U4984 (N_4984,In_2404,In_271);
or U4985 (N_4985,In_2359,In_139);
nand U4986 (N_4986,In_2805,In_2406);
nand U4987 (N_4987,In_349,In_1258);
or U4988 (N_4988,In_2462,In_2078);
xnor U4989 (N_4989,In_2342,In_709);
or U4990 (N_4990,In_905,In_1823);
nand U4991 (N_4991,In_1075,In_1567);
or U4992 (N_4992,In_176,In_146);
xnor U4993 (N_4993,In_339,In_2193);
nand U4994 (N_4994,In_1731,In_1344);
and U4995 (N_4995,In_234,In_1123);
nor U4996 (N_4996,In_1419,In_2216);
and U4997 (N_4997,In_833,In_2511);
or U4998 (N_4998,In_2911,In_153);
nor U4999 (N_4999,In_1887,In_287);
nor U5000 (N_5000,N_1302,N_3511);
nand U5001 (N_5001,N_4015,N_926);
nand U5002 (N_5002,N_610,N_2174);
nor U5003 (N_5003,N_4355,N_178);
xor U5004 (N_5004,N_2370,N_2221);
and U5005 (N_5005,N_2860,N_2003);
and U5006 (N_5006,N_268,N_1744);
or U5007 (N_5007,N_1992,N_75);
xor U5008 (N_5008,N_1211,N_3704);
nor U5009 (N_5009,N_4669,N_3617);
nand U5010 (N_5010,N_2757,N_3693);
xnor U5011 (N_5011,N_130,N_2711);
nor U5012 (N_5012,N_2312,N_4401);
xor U5013 (N_5013,N_4678,N_2704);
nand U5014 (N_5014,N_337,N_778);
or U5015 (N_5015,N_2377,N_2978);
nor U5016 (N_5016,N_733,N_4045);
or U5017 (N_5017,N_4309,N_4783);
nand U5018 (N_5018,N_4567,N_2976);
and U5019 (N_5019,N_3436,N_625);
nand U5020 (N_5020,N_2910,N_2036);
and U5021 (N_5021,N_3373,N_1672);
or U5022 (N_5022,N_648,N_3087);
and U5023 (N_5023,N_3493,N_1130);
nand U5024 (N_5024,N_1655,N_1541);
xnor U5025 (N_5025,N_1768,N_464);
nor U5026 (N_5026,N_3946,N_4634);
nand U5027 (N_5027,N_1021,N_2145);
or U5028 (N_5028,N_4294,N_2004);
or U5029 (N_5029,N_478,N_93);
nand U5030 (N_5030,N_3602,N_3925);
nand U5031 (N_5031,N_3923,N_3090);
nand U5032 (N_5032,N_2201,N_3042);
nand U5033 (N_5033,N_3473,N_3926);
and U5034 (N_5034,N_479,N_4810);
nand U5035 (N_5035,N_2208,N_2094);
and U5036 (N_5036,N_1917,N_2000);
and U5037 (N_5037,N_1382,N_848);
or U5038 (N_5038,N_1072,N_3469);
nor U5039 (N_5039,N_3346,N_4474);
nor U5040 (N_5040,N_1464,N_4137);
and U5041 (N_5041,N_4532,N_3124);
nand U5042 (N_5042,N_2360,N_2538);
and U5043 (N_5043,N_730,N_215);
or U5044 (N_5044,N_3580,N_3609);
xor U5045 (N_5045,N_1595,N_2886);
nand U5046 (N_5046,N_3379,N_1848);
nand U5047 (N_5047,N_1200,N_600);
or U5048 (N_5048,N_45,N_2631);
xor U5049 (N_5049,N_1964,N_737);
nand U5050 (N_5050,N_4027,N_1827);
xor U5051 (N_5051,N_4461,N_4488);
nand U5052 (N_5052,N_516,N_552);
or U5053 (N_5053,N_2903,N_1323);
nor U5054 (N_5054,N_4417,N_3355);
nor U5055 (N_5055,N_4550,N_3526);
nor U5056 (N_5056,N_3225,N_4814);
and U5057 (N_5057,N_1189,N_3770);
nor U5058 (N_5058,N_1248,N_121);
nor U5059 (N_5059,N_4667,N_314);
nand U5060 (N_5060,N_2455,N_4859);
nor U5061 (N_5061,N_4469,N_3262);
xor U5062 (N_5062,N_517,N_3534);
nand U5063 (N_5063,N_2409,N_3316);
or U5064 (N_5064,N_3447,N_2683);
xor U5065 (N_5065,N_4130,N_1071);
xnor U5066 (N_5066,N_2369,N_3688);
nor U5067 (N_5067,N_1242,N_3052);
nor U5068 (N_5068,N_3993,N_3948);
nand U5069 (N_5069,N_1013,N_294);
xor U5070 (N_5070,N_3778,N_4860);
nand U5071 (N_5071,N_3114,N_1643);
xor U5072 (N_5072,N_3844,N_1823);
nand U5073 (N_5073,N_4920,N_520);
and U5074 (N_5074,N_638,N_1257);
nor U5075 (N_5075,N_3332,N_2822);
xnor U5076 (N_5076,N_628,N_117);
or U5077 (N_5077,N_2542,N_1586);
nor U5078 (N_5078,N_1250,N_2143);
xor U5079 (N_5079,N_4371,N_1220);
and U5080 (N_5080,N_3480,N_3737);
nor U5081 (N_5081,N_781,N_4100);
or U5082 (N_5082,N_2566,N_2823);
or U5083 (N_5083,N_474,N_4608);
and U5084 (N_5084,N_3408,N_3587);
xnor U5085 (N_5085,N_1562,N_3924);
xor U5086 (N_5086,N_3307,N_4482);
or U5087 (N_5087,N_2375,N_4002);
nor U5088 (N_5088,N_2610,N_1689);
nand U5089 (N_5089,N_3951,N_1703);
or U5090 (N_5090,N_156,N_3339);
xor U5091 (N_5091,N_1022,N_2824);
and U5092 (N_5092,N_2942,N_874);
nand U5093 (N_5093,N_1237,N_1261);
nor U5094 (N_5094,N_1721,N_3936);
nor U5095 (N_5095,N_3848,N_1572);
nand U5096 (N_5096,N_4381,N_2156);
nand U5097 (N_5097,N_2282,N_4871);
nor U5098 (N_5098,N_1367,N_3880);
or U5099 (N_5099,N_4263,N_2674);
nor U5100 (N_5100,N_2906,N_2393);
nand U5101 (N_5101,N_2947,N_1331);
and U5102 (N_5102,N_2401,N_272);
nand U5103 (N_5103,N_2792,N_1436);
or U5104 (N_5104,N_2560,N_4108);
xor U5105 (N_5105,N_2698,N_4940);
xnor U5106 (N_5106,N_3930,N_1707);
nand U5107 (N_5107,N_1110,N_798);
nand U5108 (N_5108,N_3348,N_4657);
and U5109 (N_5109,N_1664,N_4833);
and U5110 (N_5110,N_2622,N_3746);
or U5111 (N_5111,N_4362,N_3264);
nand U5112 (N_5112,N_3655,N_745);
nand U5113 (N_5113,N_2289,N_4049);
and U5114 (N_5114,N_546,N_3120);
nand U5115 (N_5115,N_3518,N_1970);
xnor U5116 (N_5116,N_3658,N_3873);
and U5117 (N_5117,N_468,N_4511);
nor U5118 (N_5118,N_2376,N_460);
or U5119 (N_5119,N_3767,N_2742);
nor U5120 (N_5120,N_1428,N_3822);
or U5121 (N_5121,N_328,N_4942);
nor U5122 (N_5122,N_538,N_4785);
and U5123 (N_5123,N_4772,N_2654);
nor U5124 (N_5124,N_4046,N_168);
nor U5125 (N_5125,N_4624,N_1438);
xor U5126 (N_5126,N_21,N_870);
xnor U5127 (N_5127,N_2684,N_2091);
or U5128 (N_5128,N_2160,N_1872);
and U5129 (N_5129,N_4808,N_3649);
or U5130 (N_5130,N_2058,N_4518);
xnor U5131 (N_5131,N_1074,N_3825);
nor U5132 (N_5132,N_1080,N_2520);
and U5133 (N_5133,N_1390,N_4821);
nor U5134 (N_5134,N_2863,N_4481);
xnor U5135 (N_5135,N_476,N_2275);
and U5136 (N_5136,N_4733,N_4062);
nand U5137 (N_5137,N_3523,N_2827);
nand U5138 (N_5138,N_4190,N_3338);
xor U5139 (N_5139,N_649,N_1980);
nor U5140 (N_5140,N_3131,N_4295);
nor U5141 (N_5141,N_3459,N_2052);
nand U5142 (N_5142,N_2279,N_1141);
nand U5143 (N_5143,N_3254,N_1136);
nor U5144 (N_5144,N_3678,N_4026);
nand U5145 (N_5145,N_4186,N_4575);
or U5146 (N_5146,N_4463,N_4233);
nand U5147 (N_5147,N_1949,N_3178);
nor U5148 (N_5148,N_3369,N_2859);
or U5149 (N_5149,N_2551,N_3017);
and U5150 (N_5150,N_136,N_3078);
and U5151 (N_5151,N_2534,N_2709);
xnor U5152 (N_5152,N_3166,N_2999);
xnor U5153 (N_5153,N_2172,N_1083);
and U5154 (N_5154,N_4569,N_3304);
or U5155 (N_5155,N_2653,N_2294);
and U5156 (N_5156,N_4626,N_1737);
and U5157 (N_5157,N_1799,N_3870);
nand U5158 (N_5158,N_1445,N_3639);
and U5159 (N_5159,N_2920,N_2723);
xor U5160 (N_5160,N_1231,N_4255);
or U5161 (N_5161,N_3249,N_2006);
xnor U5162 (N_5162,N_1733,N_2437);
nor U5163 (N_5163,N_761,N_1603);
nand U5164 (N_5164,N_3489,N_262);
and U5165 (N_5165,N_3100,N_3618);
and U5166 (N_5166,N_2883,N_1521);
nand U5167 (N_5167,N_4987,N_4741);
xnor U5168 (N_5168,N_3950,N_2103);
or U5169 (N_5169,N_1734,N_2295);
xnor U5170 (N_5170,N_2801,N_2936);
xnor U5171 (N_5171,N_2894,N_2271);
and U5172 (N_5172,N_1588,N_4414);
nor U5173 (N_5173,N_2780,N_1808);
or U5174 (N_5174,N_3540,N_364);
or U5175 (N_5175,N_176,N_4531);
and U5176 (N_5176,N_373,N_4841);
nor U5177 (N_5177,N_3206,N_1125);
xnor U5178 (N_5178,N_4494,N_1955);
nor U5179 (N_5179,N_1801,N_4755);
nand U5180 (N_5180,N_1860,N_1565);
or U5181 (N_5181,N_442,N_4891);
nor U5182 (N_5182,N_1239,N_2820);
xnor U5183 (N_5183,N_3214,N_303);
xor U5184 (N_5184,N_2268,N_3958);
nor U5185 (N_5185,N_128,N_4252);
and U5186 (N_5186,N_564,N_1000);
nor U5187 (N_5187,N_3392,N_2232);
nor U5188 (N_5188,N_883,N_1101);
nor U5189 (N_5189,N_4257,N_1166);
nor U5190 (N_5190,N_4195,N_1753);
nand U5191 (N_5191,N_3119,N_3491);
nand U5192 (N_5192,N_1037,N_4903);
or U5193 (N_5193,N_3508,N_4948);
xor U5194 (N_5194,N_4549,N_456);
or U5195 (N_5195,N_3170,N_639);
and U5196 (N_5196,N_4870,N_1989);
or U5197 (N_5197,N_3322,N_2620);
nor U5198 (N_5198,N_2461,N_2380);
nand U5199 (N_5199,N_4435,N_1224);
and U5200 (N_5200,N_36,N_938);
nor U5201 (N_5201,N_680,N_1965);
nand U5202 (N_5202,N_3967,N_2239);
xor U5203 (N_5203,N_1954,N_4129);
nand U5204 (N_5204,N_4796,N_3673);
or U5205 (N_5205,N_2465,N_2356);
or U5206 (N_5206,N_772,N_3033);
xnor U5207 (N_5207,N_4054,N_2794);
xor U5208 (N_5208,N_1444,N_2612);
nor U5209 (N_5209,N_1271,N_2146);
nor U5210 (N_5210,N_821,N_1133);
or U5211 (N_5211,N_1591,N_3838);
and U5212 (N_5212,N_192,N_4168);
nand U5213 (N_5213,N_2988,N_3195);
or U5214 (N_5214,N_4237,N_2755);
nor U5215 (N_5215,N_1215,N_1184);
and U5216 (N_5216,N_487,N_3629);
or U5217 (N_5217,N_1709,N_3986);
and U5218 (N_5218,N_3600,N_1629);
and U5219 (N_5219,N_1047,N_1063);
nand U5220 (N_5220,N_1310,N_911);
nor U5221 (N_5221,N_2114,N_2243);
xor U5222 (N_5222,N_247,N_918);
nand U5223 (N_5223,N_3748,N_4153);
nor U5224 (N_5224,N_4666,N_1792);
or U5225 (N_5225,N_4754,N_1661);
or U5226 (N_5226,N_2413,N_1963);
or U5227 (N_5227,N_4197,N_3287);
nor U5228 (N_5228,N_1598,N_4932);
and U5229 (N_5229,N_742,N_3147);
nand U5230 (N_5230,N_3871,N_3862);
and U5231 (N_5231,N_4019,N_3347);
nand U5232 (N_5232,N_1087,N_4770);
and U5233 (N_5233,N_4444,N_308);
or U5234 (N_5234,N_4544,N_1175);
or U5235 (N_5235,N_1086,N_2513);
nor U5236 (N_5236,N_1046,N_1693);
xnor U5237 (N_5237,N_4954,N_3957);
or U5238 (N_5238,N_2652,N_1722);
nor U5239 (N_5239,N_2269,N_3446);
nand U5240 (N_5240,N_397,N_527);
xnor U5241 (N_5241,N_519,N_713);
xor U5242 (N_5242,N_1662,N_2442);
nor U5243 (N_5243,N_1285,N_1622);
and U5244 (N_5244,N_3468,N_4646);
nand U5245 (N_5245,N_2726,N_3814);
or U5246 (N_5246,N_774,N_979);
and U5247 (N_5247,N_3697,N_4024);
and U5248 (N_5248,N_1442,N_350);
xor U5249 (N_5249,N_3653,N_4877);
and U5250 (N_5250,N_214,N_2518);
and U5251 (N_5251,N_1781,N_640);
nand U5252 (N_5252,N_2362,N_2196);
or U5253 (N_5253,N_3519,N_4057);
nor U5254 (N_5254,N_1933,N_3263);
or U5255 (N_5255,N_270,N_170);
nor U5256 (N_5256,N_857,N_2582);
or U5257 (N_5257,N_1164,N_627);
or U5258 (N_5258,N_3572,N_4312);
nand U5259 (N_5259,N_4457,N_4768);
nand U5260 (N_5260,N_4445,N_1191);
or U5261 (N_5261,N_593,N_431);
or U5262 (N_5262,N_1497,N_4647);
nor U5263 (N_5263,N_4105,N_2429);
nor U5264 (N_5264,N_4798,N_1551);
xor U5265 (N_5265,N_4816,N_1104);
nor U5266 (N_5266,N_2167,N_380);
or U5267 (N_5267,N_4286,N_318);
and U5268 (N_5268,N_396,N_165);
or U5269 (N_5269,N_1201,N_3173);
nand U5270 (N_5270,N_271,N_1490);
and U5271 (N_5271,N_2479,N_1563);
or U5272 (N_5272,N_780,N_2186);
or U5273 (N_5273,N_2825,N_3550);
or U5274 (N_5274,N_394,N_1324);
xnor U5275 (N_5275,N_199,N_1391);
nand U5276 (N_5276,N_1385,N_788);
and U5277 (N_5277,N_3516,N_1400);
or U5278 (N_5278,N_205,N_2241);
nand U5279 (N_5279,N_2946,N_1420);
and U5280 (N_5280,N_3380,N_4432);
and U5281 (N_5281,N_3261,N_2948);
or U5282 (N_5282,N_3148,N_1472);
nand U5283 (N_5283,N_1301,N_1359);
xor U5284 (N_5284,N_2206,N_3125);
nand U5285 (N_5285,N_4075,N_177);
nand U5286 (N_5286,N_70,N_1064);
nor U5287 (N_5287,N_2943,N_4344);
xnor U5288 (N_5288,N_3185,N_2477);
nor U5289 (N_5289,N_3244,N_2561);
nor U5290 (N_5290,N_602,N_4365);
nor U5291 (N_5291,N_4221,N_3418);
or U5292 (N_5292,N_974,N_3537);
nor U5293 (N_5293,N_2682,N_1557);
and U5294 (N_5294,N_2641,N_776);
nand U5295 (N_5295,N_336,N_2981);
nor U5296 (N_5296,N_2423,N_4815);
nor U5297 (N_5297,N_4410,N_2795);
and U5298 (N_5298,N_507,N_881);
xnor U5299 (N_5299,N_2556,N_2990);
nor U5300 (N_5300,N_163,N_4340);
nand U5301 (N_5301,N_3635,N_2035);
xnor U5302 (N_5302,N_1608,N_4665);
or U5303 (N_5303,N_2591,N_2080);
or U5304 (N_5304,N_3135,N_3411);
xnor U5305 (N_5305,N_2592,N_172);
xnor U5306 (N_5306,N_1876,N_825);
nand U5307 (N_5307,N_4698,N_69);
or U5308 (N_5308,N_1415,N_3005);
nor U5309 (N_5309,N_1748,N_2899);
nor U5310 (N_5310,N_560,N_966);
or U5311 (N_5311,N_171,N_2882);
or U5312 (N_5312,N_2685,N_2833);
and U5313 (N_5313,N_55,N_2902);
nor U5314 (N_5314,N_1810,N_530);
nor U5315 (N_5315,N_2905,N_2662);
or U5316 (N_5316,N_2963,N_2300);
nor U5317 (N_5317,N_721,N_2473);
or U5318 (N_5318,N_2419,N_239);
xor U5319 (N_5319,N_945,N_3077);
or U5320 (N_5320,N_186,N_1247);
nor U5321 (N_5321,N_1784,N_3758);
and U5322 (N_5322,N_4882,N_3012);
or U5323 (N_5323,N_1858,N_349);
nand U5324 (N_5324,N_4319,N_2298);
xnor U5325 (N_5325,N_710,N_1407);
or U5326 (N_5326,N_1577,N_1619);
and U5327 (N_5327,N_412,N_3318);
xor U5328 (N_5328,N_2672,N_2839);
and U5329 (N_5329,N_1544,N_1199);
and U5330 (N_5330,N_2569,N_3744);
or U5331 (N_5331,N_1704,N_3359);
xor U5332 (N_5332,N_609,N_2418);
xnor U5333 (N_5333,N_2828,N_1156);
and U5334 (N_5334,N_4602,N_1584);
and U5335 (N_5335,N_1179,N_2655);
or U5336 (N_5336,N_376,N_1322);
or U5337 (N_5337,N_3402,N_3513);
nand U5338 (N_5338,N_1791,N_4095);
xnor U5339 (N_5339,N_4743,N_1170);
and U5340 (N_5340,N_2326,N_889);
or U5341 (N_5341,N_3046,N_4178);
nand U5342 (N_5342,N_962,N_2789);
xor U5343 (N_5343,N_1507,N_3200);
xnor U5344 (N_5344,N_2308,N_3426);
nor U5345 (N_5345,N_4889,N_4979);
nand U5346 (N_5346,N_2132,N_4396);
nand U5347 (N_5347,N_3622,N_1355);
nor U5348 (N_5348,N_722,N_2032);
nor U5349 (N_5349,N_3073,N_2918);
xor U5350 (N_5350,N_3689,N_1885);
or U5351 (N_5351,N_3080,N_2811);
nand U5352 (N_5352,N_2885,N_3840);
and U5353 (N_5353,N_559,N_2272);
xnor U5354 (N_5354,N_280,N_3495);
nand U5355 (N_5355,N_1864,N_461);
nand U5356 (N_5356,N_4266,N_3109);
and U5357 (N_5357,N_3414,N_584);
nand U5358 (N_5358,N_1216,N_3500);
or U5359 (N_5359,N_1238,N_4961);
and U5360 (N_5360,N_497,N_794);
or U5361 (N_5361,N_668,N_4538);
or U5362 (N_5362,N_2666,N_4310);
and U5363 (N_5363,N_3417,N_4786);
nor U5364 (N_5364,N_3103,N_4314);
xnor U5365 (N_5365,N_3247,N_2266);
or U5366 (N_5366,N_3852,N_3820);
nand U5367 (N_5367,N_985,N_2007);
or U5368 (N_5368,N_2987,N_1099);
nor U5369 (N_5369,N_4572,N_1794);
nand U5370 (N_5370,N_2624,N_1062);
nor U5371 (N_5371,N_3142,N_4323);
nor U5372 (N_5372,N_1399,N_2445);
nor U5373 (N_5373,N_1480,N_352);
xor U5374 (N_5374,N_3023,N_2816);
and U5375 (N_5375,N_882,N_3145);
nor U5376 (N_5376,N_4548,N_2667);
and U5377 (N_5377,N_3788,N_2057);
and U5378 (N_5378,N_2482,N_550);
nand U5379 (N_5379,N_1030,N_1460);
nor U5380 (N_5380,N_4804,N_3834);
xor U5381 (N_5381,N_1082,N_2665);
or U5382 (N_5382,N_707,N_3809);
and U5383 (N_5383,N_2777,N_106);
nor U5384 (N_5384,N_1815,N_4724);
or U5385 (N_5385,N_365,N_3096);
nor U5386 (N_5386,N_3352,N_4510);
and U5387 (N_5387,N_1764,N_2689);
xor U5388 (N_5388,N_4397,N_1633);
or U5389 (N_5389,N_2022,N_2077);
nor U5390 (N_5390,N_179,N_315);
nand U5391 (N_5391,N_1380,N_3899);
or U5392 (N_5392,N_4977,N_3740);
and U5393 (N_5393,N_2770,N_971);
and U5394 (N_5394,N_3793,N_2993);
xor U5395 (N_5395,N_4499,N_673);
or U5396 (N_5396,N_4307,N_3037);
and U5397 (N_5397,N_4235,N_4308);
and U5398 (N_5398,N_4101,N_144);
nand U5399 (N_5399,N_2932,N_44);
xnor U5400 (N_5400,N_1081,N_1332);
and U5401 (N_5401,N_3736,N_1576);
or U5402 (N_5402,N_1932,N_3279);
xnor U5403 (N_5403,N_3633,N_2512);
or U5404 (N_5404,N_4686,N_3596);
nand U5405 (N_5405,N_2962,N_3860);
or U5406 (N_5406,N_4029,N_1494);
or U5407 (N_5407,N_3623,N_3503);
nor U5408 (N_5408,N_3427,N_4082);
or U5409 (N_5409,N_4892,N_3471);
or U5410 (N_5410,N_450,N_4228);
nor U5411 (N_5411,N_2029,N_2244);
xor U5412 (N_5412,N_3014,N_3413);
and U5413 (N_5413,N_1127,N_978);
nand U5414 (N_5414,N_3309,N_3226);
nor U5415 (N_5415,N_611,N_3654);
or U5416 (N_5416,N_541,N_4507);
nor U5417 (N_5417,N_4452,N_4150);
or U5418 (N_5418,N_3533,N_3458);
and U5419 (N_5419,N_3779,N_1416);
xor U5420 (N_5420,N_4144,N_1153);
or U5421 (N_5421,N_2994,N_3650);
xor U5422 (N_5422,N_2412,N_1666);
xnor U5423 (N_5423,N_4421,N_2916);
or U5424 (N_5424,N_1979,N_3430);
or U5425 (N_5425,N_196,N_3849);
nor U5426 (N_5426,N_2112,N_1326);
and U5427 (N_5427,N_1983,N_3905);
xor U5428 (N_5428,N_4127,N_4935);
and U5429 (N_5429,N_3524,N_3105);
and U5430 (N_5430,N_1431,N_2469);
and U5431 (N_5431,N_207,N_2807);
or U5432 (N_5432,N_3079,N_2152);
xor U5433 (N_5433,N_1831,N_1800);
nor U5434 (N_5434,N_1812,N_3591);
and U5435 (N_5435,N_4508,N_4876);
xnor U5436 (N_5436,N_2304,N_3107);
xnor U5437 (N_5437,N_727,N_1531);
xor U5438 (N_5438,N_3084,N_162);
and U5439 (N_5439,N_2390,N_3889);
nor U5440 (N_5440,N_980,N_961);
nor U5441 (N_5441,N_863,N_2358);
xor U5442 (N_5442,N_1027,N_982);
or U5443 (N_5443,N_2956,N_1611);
or U5444 (N_5444,N_1600,N_2487);
nand U5445 (N_5445,N_4337,N_4491);
xor U5446 (N_5446,N_409,N_498);
xor U5447 (N_5447,N_965,N_240);
nor U5448 (N_5448,N_4149,N_2544);
or U5449 (N_5449,N_236,N_2319);
or U5450 (N_5450,N_775,N_2878);
xnor U5451 (N_5451,N_4305,N_3898);
nor U5452 (N_5452,N_4553,N_732);
or U5453 (N_5453,N_3615,N_370);
nand U5454 (N_5454,N_3644,N_4874);
and U5455 (N_5455,N_2468,N_3892);
nand U5456 (N_5456,N_3097,N_2618);
nor U5457 (N_5457,N_1229,N_2533);
and U5458 (N_5458,N_2896,N_1888);
xor U5459 (N_5459,N_3754,N_4388);
nand U5460 (N_5460,N_2848,N_443);
or U5461 (N_5461,N_2869,N_3538);
or U5462 (N_5462,N_4236,N_4119);
nand U5463 (N_5463,N_1570,N_4703);
or U5464 (N_5464,N_2164,N_2105);
or U5465 (N_5465,N_3520,N_300);
or U5466 (N_5466,N_617,N_2921);
and U5467 (N_5467,N_4503,N_3271);
xor U5468 (N_5468,N_3074,N_4866);
nor U5469 (N_5469,N_3659,N_175);
or U5470 (N_5470,N_1900,N_3841);
nor U5471 (N_5471,N_2194,N_2288);
nand U5472 (N_5472,N_2428,N_4663);
or U5473 (N_5473,N_4619,N_2026);
xor U5474 (N_5474,N_1440,N_4121);
xnor U5475 (N_5475,N_3175,N_976);
xnor U5476 (N_5476,N_2044,N_1575);
nand U5477 (N_5477,N_4566,N_4434);
nor U5478 (N_5478,N_1911,N_1914);
nand U5479 (N_5479,N_4965,N_1258);
and U5480 (N_5480,N_1388,N_1806);
xnor U5481 (N_5481,N_4854,N_4536);
or U5482 (N_5482,N_1976,N_1154);
and U5483 (N_5483,N_2458,N_1147);
nand U5484 (N_5484,N_2189,N_719);
xnor U5485 (N_5485,N_935,N_540);
nand U5486 (N_5486,N_2081,N_3202);
and U5487 (N_5487,N_3783,N_3499);
or U5488 (N_5488,N_3861,N_3728);
nor U5489 (N_5489,N_1102,N_1797);
xnor U5490 (N_5490,N_4436,N_220);
or U5491 (N_5491,N_4609,N_3323);
xnor U5492 (N_5492,N_3275,N_198);
nor U5493 (N_5493,N_581,N_4033);
xnor U5494 (N_5494,N_345,N_1902);
or U5495 (N_5495,N_3434,N_1338);
xor U5496 (N_5496,N_2635,N_4067);
and U5497 (N_5497,N_4956,N_1180);
nor U5498 (N_5498,N_906,N_151);
and U5499 (N_5499,N_2264,N_3065);
nand U5500 (N_5500,N_3296,N_3386);
or U5501 (N_5501,N_948,N_3585);
nor U5502 (N_5502,N_3611,N_2259);
xor U5503 (N_5503,N_1690,N_3762);
nand U5504 (N_5504,N_2365,N_2570);
nand U5505 (N_5505,N_1389,N_203);
and U5506 (N_5506,N_4192,N_2449);
xor U5507 (N_5507,N_2100,N_578);
nand U5508 (N_5508,N_1397,N_1972);
and U5509 (N_5509,N_555,N_4245);
and U5510 (N_5510,N_2640,N_1805);
or U5511 (N_5511,N_4296,N_4078);
or U5512 (N_5512,N_4881,N_2659);
xnor U5513 (N_5513,N_4823,N_3343);
or U5514 (N_5514,N_1910,N_4325);
and U5515 (N_5515,N_2598,N_1961);
or U5516 (N_5516,N_232,N_819);
and U5517 (N_5517,N_501,N_1899);
nor U5518 (N_5518,N_942,N_4018);
nand U5519 (N_5519,N_2519,N_4068);
xor U5520 (N_5520,N_441,N_4006);
xor U5521 (N_5521,N_1306,N_1026);
nor U5522 (N_5522,N_4280,N_417);
xor U5523 (N_5523,N_1268,N_4999);
nor U5524 (N_5524,N_4211,N_2440);
xnor U5525 (N_5525,N_1684,N_3028);
and U5526 (N_5526,N_837,N_757);
nor U5527 (N_5527,N_4400,N_1406);
xnor U5528 (N_5528,N_551,N_4927);
xor U5529 (N_5529,N_4297,N_1950);
or U5530 (N_5530,N_2451,N_923);
xnor U5531 (N_5531,N_2372,N_3305);
and U5532 (N_5532,N_675,N_2491);
nor U5533 (N_5533,N_4690,N_1923);
nor U5534 (N_5534,N_284,N_3743);
or U5535 (N_5535,N_853,N_1006);
nand U5536 (N_5536,N_3536,N_4025);
nor U5537 (N_5537,N_1403,N_4334);
nand U5538 (N_5538,N_2589,N_1962);
or U5539 (N_5539,N_493,N_4693);
or U5540 (N_5540,N_342,N_3419);
nand U5541 (N_5541,N_4443,N_2706);
nor U5542 (N_5542,N_2743,N_4957);
nor U5543 (N_5543,N_22,N_1871);
xnor U5544 (N_5544,N_2527,N_1470);
and U5545 (N_5545,N_4943,N_4593);
nand U5546 (N_5546,N_2810,N_385);
nor U5547 (N_5547,N_1886,N_3547);
nand U5548 (N_5548,N_1169,N_3808);
nor U5549 (N_5549,N_1695,N_2521);
xor U5550 (N_5550,N_3180,N_2175);
nand U5551 (N_5551,N_2462,N_437);
or U5552 (N_5552,N_4293,N_3389);
and U5553 (N_5553,N_2225,N_532);
nor U5554 (N_5554,N_3681,N_1921);
and U5555 (N_5555,N_4662,N_568);
and U5556 (N_5556,N_3568,N_3349);
xnor U5557 (N_5557,N_1475,N_4262);
nor U5558 (N_5558,N_1638,N_3344);
nand U5559 (N_5559,N_3007,N_4447);
xnor U5560 (N_5560,N_1172,N_4478);
and U5561 (N_5561,N_1554,N_4729);
nor U5562 (N_5562,N_3190,N_348);
and U5563 (N_5563,N_2911,N_553);
nor U5564 (N_5564,N_1060,N_2984);
or U5565 (N_5565,N_864,N_3823);
nand U5566 (N_5566,N_1235,N_3293);
xnor U5567 (N_5567,N_1918,N_2775);
xor U5568 (N_5568,N_4811,N_62);
and U5569 (N_5569,N_1652,N_1084);
xor U5570 (N_5570,N_403,N_696);
xor U5571 (N_5571,N_791,N_3421);
or U5572 (N_5572,N_879,N_1680);
nand U5573 (N_5573,N_1025,N_316);
and U5574 (N_5574,N_4583,N_3594);
and U5575 (N_5575,N_3057,N_3652);
xnor U5576 (N_5576,N_4519,N_1350);
or U5577 (N_5577,N_1788,N_2121);
xnor U5578 (N_5578,N_4994,N_1614);
xnor U5579 (N_5579,N_1865,N_699);
and U5580 (N_5580,N_3939,N_556);
and U5581 (N_5581,N_2056,N_152);
nor U5582 (N_5582,N_4370,N_3278);
and U5583 (N_5583,N_4456,N_3088);
nor U5584 (N_5584,N_1163,N_2411);
and U5585 (N_5585,N_3699,N_2593);
nand U5586 (N_5586,N_839,N_3733);
or U5587 (N_5587,N_26,N_2424);
nor U5588 (N_5588,N_1919,N_4291);
and U5589 (N_5589,N_2126,N_3627);
nor U5590 (N_5590,N_2502,N_912);
or U5591 (N_5591,N_2154,N_1589);
or U5592 (N_5592,N_3535,N_278);
nand U5593 (N_5593,N_679,N_2813);
xnor U5594 (N_5594,N_123,N_390);
and U5595 (N_5595,N_2128,N_505);
xor U5596 (N_5596,N_1967,N_4565);
xor U5597 (N_5597,N_445,N_1384);
and U5598 (N_5598,N_4610,N_2919);
xor U5599 (N_5599,N_1282,N_2515);
nand U5600 (N_5600,N_2730,N_1426);
nor U5601 (N_5601,N_4764,N_2484);
xnor U5602 (N_5602,N_1567,N_2671);
xnor U5603 (N_5603,N_2590,N_2082);
xnor U5604 (N_5604,N_1057,N_3076);
xor U5605 (N_5605,N_2955,N_1474);
nand U5606 (N_5606,N_880,N_1429);
nand U5607 (N_5607,N_686,N_4828);
nor U5608 (N_5608,N_1641,N_2926);
or U5609 (N_5609,N_1096,N_4249);
xnor U5610 (N_5610,N_3069,N_1887);
nand U5611 (N_5611,N_633,N_620);
nor U5612 (N_5612,N_1867,N_119);
or U5613 (N_5613,N_711,N_4715);
nor U5614 (N_5614,N_2815,N_4784);
nor U5615 (N_5615,N_4128,N_3081);
nand U5616 (N_5616,N_3203,N_4959);
nor U5617 (N_5617,N_2307,N_854);
nand U5618 (N_5618,N_1142,N_2890);
nand U5619 (N_5619,N_3735,N_1218);
nand U5620 (N_5620,N_3529,N_302);
xor U5621 (N_5621,N_660,N_2573);
and U5622 (N_5622,N_3816,N_31);
xnor U5623 (N_5623,N_4837,N_1398);
and U5624 (N_5624,N_973,N_2840);
or U5625 (N_5625,N_3867,N_4403);
nand U5626 (N_5626,N_3058,N_4473);
and U5627 (N_5627,N_3215,N_4422);
and U5628 (N_5628,N_3213,N_3301);
xnor U5629 (N_5629,N_3641,N_242);
or U5630 (N_5630,N_3391,N_1178);
xnor U5631 (N_5631,N_3186,N_2771);
nand U5632 (N_5632,N_209,N_869);
and U5633 (N_5633,N_3334,N_3932);
xnor U5634 (N_5634,N_2159,N_4366);
nor U5635 (N_5635,N_1613,N_4584);
xor U5636 (N_5636,N_2847,N_1993);
nor U5637 (N_5637,N_4901,N_1631);
or U5638 (N_5638,N_1843,N_1861);
nand U5639 (N_5639,N_2673,N_3549);
and U5640 (N_5640,N_2877,N_3657);
xnor U5641 (N_5641,N_3325,N_141);
nor U5642 (N_5642,N_3162,N_3191);
xor U5643 (N_5643,N_1290,N_1928);
nand U5644 (N_5644,N_2953,N_3406);
and U5645 (N_5645,N_665,N_1518);
nand U5646 (N_5646,N_3246,N_2923);
nand U5647 (N_5647,N_4064,N_4003);
nor U5648 (N_5648,N_4358,N_2986);
nand U5649 (N_5649,N_226,N_187);
nor U5650 (N_5650,N_3662,N_972);
and U5651 (N_5651,N_862,N_914);
and U5652 (N_5652,N_3562,N_3546);
nand U5653 (N_5653,N_4282,N_2088);
xnor U5654 (N_5654,N_2935,N_2400);
nor U5655 (N_5655,N_1755,N_2494);
or U5656 (N_5656,N_2733,N_2039);
nand U5657 (N_5657,N_4146,N_4523);
and U5658 (N_5658,N_4953,N_2609);
nand U5659 (N_5659,N_3502,N_2379);
nor U5660 (N_5660,N_4980,N_4712);
or U5661 (N_5661,N_4086,N_3008);
nand U5662 (N_5662,N_2276,N_4020);
or U5663 (N_5663,N_4215,N_2133);
xor U5664 (N_5664,N_890,N_4951);
or U5665 (N_5665,N_3713,N_4702);
nor U5666 (N_5666,N_4425,N_1205);
and U5667 (N_5667,N_1625,N_1042);
nand U5668 (N_5668,N_2602,N_1825);
nand U5669 (N_5669,N_3756,N_3253);
xor U5670 (N_5670,N_850,N_1726);
or U5671 (N_5671,N_1044,N_644);
and U5672 (N_5672,N_4380,N_526);
nand U5673 (N_5673,N_1453,N_4087);
or U5674 (N_5674,N_3601,N_2650);
and U5675 (N_5675,N_4103,N_3116);
nor U5676 (N_5676,N_1759,N_4462);
nor U5677 (N_5677,N_2929,N_4819);
xor U5678 (N_5678,N_1455,N_2835);
nor U5679 (N_5679,N_3239,N_884);
or U5680 (N_5680,N_2973,N_3115);
or U5681 (N_5681,N_697,N_2579);
and U5682 (N_5682,N_500,N_824);
xor U5683 (N_5683,N_1713,N_1210);
nor U5684 (N_5684,N_2645,N_547);
or U5685 (N_5685,N_3876,N_797);
nor U5686 (N_5686,N_173,N_4104);
or U5687 (N_5687,N_861,N_1011);
or U5688 (N_5688,N_4361,N_3672);
or U5689 (N_5689,N_311,N_3061);
and U5690 (N_5690,N_3612,N_1283);
nand U5691 (N_5691,N_4454,N_2912);
nand U5692 (N_5692,N_833,N_4756);
and U5693 (N_5693,N_2363,N_2745);
or U5694 (N_5694,N_3786,N_341);
nand U5695 (N_5695,N_3139,N_2330);
xor U5696 (N_5696,N_4123,N_2215);
xnor U5697 (N_5697,N_1893,N_2066);
nor U5698 (N_5698,N_3998,N_1002);
nand U5699 (N_5699,N_74,N_4316);
and U5700 (N_5700,N_2554,N_957);
nor U5701 (N_5701,N_1874,N_3281);
nor U5702 (N_5702,N_4004,N_3003);
and U5703 (N_5703,N_3565,N_606);
xnor U5704 (N_5704,N_4964,N_1486);
nand U5705 (N_5705,N_897,N_3571);
or U5706 (N_5706,N_2016,N_10);
nor U5707 (N_5707,N_4842,N_4080);
nand U5708 (N_5708,N_3774,N_4060);
and U5709 (N_5709,N_3686,N_2642);
and U5710 (N_5710,N_3128,N_2270);
nor U5711 (N_5711,N_2261,N_1226);
and U5712 (N_5712,N_3481,N_4470);
or U5713 (N_5713,N_4231,N_3723);
or U5714 (N_5714,N_1895,N_89);
nand U5715 (N_5715,N_1757,N_34);
and U5716 (N_5716,N_2648,N_1171);
xnor U5717 (N_5717,N_3030,N_703);
and U5718 (N_5718,N_2073,N_2897);
xor U5719 (N_5719,N_2687,N_666);
xor U5720 (N_5720,N_1566,N_132);
nand U5721 (N_5721,N_306,N_4998);
nor U5722 (N_5722,N_1994,N_1988);
nor U5723 (N_5723,N_1487,N_759);
and U5724 (N_5724,N_2209,N_613);
and U5725 (N_5725,N_354,N_3212);
and U5726 (N_5726,N_4709,N_4035);
nor U5727 (N_5727,N_2063,N_4939);
or U5728 (N_5728,N_4392,N_4813);
nor U5729 (N_5729,N_4739,N_2171);
or U5730 (N_5730,N_1982,N_765);
nor U5731 (N_5731,N_1547,N_4726);
or U5732 (N_5732,N_4921,N_1124);
and U5733 (N_5733,N_1309,N_41);
xnor U5734 (N_5734,N_667,N_3902);
or U5735 (N_5735,N_2183,N_657);
xnor U5736 (N_5736,N_4931,N_2397);
nor U5737 (N_5737,N_3132,N_87);
nor U5738 (N_5738,N_1182,N_2580);
nand U5739 (N_5739,N_276,N_812);
and U5740 (N_5740,N_388,N_4551);
or U5741 (N_5741,N_4155,N_2507);
nor U5742 (N_5742,N_1651,N_2177);
xor U5743 (N_5743,N_4831,N_3732);
xnor U5744 (N_5744,N_3716,N_1946);
xor U5745 (N_5745,N_4152,N_1192);
and U5746 (N_5746,N_4879,N_4107);
and U5747 (N_5747,N_1984,N_1348);
and U5748 (N_5748,N_1752,N_1234);
xor U5749 (N_5749,N_3111,N_3815);
and U5750 (N_5750,N_491,N_4453);
xnor U5751 (N_5751,N_4605,N_2042);
and U5752 (N_5752,N_3906,N_1945);
nand U5753 (N_5753,N_3807,N_1947);
nor U5754 (N_5754,N_4142,N_2158);
and U5755 (N_5755,N_3035,N_4411);
nand U5756 (N_5756,N_4606,N_3412);
nor U5757 (N_5757,N_3238,N_4591);
nor U5758 (N_5758,N_3223,N_508);
and U5759 (N_5759,N_427,N_1627);
and U5760 (N_5760,N_4012,N_511);
nand U5761 (N_5761,N_1802,N_4016);
xnor U5762 (N_5762,N_4063,N_2790);
nor U5763 (N_5763,N_868,N_4213);
xnor U5764 (N_5764,N_1443,N_4292);
or U5765 (N_5765,N_1699,N_513);
xnor U5766 (N_5766,N_120,N_4164);
and U5767 (N_5767,N_3482,N_4386);
nor U5768 (N_5768,N_2778,N_3324);
or U5769 (N_5769,N_3694,N_1981);
nor U5770 (N_5770,N_88,N_1370);
xnor U5771 (N_5771,N_221,N_4742);
and U5772 (N_5772,N_565,N_4946);
nand U5773 (N_5773,N_3015,N_2198);
and U5774 (N_5774,N_701,N_908);
nand U5775 (N_5775,N_522,N_2717);
nand U5776 (N_5776,N_2550,N_2753);
or U5777 (N_5777,N_4723,N_4065);
nand U5778 (N_5778,N_2568,N_1481);
nand U5779 (N_5779,N_2350,N_3040);
and U5780 (N_5780,N_33,N_4114);
and U5781 (N_5781,N_2539,N_3842);
and U5782 (N_5782,N_1905,N_1176);
and U5783 (N_5783,N_228,N_3108);
and U5784 (N_5784,N_4986,N_2384);
and U5785 (N_5785,N_1796,N_4441);
or U5786 (N_5786,N_3625,N_1371);
and U5787 (N_5787,N_3577,N_3172);
or U5788 (N_5788,N_23,N_3790);
nor U5789 (N_5789,N_1844,N_3685);
and U5790 (N_5790,N_2439,N_3054);
nor U5791 (N_5791,N_65,N_4011);
nand U5792 (N_5792,N_3257,N_574);
or U5793 (N_5793,N_2844,N_4685);
nand U5794 (N_5794,N_481,N_2280);
nand U5795 (N_5795,N_79,N_1243);
or U5796 (N_5796,N_3060,N_3945);
xor U5797 (N_5797,N_2638,N_2236);
nand U5798 (N_5798,N_2287,N_4672);
or U5799 (N_5799,N_1820,N_4423);
nor U5800 (N_5800,N_2310,N_48);
nor U5801 (N_5801,N_72,N_1112);
nor U5802 (N_5802,N_1107,N_4504);
nor U5803 (N_5803,N_4545,N_2989);
nand U5804 (N_5804,N_3026,N_4840);
and U5805 (N_5805,N_3233,N_3978);
nand U5806 (N_5806,N_4629,N_1221);
nand U5807 (N_5807,N_1512,N_1675);
nor U5808 (N_5808,N_4147,N_1639);
nor U5809 (N_5809,N_3541,N_3403);
or U5810 (N_5810,N_4925,N_706);
xnor U5811 (N_5811,N_807,N_1092);
or U5812 (N_5812,N_2265,N_3784);
and U5813 (N_5813,N_2431,N_2945);
or U5814 (N_5814,N_492,N_3781);
and U5815 (N_5815,N_2037,N_698);
nand U5816 (N_5816,N_2541,N_3574);
nor U5817 (N_5817,N_104,N_1118);
or U5818 (N_5818,N_4960,N_4559);
xnor U5819 (N_5819,N_2738,N_2759);
and U5820 (N_5820,N_258,N_3113);
or U5821 (N_5821,N_358,N_959);
xor U5822 (N_5822,N_4981,N_4328);
or U5823 (N_5823,N_577,N_4170);
and U5824 (N_5824,N_3674,N_3745);
xnor U5825 (N_5825,N_1458,N_1766);
nor U5826 (N_5826,N_2153,N_539);
nand U5827 (N_5827,N_1996,N_1841);
nand U5828 (N_5828,N_2705,N_3197);
or U5829 (N_5829,N_1404,N_3360);
and U5830 (N_5830,N_3290,N_5);
and U5831 (N_5831,N_3874,N_3647);
nor U5832 (N_5832,N_1618,N_3853);
and U5833 (N_5833,N_2135,N_406);
nor U5834 (N_5834,N_3286,N_4181);
nor U5835 (N_5835,N_2496,N_4776);
nor U5836 (N_5836,N_1187,N_1637);
or U5837 (N_5837,N_2070,N_1692);
or U5838 (N_5838,N_688,N_762);
and U5839 (N_5839,N_3241,N_4429);
or U5840 (N_5840,N_4847,N_299);
and U5841 (N_5841,N_4658,N_2707);
or U5842 (N_5842,N_2746,N_580);
nor U5843 (N_5843,N_4611,N_1289);
and U5844 (N_5844,N_1756,N_3056);
nor U5845 (N_5845,N_3828,N_4390);
nand U5846 (N_5846,N_3234,N_939);
nor U5847 (N_5847,N_2481,N_1241);
and U5848 (N_5848,N_3326,N_1240);
nand U5849 (N_5849,N_3506,N_2740);
nor U5850 (N_5850,N_2273,N_1593);
xnor U5851 (N_5851,N_3877,N_4552);
and U5852 (N_5852,N_2678,N_2047);
xnor U5853 (N_5853,N_2344,N_4749);
or U5854 (N_5854,N_3452,N_3691);
or U5855 (N_5855,N_1500,N_2838);
xor U5856 (N_5856,N_4000,N_2131);
or U5857 (N_5857,N_4800,N_561);
nand U5858 (N_5858,N_4094,N_2898);
nor U5859 (N_5859,N_4350,N_571);
and U5860 (N_5860,N_1227,N_700);
and U5861 (N_5861,N_4289,N_1543);
nor U5862 (N_5862,N_3188,N_2581);
or U5863 (N_5863,N_693,N_4010);
or U5864 (N_5864,N_149,N_4525);
or U5865 (N_5865,N_2059,N_2629);
nand U5866 (N_5866,N_111,N_1727);
nor U5867 (N_5867,N_4092,N_1421);
nor U5868 (N_5868,N_2483,N_2751);
nor U5869 (N_5869,N_1295,N_2663);
or U5870 (N_5870,N_408,N_71);
or U5871 (N_5871,N_2292,N_1767);
nor U5872 (N_5872,N_796,N_2240);
nand U5873 (N_5873,N_3396,N_2316);
and U5874 (N_5874,N_887,N_2587);
xnor U5875 (N_5875,N_1552,N_1108);
xnor U5876 (N_5876,N_3917,N_4627);
or U5877 (N_5877,N_4737,N_438);
nand U5878 (N_5878,N_4969,N_3299);
nor U5879 (N_5879,N_1372,N_2737);
and U5880 (N_5880,N_361,N_4134);
and U5881 (N_5881,N_3442,N_114);
and U5882 (N_5882,N_2291,N_1049);
nor U5883 (N_5883,N_2633,N_167);
or U5884 (N_5884,N_1542,N_2862);
and U5885 (N_5885,N_502,N_4714);
xor U5886 (N_5886,N_4767,N_1311);
nor U5887 (N_5887,N_105,N_3543);
nor U5888 (N_5888,N_3505,N_4055);
nand U5889 (N_5889,N_2020,N_3595);
nand U5890 (N_5890,N_1669,N_1432);
nand U5891 (N_5891,N_4995,N_4790);
xnor U5892 (N_5892,N_46,N_1008);
or U5893 (N_5893,N_4585,N_3631);
nor U5894 (N_5894,N_2366,N_486);
xor U5895 (N_5895,N_920,N_2939);
or U5896 (N_5896,N_597,N_1045);
xor U5897 (N_5897,N_3804,N_1657);
or U5898 (N_5898,N_2404,N_787);
xor U5899 (N_5899,N_1392,N_4736);
and U5900 (N_5900,N_3578,N_471);
nand U5901 (N_5901,N_3351,N_3071);
xnor U5902 (N_5902,N_1778,N_3776);
or U5903 (N_5903,N_3133,N_1408);
xor U5904 (N_5904,N_249,N_4577);
or U5905 (N_5905,N_2511,N_3182);
xor U5906 (N_5906,N_1364,N_2604);
and U5907 (N_5907,N_4832,N_4618);
and U5908 (N_5908,N_3830,N_61);
and U5909 (N_5909,N_621,N_1095);
nor U5910 (N_5910,N_2023,N_335);
nand U5911 (N_5911,N_3025,N_4974);
nand U5912 (N_5912,N_4747,N_4450);
and U5913 (N_5913,N_424,N_1194);
nand U5914 (N_5914,N_1813,N_3765);
and U5915 (N_5915,N_1034,N_846);
and U5916 (N_5916,N_2712,N_4047);
and U5917 (N_5917,N_3067,N_946);
and U5918 (N_5918,N_2178,N_3375);
nor U5919 (N_5919,N_4598,N_4017);
and U5920 (N_5920,N_2982,N_2529);
nor U5921 (N_5921,N_1314,N_3670);
nand U5922 (N_5922,N_190,N_4219);
nand U5923 (N_5923,N_2997,N_754);
nor U5924 (N_5924,N_155,N_4725);
nor U5925 (N_5925,N_3983,N_2176);
xor U5926 (N_5926,N_1671,N_2643);
nand U5927 (N_5927,N_2892,N_1396);
and U5928 (N_5928,N_1866,N_3742);
and U5929 (N_5929,N_3272,N_2180);
xor U5930 (N_5930,N_1254,N_2090);
xor U5931 (N_5931,N_678,N_1296);
nor U5932 (N_5932,N_591,N_3219);
nor U5933 (N_5933,N_68,N_237);
nor U5934 (N_5934,N_2278,N_4415);
nor U5935 (N_5935,N_1452,N_2254);
and U5936 (N_5936,N_99,N_2651);
or U5937 (N_5937,N_1202,N_1413);
xor U5938 (N_5938,N_2263,N_2118);
xor U5939 (N_5939,N_3302,N_346);
xor U5940 (N_5940,N_4641,N_4216);
or U5941 (N_5941,N_3193,N_1361);
or U5942 (N_5942,N_418,N_3398);
nor U5943 (N_5943,N_1269,N_3785);
nand U5944 (N_5944,N_1020,N_4332);
nand U5945 (N_5945,N_2041,N_2050);
nor U5946 (N_5946,N_4428,N_2169);
xnor U5947 (N_5947,N_2714,N_4760);
and U5948 (N_5948,N_528,N_3771);
and U5949 (N_5949,N_2583,N_3582);
nor U5950 (N_5950,N_2968,N_1508);
xnor U5951 (N_5951,N_3201,N_3780);
nand U5952 (N_5952,N_4522,N_169);
nor U5953 (N_5953,N_2396,N_3313);
nor U5954 (N_5954,N_447,N_1944);
or U5955 (N_5955,N_4895,N_2891);
nor U5956 (N_5956,N_4505,N_3295);
nor U5957 (N_5957,N_4378,N_4630);
xnor U5958 (N_5958,N_1369,N_2141);
and U5959 (N_5959,N_425,N_2446);
nand U5960 (N_5960,N_2895,N_4793);
nand U5961 (N_5961,N_1339,N_325);
nor U5962 (N_5962,N_685,N_4501);
and U5963 (N_5963,N_12,N_4458);
or U5964 (N_5964,N_1039,N_2235);
nor U5965 (N_5965,N_2454,N_4656);
and U5966 (N_5966,N_2668,N_4982);
xor U5967 (N_5967,N_1644,N_4402);
xnor U5968 (N_5968,N_3039,N_1679);
and U5969 (N_5969,N_142,N_3082);
xnor U5970 (N_5970,N_3620,N_4963);
and U5971 (N_5971,N_3049,N_4200);
nand U5972 (N_5972,N_42,N_4302);
nand U5973 (N_5973,N_2342,N_2452);
nand U5974 (N_5974,N_3251,N_1828);
xor U5975 (N_5975,N_4771,N_1924);
and U5976 (N_5976,N_4886,N_4367);
nor U5977 (N_5977,N_814,N_1630);
and U5978 (N_5978,N_4528,N_2108);
or U5979 (N_5979,N_4990,N_2480);
nand U5980 (N_5980,N_1196,N_389);
xnor U5981 (N_5981,N_1353,N_2018);
or U5982 (N_5982,N_2765,N_2313);
nand U5983 (N_5983,N_4394,N_4124);
and U5984 (N_5984,N_1351,N_1315);
nor U5985 (N_5985,N_4126,N_2497);
or U5986 (N_5986,N_1368,N_3047);
nand U5987 (N_5987,N_608,N_4844);
nand U5988 (N_5988,N_4387,N_3464);
xor U5989 (N_5989,N_4440,N_1851);
or U5990 (N_5990,N_739,N_2661);
nand U5991 (N_5991,N_1246,N_3176);
nor U5992 (N_5992,N_1230,N_1395);
xor U5993 (N_5993,N_1842,N_2102);
nor U5994 (N_5994,N_2656,N_670);
or U5995 (N_5995,N_4716,N_1024);
or U5996 (N_5996,N_3121,N_1208);
and U5997 (N_5997,N_2908,N_2691);
nand U5998 (N_5998,N_4782,N_1181);
nor U5999 (N_5999,N_2069,N_3575);
nand U6000 (N_6000,N_586,N_293);
nor U6001 (N_6001,N_1478,N_4122);
nand U6002 (N_6002,N_1150,N_847);
nor U6003 (N_6003,N_2739,N_3888);
nor U6004 (N_6004,N_2060,N_4158);
xor U6005 (N_6005,N_4717,N_320);
nor U6006 (N_6006,N_1894,N_2328);
nor U6007 (N_6007,N_1327,N_2470);
nand U6008 (N_6008,N_4984,N_4547);
xor U6009 (N_6009,N_4088,N_554);
nand U6010 (N_6010,N_3171,N_2628);
xor U6011 (N_6011,N_4616,N_2907);
xor U6012 (N_6012,N_1058,N_4581);
and U6013 (N_6013,N_4664,N_4809);
nand U6014 (N_6014,N_2245,N_3232);
nor U6015 (N_6015,N_1715,N_2137);
xor U6016 (N_6016,N_4592,N_2012);
and U6017 (N_6017,N_338,N_4765);
nor U6018 (N_6018,N_4838,N_3514);
nor U6019 (N_6019,N_1116,N_898);
and U6020 (N_6020,N_2623,N_4757);
or U6021 (N_6021,N_3532,N_3552);
nor U6022 (N_6022,N_3210,N_2964);
xnor U6023 (N_6023,N_440,N_1822);
nand U6024 (N_6024,N_2781,N_3143);
nand U6025 (N_6025,N_1634,N_1706);
nand U6026 (N_6026,N_37,N_2808);
nor U6027 (N_6027,N_3320,N_1819);
and U6028 (N_6028,N_2680,N_802);
xnor U6029 (N_6029,N_3667,N_2444);
nand U6030 (N_6030,N_246,N_1152);
nand U6031 (N_6031,N_525,N_4368);
nand U6032 (N_6032,N_3207,N_768);
or U6033 (N_6033,N_3474,N_3772);
or U6034 (N_6034,N_2253,N_4558);
or U6035 (N_6035,N_4039,N_223);
xor U6036 (N_6036,N_3554,N_2791);
nand U6037 (N_6037,N_2545,N_4516);
nor U6038 (N_6038,N_1782,N_3327);
xor U6039 (N_6039,N_3357,N_1043);
nor U6040 (N_6040,N_4557,N_2359);
nand U6041 (N_6041,N_2297,N_3235);
and U6042 (N_6042,N_4193,N_383);
or U6043 (N_6043,N_4333,N_4562);
nand U6044 (N_6044,N_3555,N_3024);
or U6045 (N_6045,N_49,N_2315);
nor U6046 (N_6046,N_3806,N_4267);
xnor U6047 (N_6047,N_4962,N_3589);
xor U6048 (N_6048,N_4182,N_3797);
nor U6049 (N_6049,N_3160,N_3092);
xor U6050 (N_6050,N_2200,N_1873);
and U6051 (N_6051,N_2686,N_4225);
nand U6052 (N_6052,N_585,N_907);
xnor U6053 (N_6053,N_766,N_4253);
nor U6054 (N_6054,N_146,N_490);
nand U6055 (N_6055,N_2710,N_102);
nor U6056 (N_6056,N_3992,N_1159);
nand U6057 (N_6057,N_1483,N_970);
xnor U6058 (N_6058,N_2399,N_434);
or U6059 (N_6059,N_30,N_2234);
or U6060 (N_6060,N_2378,N_4391);
xor U6061 (N_6061,N_694,N_4829);
and U6062 (N_6062,N_3401,N_4497);
and U6063 (N_6063,N_930,N_2450);
xnor U6064 (N_6064,N_4897,N_1729);
or U6065 (N_6065,N_2139,N_2535);
xnor U6066 (N_6066,N_4512,N_1880);
nand U6067 (N_6067,N_2657,N_3851);
nand U6068 (N_6068,N_2486,N_1550);
xnor U6069 (N_6069,N_4587,N_3504);
nand U6070 (N_6070,N_1667,N_4132);
and U6071 (N_6071,N_4090,N_283);
xor U6072 (N_6072,N_2772,N_535);
nor U6073 (N_6073,N_4071,N_2901);
nor U6074 (N_6074,N_4084,N_3448);
or U6075 (N_6075,N_3004,N_321);
or U6076 (N_6076,N_3800,N_3700);
nor U6077 (N_6077,N_2927,N_984);
and U6078 (N_6078,N_1410,N_885);
and U6079 (N_6079,N_2111,N_2876);
nor U6080 (N_6080,N_3628,N_1320);
nand U6081 (N_6081,N_81,N_1594);
or U6082 (N_6082,N_2242,N_4331);
nor U6083 (N_6083,N_4191,N_331);
nand U6084 (N_6084,N_2728,N_4997);
and U6085 (N_6085,N_4533,N_2290);
or U6086 (N_6086,N_3909,N_1362);
nor U6087 (N_6087,N_3824,N_4384);
or U6088 (N_6088,N_2516,N_1836);
xnor U6089 (N_6089,N_4204,N_3791);
xor U6090 (N_6090,N_2501,N_211);
nand U6091 (N_6091,N_4683,N_2116);
nand U6092 (N_6092,N_3072,N_729);
nand U6093 (N_6093,N_435,N_1469);
and U6094 (N_6094,N_2068,N_997);
nand U6095 (N_6095,N_4203,N_992);
nand U6096 (N_6096,N_916,N_1374);
nor U6097 (N_6097,N_2836,N_1553);
and U6098 (N_6098,N_645,N_4850);
nand U6099 (N_6099,N_3022,N_3976);
or U6100 (N_6100,N_2767,N_245);
or U6101 (N_6101,N_1754,N_2809);
nor U6102 (N_6102,N_659,N_4875);
nand U6103 (N_6103,N_3766,N_612);
or U6104 (N_6104,N_2303,N_1330);
nand U6105 (N_6105,N_3399,N_1003);
xor U6106 (N_6106,N_4668,N_277);
and U6107 (N_6107,N_2495,N_3110);
nand U6108 (N_6108,N_4554,N_1889);
nor U6109 (N_6109,N_2660,N_485);
or U6110 (N_6110,N_4418,N_3285);
nand U6111 (N_6111,N_2548,N_4301);
or U6112 (N_6112,N_836,N_92);
and U6113 (N_6113,N_3624,N_4758);
xor U6114 (N_6114,N_3985,N_3599);
nand U6115 (N_6115,N_1139,N_3884);
and U6116 (N_6116,N_2392,N_1188);
or U6117 (N_6117,N_704,N_3720);
nor U6118 (N_6118,N_457,N_2205);
or U6119 (N_6119,N_2248,N_741);
nor U6120 (N_6120,N_317,N_4311);
or U6121 (N_6121,N_436,N_1038);
nand U6122 (N_6122,N_3404,N_3340);
or U6123 (N_6123,N_3510,N_3101);
nand U6124 (N_6124,N_451,N_2277);
and U6125 (N_6125,N_298,N_134);
and U6126 (N_6126,N_4369,N_4348);
xor U6127 (N_6127,N_4883,N_4856);
and U6128 (N_6128,N_3997,N_4966);
nand U6129 (N_6129,N_4007,N_4858);
xnor U6130 (N_6130,N_2162,N_295);
nor U6131 (N_6131,N_2619,N_2842);
or U6132 (N_6132,N_2109,N_3576);
xnor U6133 (N_6133,N_2725,N_3579);
and U6134 (N_6134,N_3527,N_799);
and U6135 (N_6135,N_2038,N_251);
nand U6136 (N_6136,N_2262,N_605);
xor U6137 (N_6137,N_3354,N_3885);
nand U6138 (N_6138,N_2314,N_3690);
and U6139 (N_6139,N_3064,N_1365);
nand U6140 (N_6140,N_4973,N_994);
or U6141 (N_6141,N_623,N_2250);
or U6142 (N_6142,N_1405,N_309);
and U6143 (N_6143,N_3676,N_1207);
nor U6144 (N_6144,N_1435,N_3138);
and U6145 (N_6145,N_1581,N_1373);
and U6146 (N_6146,N_2127,N_1587);
nand U6147 (N_6147,N_1821,N_1402);
nor U6148 (N_6148,N_720,N_78);
nand U6149 (N_6149,N_960,N_135);
xnor U6150 (N_6150,N_4070,N_2009);
xnor U6151 (N_6151,N_3509,N_549);
or U6152 (N_6152,N_4855,N_3857);
xnor U6153 (N_6153,N_654,N_1253);
nor U6154 (N_6154,N_3031,N_4076);
and U6155 (N_6155,N_4041,N_2679);
nand U6156 (N_6156,N_3294,N_2900);
xnor U6157 (N_6157,N_1017,N_4416);
or U6158 (N_6158,N_2922,N_1779);
and U6159 (N_6159,N_4839,N_347);
nor U6160 (N_6160,N_2348,N_2577);
nand U6161 (N_6161,N_1280,N_2410);
xor U6162 (N_6162,N_3960,N_4677);
and U6163 (N_6163,N_1804,N_18);
nor U6164 (N_6164,N_482,N_3592);
or U6165 (N_6165,N_3169,N_1658);
or U6166 (N_6166,N_714,N_467);
nor U6167 (N_6167,N_4272,N_3962);
xor U6168 (N_6168,N_1739,N_2202);
xnor U6169 (N_6169,N_738,N_809);
xor U6170 (N_6170,N_3435,N_444);
xnor U6171 (N_6171,N_263,N_4141);
nand U6172 (N_6172,N_904,N_3050);
xnor U6173 (N_6173,N_4360,N_2354);
xnor U6174 (N_6174,N_4194,N_1582);
nor U6175 (N_6175,N_90,N_7);
xnor U6176 (N_6176,N_1838,N_459);
nor U6177 (N_6177,N_3558,N_1162);
and U6178 (N_6178,N_4991,N_3358);
and U6179 (N_6179,N_2676,N_4346);
nor U6180 (N_6180,N_1609,N_1717);
nor U6181 (N_6181,N_2812,N_3942);
or U6182 (N_6182,N_1427,N_115);
xnor U6183 (N_6183,N_3288,N_3303);
nor U6184 (N_6184,N_1760,N_2803);
or U6185 (N_6185,N_366,N_1155);
and U6186 (N_6186,N_2443,N_3661);
nor U6187 (N_6187,N_3134,N_3353);
or U6188 (N_6188,N_4455,N_3680);
and U6189 (N_6189,N_1698,N_913);
nor U6190 (N_6190,N_2625,N_1425);
xor U6191 (N_6191,N_2724,N_1573);
or U6192 (N_6192,N_2586,N_1514);
nand U6193 (N_6193,N_1131,N_783);
xor U6194 (N_6194,N_1109,N_2281);
or U6195 (N_6195,N_108,N_3001);
and U6196 (N_6196,N_225,N_1411);
nor U6197 (N_6197,N_2394,N_4534);
nor U6198 (N_6198,N_2722,N_234);
xor U6199 (N_6199,N_3854,N_1479);
and U6200 (N_6200,N_1533,N_421);
nand U6201 (N_6201,N_4139,N_3141);
or U6202 (N_6202,N_800,N_1212);
nand U6203 (N_6203,N_2785,N_4487);
nand U6204 (N_6204,N_446,N_1855);
or U6205 (N_6205,N_806,N_642);
nor U6206 (N_6206,N_3878,N_2405);
or U6207 (N_6207,N_4640,N_3944);
nor U6208 (N_6208,N_995,N_2996);
and U6209 (N_6209,N_1583,N_1001);
nor U6210 (N_6210,N_2260,N_4992);
nor U6211 (N_6211,N_3542,N_3086);
or U6212 (N_6212,N_2030,N_2447);
and U6213 (N_6213,N_253,N_1328);
nand U6214 (N_6214,N_1897,N_4218);
and U6215 (N_6215,N_1536,N_4317);
nand U6216 (N_6216,N_1793,N_1837);
and U6217 (N_6217,N_1785,N_63);
or U6218 (N_6218,N_1366,N_3912);
xnor U6219 (N_6219,N_244,N_1869);
nor U6220 (N_6220,N_3466,N_3282);
or U6221 (N_6221,N_4696,N_3423);
xnor U6222 (N_6222,N_1561,N_4273);
xnor U6223 (N_6223,N_3161,N_405);
nand U6224 (N_6224,N_2985,N_3987);
nand U6225 (N_6225,N_958,N_1029);
and U6226 (N_6226,N_3463,N_3964);
nand U6227 (N_6227,N_3168,N_4822);
nand U6228 (N_6228,N_1061,N_1731);
nand U6229 (N_6229,N_2430,N_2599);
or U6230 (N_6230,N_1647,N_1882);
nor U6231 (N_6231,N_1891,N_4799);
and U6232 (N_6232,N_662,N_96);
nand U6233 (N_6233,N_1286,N_255);
and U6234 (N_6234,N_2403,N_3331);
and U6235 (N_6235,N_1491,N_903);
xor U6236 (N_6236,N_3581,N_1904);
nor U6237 (N_6237,N_4631,N_827);
and U6238 (N_6238,N_2099,N_1450);
xor U6239 (N_6239,N_2092,N_1559);
xnor U6240 (N_6240,N_2459,N_1456);
nand U6241 (N_6241,N_4270,N_404);
or U6242 (N_6242,N_3236,N_1473);
nand U6243 (N_6243,N_3714,N_1777);
nand U6244 (N_6244,N_3475,N_1065);
nand U6245 (N_6245,N_3683,N_3451);
xnor U6246 (N_6246,N_2048,N_11);
nor U6247 (N_6247,N_256,N_180);
nand U6248 (N_6248,N_3140,N_1375);
or U6249 (N_6249,N_1,N_1346);
nand U6250 (N_6250,N_2071,N_2085);
nand U6251 (N_6251,N_2616,N_3276);
nand U6252 (N_6252,N_4061,N_2562);
xor U6253 (N_6253,N_4009,N_4563);
and U6254 (N_6254,N_197,N_2760);
nor U6255 (N_6255,N_4941,N_1870);
nor U6256 (N_6256,N_782,N_1929);
nor U6257 (N_6257,N_531,N_2123);
nand U6258 (N_6258,N_2229,N_4351);
or U6259 (N_6259,N_3229,N_767);
and U6260 (N_6260,N_1263,N_4196);
nor U6261 (N_6261,N_3927,N_2448);
nor U6262 (N_6262,N_1934,N_3989);
or U6263 (N_6263,N_4621,N_3184);
nand U6264 (N_6264,N_4794,N_637);
and U6265 (N_6265,N_3027,N_1540);
nand U6266 (N_6266,N_439,N_726);
and U6267 (N_6267,N_3560,N_3621);
nand U6268 (N_6268,N_4574,N_4468);
xor U6269 (N_6269,N_50,N_4648);
xnor U6270 (N_6270,N_804,N_415);
or U6271 (N_6271,N_4449,N_2195);
nand U6272 (N_6272,N_158,N_1056);
and U6273 (N_6273,N_3919,N_4183);
or U6274 (N_6274,N_1898,N_2193);
nor U6275 (N_6275,N_465,N_506);
nand U6276 (N_6276,N_2517,N_3157);
nand U6277 (N_6277,N_988,N_2741);
nand U6278 (N_6278,N_1670,N_2148);
or U6279 (N_6279,N_499,N_2309);
nor U6280 (N_6280,N_257,N_1461);
nor U6281 (N_6281,N_2382,N_1545);
nand U6282 (N_6282,N_2325,N_687);
and U6283 (N_6283,N_601,N_2124);
nand U6284 (N_6284,N_4722,N_103);
xor U6285 (N_6285,N_3010,N_1228);
nor U6286 (N_6286,N_3865,N_2493);
nor U6287 (N_6287,N_4830,N_3521);
nand U6288 (N_6288,N_290,N_4546);
and U6289 (N_6289,N_1659,N_822);
nor U6290 (N_6290,N_206,N_3252);
and U6291 (N_6291,N_3385,N_3453);
or U6292 (N_6292,N_3920,N_3177);
nor U6293 (N_6293,N_369,N_3258);
and U6294 (N_6294,N_2928,N_4812);
xor U6295 (N_6295,N_2708,N_1685);
and U6296 (N_6296,N_4851,N_3684);
xor U6297 (N_6297,N_2763,N_4102);
nor U6298 (N_6298,N_3345,N_407);
xor U6299 (N_6299,N_758,N_1484);
nor U6300 (N_6300,N_1160,N_4603);
nor U6301 (N_6301,N_4177,N_1642);
nor U6302 (N_6302,N_3486,N_977);
xnor U6303 (N_6303,N_4156,N_2818);
and U6304 (N_6304,N_2571,N_3933);
xnor U6305 (N_6305,N_3291,N_4356);
xor U6306 (N_6306,N_1798,N_4330);
or U6307 (N_6307,N_4259,N_3687);
and U6308 (N_6308,N_4327,N_3038);
nor U6309 (N_6309,N_4923,N_893);
or U6310 (N_6310,N_728,N_4451);
xor U6311 (N_6311,N_4201,N_2311);
nor U6312 (N_6312,N_2563,N_2944);
and U6313 (N_6313,N_2821,N_3070);
nor U6314 (N_6314,N_2834,N_634);
and U6315 (N_6315,N_4412,N_1546);
and U6316 (N_6316,N_4779,N_4579);
or U6317 (N_6317,N_2881,N_355);
and U6318 (N_6318,N_2540,N_3289);
nor U6319 (N_6319,N_2427,N_4989);
xor U6320 (N_6320,N_4978,N_4922);
or U6321 (N_6321,N_1085,N_248);
nand U6322 (N_6322,N_282,N_1465);
and U6323 (N_6323,N_2752,N_2324);
nor U6324 (N_6324,N_4419,N_4970);
or U6325 (N_6325,N_4509,N_1763);
nand U6326 (N_6326,N_2064,N_4243);
nor U6327 (N_6327,N_3832,N_2846);
xnor U6328 (N_6328,N_285,N_4513);
nand U6329 (N_6329,N_2744,N_433);
xnor U6330 (N_6330,N_2983,N_1319);
nand U6331 (N_6331,N_2467,N_576);
nand U6332 (N_6332,N_4650,N_3656);
or U6333 (N_6333,N_4490,N_368);
xnor U6334 (N_6334,N_1968,N_1140);
nand U6335 (N_6335,N_1569,N_2879);
nor U6336 (N_6336,N_116,N_3273);
or U6337 (N_6337,N_3484,N_4912);
nor U6338 (N_6338,N_16,N_2782);
xor U6339 (N_6339,N_3760,N_1439);
nor U6340 (N_6340,N_2335,N_2147);
or U6341 (N_6341,N_2889,N_1829);
nor U6342 (N_6342,N_3268,N_4298);
or U6343 (N_6343,N_1958,N_3437);
xnor U6344 (N_6344,N_860,N_2505);
xor U6345 (N_6345,N_3570,N_1342);
nand U6346 (N_6346,N_1337,N_4073);
nor U6347 (N_6347,N_3230,N_2014);
nor U6348 (N_6348,N_3706,N_2632);
nand U6349 (N_6349,N_1555,N_91);
xnor U6350 (N_6350,N_4459,N_3947);
nand U6351 (N_6351,N_1896,N_429);
nand U6352 (N_6352,N_2385,N_3112);
and U6353 (N_6353,N_1868,N_842);
or U6354 (N_6354,N_702,N_118);
or U6355 (N_6355,N_2749,N_1441);
xnor U6356 (N_6356,N_1780,N_3640);
nand U6357 (N_6357,N_1931,N_950);
xor U6358 (N_6358,N_2558,N_4878);
and U6359 (N_6359,N_2750,N_3721);
and U6360 (N_6360,N_3494,N_3669);
xnor U6361 (N_6361,N_2630,N_3117);
or U6362 (N_6362,N_1646,N_1771);
nor U6363 (N_6363,N_3461,N_1762);
and U6364 (N_6364,N_934,N_2115);
and U6365 (N_6365,N_1173,N_1298);
nand U6366 (N_6366,N_2389,N_202);
and U6367 (N_6367,N_4936,N_4713);
and U6368 (N_6368,N_975,N_3665);
or U6369 (N_6369,N_3407,N_2952);
nor U6370 (N_6370,N_0,N_3136);
and U6371 (N_6371,N_3242,N_3805);
or U6372 (N_6372,N_1632,N_1645);
or U6373 (N_6373,N_374,N_1560);
nor U6374 (N_6374,N_1409,N_2992);
nand U6375 (N_6375,N_2011,N_2537);
xnor U6376 (N_6376,N_1701,N_4933);
xor U6377 (N_6377,N_2065,N_1750);
nor U6378 (N_6378,N_4728,N_2345);
nand U6379 (N_6379,N_2832,N_494);
xnor U6380 (N_6380,N_472,N_895);
or U6381 (N_6381,N_13,N_3869);
or U6382 (N_6382,N_2958,N_956);
or U6383 (N_6383,N_3470,N_3438);
or U6384 (N_6384,N_1592,N_4032);
xnor U6385 (N_6385,N_4042,N_828);
nand U6386 (N_6386,N_3792,N_286);
and U6387 (N_6387,N_1106,N_1251);
and U6388 (N_6388,N_243,N_3472);
and U6389 (N_6389,N_3883,N_1956);
nand U6390 (N_6390,N_4797,N_4240);
or U6391 (N_6391,N_1538,N_1856);
nand U6392 (N_6392,N_4836,N_3159);
or U6393 (N_6393,N_2414,N_3773);
and U6394 (N_6394,N_301,N_4601);
or U6395 (N_6395,N_2098,N_2980);
nand U6396 (N_6396,N_2695,N_3907);
or U6397 (N_6397,N_1966,N_1660);
xor U6398 (N_6398,N_3590,N_859);
xor U6399 (N_6399,N_2991,N_4476);
nor U6400 (N_6400,N_2002,N_4632);
and U6401 (N_6401,N_2489,N_2605);
and U6402 (N_6402,N_4306,N_3707);
nand U6403 (N_6403,N_4806,N_4427);
and U6404 (N_6404,N_2329,N_4303);
and U6405 (N_6405,N_1845,N_2851);
nor U6406 (N_6406,N_2764,N_873);
and U6407 (N_6407,N_2185,N_2969);
xor U6408 (N_6408,N_777,N_748);
nor U6409 (N_6409,N_4172,N_851);
nor U6410 (N_6410,N_2915,N_455);
nor U6411 (N_6411,N_4589,N_875);
and U6412 (N_6412,N_4762,N_2284);
or U6413 (N_6413,N_4789,N_423);
and U6414 (N_6414,N_669,N_2161);
nand U6415 (N_6415,N_2574,N_731);
xor U6416 (N_6416,N_3496,N_4612);
nand U6417 (N_6417,N_428,N_3000);
xor U6418 (N_6418,N_4198,N_3881);
and U6419 (N_6419,N_222,N_4405);
xnor U6420 (N_6420,N_4890,N_4894);
xnor U6421 (N_6421,N_653,N_3753);
nor U6422 (N_6422,N_1501,N_2937);
and U6423 (N_6423,N_4279,N_3032);
or U6424 (N_6424,N_227,N_3671);
xor U6425 (N_6425,N_1761,N_4599);
and U6426 (N_6426,N_1879,N_1451);
or U6427 (N_6427,N_410,N_3063);
and U6428 (N_6428,N_2031,N_3961);
xnor U6429 (N_6429,N_1719,N_3016);
nand U6430 (N_6430,N_3217,N_273);
and U6431 (N_6431,N_4803,N_2636);
nand U6432 (N_6432,N_1515,N_4300);
nor U6433 (N_6433,N_2756,N_2293);
nor U6434 (N_6434,N_917,N_1360);
and U6435 (N_6435,N_1529,N_126);
nor U6436 (N_6436,N_2584,N_3856);
and U6437 (N_6437,N_2211,N_2368);
xnor U6438 (N_6438,N_1653,N_2826);
nand U6439 (N_6439,N_1305,N_1040);
nor U6440 (N_6440,N_1381,N_595);
xnor U6441 (N_6441,N_1668,N_1012);
or U6442 (N_6442,N_3566,N_2045);
xor U6443 (N_6443,N_663,N_3034);
xor U6444 (N_6444,N_3104,N_1724);
nand U6445 (N_6445,N_1051,N_1143);
and U6446 (N_6446,N_1333,N_3137);
xor U6447 (N_6447,N_3337,N_888);
nor U6448 (N_6448,N_835,N_2472);
or U6449 (N_6449,N_3368,N_4278);
nor U6450 (N_6450,N_2549,N_4824);
and U6451 (N_6451,N_1524,N_3759);
xor U6452 (N_6452,N_3569,N_4744);
nand U6453 (N_6453,N_3221,N_3280);
xor U6454 (N_6454,N_1462,N_514);
nand U6455 (N_6455,N_4354,N_3443);
xnor U6456 (N_6456,N_2228,N_3266);
nand U6457 (N_6457,N_4111,N_2884);
nand U6458 (N_6458,N_3528,N_1978);
xnor U6459 (N_6459,N_1616,N_3130);
and U6460 (N_6460,N_2611,N_67);
xor U6461 (N_6461,N_1696,N_967);
xnor U6462 (N_6462,N_1053,N_2607);
or U6463 (N_6463,N_3045,N_4227);
nand U6464 (N_6464,N_2173,N_2664);
or U6465 (N_6465,N_19,N_953);
and U6466 (N_6466,N_900,N_420);
and U6467 (N_6467,N_789,N_1294);
and U6468 (N_6468,N_3891,N_3799);
or U6469 (N_6469,N_413,N_816);
and U6470 (N_6470,N_230,N_4561);
or U6471 (N_6471,N_3333,N_1174);
nand U6472 (N_6472,N_4671,N_1186);
nor U6473 (N_6473,N_4322,N_4681);
xor U6474 (N_6474,N_153,N_1558);
nand U6475 (N_6475,N_2096,N_2336);
nand U6476 (N_6476,N_2805,N_2347);
or U6477 (N_6477,N_1712,N_3727);
nor U6478 (N_6478,N_1203,N_1098);
xor U6479 (N_6479,N_448,N_1604);
xor U6480 (N_6480,N_2338,N_1942);
and U6481 (N_6481,N_1773,N_1236);
and U6482 (N_6482,N_386,N_2731);
xor U6483 (N_6483,N_1688,N_3630);
nand U6484 (N_6484,N_968,N_2858);
or U6485 (N_6485,N_2506,N_1953);
xnor U6486 (N_6486,N_4687,N_2079);
or U6487 (N_6487,N_252,N_3220);
nor U6488 (N_6488,N_1297,N_4407);
nor U6489 (N_6489,N_3377,N_4053);
and U6490 (N_6490,N_414,N_193);
nor U6491 (N_6491,N_932,N_3415);
and U6492 (N_6492,N_483,N_1477);
nand U6493 (N_6493,N_3441,N_674);
or U6494 (N_6494,N_1459,N_1786);
xor U6495 (N_6495,N_1830,N_2075);
nand U6496 (N_6496,N_3730,N_4109);
nand U6497 (N_6497,N_343,N_411);
nand U6498 (N_6498,N_4106,N_391);
nor U6499 (N_6499,N_1356,N_1394);
and U6500 (N_6500,N_3433,N_4795);
or U6501 (N_6501,N_80,N_2061);
and U6502 (N_6502,N_3710,N_954);
nand U6503 (N_6503,N_305,N_2210);
nor U6504 (N_6504,N_4372,N_1498);
or U6505 (N_6505,N_813,N_2110);
and U6506 (N_6506,N_51,N_2341);
or U6507 (N_6507,N_3416,N_4689);
and U6508 (N_6508,N_217,N_1093);
nand U6509 (N_6509,N_4489,N_4926);
or U6510 (N_6510,N_3095,N_250);
xor U6511 (N_6511,N_4929,N_4857);
or U6512 (N_6512,N_795,N_3619);
nor U6513 (N_6513,N_4013,N_4148);
nor U6514 (N_6514,N_401,N_1971);
xnor U6515 (N_6515,N_3383,N_4908);
nor U6516 (N_6516,N_1511,N_1259);
xnor U6517 (N_6517,N_2192,N_379);
or U6518 (N_6518,N_3209,N_1977);
xnor U6519 (N_6519,N_803,N_830);
and U6520 (N_6520,N_66,N_2351);
or U6521 (N_6521,N_4324,N_1209);
nor U6522 (N_6522,N_3940,N_2797);
or U6523 (N_6523,N_4460,N_2617);
nor U6524 (N_6524,N_4315,N_3018);
and U6525 (N_6525,N_384,N_3228);
nor U6526 (N_6526,N_129,N_4817);
nand U6527 (N_6527,N_1383,N_4261);
or U6528 (N_6528,N_4485,N_4285);
and U6529 (N_6529,N_1197,N_661);
xor U6530 (N_6530,N_998,N_4682);
nor U6531 (N_6531,N_3973,N_2320);
xor U6532 (N_6532,N_3393,N_475);
and U6533 (N_6533,N_3991,N_4382);
nor U6534 (N_6534,N_769,N_3928);
nand U6535 (N_6535,N_4802,N_2788);
nor U6536 (N_6536,N_4778,N_509);
nor U6537 (N_6537,N_2062,N_1975);
xnor U6538 (N_6538,N_1686,N_2286);
and U6539 (N_6539,N_4467,N_944);
and U6540 (N_6540,N_3564,N_4031);
nand U6541 (N_6541,N_3738,N_4406);
and U6542 (N_6542,N_3256,N_894);
nor U6543 (N_6543,N_4059,N_2331);
nand U6544 (N_6544,N_925,N_4861);
and U6545 (N_6545,N_32,N_2597);
nor U6546 (N_6546,N_4775,N_2930);
xor U6547 (N_6547,N_747,N_4268);
xnor U6548 (N_6548,N_4862,N_4304);
or U6549 (N_6549,N_3051,N_3479);
nor U6550 (N_6550,N_521,N_943);
and U6551 (N_6551,N_1463,N_3091);
xor U6552 (N_6552,N_4349,N_2076);
xnor U6553 (N_6553,N_1325,N_1623);
xnor U6554 (N_6554,N_4653,N_716);
nor U6555 (N_6555,N_1585,N_2552);
xnor U6556 (N_6556,N_3497,N_2748);
nor U6557 (N_6557,N_2594,N_2087);
xnor U6558 (N_6558,N_1274,N_2498);
and U6559 (N_6559,N_4872,N_4260);
and U6560 (N_6560,N_4466,N_2203);
xnor U6561 (N_6561,N_3312,N_3363);
xnor U6562 (N_6562,N_1714,N_359);
nor U6563 (N_6563,N_3102,N_2078);
nor U6564 (N_6564,N_4326,N_3974);
xnor U6565 (N_6565,N_4264,N_1502);
xnor U6566 (N_6566,N_1807,N_3606);
nor U6567 (N_6567,N_332,N_3477);
or U6568 (N_6568,N_3999,N_4524);
nand U6569 (N_6569,N_891,N_2119);
and U6570 (N_6570,N_1266,N_3965);
xor U6571 (N_6571,N_820,N_2720);
nand U6572 (N_6572,N_3292,N_2485);
xor U6573 (N_6573,N_4479,N_2386);
and U6574 (N_6574,N_4167,N_1530);
and U6575 (N_6575,N_1225,N_2977);
nand U6576 (N_6576,N_4180,N_2256);
xnor U6577 (N_6577,N_2321,N_1321);
or U6578 (N_6578,N_2831,N_1287);
or U6579 (N_6579,N_4097,N_1991);
xnor U6580 (N_6580,N_3757,N_2474);
and U6581 (N_6581,N_3812,N_2438);
xnor U6582 (N_6582,N_1912,N_815);
nand U6583 (N_6583,N_4099,N_4761);
or U6584 (N_6584,N_1986,N_866);
nand U6585 (N_6585,N_3378,N_1354);
or U6586 (N_6586,N_2523,N_3341);
xor U6587 (N_6587,N_619,N_3977);
nor U6588 (N_6588,N_4188,N_1605);
or U6589 (N_6589,N_4404,N_1676);
nor U6590 (N_6590,N_4655,N_764);
or U6591 (N_6591,N_3155,N_6);
xnor U6592 (N_6592,N_3846,N_4037);
and U6593 (N_6593,N_3265,N_562);
nand U6594 (N_6594,N_2634,N_1883);
and U6595 (N_6595,N_1920,N_3328);
nor U6596 (N_6596,N_604,N_1005);
and U6597 (N_6597,N_1376,N_3955);
or U6598 (N_6598,N_618,N_2917);
xnor U6599 (N_6599,N_1574,N_356);
and U6600 (N_6600,N_147,N_1656);
and U6601 (N_6601,N_4210,N_3544);
or U6602 (N_6602,N_4242,N_872);
or U6603 (N_6603,N_184,N_1943);
nand U6604 (N_6604,N_4911,N_2941);
nand U6605 (N_6605,N_1291,N_1922);
xnor U6606 (N_6606,N_1105,N_1219);
xor U6607 (N_6607,N_3827,N_3789);
nor U6608 (N_6608,N_3283,N_3715);
and U6609 (N_6609,N_3701,N_3041);
and U6610 (N_6610,N_4588,N_2875);
and U6611 (N_6611,N_4465,N_3915);
and U6612 (N_6612,N_95,N_2227);
nand U6613 (N_6613,N_3267,N_3154);
or U6614 (N_6614,N_2716,N_2914);
and U6615 (N_6615,N_4694,N_4374);
nand U6616 (N_6616,N_1795,N_2134);
or U6617 (N_6617,N_1378,N_3156);
and U6618 (N_6618,N_3811,N_2478);
or U6619 (N_6619,N_4985,N_2136);
nor U6620 (N_6620,N_4623,N_3980);
nand U6621 (N_6621,N_1050,N_1772);
or U6622 (N_6622,N_2713,N_4968);
nor U6623 (N_6623,N_2040,N_2187);
nand U6624 (N_6624,N_2874,N_708);
and U6625 (N_6625,N_4408,N_3810);
xor U6626 (N_6626,N_4159,N_3610);
nor U6627 (N_6627,N_4248,N_570);
and U6628 (N_6628,N_4843,N_3431);
and U6629 (N_6629,N_3192,N_4014);
and U6630 (N_6630,N_2998,N_1341);
or U6631 (N_6631,N_2888,N_3317);
xor U6632 (N_6632,N_1300,N_736);
nand U6633 (N_6633,N_4008,N_1884);
nand U6634 (N_6634,N_4615,N_1839);
or U6635 (N_6635,N_1016,N_2925);
nand U6636 (N_6636,N_3893,N_3593);
xnor U6637 (N_6637,N_544,N_4594);
and U6638 (N_6638,N_3818,N_4930);
or U6639 (N_6639,N_2113,N_1279);
or U6640 (N_6640,N_3372,N_367);
and U6641 (N_6641,N_3364,N_3975);
nand U6642 (N_6642,N_4710,N_4751);
or U6643 (N_6643,N_1878,N_2466);
nand U6644 (N_6644,N_1111,N_4287);
nor U6645 (N_6645,N_1041,N_3938);
nor U6646 (N_6646,N_1999,N_3984);
xor U6647 (N_6647,N_1312,N_543);
or U6648 (N_6648,N_4805,N_2251);
xor U6649 (N_6649,N_4719,N_2995);
or U6650 (N_6650,N_843,N_921);
and U6651 (N_6651,N_3428,N_387);
and U6652 (N_6652,N_4604,N_2151);
xnor U6653 (N_6653,N_4780,N_54);
nor U6654 (N_6654,N_3750,N_2762);
nor U6655 (N_6655,N_664,N_297);
or U6656 (N_6656,N_753,N_3420);
nor U6657 (N_6657,N_510,N_1635);
nor U6658 (N_6658,N_1089,N_1673);
nand U6659 (N_6659,N_1578,N_4383);
nor U6660 (N_6660,N_4537,N_1677);
and U6661 (N_6661,N_2371,N_101);
nand U6662 (N_6662,N_4336,N_1769);
and U6663 (N_6663,N_3515,N_1617);
nand U6664 (N_6664,N_1115,N_1048);
and U6665 (N_6665,N_216,N_4607);
and U6666 (N_6666,N_2138,N_1742);
or U6667 (N_6667,N_1640,N_2432);
or U6668 (N_6668,N_4173,N_3361);
and U6669 (N_6669,N_3584,N_3952);
or U6670 (N_6670,N_1167,N_2887);
or U6671 (N_6671,N_786,N_3194);
or U6672 (N_6672,N_4161,N_327);
nor U6673 (N_6673,N_24,N_4834);
nor U6674 (N_6674,N_3677,N_4541);
nor U6675 (N_6675,N_1847,N_3439);
nor U6676 (N_6676,N_4636,N_1422);
or U6677 (N_6677,N_1135,N_3498);
and U6678 (N_6678,N_363,N_876);
or U6679 (N_6679,N_2849,N_3831);
nor U6680 (N_6680,N_643,N_616);
and U6681 (N_6681,N_4692,N_1513);
nor U6682 (N_6682,N_3954,N_656);
and U6683 (N_6683,N_3429,N_4555);
nor U6684 (N_6684,N_4030,N_3270);
nand U6685 (N_6685,N_1941,N_1363);
or U6686 (N_6686,N_4972,N_1434);
xor U6687 (N_6687,N_4905,N_1527);
nand U6688 (N_6688,N_1183,N_4596);
or U6689 (N_6689,N_148,N_3968);
xor U6690 (N_6690,N_1916,N_2408);
nor U6691 (N_6691,N_4864,N_3367);
and U6692 (N_6692,N_3703,N_3330);
and U6693 (N_6693,N_289,N_3642);
xor U6694 (N_6694,N_4115,N_480);
or U6695 (N_6695,N_763,N_1214);
xnor U6696 (N_6696,N_2267,N_452);
xor U6697 (N_6697,N_2049,N_1288);
and U6698 (N_6698,N_2237,N_3752);
or U6699 (N_6699,N_1850,N_2157);
xnor U6700 (N_6700,N_2855,N_2019);
nand U6701 (N_6701,N_3405,N_1260);
and U6702 (N_6702,N_810,N_1223);
nor U6703 (N_6703,N_1256,N_1520);
and U6704 (N_6704,N_4254,N_1313);
nand U6705 (N_6705,N_4133,N_655);
or U6706 (N_6706,N_1264,N_3);
nor U6707 (N_6707,N_131,N_4038);
xnor U6708 (N_6708,N_582,N_4885);
and U6709 (N_6709,N_4568,N_3551);
xnor U6710 (N_6710,N_3863,N_855);
xor U6711 (N_6711,N_1278,N_3586);
and U6712 (N_6712,N_4176,N_3122);
xnor U6713 (N_6713,N_4766,N_4578);
nor U6714 (N_6714,N_2967,N_1909);
and U6715 (N_6715,N_2054,N_805);
xor U6716 (N_6716,N_2867,N_1528);
or U6717 (N_6717,N_3908,N_771);
or U6718 (N_6718,N_1809,N_14);
xnor U6719 (N_6719,N_194,N_3274);
xor U6720 (N_6720,N_840,N_512);
nor U6721 (N_6721,N_4353,N_3872);
and U6722 (N_6722,N_4347,N_4112);
or U6723 (N_6723,N_1454,N_1580);
xnor U6724 (N_6724,N_823,N_4675);
nor U6725 (N_6725,N_4691,N_1620);
or U6726 (N_6726,N_2129,N_1549);
or U6727 (N_6727,N_2107,N_749);
nand U6728 (N_6728,N_4143,N_3692);
nor U6729 (N_6729,N_362,N_4701);
nand U6730 (N_6730,N_3666,N_3362);
or U6731 (N_6731,N_1751,N_4918);
nand U6732 (N_6732,N_296,N_4044);
xor U6733 (N_6733,N_4652,N_1960);
and U6734 (N_6734,N_1890,N_4928);
or U6735 (N_6735,N_477,N_1485);
or U6736 (N_6736,N_1217,N_2845);
xnor U6737 (N_6737,N_4781,N_4752);
nor U6738 (N_6738,N_4660,N_1055);
xnor U6739 (N_6739,N_85,N_2868);
and U6740 (N_6740,N_2872,N_3129);
and U6741 (N_6741,N_2531,N_545);
nand U6742 (N_6742,N_2647,N_4902);
and U6743 (N_6743,N_484,N_4705);
nand U6744 (N_6744,N_1284,N_695);
and U6745 (N_6745,N_933,N_4246);
or U6746 (N_6746,N_877,N_3695);
nand U6747 (N_6747,N_1789,N_3525);
or U6748 (N_6748,N_4731,N_4868);
nand U6749 (N_6749,N_4914,N_4644);
xnor U6750 (N_6750,N_4639,N_2796);
nand U6751 (N_6751,N_2252,N_1424);
nor U6752 (N_6752,N_3153,N_3921);
xor U6753 (N_6753,N_4642,N_630);
nor U6754 (N_6754,N_937,N_3847);
nand U6755 (N_6755,N_902,N_488);
xor U6756 (N_6756,N_4700,N_2957);
and U6757 (N_6757,N_4827,N_3277);
nand U6758 (N_6758,N_59,N_3769);
nor U6759 (N_6759,N_1493,N_1075);
nor U6760 (N_6760,N_2546,N_4820);
xor U6761 (N_6761,N_2938,N_4967);
or U6762 (N_6762,N_3613,N_4299);
xor U6763 (N_6763,N_2084,N_2601);
and U6764 (N_6764,N_1596,N_3718);
or U6765 (N_6765,N_1070,N_2702);
or U6766 (N_6766,N_473,N_4988);
or U6767 (N_6767,N_715,N_2299);
nor U6768 (N_6768,N_267,N_1854);
nand U6769 (N_6769,N_3616,N_3868);
nand U6770 (N_6770,N_1466,N_4430);
or U6771 (N_6771,N_231,N_3205);
nor U6772 (N_6772,N_3089,N_4748);
nand U6773 (N_6773,N_4721,N_1489);
nand U6774 (N_6774,N_3539,N_238);
and U6775 (N_6775,N_1700,N_3747);
nor U6776 (N_6776,N_723,N_2456);
nand U6777 (N_6777,N_677,N_288);
or U6778 (N_6778,N_1938,N_1316);
xnor U6779 (N_6779,N_1132,N_2639);
nor U6780 (N_6780,N_1329,N_3370);
and U6781 (N_6781,N_2191,N_1433);
nor U6782 (N_6782,N_4472,N_4543);
nor U6783 (N_6783,N_2024,N_1157);
xnor U6784 (N_6784,N_1158,N_3953);
and U6785 (N_6785,N_2572,N_60);
nand U6786 (N_6786,N_2786,N_579);
nand U6787 (N_6787,N_2960,N_82);
nand U6788 (N_6788,N_2104,N_2954);
nor U6789 (N_6789,N_1877,N_3796);
xnor U6790 (N_6790,N_1032,N_3044);
nor U6791 (N_6791,N_2415,N_3384);
and U6792 (N_6792,N_1467,N_676);
nand U6793 (N_6793,N_3118,N_2181);
nor U6794 (N_6794,N_3181,N_3410);
and U6795 (N_6795,N_3882,N_924);
nor U6796 (N_6796,N_3335,N_4034);
nor U6797 (N_6797,N_1534,N_4091);
xor U6798 (N_6798,N_4590,N_2067);
nor U6799 (N_6799,N_3724,N_122);
nand U6800 (N_6800,N_1014,N_4697);
and U6801 (N_6801,N_399,N_919);
xor U6802 (N_6802,N_4363,N_4600);
or U6803 (N_6803,N_98,N_4184);
and U6804 (N_6804,N_2230,N_4256);
nor U6805 (N_6805,N_983,N_4735);
nor U6806 (N_6806,N_3897,N_1907);
nand U6807 (N_6807,N_2864,N_1272);
xnor U6808 (N_6808,N_4023,N_3559);
or U6809 (N_6809,N_1532,N_801);
and U6810 (N_6810,N_1775,N_4359);
or U6811 (N_6811,N_515,N_4539);
nand U6812 (N_6812,N_3979,N_3708);
nor U6813 (N_6813,N_709,N_1738);
nor U6814 (N_6814,N_1430,N_3308);
xor U6815 (N_6815,N_470,N_4022);
or U6816 (N_6816,N_1161,N_4251);
xor U6817 (N_6817,N_395,N_4526);
xor U6818 (N_6818,N_1747,N_845);
nor U6819 (N_6819,N_1019,N_2220);
nor U6820 (N_6820,N_2970,N_1683);
or U6821 (N_6821,N_4345,N_2340);
nand U6822 (N_6822,N_1833,N_4117);
or U6823 (N_6823,N_4849,N_360);
nor U6824 (N_6824,N_3775,N_3314);
xnor U6825 (N_6825,N_2488,N_537);
and U6826 (N_6826,N_940,N_4955);
nor U6827 (N_6827,N_2339,N_3875);
nand U6828 (N_6828,N_2600,N_2802);
xnor U6829 (N_6829,N_4214,N_4313);
and U6830 (N_6830,N_3761,N_3440);
xnor U6831 (N_6831,N_3836,N_603);
nor U6832 (N_6832,N_2355,N_241);
nand U6833 (N_6833,N_4083,N_4269);
and U6834 (N_6834,N_2391,N_4720);
and U6835 (N_6835,N_1419,N_3604);
or U6836 (N_6836,N_2258,N_4944);
and U6837 (N_6837,N_1725,N_27);
nand U6838 (N_6838,N_936,N_1222);
or U6839 (N_6839,N_127,N_1548);
and U6840 (N_6840,N_652,N_3211);
nand U6841 (N_6841,N_1307,N_1004);
nor U6842 (N_6842,N_1730,N_3310);
and U6843 (N_6843,N_1177,N_4085);
and U6844 (N_6844,N_382,N_2028);
xor U6845 (N_6845,N_4614,N_901);
or U6846 (N_6846,N_744,N_4271);
nor U6847 (N_6847,N_4492,N_4643);
nor U6848 (N_6848,N_188,N_2257);
xnor U6849 (N_6849,N_2188,N_4993);
and U6850 (N_6850,N_3029,N_2578);
and U6851 (N_6851,N_1308,N_164);
xor U6852 (N_6852,N_1997,N_326);
nand U6853 (N_6853,N_4899,N_329);
nand U6854 (N_6854,N_313,N_2387);
nand U6855 (N_6855,N_3055,N_4072);
and U6856 (N_6856,N_1492,N_4573);
nand U6857 (N_6857,N_160,N_773);
nand U6858 (N_6858,N_963,N_4651);
nand U6859 (N_6859,N_2595,N_3605);
and U6860 (N_6860,N_4342,N_1718);
or U6861 (N_6861,N_651,N_1437);
nand U6862 (N_6862,N_1471,N_4110);
and U6863 (N_6863,N_981,N_1987);
nor U6864 (N_6864,N_1758,N_4229);
nor U6865 (N_6865,N_3850,N_292);
and U6866 (N_6866,N_4125,N_3187);
nor U6867 (N_6867,N_856,N_3734);
and U6868 (N_6868,N_1740,N_4645);
or U6869 (N_6869,N_3971,N_4145);
xnor U6870 (N_6870,N_3651,N_3260);
nor U6871 (N_6871,N_838,N_1028);
nand U6872 (N_6872,N_3231,N_265);
nand U6873 (N_6873,N_3583,N_3476);
xor U6874 (N_6874,N_1517,N_951);
nor U6875 (N_6875,N_4480,N_3478);
or U6876 (N_6876,N_140,N_462);
or U6877 (N_6877,N_453,N_2837);
and U6878 (N_6878,N_1505,N_2747);
xor U6879 (N_6879,N_3224,N_567);
and U6880 (N_6880,N_323,N_2800);
nor U6881 (N_6881,N_536,N_3837);
or U6882 (N_6882,N_3829,N_3972);
or U6883 (N_6883,N_1951,N_2694);
and U6884 (N_6884,N_4620,N_1650);
and U6885 (N_6885,N_2046,N_2758);
or U6886 (N_6886,N_1612,N_3150);
nor U6887 (N_6887,N_3638,N_3916);
nand U6888 (N_6888,N_3066,N_4670);
xnor U6889 (N_6889,N_109,N_137);
nand U6890 (N_6890,N_9,N_3553);
nor U6891 (N_6891,N_4413,N_1036);
or U6892 (N_6892,N_333,N_841);
and U6893 (N_6893,N_17,N_2460);
xor U6894 (N_6894,N_20,N_2013);
and U6895 (N_6895,N_77,N_1078);
and U6896 (N_6896,N_2734,N_2866);
or U6897 (N_6897,N_1539,N_2219);
or U6898 (N_6898,N_4223,N_1915);
nand U6899 (N_6899,N_2690,N_4718);
xor U6900 (N_6900,N_650,N_991);
or U6901 (N_6901,N_4135,N_3019);
nand U6902 (N_6902,N_2327,N_4495);
nand U6903 (N_6903,N_3726,N_792);
nor U6904 (N_6904,N_929,N_1952);
nor U6905 (N_6905,N_503,N_4773);
or U6906 (N_6906,N_2492,N_2933);
xnor U6907 (N_6907,N_351,N_3311);
xor U6908 (N_6908,N_1681,N_2971);
xor U6909 (N_6909,N_4081,N_4826);
or U6910 (N_6910,N_419,N_3342);
or U6911 (N_6911,N_2861,N_1624);
and U6912 (N_6912,N_2471,N_4576);
and U6913 (N_6913,N_3432,N_3306);
xnor U6914 (N_6914,N_4521,N_4);
nor U6915 (N_6915,N_4695,N_3922);
and U6916 (N_6916,N_2233,N_2204);
xor U6917 (N_6917,N_626,N_39);
nor U6918 (N_6918,N_2857,N_3020);
nand U6919 (N_6919,N_4947,N_589);
nor U6920 (N_6920,N_2318,N_3269);
or U6921 (N_6921,N_4887,N_1926);
nor U6922 (N_6922,N_1476,N_3988);
xnor U6923 (N_6923,N_1516,N_3248);
and U6924 (N_6924,N_4869,N_4089);
nor U6925 (N_6925,N_4976,N_2005);
nor U6926 (N_6926,N_2856,N_4448);
or U6927 (N_6927,N_1114,N_2357);
and U6928 (N_6928,N_2693,N_1423);
nand U6929 (N_6929,N_4791,N_1010);
or U6930 (N_6930,N_3059,N_4433);
nor U6931 (N_6931,N_4835,N_1770);
and U6932 (N_6932,N_2773,N_233);
and U6933 (N_6933,N_2407,N_4484);
and U6934 (N_6934,N_2779,N_157);
or U6935 (N_6935,N_3996,N_4706);
xnor U6936 (N_6936,N_4934,N_3675);
nor U6937 (N_6937,N_2499,N_1144);
or U6938 (N_6938,N_3886,N_1535);
and U6939 (N_6939,N_1352,N_3126);
nand U6940 (N_6940,N_261,N_1519);
xor U6941 (N_6941,N_817,N_2199);
and U6942 (N_6942,N_3152,N_2420);
nor U6943 (N_6943,N_834,N_235);
xor U6944 (N_6944,N_3530,N_4341);
and U6945 (N_6945,N_2565,N_2053);
or U6946 (N_6946,N_3819,N_2528);
or U6947 (N_6947,N_2086,N_4498);
or U6948 (N_6948,N_1292,N_2646);
xor U6949 (N_6949,N_4426,N_1126);
and U6950 (N_6950,N_1735,N_725);
xor U6951 (N_6951,N_2627,N_4393);
nand U6952 (N_6952,N_4777,N_183);
and U6953 (N_6953,N_2212,N_3382);
or U6954 (N_6954,N_1859,N_3896);
and U6955 (N_6955,N_1097,N_4542);
or U6956 (N_6956,N_4595,N_1134);
nand U6957 (N_6957,N_3492,N_189);
nand U6958 (N_6958,N_3099,N_4654);
and U6959 (N_6959,N_1009,N_755);
nand U6960 (N_6960,N_4888,N_558);
and U6961 (N_6961,N_3199,N_607);
xnor U6962 (N_6962,N_4730,N_1447);
nand U6963 (N_6963,N_4746,N_3634);
nand U6964 (N_6964,N_4910,N_4375);
and U6965 (N_6965,N_2301,N_1018);
nor U6966 (N_6966,N_3573,N_2670);
xor U6967 (N_6967,N_2793,N_2761);
and U6968 (N_6968,N_1816,N_793);
nor U6969 (N_6969,N_2457,N_1875);
nor U6970 (N_6970,N_2766,N_3887);
and U6971 (N_6971,N_3913,N_2553);
nor U6972 (N_6972,N_2972,N_2306);
and U6973 (N_6973,N_1818,N_1564);
nand U6974 (N_6974,N_3449,N_1069);
xnor U6975 (N_6975,N_1318,N_218);
xnor U6976 (N_6976,N_4040,N_3719);
nand U6977 (N_6977,N_2596,N_1906);
and U6978 (N_6978,N_3749,N_1710);
nor U6979 (N_6979,N_3725,N_1113);
xor U6980 (N_6980,N_4597,N_615);
nor U6981 (N_6981,N_4958,N_563);
nor U6982 (N_6982,N_3165,N_1674);
or U6983 (N_6983,N_4622,N_4907);
xor U6984 (N_6984,N_1774,N_182);
xnor U6985 (N_6985,N_4234,N_4486);
nor U6986 (N_6986,N_1973,N_3717);
or U6987 (N_6987,N_2504,N_2543);
or U6988 (N_6988,N_717,N_400);
or U6989 (N_6989,N_1702,N_2223);
xnor U6990 (N_6990,N_86,N_4759);
and U6991 (N_6991,N_2025,N_4661);
or U6992 (N_6992,N_1716,N_1495);
xnor U6993 (N_6993,N_1892,N_523);
or U6994 (N_6994,N_4916,N_2510);
nor U6995 (N_6995,N_4376,N_4975);
nor U6996 (N_6996,N_2806,N_3151);
xnor U6997 (N_6997,N_4477,N_4335);
nand U6998 (N_6998,N_1206,N_4734);
nor U6999 (N_6999,N_4896,N_3614);
and U7000 (N_7000,N_4379,N_829);
or U7001 (N_7001,N_201,N_1094);
xor U7002 (N_7002,N_3376,N_138);
or U7003 (N_7003,N_3679,N_1602);
nand U7004 (N_7004,N_2508,N_3914);
xnor U7005 (N_7005,N_1935,N_905);
and U7006 (N_7006,N_832,N_1088);
xnor U7007 (N_7007,N_831,N_3787);
xnor U7008 (N_7008,N_469,N_3512);
xnor U7009 (N_7009,N_1537,N_1468);
nor U7010 (N_7010,N_4151,N_575);
and U7011 (N_7011,N_3949,N_229);
and U7012 (N_7012,N_2435,N_1195);
or U7013 (N_7013,N_3196,N_2010);
nor U7014 (N_7014,N_1509,N_4496);
or U7015 (N_7015,N_4329,N_1525);
nor U7016 (N_7016,N_4853,N_1336);
xor U7017 (N_7017,N_2909,N_3501);
or U7018 (N_7018,N_4517,N_2218);
nand U7019 (N_7019,N_941,N_3935);
and U7020 (N_7020,N_4224,N_790);
or U7021 (N_7021,N_590,N_1995);
and U7022 (N_7022,N_43,N_4909);
and U7023 (N_7023,N_1745,N_2101);
xor U7024 (N_7024,N_2880,N_4321);
and U7025 (N_7025,N_4983,N_166);
nand U7026 (N_7026,N_2274,N_3297);
or U7027 (N_7027,N_2433,N_3663);
nor U7028 (N_7028,N_2530,N_658);
nand U7029 (N_7029,N_2395,N_402);
nand U7030 (N_7030,N_2769,N_2637);
nor U7031 (N_7031,N_2168,N_3208);
and U7032 (N_7032,N_2373,N_3485);
or U7033 (N_7033,N_1193,N_529);
nor U7034 (N_7034,N_2966,N_3424);
nand U7035 (N_7035,N_3450,N_3259);
xor U7036 (N_7036,N_4283,N_3350);
nor U7037 (N_7037,N_3941,N_4212);
and U7038 (N_7038,N_4136,N_76);
or U7039 (N_7039,N_986,N_4281);
or U7040 (N_7040,N_224,N_4738);
or U7041 (N_7041,N_4475,N_25);
and U7042 (N_7042,N_1334,N_2974);
and U7043 (N_7043,N_592,N_4580);
nand U7044 (N_7044,N_2163,N_3329);
xor U7045 (N_7045,N_2675,N_2735);
xnor U7046 (N_7046,N_1103,N_2536);
and U7047 (N_7047,N_1276,N_1663);
nor U7048 (N_7048,N_181,N_3093);
or U7049 (N_7049,N_3204,N_1335);
xnor U7050 (N_7050,N_3456,N_1705);
or U7051 (N_7051,N_4704,N_2352);
or U7052 (N_7052,N_1862,N_3011);
nor U7053 (N_7053,N_1137,N_3048);
nor U7054 (N_7054,N_2613,N_4398);
nor U7055 (N_7055,N_1817,N_3561);
nand U7056 (N_7056,N_4166,N_4464);
or U7057 (N_7057,N_1678,N_2871);
nand U7058 (N_7058,N_1386,N_1304);
xnor U7059 (N_7059,N_1117,N_2606);
nand U7060 (N_7060,N_3843,N_1145);
nor U7061 (N_7061,N_2865,N_4258);
nor U7062 (N_7062,N_1273,N_2817);
or U7063 (N_7063,N_3795,N_4937);
or U7064 (N_7064,N_3864,N_2701);
nor U7065 (N_7065,N_4189,N_587);
or U7066 (N_7066,N_2055,N_4241);
nor U7067 (N_7067,N_2798,N_2524);
nand U7068 (N_7068,N_1522,N_2799);
and U7069 (N_7069,N_4530,N_1723);
and U7070 (N_7070,N_264,N_1832);
xnor U7071 (N_7071,N_1357,N_2509);
xor U7072 (N_7072,N_4079,N_3608);
and U7073 (N_7073,N_647,N_4096);
and U7074 (N_7074,N_200,N_4093);
nand U7075 (N_7075,N_4179,N_2333);
nor U7076 (N_7076,N_3394,N_1303);
nor U7077 (N_7077,N_3660,N_1556);
nand U7078 (N_7078,N_2774,N_4556);
or U7079 (N_7079,N_4318,N_2850);
xor U7080 (N_7080,N_2425,N_1233);
nand U7081 (N_7081,N_2614,N_1146);
xor U7082 (N_7082,N_287,N_1526);
nor U7083 (N_7083,N_2776,N_4769);
xnor U7084 (N_7084,N_3664,N_4676);
xor U7085 (N_7085,N_3929,N_3963);
or U7086 (N_7086,N_1245,N_785);
nand U7087 (N_7087,N_4431,N_4865);
and U7088 (N_7088,N_2644,N_4420);
nor U7089 (N_7089,N_3904,N_3490);
nand U7090 (N_7090,N_4209,N_1863);
or U7091 (N_7091,N_113,N_1741);
nand U7092 (N_7092,N_2979,N_3969);
nor U7093 (N_7093,N_1913,N_548);
nor U7094 (N_7094,N_3237,N_583);
xor U7095 (N_7095,N_159,N_2214);
or U7096 (N_7096,N_2841,N_2564);
and U7097 (N_7097,N_254,N_1076);
nand U7098 (N_7098,N_4052,N_4674);
nor U7099 (N_7099,N_3395,N_2904);
and U7100 (N_7100,N_1503,N_185);
nand U7101 (N_7101,N_4171,N_3243);
or U7102 (N_7102,N_4570,N_1803);
nor U7103 (N_7103,N_3597,N_1682);
or U7104 (N_7104,N_1393,N_2422);
nor U7105 (N_7105,N_4788,N_107);
and U7106 (N_7106,N_4852,N_1940);
or U7107 (N_7107,N_4288,N_1121);
and U7108 (N_7108,N_2804,N_1590);
nand U7109 (N_7109,N_3956,N_1776);
nor U7110 (N_7110,N_489,N_2852);
nor U7111 (N_7111,N_3388,N_100);
or U7112 (N_7112,N_2490,N_2547);
and U7113 (N_7113,N_4898,N_1936);
or U7114 (N_7114,N_110,N_641);
or U7115 (N_7115,N_3068,N_557);
and U7116 (N_7116,N_4659,N_4699);
xnor U7117 (N_7117,N_4157,N_3729);
xor U7118 (N_7118,N_672,N_1277);
nand U7119 (N_7119,N_3381,N_1059);
or U7120 (N_7120,N_2854,N_1148);
nand U7121 (N_7121,N_867,N_886);
or U7122 (N_7122,N_2729,N_3487);
nor U7123 (N_7123,N_1568,N_3598);
or U7124 (N_7124,N_2621,N_4165);
and U7125 (N_7125,N_2334,N_4364);
nor U7126 (N_7126,N_330,N_291);
xor U7127 (N_7127,N_1255,N_4732);
xnor U7128 (N_7128,N_1790,N_2150);
and U7129 (N_7129,N_340,N_750);
nand U7130 (N_7130,N_4160,N_2034);
or U7131 (N_7131,N_689,N_398);
nand U7132 (N_7132,N_724,N_1275);
and U7133 (N_7133,N_746,N_4807);
or U7134 (N_7134,N_2,N_2089);
or U7135 (N_7135,N_4638,N_4357);
or U7136 (N_7136,N_94,N_594);
xnor U7137 (N_7137,N_818,N_212);
and U7138 (N_7138,N_4906,N_4515);
nand U7139 (N_7139,N_3222,N_4051);
or U7140 (N_7140,N_1054,N_4863);
nand U7141 (N_7141,N_3903,N_2285);
and U7142 (N_7142,N_3937,N_4635);
nor U7143 (N_7143,N_2532,N_779);
nor U7144 (N_7144,N_1035,N_1504);
or U7145 (N_7145,N_4483,N_4131);
nand U7146 (N_7146,N_4637,N_2296);
or U7147 (N_7147,N_2283,N_1244);
nor U7148 (N_7148,N_1783,N_2246);
nand U7149 (N_7149,N_2072,N_4021);
or U7150 (N_7150,N_760,N_1270);
or U7151 (N_7151,N_4320,N_2853);
and U7152 (N_7152,N_4399,N_1814);
xnor U7153 (N_7153,N_334,N_53);
xor U7154 (N_7154,N_4275,N_195);
nand U7155 (N_7155,N_2700,N_2343);
xor U7156 (N_7156,N_1129,N_3365);
xnor U7157 (N_7157,N_1811,N_2814);
or U7158 (N_7158,N_191,N_3189);
nand U7159 (N_7159,N_1654,N_2959);
nand U7160 (N_7160,N_4116,N_2402);
and U7161 (N_7161,N_2649,N_2727);
and U7162 (N_7162,N_3517,N_4162);
xnor U7163 (N_7163,N_3075,N_4199);
nand U7164 (N_7164,N_307,N_4845);
xnor U7165 (N_7165,N_2426,N_4707);
and U7166 (N_7166,N_1571,N_2949);
xnor U7167 (N_7167,N_3755,N_2353);
xnor U7168 (N_7168,N_2721,N_1031);
xnor U7169 (N_7169,N_4514,N_3859);
or U7170 (N_7170,N_4684,N_534);
xor U7171 (N_7171,N_3284,N_2514);
and U7172 (N_7172,N_588,N_378);
or U7173 (N_7173,N_3900,N_1824);
nand U7174 (N_7174,N_3123,N_622);
or U7175 (N_7175,N_1708,N_3839);
nand U7176 (N_7176,N_3454,N_631);
and U7177 (N_7177,N_266,N_3183);
nand U7178 (N_7178,N_377,N_712);
nor U7179 (N_7179,N_1610,N_2557);
nor U7180 (N_7180,N_1446,N_4265);
or U7181 (N_7181,N_4338,N_3959);
and U7182 (N_7182,N_4996,N_1293);
and U7183 (N_7183,N_3465,N_2106);
nand U7184 (N_7184,N_4066,N_2021);
and U7185 (N_7185,N_3794,N_2736);
nand U7186 (N_7186,N_915,N_426);
xor U7187 (N_7187,N_4120,N_1749);
or U7188 (N_7188,N_2122,N_3374);
xor U7189 (N_7189,N_949,N_3098);
nand U7190 (N_7190,N_2033,N_3488);
xor U7191 (N_7191,N_125,N_4239);
nand U7192 (N_7192,N_632,N_4917);
xor U7193 (N_7193,N_2349,N_161);
nor U7194 (N_7194,N_1881,N_2732);
or U7195 (N_7195,N_3588,N_2364);
nand U7196 (N_7196,N_1052,N_4424);
nor U7197 (N_7197,N_705,N_4377);
xnor U7198 (N_7198,N_274,N_3739);
xor U7199 (N_7199,N_29,N_572);
nand U7200 (N_7200,N_3158,N_1496);
xor U7201 (N_7201,N_4290,N_1985);
nand U7202 (N_7202,N_2567,N_47);
nor U7203 (N_7203,N_1523,N_2719);
nor U7204 (N_7204,N_3053,N_2463);
xnor U7205 (N_7205,N_3995,N_4801);
nor U7206 (N_7206,N_57,N_1579);
or U7207 (N_7207,N_2500,N_740);
nor U7208 (N_7208,N_2184,N_3036);
nand U7209 (N_7209,N_2934,N_2703);
and U7210 (N_7210,N_3531,N_2217);
and U7211 (N_7211,N_1122,N_1100);
nor U7212 (N_7212,N_1068,N_210);
nand U7213 (N_7213,N_2130,N_3563);
xnor U7214 (N_7214,N_3768,N_1232);
or U7215 (N_7215,N_784,N_4904);
and U7216 (N_7216,N_1728,N_1711);
and U7217 (N_7217,N_4163,N_4373);
xor U7218 (N_7218,N_3826,N_2441);
or U7219 (N_7219,N_2893,N_28);
nand U7220 (N_7220,N_3146,N_466);
nor U7221 (N_7221,N_3522,N_3731);
nand U7222 (N_7222,N_3567,N_4056);
and U7223 (N_7223,N_3966,N_4535);
nand U7224 (N_7224,N_844,N_1340);
nand U7225 (N_7225,N_3422,N_1414);
and U7226 (N_7226,N_304,N_2503);
and U7227 (N_7227,N_3777,N_2144);
and U7228 (N_7228,N_4226,N_811);
or U7229 (N_7229,N_3637,N_4848);
or U7230 (N_7230,N_4284,N_1149);
nor U7231 (N_7231,N_73,N_3764);
nand U7232 (N_7232,N_3636,N_97);
or U7233 (N_7233,N_4938,N_1908);
xor U7234 (N_7234,N_3943,N_2961);
nand U7235 (N_7235,N_4520,N_4617);
and U7236 (N_7236,N_143,N_1930);
nor U7237 (N_7237,N_3457,N_2323);
and U7238 (N_7238,N_4232,N_3409);
and U7239 (N_7239,N_4395,N_3722);
xnor U7240 (N_7240,N_2406,N_2140);
nand U7241 (N_7241,N_1835,N_3698);
nor U7242 (N_7242,N_1969,N_2522);
and U7243 (N_7243,N_1190,N_4971);
nand U7244 (N_7244,N_2302,N_3462);
and U7245 (N_7245,N_1852,N_2559);
xnor U7246 (N_7246,N_64,N_4438);
nor U7247 (N_7247,N_279,N_2416);
nor U7248 (N_7248,N_2608,N_692);
and U7249 (N_7249,N_213,N_2696);
or U7250 (N_7250,N_2332,N_3444);
or U7251 (N_7251,N_133,N_1974);
nor U7252 (N_7252,N_2975,N_3702);
nand U7253 (N_7253,N_1499,N_996);
nor U7254 (N_7254,N_596,N_598);
and U7255 (N_7255,N_3043,N_2819);
and U7256 (N_7256,N_2951,N_1736);
nand U7257 (N_7257,N_1067,N_4206);
and U7258 (N_7258,N_952,N_344);
nand U7259 (N_7259,N_2692,N_310);
nand U7260 (N_7260,N_1840,N_690);
nand U7261 (N_7261,N_1626,N_4880);
nand U7262 (N_7262,N_2388,N_3216);
or U7263 (N_7263,N_4343,N_3879);
and U7264 (N_7264,N_15,N_2197);
and U7265 (N_7265,N_1990,N_2843);
nor U7266 (N_7266,N_947,N_1165);
nand U7267 (N_7267,N_3319,N_4649);
nand U7268 (N_7268,N_756,N_3371);
and U7269 (N_7269,N_4818,N_1691);
and U7270 (N_7270,N_849,N_2207);
and U7271 (N_7271,N_3083,N_3803);
nand U7272 (N_7272,N_454,N_3911);
or U7273 (N_7273,N_84,N_2434);
or U7274 (N_7274,N_1849,N_2361);
and U7275 (N_7275,N_1387,N_2216);
nand U7276 (N_7276,N_4230,N_2015);
nor U7277 (N_7277,N_1344,N_671);
nor U7278 (N_7278,N_4952,N_1066);
nand U7279 (N_7279,N_4825,N_3918);
and U7280 (N_7280,N_3106,N_2464);
or U7281 (N_7281,N_3163,N_1317);
nand U7282 (N_7282,N_3013,N_150);
or U7283 (N_7283,N_38,N_4217);
xnor U7284 (N_7284,N_2125,N_1349);
xnor U7285 (N_7285,N_1925,N_852);
nor U7286 (N_7286,N_1457,N_2182);
xor U7287 (N_7287,N_2337,N_3648);
nor U7288 (N_7288,N_416,N_2322);
nand U7289 (N_7289,N_928,N_3085);
nor U7290 (N_7290,N_2117,N_1853);
nand U7291 (N_7291,N_2149,N_4471);
and U7292 (N_7292,N_1265,N_542);
and U7293 (N_7293,N_1746,N_2231);
or U7294 (N_7294,N_393,N_1488);
nand U7295 (N_7295,N_2436,N_2603);
xnor U7296 (N_7296,N_635,N_3705);
or U7297 (N_7297,N_2317,N_3643);
nor U7298 (N_7298,N_566,N_4098);
nor U7299 (N_7299,N_896,N_770);
nor U7300 (N_7300,N_3646,N_2615);
nand U7301 (N_7301,N_3845,N_4048);
or U7302 (N_7302,N_2093,N_4628);
nand U7303 (N_7303,N_2688,N_4220);
nor U7304 (N_7304,N_3712,N_1418);
or U7305 (N_7305,N_1249,N_1597);
and U7306 (N_7306,N_2226,N_533);
and U7307 (N_7307,N_990,N_3127);
nand U7308 (N_7308,N_3632,N_3866);
and U7309 (N_7309,N_1138,N_614);
and U7310 (N_7310,N_4582,N_3833);
nor U7311 (N_7311,N_2142,N_357);
and U7312 (N_7312,N_1687,N_4527);
nand U7313 (N_7313,N_174,N_4277);
and U7314 (N_7314,N_1119,N_2155);
xor U7315 (N_7315,N_573,N_56);
and U7316 (N_7316,N_2829,N_371);
nor U7317 (N_7317,N_4915,N_2222);
nor U7318 (N_7318,N_2784,N_931);
or U7319 (N_7319,N_4708,N_2525);
nand U7320 (N_7320,N_1377,N_1720);
xnor U7321 (N_7321,N_2658,N_2043);
nand U7322 (N_7322,N_4138,N_430);
and U7323 (N_7323,N_2305,N_3179);
nor U7324 (N_7324,N_2870,N_375);
xor U7325 (N_7325,N_3802,N_3250);
nand U7326 (N_7326,N_3240,N_1120);
xnor U7327 (N_7327,N_4792,N_4586);
and U7328 (N_7328,N_4077,N_1123);
nand U7329 (N_7329,N_1697,N_955);
nand U7330 (N_7330,N_4069,N_496);
nand U7331 (N_7331,N_2830,N_4250);
nor U7332 (N_7332,N_1090,N_2526);
or U7333 (N_7333,N_3002,N_319);
xnor U7334 (N_7334,N_1834,N_3321);
and U7335 (N_7335,N_735,N_2238);
xnor U7336 (N_7336,N_3813,N_4774);
nand U7337 (N_7337,N_3934,N_878);
xnor U7338 (N_7338,N_3798,N_4437);
xor U7339 (N_7339,N_4867,N_1007);
nor U7340 (N_7340,N_624,N_2383);
nor U7341 (N_7341,N_4679,N_4571);
nor U7342 (N_7342,N_3390,N_3548);
xnor U7343 (N_7343,N_1204,N_504);
nor U7344 (N_7344,N_2074,N_3094);
and U7345 (N_7345,N_2924,N_1482);
nor U7346 (N_7346,N_4446,N_3990);
nor U7347 (N_7347,N_2475,N_1957);
nand U7348 (N_7348,N_4633,N_4500);
and U7349 (N_7349,N_3467,N_260);
nand U7350 (N_7350,N_2931,N_4924);
or U7351 (N_7351,N_4727,N_743);
and U7352 (N_7352,N_1358,N_4688);
nand U7353 (N_7353,N_2421,N_2588);
or U7354 (N_7354,N_2718,N_3696);
xnor U7355 (N_7355,N_2120,N_2165);
or U7356 (N_7356,N_684,N_3607);
or U7357 (N_7357,N_4169,N_808);
xor U7358 (N_7358,N_993,N_1379);
nor U7359 (N_7359,N_2001,N_3227);
nor U7360 (N_7360,N_8,N_4028);
nor U7361 (N_7361,N_1621,N_734);
xnor U7362 (N_7362,N_3782,N_1262);
nand U7363 (N_7363,N_1412,N_3483);
nor U7364 (N_7364,N_1599,N_636);
xor U7365 (N_7365,N_4884,N_1401);
and U7366 (N_7366,N_4043,N_4222);
or U7367 (N_7367,N_4036,N_1846);
nor U7368 (N_7368,N_4207,N_1299);
nor U7369 (N_7369,N_2367,N_3645);
or U7370 (N_7370,N_2783,N_1417);
nor U7371 (N_7371,N_3751,N_381);
nor U7372 (N_7372,N_3894,N_275);
nor U7373 (N_7373,N_3895,N_4202);
and U7374 (N_7374,N_1939,N_154);
and U7375 (N_7375,N_3062,N_2097);
nand U7376 (N_7376,N_2669,N_1033);
xor U7377 (N_7377,N_1901,N_2083);
or U7378 (N_7378,N_208,N_3366);
nand U7379 (N_7379,N_4753,N_3315);
nor U7380 (N_7380,N_2950,N_145);
and U7381 (N_7381,N_4439,N_458);
xor U7382 (N_7382,N_2179,N_4711);
xor U7383 (N_7383,N_259,N_1077);
nand U7384 (N_7384,N_2787,N_422);
or U7385 (N_7385,N_4074,N_646);
nor U7386 (N_7386,N_3455,N_1937);
nand U7387 (N_7387,N_4175,N_1168);
and U7388 (N_7388,N_2398,N_353);
nor U7389 (N_7389,N_2965,N_4187);
xnor U7390 (N_7390,N_3445,N_4564);
or U7391 (N_7391,N_1665,N_3821);
nor U7392 (N_7392,N_4001,N_392);
xnor U7393 (N_7393,N_3460,N_999);
nand U7394 (N_7394,N_3149,N_3982);
xor U7395 (N_7395,N_3858,N_1903);
and U7396 (N_7396,N_4680,N_4846);
or U7397 (N_7397,N_1213,N_4900);
xnor U7398 (N_7398,N_281,N_909);
xnor U7399 (N_7399,N_322,N_1267);
or U7400 (N_7400,N_4274,N_2417);
nand U7401 (N_7401,N_4750,N_3890);
xor U7402 (N_7402,N_691,N_2255);
or U7403 (N_7403,N_1347,N_3167);
xor U7404 (N_7404,N_3006,N_1079);
xor U7405 (N_7405,N_899,N_2585);
nor U7406 (N_7406,N_2224,N_3557);
nor U7407 (N_7407,N_4385,N_1787);
and U7408 (N_7408,N_826,N_987);
or U7409 (N_7409,N_4787,N_4560);
xor U7410 (N_7410,N_682,N_910);
xor U7411 (N_7411,N_2374,N_2453);
nor U7412 (N_7412,N_1449,N_1281);
nor U7413 (N_7413,N_3245,N_112);
nor U7414 (N_7414,N_4247,N_2873);
nor U7415 (N_7415,N_52,N_2697);
and U7416 (N_7416,N_4389,N_124);
or U7417 (N_7417,N_4442,N_3603);
nand U7418 (N_7418,N_1185,N_1948);
nand U7419 (N_7419,N_3387,N_3218);
xnor U7420 (N_7420,N_3009,N_4050);
and U7421 (N_7421,N_3300,N_3981);
nand U7422 (N_7422,N_1198,N_4540);
nand U7423 (N_7423,N_4919,N_269);
or U7424 (N_7424,N_4208,N_2008);
or U7425 (N_7425,N_1343,N_629);
nand U7426 (N_7426,N_35,N_4409);
nand U7427 (N_7427,N_3970,N_3817);
nor U7428 (N_7428,N_922,N_495);
or U7429 (N_7429,N_4174,N_3400);
nand U7430 (N_7430,N_2555,N_339);
nand U7431 (N_7431,N_681,N_3855);
nor U7432 (N_7432,N_2626,N_1998);
nand U7433 (N_7433,N_2913,N_4276);
xnor U7434 (N_7434,N_2476,N_3741);
nand U7435 (N_7435,N_752,N_1015);
or U7436 (N_7436,N_2249,N_2017);
or U7437 (N_7437,N_1743,N_2166);
nor U7438 (N_7438,N_1073,N_4502);
xor U7439 (N_7439,N_1649,N_1510);
nand U7440 (N_7440,N_83,N_2027);
and U7441 (N_7441,N_569,N_3425);
nand U7442 (N_7442,N_4493,N_2213);
xor U7443 (N_7443,N_432,N_40);
xnor U7444 (N_7444,N_892,N_4339);
and U7445 (N_7445,N_858,N_4745);
xor U7446 (N_7446,N_3397,N_4154);
xor U7447 (N_7447,N_3626,N_58);
and U7448 (N_7448,N_2754,N_1606);
nor U7449 (N_7449,N_2715,N_139);
or U7450 (N_7450,N_4625,N_4763);
and U7451 (N_7451,N_3545,N_1615);
nand U7452 (N_7452,N_3709,N_3174);
or U7453 (N_7453,N_1648,N_1506);
and U7454 (N_7454,N_4113,N_969);
nor U7455 (N_7455,N_2381,N_4506);
and U7456 (N_7456,N_463,N_3931);
xnor U7457 (N_7457,N_865,N_3021);
and U7458 (N_7458,N_524,N_2095);
nor U7459 (N_7459,N_219,N_1826);
xor U7460 (N_7460,N_2576,N_1448);
nor U7461 (N_7461,N_4205,N_1694);
nand U7462 (N_7462,N_1151,N_683);
and U7463 (N_7463,N_4244,N_2051);
and U7464 (N_7464,N_4893,N_1607);
nand U7465 (N_7465,N_2247,N_1252);
nor U7466 (N_7466,N_927,N_449);
nand U7467 (N_7467,N_3298,N_4673);
nand U7468 (N_7468,N_1628,N_2699);
nand U7469 (N_7469,N_3144,N_2575);
and U7470 (N_7470,N_4950,N_964);
nor U7471 (N_7471,N_3556,N_1857);
xnor U7472 (N_7472,N_2681,N_324);
or U7473 (N_7473,N_3356,N_204);
or U7474 (N_7474,N_1636,N_2940);
nor U7475 (N_7475,N_3763,N_718);
nor U7476 (N_7476,N_4005,N_2677);
xnor U7477 (N_7477,N_4529,N_3994);
or U7478 (N_7478,N_2170,N_4118);
or U7479 (N_7479,N_3835,N_751);
nand U7480 (N_7480,N_4873,N_1959);
xnor U7481 (N_7481,N_1765,N_871);
nand U7482 (N_7482,N_4945,N_1091);
xor U7483 (N_7483,N_1732,N_4949);
nor U7484 (N_7484,N_312,N_3255);
and U7485 (N_7485,N_1023,N_4352);
nand U7486 (N_7486,N_3910,N_3801);
nor U7487 (N_7487,N_4140,N_2768);
nor U7488 (N_7488,N_1345,N_2190);
and U7489 (N_7489,N_599,N_3668);
and U7490 (N_7490,N_3198,N_4238);
xnor U7491 (N_7491,N_1128,N_4613);
nand U7492 (N_7492,N_989,N_1927);
or U7493 (N_7493,N_3682,N_3901);
xor U7494 (N_7494,N_4740,N_3336);
xor U7495 (N_7495,N_1601,N_4185);
xor U7496 (N_7496,N_3164,N_4913);
or U7497 (N_7497,N_3507,N_372);
nand U7498 (N_7498,N_518,N_3711);
nand U7499 (N_7499,N_2346,N_4058);
xor U7500 (N_7500,N_849,N_3740);
xor U7501 (N_7501,N_57,N_627);
or U7502 (N_7502,N_3049,N_74);
xor U7503 (N_7503,N_3564,N_3755);
nand U7504 (N_7504,N_849,N_3904);
and U7505 (N_7505,N_150,N_2152);
and U7506 (N_7506,N_3471,N_1745);
nand U7507 (N_7507,N_1498,N_3840);
and U7508 (N_7508,N_793,N_3034);
and U7509 (N_7509,N_3764,N_3497);
xor U7510 (N_7510,N_1942,N_3110);
and U7511 (N_7511,N_4321,N_457);
or U7512 (N_7512,N_501,N_2615);
xnor U7513 (N_7513,N_2137,N_3623);
nor U7514 (N_7514,N_1383,N_1535);
or U7515 (N_7515,N_538,N_260);
and U7516 (N_7516,N_4952,N_4572);
or U7517 (N_7517,N_4309,N_3252);
nor U7518 (N_7518,N_3829,N_3163);
or U7519 (N_7519,N_4125,N_2708);
nor U7520 (N_7520,N_4783,N_2111);
nor U7521 (N_7521,N_4049,N_1475);
nand U7522 (N_7522,N_4916,N_2512);
or U7523 (N_7523,N_1421,N_4610);
and U7524 (N_7524,N_3426,N_4357);
nand U7525 (N_7525,N_2923,N_634);
and U7526 (N_7526,N_1631,N_2523);
or U7527 (N_7527,N_917,N_1968);
nor U7528 (N_7528,N_1651,N_2198);
xnor U7529 (N_7529,N_4575,N_4296);
xor U7530 (N_7530,N_1366,N_3493);
and U7531 (N_7531,N_4717,N_2226);
xnor U7532 (N_7532,N_2032,N_1657);
nor U7533 (N_7533,N_4750,N_2862);
or U7534 (N_7534,N_1527,N_808);
and U7535 (N_7535,N_2468,N_2961);
nand U7536 (N_7536,N_3071,N_180);
nand U7537 (N_7537,N_1941,N_1169);
and U7538 (N_7538,N_2461,N_951);
nand U7539 (N_7539,N_4796,N_951);
xnor U7540 (N_7540,N_556,N_4236);
or U7541 (N_7541,N_2571,N_3754);
nor U7542 (N_7542,N_206,N_3598);
nor U7543 (N_7543,N_2619,N_1697);
nand U7544 (N_7544,N_3815,N_4550);
nor U7545 (N_7545,N_3690,N_2472);
xor U7546 (N_7546,N_3797,N_1511);
or U7547 (N_7547,N_482,N_4460);
nand U7548 (N_7548,N_4435,N_3379);
nor U7549 (N_7549,N_4286,N_3663);
nand U7550 (N_7550,N_2309,N_731);
and U7551 (N_7551,N_144,N_65);
nor U7552 (N_7552,N_1264,N_3174);
and U7553 (N_7553,N_4598,N_2882);
and U7554 (N_7554,N_4415,N_917);
nor U7555 (N_7555,N_3103,N_2272);
nor U7556 (N_7556,N_4440,N_1906);
nor U7557 (N_7557,N_3929,N_2483);
xor U7558 (N_7558,N_751,N_4596);
nand U7559 (N_7559,N_482,N_4353);
xnor U7560 (N_7560,N_3,N_3620);
xnor U7561 (N_7561,N_631,N_3304);
nand U7562 (N_7562,N_2681,N_3088);
nand U7563 (N_7563,N_236,N_3491);
nor U7564 (N_7564,N_2234,N_3040);
and U7565 (N_7565,N_1283,N_4472);
nor U7566 (N_7566,N_4256,N_3708);
and U7567 (N_7567,N_4753,N_333);
nor U7568 (N_7568,N_2889,N_1987);
nand U7569 (N_7569,N_834,N_1736);
nand U7570 (N_7570,N_1148,N_3852);
xnor U7571 (N_7571,N_4986,N_304);
nor U7572 (N_7572,N_2136,N_3439);
nand U7573 (N_7573,N_508,N_4578);
nor U7574 (N_7574,N_626,N_783);
or U7575 (N_7575,N_2982,N_2446);
nand U7576 (N_7576,N_3889,N_1471);
nand U7577 (N_7577,N_715,N_119);
nand U7578 (N_7578,N_862,N_3354);
and U7579 (N_7579,N_3588,N_4774);
and U7580 (N_7580,N_3089,N_623);
nand U7581 (N_7581,N_1053,N_2583);
and U7582 (N_7582,N_4090,N_2274);
nand U7583 (N_7583,N_562,N_4306);
nand U7584 (N_7584,N_1754,N_4434);
nand U7585 (N_7585,N_2132,N_4297);
nand U7586 (N_7586,N_2454,N_1034);
nand U7587 (N_7587,N_3412,N_4267);
or U7588 (N_7588,N_1629,N_1136);
nand U7589 (N_7589,N_3450,N_1273);
nand U7590 (N_7590,N_2741,N_4091);
or U7591 (N_7591,N_2097,N_2656);
and U7592 (N_7592,N_4521,N_2858);
nor U7593 (N_7593,N_3693,N_2399);
and U7594 (N_7594,N_139,N_4464);
or U7595 (N_7595,N_3361,N_3119);
nand U7596 (N_7596,N_4585,N_848);
nor U7597 (N_7597,N_1275,N_162);
nand U7598 (N_7598,N_4216,N_865);
nand U7599 (N_7599,N_1857,N_2468);
xnor U7600 (N_7600,N_1465,N_1573);
or U7601 (N_7601,N_1962,N_4372);
xor U7602 (N_7602,N_4110,N_154);
xnor U7603 (N_7603,N_4019,N_1058);
or U7604 (N_7604,N_722,N_3764);
nor U7605 (N_7605,N_555,N_2550);
nand U7606 (N_7606,N_391,N_2945);
nor U7607 (N_7607,N_2381,N_4902);
nand U7608 (N_7608,N_3751,N_362);
and U7609 (N_7609,N_2210,N_1989);
xor U7610 (N_7610,N_2683,N_3222);
and U7611 (N_7611,N_2521,N_784);
xnor U7612 (N_7612,N_1215,N_2548);
or U7613 (N_7613,N_1366,N_3245);
nor U7614 (N_7614,N_4455,N_268);
nand U7615 (N_7615,N_3431,N_2660);
or U7616 (N_7616,N_1953,N_3945);
and U7617 (N_7617,N_2806,N_4852);
xor U7618 (N_7618,N_157,N_4069);
and U7619 (N_7619,N_1548,N_685);
nor U7620 (N_7620,N_4166,N_1259);
nand U7621 (N_7621,N_3901,N_6);
or U7622 (N_7622,N_2076,N_2646);
nor U7623 (N_7623,N_455,N_143);
and U7624 (N_7624,N_4350,N_1420);
nor U7625 (N_7625,N_1313,N_3355);
or U7626 (N_7626,N_3610,N_4066);
xor U7627 (N_7627,N_3369,N_3901);
nor U7628 (N_7628,N_4147,N_2549);
xor U7629 (N_7629,N_4051,N_2614);
nor U7630 (N_7630,N_862,N_4926);
and U7631 (N_7631,N_1262,N_4223);
xnor U7632 (N_7632,N_4143,N_4997);
nor U7633 (N_7633,N_1347,N_2892);
and U7634 (N_7634,N_3278,N_1924);
or U7635 (N_7635,N_4358,N_4050);
and U7636 (N_7636,N_2491,N_2407);
and U7637 (N_7637,N_2223,N_69);
nand U7638 (N_7638,N_2659,N_3563);
nor U7639 (N_7639,N_728,N_3003);
or U7640 (N_7640,N_4772,N_3416);
xor U7641 (N_7641,N_4552,N_2288);
nor U7642 (N_7642,N_3182,N_2200);
nor U7643 (N_7643,N_4064,N_1542);
xor U7644 (N_7644,N_2788,N_3455);
or U7645 (N_7645,N_4281,N_4696);
xnor U7646 (N_7646,N_3179,N_670);
nand U7647 (N_7647,N_752,N_4361);
xnor U7648 (N_7648,N_4369,N_2258);
nand U7649 (N_7649,N_4601,N_242);
nand U7650 (N_7650,N_4573,N_2991);
xnor U7651 (N_7651,N_1721,N_403);
nand U7652 (N_7652,N_2226,N_3961);
or U7653 (N_7653,N_217,N_4254);
xor U7654 (N_7654,N_4678,N_833);
xor U7655 (N_7655,N_1853,N_1729);
and U7656 (N_7656,N_3716,N_3011);
nand U7657 (N_7657,N_4735,N_1638);
xnor U7658 (N_7658,N_96,N_575);
nand U7659 (N_7659,N_2197,N_949);
nand U7660 (N_7660,N_1338,N_2524);
nor U7661 (N_7661,N_4624,N_1907);
xor U7662 (N_7662,N_527,N_54);
nand U7663 (N_7663,N_3083,N_4815);
nand U7664 (N_7664,N_1430,N_4767);
or U7665 (N_7665,N_1788,N_472);
nand U7666 (N_7666,N_3033,N_3193);
or U7667 (N_7667,N_4968,N_1752);
nand U7668 (N_7668,N_866,N_684);
nand U7669 (N_7669,N_1744,N_3310);
or U7670 (N_7670,N_2279,N_4984);
and U7671 (N_7671,N_151,N_3770);
xor U7672 (N_7672,N_275,N_3694);
nor U7673 (N_7673,N_4923,N_2213);
nand U7674 (N_7674,N_3657,N_2321);
and U7675 (N_7675,N_2066,N_1293);
nand U7676 (N_7676,N_2819,N_4694);
and U7677 (N_7677,N_2958,N_4756);
nor U7678 (N_7678,N_1272,N_253);
nor U7679 (N_7679,N_2657,N_1763);
xor U7680 (N_7680,N_1722,N_4216);
nand U7681 (N_7681,N_3372,N_248);
or U7682 (N_7682,N_900,N_275);
or U7683 (N_7683,N_2899,N_2770);
xnor U7684 (N_7684,N_3771,N_1901);
xor U7685 (N_7685,N_2959,N_552);
nand U7686 (N_7686,N_215,N_3571);
nor U7687 (N_7687,N_2500,N_1208);
or U7688 (N_7688,N_2766,N_3884);
and U7689 (N_7689,N_3663,N_834);
nor U7690 (N_7690,N_851,N_3219);
nor U7691 (N_7691,N_1372,N_74);
nor U7692 (N_7692,N_4528,N_2072);
and U7693 (N_7693,N_1032,N_903);
or U7694 (N_7694,N_1256,N_2061);
nand U7695 (N_7695,N_2790,N_1556);
and U7696 (N_7696,N_833,N_3723);
nor U7697 (N_7697,N_3919,N_4493);
or U7698 (N_7698,N_2083,N_41);
nand U7699 (N_7699,N_1049,N_1086);
nand U7700 (N_7700,N_2105,N_622);
nor U7701 (N_7701,N_4251,N_2932);
and U7702 (N_7702,N_2366,N_4784);
xor U7703 (N_7703,N_4103,N_3095);
and U7704 (N_7704,N_4326,N_4484);
and U7705 (N_7705,N_2251,N_1333);
nand U7706 (N_7706,N_3468,N_1266);
and U7707 (N_7707,N_2418,N_2443);
and U7708 (N_7708,N_4325,N_4331);
nor U7709 (N_7709,N_2364,N_4973);
or U7710 (N_7710,N_1176,N_923);
nand U7711 (N_7711,N_4340,N_3992);
nor U7712 (N_7712,N_2515,N_1920);
and U7713 (N_7713,N_4949,N_2771);
nor U7714 (N_7714,N_4657,N_2835);
and U7715 (N_7715,N_1483,N_4226);
nor U7716 (N_7716,N_242,N_3525);
xnor U7717 (N_7717,N_845,N_4403);
or U7718 (N_7718,N_3934,N_1990);
and U7719 (N_7719,N_1947,N_1240);
xor U7720 (N_7720,N_2317,N_1299);
xor U7721 (N_7721,N_1848,N_300);
or U7722 (N_7722,N_2110,N_4683);
xor U7723 (N_7723,N_4141,N_2919);
xnor U7724 (N_7724,N_393,N_960);
xor U7725 (N_7725,N_732,N_163);
xor U7726 (N_7726,N_99,N_4039);
nor U7727 (N_7727,N_2613,N_2286);
nor U7728 (N_7728,N_1560,N_1753);
or U7729 (N_7729,N_576,N_4226);
nand U7730 (N_7730,N_295,N_4893);
and U7731 (N_7731,N_4763,N_1046);
or U7732 (N_7732,N_437,N_2541);
nand U7733 (N_7733,N_1094,N_1757);
and U7734 (N_7734,N_2323,N_872);
nand U7735 (N_7735,N_3831,N_342);
xnor U7736 (N_7736,N_3613,N_4469);
nor U7737 (N_7737,N_4623,N_2076);
and U7738 (N_7738,N_4526,N_280);
nand U7739 (N_7739,N_1584,N_801);
xnor U7740 (N_7740,N_2175,N_2967);
or U7741 (N_7741,N_1629,N_3377);
xor U7742 (N_7742,N_2185,N_4790);
nor U7743 (N_7743,N_4465,N_4105);
xor U7744 (N_7744,N_3866,N_4573);
and U7745 (N_7745,N_301,N_3424);
nor U7746 (N_7746,N_4179,N_696);
xnor U7747 (N_7747,N_1813,N_3434);
nand U7748 (N_7748,N_2592,N_4402);
nand U7749 (N_7749,N_3528,N_4214);
nand U7750 (N_7750,N_114,N_3443);
nand U7751 (N_7751,N_1791,N_1941);
and U7752 (N_7752,N_1167,N_4507);
nand U7753 (N_7753,N_3761,N_822);
or U7754 (N_7754,N_17,N_353);
nor U7755 (N_7755,N_223,N_4397);
xor U7756 (N_7756,N_4009,N_2309);
or U7757 (N_7757,N_4491,N_4796);
and U7758 (N_7758,N_2179,N_4445);
and U7759 (N_7759,N_370,N_4761);
nand U7760 (N_7760,N_2463,N_4815);
and U7761 (N_7761,N_872,N_207);
or U7762 (N_7762,N_2682,N_338);
and U7763 (N_7763,N_3350,N_2800);
xnor U7764 (N_7764,N_4973,N_234);
or U7765 (N_7765,N_4432,N_4460);
xor U7766 (N_7766,N_1638,N_2197);
or U7767 (N_7767,N_4262,N_3912);
xor U7768 (N_7768,N_399,N_462);
nor U7769 (N_7769,N_2225,N_2082);
or U7770 (N_7770,N_1449,N_2293);
nor U7771 (N_7771,N_3618,N_2211);
and U7772 (N_7772,N_2981,N_2002);
nor U7773 (N_7773,N_805,N_3066);
nand U7774 (N_7774,N_101,N_836);
and U7775 (N_7775,N_1930,N_237);
nor U7776 (N_7776,N_4810,N_4746);
and U7777 (N_7777,N_3446,N_2752);
xnor U7778 (N_7778,N_3743,N_4881);
or U7779 (N_7779,N_825,N_4689);
nand U7780 (N_7780,N_2244,N_1085);
and U7781 (N_7781,N_404,N_4633);
or U7782 (N_7782,N_1724,N_651);
or U7783 (N_7783,N_4713,N_3264);
or U7784 (N_7784,N_796,N_3276);
nor U7785 (N_7785,N_291,N_1779);
xnor U7786 (N_7786,N_4173,N_293);
or U7787 (N_7787,N_3310,N_991);
nor U7788 (N_7788,N_1165,N_2477);
xnor U7789 (N_7789,N_1434,N_856);
and U7790 (N_7790,N_1055,N_2638);
or U7791 (N_7791,N_3792,N_1699);
or U7792 (N_7792,N_2573,N_4829);
or U7793 (N_7793,N_4970,N_2187);
nor U7794 (N_7794,N_222,N_2679);
nor U7795 (N_7795,N_3638,N_4553);
xnor U7796 (N_7796,N_3257,N_1049);
nand U7797 (N_7797,N_2136,N_304);
and U7798 (N_7798,N_2163,N_4727);
or U7799 (N_7799,N_1894,N_1282);
nor U7800 (N_7800,N_3753,N_2322);
and U7801 (N_7801,N_2704,N_1312);
and U7802 (N_7802,N_2790,N_2786);
nand U7803 (N_7803,N_3440,N_2997);
xor U7804 (N_7804,N_3273,N_4214);
nand U7805 (N_7805,N_2832,N_567);
nand U7806 (N_7806,N_4464,N_2928);
and U7807 (N_7807,N_2893,N_3147);
nand U7808 (N_7808,N_1349,N_1082);
xnor U7809 (N_7809,N_1386,N_4564);
nand U7810 (N_7810,N_3304,N_84);
nand U7811 (N_7811,N_1548,N_3947);
xor U7812 (N_7812,N_4081,N_3104);
xnor U7813 (N_7813,N_4737,N_1558);
xnor U7814 (N_7814,N_1754,N_1446);
nor U7815 (N_7815,N_2944,N_3911);
nand U7816 (N_7816,N_3546,N_1426);
and U7817 (N_7817,N_2855,N_2032);
nor U7818 (N_7818,N_4462,N_740);
or U7819 (N_7819,N_1980,N_580);
and U7820 (N_7820,N_2868,N_1910);
or U7821 (N_7821,N_2046,N_4541);
or U7822 (N_7822,N_2535,N_4912);
or U7823 (N_7823,N_249,N_1611);
xnor U7824 (N_7824,N_871,N_3668);
xor U7825 (N_7825,N_4994,N_3843);
nor U7826 (N_7826,N_3778,N_2534);
nand U7827 (N_7827,N_4346,N_2469);
xnor U7828 (N_7828,N_709,N_3848);
xor U7829 (N_7829,N_4458,N_4638);
and U7830 (N_7830,N_737,N_3517);
xor U7831 (N_7831,N_2724,N_418);
nand U7832 (N_7832,N_3156,N_4802);
nor U7833 (N_7833,N_69,N_3751);
or U7834 (N_7834,N_4225,N_4493);
and U7835 (N_7835,N_588,N_1644);
and U7836 (N_7836,N_2817,N_1191);
or U7837 (N_7837,N_2942,N_1575);
nand U7838 (N_7838,N_2542,N_3802);
xor U7839 (N_7839,N_958,N_4689);
nand U7840 (N_7840,N_486,N_1589);
nand U7841 (N_7841,N_3928,N_4935);
and U7842 (N_7842,N_4564,N_4848);
nand U7843 (N_7843,N_200,N_3602);
or U7844 (N_7844,N_2015,N_3042);
nor U7845 (N_7845,N_4581,N_2246);
or U7846 (N_7846,N_3437,N_2397);
nor U7847 (N_7847,N_3409,N_2525);
xnor U7848 (N_7848,N_4288,N_1899);
xnor U7849 (N_7849,N_4738,N_3173);
nor U7850 (N_7850,N_774,N_2972);
xnor U7851 (N_7851,N_2338,N_1630);
and U7852 (N_7852,N_3358,N_4588);
or U7853 (N_7853,N_3398,N_4782);
and U7854 (N_7854,N_172,N_4606);
and U7855 (N_7855,N_402,N_755);
and U7856 (N_7856,N_1502,N_896);
nand U7857 (N_7857,N_2566,N_4043);
nor U7858 (N_7858,N_4088,N_3136);
and U7859 (N_7859,N_4762,N_1273);
or U7860 (N_7860,N_3232,N_2746);
xnor U7861 (N_7861,N_2843,N_141);
or U7862 (N_7862,N_1573,N_4399);
or U7863 (N_7863,N_3107,N_2583);
nand U7864 (N_7864,N_3943,N_2119);
nor U7865 (N_7865,N_2935,N_2641);
nor U7866 (N_7866,N_4735,N_951);
nor U7867 (N_7867,N_1187,N_1235);
xor U7868 (N_7868,N_260,N_769);
nor U7869 (N_7869,N_4559,N_4509);
nand U7870 (N_7870,N_1243,N_1624);
nor U7871 (N_7871,N_3535,N_2281);
xor U7872 (N_7872,N_284,N_3981);
and U7873 (N_7873,N_2917,N_4872);
nand U7874 (N_7874,N_1467,N_4973);
and U7875 (N_7875,N_2561,N_2400);
or U7876 (N_7876,N_3028,N_1755);
or U7877 (N_7877,N_27,N_3512);
nand U7878 (N_7878,N_3152,N_2994);
xor U7879 (N_7879,N_2588,N_2194);
and U7880 (N_7880,N_4471,N_500);
nand U7881 (N_7881,N_1952,N_2229);
nor U7882 (N_7882,N_4687,N_0);
and U7883 (N_7883,N_3858,N_3759);
nand U7884 (N_7884,N_2683,N_3709);
or U7885 (N_7885,N_3381,N_4652);
nor U7886 (N_7886,N_2768,N_3789);
and U7887 (N_7887,N_3053,N_4396);
xor U7888 (N_7888,N_2719,N_452);
and U7889 (N_7889,N_1800,N_4239);
or U7890 (N_7890,N_2513,N_3019);
xnor U7891 (N_7891,N_3665,N_3544);
and U7892 (N_7892,N_2562,N_1875);
nand U7893 (N_7893,N_980,N_408);
nor U7894 (N_7894,N_272,N_731);
xor U7895 (N_7895,N_2672,N_1005);
nand U7896 (N_7896,N_753,N_1774);
nor U7897 (N_7897,N_4994,N_2339);
nand U7898 (N_7898,N_2487,N_366);
and U7899 (N_7899,N_1269,N_4972);
xor U7900 (N_7900,N_1282,N_3449);
nand U7901 (N_7901,N_4114,N_1977);
nand U7902 (N_7902,N_3917,N_1398);
nor U7903 (N_7903,N_260,N_3043);
nand U7904 (N_7904,N_3116,N_2366);
and U7905 (N_7905,N_2003,N_746);
xor U7906 (N_7906,N_1738,N_375);
and U7907 (N_7907,N_284,N_2470);
or U7908 (N_7908,N_2240,N_1738);
xnor U7909 (N_7909,N_4384,N_1333);
nor U7910 (N_7910,N_366,N_2083);
and U7911 (N_7911,N_2000,N_3384);
or U7912 (N_7912,N_4102,N_4756);
xor U7913 (N_7913,N_4402,N_3329);
nand U7914 (N_7914,N_2234,N_4545);
and U7915 (N_7915,N_1413,N_2349);
and U7916 (N_7916,N_125,N_1522);
or U7917 (N_7917,N_2965,N_3573);
nor U7918 (N_7918,N_2670,N_849);
nor U7919 (N_7919,N_4886,N_2193);
nand U7920 (N_7920,N_2982,N_1851);
nor U7921 (N_7921,N_4765,N_284);
and U7922 (N_7922,N_4048,N_3170);
and U7923 (N_7923,N_3108,N_3325);
nand U7924 (N_7924,N_2343,N_540);
xnor U7925 (N_7925,N_3721,N_1537);
nand U7926 (N_7926,N_536,N_610);
or U7927 (N_7927,N_1170,N_579);
and U7928 (N_7928,N_2733,N_3302);
nor U7929 (N_7929,N_2216,N_2328);
xnor U7930 (N_7930,N_30,N_4708);
xor U7931 (N_7931,N_4934,N_3800);
nor U7932 (N_7932,N_4753,N_179);
xnor U7933 (N_7933,N_2997,N_2462);
or U7934 (N_7934,N_3416,N_335);
nand U7935 (N_7935,N_4532,N_2734);
nor U7936 (N_7936,N_2525,N_483);
and U7937 (N_7937,N_3275,N_516);
nand U7938 (N_7938,N_3,N_3245);
xor U7939 (N_7939,N_3470,N_1543);
or U7940 (N_7940,N_3180,N_3182);
xor U7941 (N_7941,N_4733,N_2877);
and U7942 (N_7942,N_3881,N_4012);
and U7943 (N_7943,N_1393,N_2937);
nand U7944 (N_7944,N_3078,N_3191);
xor U7945 (N_7945,N_91,N_4478);
or U7946 (N_7946,N_2947,N_1214);
xor U7947 (N_7947,N_3106,N_961);
nand U7948 (N_7948,N_4633,N_234);
and U7949 (N_7949,N_1488,N_4418);
or U7950 (N_7950,N_1657,N_4757);
nand U7951 (N_7951,N_4300,N_238);
nor U7952 (N_7952,N_2282,N_4438);
and U7953 (N_7953,N_966,N_3666);
or U7954 (N_7954,N_1034,N_3192);
nor U7955 (N_7955,N_2931,N_1832);
nor U7956 (N_7956,N_1563,N_1634);
nand U7957 (N_7957,N_4729,N_237);
nand U7958 (N_7958,N_1599,N_3260);
xor U7959 (N_7959,N_2920,N_563);
or U7960 (N_7960,N_3935,N_4300);
xnor U7961 (N_7961,N_3131,N_4639);
or U7962 (N_7962,N_2426,N_1450);
nand U7963 (N_7963,N_3665,N_4626);
nand U7964 (N_7964,N_694,N_4074);
and U7965 (N_7965,N_561,N_3131);
and U7966 (N_7966,N_3807,N_1669);
or U7967 (N_7967,N_4908,N_2157);
or U7968 (N_7968,N_4269,N_327);
nand U7969 (N_7969,N_3803,N_4106);
and U7970 (N_7970,N_3143,N_3289);
nand U7971 (N_7971,N_1730,N_1829);
nor U7972 (N_7972,N_2803,N_2785);
nand U7973 (N_7973,N_4606,N_2668);
and U7974 (N_7974,N_3937,N_618);
nand U7975 (N_7975,N_2206,N_4760);
xor U7976 (N_7976,N_1986,N_1008);
or U7977 (N_7977,N_2222,N_3573);
xnor U7978 (N_7978,N_4581,N_3775);
or U7979 (N_7979,N_1754,N_679);
or U7980 (N_7980,N_4117,N_4336);
xor U7981 (N_7981,N_3755,N_726);
and U7982 (N_7982,N_4063,N_4216);
or U7983 (N_7983,N_1532,N_1817);
and U7984 (N_7984,N_2406,N_2144);
nor U7985 (N_7985,N_4066,N_2039);
and U7986 (N_7986,N_1848,N_653);
nor U7987 (N_7987,N_2541,N_4048);
or U7988 (N_7988,N_2903,N_1253);
nand U7989 (N_7989,N_3344,N_2366);
nand U7990 (N_7990,N_205,N_573);
nand U7991 (N_7991,N_3088,N_3530);
xor U7992 (N_7992,N_4624,N_4173);
and U7993 (N_7993,N_4869,N_640);
and U7994 (N_7994,N_4086,N_2720);
and U7995 (N_7995,N_795,N_339);
xor U7996 (N_7996,N_2378,N_912);
or U7997 (N_7997,N_373,N_145);
nor U7998 (N_7998,N_1346,N_1640);
xor U7999 (N_7999,N_2218,N_1298);
xor U8000 (N_8000,N_4967,N_4668);
or U8001 (N_8001,N_4770,N_4649);
or U8002 (N_8002,N_4926,N_363);
xor U8003 (N_8003,N_350,N_37);
nor U8004 (N_8004,N_1740,N_1562);
xnor U8005 (N_8005,N_459,N_4116);
nand U8006 (N_8006,N_2965,N_4828);
nor U8007 (N_8007,N_3181,N_4985);
or U8008 (N_8008,N_3051,N_1803);
or U8009 (N_8009,N_3371,N_4629);
xor U8010 (N_8010,N_425,N_886);
nor U8011 (N_8011,N_3425,N_184);
xor U8012 (N_8012,N_389,N_956);
nor U8013 (N_8013,N_4731,N_1393);
nor U8014 (N_8014,N_2905,N_2559);
and U8015 (N_8015,N_1458,N_2973);
and U8016 (N_8016,N_4948,N_518);
and U8017 (N_8017,N_2129,N_2959);
xnor U8018 (N_8018,N_4733,N_577);
nand U8019 (N_8019,N_2441,N_2894);
nor U8020 (N_8020,N_1310,N_4665);
xnor U8021 (N_8021,N_504,N_4802);
or U8022 (N_8022,N_27,N_4612);
xor U8023 (N_8023,N_922,N_2179);
nor U8024 (N_8024,N_3924,N_3760);
nor U8025 (N_8025,N_4848,N_4447);
or U8026 (N_8026,N_1941,N_4690);
and U8027 (N_8027,N_4173,N_3348);
nand U8028 (N_8028,N_4086,N_4188);
xnor U8029 (N_8029,N_2289,N_1115);
xor U8030 (N_8030,N_222,N_1103);
or U8031 (N_8031,N_2106,N_479);
xor U8032 (N_8032,N_3265,N_88);
nand U8033 (N_8033,N_3718,N_2050);
and U8034 (N_8034,N_829,N_1146);
nor U8035 (N_8035,N_2511,N_1409);
or U8036 (N_8036,N_822,N_1627);
xnor U8037 (N_8037,N_3058,N_1450);
xor U8038 (N_8038,N_528,N_2385);
and U8039 (N_8039,N_1374,N_4196);
xnor U8040 (N_8040,N_3170,N_3561);
or U8041 (N_8041,N_2082,N_3446);
nand U8042 (N_8042,N_1308,N_4747);
nand U8043 (N_8043,N_1561,N_4551);
and U8044 (N_8044,N_3058,N_1737);
nor U8045 (N_8045,N_4704,N_949);
xnor U8046 (N_8046,N_3593,N_974);
and U8047 (N_8047,N_3830,N_1788);
xnor U8048 (N_8048,N_812,N_3816);
or U8049 (N_8049,N_4274,N_489);
or U8050 (N_8050,N_3677,N_3320);
or U8051 (N_8051,N_1035,N_313);
nand U8052 (N_8052,N_1792,N_2190);
nor U8053 (N_8053,N_263,N_1544);
and U8054 (N_8054,N_4864,N_1955);
nand U8055 (N_8055,N_108,N_3276);
or U8056 (N_8056,N_1233,N_1398);
nand U8057 (N_8057,N_782,N_2939);
xnor U8058 (N_8058,N_2223,N_2778);
or U8059 (N_8059,N_316,N_51);
nor U8060 (N_8060,N_1705,N_714);
or U8061 (N_8061,N_3682,N_4635);
xor U8062 (N_8062,N_1979,N_616);
nor U8063 (N_8063,N_487,N_3319);
xor U8064 (N_8064,N_1936,N_2147);
xnor U8065 (N_8065,N_300,N_804);
nand U8066 (N_8066,N_4191,N_1031);
nor U8067 (N_8067,N_2968,N_758);
and U8068 (N_8068,N_4756,N_1069);
xnor U8069 (N_8069,N_126,N_4473);
nor U8070 (N_8070,N_40,N_194);
and U8071 (N_8071,N_2878,N_4688);
xor U8072 (N_8072,N_4069,N_4885);
or U8073 (N_8073,N_2187,N_4815);
xor U8074 (N_8074,N_496,N_2777);
nor U8075 (N_8075,N_220,N_621);
nor U8076 (N_8076,N_797,N_2896);
nand U8077 (N_8077,N_875,N_4103);
and U8078 (N_8078,N_4746,N_3072);
xor U8079 (N_8079,N_3990,N_2773);
nand U8080 (N_8080,N_2139,N_3589);
nor U8081 (N_8081,N_808,N_4355);
nand U8082 (N_8082,N_4669,N_206);
and U8083 (N_8083,N_1389,N_4307);
xor U8084 (N_8084,N_1263,N_3134);
nand U8085 (N_8085,N_3665,N_111);
nor U8086 (N_8086,N_3684,N_4924);
xnor U8087 (N_8087,N_2958,N_2979);
and U8088 (N_8088,N_2625,N_807);
nor U8089 (N_8089,N_2034,N_3445);
nand U8090 (N_8090,N_4279,N_2088);
nor U8091 (N_8091,N_4439,N_3420);
and U8092 (N_8092,N_437,N_1239);
xor U8093 (N_8093,N_3435,N_2259);
nor U8094 (N_8094,N_795,N_1838);
nand U8095 (N_8095,N_4519,N_570);
and U8096 (N_8096,N_1650,N_3193);
xor U8097 (N_8097,N_283,N_3450);
and U8098 (N_8098,N_4296,N_4394);
nand U8099 (N_8099,N_1100,N_4092);
and U8100 (N_8100,N_1317,N_2639);
nor U8101 (N_8101,N_3016,N_1359);
xor U8102 (N_8102,N_2115,N_23);
and U8103 (N_8103,N_3975,N_552);
nand U8104 (N_8104,N_4708,N_3090);
nand U8105 (N_8105,N_1576,N_321);
and U8106 (N_8106,N_3050,N_270);
nand U8107 (N_8107,N_3604,N_2145);
nand U8108 (N_8108,N_1914,N_4312);
nand U8109 (N_8109,N_730,N_3997);
xor U8110 (N_8110,N_3780,N_1880);
nand U8111 (N_8111,N_99,N_1402);
and U8112 (N_8112,N_4136,N_4816);
xor U8113 (N_8113,N_1660,N_1757);
nor U8114 (N_8114,N_489,N_2400);
xor U8115 (N_8115,N_4265,N_1170);
nand U8116 (N_8116,N_2850,N_1247);
xor U8117 (N_8117,N_4267,N_2221);
xnor U8118 (N_8118,N_533,N_2115);
nor U8119 (N_8119,N_1435,N_2990);
xnor U8120 (N_8120,N_4065,N_753);
or U8121 (N_8121,N_1712,N_4399);
nand U8122 (N_8122,N_194,N_4055);
or U8123 (N_8123,N_1184,N_444);
or U8124 (N_8124,N_3672,N_3750);
nor U8125 (N_8125,N_4309,N_4185);
or U8126 (N_8126,N_4586,N_589);
or U8127 (N_8127,N_3463,N_963);
or U8128 (N_8128,N_3072,N_1519);
nand U8129 (N_8129,N_3463,N_2621);
nor U8130 (N_8130,N_1706,N_2463);
or U8131 (N_8131,N_1191,N_3236);
and U8132 (N_8132,N_4373,N_542);
nand U8133 (N_8133,N_3741,N_1181);
nor U8134 (N_8134,N_4839,N_3158);
or U8135 (N_8135,N_446,N_3688);
nand U8136 (N_8136,N_4852,N_1693);
nor U8137 (N_8137,N_2428,N_4588);
nand U8138 (N_8138,N_1668,N_3938);
nand U8139 (N_8139,N_1864,N_441);
and U8140 (N_8140,N_2203,N_853);
and U8141 (N_8141,N_3450,N_4279);
or U8142 (N_8142,N_664,N_4427);
and U8143 (N_8143,N_3268,N_3043);
nor U8144 (N_8144,N_3225,N_1330);
nor U8145 (N_8145,N_1226,N_4675);
xnor U8146 (N_8146,N_4501,N_4913);
nor U8147 (N_8147,N_4092,N_3034);
xor U8148 (N_8148,N_837,N_453);
or U8149 (N_8149,N_2569,N_1033);
nor U8150 (N_8150,N_1188,N_668);
xnor U8151 (N_8151,N_466,N_4484);
nor U8152 (N_8152,N_397,N_1000);
xor U8153 (N_8153,N_545,N_637);
and U8154 (N_8154,N_2743,N_1005);
xor U8155 (N_8155,N_3989,N_687);
and U8156 (N_8156,N_120,N_1048);
xor U8157 (N_8157,N_1562,N_450);
xnor U8158 (N_8158,N_1482,N_2016);
xor U8159 (N_8159,N_346,N_4489);
xnor U8160 (N_8160,N_3047,N_2998);
or U8161 (N_8161,N_3582,N_268);
or U8162 (N_8162,N_4719,N_1629);
or U8163 (N_8163,N_4933,N_988);
and U8164 (N_8164,N_2799,N_1940);
or U8165 (N_8165,N_191,N_3138);
nand U8166 (N_8166,N_4277,N_4172);
and U8167 (N_8167,N_1691,N_4564);
or U8168 (N_8168,N_2855,N_2676);
nand U8169 (N_8169,N_4142,N_4806);
xor U8170 (N_8170,N_466,N_1432);
and U8171 (N_8171,N_4761,N_1889);
nor U8172 (N_8172,N_467,N_2626);
nor U8173 (N_8173,N_1629,N_4768);
xor U8174 (N_8174,N_1281,N_2800);
xor U8175 (N_8175,N_4197,N_1044);
nand U8176 (N_8176,N_2788,N_2265);
or U8177 (N_8177,N_1920,N_4102);
or U8178 (N_8178,N_3055,N_3504);
nor U8179 (N_8179,N_4696,N_3004);
and U8180 (N_8180,N_3166,N_996);
and U8181 (N_8181,N_78,N_820);
xor U8182 (N_8182,N_771,N_3366);
or U8183 (N_8183,N_1590,N_3334);
nor U8184 (N_8184,N_3237,N_2411);
nand U8185 (N_8185,N_4461,N_2843);
and U8186 (N_8186,N_3610,N_752);
or U8187 (N_8187,N_4599,N_215);
nand U8188 (N_8188,N_3789,N_756);
nor U8189 (N_8189,N_2570,N_4724);
xor U8190 (N_8190,N_3548,N_3612);
nand U8191 (N_8191,N_3904,N_547);
nand U8192 (N_8192,N_1448,N_4662);
nor U8193 (N_8193,N_3930,N_3264);
and U8194 (N_8194,N_3828,N_1672);
and U8195 (N_8195,N_2453,N_714);
nor U8196 (N_8196,N_2873,N_4460);
or U8197 (N_8197,N_1435,N_3791);
or U8198 (N_8198,N_3287,N_503);
nand U8199 (N_8199,N_1392,N_4183);
or U8200 (N_8200,N_3946,N_4592);
and U8201 (N_8201,N_239,N_2414);
nor U8202 (N_8202,N_499,N_2736);
xnor U8203 (N_8203,N_134,N_402);
xor U8204 (N_8204,N_2011,N_3930);
nor U8205 (N_8205,N_4403,N_4627);
and U8206 (N_8206,N_930,N_2381);
and U8207 (N_8207,N_2676,N_1126);
xor U8208 (N_8208,N_783,N_2006);
or U8209 (N_8209,N_1130,N_3737);
xor U8210 (N_8210,N_2608,N_3168);
nand U8211 (N_8211,N_62,N_1717);
nand U8212 (N_8212,N_985,N_105);
nand U8213 (N_8213,N_2320,N_2696);
and U8214 (N_8214,N_1944,N_196);
nor U8215 (N_8215,N_3318,N_4378);
nor U8216 (N_8216,N_948,N_1885);
or U8217 (N_8217,N_3595,N_4863);
xnor U8218 (N_8218,N_4749,N_298);
and U8219 (N_8219,N_4113,N_1118);
and U8220 (N_8220,N_4167,N_4061);
xnor U8221 (N_8221,N_1373,N_4288);
and U8222 (N_8222,N_4276,N_4041);
nor U8223 (N_8223,N_237,N_4792);
xnor U8224 (N_8224,N_918,N_4443);
xor U8225 (N_8225,N_1566,N_1163);
or U8226 (N_8226,N_239,N_971);
nor U8227 (N_8227,N_1652,N_183);
xnor U8228 (N_8228,N_4332,N_780);
or U8229 (N_8229,N_732,N_2831);
xnor U8230 (N_8230,N_4349,N_3885);
xor U8231 (N_8231,N_4659,N_4587);
nor U8232 (N_8232,N_2985,N_2668);
nand U8233 (N_8233,N_4231,N_3132);
nand U8234 (N_8234,N_1952,N_3668);
nor U8235 (N_8235,N_4887,N_4102);
xnor U8236 (N_8236,N_175,N_3474);
xnor U8237 (N_8237,N_2283,N_3344);
nor U8238 (N_8238,N_2809,N_2646);
xnor U8239 (N_8239,N_1290,N_4389);
xor U8240 (N_8240,N_1349,N_3692);
nor U8241 (N_8241,N_1880,N_829);
nand U8242 (N_8242,N_4888,N_4969);
or U8243 (N_8243,N_746,N_4326);
or U8244 (N_8244,N_686,N_4254);
and U8245 (N_8245,N_4987,N_3360);
nand U8246 (N_8246,N_3509,N_2143);
xnor U8247 (N_8247,N_2016,N_4094);
or U8248 (N_8248,N_4477,N_2218);
nand U8249 (N_8249,N_3258,N_2188);
xnor U8250 (N_8250,N_3930,N_3219);
nor U8251 (N_8251,N_1999,N_16);
xor U8252 (N_8252,N_1076,N_4326);
nor U8253 (N_8253,N_3207,N_4400);
and U8254 (N_8254,N_2672,N_4580);
xor U8255 (N_8255,N_4798,N_2600);
and U8256 (N_8256,N_504,N_3428);
xnor U8257 (N_8257,N_959,N_231);
or U8258 (N_8258,N_3568,N_484);
xnor U8259 (N_8259,N_2352,N_1507);
and U8260 (N_8260,N_1707,N_895);
xnor U8261 (N_8261,N_431,N_3603);
nand U8262 (N_8262,N_238,N_1068);
nand U8263 (N_8263,N_2352,N_2619);
nand U8264 (N_8264,N_2152,N_2590);
and U8265 (N_8265,N_3692,N_570);
nand U8266 (N_8266,N_330,N_3989);
nand U8267 (N_8267,N_457,N_3346);
nand U8268 (N_8268,N_983,N_4712);
or U8269 (N_8269,N_3029,N_1207);
or U8270 (N_8270,N_1082,N_3216);
and U8271 (N_8271,N_1966,N_1073);
or U8272 (N_8272,N_2445,N_4669);
nand U8273 (N_8273,N_4477,N_704);
nand U8274 (N_8274,N_4881,N_2965);
xor U8275 (N_8275,N_4773,N_2440);
xnor U8276 (N_8276,N_4241,N_876);
nand U8277 (N_8277,N_2432,N_1352);
or U8278 (N_8278,N_4223,N_3355);
xor U8279 (N_8279,N_32,N_3170);
and U8280 (N_8280,N_4300,N_1349);
nor U8281 (N_8281,N_4306,N_2704);
xnor U8282 (N_8282,N_12,N_278);
nor U8283 (N_8283,N_3326,N_3501);
xnor U8284 (N_8284,N_548,N_1083);
nand U8285 (N_8285,N_2047,N_4924);
nor U8286 (N_8286,N_3769,N_2148);
and U8287 (N_8287,N_4858,N_4427);
or U8288 (N_8288,N_3801,N_3211);
nand U8289 (N_8289,N_903,N_514);
nor U8290 (N_8290,N_1466,N_2176);
or U8291 (N_8291,N_4644,N_1686);
xor U8292 (N_8292,N_141,N_3397);
and U8293 (N_8293,N_3136,N_4297);
or U8294 (N_8294,N_3702,N_2925);
xnor U8295 (N_8295,N_1138,N_334);
and U8296 (N_8296,N_2723,N_3365);
xnor U8297 (N_8297,N_4469,N_4015);
or U8298 (N_8298,N_2907,N_1874);
nor U8299 (N_8299,N_123,N_2569);
xor U8300 (N_8300,N_4783,N_4125);
nand U8301 (N_8301,N_2182,N_3417);
and U8302 (N_8302,N_4218,N_4900);
nand U8303 (N_8303,N_1795,N_2420);
nand U8304 (N_8304,N_2135,N_1342);
or U8305 (N_8305,N_2099,N_1336);
nand U8306 (N_8306,N_3127,N_2650);
xor U8307 (N_8307,N_940,N_256);
xor U8308 (N_8308,N_4228,N_1033);
or U8309 (N_8309,N_2333,N_3398);
nand U8310 (N_8310,N_1014,N_537);
nor U8311 (N_8311,N_1396,N_4227);
nand U8312 (N_8312,N_1161,N_4831);
nor U8313 (N_8313,N_71,N_4768);
xnor U8314 (N_8314,N_2907,N_3340);
xnor U8315 (N_8315,N_652,N_290);
xnor U8316 (N_8316,N_3464,N_2161);
nand U8317 (N_8317,N_1819,N_3060);
or U8318 (N_8318,N_3649,N_2774);
nand U8319 (N_8319,N_3812,N_3955);
nand U8320 (N_8320,N_1003,N_2997);
xor U8321 (N_8321,N_984,N_3183);
nor U8322 (N_8322,N_2652,N_158);
and U8323 (N_8323,N_893,N_3887);
nor U8324 (N_8324,N_1527,N_2726);
nor U8325 (N_8325,N_2386,N_1795);
and U8326 (N_8326,N_2095,N_1046);
and U8327 (N_8327,N_1189,N_1143);
xor U8328 (N_8328,N_4937,N_4497);
nor U8329 (N_8329,N_4822,N_4291);
xor U8330 (N_8330,N_1769,N_4988);
xnor U8331 (N_8331,N_3463,N_2932);
nor U8332 (N_8332,N_2718,N_3302);
xnor U8333 (N_8333,N_4649,N_762);
nor U8334 (N_8334,N_3463,N_803);
and U8335 (N_8335,N_4663,N_4579);
nand U8336 (N_8336,N_1787,N_3127);
and U8337 (N_8337,N_3972,N_1871);
nand U8338 (N_8338,N_4762,N_3571);
and U8339 (N_8339,N_583,N_914);
or U8340 (N_8340,N_3149,N_1912);
and U8341 (N_8341,N_3056,N_2756);
xor U8342 (N_8342,N_1720,N_1612);
or U8343 (N_8343,N_4085,N_3789);
or U8344 (N_8344,N_3820,N_4180);
or U8345 (N_8345,N_3121,N_4668);
xnor U8346 (N_8346,N_1282,N_3223);
nand U8347 (N_8347,N_4958,N_4763);
nor U8348 (N_8348,N_3233,N_2500);
and U8349 (N_8349,N_1979,N_3422);
or U8350 (N_8350,N_3178,N_3691);
xor U8351 (N_8351,N_660,N_185);
xnor U8352 (N_8352,N_2173,N_3433);
and U8353 (N_8353,N_3182,N_4908);
and U8354 (N_8354,N_2759,N_1510);
xnor U8355 (N_8355,N_939,N_3252);
xnor U8356 (N_8356,N_359,N_4371);
or U8357 (N_8357,N_4407,N_3154);
nand U8358 (N_8358,N_1719,N_790);
xor U8359 (N_8359,N_4446,N_3472);
nand U8360 (N_8360,N_4061,N_693);
nor U8361 (N_8361,N_3016,N_3690);
nor U8362 (N_8362,N_3515,N_3864);
nand U8363 (N_8363,N_4126,N_3279);
nand U8364 (N_8364,N_1638,N_504);
nor U8365 (N_8365,N_2700,N_2213);
nand U8366 (N_8366,N_3322,N_2385);
and U8367 (N_8367,N_1145,N_313);
nor U8368 (N_8368,N_3611,N_808);
and U8369 (N_8369,N_2300,N_2531);
or U8370 (N_8370,N_4548,N_1326);
nand U8371 (N_8371,N_149,N_3936);
xnor U8372 (N_8372,N_1151,N_2965);
xor U8373 (N_8373,N_1327,N_2748);
xnor U8374 (N_8374,N_1725,N_4645);
or U8375 (N_8375,N_3176,N_3768);
xor U8376 (N_8376,N_647,N_3309);
nand U8377 (N_8377,N_573,N_753);
xnor U8378 (N_8378,N_2094,N_315);
or U8379 (N_8379,N_530,N_1839);
nand U8380 (N_8380,N_4362,N_4862);
or U8381 (N_8381,N_4406,N_1470);
nand U8382 (N_8382,N_3260,N_4800);
xnor U8383 (N_8383,N_4646,N_4722);
xor U8384 (N_8384,N_2282,N_3953);
or U8385 (N_8385,N_1980,N_4527);
or U8386 (N_8386,N_1163,N_4877);
nor U8387 (N_8387,N_1805,N_4463);
xnor U8388 (N_8388,N_4996,N_2144);
nor U8389 (N_8389,N_1800,N_2186);
nor U8390 (N_8390,N_4395,N_257);
or U8391 (N_8391,N_3765,N_3483);
xnor U8392 (N_8392,N_965,N_3276);
or U8393 (N_8393,N_4949,N_4513);
nor U8394 (N_8394,N_3494,N_4795);
nand U8395 (N_8395,N_139,N_1894);
nor U8396 (N_8396,N_4697,N_2563);
or U8397 (N_8397,N_3860,N_3829);
nand U8398 (N_8398,N_2682,N_4620);
nor U8399 (N_8399,N_3588,N_1715);
nand U8400 (N_8400,N_2249,N_1274);
xor U8401 (N_8401,N_3040,N_2819);
xnor U8402 (N_8402,N_4007,N_1734);
nand U8403 (N_8403,N_3943,N_3550);
nand U8404 (N_8404,N_2104,N_1588);
nand U8405 (N_8405,N_4669,N_4619);
xor U8406 (N_8406,N_1042,N_686);
nand U8407 (N_8407,N_761,N_3127);
or U8408 (N_8408,N_1865,N_3822);
and U8409 (N_8409,N_2117,N_1486);
xnor U8410 (N_8410,N_2520,N_4817);
xor U8411 (N_8411,N_2738,N_2670);
nand U8412 (N_8412,N_691,N_4055);
xnor U8413 (N_8413,N_3300,N_1165);
nor U8414 (N_8414,N_178,N_924);
and U8415 (N_8415,N_4339,N_4372);
nor U8416 (N_8416,N_4161,N_2132);
or U8417 (N_8417,N_4285,N_4807);
or U8418 (N_8418,N_2720,N_791);
nor U8419 (N_8419,N_4958,N_4858);
nand U8420 (N_8420,N_4275,N_3449);
nand U8421 (N_8421,N_2281,N_4512);
and U8422 (N_8422,N_1494,N_65);
or U8423 (N_8423,N_1593,N_4981);
nor U8424 (N_8424,N_1743,N_681);
nor U8425 (N_8425,N_2037,N_3269);
nand U8426 (N_8426,N_1025,N_3089);
nand U8427 (N_8427,N_210,N_3522);
nand U8428 (N_8428,N_1490,N_2067);
and U8429 (N_8429,N_2774,N_4652);
nor U8430 (N_8430,N_1257,N_33);
xnor U8431 (N_8431,N_3334,N_776);
xor U8432 (N_8432,N_2152,N_1283);
or U8433 (N_8433,N_320,N_822);
nand U8434 (N_8434,N_1817,N_842);
xor U8435 (N_8435,N_1701,N_1511);
or U8436 (N_8436,N_2413,N_4776);
nand U8437 (N_8437,N_1904,N_3093);
and U8438 (N_8438,N_1585,N_1350);
xnor U8439 (N_8439,N_1001,N_2184);
or U8440 (N_8440,N_2103,N_1105);
or U8441 (N_8441,N_3822,N_1097);
xnor U8442 (N_8442,N_666,N_2653);
nor U8443 (N_8443,N_2073,N_189);
nor U8444 (N_8444,N_1348,N_3841);
nand U8445 (N_8445,N_3973,N_1940);
xnor U8446 (N_8446,N_3360,N_2442);
xor U8447 (N_8447,N_155,N_490);
nand U8448 (N_8448,N_1615,N_1060);
and U8449 (N_8449,N_3614,N_355);
or U8450 (N_8450,N_4560,N_1929);
nor U8451 (N_8451,N_2113,N_2869);
or U8452 (N_8452,N_3695,N_1215);
xnor U8453 (N_8453,N_1333,N_2164);
and U8454 (N_8454,N_3263,N_2289);
or U8455 (N_8455,N_3616,N_2840);
nand U8456 (N_8456,N_1430,N_416);
nor U8457 (N_8457,N_341,N_1840);
xor U8458 (N_8458,N_4549,N_3476);
nand U8459 (N_8459,N_2801,N_3204);
nand U8460 (N_8460,N_450,N_1296);
and U8461 (N_8461,N_4592,N_2092);
xor U8462 (N_8462,N_4177,N_4305);
nand U8463 (N_8463,N_414,N_48);
or U8464 (N_8464,N_2855,N_1012);
and U8465 (N_8465,N_1847,N_2100);
or U8466 (N_8466,N_3801,N_2200);
nor U8467 (N_8467,N_369,N_4920);
and U8468 (N_8468,N_1585,N_4769);
xnor U8469 (N_8469,N_3149,N_4594);
and U8470 (N_8470,N_3974,N_607);
nand U8471 (N_8471,N_4155,N_772);
nand U8472 (N_8472,N_3508,N_2331);
nand U8473 (N_8473,N_3688,N_734);
xor U8474 (N_8474,N_1143,N_4113);
nand U8475 (N_8475,N_3049,N_1224);
or U8476 (N_8476,N_3022,N_2487);
or U8477 (N_8477,N_2916,N_4827);
nand U8478 (N_8478,N_135,N_3694);
nand U8479 (N_8479,N_3152,N_3196);
nor U8480 (N_8480,N_1169,N_2383);
nor U8481 (N_8481,N_1068,N_2671);
nor U8482 (N_8482,N_4420,N_3170);
and U8483 (N_8483,N_3272,N_1593);
and U8484 (N_8484,N_2051,N_4802);
nor U8485 (N_8485,N_4562,N_265);
and U8486 (N_8486,N_4868,N_1172);
or U8487 (N_8487,N_429,N_4165);
xor U8488 (N_8488,N_2972,N_604);
nor U8489 (N_8489,N_2430,N_4589);
and U8490 (N_8490,N_3062,N_1578);
or U8491 (N_8491,N_1883,N_4457);
and U8492 (N_8492,N_508,N_1245);
nor U8493 (N_8493,N_2908,N_3546);
xor U8494 (N_8494,N_3748,N_1199);
and U8495 (N_8495,N_216,N_865);
and U8496 (N_8496,N_2284,N_645);
xor U8497 (N_8497,N_4070,N_1513);
nand U8498 (N_8498,N_385,N_60);
nor U8499 (N_8499,N_543,N_1330);
xor U8500 (N_8500,N_1359,N_4439);
xor U8501 (N_8501,N_4491,N_840);
or U8502 (N_8502,N_4726,N_2825);
xnor U8503 (N_8503,N_2480,N_4665);
nand U8504 (N_8504,N_4050,N_4747);
and U8505 (N_8505,N_204,N_3767);
nor U8506 (N_8506,N_4311,N_3858);
or U8507 (N_8507,N_1518,N_4651);
nor U8508 (N_8508,N_2941,N_3589);
and U8509 (N_8509,N_3265,N_4205);
or U8510 (N_8510,N_2494,N_519);
nor U8511 (N_8511,N_2159,N_3223);
nor U8512 (N_8512,N_881,N_8);
and U8513 (N_8513,N_2246,N_2770);
xor U8514 (N_8514,N_3334,N_2410);
and U8515 (N_8515,N_238,N_3401);
or U8516 (N_8516,N_709,N_2326);
nor U8517 (N_8517,N_2185,N_115);
xor U8518 (N_8518,N_46,N_4030);
xnor U8519 (N_8519,N_2778,N_3805);
or U8520 (N_8520,N_4289,N_3755);
nor U8521 (N_8521,N_796,N_832);
and U8522 (N_8522,N_820,N_652);
or U8523 (N_8523,N_2653,N_2680);
or U8524 (N_8524,N_4008,N_4678);
or U8525 (N_8525,N_4706,N_350);
nand U8526 (N_8526,N_109,N_426);
and U8527 (N_8527,N_14,N_752);
nand U8528 (N_8528,N_3127,N_4573);
nand U8529 (N_8529,N_1388,N_1507);
and U8530 (N_8530,N_3507,N_321);
nor U8531 (N_8531,N_542,N_4603);
xnor U8532 (N_8532,N_975,N_4274);
or U8533 (N_8533,N_893,N_353);
nor U8534 (N_8534,N_724,N_4112);
nor U8535 (N_8535,N_2046,N_2362);
nand U8536 (N_8536,N_2071,N_2988);
or U8537 (N_8537,N_669,N_701);
or U8538 (N_8538,N_176,N_4584);
xor U8539 (N_8539,N_4471,N_437);
and U8540 (N_8540,N_875,N_3848);
or U8541 (N_8541,N_2887,N_2878);
nand U8542 (N_8542,N_4254,N_3789);
nand U8543 (N_8543,N_4081,N_4817);
nor U8544 (N_8544,N_2161,N_4877);
and U8545 (N_8545,N_4838,N_4320);
and U8546 (N_8546,N_4001,N_307);
xnor U8547 (N_8547,N_3569,N_3424);
and U8548 (N_8548,N_1625,N_1518);
xor U8549 (N_8549,N_4268,N_799);
and U8550 (N_8550,N_2358,N_1851);
xnor U8551 (N_8551,N_4565,N_522);
or U8552 (N_8552,N_4359,N_1698);
or U8553 (N_8553,N_2976,N_616);
xor U8554 (N_8554,N_1080,N_3073);
nor U8555 (N_8555,N_738,N_3459);
or U8556 (N_8556,N_4508,N_3659);
nand U8557 (N_8557,N_4270,N_4972);
nor U8558 (N_8558,N_1581,N_2300);
or U8559 (N_8559,N_2078,N_4814);
nor U8560 (N_8560,N_2600,N_3536);
xor U8561 (N_8561,N_4121,N_4270);
and U8562 (N_8562,N_3967,N_1490);
nor U8563 (N_8563,N_2896,N_4930);
xnor U8564 (N_8564,N_2989,N_1603);
or U8565 (N_8565,N_3963,N_4298);
nor U8566 (N_8566,N_2871,N_1118);
nor U8567 (N_8567,N_3802,N_4486);
or U8568 (N_8568,N_86,N_4705);
xnor U8569 (N_8569,N_3389,N_528);
nand U8570 (N_8570,N_4841,N_2083);
xor U8571 (N_8571,N_2263,N_4300);
or U8572 (N_8572,N_1336,N_1485);
xor U8573 (N_8573,N_3710,N_4588);
nor U8574 (N_8574,N_2208,N_1072);
and U8575 (N_8575,N_1026,N_1314);
nand U8576 (N_8576,N_3552,N_1343);
or U8577 (N_8577,N_2691,N_4125);
nor U8578 (N_8578,N_4073,N_454);
xnor U8579 (N_8579,N_4269,N_4666);
nand U8580 (N_8580,N_862,N_39);
xor U8581 (N_8581,N_393,N_4078);
nor U8582 (N_8582,N_2411,N_535);
or U8583 (N_8583,N_4543,N_3698);
and U8584 (N_8584,N_2373,N_3675);
nor U8585 (N_8585,N_2060,N_240);
or U8586 (N_8586,N_2171,N_4646);
xnor U8587 (N_8587,N_1848,N_2952);
nor U8588 (N_8588,N_745,N_812);
nor U8589 (N_8589,N_4252,N_3057);
xor U8590 (N_8590,N_3544,N_758);
or U8591 (N_8591,N_1046,N_2426);
nand U8592 (N_8592,N_3473,N_2646);
xor U8593 (N_8593,N_329,N_2163);
xor U8594 (N_8594,N_1923,N_1067);
xor U8595 (N_8595,N_3858,N_511);
nor U8596 (N_8596,N_357,N_1768);
nand U8597 (N_8597,N_599,N_308);
nor U8598 (N_8598,N_2421,N_4348);
nand U8599 (N_8599,N_4501,N_1794);
and U8600 (N_8600,N_3359,N_3574);
or U8601 (N_8601,N_4545,N_2098);
nand U8602 (N_8602,N_726,N_29);
nor U8603 (N_8603,N_470,N_1467);
nor U8604 (N_8604,N_696,N_3580);
xnor U8605 (N_8605,N_4998,N_110);
nand U8606 (N_8606,N_3844,N_2764);
and U8607 (N_8607,N_4151,N_3089);
or U8608 (N_8608,N_3240,N_2938);
nand U8609 (N_8609,N_4951,N_4510);
or U8610 (N_8610,N_716,N_1016);
nand U8611 (N_8611,N_2515,N_1342);
and U8612 (N_8612,N_4088,N_4711);
and U8613 (N_8613,N_1245,N_3630);
nor U8614 (N_8614,N_4246,N_439);
xnor U8615 (N_8615,N_3988,N_2861);
nor U8616 (N_8616,N_4100,N_1480);
and U8617 (N_8617,N_959,N_4663);
xnor U8618 (N_8618,N_2663,N_3759);
or U8619 (N_8619,N_383,N_375);
nand U8620 (N_8620,N_2640,N_3129);
xnor U8621 (N_8621,N_228,N_3734);
or U8622 (N_8622,N_2810,N_3496);
nor U8623 (N_8623,N_877,N_274);
or U8624 (N_8624,N_4218,N_781);
and U8625 (N_8625,N_944,N_4167);
or U8626 (N_8626,N_3279,N_4454);
xor U8627 (N_8627,N_3515,N_455);
and U8628 (N_8628,N_4841,N_1735);
nor U8629 (N_8629,N_2597,N_435);
nor U8630 (N_8630,N_223,N_3987);
and U8631 (N_8631,N_1532,N_2786);
xnor U8632 (N_8632,N_1909,N_4806);
nor U8633 (N_8633,N_154,N_3654);
and U8634 (N_8634,N_3826,N_2554);
or U8635 (N_8635,N_3548,N_1782);
nor U8636 (N_8636,N_3077,N_502);
xor U8637 (N_8637,N_1216,N_3972);
or U8638 (N_8638,N_4719,N_1914);
and U8639 (N_8639,N_1732,N_4744);
nor U8640 (N_8640,N_1481,N_1831);
nand U8641 (N_8641,N_1763,N_4590);
nor U8642 (N_8642,N_1602,N_1149);
and U8643 (N_8643,N_4244,N_200);
or U8644 (N_8644,N_107,N_3046);
xnor U8645 (N_8645,N_4362,N_3663);
nand U8646 (N_8646,N_2051,N_4278);
and U8647 (N_8647,N_1595,N_621);
nand U8648 (N_8648,N_2367,N_2480);
and U8649 (N_8649,N_1944,N_1785);
xor U8650 (N_8650,N_4279,N_4822);
nor U8651 (N_8651,N_456,N_2862);
nand U8652 (N_8652,N_2989,N_1181);
nor U8653 (N_8653,N_4153,N_2744);
or U8654 (N_8654,N_737,N_2545);
and U8655 (N_8655,N_399,N_2820);
and U8656 (N_8656,N_88,N_644);
xor U8657 (N_8657,N_1947,N_102);
or U8658 (N_8658,N_4349,N_2288);
or U8659 (N_8659,N_3100,N_164);
nand U8660 (N_8660,N_3613,N_1306);
or U8661 (N_8661,N_3347,N_176);
and U8662 (N_8662,N_1034,N_298);
and U8663 (N_8663,N_4146,N_2169);
nand U8664 (N_8664,N_2773,N_2093);
or U8665 (N_8665,N_1743,N_2136);
or U8666 (N_8666,N_665,N_3833);
xor U8667 (N_8667,N_2618,N_2828);
or U8668 (N_8668,N_490,N_1224);
and U8669 (N_8669,N_918,N_185);
xor U8670 (N_8670,N_250,N_2584);
xor U8671 (N_8671,N_3094,N_2139);
nand U8672 (N_8672,N_1514,N_23);
nor U8673 (N_8673,N_4804,N_1155);
nand U8674 (N_8674,N_2903,N_4961);
or U8675 (N_8675,N_4357,N_333);
xor U8676 (N_8676,N_2728,N_3250);
or U8677 (N_8677,N_4657,N_3592);
nor U8678 (N_8678,N_100,N_4204);
or U8679 (N_8679,N_2251,N_4740);
nor U8680 (N_8680,N_2069,N_4478);
or U8681 (N_8681,N_3175,N_1014);
nor U8682 (N_8682,N_601,N_4966);
or U8683 (N_8683,N_2517,N_2662);
nor U8684 (N_8684,N_548,N_3344);
and U8685 (N_8685,N_347,N_3036);
nor U8686 (N_8686,N_3729,N_676);
xor U8687 (N_8687,N_867,N_1728);
and U8688 (N_8688,N_1519,N_882);
xnor U8689 (N_8689,N_2557,N_2302);
and U8690 (N_8690,N_2856,N_2834);
xnor U8691 (N_8691,N_4656,N_1507);
xor U8692 (N_8692,N_3093,N_131);
or U8693 (N_8693,N_4905,N_4569);
or U8694 (N_8694,N_54,N_4892);
xor U8695 (N_8695,N_2141,N_987);
nor U8696 (N_8696,N_1896,N_1658);
and U8697 (N_8697,N_4893,N_517);
nand U8698 (N_8698,N_2215,N_3581);
or U8699 (N_8699,N_172,N_2263);
or U8700 (N_8700,N_1030,N_756);
and U8701 (N_8701,N_1735,N_285);
or U8702 (N_8702,N_708,N_1316);
nand U8703 (N_8703,N_1263,N_2615);
and U8704 (N_8704,N_2455,N_4071);
and U8705 (N_8705,N_1767,N_3057);
or U8706 (N_8706,N_3756,N_4490);
and U8707 (N_8707,N_592,N_2375);
xor U8708 (N_8708,N_3300,N_1060);
or U8709 (N_8709,N_1300,N_2556);
nand U8710 (N_8710,N_4477,N_3876);
nor U8711 (N_8711,N_3682,N_56);
xor U8712 (N_8712,N_963,N_1300);
xor U8713 (N_8713,N_2107,N_4606);
and U8714 (N_8714,N_4340,N_1038);
nand U8715 (N_8715,N_1283,N_1941);
xnor U8716 (N_8716,N_1540,N_810);
nor U8717 (N_8717,N_2714,N_174);
nor U8718 (N_8718,N_617,N_1171);
or U8719 (N_8719,N_229,N_1689);
or U8720 (N_8720,N_1167,N_287);
or U8721 (N_8721,N_436,N_607);
or U8722 (N_8722,N_330,N_2023);
nor U8723 (N_8723,N_2398,N_2624);
xor U8724 (N_8724,N_275,N_4971);
nor U8725 (N_8725,N_3349,N_333);
or U8726 (N_8726,N_919,N_1632);
and U8727 (N_8727,N_2945,N_3110);
nand U8728 (N_8728,N_4625,N_1532);
nand U8729 (N_8729,N_3765,N_3318);
xnor U8730 (N_8730,N_4318,N_3781);
xor U8731 (N_8731,N_974,N_184);
nor U8732 (N_8732,N_3493,N_2308);
and U8733 (N_8733,N_1287,N_4949);
nor U8734 (N_8734,N_3384,N_1275);
nor U8735 (N_8735,N_1009,N_2796);
and U8736 (N_8736,N_3335,N_2670);
or U8737 (N_8737,N_991,N_371);
or U8738 (N_8738,N_1642,N_3432);
nand U8739 (N_8739,N_633,N_4945);
nor U8740 (N_8740,N_3698,N_4825);
or U8741 (N_8741,N_4200,N_1595);
and U8742 (N_8742,N_1510,N_866);
nand U8743 (N_8743,N_2833,N_2444);
and U8744 (N_8744,N_2560,N_1685);
nand U8745 (N_8745,N_130,N_2574);
or U8746 (N_8746,N_4089,N_342);
or U8747 (N_8747,N_1646,N_601);
or U8748 (N_8748,N_3439,N_1547);
xnor U8749 (N_8749,N_1336,N_2920);
nor U8750 (N_8750,N_869,N_1786);
or U8751 (N_8751,N_1164,N_481);
and U8752 (N_8752,N_4243,N_950);
xor U8753 (N_8753,N_2656,N_4433);
nor U8754 (N_8754,N_375,N_995);
and U8755 (N_8755,N_2491,N_152);
xor U8756 (N_8756,N_4901,N_68);
nand U8757 (N_8757,N_3789,N_2870);
and U8758 (N_8758,N_4520,N_327);
nor U8759 (N_8759,N_167,N_906);
or U8760 (N_8760,N_758,N_2662);
nand U8761 (N_8761,N_1528,N_2107);
nor U8762 (N_8762,N_2743,N_4425);
and U8763 (N_8763,N_2968,N_2451);
and U8764 (N_8764,N_3556,N_2624);
and U8765 (N_8765,N_1676,N_890);
nand U8766 (N_8766,N_1348,N_525);
xor U8767 (N_8767,N_3338,N_2312);
nand U8768 (N_8768,N_4043,N_2360);
nand U8769 (N_8769,N_3015,N_3183);
xor U8770 (N_8770,N_1571,N_1106);
nand U8771 (N_8771,N_1021,N_3410);
nor U8772 (N_8772,N_1203,N_4131);
nor U8773 (N_8773,N_2923,N_4112);
xor U8774 (N_8774,N_4463,N_2294);
xnor U8775 (N_8775,N_3556,N_2671);
nor U8776 (N_8776,N_934,N_1662);
xnor U8777 (N_8777,N_816,N_3144);
nand U8778 (N_8778,N_1008,N_4728);
and U8779 (N_8779,N_394,N_3926);
xor U8780 (N_8780,N_4709,N_4832);
and U8781 (N_8781,N_3072,N_4739);
and U8782 (N_8782,N_2185,N_4792);
nand U8783 (N_8783,N_2101,N_2125);
or U8784 (N_8784,N_3266,N_76);
xor U8785 (N_8785,N_3884,N_4303);
xnor U8786 (N_8786,N_1274,N_4022);
nor U8787 (N_8787,N_4747,N_4426);
or U8788 (N_8788,N_4477,N_1757);
xor U8789 (N_8789,N_4886,N_75);
and U8790 (N_8790,N_1990,N_2139);
nand U8791 (N_8791,N_4714,N_338);
nand U8792 (N_8792,N_4903,N_3531);
xnor U8793 (N_8793,N_3318,N_102);
nor U8794 (N_8794,N_369,N_947);
and U8795 (N_8795,N_97,N_2831);
nand U8796 (N_8796,N_3259,N_246);
or U8797 (N_8797,N_4550,N_2851);
or U8798 (N_8798,N_892,N_4866);
nor U8799 (N_8799,N_3533,N_3034);
or U8800 (N_8800,N_348,N_2736);
xor U8801 (N_8801,N_2478,N_503);
and U8802 (N_8802,N_1455,N_929);
and U8803 (N_8803,N_4363,N_3856);
and U8804 (N_8804,N_3470,N_2196);
xnor U8805 (N_8805,N_2497,N_1258);
nand U8806 (N_8806,N_139,N_131);
xnor U8807 (N_8807,N_3098,N_1037);
and U8808 (N_8808,N_2157,N_772);
nor U8809 (N_8809,N_4211,N_898);
xor U8810 (N_8810,N_4519,N_290);
or U8811 (N_8811,N_3083,N_178);
xnor U8812 (N_8812,N_1118,N_643);
nor U8813 (N_8813,N_3837,N_3692);
nand U8814 (N_8814,N_242,N_3970);
and U8815 (N_8815,N_1759,N_630);
nor U8816 (N_8816,N_3581,N_2736);
nand U8817 (N_8817,N_4952,N_1156);
nand U8818 (N_8818,N_2428,N_4944);
nor U8819 (N_8819,N_158,N_2);
and U8820 (N_8820,N_2354,N_4224);
nor U8821 (N_8821,N_132,N_3526);
nand U8822 (N_8822,N_3092,N_4640);
xor U8823 (N_8823,N_1996,N_4838);
and U8824 (N_8824,N_281,N_2234);
and U8825 (N_8825,N_2510,N_97);
xor U8826 (N_8826,N_199,N_131);
and U8827 (N_8827,N_1168,N_953);
nor U8828 (N_8828,N_4004,N_3225);
nor U8829 (N_8829,N_3137,N_2243);
or U8830 (N_8830,N_1865,N_3516);
nor U8831 (N_8831,N_3773,N_597);
nand U8832 (N_8832,N_4387,N_1614);
nor U8833 (N_8833,N_100,N_981);
nor U8834 (N_8834,N_3423,N_1526);
and U8835 (N_8835,N_1782,N_4402);
nand U8836 (N_8836,N_3022,N_2912);
nand U8837 (N_8837,N_1649,N_3993);
or U8838 (N_8838,N_1681,N_2828);
xor U8839 (N_8839,N_312,N_1093);
or U8840 (N_8840,N_2487,N_2965);
and U8841 (N_8841,N_4917,N_777);
or U8842 (N_8842,N_2699,N_1534);
nor U8843 (N_8843,N_1089,N_2786);
nor U8844 (N_8844,N_336,N_2410);
nor U8845 (N_8845,N_2997,N_196);
and U8846 (N_8846,N_3679,N_245);
nand U8847 (N_8847,N_2694,N_3540);
nand U8848 (N_8848,N_1867,N_3779);
or U8849 (N_8849,N_1465,N_3802);
and U8850 (N_8850,N_2211,N_2653);
nand U8851 (N_8851,N_3868,N_3283);
and U8852 (N_8852,N_261,N_3952);
nor U8853 (N_8853,N_285,N_1049);
and U8854 (N_8854,N_584,N_1178);
and U8855 (N_8855,N_2560,N_2889);
xor U8856 (N_8856,N_4178,N_4245);
or U8857 (N_8857,N_4998,N_4930);
xnor U8858 (N_8858,N_4514,N_3588);
xor U8859 (N_8859,N_663,N_1570);
xor U8860 (N_8860,N_30,N_4304);
xnor U8861 (N_8861,N_621,N_2649);
xor U8862 (N_8862,N_996,N_1392);
and U8863 (N_8863,N_4011,N_1422);
or U8864 (N_8864,N_2559,N_4584);
or U8865 (N_8865,N_412,N_1932);
nand U8866 (N_8866,N_2603,N_4409);
and U8867 (N_8867,N_4303,N_4682);
xor U8868 (N_8868,N_1699,N_1206);
nand U8869 (N_8869,N_94,N_3299);
xnor U8870 (N_8870,N_2887,N_4341);
nor U8871 (N_8871,N_3000,N_591);
nand U8872 (N_8872,N_1708,N_1242);
nor U8873 (N_8873,N_4125,N_3517);
nand U8874 (N_8874,N_4607,N_1766);
or U8875 (N_8875,N_2126,N_3324);
nand U8876 (N_8876,N_3320,N_3054);
xnor U8877 (N_8877,N_1785,N_4213);
or U8878 (N_8878,N_2883,N_997);
and U8879 (N_8879,N_3989,N_3951);
or U8880 (N_8880,N_760,N_3414);
xor U8881 (N_8881,N_216,N_4782);
or U8882 (N_8882,N_3021,N_623);
nor U8883 (N_8883,N_1886,N_0);
or U8884 (N_8884,N_3862,N_400);
and U8885 (N_8885,N_335,N_3783);
xnor U8886 (N_8886,N_2216,N_1000);
nand U8887 (N_8887,N_2673,N_4064);
and U8888 (N_8888,N_1546,N_2255);
and U8889 (N_8889,N_4515,N_441);
nand U8890 (N_8890,N_167,N_4824);
nand U8891 (N_8891,N_3368,N_1209);
nor U8892 (N_8892,N_1504,N_2535);
nor U8893 (N_8893,N_739,N_1385);
nand U8894 (N_8894,N_168,N_2481);
xor U8895 (N_8895,N_4670,N_1852);
or U8896 (N_8896,N_2520,N_1851);
nand U8897 (N_8897,N_3334,N_1609);
nor U8898 (N_8898,N_200,N_2411);
or U8899 (N_8899,N_3562,N_3305);
xor U8900 (N_8900,N_3806,N_1687);
nor U8901 (N_8901,N_4841,N_3507);
nand U8902 (N_8902,N_4638,N_2166);
xor U8903 (N_8903,N_1101,N_3790);
or U8904 (N_8904,N_773,N_3947);
or U8905 (N_8905,N_1408,N_100);
nand U8906 (N_8906,N_4565,N_2616);
xnor U8907 (N_8907,N_235,N_4461);
nor U8908 (N_8908,N_1014,N_3273);
and U8909 (N_8909,N_915,N_1846);
nand U8910 (N_8910,N_3454,N_2207);
nor U8911 (N_8911,N_1172,N_723);
nor U8912 (N_8912,N_3330,N_4804);
nor U8913 (N_8913,N_1829,N_390);
nor U8914 (N_8914,N_4807,N_1396);
nor U8915 (N_8915,N_1876,N_2832);
nand U8916 (N_8916,N_2320,N_2190);
nor U8917 (N_8917,N_492,N_4521);
xnor U8918 (N_8918,N_1840,N_548);
or U8919 (N_8919,N_4975,N_1553);
nor U8920 (N_8920,N_3775,N_1146);
nor U8921 (N_8921,N_63,N_200);
and U8922 (N_8922,N_3479,N_3977);
and U8923 (N_8923,N_796,N_4118);
nand U8924 (N_8924,N_2642,N_2139);
xor U8925 (N_8925,N_1140,N_3478);
and U8926 (N_8926,N_4762,N_4735);
xnor U8927 (N_8927,N_1806,N_326);
and U8928 (N_8928,N_3411,N_1671);
nand U8929 (N_8929,N_2099,N_3645);
xor U8930 (N_8930,N_373,N_4620);
or U8931 (N_8931,N_572,N_4162);
nor U8932 (N_8932,N_4299,N_4120);
nor U8933 (N_8933,N_3737,N_3465);
xnor U8934 (N_8934,N_1439,N_3940);
or U8935 (N_8935,N_1254,N_4746);
or U8936 (N_8936,N_4009,N_4892);
or U8937 (N_8937,N_4186,N_1607);
and U8938 (N_8938,N_344,N_156);
nor U8939 (N_8939,N_3915,N_14);
or U8940 (N_8940,N_4072,N_4619);
or U8941 (N_8941,N_4698,N_2398);
and U8942 (N_8942,N_380,N_4327);
nor U8943 (N_8943,N_1525,N_3252);
and U8944 (N_8944,N_1858,N_508);
xor U8945 (N_8945,N_3677,N_1656);
and U8946 (N_8946,N_2086,N_4050);
or U8947 (N_8947,N_2055,N_2628);
nand U8948 (N_8948,N_417,N_4403);
xnor U8949 (N_8949,N_2598,N_879);
or U8950 (N_8950,N_988,N_4520);
nor U8951 (N_8951,N_520,N_4966);
and U8952 (N_8952,N_547,N_3654);
nand U8953 (N_8953,N_2307,N_243);
xnor U8954 (N_8954,N_2782,N_1553);
nor U8955 (N_8955,N_1866,N_3555);
xnor U8956 (N_8956,N_720,N_1752);
nand U8957 (N_8957,N_4676,N_4446);
nor U8958 (N_8958,N_4915,N_4763);
nor U8959 (N_8959,N_2746,N_4007);
nand U8960 (N_8960,N_3373,N_1829);
and U8961 (N_8961,N_132,N_910);
and U8962 (N_8962,N_1640,N_2181);
or U8963 (N_8963,N_968,N_4191);
nand U8964 (N_8964,N_1164,N_2934);
or U8965 (N_8965,N_364,N_679);
xnor U8966 (N_8966,N_2274,N_2159);
nor U8967 (N_8967,N_900,N_1006);
and U8968 (N_8968,N_906,N_2566);
and U8969 (N_8969,N_4518,N_4469);
or U8970 (N_8970,N_2434,N_3162);
and U8971 (N_8971,N_860,N_1155);
and U8972 (N_8972,N_2688,N_4185);
nand U8973 (N_8973,N_723,N_1154);
and U8974 (N_8974,N_1928,N_3634);
or U8975 (N_8975,N_2463,N_4524);
nor U8976 (N_8976,N_66,N_1154);
or U8977 (N_8977,N_3986,N_3044);
and U8978 (N_8978,N_3739,N_791);
xnor U8979 (N_8979,N_1687,N_553);
nand U8980 (N_8980,N_3611,N_4368);
xor U8981 (N_8981,N_3289,N_2391);
nand U8982 (N_8982,N_134,N_1744);
nor U8983 (N_8983,N_3713,N_1451);
or U8984 (N_8984,N_2056,N_4210);
nand U8985 (N_8985,N_3518,N_424);
nand U8986 (N_8986,N_545,N_4520);
nand U8987 (N_8987,N_959,N_3601);
or U8988 (N_8988,N_1911,N_1921);
and U8989 (N_8989,N_3731,N_508);
nor U8990 (N_8990,N_1137,N_1444);
nor U8991 (N_8991,N_3831,N_3308);
or U8992 (N_8992,N_1281,N_4057);
or U8993 (N_8993,N_3068,N_4184);
xnor U8994 (N_8994,N_3212,N_3572);
or U8995 (N_8995,N_670,N_3886);
nor U8996 (N_8996,N_3722,N_1243);
and U8997 (N_8997,N_1963,N_4111);
nor U8998 (N_8998,N_538,N_815);
nor U8999 (N_8999,N_1824,N_4229);
xor U9000 (N_9000,N_1153,N_4142);
nor U9001 (N_9001,N_73,N_3575);
and U9002 (N_9002,N_6,N_1309);
xnor U9003 (N_9003,N_295,N_3245);
and U9004 (N_9004,N_518,N_2206);
xnor U9005 (N_9005,N_4647,N_1833);
and U9006 (N_9006,N_4165,N_760);
and U9007 (N_9007,N_4600,N_1452);
nand U9008 (N_9008,N_789,N_3004);
and U9009 (N_9009,N_1774,N_830);
or U9010 (N_9010,N_3753,N_391);
nand U9011 (N_9011,N_486,N_1673);
nor U9012 (N_9012,N_3490,N_2654);
and U9013 (N_9013,N_2600,N_2570);
nand U9014 (N_9014,N_544,N_2552);
xor U9015 (N_9015,N_771,N_79);
or U9016 (N_9016,N_3573,N_2926);
nor U9017 (N_9017,N_1649,N_4103);
and U9018 (N_9018,N_4728,N_1050);
nand U9019 (N_9019,N_3098,N_3551);
and U9020 (N_9020,N_3359,N_1099);
and U9021 (N_9021,N_1270,N_4632);
or U9022 (N_9022,N_2584,N_1795);
and U9023 (N_9023,N_2225,N_892);
or U9024 (N_9024,N_2982,N_3737);
and U9025 (N_9025,N_4536,N_2777);
nor U9026 (N_9026,N_4131,N_1583);
nand U9027 (N_9027,N_4481,N_4598);
xor U9028 (N_9028,N_526,N_3);
nor U9029 (N_9029,N_1227,N_4186);
nand U9030 (N_9030,N_978,N_4025);
nand U9031 (N_9031,N_1747,N_3327);
and U9032 (N_9032,N_2960,N_1496);
or U9033 (N_9033,N_2945,N_988);
or U9034 (N_9034,N_855,N_2382);
nand U9035 (N_9035,N_1337,N_4094);
xnor U9036 (N_9036,N_356,N_3208);
and U9037 (N_9037,N_2817,N_2961);
or U9038 (N_9038,N_4084,N_1184);
and U9039 (N_9039,N_1143,N_2632);
and U9040 (N_9040,N_1436,N_92);
or U9041 (N_9041,N_2409,N_2628);
xnor U9042 (N_9042,N_886,N_645);
or U9043 (N_9043,N_3813,N_426);
nor U9044 (N_9044,N_1569,N_3128);
nor U9045 (N_9045,N_2143,N_2934);
and U9046 (N_9046,N_2562,N_1991);
or U9047 (N_9047,N_2264,N_242);
and U9048 (N_9048,N_4609,N_2595);
xnor U9049 (N_9049,N_1002,N_638);
or U9050 (N_9050,N_645,N_545);
or U9051 (N_9051,N_4223,N_3789);
xor U9052 (N_9052,N_3122,N_2704);
and U9053 (N_9053,N_975,N_202);
or U9054 (N_9054,N_4660,N_801);
or U9055 (N_9055,N_839,N_299);
xnor U9056 (N_9056,N_885,N_15);
nand U9057 (N_9057,N_3221,N_1307);
nand U9058 (N_9058,N_2961,N_3023);
and U9059 (N_9059,N_1665,N_3834);
nand U9060 (N_9060,N_1802,N_437);
and U9061 (N_9061,N_2223,N_3552);
nand U9062 (N_9062,N_101,N_4265);
and U9063 (N_9063,N_4465,N_1708);
xnor U9064 (N_9064,N_1059,N_3842);
nand U9065 (N_9065,N_4182,N_3384);
or U9066 (N_9066,N_4314,N_4770);
xor U9067 (N_9067,N_929,N_2686);
nand U9068 (N_9068,N_939,N_2449);
nand U9069 (N_9069,N_3344,N_770);
nor U9070 (N_9070,N_1257,N_919);
nor U9071 (N_9071,N_387,N_221);
nor U9072 (N_9072,N_4997,N_2897);
and U9073 (N_9073,N_3909,N_2713);
and U9074 (N_9074,N_1931,N_95);
nor U9075 (N_9075,N_1261,N_1850);
and U9076 (N_9076,N_1171,N_2783);
nor U9077 (N_9077,N_1876,N_848);
xor U9078 (N_9078,N_3060,N_2432);
xor U9079 (N_9079,N_1472,N_1401);
nor U9080 (N_9080,N_4413,N_4877);
nor U9081 (N_9081,N_1295,N_3321);
or U9082 (N_9082,N_385,N_2288);
and U9083 (N_9083,N_2000,N_4240);
and U9084 (N_9084,N_3327,N_483);
nand U9085 (N_9085,N_3141,N_4514);
nor U9086 (N_9086,N_3379,N_20);
nor U9087 (N_9087,N_1896,N_1144);
and U9088 (N_9088,N_903,N_273);
xor U9089 (N_9089,N_208,N_55);
nand U9090 (N_9090,N_2860,N_2956);
and U9091 (N_9091,N_60,N_3059);
or U9092 (N_9092,N_1803,N_22);
and U9093 (N_9093,N_2941,N_4608);
xor U9094 (N_9094,N_2365,N_3706);
nand U9095 (N_9095,N_4718,N_2127);
and U9096 (N_9096,N_3623,N_3551);
xor U9097 (N_9097,N_1426,N_4880);
and U9098 (N_9098,N_2014,N_4551);
or U9099 (N_9099,N_3638,N_558);
nand U9100 (N_9100,N_3207,N_3092);
nor U9101 (N_9101,N_1231,N_3500);
or U9102 (N_9102,N_4566,N_4712);
or U9103 (N_9103,N_2301,N_2613);
and U9104 (N_9104,N_952,N_4903);
and U9105 (N_9105,N_4403,N_3264);
nor U9106 (N_9106,N_1373,N_2530);
nand U9107 (N_9107,N_1102,N_2345);
nor U9108 (N_9108,N_3329,N_2050);
or U9109 (N_9109,N_1342,N_4215);
xnor U9110 (N_9110,N_2332,N_830);
nand U9111 (N_9111,N_4659,N_2367);
nand U9112 (N_9112,N_4302,N_4667);
or U9113 (N_9113,N_4282,N_888);
nor U9114 (N_9114,N_772,N_228);
or U9115 (N_9115,N_2895,N_3028);
and U9116 (N_9116,N_833,N_84);
or U9117 (N_9117,N_1368,N_2860);
xor U9118 (N_9118,N_613,N_1847);
and U9119 (N_9119,N_725,N_1540);
xnor U9120 (N_9120,N_3694,N_3682);
nand U9121 (N_9121,N_522,N_4000);
nand U9122 (N_9122,N_123,N_172);
xnor U9123 (N_9123,N_3890,N_2961);
and U9124 (N_9124,N_1479,N_798);
nor U9125 (N_9125,N_3047,N_4083);
xor U9126 (N_9126,N_984,N_3470);
nor U9127 (N_9127,N_2954,N_4213);
nand U9128 (N_9128,N_4972,N_2537);
xnor U9129 (N_9129,N_3743,N_3046);
or U9130 (N_9130,N_858,N_3633);
and U9131 (N_9131,N_2301,N_553);
nor U9132 (N_9132,N_1389,N_4162);
and U9133 (N_9133,N_2143,N_1626);
nor U9134 (N_9134,N_2367,N_3222);
nor U9135 (N_9135,N_3709,N_1313);
xnor U9136 (N_9136,N_4147,N_1235);
nor U9137 (N_9137,N_4673,N_2079);
and U9138 (N_9138,N_2751,N_4906);
and U9139 (N_9139,N_4578,N_2598);
nand U9140 (N_9140,N_4102,N_1779);
and U9141 (N_9141,N_1893,N_3178);
nand U9142 (N_9142,N_3920,N_1501);
nand U9143 (N_9143,N_2796,N_3753);
xnor U9144 (N_9144,N_3405,N_3292);
nor U9145 (N_9145,N_1863,N_4029);
or U9146 (N_9146,N_3506,N_11);
nand U9147 (N_9147,N_1833,N_1584);
or U9148 (N_9148,N_1072,N_3094);
xor U9149 (N_9149,N_3426,N_679);
nand U9150 (N_9150,N_2438,N_127);
nand U9151 (N_9151,N_967,N_849);
and U9152 (N_9152,N_1623,N_841);
nor U9153 (N_9153,N_4016,N_1426);
nand U9154 (N_9154,N_2558,N_252);
nor U9155 (N_9155,N_1320,N_1600);
nor U9156 (N_9156,N_173,N_1104);
and U9157 (N_9157,N_3323,N_3605);
or U9158 (N_9158,N_1518,N_670);
or U9159 (N_9159,N_2138,N_528);
nor U9160 (N_9160,N_3967,N_1135);
xor U9161 (N_9161,N_1718,N_2859);
nor U9162 (N_9162,N_4402,N_1207);
nor U9163 (N_9163,N_4153,N_2909);
and U9164 (N_9164,N_4144,N_4066);
nand U9165 (N_9165,N_300,N_4412);
nand U9166 (N_9166,N_118,N_761);
nor U9167 (N_9167,N_1140,N_4062);
or U9168 (N_9168,N_353,N_3465);
nand U9169 (N_9169,N_4887,N_3507);
nand U9170 (N_9170,N_3839,N_798);
xnor U9171 (N_9171,N_1099,N_4939);
nor U9172 (N_9172,N_2713,N_4874);
and U9173 (N_9173,N_2516,N_2258);
nor U9174 (N_9174,N_3981,N_2974);
nor U9175 (N_9175,N_2551,N_499);
xor U9176 (N_9176,N_2220,N_3359);
xnor U9177 (N_9177,N_61,N_689);
nor U9178 (N_9178,N_3457,N_2248);
xnor U9179 (N_9179,N_1286,N_2214);
xor U9180 (N_9180,N_1899,N_1454);
nand U9181 (N_9181,N_2842,N_212);
nor U9182 (N_9182,N_3919,N_3004);
xnor U9183 (N_9183,N_3106,N_2057);
nor U9184 (N_9184,N_4580,N_4023);
nand U9185 (N_9185,N_3015,N_2562);
and U9186 (N_9186,N_2953,N_3427);
nor U9187 (N_9187,N_3003,N_3868);
or U9188 (N_9188,N_415,N_3990);
or U9189 (N_9189,N_3083,N_1811);
nand U9190 (N_9190,N_526,N_2452);
and U9191 (N_9191,N_4105,N_414);
or U9192 (N_9192,N_217,N_2683);
nand U9193 (N_9193,N_928,N_4905);
xnor U9194 (N_9194,N_4437,N_1834);
nor U9195 (N_9195,N_3771,N_3156);
and U9196 (N_9196,N_1854,N_2313);
and U9197 (N_9197,N_1289,N_3203);
nand U9198 (N_9198,N_53,N_1276);
and U9199 (N_9199,N_223,N_4508);
nor U9200 (N_9200,N_2780,N_3602);
xnor U9201 (N_9201,N_1263,N_2970);
and U9202 (N_9202,N_1325,N_3041);
nor U9203 (N_9203,N_4874,N_1150);
and U9204 (N_9204,N_693,N_4559);
and U9205 (N_9205,N_419,N_3657);
or U9206 (N_9206,N_4629,N_1687);
nand U9207 (N_9207,N_4459,N_628);
nand U9208 (N_9208,N_3743,N_2386);
xnor U9209 (N_9209,N_1757,N_3512);
nand U9210 (N_9210,N_4188,N_2297);
and U9211 (N_9211,N_4414,N_503);
nor U9212 (N_9212,N_54,N_4393);
and U9213 (N_9213,N_1066,N_2815);
and U9214 (N_9214,N_3372,N_3848);
and U9215 (N_9215,N_4875,N_4245);
nor U9216 (N_9216,N_723,N_4704);
and U9217 (N_9217,N_601,N_2851);
and U9218 (N_9218,N_232,N_4445);
nor U9219 (N_9219,N_2737,N_2937);
nor U9220 (N_9220,N_3541,N_268);
or U9221 (N_9221,N_1677,N_1713);
or U9222 (N_9222,N_3937,N_3416);
nand U9223 (N_9223,N_108,N_2323);
and U9224 (N_9224,N_633,N_1614);
nand U9225 (N_9225,N_3356,N_267);
nor U9226 (N_9226,N_2726,N_1742);
or U9227 (N_9227,N_123,N_3505);
or U9228 (N_9228,N_2358,N_1843);
and U9229 (N_9229,N_1836,N_1734);
xnor U9230 (N_9230,N_2656,N_4336);
and U9231 (N_9231,N_2633,N_473);
nand U9232 (N_9232,N_523,N_1706);
and U9233 (N_9233,N_3134,N_1566);
nand U9234 (N_9234,N_4670,N_3883);
and U9235 (N_9235,N_3427,N_1379);
and U9236 (N_9236,N_3901,N_1553);
nand U9237 (N_9237,N_3176,N_260);
xnor U9238 (N_9238,N_2500,N_4878);
and U9239 (N_9239,N_1479,N_2456);
or U9240 (N_9240,N_2881,N_4760);
or U9241 (N_9241,N_2687,N_4943);
nor U9242 (N_9242,N_2277,N_469);
nand U9243 (N_9243,N_3227,N_3434);
and U9244 (N_9244,N_3866,N_2758);
or U9245 (N_9245,N_3360,N_4475);
xnor U9246 (N_9246,N_1332,N_2706);
nand U9247 (N_9247,N_3752,N_2360);
nand U9248 (N_9248,N_3228,N_3472);
or U9249 (N_9249,N_2338,N_2318);
xnor U9250 (N_9250,N_1989,N_880);
xnor U9251 (N_9251,N_70,N_3437);
and U9252 (N_9252,N_4447,N_1251);
or U9253 (N_9253,N_2631,N_412);
xnor U9254 (N_9254,N_4768,N_2734);
or U9255 (N_9255,N_3573,N_241);
xor U9256 (N_9256,N_2036,N_1026);
xnor U9257 (N_9257,N_4596,N_2225);
xnor U9258 (N_9258,N_767,N_3166);
and U9259 (N_9259,N_1310,N_2125);
xor U9260 (N_9260,N_602,N_4962);
nor U9261 (N_9261,N_1262,N_3299);
and U9262 (N_9262,N_1613,N_2285);
nand U9263 (N_9263,N_925,N_354);
and U9264 (N_9264,N_3690,N_469);
nand U9265 (N_9265,N_3259,N_3476);
xor U9266 (N_9266,N_4714,N_3841);
nor U9267 (N_9267,N_4497,N_2665);
nor U9268 (N_9268,N_4057,N_3589);
or U9269 (N_9269,N_2549,N_25);
or U9270 (N_9270,N_1491,N_4415);
nor U9271 (N_9271,N_3017,N_382);
nand U9272 (N_9272,N_2793,N_2861);
xnor U9273 (N_9273,N_2580,N_4011);
and U9274 (N_9274,N_3191,N_3927);
or U9275 (N_9275,N_967,N_3532);
nand U9276 (N_9276,N_1381,N_3210);
nand U9277 (N_9277,N_834,N_4472);
xor U9278 (N_9278,N_3029,N_3080);
and U9279 (N_9279,N_901,N_2040);
nor U9280 (N_9280,N_1506,N_1995);
nand U9281 (N_9281,N_852,N_3656);
or U9282 (N_9282,N_1793,N_2882);
and U9283 (N_9283,N_1532,N_1584);
and U9284 (N_9284,N_3428,N_1491);
and U9285 (N_9285,N_3949,N_3707);
or U9286 (N_9286,N_3086,N_4492);
and U9287 (N_9287,N_3396,N_2724);
xor U9288 (N_9288,N_2842,N_950);
nor U9289 (N_9289,N_796,N_2031);
nor U9290 (N_9290,N_172,N_1967);
nand U9291 (N_9291,N_4567,N_848);
and U9292 (N_9292,N_3149,N_2371);
and U9293 (N_9293,N_3240,N_4564);
xor U9294 (N_9294,N_1948,N_2829);
nand U9295 (N_9295,N_4350,N_2468);
and U9296 (N_9296,N_452,N_2391);
or U9297 (N_9297,N_1685,N_1989);
nor U9298 (N_9298,N_2317,N_679);
and U9299 (N_9299,N_4657,N_4232);
nor U9300 (N_9300,N_3418,N_3044);
or U9301 (N_9301,N_2000,N_4715);
and U9302 (N_9302,N_308,N_1728);
nor U9303 (N_9303,N_1749,N_878);
nor U9304 (N_9304,N_1618,N_4832);
and U9305 (N_9305,N_55,N_4793);
nand U9306 (N_9306,N_1323,N_838);
xnor U9307 (N_9307,N_3731,N_239);
xnor U9308 (N_9308,N_1957,N_3274);
nor U9309 (N_9309,N_533,N_769);
or U9310 (N_9310,N_2708,N_408);
nor U9311 (N_9311,N_614,N_4430);
nor U9312 (N_9312,N_716,N_1944);
nor U9313 (N_9313,N_241,N_2940);
xor U9314 (N_9314,N_2650,N_864);
nand U9315 (N_9315,N_2575,N_2006);
nand U9316 (N_9316,N_988,N_3895);
nor U9317 (N_9317,N_693,N_119);
or U9318 (N_9318,N_1164,N_2752);
xnor U9319 (N_9319,N_3799,N_3946);
and U9320 (N_9320,N_1992,N_809);
or U9321 (N_9321,N_3669,N_4920);
nand U9322 (N_9322,N_4615,N_1978);
and U9323 (N_9323,N_1942,N_116);
nand U9324 (N_9324,N_2472,N_2143);
and U9325 (N_9325,N_2572,N_422);
and U9326 (N_9326,N_4083,N_2162);
nand U9327 (N_9327,N_3737,N_4795);
xor U9328 (N_9328,N_1953,N_2713);
or U9329 (N_9329,N_3160,N_3238);
or U9330 (N_9330,N_3964,N_2443);
nand U9331 (N_9331,N_876,N_1440);
and U9332 (N_9332,N_4355,N_2652);
and U9333 (N_9333,N_766,N_1950);
nand U9334 (N_9334,N_1150,N_633);
nor U9335 (N_9335,N_1175,N_1776);
and U9336 (N_9336,N_1406,N_2385);
or U9337 (N_9337,N_2669,N_1893);
xnor U9338 (N_9338,N_2431,N_4248);
nand U9339 (N_9339,N_3166,N_1182);
xor U9340 (N_9340,N_3063,N_3081);
nor U9341 (N_9341,N_948,N_2714);
xnor U9342 (N_9342,N_279,N_3933);
nand U9343 (N_9343,N_1278,N_1745);
and U9344 (N_9344,N_2737,N_3531);
nand U9345 (N_9345,N_1677,N_2017);
or U9346 (N_9346,N_830,N_3340);
and U9347 (N_9347,N_2202,N_2674);
nor U9348 (N_9348,N_3201,N_4697);
nor U9349 (N_9349,N_3205,N_2194);
nand U9350 (N_9350,N_2772,N_1420);
nor U9351 (N_9351,N_940,N_3309);
nand U9352 (N_9352,N_3251,N_1120);
nand U9353 (N_9353,N_3477,N_2410);
nand U9354 (N_9354,N_3434,N_1055);
or U9355 (N_9355,N_4161,N_605);
and U9356 (N_9356,N_26,N_3017);
and U9357 (N_9357,N_4259,N_3876);
xnor U9358 (N_9358,N_1143,N_4581);
nand U9359 (N_9359,N_2433,N_1178);
and U9360 (N_9360,N_3546,N_240);
nor U9361 (N_9361,N_2272,N_3007);
nand U9362 (N_9362,N_289,N_133);
xor U9363 (N_9363,N_457,N_2737);
nor U9364 (N_9364,N_1583,N_2434);
nor U9365 (N_9365,N_1767,N_1413);
or U9366 (N_9366,N_3926,N_4232);
or U9367 (N_9367,N_427,N_2103);
xor U9368 (N_9368,N_1273,N_3840);
nand U9369 (N_9369,N_2057,N_3705);
nand U9370 (N_9370,N_2128,N_4330);
nor U9371 (N_9371,N_3564,N_273);
nand U9372 (N_9372,N_1202,N_1183);
or U9373 (N_9373,N_1923,N_1454);
xnor U9374 (N_9374,N_4288,N_4607);
nand U9375 (N_9375,N_328,N_3229);
xnor U9376 (N_9376,N_3780,N_2080);
or U9377 (N_9377,N_2051,N_3926);
nor U9378 (N_9378,N_1164,N_1589);
or U9379 (N_9379,N_2843,N_3217);
xnor U9380 (N_9380,N_4752,N_302);
and U9381 (N_9381,N_3101,N_4546);
nand U9382 (N_9382,N_3401,N_2229);
and U9383 (N_9383,N_83,N_202);
and U9384 (N_9384,N_266,N_962);
nor U9385 (N_9385,N_1753,N_3700);
xor U9386 (N_9386,N_624,N_4874);
xnor U9387 (N_9387,N_1056,N_3928);
or U9388 (N_9388,N_538,N_82);
xnor U9389 (N_9389,N_1874,N_1898);
nand U9390 (N_9390,N_4929,N_4347);
nor U9391 (N_9391,N_704,N_3679);
and U9392 (N_9392,N_1688,N_1765);
and U9393 (N_9393,N_1689,N_4892);
and U9394 (N_9394,N_508,N_3079);
xnor U9395 (N_9395,N_3312,N_559);
and U9396 (N_9396,N_1152,N_643);
and U9397 (N_9397,N_2099,N_2961);
nor U9398 (N_9398,N_2842,N_2206);
nand U9399 (N_9399,N_3461,N_3134);
or U9400 (N_9400,N_1358,N_4);
nor U9401 (N_9401,N_585,N_3412);
or U9402 (N_9402,N_642,N_3752);
nand U9403 (N_9403,N_4041,N_4542);
nand U9404 (N_9404,N_1277,N_1255);
xnor U9405 (N_9405,N_2148,N_2061);
nand U9406 (N_9406,N_2603,N_4043);
nand U9407 (N_9407,N_4830,N_3298);
nand U9408 (N_9408,N_1956,N_2821);
xnor U9409 (N_9409,N_2340,N_3039);
or U9410 (N_9410,N_2080,N_1177);
xor U9411 (N_9411,N_303,N_872);
nor U9412 (N_9412,N_1447,N_1984);
and U9413 (N_9413,N_2503,N_3496);
or U9414 (N_9414,N_4521,N_683);
xnor U9415 (N_9415,N_2104,N_3024);
or U9416 (N_9416,N_605,N_4368);
or U9417 (N_9417,N_369,N_4593);
and U9418 (N_9418,N_165,N_2704);
nand U9419 (N_9419,N_4185,N_1315);
and U9420 (N_9420,N_3173,N_3615);
nor U9421 (N_9421,N_3113,N_4448);
xnor U9422 (N_9422,N_1829,N_1340);
or U9423 (N_9423,N_2826,N_4135);
and U9424 (N_9424,N_1954,N_3169);
nor U9425 (N_9425,N_3309,N_4620);
xor U9426 (N_9426,N_4598,N_1021);
or U9427 (N_9427,N_2684,N_319);
nor U9428 (N_9428,N_2757,N_213);
and U9429 (N_9429,N_3564,N_1722);
xnor U9430 (N_9430,N_598,N_112);
nand U9431 (N_9431,N_4701,N_522);
or U9432 (N_9432,N_4811,N_2845);
nor U9433 (N_9433,N_1050,N_1490);
and U9434 (N_9434,N_783,N_4231);
or U9435 (N_9435,N_2998,N_1239);
and U9436 (N_9436,N_2669,N_1915);
xor U9437 (N_9437,N_3633,N_4880);
or U9438 (N_9438,N_3030,N_1206);
and U9439 (N_9439,N_65,N_3233);
or U9440 (N_9440,N_2382,N_3775);
nand U9441 (N_9441,N_154,N_1455);
nor U9442 (N_9442,N_1166,N_313);
and U9443 (N_9443,N_1627,N_3912);
and U9444 (N_9444,N_1168,N_2379);
nor U9445 (N_9445,N_3932,N_467);
nor U9446 (N_9446,N_1939,N_381);
nor U9447 (N_9447,N_2449,N_43);
nor U9448 (N_9448,N_4544,N_3601);
or U9449 (N_9449,N_1495,N_2093);
and U9450 (N_9450,N_619,N_485);
or U9451 (N_9451,N_3742,N_1152);
xnor U9452 (N_9452,N_1475,N_1914);
nor U9453 (N_9453,N_2129,N_3272);
xor U9454 (N_9454,N_4348,N_4681);
or U9455 (N_9455,N_49,N_3166);
or U9456 (N_9456,N_740,N_1626);
and U9457 (N_9457,N_3713,N_3619);
nor U9458 (N_9458,N_1643,N_1640);
and U9459 (N_9459,N_2167,N_2300);
or U9460 (N_9460,N_887,N_3982);
or U9461 (N_9461,N_4980,N_1172);
nor U9462 (N_9462,N_3518,N_4420);
or U9463 (N_9463,N_4091,N_1560);
and U9464 (N_9464,N_2680,N_59);
and U9465 (N_9465,N_1237,N_4606);
nand U9466 (N_9466,N_989,N_3807);
nand U9467 (N_9467,N_458,N_3182);
nand U9468 (N_9468,N_2834,N_2102);
nand U9469 (N_9469,N_1838,N_1045);
and U9470 (N_9470,N_4042,N_3194);
xor U9471 (N_9471,N_3372,N_2836);
xnor U9472 (N_9472,N_1952,N_253);
or U9473 (N_9473,N_1892,N_4607);
xnor U9474 (N_9474,N_4048,N_2134);
nor U9475 (N_9475,N_850,N_4097);
nand U9476 (N_9476,N_4113,N_285);
nand U9477 (N_9477,N_56,N_2141);
xor U9478 (N_9478,N_4075,N_1700);
and U9479 (N_9479,N_3889,N_121);
and U9480 (N_9480,N_818,N_2404);
nor U9481 (N_9481,N_1427,N_2950);
nor U9482 (N_9482,N_4718,N_3519);
xor U9483 (N_9483,N_2193,N_3344);
nor U9484 (N_9484,N_3500,N_2873);
nand U9485 (N_9485,N_4883,N_3794);
nand U9486 (N_9486,N_213,N_2232);
nand U9487 (N_9487,N_4185,N_1123);
or U9488 (N_9488,N_261,N_4445);
nor U9489 (N_9489,N_4676,N_1470);
xor U9490 (N_9490,N_3671,N_3733);
xnor U9491 (N_9491,N_1953,N_763);
and U9492 (N_9492,N_3185,N_3736);
xnor U9493 (N_9493,N_4119,N_4027);
nor U9494 (N_9494,N_3052,N_2805);
nor U9495 (N_9495,N_3011,N_4791);
nor U9496 (N_9496,N_2864,N_449);
nor U9497 (N_9497,N_4365,N_525);
nand U9498 (N_9498,N_2636,N_3047);
or U9499 (N_9499,N_919,N_3792);
nor U9500 (N_9500,N_1154,N_658);
and U9501 (N_9501,N_4757,N_4667);
or U9502 (N_9502,N_2453,N_2812);
or U9503 (N_9503,N_3894,N_350);
or U9504 (N_9504,N_1683,N_2468);
nor U9505 (N_9505,N_2950,N_2295);
nor U9506 (N_9506,N_1007,N_4725);
nand U9507 (N_9507,N_3932,N_1755);
nand U9508 (N_9508,N_2053,N_2387);
or U9509 (N_9509,N_2556,N_4480);
or U9510 (N_9510,N_3051,N_3902);
or U9511 (N_9511,N_2833,N_22);
xor U9512 (N_9512,N_2429,N_763);
nand U9513 (N_9513,N_2764,N_3541);
and U9514 (N_9514,N_4664,N_3338);
nand U9515 (N_9515,N_4452,N_1467);
nor U9516 (N_9516,N_3597,N_803);
and U9517 (N_9517,N_2456,N_1900);
nand U9518 (N_9518,N_948,N_1576);
nor U9519 (N_9519,N_4249,N_2065);
or U9520 (N_9520,N_3891,N_881);
nor U9521 (N_9521,N_2476,N_3828);
and U9522 (N_9522,N_2222,N_4714);
xor U9523 (N_9523,N_2216,N_3774);
nor U9524 (N_9524,N_3014,N_2815);
nor U9525 (N_9525,N_3516,N_3416);
xnor U9526 (N_9526,N_2971,N_294);
or U9527 (N_9527,N_4459,N_511);
and U9528 (N_9528,N_3740,N_2659);
nor U9529 (N_9529,N_723,N_1150);
or U9530 (N_9530,N_2375,N_648);
or U9531 (N_9531,N_2522,N_2323);
and U9532 (N_9532,N_2263,N_4237);
nand U9533 (N_9533,N_472,N_869);
xnor U9534 (N_9534,N_1336,N_3387);
nand U9535 (N_9535,N_2415,N_1377);
or U9536 (N_9536,N_1021,N_3529);
nor U9537 (N_9537,N_133,N_1642);
and U9538 (N_9538,N_1389,N_455);
nor U9539 (N_9539,N_150,N_2410);
or U9540 (N_9540,N_1178,N_285);
nor U9541 (N_9541,N_1177,N_3419);
or U9542 (N_9542,N_750,N_688);
or U9543 (N_9543,N_1939,N_1068);
xnor U9544 (N_9544,N_1464,N_1878);
and U9545 (N_9545,N_224,N_3089);
nor U9546 (N_9546,N_4601,N_1691);
and U9547 (N_9547,N_180,N_543);
and U9548 (N_9548,N_2061,N_873);
xnor U9549 (N_9549,N_2780,N_3723);
nor U9550 (N_9550,N_369,N_3197);
nand U9551 (N_9551,N_1544,N_2351);
xor U9552 (N_9552,N_2310,N_2673);
nor U9553 (N_9553,N_3415,N_2380);
xor U9554 (N_9554,N_4905,N_1983);
nand U9555 (N_9555,N_451,N_679);
or U9556 (N_9556,N_1786,N_897);
and U9557 (N_9557,N_2272,N_20);
xnor U9558 (N_9558,N_3330,N_4659);
or U9559 (N_9559,N_2563,N_1705);
nand U9560 (N_9560,N_3660,N_4711);
or U9561 (N_9561,N_2859,N_1216);
nor U9562 (N_9562,N_722,N_4553);
xnor U9563 (N_9563,N_984,N_3740);
nand U9564 (N_9564,N_318,N_4593);
xor U9565 (N_9565,N_2804,N_1345);
and U9566 (N_9566,N_2649,N_4006);
xor U9567 (N_9567,N_866,N_1980);
xor U9568 (N_9568,N_2300,N_2690);
and U9569 (N_9569,N_2422,N_2722);
nor U9570 (N_9570,N_4113,N_719);
and U9571 (N_9571,N_3783,N_4086);
or U9572 (N_9572,N_2356,N_263);
xnor U9573 (N_9573,N_4499,N_4324);
nand U9574 (N_9574,N_649,N_4516);
nand U9575 (N_9575,N_1312,N_1879);
or U9576 (N_9576,N_1814,N_2122);
nand U9577 (N_9577,N_500,N_2893);
xor U9578 (N_9578,N_3073,N_3918);
and U9579 (N_9579,N_2303,N_1110);
nand U9580 (N_9580,N_4736,N_4053);
xnor U9581 (N_9581,N_4399,N_4078);
or U9582 (N_9582,N_1255,N_1946);
xnor U9583 (N_9583,N_1808,N_1418);
nor U9584 (N_9584,N_3177,N_4689);
or U9585 (N_9585,N_2271,N_3215);
nand U9586 (N_9586,N_3951,N_3088);
xnor U9587 (N_9587,N_1404,N_3822);
and U9588 (N_9588,N_541,N_2830);
xnor U9589 (N_9589,N_4840,N_1952);
and U9590 (N_9590,N_1436,N_2509);
xnor U9591 (N_9591,N_3154,N_2738);
xor U9592 (N_9592,N_1275,N_2870);
nand U9593 (N_9593,N_310,N_2386);
nor U9594 (N_9594,N_4673,N_3143);
xor U9595 (N_9595,N_794,N_4941);
or U9596 (N_9596,N_4023,N_4694);
and U9597 (N_9597,N_2478,N_1024);
or U9598 (N_9598,N_2847,N_280);
nor U9599 (N_9599,N_3724,N_837);
nor U9600 (N_9600,N_279,N_1792);
or U9601 (N_9601,N_2629,N_4054);
xnor U9602 (N_9602,N_1331,N_4791);
nor U9603 (N_9603,N_3715,N_4338);
xnor U9604 (N_9604,N_1202,N_1678);
xnor U9605 (N_9605,N_1900,N_3494);
or U9606 (N_9606,N_3153,N_3306);
and U9607 (N_9607,N_4100,N_4080);
xnor U9608 (N_9608,N_4199,N_887);
nand U9609 (N_9609,N_3645,N_2781);
nand U9610 (N_9610,N_1301,N_499);
and U9611 (N_9611,N_3357,N_877);
or U9612 (N_9612,N_473,N_3968);
and U9613 (N_9613,N_4646,N_3320);
nand U9614 (N_9614,N_1819,N_2260);
and U9615 (N_9615,N_3067,N_494);
and U9616 (N_9616,N_2493,N_2131);
xnor U9617 (N_9617,N_4146,N_1267);
nand U9618 (N_9618,N_3146,N_1101);
xnor U9619 (N_9619,N_2644,N_2696);
nor U9620 (N_9620,N_3080,N_1701);
nand U9621 (N_9621,N_1801,N_989);
or U9622 (N_9622,N_848,N_2177);
or U9623 (N_9623,N_1088,N_2308);
nor U9624 (N_9624,N_18,N_503);
nand U9625 (N_9625,N_4276,N_2061);
or U9626 (N_9626,N_2973,N_1035);
and U9627 (N_9627,N_4626,N_3440);
nand U9628 (N_9628,N_1637,N_2355);
nor U9629 (N_9629,N_4447,N_1305);
or U9630 (N_9630,N_3856,N_1839);
nand U9631 (N_9631,N_1571,N_1361);
nor U9632 (N_9632,N_2734,N_1969);
nand U9633 (N_9633,N_1409,N_96);
and U9634 (N_9634,N_1265,N_2574);
nor U9635 (N_9635,N_3056,N_2254);
nand U9636 (N_9636,N_561,N_1153);
and U9637 (N_9637,N_2380,N_876);
xor U9638 (N_9638,N_3483,N_1741);
nor U9639 (N_9639,N_4783,N_1379);
and U9640 (N_9640,N_4183,N_2548);
xor U9641 (N_9641,N_1152,N_3183);
and U9642 (N_9642,N_3058,N_2981);
xor U9643 (N_9643,N_1883,N_4613);
or U9644 (N_9644,N_4140,N_229);
nor U9645 (N_9645,N_1348,N_3057);
and U9646 (N_9646,N_542,N_399);
nor U9647 (N_9647,N_1371,N_2966);
and U9648 (N_9648,N_4288,N_3103);
nor U9649 (N_9649,N_2653,N_3165);
xnor U9650 (N_9650,N_4700,N_2007);
or U9651 (N_9651,N_715,N_4559);
xor U9652 (N_9652,N_931,N_4385);
xnor U9653 (N_9653,N_1911,N_647);
xnor U9654 (N_9654,N_44,N_48);
nor U9655 (N_9655,N_2242,N_3490);
or U9656 (N_9656,N_4192,N_3190);
nand U9657 (N_9657,N_4330,N_641);
nor U9658 (N_9658,N_874,N_2831);
or U9659 (N_9659,N_4690,N_1133);
nor U9660 (N_9660,N_4075,N_1937);
nor U9661 (N_9661,N_579,N_1581);
and U9662 (N_9662,N_4217,N_4323);
nor U9663 (N_9663,N_379,N_1213);
xnor U9664 (N_9664,N_1638,N_4106);
nand U9665 (N_9665,N_4950,N_2928);
or U9666 (N_9666,N_2959,N_3003);
or U9667 (N_9667,N_4166,N_159);
nor U9668 (N_9668,N_813,N_3642);
and U9669 (N_9669,N_174,N_4554);
or U9670 (N_9670,N_1560,N_1309);
or U9671 (N_9671,N_2831,N_4570);
nor U9672 (N_9672,N_2188,N_1696);
and U9673 (N_9673,N_791,N_823);
xor U9674 (N_9674,N_2002,N_3191);
xnor U9675 (N_9675,N_3315,N_4589);
nor U9676 (N_9676,N_1274,N_96);
and U9677 (N_9677,N_2955,N_2072);
nand U9678 (N_9678,N_2433,N_3772);
nand U9679 (N_9679,N_1528,N_3885);
xnor U9680 (N_9680,N_4860,N_3898);
nor U9681 (N_9681,N_1450,N_3432);
nand U9682 (N_9682,N_3905,N_953);
xnor U9683 (N_9683,N_1298,N_295);
xor U9684 (N_9684,N_4857,N_3649);
or U9685 (N_9685,N_4833,N_1511);
nor U9686 (N_9686,N_1893,N_4000);
and U9687 (N_9687,N_1121,N_3589);
or U9688 (N_9688,N_3634,N_2049);
xor U9689 (N_9689,N_2902,N_432);
and U9690 (N_9690,N_3217,N_2496);
nand U9691 (N_9691,N_2241,N_2366);
nand U9692 (N_9692,N_4195,N_2405);
and U9693 (N_9693,N_2136,N_4563);
or U9694 (N_9694,N_1769,N_2628);
nand U9695 (N_9695,N_523,N_311);
or U9696 (N_9696,N_3045,N_3159);
nand U9697 (N_9697,N_4060,N_2274);
nor U9698 (N_9698,N_4734,N_2846);
or U9699 (N_9699,N_2917,N_4960);
and U9700 (N_9700,N_3441,N_243);
and U9701 (N_9701,N_2269,N_4142);
xor U9702 (N_9702,N_2312,N_688);
nand U9703 (N_9703,N_2413,N_387);
or U9704 (N_9704,N_2404,N_3772);
or U9705 (N_9705,N_3056,N_2423);
nor U9706 (N_9706,N_1672,N_2631);
nor U9707 (N_9707,N_3001,N_4502);
and U9708 (N_9708,N_3573,N_511);
xor U9709 (N_9709,N_3341,N_930);
nor U9710 (N_9710,N_2756,N_3503);
or U9711 (N_9711,N_1722,N_1473);
xor U9712 (N_9712,N_3021,N_312);
xnor U9713 (N_9713,N_2645,N_615);
and U9714 (N_9714,N_3175,N_897);
nor U9715 (N_9715,N_3267,N_4197);
nor U9716 (N_9716,N_1128,N_2368);
xor U9717 (N_9717,N_2336,N_4901);
xnor U9718 (N_9718,N_1659,N_1802);
nand U9719 (N_9719,N_4103,N_551);
nor U9720 (N_9720,N_9,N_334);
and U9721 (N_9721,N_4886,N_62);
or U9722 (N_9722,N_2003,N_1388);
nand U9723 (N_9723,N_492,N_3650);
nand U9724 (N_9724,N_1942,N_3994);
xor U9725 (N_9725,N_2063,N_454);
nand U9726 (N_9726,N_1685,N_1257);
and U9727 (N_9727,N_4665,N_1964);
nand U9728 (N_9728,N_1080,N_4823);
or U9729 (N_9729,N_852,N_3802);
nor U9730 (N_9730,N_4392,N_3249);
nor U9731 (N_9731,N_4199,N_1997);
xor U9732 (N_9732,N_2881,N_2157);
and U9733 (N_9733,N_3229,N_2668);
xor U9734 (N_9734,N_3853,N_4230);
or U9735 (N_9735,N_4520,N_1450);
and U9736 (N_9736,N_3361,N_2499);
nor U9737 (N_9737,N_1954,N_2894);
nor U9738 (N_9738,N_2912,N_1515);
and U9739 (N_9739,N_4261,N_504);
nor U9740 (N_9740,N_2675,N_3201);
xnor U9741 (N_9741,N_4606,N_4361);
nor U9742 (N_9742,N_2670,N_13);
and U9743 (N_9743,N_2867,N_1488);
xnor U9744 (N_9744,N_3736,N_3084);
and U9745 (N_9745,N_2340,N_3131);
nand U9746 (N_9746,N_1477,N_4320);
and U9747 (N_9747,N_3287,N_836);
nor U9748 (N_9748,N_2619,N_2296);
nor U9749 (N_9749,N_2043,N_1539);
and U9750 (N_9750,N_2027,N_853);
nand U9751 (N_9751,N_2316,N_4313);
nor U9752 (N_9752,N_4281,N_2975);
and U9753 (N_9753,N_2982,N_2875);
nor U9754 (N_9754,N_2407,N_4544);
and U9755 (N_9755,N_2319,N_3493);
xor U9756 (N_9756,N_2053,N_2336);
or U9757 (N_9757,N_3614,N_655);
nor U9758 (N_9758,N_738,N_2218);
nand U9759 (N_9759,N_4585,N_4727);
or U9760 (N_9760,N_4868,N_1039);
xnor U9761 (N_9761,N_3996,N_4409);
xnor U9762 (N_9762,N_2017,N_3622);
or U9763 (N_9763,N_3228,N_2661);
nand U9764 (N_9764,N_375,N_4847);
nor U9765 (N_9765,N_4358,N_4761);
or U9766 (N_9766,N_554,N_4595);
xnor U9767 (N_9767,N_3561,N_1194);
or U9768 (N_9768,N_1121,N_2417);
or U9769 (N_9769,N_1670,N_2234);
and U9770 (N_9770,N_203,N_2061);
and U9771 (N_9771,N_1789,N_2357);
nor U9772 (N_9772,N_3126,N_1775);
xor U9773 (N_9773,N_1355,N_1959);
or U9774 (N_9774,N_219,N_4345);
and U9775 (N_9775,N_1509,N_932);
and U9776 (N_9776,N_3115,N_2161);
nor U9777 (N_9777,N_2326,N_1930);
nand U9778 (N_9778,N_153,N_1353);
nand U9779 (N_9779,N_273,N_3595);
nand U9780 (N_9780,N_1134,N_1445);
or U9781 (N_9781,N_238,N_4775);
nand U9782 (N_9782,N_3094,N_4861);
nand U9783 (N_9783,N_2904,N_3600);
nor U9784 (N_9784,N_475,N_3334);
or U9785 (N_9785,N_294,N_1402);
nor U9786 (N_9786,N_1728,N_3634);
xnor U9787 (N_9787,N_4186,N_1213);
or U9788 (N_9788,N_4821,N_2831);
nor U9789 (N_9789,N_2870,N_614);
or U9790 (N_9790,N_1658,N_140);
nor U9791 (N_9791,N_1759,N_2277);
or U9792 (N_9792,N_2328,N_3232);
or U9793 (N_9793,N_2916,N_118);
xnor U9794 (N_9794,N_3548,N_3706);
or U9795 (N_9795,N_4337,N_4533);
and U9796 (N_9796,N_2399,N_1053);
nor U9797 (N_9797,N_4380,N_966);
xnor U9798 (N_9798,N_269,N_1201);
and U9799 (N_9799,N_3587,N_1453);
nor U9800 (N_9800,N_971,N_2580);
and U9801 (N_9801,N_3695,N_4696);
or U9802 (N_9802,N_4539,N_147);
or U9803 (N_9803,N_3513,N_900);
xor U9804 (N_9804,N_167,N_1277);
xnor U9805 (N_9805,N_131,N_1165);
nand U9806 (N_9806,N_2545,N_2193);
or U9807 (N_9807,N_129,N_3557);
and U9808 (N_9808,N_2492,N_1629);
or U9809 (N_9809,N_1047,N_953);
or U9810 (N_9810,N_4046,N_4979);
nor U9811 (N_9811,N_4511,N_975);
xor U9812 (N_9812,N_3808,N_4411);
nor U9813 (N_9813,N_4085,N_950);
xnor U9814 (N_9814,N_4073,N_4052);
or U9815 (N_9815,N_4183,N_2239);
nor U9816 (N_9816,N_1543,N_2184);
xnor U9817 (N_9817,N_3147,N_2554);
nor U9818 (N_9818,N_886,N_4962);
nand U9819 (N_9819,N_2166,N_2752);
xor U9820 (N_9820,N_2350,N_1473);
xor U9821 (N_9821,N_3209,N_2862);
xor U9822 (N_9822,N_3647,N_3223);
and U9823 (N_9823,N_4804,N_3587);
or U9824 (N_9824,N_2141,N_959);
xor U9825 (N_9825,N_2117,N_3535);
nor U9826 (N_9826,N_4110,N_1334);
nor U9827 (N_9827,N_1366,N_2435);
nor U9828 (N_9828,N_4905,N_1985);
and U9829 (N_9829,N_3883,N_1767);
and U9830 (N_9830,N_4588,N_649);
and U9831 (N_9831,N_4619,N_3628);
nand U9832 (N_9832,N_3065,N_1355);
nor U9833 (N_9833,N_1019,N_2174);
or U9834 (N_9834,N_23,N_3222);
nand U9835 (N_9835,N_2323,N_3765);
nor U9836 (N_9836,N_4992,N_3534);
nor U9837 (N_9837,N_4653,N_306);
xnor U9838 (N_9838,N_3490,N_1351);
nor U9839 (N_9839,N_4662,N_1706);
or U9840 (N_9840,N_3247,N_4297);
nand U9841 (N_9841,N_4184,N_2589);
nand U9842 (N_9842,N_3670,N_4356);
nor U9843 (N_9843,N_4893,N_4173);
xor U9844 (N_9844,N_919,N_4700);
and U9845 (N_9845,N_956,N_3833);
xor U9846 (N_9846,N_184,N_1580);
nand U9847 (N_9847,N_979,N_3788);
nand U9848 (N_9848,N_3517,N_4268);
nand U9849 (N_9849,N_119,N_3989);
or U9850 (N_9850,N_1716,N_4686);
nand U9851 (N_9851,N_4871,N_3636);
nor U9852 (N_9852,N_83,N_3729);
nor U9853 (N_9853,N_4733,N_2265);
nor U9854 (N_9854,N_1065,N_2119);
nand U9855 (N_9855,N_3908,N_1963);
nand U9856 (N_9856,N_1032,N_3522);
and U9857 (N_9857,N_3763,N_3063);
nor U9858 (N_9858,N_2202,N_1952);
or U9859 (N_9859,N_3552,N_3612);
and U9860 (N_9860,N_3766,N_2176);
and U9861 (N_9861,N_997,N_287);
nand U9862 (N_9862,N_147,N_1493);
and U9863 (N_9863,N_844,N_867);
or U9864 (N_9864,N_2722,N_1823);
xor U9865 (N_9865,N_689,N_4509);
or U9866 (N_9866,N_1076,N_976);
or U9867 (N_9867,N_2532,N_3013);
xor U9868 (N_9868,N_4138,N_433);
nand U9869 (N_9869,N_679,N_4108);
xnor U9870 (N_9870,N_4132,N_2050);
nor U9871 (N_9871,N_1119,N_2280);
or U9872 (N_9872,N_2387,N_1872);
xnor U9873 (N_9873,N_2124,N_3343);
nor U9874 (N_9874,N_115,N_3850);
nor U9875 (N_9875,N_2446,N_759);
nor U9876 (N_9876,N_325,N_243);
nor U9877 (N_9877,N_1754,N_1751);
nand U9878 (N_9878,N_4422,N_2473);
nor U9879 (N_9879,N_479,N_1904);
and U9880 (N_9880,N_3660,N_384);
xnor U9881 (N_9881,N_2621,N_2511);
and U9882 (N_9882,N_629,N_4720);
and U9883 (N_9883,N_4756,N_4380);
nand U9884 (N_9884,N_1504,N_3);
xor U9885 (N_9885,N_4294,N_551);
or U9886 (N_9886,N_1793,N_172);
or U9887 (N_9887,N_4795,N_4550);
nand U9888 (N_9888,N_2396,N_4701);
nor U9889 (N_9889,N_177,N_111);
xnor U9890 (N_9890,N_3647,N_3399);
nand U9891 (N_9891,N_1674,N_2839);
nand U9892 (N_9892,N_1702,N_1937);
xor U9893 (N_9893,N_1983,N_1389);
xor U9894 (N_9894,N_3765,N_127);
nor U9895 (N_9895,N_2010,N_1169);
nand U9896 (N_9896,N_3302,N_1902);
and U9897 (N_9897,N_2183,N_2947);
or U9898 (N_9898,N_3697,N_4497);
or U9899 (N_9899,N_565,N_2110);
and U9900 (N_9900,N_2312,N_1936);
xor U9901 (N_9901,N_2713,N_4382);
nand U9902 (N_9902,N_503,N_2641);
xor U9903 (N_9903,N_922,N_3099);
and U9904 (N_9904,N_2943,N_4863);
nor U9905 (N_9905,N_4034,N_376);
xnor U9906 (N_9906,N_3765,N_1748);
nor U9907 (N_9907,N_3666,N_3232);
and U9908 (N_9908,N_3566,N_4004);
and U9909 (N_9909,N_4599,N_3674);
nand U9910 (N_9910,N_2930,N_1782);
and U9911 (N_9911,N_1093,N_4005);
or U9912 (N_9912,N_761,N_4087);
nand U9913 (N_9913,N_4917,N_1069);
nor U9914 (N_9914,N_4114,N_4653);
nor U9915 (N_9915,N_4039,N_3794);
and U9916 (N_9916,N_2812,N_1963);
or U9917 (N_9917,N_4221,N_3092);
xor U9918 (N_9918,N_4498,N_1007);
or U9919 (N_9919,N_1691,N_254);
or U9920 (N_9920,N_308,N_2584);
or U9921 (N_9921,N_2341,N_4903);
or U9922 (N_9922,N_1635,N_4251);
and U9923 (N_9923,N_2563,N_475);
nor U9924 (N_9924,N_4649,N_850);
and U9925 (N_9925,N_4259,N_1012);
xor U9926 (N_9926,N_275,N_2550);
xor U9927 (N_9927,N_562,N_3165);
xnor U9928 (N_9928,N_2855,N_2805);
and U9929 (N_9929,N_3683,N_2954);
xor U9930 (N_9930,N_1981,N_4633);
nand U9931 (N_9931,N_1552,N_4479);
nor U9932 (N_9932,N_1293,N_2549);
nor U9933 (N_9933,N_4208,N_4205);
nor U9934 (N_9934,N_4609,N_1523);
nand U9935 (N_9935,N_3351,N_1720);
and U9936 (N_9936,N_3576,N_3182);
and U9937 (N_9937,N_4938,N_4890);
nor U9938 (N_9938,N_1373,N_2553);
and U9939 (N_9939,N_3250,N_4013);
and U9940 (N_9940,N_2071,N_4628);
and U9941 (N_9941,N_4379,N_1157);
and U9942 (N_9942,N_2972,N_3184);
and U9943 (N_9943,N_4635,N_1567);
and U9944 (N_9944,N_82,N_1873);
xnor U9945 (N_9945,N_2521,N_4817);
xnor U9946 (N_9946,N_4022,N_219);
or U9947 (N_9947,N_166,N_2241);
and U9948 (N_9948,N_668,N_785);
xnor U9949 (N_9949,N_444,N_3598);
and U9950 (N_9950,N_4612,N_4992);
xnor U9951 (N_9951,N_3104,N_4011);
or U9952 (N_9952,N_4902,N_1913);
and U9953 (N_9953,N_4681,N_3065);
xor U9954 (N_9954,N_146,N_1849);
nor U9955 (N_9955,N_3707,N_1252);
nor U9956 (N_9956,N_4127,N_4950);
or U9957 (N_9957,N_1254,N_1336);
and U9958 (N_9958,N_152,N_3665);
nand U9959 (N_9959,N_1173,N_2181);
nand U9960 (N_9960,N_2241,N_3966);
nor U9961 (N_9961,N_1251,N_4650);
xor U9962 (N_9962,N_2391,N_4532);
and U9963 (N_9963,N_2654,N_3376);
and U9964 (N_9964,N_464,N_2087);
nor U9965 (N_9965,N_1587,N_970);
and U9966 (N_9966,N_615,N_44);
nor U9967 (N_9967,N_489,N_1622);
nand U9968 (N_9968,N_2662,N_2177);
nand U9969 (N_9969,N_2318,N_4864);
nand U9970 (N_9970,N_2343,N_2634);
xnor U9971 (N_9971,N_3086,N_514);
nor U9972 (N_9972,N_3695,N_4879);
nor U9973 (N_9973,N_1901,N_2308);
or U9974 (N_9974,N_3380,N_2958);
nor U9975 (N_9975,N_1942,N_1994);
nor U9976 (N_9976,N_1508,N_4567);
and U9977 (N_9977,N_309,N_2436);
nand U9978 (N_9978,N_1455,N_856);
or U9979 (N_9979,N_74,N_4987);
or U9980 (N_9980,N_4710,N_1299);
nor U9981 (N_9981,N_1755,N_1797);
or U9982 (N_9982,N_2453,N_2459);
nor U9983 (N_9983,N_730,N_2885);
nor U9984 (N_9984,N_3300,N_771);
xor U9985 (N_9985,N_3250,N_4633);
nand U9986 (N_9986,N_2395,N_797);
and U9987 (N_9987,N_3589,N_2203);
xor U9988 (N_9988,N_3145,N_642);
and U9989 (N_9989,N_4613,N_4135);
or U9990 (N_9990,N_2669,N_4589);
nand U9991 (N_9991,N_2857,N_678);
xnor U9992 (N_9992,N_1765,N_2429);
nor U9993 (N_9993,N_1319,N_4043);
and U9994 (N_9994,N_1082,N_3997);
and U9995 (N_9995,N_1228,N_4026);
nor U9996 (N_9996,N_120,N_4034);
and U9997 (N_9997,N_3851,N_840);
or U9998 (N_9998,N_2966,N_4246);
or U9999 (N_9999,N_122,N_1199);
nor U10000 (N_10000,N_8096,N_8297);
and U10001 (N_10001,N_9198,N_7644);
and U10002 (N_10002,N_9739,N_9842);
nand U10003 (N_10003,N_9599,N_8550);
nor U10004 (N_10004,N_7535,N_7160);
nand U10005 (N_10005,N_9833,N_8959);
or U10006 (N_10006,N_5054,N_5042);
xnor U10007 (N_10007,N_5929,N_6137);
xnor U10008 (N_10008,N_5138,N_6868);
nor U10009 (N_10009,N_9377,N_6419);
xnor U10010 (N_10010,N_9341,N_7309);
nand U10011 (N_10011,N_5649,N_7020);
or U10012 (N_10012,N_7257,N_6912);
nand U10013 (N_10013,N_6220,N_8926);
nand U10014 (N_10014,N_9935,N_6946);
xor U10015 (N_10015,N_5920,N_5513);
nand U10016 (N_10016,N_5095,N_8692);
nor U10017 (N_10017,N_7960,N_5029);
nor U10018 (N_10018,N_5990,N_6064);
nand U10019 (N_10019,N_9468,N_7650);
nor U10020 (N_10020,N_6654,N_9572);
nor U10021 (N_10021,N_6798,N_7864);
nor U10022 (N_10022,N_5177,N_9230);
xor U10023 (N_10023,N_6254,N_8325);
and U10024 (N_10024,N_5001,N_7948);
xor U10025 (N_10025,N_7396,N_8215);
nor U10026 (N_10026,N_6745,N_7176);
nand U10027 (N_10027,N_6392,N_7943);
nor U10028 (N_10028,N_5952,N_6151);
or U10029 (N_10029,N_7800,N_9699);
xor U10030 (N_10030,N_5201,N_8431);
nand U10031 (N_10031,N_9964,N_6205);
nand U10032 (N_10032,N_8988,N_7829);
and U10033 (N_10033,N_9414,N_5287);
nand U10034 (N_10034,N_9937,N_9413);
xnor U10035 (N_10035,N_5324,N_9531);
nand U10036 (N_10036,N_9322,N_7271);
nor U10037 (N_10037,N_9149,N_8985);
xor U10038 (N_10038,N_9951,N_7277);
nor U10039 (N_10039,N_8013,N_7456);
xnor U10040 (N_10040,N_8420,N_5101);
or U10041 (N_10041,N_6449,N_6674);
and U10042 (N_10042,N_8669,N_6863);
nor U10043 (N_10043,N_6425,N_5963);
and U10044 (N_10044,N_5310,N_5272);
and U10045 (N_10045,N_8974,N_6832);
nand U10046 (N_10046,N_6242,N_8544);
and U10047 (N_10047,N_8484,N_9484);
and U10048 (N_10048,N_8520,N_5150);
or U10049 (N_10049,N_7006,N_9718);
and U10050 (N_10050,N_8630,N_9002);
or U10051 (N_10051,N_6129,N_5006);
nand U10052 (N_10052,N_8425,N_9271);
or U10053 (N_10053,N_8643,N_7435);
and U10054 (N_10054,N_9005,N_9985);
nor U10055 (N_10055,N_8745,N_5947);
nand U10056 (N_10056,N_8180,N_5521);
xnor U10057 (N_10057,N_5615,N_6616);
or U10058 (N_10058,N_9009,N_9034);
nor U10059 (N_10059,N_9956,N_5240);
and U10060 (N_10060,N_5664,N_5304);
xnor U10061 (N_10061,N_9229,N_6368);
and U10062 (N_10062,N_8638,N_8913);
xor U10063 (N_10063,N_8558,N_7298);
xnor U10064 (N_10064,N_5793,N_5917);
or U10065 (N_10065,N_6700,N_5779);
xnor U10066 (N_10066,N_8277,N_7091);
nor U10067 (N_10067,N_6742,N_5005);
and U10068 (N_10068,N_9757,N_8562);
nand U10069 (N_10069,N_6640,N_7621);
nand U10070 (N_10070,N_9061,N_6145);
nand U10071 (N_10071,N_7063,N_8035);
nand U10072 (N_10072,N_5209,N_9140);
or U10073 (N_10073,N_9633,N_6716);
and U10074 (N_10074,N_5506,N_8938);
xor U10075 (N_10075,N_6057,N_5372);
nand U10076 (N_10076,N_7686,N_6202);
nor U10077 (N_10077,N_5192,N_6572);
nand U10078 (N_10078,N_5485,N_6394);
or U10079 (N_10079,N_7178,N_9277);
nor U10080 (N_10080,N_9037,N_5489);
nor U10081 (N_10081,N_7842,N_7598);
and U10082 (N_10082,N_6929,N_9035);
nand U10083 (N_10083,N_6257,N_7990);
nor U10084 (N_10084,N_5044,N_6289);
nor U10085 (N_10085,N_9696,N_5910);
or U10086 (N_10086,N_9418,N_5741);
and U10087 (N_10087,N_7744,N_6653);
and U10088 (N_10088,N_8504,N_7515);
or U10089 (N_10089,N_8012,N_5366);
or U10090 (N_10090,N_7014,N_7916);
nand U10091 (N_10091,N_5239,N_7734);
nand U10092 (N_10092,N_8709,N_6731);
and U10093 (N_10093,N_8819,N_8691);
or U10094 (N_10094,N_6917,N_6315);
nand U10095 (N_10095,N_9378,N_7290);
nand U10096 (N_10096,N_7081,N_7693);
and U10097 (N_10097,N_6194,N_6577);
xor U10098 (N_10098,N_8730,N_5255);
nor U10099 (N_10099,N_8775,N_9219);
and U10100 (N_10100,N_8127,N_7062);
nor U10101 (N_10101,N_8972,N_9383);
or U10102 (N_10102,N_6104,N_5801);
nand U10103 (N_10103,N_8479,N_6106);
xor U10104 (N_10104,N_9578,N_9285);
or U10105 (N_10105,N_9183,N_9530);
xor U10106 (N_10106,N_8905,N_7614);
xnor U10107 (N_10107,N_7626,N_8169);
xnor U10108 (N_10108,N_5979,N_9952);
nor U10109 (N_10109,N_8024,N_8718);
nor U10110 (N_10110,N_9128,N_6432);
xnor U10111 (N_10111,N_5724,N_8073);
nand U10112 (N_10112,N_8859,N_9724);
and U10113 (N_10113,N_8700,N_8351);
xnor U10114 (N_10114,N_5523,N_8327);
and U10115 (N_10115,N_9697,N_7319);
or U10116 (N_10116,N_9958,N_9591);
nand U10117 (N_10117,N_7170,N_6322);
and U10118 (N_10118,N_6045,N_8057);
or U10119 (N_10119,N_6418,N_8538);
nor U10120 (N_10120,N_9488,N_6527);
and U10121 (N_10121,N_9154,N_8768);
or U10122 (N_10122,N_8921,N_7712);
xor U10123 (N_10123,N_9018,N_9090);
nor U10124 (N_10124,N_7600,N_7302);
xor U10125 (N_10125,N_5644,N_6559);
xnor U10126 (N_10126,N_5866,N_7975);
or U10127 (N_10127,N_6113,N_6105);
nand U10128 (N_10128,N_6316,N_8069);
or U10129 (N_10129,N_7871,N_5079);
and U10130 (N_10130,N_7415,N_8660);
and U10131 (N_10131,N_7635,N_7487);
nor U10132 (N_10132,N_8023,N_8843);
xor U10133 (N_10133,N_6152,N_5211);
nor U10134 (N_10134,N_6850,N_7323);
or U10135 (N_10135,N_6567,N_6496);
nor U10136 (N_10136,N_6818,N_5157);
and U10137 (N_10137,N_8901,N_7446);
nand U10138 (N_10138,N_7459,N_5110);
nor U10139 (N_10139,N_7304,N_5625);
xor U10140 (N_10140,N_6763,N_9924);
nor U10141 (N_10141,N_8152,N_6372);
or U10142 (N_10142,N_6177,N_9839);
nor U10143 (N_10143,N_6204,N_9595);
xnor U10144 (N_10144,N_8195,N_7776);
xnor U10145 (N_10145,N_6494,N_5322);
or U10146 (N_10146,N_6748,N_5752);
nand U10147 (N_10147,N_5817,N_7254);
xnor U10148 (N_10148,N_5340,N_9917);
xor U10149 (N_10149,N_7389,N_9922);
and U10150 (N_10150,N_7291,N_9071);
nand U10151 (N_10151,N_9346,N_8375);
nor U10152 (N_10152,N_9016,N_5773);
xor U10153 (N_10153,N_6846,N_9225);
and U10154 (N_10154,N_8248,N_7008);
or U10155 (N_10155,N_7153,N_6490);
nor U10156 (N_10156,N_6085,N_7763);
xor U10157 (N_10157,N_6050,N_8551);
or U10158 (N_10158,N_5934,N_5977);
nand U10159 (N_10159,N_9705,N_8072);
or U10160 (N_10160,N_8896,N_5700);
nor U10161 (N_10161,N_9355,N_5417);
nand U10162 (N_10162,N_8486,N_8311);
and U10163 (N_10163,N_6142,N_8089);
or U10164 (N_10164,N_7995,N_6150);
xor U10165 (N_10165,N_6859,N_5620);
and U10166 (N_10166,N_5124,N_7764);
and U10167 (N_10167,N_6463,N_6968);
nor U10168 (N_10168,N_8377,N_6361);
xnor U10169 (N_10169,N_9182,N_7993);
nand U10170 (N_10170,N_9542,N_5422);
nand U10171 (N_10171,N_9084,N_7998);
nor U10172 (N_10172,N_6634,N_6026);
and U10173 (N_10173,N_8061,N_6061);
nor U10174 (N_10174,N_8742,N_9695);
nor U10175 (N_10175,N_6582,N_5196);
or U10176 (N_10176,N_8727,N_7834);
and U10177 (N_10177,N_7891,N_7608);
xnor U10178 (N_10178,N_5305,N_9963);
nand U10179 (N_10179,N_5348,N_6979);
and U10180 (N_10180,N_8744,N_7582);
or U10181 (N_10181,N_5659,N_5732);
nor U10182 (N_10182,N_6556,N_6816);
and U10183 (N_10183,N_8565,N_6510);
and U10184 (N_10184,N_6560,N_9682);
or U10185 (N_10185,N_6153,N_8365);
and U10186 (N_10186,N_6858,N_5785);
and U10187 (N_10187,N_6771,N_7168);
nand U10188 (N_10188,N_6903,N_8508);
and U10189 (N_10189,N_7468,N_9123);
or U10190 (N_10190,N_6423,N_6337);
nand U10191 (N_10191,N_7620,N_5195);
nand U10192 (N_10192,N_9385,N_5872);
or U10193 (N_10193,N_8689,N_7550);
nor U10194 (N_10194,N_9957,N_7890);
xnor U10195 (N_10195,N_6787,N_7991);
xnor U10196 (N_10196,N_8029,N_9515);
nand U10197 (N_10197,N_8624,N_6678);
xor U10198 (N_10198,N_9000,N_8791);
or U10199 (N_10199,N_8392,N_9597);
nand U10200 (N_10200,N_9946,N_6893);
nor U10201 (N_10201,N_9487,N_9867);
nand U10202 (N_10202,N_7407,N_7833);
nand U10203 (N_10203,N_7966,N_5944);
or U10204 (N_10204,N_5337,N_7819);
or U10205 (N_10205,N_8289,N_5269);
nand U10206 (N_10206,N_8906,N_5013);
nor U10207 (N_10207,N_6226,N_6428);
or U10208 (N_10208,N_9081,N_9345);
xor U10209 (N_10209,N_8793,N_7606);
and U10210 (N_10210,N_9527,N_6797);
or U10211 (N_10211,N_8561,N_5574);
nand U10212 (N_10212,N_5321,N_6112);
or U10213 (N_10213,N_7882,N_6073);
and U10214 (N_10214,N_6053,N_9437);
nor U10215 (N_10215,N_7034,N_5015);
and U10216 (N_10216,N_5887,N_5774);
nand U10217 (N_10217,N_7884,N_7426);
xnor U10218 (N_10218,N_7245,N_9897);
or U10219 (N_10219,N_7520,N_5378);
nor U10220 (N_10220,N_7959,N_8134);
nor U10221 (N_10221,N_8296,N_9478);
xor U10222 (N_10222,N_9275,N_6525);
or U10223 (N_10223,N_7240,N_6707);
xnor U10224 (N_10224,N_6025,N_8903);
or U10225 (N_10225,N_6982,N_9569);
xor U10226 (N_10226,N_9805,N_6318);
or U10227 (N_10227,N_7317,N_6051);
nand U10228 (N_10228,N_6348,N_7102);
nor U10229 (N_10229,N_6002,N_9004);
nor U10230 (N_10230,N_5745,N_5263);
or U10231 (N_10231,N_7641,N_9232);
nor U10232 (N_10232,N_8795,N_8383);
or U10233 (N_10233,N_7911,N_6238);
nor U10234 (N_10234,N_5188,N_8402);
nand U10235 (N_10235,N_9169,N_7156);
nor U10236 (N_10236,N_6028,N_8876);
or U10237 (N_10237,N_9580,N_8036);
and U10238 (N_10238,N_9774,N_5014);
xnor U10239 (N_10239,N_8338,N_9499);
nor U10240 (N_10240,N_7836,N_7397);
and U10241 (N_10241,N_7775,N_8542);
xnor U10242 (N_10242,N_8199,N_6311);
and U10243 (N_10243,N_9312,N_8173);
nand U10244 (N_10244,N_6273,N_6340);
or U10245 (N_10245,N_5469,N_8320);
xor U10246 (N_10246,N_6324,N_8713);
nor U10247 (N_10247,N_7767,N_7611);
and U10248 (N_10248,N_8919,N_8010);
nor U10249 (N_10249,N_7452,N_6649);
and U10250 (N_10250,N_5345,N_8715);
or U10251 (N_10251,N_5257,N_5915);
nand U10252 (N_10252,N_7703,N_5077);
and U10253 (N_10253,N_7726,N_9574);
nor U10254 (N_10254,N_5679,N_7771);
nand U10255 (N_10255,N_6648,N_8039);
nor U10256 (N_10256,N_9282,N_7258);
or U10257 (N_10257,N_6391,N_9047);
and U10258 (N_10258,N_6139,N_7722);
or U10259 (N_10259,N_9781,N_7964);
or U10260 (N_10260,N_6079,N_9814);
nand U10261 (N_10261,N_5039,N_8231);
and U10262 (N_10262,N_6970,N_5285);
and U10263 (N_10263,N_5733,N_6939);
nand U10264 (N_10264,N_9129,N_5823);
and U10265 (N_10265,N_9589,N_8917);
and U10266 (N_10266,N_8610,N_5181);
nand U10267 (N_10267,N_9191,N_9262);
xnor U10268 (N_10268,N_7144,N_7560);
xor U10269 (N_10269,N_5657,N_6455);
and U10270 (N_10270,N_7559,N_6218);
nand U10271 (N_10271,N_9801,N_5692);
and U10272 (N_10272,N_6453,N_5302);
nor U10273 (N_10273,N_9729,N_7066);
nor U10274 (N_10274,N_5671,N_9222);
nor U10275 (N_10275,N_6692,N_5163);
or U10276 (N_10276,N_9715,N_7113);
nor U10277 (N_10277,N_7795,N_6937);
and U10278 (N_10278,N_9541,N_8342);
and U10279 (N_10279,N_9110,N_6127);
and U10280 (N_10280,N_5935,N_6883);
nor U10281 (N_10281,N_7162,N_6346);
and U10282 (N_10282,N_6377,N_9506);
nor U10283 (N_10283,N_8279,N_9280);
xnor U10284 (N_10284,N_9480,N_7401);
and U10285 (N_10285,N_7813,N_8858);
nand U10286 (N_10286,N_5284,N_7280);
nor U10287 (N_10287,N_9051,N_9315);
xor U10288 (N_10288,N_9775,N_9650);
xor U10289 (N_10289,N_7430,N_6784);
nand U10290 (N_10290,N_7080,N_7869);
or U10291 (N_10291,N_6591,N_7876);
nor U10292 (N_10292,N_7649,N_5590);
xnor U10293 (N_10293,N_5207,N_9142);
xnor U10294 (N_10294,N_6248,N_7896);
xor U10295 (N_10295,N_7410,N_5791);
nand U10296 (N_10296,N_7222,N_7075);
xor U10297 (N_10297,N_7759,N_8577);
and U10298 (N_10298,N_7194,N_5000);
and U10299 (N_10299,N_9773,N_7538);
xor U10300 (N_10300,N_6600,N_9932);
nand U10301 (N_10301,N_7749,N_9570);
xnor U10302 (N_10302,N_9253,N_9927);
nand U10303 (N_10303,N_9422,N_9745);
and U10304 (N_10304,N_9294,N_9746);
nor U10305 (N_10305,N_9099,N_5580);
or U10306 (N_10306,N_9658,N_5190);
nor U10307 (N_10307,N_7227,N_6972);
and U10308 (N_10308,N_9489,N_8712);
xnor U10309 (N_10309,N_7847,N_8763);
xor U10310 (N_10310,N_5125,N_7088);
and U10311 (N_10311,N_6872,N_7601);
and U10312 (N_10312,N_6470,N_7669);
or U10313 (N_10313,N_6468,N_8841);
and U10314 (N_10314,N_9333,N_5879);
nand U10315 (N_10315,N_7332,N_8470);
and U10316 (N_10316,N_7566,N_9211);
or U10317 (N_10317,N_7129,N_6799);
or U10318 (N_10318,N_6536,N_7053);
xnor U10319 (N_10319,N_5666,N_8453);
or U10320 (N_10320,N_7574,N_7778);
or U10321 (N_10321,N_9108,N_9614);
nor U10322 (N_10322,N_7355,N_9810);
nand U10323 (N_10323,N_8506,N_8942);
or U10324 (N_10324,N_9868,N_9025);
nand U10325 (N_10325,N_8051,N_6495);
nor U10326 (N_10326,N_6301,N_5156);
or U10327 (N_10327,N_5706,N_8464);
or U10328 (N_10328,N_7903,N_8958);
nor U10329 (N_10329,N_5481,N_7307);
nand U10330 (N_10330,N_8009,N_8509);
xor U10331 (N_10331,N_9670,N_6664);
xnor U10332 (N_10332,N_7682,N_6158);
or U10333 (N_10333,N_6758,N_8754);
xnor U10334 (N_10334,N_5460,N_6269);
xnor U10335 (N_10335,N_6733,N_9258);
xor U10336 (N_10336,N_7447,N_7656);
nand U10337 (N_10337,N_8167,N_8295);
nand U10338 (N_10338,N_8908,N_5600);
nor U10339 (N_10339,N_6222,N_7138);
nand U10340 (N_10340,N_9238,N_7386);
nand U10341 (N_10341,N_7770,N_9425);
nor U10342 (N_10342,N_5056,N_8871);
xnor U10343 (N_10343,N_9159,N_6213);
nor U10344 (N_10344,N_6189,N_9762);
and U10345 (N_10345,N_6909,N_6895);
nor U10346 (N_10346,N_7612,N_6545);
and U10347 (N_10347,N_5122,N_6951);
or U10348 (N_10348,N_9862,N_9357);
nand U10349 (N_10349,N_8306,N_8976);
nand U10350 (N_10350,N_9244,N_6302);
nor U10351 (N_10351,N_9075,N_8068);
nor U10352 (N_10352,N_5820,N_9539);
nand U10353 (N_10353,N_8547,N_5547);
and U10354 (N_10354,N_6041,N_9701);
and U10355 (N_10355,N_8397,N_7076);
and U10356 (N_10356,N_7195,N_9826);
nand U10357 (N_10357,N_8825,N_5711);
nand U10358 (N_10358,N_9903,N_8198);
nor U10359 (N_10359,N_7630,N_7275);
nor U10360 (N_10360,N_6842,N_7248);
nand U10361 (N_10361,N_6056,N_7269);
nor U10362 (N_10362,N_8501,N_5584);
and U10363 (N_10363,N_7753,N_8472);
nor U10364 (N_10364,N_5396,N_9406);
or U10365 (N_10365,N_9206,N_6224);
xor U10366 (N_10366,N_5176,N_7278);
nand U10367 (N_10367,N_8326,N_6760);
nor U10368 (N_10368,N_9509,N_8851);
and U10369 (N_10369,N_8185,N_8787);
and U10370 (N_10370,N_8609,N_7958);
and U10371 (N_10371,N_9237,N_9331);
and U10372 (N_10372,N_6702,N_5282);
and U10373 (N_10373,N_8373,N_7537);
nor U10374 (N_10374,N_9470,N_6303);
nor U10375 (N_10375,N_5888,N_9021);
nand U10376 (N_10376,N_5640,N_9843);
or U10377 (N_10377,N_9521,N_9223);
or U10378 (N_10378,N_8150,N_5402);
and U10379 (N_10379,N_5058,N_9716);
nand U10380 (N_10380,N_8681,N_7521);
nand U10381 (N_10381,N_6483,N_9390);
nor U10382 (N_10382,N_7161,N_5486);
nand U10383 (N_10383,N_6570,N_9571);
nand U10384 (N_10384,N_9813,N_9749);
nor U10385 (N_10385,N_8019,N_9150);
xnor U10386 (N_10386,N_9319,N_9038);
nor U10387 (N_10387,N_7547,N_6888);
nor U10388 (N_10388,N_6331,N_9343);
and U10389 (N_10389,N_7653,N_6395);
and U10390 (N_10390,N_7181,N_9665);
nor U10391 (N_10391,N_9027,N_6004);
nand U10392 (N_10392,N_5464,N_6091);
nor U10393 (N_10393,N_9329,N_5650);
and U10394 (N_10394,N_8154,N_7617);
nor U10395 (N_10395,N_6170,N_9712);
or U10396 (N_10396,N_6610,N_5877);
nor U10397 (N_10397,N_9876,N_6550);
nand U10398 (N_10398,N_7388,N_6681);
nor U10399 (N_10399,N_5946,N_9153);
and U10400 (N_10400,N_8418,N_5660);
nand U10401 (N_10401,N_5716,N_9247);
or U10402 (N_10402,N_6407,N_9114);
or U10403 (N_10403,N_9330,N_8194);
and U10404 (N_10404,N_5012,N_9864);
nor U10405 (N_10405,N_5844,N_6845);
or U10406 (N_10406,N_8065,N_9395);
xnor U10407 (N_10407,N_7544,N_8507);
and U10408 (N_10408,N_6499,N_7673);
nor U10409 (N_10409,N_9994,N_5045);
nor U10410 (N_10410,N_8478,N_8641);
nand U10411 (N_10411,N_8552,N_5379);
and U10412 (N_10412,N_6985,N_6534);
nor U10413 (N_10413,N_5592,N_6978);
nand U10414 (N_10414,N_8640,N_8469);
or U10415 (N_10415,N_7820,N_7804);
nor U10416 (N_10416,N_7470,N_6304);
nor U10417 (N_10417,N_5373,N_6141);
xnor U10418 (N_10418,N_9006,N_8126);
nor U10419 (N_10419,N_5756,N_6877);
nor U10420 (N_10420,N_6628,N_8725);
nand U10421 (N_10421,N_7992,N_8576);
nor U10422 (N_10422,N_7143,N_5748);
or U10423 (N_10423,N_7745,N_6245);
nand U10424 (N_10424,N_8879,N_5669);
nor U10425 (N_10425,N_9832,N_7262);
nand U10426 (N_10426,N_6469,N_7368);
nor U10427 (N_10427,N_9296,N_8457);
and U10428 (N_10428,N_7562,N_5404);
nor U10429 (N_10429,N_8444,N_7888);
xnor U10430 (N_10430,N_8933,N_9190);
nor U10431 (N_10431,N_6360,N_6488);
nor U10432 (N_10432,N_7904,N_5758);
xnor U10433 (N_10433,N_9646,N_8502);
nand U10434 (N_10434,N_8189,N_8695);
nor U10435 (N_10435,N_8849,N_8541);
nand U10436 (N_10436,N_6861,N_9185);
nand U10437 (N_10437,N_7223,N_5298);
nand U10438 (N_10438,N_5374,N_5071);
or U10439 (N_10439,N_7528,N_6711);
nor U10440 (N_10440,N_8534,N_9420);
nor U10441 (N_10441,N_5290,N_6624);
nor U10442 (N_10442,N_8158,N_5767);
nand U10443 (N_10443,N_8894,N_6677);
nor U10444 (N_10444,N_9399,N_9626);
nor U10445 (N_10445,N_9988,N_8644);
nand U10446 (N_10446,N_8612,N_8485);
xnor U10447 (N_10447,N_8042,N_9717);
or U10448 (N_10448,N_6867,N_7482);
xor U10449 (N_10449,N_9885,N_7228);
or U10450 (N_10450,N_7343,N_8855);
or U10451 (N_10451,N_5160,N_8663);
or U10452 (N_10452,N_7706,N_7367);
nand U10453 (N_10453,N_7557,N_6708);
nand U10454 (N_10454,N_6427,N_6699);
nand U10455 (N_10455,N_5693,N_7879);
and U10456 (N_10456,N_8814,N_8053);
xor U10457 (N_10457,N_8877,N_5972);
xnor U10458 (N_10458,N_7377,N_6014);
nand U10459 (N_10459,N_6879,N_8468);
and U10460 (N_10460,N_6336,N_9264);
and U10461 (N_10461,N_9836,N_6905);
xor U10462 (N_10462,N_8521,N_9251);
nor U10463 (N_10463,N_9165,N_9560);
nand U10464 (N_10464,N_8001,N_8459);
or U10465 (N_10465,N_6990,N_6179);
nand U10466 (N_10466,N_6706,N_7233);
nand U10467 (N_10467,N_7460,N_5841);
or U10468 (N_10468,N_5334,N_9293);
nor U10469 (N_10469,N_5357,N_5041);
nor U10470 (N_10470,N_9166,N_8466);
nor U10471 (N_10471,N_9608,N_6434);
and U10472 (N_10472,N_6575,N_9848);
xor U10473 (N_10473,N_9397,N_5661);
nor U10474 (N_10474,N_5397,N_7963);
nor U10475 (N_10475,N_7524,N_7512);
or U10476 (N_10476,N_8266,N_7112);
nor U10477 (N_10477,N_5870,N_7919);
xor U10478 (N_10478,N_9783,N_8137);
and U10479 (N_10479,N_9620,N_8164);
nor U10480 (N_10480,N_5968,N_6639);
nor U10481 (N_10481,N_6590,N_7180);
nor U10482 (N_10482,N_6751,N_6622);
and U10483 (N_10483,N_7742,N_8621);
or U10484 (N_10484,N_6436,N_6408);
nor U10485 (N_10485,N_6857,N_5094);
nor U10486 (N_10486,N_5172,N_5320);
nor U10487 (N_10487,N_6197,N_9112);
xor U10488 (N_10488,N_9637,N_8586);
xor U10489 (N_10489,N_6107,N_6251);
nand U10490 (N_10490,N_7725,N_8625);
and U10491 (N_10491,N_7675,N_6523);
xnor U10492 (N_10492,N_8614,N_7321);
or U10493 (N_10493,N_5368,N_5258);
nor U10494 (N_10494,N_9217,N_5864);
and U10495 (N_10495,N_9485,N_6344);
nor U10496 (N_10496,N_5007,N_9849);
or U10497 (N_10497,N_8344,N_6843);
or U10498 (N_10498,N_5818,N_6612);
xnor U10499 (N_10499,N_7352,N_6435);
xnor U10500 (N_10500,N_8087,N_7501);
nor U10501 (N_10501,N_8493,N_9243);
nor U10502 (N_10502,N_7818,N_7167);
and U10503 (N_10503,N_8671,N_9700);
nor U10504 (N_10504,N_8109,N_7625);
and U10505 (N_10505,N_7652,N_5468);
xor U10506 (N_10506,N_9962,N_6999);
xor U10507 (N_10507,N_9339,N_7431);
nand U10508 (N_10508,N_8531,N_7106);
and U10509 (N_10509,N_8267,N_6080);
and U10510 (N_10510,N_8208,N_8655);
or U10511 (N_10511,N_9146,N_9281);
or U10512 (N_10512,N_6767,N_5558);
xor U10513 (N_10513,N_7107,N_7824);
nand U10514 (N_10514,N_7509,N_7433);
and U10515 (N_10515,N_8462,N_8082);
xor U10516 (N_10516,N_5674,N_6446);
xnor U10517 (N_10517,N_8362,N_6086);
or U10518 (N_10518,N_9995,N_6549);
nor U10519 (N_10519,N_8622,N_5410);
or U10520 (N_10520,N_5822,N_6504);
nand U10521 (N_10521,N_5147,N_8888);
nand U10522 (N_10522,N_6657,N_9629);
nand U10523 (N_10523,N_8423,N_9960);
nand U10524 (N_10524,N_9226,N_6313);
xor U10525 (N_10525,N_8105,N_6393);
or U10526 (N_10526,N_5222,N_8390);
xor U10527 (N_10527,N_7555,N_5136);
nor U10528 (N_10528,N_6960,N_8143);
xnor U10529 (N_10529,N_9544,N_9070);
and U10530 (N_10530,N_7184,N_6363);
nor U10531 (N_10531,N_6460,N_9501);
or U10532 (N_10532,N_8230,N_9981);
nand U10533 (N_10533,N_9577,N_9847);
nand U10534 (N_10534,N_6035,N_7956);
nor U10535 (N_10535,N_6529,N_8074);
and U10536 (N_10536,N_6796,N_9122);
nor U10537 (N_10537,N_8247,N_5699);
and U10538 (N_10538,N_8834,N_6431);
xnor U10539 (N_10539,N_7880,N_8719);
xnor U10540 (N_10540,N_9250,N_6566);
and U10541 (N_10541,N_6696,N_9164);
nand U10542 (N_10542,N_5279,N_5966);
nand U10543 (N_10543,N_8460,N_7255);
xnor U10544 (N_10544,N_8037,N_5663);
or U10545 (N_10545,N_9064,N_5882);
and U10546 (N_10546,N_7001,N_6356);
and U10547 (N_10547,N_5548,N_9055);
nand U10548 (N_10548,N_7357,N_6038);
or U10549 (N_10549,N_5965,N_8439);
xor U10550 (N_10550,N_7187,N_8887);
nand U10551 (N_10551,N_5245,N_9708);
xnor U10552 (N_10552,N_8401,N_9893);
and U10553 (N_10553,N_9852,N_7704);
and U10554 (N_10554,N_6530,N_5052);
nor U10555 (N_10555,N_6070,N_6598);
nand U10556 (N_10556,N_6548,N_7865);
nor U10557 (N_10557,N_9207,N_6975);
and U10558 (N_10558,N_9661,N_5243);
nor U10559 (N_10559,N_8251,N_8437);
or U10560 (N_10560,N_9575,N_9835);
nor U10561 (N_10561,N_5763,N_9940);
nand U10562 (N_10562,N_7905,N_5677);
xor U10563 (N_10563,N_5593,N_8571);
nor U10564 (N_10564,N_8907,N_7422);
nand U10565 (N_10565,N_6997,N_6558);
nor U10566 (N_10566,N_9491,N_7531);
or U10567 (N_10567,N_6701,N_5876);
nand U10568 (N_10568,N_6310,N_8801);
and U10569 (N_10569,N_6643,N_8234);
and U10570 (N_10570,N_6186,N_7640);
nand U10571 (N_10571,N_8852,N_7940);
xor U10572 (N_10572,N_7079,N_5339);
and U10573 (N_10573,N_9187,N_8161);
xor U10574 (N_10574,N_7755,N_5206);
nor U10575 (N_10575,N_8818,N_9857);
or U10576 (N_10576,N_5543,N_8676);
nand U10577 (N_10577,N_9486,N_6710);
nand U10578 (N_10578,N_8983,N_7583);
or U10579 (N_10579,N_7217,N_7667);
and U10580 (N_10580,N_9174,N_6924);
or U10581 (N_10581,N_8465,N_8675);
and U10582 (N_10582,N_7134,N_9023);
or U10583 (N_10583,N_6239,N_6870);
and U10584 (N_10584,N_8603,N_9233);
nor U10585 (N_10585,N_9576,N_7120);
nand U10586 (N_10586,N_9060,N_6963);
nand U10587 (N_10587,N_9384,N_7942);
and U10588 (N_10588,N_9131,N_9618);
xor U10589 (N_10589,N_9479,N_5566);
nor U10590 (N_10590,N_9684,N_7857);
nand U10591 (N_10591,N_8442,N_8774);
nand U10592 (N_10592,N_8751,N_5654);
xor U10593 (N_10593,N_9563,N_9147);
or U10594 (N_10594,N_9533,N_9189);
nor U10595 (N_10595,N_5687,N_6786);
xnor U10596 (N_10596,N_7165,N_7519);
and U10597 (N_10597,N_8623,N_7505);
nand U10598 (N_10598,N_5499,N_7274);
nand U10599 (N_10599,N_8004,N_5609);
nand U10600 (N_10600,N_6949,N_8982);
nor U10601 (N_10601,N_7127,N_8902);
xor U10602 (N_10602,N_9461,N_7709);
or U10603 (N_10603,N_7955,N_9792);
xor U10604 (N_10604,N_9184,N_7467);
nand U10605 (N_10605,N_6265,N_7328);
nand U10606 (N_10606,N_7518,N_5672);
or U10607 (N_10607,N_8613,N_5769);
nand U10608 (N_10608,N_9777,N_7886);
nor U10609 (N_10609,N_7586,N_7633);
or U10610 (N_10610,N_5223,N_6497);
or U10611 (N_10611,N_7728,N_6747);
xor U10612 (N_10612,N_9421,N_5681);
or U10613 (N_10613,N_7239,N_6444);
and U10614 (N_10614,N_9504,N_6279);
xnor U10615 (N_10615,N_6409,N_9297);
nand U10616 (N_10616,N_6683,N_9170);
or U10617 (N_10617,N_6201,N_8540);
or U10618 (N_10618,N_8498,N_7738);
nor U10619 (N_10619,N_6641,N_7037);
and U10620 (N_10620,N_5563,N_6588);
and U10621 (N_10621,N_7750,N_9113);
or U10622 (N_10622,N_8922,N_7986);
nor U10623 (N_10623,N_6730,N_7412);
nor U10624 (N_10624,N_6722,N_9148);
or U10625 (N_10625,N_7264,N_8648);
xor U10626 (N_10626,N_9588,N_9303);
nor U10627 (N_10627,N_8885,N_5383);
xnor U10628 (N_10628,N_8144,N_7171);
xnor U10629 (N_10629,N_7576,N_7540);
or U10630 (N_10630,N_6886,N_7032);
nor U10631 (N_10631,N_5491,N_6777);
or U10632 (N_10632,N_9430,N_7199);
nand U10633 (N_10633,N_5498,N_6578);
or U10634 (N_10634,N_6062,N_5710);
and U10635 (N_10635,N_7768,N_8846);
or U10636 (N_10636,N_5115,N_6252);
nand U10637 (N_10637,N_7242,N_5731);
nand U10638 (N_10638,N_5107,N_5742);
nor U10639 (N_10639,N_8264,N_8183);
and U10640 (N_10640,N_5317,N_9089);
and U10641 (N_10641,N_7936,N_5229);
nor U10642 (N_10642,N_8020,N_9858);
or U10643 (N_10643,N_6986,N_8333);
nor U10644 (N_10644,N_8723,N_6569);
and U10645 (N_10645,N_8993,N_5277);
and U10646 (N_10646,N_6325,N_8254);
or U10647 (N_10647,N_5770,N_7141);
nand U10648 (N_10648,N_7972,N_5021);
xor U10649 (N_10649,N_9660,N_9944);
nor U10650 (N_10650,N_7893,N_7832);
xor U10651 (N_10651,N_7881,N_7954);
nand U10652 (N_10652,N_8361,N_9933);
nor U10653 (N_10653,N_8652,N_9417);
nor U10654 (N_10654,N_7457,N_8131);
xnor U10655 (N_10655,N_5436,N_8526);
and U10656 (N_10656,N_8323,N_9136);
nor U10657 (N_10657,N_6589,N_9288);
and U10658 (N_10658,N_8011,N_5750);
nor U10659 (N_10659,N_5783,N_7788);
xnor U10660 (N_10660,N_9525,N_7003);
and U10661 (N_10661,N_5611,N_7436);
nor U10662 (N_10662,N_5241,N_8762);
or U10663 (N_10663,N_7266,N_9954);
nor U10664 (N_10664,N_8110,N_8302);
xor U10665 (N_10665,N_5335,N_5262);
or U10666 (N_10666,N_8794,N_5740);
nor U10667 (N_10667,N_6994,N_5914);
or U10668 (N_10668,N_5069,N_9791);
or U10669 (N_10669,N_5958,N_5353);
nor U10670 (N_10670,N_5119,N_5549);
xnor U10671 (N_10671,N_9891,N_7114);
nor U10672 (N_10672,N_5040,N_9203);
nor U10673 (N_10673,N_5085,N_6892);
nor U10674 (N_10674,N_6159,N_9945);
xnor U10675 (N_10675,N_8312,N_9851);
nor U10676 (N_10676,N_7705,N_5244);
or U10677 (N_10677,N_8121,N_8587);
and U10678 (N_10678,N_9435,N_5011);
and U10679 (N_10679,N_6916,N_8656);
or U10680 (N_10680,N_5826,N_8799);
xnor U10681 (N_10681,N_8141,N_8945);
xor U10682 (N_10682,N_9049,N_5771);
nor U10683 (N_10683,N_7854,N_7263);
nand U10684 (N_10684,N_5159,N_6750);
or U10685 (N_10685,N_7743,N_9337);
nand U10686 (N_10686,N_7340,N_7050);
or U10687 (N_10687,N_9359,N_9654);
nand U10688 (N_10688,N_8201,N_7480);
nor U10689 (N_10689,N_8160,N_9261);
and U10690 (N_10690,N_8130,N_6264);
xor U10691 (N_10691,N_9382,N_9825);
or U10692 (N_10692,N_6568,N_6185);
nand U10693 (N_10693,N_8220,N_9407);
xnor U10694 (N_10694,N_5099,N_8305);
and U10695 (N_10695,N_9124,N_8733);
nand U10696 (N_10696,N_9540,N_5781);
nor U10697 (N_10697,N_5105,N_5511);
xor U10698 (N_10698,N_7432,N_5359);
or U10699 (N_10699,N_5516,N_5433);
nand U10700 (N_10700,N_7720,N_7192);
and U10701 (N_10701,N_7623,N_7732);
nor U10702 (N_10702,N_8481,N_9806);
and U10703 (N_10703,N_7639,N_8269);
xnor U10704 (N_10704,N_6608,N_9898);
nand U10705 (N_10705,N_5670,N_8257);
and U10706 (N_10706,N_6190,N_6967);
and U10707 (N_10707,N_8003,N_6538);
xnor U10708 (N_10708,N_9419,N_5825);
nand U10709 (N_10709,N_5022,N_7711);
nor U10710 (N_10710,N_5714,N_8683);
or U10711 (N_10711,N_9989,N_6526);
and U10712 (N_10712,N_6128,N_6305);
nor U10713 (N_10713,N_9205,N_8658);
nor U10714 (N_10714,N_9252,N_7603);
or U10715 (N_10715,N_8098,N_5564);
and U10716 (N_10716,N_7688,N_7602);
nor U10717 (N_10717,N_9062,N_5544);
and U10718 (N_10718,N_9094,N_6919);
nand U10719 (N_10719,N_5751,N_6800);
and U10720 (N_10720,N_7204,N_6953);
or U10721 (N_10721,N_5969,N_8601);
nand U10722 (N_10722,N_9581,N_8978);
xnor U10723 (N_10723,N_6714,N_7495);
or U10724 (N_10724,N_7937,N_7638);
nand U10725 (N_10725,N_9884,N_7220);
xnor U10726 (N_10726,N_7166,N_7016);
nor U10727 (N_10727,N_7808,N_5092);
nor U10728 (N_10728,N_5939,N_6603);
or U10729 (N_10729,N_7219,N_9953);
nor U10730 (N_10730,N_6727,N_5905);
or U10731 (N_10731,N_9820,N_9744);
nand U10732 (N_10732,N_9613,N_7761);
nor U10733 (N_10733,N_7119,N_5346);
and U10734 (N_10734,N_7866,N_8032);
or U10735 (N_10735,N_8233,N_6776);
nor U10736 (N_10736,N_5178,N_7513);
or U10737 (N_10737,N_6703,N_5363);
xnor U10738 (N_10738,N_6599,N_8898);
and U10739 (N_10739,N_5986,N_8210);
nor U10740 (N_10740,N_7137,N_6882);
or U10741 (N_10741,N_5063,N_9753);
and U10742 (N_10742,N_7488,N_5098);
or U10743 (N_10743,N_8914,N_7914);
nor U10744 (N_10744,N_8867,N_7812);
or U10745 (N_10745,N_9609,N_9471);
nor U10746 (N_10746,N_6275,N_8050);
nand U10747 (N_10747,N_6121,N_9350);
and U10748 (N_10748,N_7179,N_9841);
xnor U10749 (N_10749,N_8404,N_7413);
and U10750 (N_10750,N_7811,N_9721);
nand U10751 (N_10751,N_8738,N_6484);
nor U10752 (N_10752,N_6615,N_7977);
and U10753 (N_10753,N_6514,N_8491);
nor U10754 (N_10754,N_7792,N_7152);
nor U10755 (N_10755,N_6554,N_9118);
xor U10756 (N_10756,N_7883,N_5981);
xor U10757 (N_10757,N_8714,N_9008);
nor U10758 (N_10758,N_9765,N_5658);
nand U10759 (N_10759,N_5588,N_6768);
and U10760 (N_10760,N_5198,N_6511);
nand U10761 (N_10761,N_8618,N_7947);
xor U10762 (N_10762,N_6931,N_7710);
and U10763 (N_10763,N_8990,N_6631);
or U10764 (N_10764,N_6652,N_9782);
nand U10765 (N_10765,N_8597,N_6811);
xor U10766 (N_10766,N_6386,N_7492);
nand U10767 (N_10767,N_6327,N_9046);
and U10768 (N_10768,N_6881,N_6595);
and U10769 (N_10769,N_9126,N_5380);
and U10770 (N_10770,N_6007,N_9647);
and U10771 (N_10771,N_5409,N_8005);
and U10772 (N_10772,N_5431,N_6308);
nor U10773 (N_10773,N_6146,N_5578);
nor U10774 (N_10774,N_7384,N_7481);
or U10775 (N_10775,N_6995,N_5684);
nand U10776 (N_10776,N_7499,N_9516);
or U10777 (N_10777,N_9394,N_5097);
xor U10778 (N_10778,N_7791,N_9227);
or U10779 (N_10779,N_7558,N_9905);
or U10780 (N_10780,N_7077,N_8892);
nand U10781 (N_10781,N_7758,N_7950);
xor U10782 (N_10782,N_7760,N_5725);
xor U10783 (N_10783,N_8928,N_7752);
xor U10784 (N_10784,N_8979,N_5662);
nor U10785 (N_10785,N_5504,N_5415);
xnor U10786 (N_10786,N_7867,N_6672);
nand U10787 (N_10787,N_5133,N_9310);
or U10788 (N_10788,N_6433,N_6865);
nor U10789 (N_10789,N_7369,N_9722);
or U10790 (N_10790,N_5398,N_5430);
and U10791 (N_10791,N_8112,N_7054);
and U10792 (N_10792,N_8749,N_7015);
and U10793 (N_10793,N_7453,N_5009);
or U10794 (N_10794,N_9769,N_8968);
nand U10795 (N_10795,N_8303,N_7679);
nand U10796 (N_10796,N_5050,N_6521);
and U10797 (N_10797,N_8014,N_9138);
and U10798 (N_10798,N_6860,N_9116);
and U10799 (N_10799,N_5778,N_9092);
nand U10800 (N_10800,N_7699,N_8516);
and U10801 (N_10801,N_6940,N_7358);
or U10802 (N_10802,N_8706,N_7090);
nor U10803 (N_10803,N_5943,N_5542);
or U10804 (N_10804,N_5613,N_9667);
nor U10805 (N_10805,N_7949,N_7265);
or U10806 (N_10806,N_5597,N_9152);
nand U10807 (N_10807,N_6456,N_5440);
nand U10808 (N_10808,N_7101,N_5248);
and U10809 (N_10809,N_9267,N_5667);
nand U10810 (N_10810,N_9887,N_7177);
nor U10811 (N_10811,N_8102,N_6759);
nor U10812 (N_10812,N_9380,N_8041);
xor U10813 (N_10813,N_5082,N_6068);
or U10814 (N_10814,N_5173,N_8769);
xor U10815 (N_10815,N_6749,N_6913);
nand U10816 (N_10816,N_7209,N_7853);
nand U10817 (N_10817,N_5526,N_8703);
xor U10818 (N_10818,N_8777,N_6208);
and U10819 (N_10819,N_6165,N_7915);
or U10820 (N_10820,N_5754,N_9562);
nand U10821 (N_10821,N_8869,N_9415);
xnor U10822 (N_10822,N_8353,N_9547);
and U10823 (N_10823,N_5200,N_7663);
xor U10824 (N_10824,N_9798,N_8927);
xnor U10825 (N_10825,N_5623,N_5034);
nor U10826 (N_10826,N_9617,N_9949);
xnor U10827 (N_10827,N_7999,N_7592);
nand U10828 (N_10828,N_6022,N_7698);
and U10829 (N_10829,N_9220,N_9663);
nor U10830 (N_10830,N_8893,N_7491);
and U10831 (N_10831,N_9449,N_9513);
nor U10832 (N_10832,N_8568,N_9242);
nand U10833 (N_10833,N_7897,N_6110);
or U10834 (N_10834,N_8770,N_5576);
xnor U10835 (N_10835,N_5443,N_9249);
and U10836 (N_10836,N_6115,N_9678);
xnor U10837 (N_10837,N_8844,N_7379);
or U10838 (N_10838,N_9584,N_5554);
and U10839 (N_10839,N_9830,N_6102);
xnor U10840 (N_10840,N_7967,N_8308);
nand U10841 (N_10841,N_8054,N_8930);
or U10842 (N_10842,N_9641,N_8653);
nor U10843 (N_10843,N_6016,N_8148);
nand U10844 (N_10844,N_9349,N_6355);
nor U10845 (N_10845,N_9265,N_6921);
nor U10846 (N_10846,N_7932,N_5909);
or U10847 (N_10847,N_7203,N_8937);
or U10848 (N_10848,N_6378,N_6594);
or U10849 (N_10849,N_7289,N_9042);
and U10850 (N_10850,N_9543,N_8872);
xor U10851 (N_10851,N_9101,N_5185);
nor U10852 (N_10852,N_7342,N_8863);
nand U10853 (N_10853,N_8341,N_6907);
and U10854 (N_10854,N_7338,N_9943);
nand U10855 (N_10855,N_7736,N_6925);
nor U10856 (N_10856,N_7084,N_6632);
nor U10857 (N_10857,N_7532,N_6680);
and U10858 (N_10858,N_7668,N_8422);
nor U10859 (N_10859,N_7545,N_5839);
and U10860 (N_10860,N_6388,N_9579);
xnor U10861 (N_10861,N_8750,N_8283);
xnor U10862 (N_10862,N_5367,N_9104);
nand U10863 (N_10863,N_5246,N_5830);
and U10864 (N_10864,N_8451,N_7737);
xor U10865 (N_10865,N_7051,N_9916);
and U10866 (N_10866,N_6405,N_6126);
nand U10867 (N_10867,N_6828,N_9967);
or U10868 (N_10868,N_8813,N_9272);
or U10869 (N_10869,N_6306,N_7142);
or U10870 (N_10870,N_7320,N_9587);
and U10871 (N_10871,N_7624,N_5472);
xor U10872 (N_10872,N_8817,N_7438);
or U10873 (N_10873,N_7894,N_9784);
and U10874 (N_10874,N_9987,N_9711);
nand U10875 (N_10875,N_9959,N_8026);
xnor U10876 (N_10876,N_6627,N_6630);
and U10877 (N_10877,N_8584,N_9321);
and U10878 (N_10878,N_8772,N_7334);
nor U10879 (N_10879,N_6397,N_5425);
and U10880 (N_10880,N_6783,N_7909);
nand U10881 (N_10881,N_7157,N_5984);
nand U10882 (N_10882,N_7933,N_6130);
nand U10883 (N_10883,N_9072,N_5555);
or U10884 (N_10884,N_8518,N_6250);
or U10885 (N_10885,N_5955,N_8780);
or U10886 (N_10886,N_9367,N_9052);
nor U10887 (N_10887,N_6959,N_9065);
or U10888 (N_10888,N_7769,N_6992);
and U10889 (N_10889,N_7005,N_6439);
xor U10890 (N_10890,N_9750,N_7780);
xnor U10891 (N_10891,N_5247,N_8429);
xnor U10892 (N_10892,N_8845,N_6543);
and U10893 (N_10893,N_8117,N_5231);
nor U10894 (N_10894,N_5233,N_6837);
nand U10895 (N_10895,N_8033,N_6686);
xor U10896 (N_10896,N_6276,N_5032);
nor U10897 (N_10897,N_6231,N_6096);
nor U10898 (N_10898,N_9360,N_5458);
or U10899 (N_10899,N_9631,N_8950);
and U10900 (N_10900,N_9566,N_7373);
and U10901 (N_10901,N_8398,N_9197);
or U10902 (N_10902,N_8080,N_8946);
and U10903 (N_10903,N_7363,N_8118);
nor U10904 (N_10904,N_8440,N_9212);
nor U10905 (N_10905,N_8523,N_7325);
xor U10906 (N_10906,N_9606,N_8746);
or U10907 (N_10907,N_7061,N_9467);
xor U10908 (N_10908,N_6576,N_7870);
nor U10909 (N_10909,N_7423,N_7025);
and U10910 (N_10910,N_7494,N_8857);
and U10911 (N_10911,N_7962,N_9931);
xnor U10912 (N_10912,N_8489,N_9391);
xnor U10913 (N_10913,N_6309,N_8886);
nor U10914 (N_10914,N_6932,N_9438);
and U10915 (N_10915,N_5390,N_5885);
nor U10916 (N_10916,N_6320,N_5606);
nor U10917 (N_10917,N_7859,N_9834);
and U10918 (N_10918,N_8899,N_6662);
nor U10919 (N_10919,N_6505,N_8163);
or U10920 (N_10920,N_8731,N_6945);
nor U10921 (N_10921,N_9352,N_7365);
xor U10922 (N_10922,N_8170,N_7875);
xnor U10923 (N_10923,N_7714,N_5737);
nand U10924 (N_10924,N_5975,N_5414);
and U10925 (N_10925,N_8474,N_9375);
and U10926 (N_10926,N_6319,N_6065);
and U10927 (N_10927,N_8186,N_9117);
xor U10928 (N_10928,N_6873,N_9778);
nor U10929 (N_10929,N_8108,N_6725);
xor U10930 (N_10930,N_7155,N_8171);
nor U10931 (N_10931,N_6517,N_7735);
nor U10932 (N_10932,N_8007,N_7594);
and U10933 (N_10933,N_6552,N_8226);
xor U10934 (N_10934,N_7326,N_6920);
or U10935 (N_10935,N_9780,N_6461);
and U10936 (N_10936,N_6387,N_9151);
nand U10937 (N_10937,N_6753,N_9313);
and U10938 (N_10938,N_9794,N_7072);
nor U10939 (N_10939,N_8861,N_6076);
or U10940 (N_10940,N_7200,N_6821);
nor U10941 (N_10941,N_7354,N_5983);
nand U10942 (N_10942,N_5155,N_5158);
nand U10943 (N_10943,N_6825,N_5429);
xnor U10944 (N_10944,N_5988,N_7043);
nand U10945 (N_10945,N_6420,N_9268);
nor U10946 (N_10946,N_8182,N_7828);
nand U10947 (N_10947,N_6950,N_9011);
nand U10948 (N_10948,N_5466,N_9400);
nor U10949 (N_10949,N_5922,N_6181);
or U10950 (N_10950,N_6182,N_6775);
or U10951 (N_10951,N_8524,N_9214);
or U10952 (N_10952,N_7443,N_5795);
nand U10953 (N_10953,N_6935,N_8890);
xnor U10954 (N_10954,N_6422,N_8936);
nor U10955 (N_10955,N_8690,N_7123);
nand U10956 (N_10956,N_8548,N_9393);
nor U10957 (N_10957,N_8207,N_9831);
or U10958 (N_10958,N_8372,N_5850);
or U10959 (N_10959,N_6069,N_5266);
or U10960 (N_10960,N_6024,N_8816);
or U10961 (N_10961,N_5395,N_8741);
xnor U10962 (N_10962,N_9645,N_9464);
or U10963 (N_10963,N_6849,N_7981);
and U10964 (N_10964,N_8944,N_9503);
nand U10965 (N_10965,N_5362,N_7163);
and U10966 (N_10966,N_7683,N_7810);
nor U10967 (N_10967,N_5907,N_6018);
nand U10968 (N_10968,N_5831,N_7564);
and U10969 (N_10969,N_5297,N_5218);
or U10970 (N_10970,N_9416,N_5921);
nand U10971 (N_10971,N_6571,N_6732);
xor U10972 (N_10972,N_6083,N_9528);
xor U10973 (N_10973,N_9103,N_5477);
and U10974 (N_10974,N_9991,N_6124);
nor U10975 (N_10975,N_9761,N_9125);
and U10976 (N_10976,N_7299,N_9719);
and U10977 (N_10977,N_7057,N_9409);
nor U10978 (N_10978,N_9245,N_9100);
xor U10979 (N_10979,N_5964,N_7346);
xor U10980 (N_10980,N_7126,N_9980);
nor U10981 (N_10981,N_6862,N_6553);
and U10982 (N_10982,N_6390,N_5350);
nand U10983 (N_10983,N_8192,N_8379);
nand U10984 (N_10984,N_9290,N_8607);
nand U10985 (N_10985,N_6351,N_7549);
or U10986 (N_10986,N_9755,N_7173);
nand U10987 (N_10987,N_9567,N_9063);
xor U10988 (N_10988,N_7719,N_5987);
nor U10989 (N_10989,N_9561,N_7724);
and U10990 (N_10990,N_7821,N_9241);
xnor U10991 (N_10991,N_5461,N_7787);
or U10992 (N_10992,N_6122,N_5804);
or U10993 (N_10993,N_8128,N_5709);
and U10994 (N_10994,N_9144,N_9546);
nand U10995 (N_10995,N_8006,N_7500);
and U10996 (N_10996,N_6385,N_8953);
nor U10997 (N_10997,N_7201,N_6809);
xor U10998 (N_10998,N_9929,N_8076);
or U10999 (N_10999,N_5954,N_6219);
and U11000 (N_11000,N_6522,N_8580);
or U11001 (N_11001,N_5017,N_5065);
nand U11002 (N_11002,N_7253,N_8394);
nor U11003 (N_11003,N_6878,N_5361);
nand U11004 (N_11004,N_6852,N_7533);
xnor U11005 (N_11005,N_9779,N_6736);
xor U11006 (N_11006,N_8332,N_6980);
nand U11007 (N_11007,N_5137,N_7417);
xor U11008 (N_11008,N_6876,N_7390);
xor U11009 (N_11009,N_6017,N_5393);
nor U11010 (N_11010,N_7182,N_6039);
xor U11011 (N_11011,N_9552,N_9324);
and U11012 (N_11012,N_8224,N_8948);
nor U11013 (N_11013,N_7296,N_5727);
xnor U11014 (N_11014,N_6266,N_5816);
nor U11015 (N_11015,N_7213,N_9168);
nor U11016 (N_11016,N_9616,N_5306);
nand U11017 (N_11017,N_7845,N_5112);
and U11018 (N_11018,N_6626,N_8513);
nor U11019 (N_11019,N_7175,N_5073);
and U11020 (N_11020,N_5744,N_7133);
and U11021 (N_11021,N_8590,N_7448);
and U11022 (N_11022,N_8049,N_8832);
and U11023 (N_11023,N_7793,N_8221);
or U11024 (N_11024,N_9379,N_6848);
nand U11025 (N_11025,N_5482,N_9615);
nor U11026 (N_11026,N_5813,N_6207);
and U11027 (N_11027,N_5479,N_7873);
nor U11028 (N_11028,N_7118,N_7930);
xor U11029 (N_11029,N_7541,N_6429);
or U11030 (N_11030,N_5074,N_6956);
and U11031 (N_11031,N_6586,N_7794);
or U11032 (N_11032,N_5886,N_5853);
nand U11033 (N_11033,N_6754,N_7322);
nor U11034 (N_11034,N_7604,N_9200);
and U11035 (N_11035,N_6583,N_9424);
xnor U11036 (N_11036,N_7987,N_8386);
and U11037 (N_11037,N_8792,N_8496);
or U11038 (N_11038,N_8396,N_9336);
nand U11039 (N_11039,N_6241,N_6063);
nand U11040 (N_11040,N_7609,N_5527);
nor U11041 (N_11041,N_5484,N_5553);
and U11042 (N_11042,N_9688,N_5858);
or U11043 (N_11043,N_8250,N_8104);
nor U11044 (N_11044,N_6629,N_9254);
xor U11045 (N_11045,N_8356,N_9362);
xnor U11046 (N_11046,N_5296,N_8093);
and U11047 (N_11047,N_7825,N_7485);
nand U11048 (N_11048,N_8157,N_8473);
and U11049 (N_11049,N_8411,N_9526);
and U11050 (N_11050,N_8490,N_7627);
nor U11051 (N_11051,N_7359,N_6172);
and U11052 (N_11052,N_9756,N_8599);
nand U11053 (N_11053,N_8449,N_6317);
and U11054 (N_11054,N_6236,N_7339);
nor U11055 (N_11055,N_7899,N_8668);
nor U11056 (N_11056,N_6688,N_8664);
xor U11057 (N_11057,N_6036,N_5936);
nand U11058 (N_11058,N_8145,N_5833);
and U11059 (N_11059,N_8605,N_6646);
nand U11060 (N_11060,N_8205,N_6579);
or U11061 (N_11061,N_5806,N_8619);
nor U11062 (N_11062,N_5132,N_9664);
nor U11063 (N_11063,N_8840,N_7944);
nand U11064 (N_11064,N_5066,N_9977);
nand U11065 (N_11065,N_7816,N_5490);
nand U11066 (N_11066,N_5349,N_8812);
xor U11067 (N_11067,N_5329,N_6246);
nand U11068 (N_11068,N_6209,N_9332);
and U11069 (N_11069,N_6597,N_7444);
or U11070 (N_11070,N_5509,N_8446);
or U11071 (N_11071,N_7934,N_8115);
or U11072 (N_11072,N_8827,N_8290);
and U11073 (N_11073,N_9444,N_6335);
nor U11074 (N_11074,N_8704,N_7064);
nor U11075 (N_11075,N_7840,N_6824);
or U11076 (N_11076,N_7327,N_6834);
nor U11077 (N_11077,N_6513,N_6509);
xor U11078 (N_11078,N_9996,N_5903);
xor U11079 (N_11079,N_9455,N_6261);
and U11080 (N_11080,N_7980,N_9239);
nor U11081 (N_11081,N_7983,N_9710);
xor U11082 (N_11082,N_8419,N_5212);
or U11083 (N_11083,N_9246,N_6023);
or U11084 (N_11084,N_9269,N_6541);
and U11085 (N_11085,N_8900,N_8162);
xor U11086 (N_11086,N_6715,N_6491);
and U11087 (N_11087,N_8046,N_6817);
xor U11088 (N_11088,N_8864,N_9193);
and U11089 (N_11089,N_8808,N_7078);
or U11090 (N_11090,N_9328,N_9160);
nor U11091 (N_11091,N_7011,N_8239);
nand U11092 (N_11092,N_7629,N_8299);
and U11093 (N_11093,N_8364,N_8317);
or U11094 (N_11094,N_6237,N_8138);
nor U11095 (N_11095,N_7680,N_8293);
and U11096 (N_11096,N_5254,N_5288);
or U11097 (N_11097,N_6620,N_5232);
nor U11098 (N_11098,N_8838,N_5608);
nand U11099 (N_11099,N_5221,N_8595);
xor U11100 (N_11100,N_8755,N_8539);
xor U11101 (N_11101,N_9534,N_5522);
xor U11102 (N_11102,N_5216,N_7830);
nor U11103 (N_11103,N_9188,N_8581);
and U11104 (N_11104,N_6819,N_7848);
nand U11105 (N_11105,N_6647,N_8427);
nor U11106 (N_11106,N_6969,N_9904);
nor U11107 (N_11107,N_7801,N_9619);
and U11108 (N_11108,N_5381,N_8891);
nor U11109 (N_11109,N_8211,N_8380);
or U11110 (N_11110,N_6430,N_7212);
or U11111 (N_11111,N_7527,N_5309);
nand U11112 (N_11112,N_5236,N_5293);
and U11113 (N_11113,N_5171,N_8022);
and U11114 (N_11114,N_5873,N_5059);
xnor U11115 (N_11115,N_7230,N_9007);
or U11116 (N_11116,N_7028,N_9502);
or U11117 (N_11117,N_5957,N_8241);
or U11118 (N_11118,N_9511,N_5318);
or U11119 (N_11119,N_8273,N_5811);
and U11120 (N_11120,N_5483,N_5411);
and U11121 (N_11121,N_6606,N_9797);
xnor U11122 (N_11122,N_7387,N_5108);
nor U11123 (N_11123,N_7570,N_6353);
xor U11124 (N_11124,N_6374,N_6890);
nor U11125 (N_11125,N_6403,N_7026);
nand U11126 (N_11126,N_8370,N_5708);
and U11127 (N_11127,N_8593,N_6216);
nand U11128 (N_11128,N_5292,N_7493);
nand U11129 (N_11129,N_5805,N_6621);
xnor U11130 (N_11130,N_7193,N_6440);
nand U11131 (N_11131,N_8839,N_6915);
xnor U11132 (N_11132,N_9741,N_6233);
xnor U11133 (N_11133,N_6401,N_5632);
nand U11134 (N_11134,N_5228,N_7048);
nand U11135 (N_11135,N_9881,N_8815);
and U11136 (N_11136,N_7347,N_9720);
and U11137 (N_11137,N_7139,N_5836);
and U11138 (N_11138,N_6955,N_8511);
and U11139 (N_11139,N_6729,N_7901);
and U11140 (N_11140,N_6655,N_7757);
nor U11141 (N_11141,N_9050,N_7335);
xor U11142 (N_11142,N_6889,N_8384);
nor U11143 (N_11143,N_6451,N_5539);
nand U11144 (N_11144,N_6350,N_5739);
or U11145 (N_11145,N_5616,N_9410);
xor U11146 (N_11146,N_5572,N_9551);
nand U11147 (N_11147,N_5268,N_8729);
or U11148 (N_11148,N_8962,N_8865);
xnor U11149 (N_11149,N_9127,N_5941);
nor U11150 (N_11150,N_5579,N_9853);
xor U11151 (N_11151,N_7475,N_6160);
nand U11152 (N_11152,N_6479,N_8153);
and U11153 (N_11153,N_8596,N_6984);
xnor U11154 (N_11154,N_9133,N_9638);
nor U11155 (N_11155,N_6258,N_9492);
xnor U11156 (N_11156,N_5982,N_7953);
and U11157 (N_11157,N_9759,N_6839);
nor U11158 (N_11158,N_8971,N_7115);
xor U11159 (N_11159,N_7941,N_9045);
xor U11160 (N_11160,N_5680,N_7017);
or U11161 (N_11161,N_6389,N_8350);
and U11162 (N_11162,N_7590,N_9338);
and U11163 (N_11163,N_8833,N_9439);
and U11164 (N_11164,N_5399,N_6095);
nand U11165 (N_11165,N_5448,N_6853);
or U11166 (N_11166,N_8659,N_8133);
and U11167 (N_11167,N_6471,N_6537);
xnor U11168 (N_11168,N_8889,N_5761);
nor U11169 (N_11169,N_9890,N_9143);
and U11170 (N_11170,N_8434,N_5441);
and U11171 (N_11171,N_5577,N_7969);
or U11172 (N_11172,N_7301,N_6694);
or U11173 (N_11173,N_6954,N_6078);
nor U11174 (N_11174,N_5487,N_7031);
or U11175 (N_11175,N_8156,N_9677);
or U11176 (N_11176,N_5235,N_6705);
xor U11177 (N_11177,N_6199,N_7311);
and U11178 (N_11178,N_9740,N_8529);
or U11179 (N_11179,N_9309,N_5533);
xnor U11180 (N_11180,N_9508,N_8608);
or U11181 (N_11181,N_8197,N_5256);
or U11182 (N_11182,N_7925,N_9804);
and U11183 (N_11183,N_7029,N_9734);
or U11184 (N_11184,N_9255,N_8776);
or U11185 (N_11185,N_8288,N_9966);
and U11186 (N_11186,N_7049,N_8091);
nand U11187 (N_11187,N_6642,N_8300);
nor U11188 (N_11188,N_8680,N_5303);
and U11189 (N_11189,N_7878,N_9520);
nor U11190 (N_11190,N_7450,N_8443);
nand U11191 (N_11191,N_9069,N_9266);
nand U11192 (N_11192,N_6944,N_7408);
or U11193 (N_11193,N_6140,N_7116);
nand U11194 (N_11194,N_6371,N_6263);
xor U11195 (N_11195,N_9208,N_7861);
and U11196 (N_11196,N_7961,N_5835);
nor U11197 (N_11197,N_8285,N_5186);
or U11198 (N_11198,N_8067,N_6109);
or U11199 (N_11199,N_8139,N_7610);
nor U11200 (N_11200,N_8802,N_7809);
and U11201 (N_11201,N_5180,N_7099);
and U11202 (N_11202,N_6438,N_8724);
nand U11203 (N_11203,N_9474,N_9555);
nand U11204 (N_11204,N_8616,N_6981);
nor U11205 (N_11205,N_9202,N_7837);
nor U11206 (N_11206,N_6902,N_9666);
xnor U11207 (N_11207,N_9308,N_5538);
nand U11208 (N_11208,N_5518,N_5388);
or U11209 (N_11209,N_6291,N_9992);
nand U11210 (N_11210,N_9053,N_7874);
and U11211 (N_11211,N_5238,N_7159);
or U11212 (N_11212,N_8761,N_8214);
nor U11213 (N_11213,N_6851,N_6805);
and U11214 (N_11214,N_8494,N_7802);
nor U11215 (N_11215,N_5862,N_5898);
xor U11216 (N_11216,N_7517,N_9354);
xnor U11217 (N_11217,N_8941,N_8759);
xor U11218 (N_11218,N_6778,N_7676);
and U11219 (N_11219,N_7689,N_7132);
nor U11220 (N_11220,N_9872,N_6214);
nand U11221 (N_11221,N_7010,N_6773);
and U11222 (N_11222,N_5713,N_5096);
or U11223 (N_11223,N_6478,N_9907);
or U11224 (N_11224,N_7587,N_8184);
nand U11225 (N_11225,N_9304,N_8114);
nor U11226 (N_11226,N_6737,N_7665);
nand U11227 (N_11227,N_7148,N_5581);
xnor U11228 (N_11228,N_9692,N_9019);
nor U11229 (N_11229,N_6093,N_8748);
or U11230 (N_11230,N_8830,N_8822);
nor U11231 (N_11231,N_5308,N_7708);
or U11232 (N_11232,N_6075,N_8455);
and U11233 (N_11233,N_7247,N_8122);
nor U11234 (N_11234,N_6006,N_5829);
or U11235 (N_11235,N_5264,N_9590);
or U11236 (N_11236,N_6835,N_5626);
nand U11237 (N_11237,N_6613,N_5591);
nor U11238 (N_11238,N_7503,N_9859);
nor U11239 (N_11239,N_9192,N_7946);
nand U11240 (N_11240,N_6298,N_9494);
nor U11241 (N_11241,N_8310,N_5338);
or U11242 (N_11242,N_7872,N_8413);
and U11243 (N_11243,N_7121,N_9077);
nor U11244 (N_11244,N_8216,N_5610);
or U11245 (N_11245,N_8236,N_7851);
xor U11246 (N_11246,N_9675,N_5327);
nand U11247 (N_11247,N_5602,N_8620);
nand U11248 (N_11248,N_7385,N_9748);
nand U11249 (N_11249,N_9162,N_6030);
and U11250 (N_11250,N_9865,N_8739);
nor U11251 (N_11251,N_7243,N_7150);
or U11252 (N_11252,N_9585,N_7058);
nor U11253 (N_11253,N_6755,N_5568);
or U11254 (N_11254,N_5893,N_9015);
or U11255 (N_11255,N_9139,N_8229);
xnor U11256 (N_11256,N_8203,N_7416);
and U11257 (N_11257,N_8635,N_8604);
xnor U11258 (N_11258,N_8172,N_9737);
xnor U11259 (N_11259,N_8428,N_8256);
nor U11260 (N_11260,N_7440,N_9299);
xnor U11261 (N_11261,N_6136,N_9300);
nor U11262 (N_11262,N_8092,N_5220);
and U11263 (N_11263,N_5760,N_9706);
or U11264 (N_11264,N_6520,N_9224);
and U11265 (N_11265,N_7314,N_5250);
and U11266 (N_11266,N_8782,N_7140);
nand U11267 (N_11267,N_5603,N_8661);
nand U11268 (N_11268,N_8566,N_6118);
nor U11269 (N_11269,N_8147,N_8368);
nand U11270 (N_11270,N_7035,N_7994);
nand U11271 (N_11271,N_5113,N_7581);
nand U11272 (N_11272,N_6143,N_7596);
nand U11273 (N_11273,N_9079,N_7033);
and U11274 (N_11274,N_7731,N_8426);
and U11275 (N_11275,N_9465,N_6187);
or U11276 (N_11276,N_7351,N_9648);
and U11277 (N_11277,N_6564,N_5326);
and U11278 (N_11278,N_9691,N_7333);
nand U11279 (N_11279,N_7730,N_7965);
nand U11280 (N_11280,N_9743,N_5535);
or U11281 (N_11281,N_5765,N_9392);
nor U11282 (N_11282,N_7938,N_5439);
and U11283 (N_11283,N_9796,N_5612);
or U11284 (N_11284,N_7672,N_7588);
and U11285 (N_11285,N_7895,N_9625);
nand U11286 (N_11286,N_9041,N_5023);
and U11287 (N_11287,N_6380,N_9186);
and U11288 (N_11288,N_6217,N_8044);
or U11289 (N_11289,N_8000,N_9882);
or U11290 (N_11290,N_8575,N_7439);
nand U11291 (N_11291,N_7920,N_5259);
or U11292 (N_11292,N_5843,N_8870);
nand U11293 (N_11293,N_8339,N_9902);
nand U11294 (N_11294,N_5894,N_6829);
or U11295 (N_11295,N_5051,N_5502);
or U11296 (N_11296,N_7721,N_8307);
nand U11297 (N_11297,N_6524,N_9961);
nand U11298 (N_11298,N_7534,N_5594);
and U11299 (N_11299,N_9892,N_5953);
nand U11300 (N_11300,N_9109,N_7103);
or U11301 (N_11301,N_6911,N_6887);
nand U11302 (N_11302,N_8246,N_8309);
nor U11303 (N_11303,N_7315,N_6163);
nor U11304 (N_11304,N_9568,N_8263);
xor U11305 (N_11305,N_7526,N_5874);
xor U11306 (N_11306,N_6546,N_9178);
and U11307 (N_11307,N_9176,N_5583);
and U11308 (N_11308,N_8579,N_8132);
and U11309 (N_11309,N_7529,N_8025);
nand U11310 (N_11310,N_9941,N_6752);
xor U11311 (N_11311,N_9403,N_5619);
and U11312 (N_11312,N_7082,N_7924);
nor U11313 (N_11313,N_7789,N_8448);
xnor U11314 (N_11314,N_6296,N_5702);
and U11315 (N_11315,N_8142,N_5962);
nand U11316 (N_11316,N_5203,N_5712);
or U11317 (N_11317,N_6123,N_8227);
and U11318 (N_11318,N_8094,N_8966);
nand U11319 (N_11319,N_6609,N_8956);
or U11320 (N_11320,N_5407,N_6154);
nand U11321 (N_11321,N_8829,N_7476);
nand U11322 (N_11322,N_6417,N_6290);
nand U11323 (N_11323,N_9920,N_6844);
and U11324 (N_11324,N_8810,N_9498);
or U11325 (N_11325,N_8847,N_5384);
and U11326 (N_11326,N_7822,N_5420);
nor U11327 (N_11327,N_8276,N_9861);
or U11328 (N_11328,N_5867,N_5168);
or U11329 (N_11329,N_6841,N_6790);
nor U11330 (N_11330,N_7827,N_7814);
nand U11331 (N_11331,N_7506,N_6339);
or U11332 (N_11332,N_7659,N_8101);
nor U11333 (N_11333,N_8393,N_8238);
and U11334 (N_11334,N_8820,N_5560);
or U11335 (N_11335,N_8536,N_6117);
nor U11336 (N_11336,N_9210,N_5728);
xor U11337 (N_11337,N_7310,N_7985);
nand U11338 (N_11338,N_6454,N_5261);
nor U11339 (N_11339,N_6977,N_6671);
or U11340 (N_11340,N_5510,N_8710);
nor U11341 (N_11341,N_7404,N_5141);
or U11342 (N_11342,N_8883,N_9669);
nand U11343 (N_11343,N_8452,N_5493);
or U11344 (N_11344,N_7411,N_8991);
nor U11345 (N_11345,N_7272,N_9999);
nor U11346 (N_11346,N_5971,N_7226);
xor U11347 (N_11347,N_6958,N_5064);
and U11348 (N_11348,N_7329,N_5824);
or U11349 (N_11349,N_6067,N_6735);
and U11350 (N_11350,N_6349,N_9196);
nand U11351 (N_11351,N_5582,N_5772);
nor U11352 (N_11352,N_9622,N_7382);
and U11353 (N_11353,N_8409,N_6054);
or U11354 (N_11354,N_9912,N_6808);
and U11355 (N_11355,N_6088,N_5331);
nand U11356 (N_11356,N_6605,N_9020);
nor U11357 (N_11357,N_9082,N_6989);
xor U11358 (N_11358,N_6820,N_9689);
nand U11359 (N_11359,N_7543,N_8055);
xor U11360 (N_11360,N_9997,N_8304);
and U11361 (N_11361,N_6884,N_5515);
xnor U11362 (N_11362,N_5123,N_7912);
nor U11363 (N_11363,N_8728,N_7473);
xnor U11364 (N_11364,N_9057,N_9344);
nor U11365 (N_11365,N_7951,N_5265);
or U11366 (N_11366,N_5135,N_8786);
and U11367 (N_11367,N_5642,N_8209);
nand U11368 (N_11368,N_5294,N_5960);
xnor U11369 (N_11369,N_8722,N_7060);
nor U11370 (N_11370,N_7024,N_9788);
xnor U11371 (N_11371,N_5865,N_5796);
or U11372 (N_11372,N_5519,N_8070);
and U11373 (N_11373,N_8487,N_9098);
and U11374 (N_11374,N_8178,N_6229);
nand U11375 (N_11375,N_5330,N_6611);
xnor U11376 (N_11376,N_6719,N_6412);
nor U11377 (N_11377,N_7516,N_9556);
and U11378 (N_11378,N_7300,N_5090);
and U11379 (N_11379,N_8435,N_6489);
nor U11380 (N_11380,N_6162,N_5120);
nand U11381 (N_11381,N_8583,N_8935);
or U11382 (N_11382,N_5567,N_6287);
and U11383 (N_11383,N_6934,N_8545);
nor U11384 (N_11384,N_5419,N_6381);
xnor U11385 (N_11385,N_5652,N_5676);
xnor U11386 (N_11386,N_5891,N_6011);
nor U11387 (N_11387,N_7197,N_7508);
or U11388 (N_11388,N_6540,N_8522);
and U11389 (N_11389,N_5114,N_8672);
and U11390 (N_11390,N_8556,N_7104);
nor U11391 (N_11391,N_5076,N_6046);
xor U11392 (N_11392,N_6899,N_5030);
or U11393 (N_11393,N_9179,N_7466);
or U11394 (N_11394,N_5167,N_7729);
nor U11395 (N_11395,N_7474,N_9446);
nor U11396 (N_11396,N_7318,N_7862);
xor U11397 (N_11397,N_9209,N_5501);
and U11398 (N_11398,N_7215,N_5821);
and U11399 (N_11399,N_6709,N_8912);
nand U11400 (N_11400,N_7378,N_8146);
xor U11401 (N_11401,N_6293,N_8346);
nor U11402 (N_11402,N_9672,N_7019);
and U11403 (N_11403,N_7553,N_9105);
nor U11404 (N_11404,N_9725,N_8778);
nor U11405 (N_11405,N_9632,N_8063);
and U11406 (N_11406,N_8187,N_6885);
or U11407 (N_11407,N_9096,N_8514);
nand U11408 (N_11408,N_5589,N_8232);
and U11409 (N_11409,N_8992,N_5048);
nor U11410 (N_11410,N_5694,N_9298);
and U11411 (N_11411,N_5260,N_7105);
nor U11412 (N_11412,N_9263,N_7337);
or U11413 (N_11413,N_6058,N_5718);
nor U11414 (N_11414,N_9340,N_6565);
xnor U11415 (N_11415,N_8697,N_9472);
and U11416 (N_11416,N_5925,N_8528);
and U11417 (N_11417,N_9727,N_8319);
and U11418 (N_11418,N_5629,N_5129);
nor U11419 (N_11419,N_8850,N_6869);
and U11420 (N_11420,N_7305,N_9078);
nor U11421 (N_11421,N_8058,N_7939);
or U11422 (N_11422,N_9624,N_5031);
xor U11423 (N_11423,N_9173,N_6793);
and U11424 (N_11424,N_7218,N_5997);
nand U11425 (N_11425,N_9457,N_6679);
or U11426 (N_11426,N_6482,N_8517);
and U11427 (N_11427,N_9448,N_8354);
xor U11428 (N_11428,N_7282,N_6475);
nand U11429 (N_11429,N_6826,N_6833);
and U11430 (N_11430,N_5370,N_8225);
xor U11431 (N_11431,N_8016,N_8318);
nand U11432 (N_11432,N_5109,N_9877);
xor U11433 (N_11433,N_7525,N_7285);
nor U11434 (N_11434,N_6544,N_5598);
nor U11435 (N_11435,N_8642,N_6744);
and U11436 (N_11436,N_6292,N_5033);
xor U11437 (N_11437,N_8929,N_7907);
xnor U11438 (N_11438,N_9827,N_5550);
and U11439 (N_11439,N_6262,N_9458);
or U11440 (N_11440,N_5016,N_9993);
xor U11441 (N_11441,N_5790,N_6856);
nand U11442 (N_11442,N_6555,N_6503);
nor U11443 (N_11443,N_8436,N_9402);
nor U11444 (N_11444,N_6506,N_7268);
or U11445 (N_11445,N_5630,N_8532);
nor U11446 (N_11446,N_8030,N_7613);
nand U11447 (N_11447,N_5840,N_9270);
and U11448 (N_11448,N_9809,N_5170);
nor U11449 (N_11449,N_5786,N_6964);
xnor U11450 (N_11450,N_7906,N_8967);
or U11451 (N_11451,N_7044,N_6450);
nand U11452 (N_11452,N_9702,N_7039);
or U11453 (N_11453,N_6539,N_5757);
and U11454 (N_11454,N_7164,N_6660);
xnor U11455 (N_11455,N_5087,N_5213);
or U11456 (N_11456,N_7766,N_5647);
xnor U11457 (N_11457,N_6174,N_8471);
xor U11458 (N_11458,N_9982,N_6044);
or U11459 (N_11459,N_7561,N_8543);
or U11460 (N_11460,N_9636,N_8193);
xnor U11461 (N_11461,N_6516,N_9234);
xnor U11462 (N_11462,N_8052,N_6019);
and U11463 (N_11463,N_7733,N_7128);
xnor U11464 (N_11464,N_6321,N_5126);
and U11465 (N_11465,N_5949,N_7125);
xor U11466 (N_11466,N_7259,N_7826);
and U11467 (N_11467,N_5512,N_9497);
nor U11468 (N_11468,N_6206,N_6584);
nor U11469 (N_11469,N_6762,N_7012);
or U11470 (N_11470,N_7643,N_8717);
and U11471 (N_11471,N_9454,N_5849);
nand U11472 (N_11472,N_5067,N_6619);
xnor U11473 (N_11473,N_9459,N_5912);
and U11474 (N_11474,N_6467,N_6271);
xor U11475 (N_11475,N_8969,N_5328);
or U11476 (N_11476,N_6232,N_9278);
nand U11477 (N_11477,N_9644,N_5139);
xor U11478 (N_11478,N_7971,N_6712);
nand U11479 (N_11479,N_6294,N_8687);
nand U11480 (N_11480,N_7231,N_8107);
xor U11481 (N_11481,N_6668,N_5354);
nor U11482 (N_11482,N_6724,N_7395);
or U11483 (N_11483,N_9163,N_8873);
or U11484 (N_11484,N_8764,N_6406);
and U11485 (N_11485,N_9095,N_7697);
xnor U11486 (N_11486,N_8925,N_5450);
nand U11487 (N_11487,N_9869,N_9473);
and U11488 (N_11488,N_7727,N_6370);
and U11489 (N_11489,N_9972,N_7511);
nand U11490 (N_11490,N_7205,N_6623);
or U11491 (N_11491,N_8218,N_8056);
nor U11492 (N_11492,N_9634,N_6904);
nor U11493 (N_11493,N_6367,N_8432);
or U11494 (N_11494,N_6323,N_7580);
and U11495 (N_11495,N_7774,N_7095);
or U11496 (N_11496,N_5705,N_8077);
nand U11497 (N_11497,N_5933,N_9469);
nor U11498 (N_11498,N_9789,N_6188);
or U11499 (N_11499,N_8271,N_6156);
nand U11500 (N_11500,N_7428,N_7224);
xnor U11501 (N_11501,N_6211,N_5978);
nand U11502 (N_11502,N_8954,N_7754);
xor U11503 (N_11503,N_7111,N_5540);
or U11504 (N_11504,N_9033,N_5149);
and U11505 (N_11505,N_7089,N_7551);
and U11506 (N_11506,N_7238,N_5557);
xnor U11507 (N_11507,N_7926,N_7174);
xnor U11508 (N_11508,N_5945,N_5800);
or U11509 (N_11509,N_8298,N_7270);
xnor U11510 (N_11510,N_7047,N_9911);
xor U11511 (N_11511,N_6090,N_7344);
xnor U11512 (N_11512,N_8355,N_6212);
xnor U11513 (N_11513,N_5325,N_8650);
and U11514 (N_11514,N_7777,N_7927);
xor U11515 (N_11515,N_5315,N_7464);
nand U11516 (N_11516,N_5847,N_9671);
and U11517 (N_11517,N_7074,N_5494);
or U11518 (N_11518,N_6074,N_9058);
or U11519 (N_11519,N_7957,N_9976);
or U11520 (N_11520,N_6810,N_6636);
or U11521 (N_11521,N_5360,N_9387);
nand U11522 (N_11522,N_9565,N_8174);
and U11523 (N_11523,N_9925,N_5224);
xnor U11524 (N_11524,N_8450,N_7569);
xnor U11525 (N_11525,N_6512,N_5131);
and U11526 (N_11526,N_7707,N_5994);
nand U11527 (N_11527,N_7068,N_6373);
nand U11528 (N_11528,N_5199,N_9866);
xnor U11529 (N_11529,N_9450,N_6375);
or U11530 (N_11530,N_9747,N_5950);
and U11531 (N_11531,N_9404,N_5628);
xor U11532 (N_11532,N_9818,N_9423);
or U11533 (N_11533,N_8743,N_9171);
and U11534 (N_11534,N_7198,N_5868);
xor U11535 (N_11535,N_8497,N_6487);
nor U11536 (N_11536,N_9986,N_8975);
and U11537 (N_11537,N_7803,N_6687);
nor U11538 (N_11538,N_6384,N_9452);
nor U11539 (N_11539,N_8500,N_6473);
and U11540 (N_11540,N_6988,N_8352);
nor U11541 (N_11541,N_8699,N_8679);
and U11542 (N_11542,N_6343,N_7244);
or U11543 (N_11543,N_5736,N_5495);
nand U11544 (N_11544,N_7018,N_5617);
xor U11545 (N_11545,N_8505,N_8981);
nor U11546 (N_11546,N_7136,N_7400);
xnor U11547 (N_11547,N_9668,N_8995);
nor U11548 (N_11548,N_7149,N_8970);
nand U11549 (N_11549,N_7575,N_6815);
and U11550 (N_11550,N_5614,N_9895);
xor U11551 (N_11551,N_8828,N_5863);
and U11552 (N_11552,N_9032,N_9132);
nor U11553 (N_11553,N_7918,N_6900);
nand U11554 (N_11554,N_8200,N_7210);
nand U11555 (N_11555,N_6772,N_8651);
and U11556 (N_11556,N_6633,N_8923);
xor U11557 (N_11557,N_9495,N_6111);
and U11558 (N_11558,N_8018,N_8176);
nand U11559 (N_11559,N_9348,N_5142);
nor U11560 (N_11560,N_6477,N_9816);
and U11561 (N_11561,N_6765,N_6286);
nor U11562 (N_11562,N_9317,N_9389);
nand U11563 (N_11563,N_5860,N_9602);
xor U11564 (N_11564,N_7739,N_6285);
xnor U11565 (N_11565,N_5722,N_6155);
or U11566 (N_11566,N_7618,N_9289);
or U11567 (N_11567,N_7619,N_7183);
and U11568 (N_11568,N_6807,N_5762);
nor U11569 (N_11569,N_7286,N_5311);
nor U11570 (N_11570,N_5342,N_6166);
or U11571 (N_11571,N_9878,N_8259);
xor U11572 (N_11572,N_6788,N_9653);
nor U11573 (N_11573,N_8525,N_6442);
and U11574 (N_11574,N_8924,N_5344);
nor U11575 (N_11575,N_9482,N_7779);
and U11576 (N_11576,N_6230,N_7716);
nor U11577 (N_11577,N_6689,N_6864);
xnor U11578 (N_11578,N_5323,N_8634);
and U11579 (N_11579,N_6625,N_7913);
nor U11580 (N_11580,N_6580,N_6443);
or U11581 (N_11581,N_9554,N_8378);
nor U11582 (N_11582,N_6936,N_5562);
nor U11583 (N_11583,N_6169,N_6354);
xor U11584 (N_11584,N_5471,N_8785);
or U11585 (N_11585,N_8395,N_5721);
or U11586 (N_11586,N_9175,N_6695);
nand U11587 (N_11587,N_8804,N_6396);
nand U11588 (N_11588,N_7225,N_8646);
xor U11589 (N_11589,N_6802,N_6280);
nand U11590 (N_11590,N_7835,N_6299);
nor U11591 (N_11591,N_6574,N_8140);
nor U11592 (N_11592,N_5991,N_9301);
nand U11593 (N_11593,N_5828,N_9889);
xnor U11594 (N_11594,N_6114,N_8291);
and U11595 (N_11595,N_5475,N_7023);
nand U11596 (N_11596,N_9855,N_6991);
or U11597 (N_11597,N_9548,N_6108);
xnor U11598 (N_11598,N_6928,N_8281);
nand U11599 (N_11599,N_7654,N_7437);
or U11600 (N_11600,N_9913,N_9256);
xnor U11601 (N_11601,N_5596,N_9371);
xnor U11602 (N_11602,N_7292,N_9698);
xnor U11603 (N_11603,N_5275,N_6032);
or U11604 (N_11604,N_6535,N_5685);
nor U11605 (N_11605,N_8031,N_9291);
xnor U11606 (N_11606,N_6066,N_7591);
or U11607 (N_11607,N_6675,N_8527);
nor U11608 (N_11608,N_6000,N_5271);
and U11609 (N_11609,N_7796,N_8934);
nand U11610 (N_11610,N_6682,N_6717);
and U11611 (N_11611,N_7539,N_7908);
xnor U11612 (N_11612,N_5480,N_6987);
nor U11613 (N_11613,N_9844,N_7657);
nand U11614 (N_11614,N_9199,N_9155);
nand U11615 (N_11615,N_6563,N_9919);
nand U11616 (N_11616,N_7191,N_6651);
or U11617 (N_11617,N_6779,N_6721);
or U11618 (N_11618,N_6283,N_9260);
nand U11619 (N_11619,N_5046,N_7445);
nor U11620 (N_11620,N_8654,N_9201);
nand U11621 (N_11621,N_7945,N_9767);
and U11622 (N_11622,N_5427,N_9770);
and U11623 (N_11623,N_8515,N_5435);
or U11624 (N_11624,N_5270,N_9642);
and U11625 (N_11625,N_8381,N_6342);
or U11626 (N_11626,N_5154,N_6448);
nor U11627 (N_11627,N_6918,N_9043);
and U11628 (N_11628,N_7135,N_9014);
nor U11629 (N_11629,N_6060,N_9323);
and U11630 (N_11630,N_8245,N_6037);
xnor U11631 (N_11631,N_5352,N_5794);
xor U11632 (N_11632,N_9276,N_5438);
nor U11633 (N_11633,N_5930,N_9752);
and U11634 (N_11634,N_5808,N_9901);
nand U11635 (N_11635,N_8868,N_9573);
nor U11636 (N_11636,N_7469,N_6840);
nor U11637 (N_11637,N_9248,N_8598);
and U11638 (N_11638,N_7122,N_7717);
nand U11639 (N_11639,N_6638,N_9003);
nor U11640 (N_11640,N_8589,N_5845);
xnor U11641 (N_11641,N_9621,N_7579);
or U11642 (N_11642,N_5901,N_6774);
or U11643 (N_11643,N_8779,N_8113);
nand U11644 (N_11644,N_9523,N_7350);
and U11645 (N_11645,N_9703,N_6094);
or U11646 (N_11646,N_8949,N_8190);
or U11647 (N_11647,N_5184,N_7009);
and U11648 (N_11648,N_8678,N_8677);
xor U11649 (N_11649,N_7658,N_8835);
or U11650 (N_11650,N_9536,N_8726);
xnor U11651 (N_11651,N_9048,N_9181);
nor U11652 (N_11652,N_8760,N_8391);
or U11653 (N_11653,N_5312,N_8017);
or U11654 (N_11654,N_8188,N_5812);
and U11655 (N_11655,N_6277,N_8533);
or U11656 (N_11656,N_9028,N_7463);
and U11657 (N_11657,N_7785,N_6617);
nor U11658 (N_11658,N_8574,N_6352);
or U11659 (N_11659,N_9640,N_7391);
nand U11660 (N_11660,N_5205,N_8235);
nand U11661 (N_11661,N_7370,N_7747);
nand U11662 (N_11662,N_5688,N_8753);
or U11663 (N_11663,N_9545,N_6173);
nand U11664 (N_11664,N_6801,N_9158);
nor U11665 (N_11665,N_5319,N_6415);
xnor U11666 (N_11666,N_7403,N_8242);
xor U11667 (N_11667,N_6943,N_8400);
and U11668 (N_11668,N_9366,N_6585);
nand U11669 (N_11669,N_8175,N_9086);
nor U11670 (N_11670,N_5651,N_7056);
or U11671 (N_11671,N_5214,N_7839);
and U11672 (N_11672,N_9141,N_9088);
or U11673 (N_11673,N_9596,N_5735);
or U11674 (N_11674,N_6314,N_9532);
nor U11675 (N_11675,N_6012,N_5932);
nand U11676 (N_11676,N_8796,N_6120);
nand U11677 (N_11677,N_9707,N_9054);
xnor U11678 (N_11678,N_8405,N_6847);
nand U11679 (N_11679,N_9693,N_7889);
or U11680 (N_11680,N_6933,N_8800);
nand U11681 (N_11681,N_8952,N_7462);
and U11682 (N_11682,N_5675,N_7013);
nand U11683 (N_11683,N_6875,N_8986);
xor U11684 (N_11684,N_9447,N_8519);
and U11685 (N_11685,N_5187,N_8939);
nor U11686 (N_11686,N_8649,N_9538);
xnor U11687 (N_11687,N_8570,N_6200);
or U11688 (N_11688,N_7542,N_7154);
and U11689 (N_11689,N_5356,N_8388);
or U11690 (N_11690,N_7607,N_8788);
or U11691 (N_11691,N_7214,N_5230);
nand U11692 (N_11692,N_6942,N_9918);
or U11693 (N_11693,N_9635,N_8530);
nor U11694 (N_11694,N_7922,N_5083);
xor U11695 (N_11695,N_8086,N_7935);
or U11696 (N_11696,N_8555,N_5759);
and U11697 (N_11697,N_5992,N_5697);
or U11698 (N_11698,N_7235,N_5861);
and U11699 (N_11699,N_8546,N_5462);
or U11700 (N_11700,N_8123,N_8897);
and U11701 (N_11701,N_9514,N_9236);
or U11702 (N_11702,N_7974,N_5106);
and U11703 (N_11703,N_8260,N_5474);
xor U11704 (N_11704,N_5507,N_9091);
and U11705 (N_11705,N_7371,N_9279);
xor U11706 (N_11706,N_5707,N_5998);
nor U11707 (N_11707,N_5719,N_6020);
nor U11708 (N_11708,N_8168,N_6684);
xnor U11709 (N_11709,N_5447,N_7996);
and U11710 (N_11710,N_5683,N_6031);
nand U11711 (N_11711,N_5197,N_6333);
xor U11712 (N_11712,N_7004,N_9910);
or U11713 (N_11713,N_5428,N_9754);
nand U11714 (N_11714,N_6769,N_7973);
nand U11715 (N_11715,N_8720,N_6894);
nand U11716 (N_11716,N_7910,N_9840);
nand U11717 (N_11717,N_5055,N_5575);
xnor U11718 (N_11718,N_7002,N_7206);
and U11719 (N_11719,N_5061,N_7748);
and U11720 (N_11720,N_5570,N_9772);
xnor U11721 (N_11721,N_8557,N_6005);
nor U11722 (N_11722,N_6087,N_6092);
and U11723 (N_11723,N_9363,N_5780);
or U11724 (N_11724,N_7483,N_5421);
nand U11725 (N_11725,N_5376,N_9325);
and U11726 (N_11726,N_7399,N_6693);
and U11727 (N_11727,N_8071,N_7421);
xnor U11728 (N_11728,N_9694,N_7294);
nand U11729 (N_11729,N_9594,N_5130);
nor U11730 (N_11730,N_9453,N_7929);
xnor U11731 (N_11731,N_6587,N_7694);
or U11732 (N_11732,N_6272,N_9026);
nand U11733 (N_11733,N_8932,N_6781);
or U11734 (N_11734,N_9736,N_6424);
nor U11735 (N_11735,N_5369,N_7715);
and U11736 (N_11736,N_8947,N_5717);
xnor U11737 (N_11737,N_6027,N_6416);
nor U11738 (N_11738,N_8135,N_5273);
nand U11739 (N_11739,N_8594,N_5571);
and U11740 (N_11740,N_9735,N_5300);
nand U11741 (N_11741,N_6125,N_7267);
nor U11742 (N_11742,N_8702,N_9334);
or U11743 (N_11743,N_9656,N_8369);
nor U11744 (N_11744,N_5144,N_7221);
or U11745 (N_11745,N_6307,N_8165);
or U11746 (N_11746,N_6855,N_5336);
nor U11747 (N_11747,N_8043,N_5406);
nand U11748 (N_11748,N_6508,N_8564);
and U11749 (N_11749,N_9683,N_8083);
or U11750 (N_11750,N_8329,N_7762);
and U11751 (N_11751,N_5377,N_6957);
nor U11752 (N_11752,N_5189,N_9923);
xnor U11753 (N_11753,N_5690,N_5242);
or U11754 (N_11754,N_5639,N_7615);
xnor U11755 (N_11755,N_9639,N_5182);
nand U11756 (N_11756,N_7678,N_5075);
xor U11757 (N_11757,N_9369,N_7130);
or U11758 (N_11758,N_9610,N_9039);
nor U11759 (N_11759,N_5449,N_9405);
nand U11760 (N_11760,N_9821,N_8358);
xnor U11761 (N_11761,N_7145,N_7383);
nand U11762 (N_11762,N_6782,N_8826);
or U11763 (N_11763,N_7246,N_8994);
or U11764 (N_11764,N_9906,N_7631);
and U11765 (N_11765,N_9947,N_9955);
nor U11766 (N_11766,N_9680,N_9829);
and U11767 (N_11767,N_7374,N_7504);
nand U11768 (N_11768,N_7921,N_5020);
and U11769 (N_11769,N_5403,N_9819);
or U11770 (N_11770,N_8842,N_7336);
and U11771 (N_11771,N_7252,N_5100);
and U11772 (N_11772,N_8315,N_8973);
xnor U11773 (N_11773,N_9401,N_8572);
or U11774 (N_11774,N_8537,N_7348);
nor U11775 (N_11775,N_7988,N_5446);
xnor U11776 (N_11776,N_9374,N_6726);
nor U11777 (N_11777,N_8920,N_9080);
xor U11778 (N_11778,N_9601,N_9627);
nand U11779 (N_11779,N_9728,N_5432);
or U11780 (N_11780,N_7073,N_7250);
xnor U11781 (N_11781,N_5333,N_9607);
and U11782 (N_11782,N_9274,N_5111);
nand U11783 (N_11783,N_9965,N_7449);
or U11784 (N_11784,N_5251,N_6515);
xor U11785 (N_11785,N_9828,N_7067);
xor U11786 (N_11786,N_5656,N_9685);
nand U11787 (N_11787,N_9068,N_6192);
nor U11788 (N_11788,N_9215,N_7815);
nor U11789 (N_11789,N_9130,N_5444);
and U11790 (N_11790,N_9451,N_5025);
and U11791 (N_11791,N_7573,N_5890);
nor U11792 (N_11792,N_8166,N_7276);
or U11793 (N_11793,N_6741,N_9564);
and U11794 (N_11794,N_5078,N_7281);
and U11795 (N_11795,N_8698,N_8809);
nand U11796 (N_11796,N_8752,N_5166);
xnor U11797 (N_11797,N_5854,N_5068);
xor U11798 (N_11798,N_8085,N_6542);
or U11799 (N_11799,N_5569,N_9790);
and U11800 (N_11800,N_7419,N_8081);
nor U11801 (N_11801,N_8882,N_9240);
and U11802 (N_11802,N_6663,N_8045);
or U11803 (N_11803,N_9655,N_5884);
nor U11804 (N_11804,N_6803,N_9031);
and U11805 (N_11805,N_9908,N_6049);
or U11806 (N_11806,N_9883,N_8685);
xnor U11807 (N_11807,N_9445,N_8021);
nand U11808 (N_11808,N_6792,N_8228);
or U11809 (N_11809,N_7229,N_8313);
and U11810 (N_11810,N_7858,N_6926);
and U11811 (N_11811,N_6365,N_9111);
and U11812 (N_11812,N_6697,N_8360);
or U11813 (N_11813,N_5928,N_7313);
xor U11814 (N_11814,N_8268,N_6338);
or U11815 (N_11815,N_6757,N_8222);
or U11816 (N_11816,N_8349,N_7756);
or U11817 (N_11817,N_9216,N_5973);
xor U11818 (N_11818,N_8376,N_7546);
nand U11819 (N_11819,N_6033,N_7303);
and U11820 (N_11820,N_9036,N_5169);
nor U11821 (N_11821,N_7065,N_5852);
nor U11822 (N_11822,N_9327,N_6295);
nor U11823 (N_11823,N_5703,N_8403);
nand U11824 (N_11824,N_8989,N_6593);
xnor U11825 (N_11825,N_5343,N_8240);
nor U11826 (N_11826,N_9793,N_5856);
nor U11827 (N_11827,N_5904,N_5118);
or U11828 (N_11828,N_9760,N_9115);
nor U11829 (N_11829,N_7585,N_8592);
nor U11830 (N_11830,N_5004,N_5057);
and U11831 (N_11831,N_5634,N_5799);
and U11832 (N_11832,N_8806,N_6983);
xnor U11833 (N_11833,N_8196,N_9968);
xnor U11834 (N_11834,N_8060,N_5895);
nor U11835 (N_11835,N_6359,N_8600);
nand U11836 (N_11836,N_9431,N_9283);
and U11837 (N_11837,N_5175,N_6100);
and U11838 (N_11838,N_8807,N_8324);
and U11839 (N_11839,N_8682,N_9598);
nor U11840 (N_11840,N_6673,N_5970);
xor U11841 (N_11841,N_8078,N_8734);
nor U11842 (N_11842,N_5316,N_9429);
xor U11843 (N_11843,N_8615,N_5267);
nor U11844 (N_11844,N_9180,N_7982);
xor U11845 (N_11845,N_8701,N_7605);
nand U11846 (N_11846,N_5102,N_9386);
or U11847 (N_11847,N_6770,N_7169);
or U11848 (N_11848,N_5919,N_6794);
or U11849 (N_11849,N_6667,N_8047);
or U11850 (N_11850,N_8495,N_9612);
nor U11851 (N_11851,N_6042,N_8585);
nand U11852 (N_11852,N_5842,N_9102);
and U11853 (N_11853,N_5961,N_5789);
xor U11854 (N_11854,N_7284,N_7496);
xor U11855 (N_11855,N_5537,N_9320);
or U11856 (N_11856,N_8874,N_5434);
nor U11857 (N_11857,N_5019,N_9134);
and U11858 (N_11858,N_6402,N_8282);
and U11859 (N_11859,N_7632,N_5645);
nor U11860 (N_11860,N_8997,N_9909);
and U11861 (N_11861,N_7071,N_9983);
nor U11862 (N_11862,N_5291,N_6009);
nand U11863 (N_11863,N_6215,N_7477);
xnor U11864 (N_11864,N_6930,N_7471);
nor U11865 (N_11865,N_5174,N_8856);
xnor U11866 (N_11866,N_9758,N_8424);
or U11867 (N_11867,N_9120,N_9505);
and U11868 (N_11868,N_8357,N_6191);
nand U11869 (N_11869,N_7565,N_5459);
xnor U11870 (N_11870,N_7622,N_5855);
nand U11871 (N_11871,N_5437,N_7394);
or U11872 (N_11872,N_6284,N_9510);
nor U11873 (N_11873,N_8410,N_7548);
nand U11874 (N_11874,N_6099,N_7097);
or U11875 (N_11875,N_7324,N_8416);
nor U11876 (N_11876,N_8918,N_7406);
xnor U11877 (N_11877,N_9811,N_5776);
nor U11878 (N_11878,N_9302,N_5161);
and U11879 (N_11879,N_8639,N_5276);
or U11880 (N_11880,N_8909,N_8034);
or U11881 (N_11881,N_9221,N_9845);
or U11882 (N_11882,N_5993,N_8492);
or U11883 (N_11883,N_7251,N_5996);
xnor U11884 (N_11884,N_8002,N_5086);
nor U11885 (N_11885,N_8784,N_6221);
xnor U11886 (N_11886,N_6618,N_5980);
or U11887 (N_11887,N_5788,N_7976);
nor U11888 (N_11888,N_6573,N_9428);
xor U11889 (N_11889,N_7979,N_5053);
nand U11890 (N_11890,N_8008,N_7409);
xnor U11891 (N_11891,N_5880,N_6047);
nand U11892 (N_11892,N_9119,N_7628);
or U11893 (N_11893,N_9863,N_9738);
and U11894 (N_11894,N_7782,N_6398);
xor U11895 (N_11895,N_7283,N_9335);
nor U11896 (N_11896,N_7571,N_8884);
nand U11897 (N_11897,N_6785,N_6282);
and U11898 (N_11898,N_6791,N_9442);
and U11899 (N_11899,N_8399,N_6528);
nand U11900 (N_11900,N_5400,N_5552);
nor U11901 (N_11901,N_8535,N_7279);
xor U11902 (N_11902,N_7645,N_5148);
nor U11903 (N_11903,N_9679,N_8591);
or U11904 (N_11904,N_7109,N_9373);
nor U11905 (N_11905,N_8219,N_7877);
or U11906 (N_11906,N_8637,N_7256);
xnor U11907 (N_11907,N_7007,N_5989);
nor U11908 (N_11908,N_7059,N_6962);
or U11909 (N_11909,N_8666,N_9030);
nor U11910 (N_11910,N_9481,N_6223);
nor U11911 (N_11911,N_7648,N_8965);
nor U11912 (N_11912,N_9460,N_6034);
nand U11913 (N_11913,N_7902,N_5093);
nand U11914 (N_11914,N_8270,N_5815);
nand U11915 (N_11915,N_5505,N_7484);
and U11916 (N_11916,N_5924,N_8499);
xnor U11917 (N_11917,N_9603,N_9426);
nor U11918 (N_11918,N_8385,N_8943);
and U11919 (N_11919,N_6650,N_9817);
nand U11920 (N_11920,N_5927,N_6347);
or U11921 (N_11921,N_8202,N_6081);
or U11922 (N_11922,N_8960,N_8181);
xor U11923 (N_11923,N_5556,N_5896);
nor U11924 (N_11924,N_7293,N_6097);
xor U11925 (N_11925,N_8280,N_7188);
xnor U11926 (N_11926,N_8998,N_6029);
nor U11927 (N_11927,N_8417,N_9886);
nand U11928 (N_11928,N_8119,N_8387);
and U11929 (N_11929,N_8286,N_7554);
xor U11930 (N_11930,N_7312,N_8129);
xor U11931 (N_11931,N_6927,N_8797);
and U11932 (N_11932,N_9733,N_6329);
or U11933 (N_11933,N_6993,N_5351);
nor U11934 (N_11934,N_8237,N_6676);
xnor U11935 (N_11935,N_5749,N_5528);
nand U11936 (N_11936,N_9001,N_5633);
nand U11937 (N_11937,N_6249,N_9558);
nor U11938 (N_11938,N_6164,N_5956);
or U11939 (N_11939,N_6656,N_7479);
or U11940 (N_11940,N_5959,N_8686);
nor U11941 (N_11941,N_7287,N_7345);
nand U11942 (N_11942,N_6533,N_9582);
xor U11943 (N_11943,N_6670,N_6485);
or U11944 (N_11944,N_9764,N_8027);
nand U11945 (N_11945,N_6898,N_6874);
xnor U11946 (N_11946,N_8673,N_8647);
xnor U11947 (N_11947,N_8716,N_6908);
xor U11948 (N_11948,N_6866,N_6481);
nand U11949 (N_11949,N_5627,N_9553);
xnor U11950 (N_11950,N_9537,N_5902);
nand U11951 (N_11951,N_5488,N_7458);
nand U11952 (N_11952,N_9978,N_9643);
and U11953 (N_11953,N_5179,N_9930);
xnor U11954 (N_11954,N_5565,N_6938);
or U11955 (N_11955,N_7261,N_5985);
xor U11956 (N_11956,N_8253,N_7692);
and U11957 (N_11957,N_6996,N_7249);
or U11958 (N_11958,N_5723,N_8823);
nor U11959 (N_11959,N_5070,N_7952);
nor U11960 (N_11960,N_9365,N_5313);
or U11961 (N_11961,N_7616,N_8915);
and U11962 (N_11962,N_5881,N_6814);
nor U11963 (N_11963,N_6364,N_8688);
nor U11964 (N_11964,N_5364,N_5358);
nand U11965 (N_11965,N_5976,N_6414);
and U11966 (N_11966,N_8433,N_8048);
and U11967 (N_11967,N_6013,N_6551);
nor U11968 (N_11968,N_7677,N_8996);
nand U11969 (N_11969,N_9012,N_6098);
and U11970 (N_11970,N_7784,N_5698);
and U11971 (N_11971,N_5152,N_8294);
xor U11972 (N_11972,N_6836,N_5777);
nand U11973 (N_11973,N_9475,N_9307);
xor U11974 (N_11974,N_6103,N_8278);
and U11975 (N_11975,N_5062,N_5341);
nor U11976 (N_11976,N_6766,N_8406);
xor U11977 (N_11977,N_7376,N_7831);
nand U11978 (N_11978,N_7306,N_7662);
nor U11979 (N_11979,N_7236,N_7931);
nor U11980 (N_11980,N_7846,N_7330);
xnor U11981 (N_11981,N_8940,N_7790);
and U11982 (N_11982,N_9314,N_5476);
nand U11983 (N_11983,N_6048,N_9107);
xnor U11984 (N_11984,N_8331,N_8447);
or U11985 (N_11985,N_7353,N_5792);
and U11986 (N_11986,N_7660,N_5413);
xnor U11987 (N_11987,N_8407,N_8408);
nand U11988 (N_11988,N_9823,N_9600);
or U11989 (N_11989,N_6228,N_7398);
nor U11990 (N_11990,N_6135,N_6812);
and U11991 (N_11991,N_8252,N_8617);
nand U11992 (N_11992,N_7781,N_5314);
and U11993 (N_11993,N_8301,N_6780);
nor U11994 (N_11994,N_6345,N_5453);
or U11995 (N_11995,N_5456,N_6476);
or U11996 (N_11996,N_6255,N_5503);
or U11997 (N_11997,N_7040,N_8412);
nand U11998 (N_11998,N_9056,N_5859);
and U11999 (N_11999,N_5913,N_6823);
nor U12000 (N_12000,N_9942,N_6592);
and U12001 (N_12001,N_8931,N_6357);
or U12002 (N_12002,N_8831,N_6052);
xor U12003 (N_12003,N_8328,N_9950);
and U12004 (N_12004,N_5878,N_7849);
xor U12005 (N_12005,N_9273,N_9870);
xnor U12006 (N_12006,N_7036,N_8670);
xor U12007 (N_12007,N_8275,N_8336);
or U12008 (N_12008,N_8860,N_5532);
xor U12009 (N_12009,N_8103,N_7288);
and U12010 (N_12010,N_5470,N_6196);
nand U12011 (N_12011,N_7110,N_5834);
xor U12012 (N_12012,N_9145,N_5621);
or U12013 (N_12013,N_5457,N_9776);
nand U12014 (N_12014,N_6001,N_5585);
or U12015 (N_12015,N_7502,N_6713);
or U12016 (N_12016,N_5931,N_5424);
or U12017 (N_12017,N_8475,N_9586);
and U12018 (N_12018,N_8213,N_5249);
xnor U12019 (N_12019,N_7997,N_6635);
xnor U12020 (N_12020,N_5253,N_7478);
nand U12021 (N_12021,N_7863,N_8097);
and U12022 (N_12022,N_5002,N_9286);
xor U12023 (N_12023,N_7486,N_8821);
or U12024 (N_12024,N_7297,N_7536);
nand U12025 (N_12025,N_6059,N_5587);
nor U12026 (N_12026,N_6831,N_9888);
nand U12027 (N_12027,N_6071,N_8347);
nor U12028 (N_12028,N_7361,N_6297);
and U12029 (N_12029,N_9649,N_9611);
or U12030 (N_12030,N_6134,N_7684);
and U12031 (N_12031,N_9802,N_5465);
nor U12032 (N_12032,N_8414,N_9529);
nor U12033 (N_12033,N_8569,N_6379);
or U12034 (N_12034,N_5365,N_8111);
or U12035 (N_12035,N_8559,N_5775);
nor U12036 (N_12036,N_8488,N_9800);
and U12037 (N_12037,N_5210,N_6685);
xor U12038 (N_12038,N_8854,N_5846);
or U12039 (N_12039,N_6341,N_7841);
xor U12040 (N_12040,N_8636,N_7465);
and U12041 (N_12041,N_6665,N_7030);
and U12042 (N_12042,N_8503,N_8367);
or U12043 (N_12043,N_8345,N_7117);
or U12044 (N_12044,N_7807,N_8895);
and U12045 (N_12045,N_6334,N_6458);
xnor U12046 (N_12046,N_7700,N_6362);
xnor U12047 (N_12047,N_5295,N_9137);
nor U12048 (N_12048,N_6268,N_5405);
or U12049 (N_12049,N_8476,N_8881);
nor U12050 (N_12050,N_7405,N_7695);
nand U12051 (N_12051,N_9990,N_6596);
and U12052 (N_12052,N_6604,N_8334);
xor U12053 (N_12053,N_6445,N_9218);
nor U12054 (N_12054,N_6452,N_7530);
or U12055 (N_12055,N_5755,N_6131);
nor U12056 (N_12056,N_9592,N_5536);
nor U12057 (N_12057,N_8582,N_9361);
xnor U12058 (N_12058,N_7372,N_5524);
nor U12059 (N_12059,N_6161,N_7868);
nand U12060 (N_12060,N_8483,N_6669);
and U12061 (N_12061,N_9657,N_6966);
and U12062 (N_12062,N_5037,N_6021);
nand U12063 (N_12063,N_8573,N_7674);
and U12064 (N_12064,N_5088,N_8790);
nand U12065 (N_12065,N_7578,N_6244);
or U12066 (N_12066,N_6822,N_5386);
or U12067 (N_12067,N_5604,N_5636);
xor U12068 (N_12068,N_5010,N_7308);
nor U12069 (N_12069,N_5766,N_7751);
nor U12070 (N_12070,N_9934,N_9318);
or U12071 (N_12071,N_7424,N_7093);
nor U12072 (N_12072,N_5999,N_5418);
nor U12073 (N_12073,N_8781,N_9257);
nor U12074 (N_12074,N_7041,N_8079);
or U12075 (N_12075,N_5686,N_9822);
nor U12076 (N_12076,N_5926,N_8578);
and U12077 (N_12077,N_8980,N_7522);
nand U12078 (N_12078,N_7027,N_8095);
nand U12079 (N_12079,N_7741,N_9550);
xor U12080 (N_12080,N_7461,N_5546);
xnor U12081 (N_12081,N_6198,N_7202);
xnor U12082 (N_12082,N_5104,N_7786);
nor U12083 (N_12083,N_6723,N_9837);
xor U12084 (N_12084,N_9194,N_6132);
xor U12085 (N_12085,N_5743,N_7108);
xor U12086 (N_12086,N_6480,N_9522);
nand U12087 (N_12087,N_8711,N_9899);
and U12088 (N_12088,N_5797,N_6897);
nor U12089 (N_12089,N_9786,N_8463);
xnor U12090 (N_12090,N_9676,N_9593);
nor U12091 (N_12091,N_7042,N_8611);
nor U12092 (N_12092,N_6168,N_5445);
nand U12093 (N_12093,N_7381,N_5027);
and U12094 (N_12094,N_5286,N_9874);
nor U12095 (N_12095,N_5307,N_5787);
xnor U12096 (N_12096,N_8064,N_9436);
nor U12097 (N_12097,N_7038,N_6531);
nor U12098 (N_12098,N_6720,N_5738);
xor U12099 (N_12099,N_6896,N_5937);
nor U12100 (N_12100,N_5631,N_7690);
xor U12101 (N_12101,N_8955,N_5807);
or U12102 (N_12102,N_7723,N_9462);
nand U12103 (N_12103,N_7661,N_7510);
or U12104 (N_12104,N_5701,N_7393);
xor U12105 (N_12105,N_8705,N_9896);
xor U12106 (N_12106,N_7331,N_7595);
nor U12107 (N_12107,N_7817,N_7567);
or U12108 (N_12108,N_9024,N_5551);
or U12109 (N_12109,N_5408,N_6382);
and U12110 (N_12110,N_9785,N_9815);
and U12111 (N_12111,N_5746,N_6040);
xor U12112 (N_12112,N_5426,N_5695);
xor U12113 (N_12113,N_6203,N_7022);
xor U12114 (N_12114,N_6901,N_8445);
or U12115 (N_12115,N_7092,N_6227);
or U12116 (N_12116,N_7718,N_7241);
or U12117 (N_12117,N_6437,N_8987);
and U12118 (N_12118,N_8348,N_9673);
xor U12119 (N_12119,N_5643,N_5140);
nor U12120 (N_12120,N_8217,N_9087);
nand U12121 (N_12121,N_8155,N_9938);
xnor U12122 (N_12122,N_8374,N_5906);
nand U12123 (N_12123,N_7823,N_6644);
nand U12124 (N_12124,N_9936,N_7052);
and U12125 (N_12125,N_6871,N_5281);
and U12126 (N_12126,N_7552,N_5838);
or U12127 (N_12127,N_8866,N_5496);
nand U12128 (N_12128,N_8284,N_7094);
nor U12129 (N_12129,N_5517,N_5274);
or U12130 (N_12130,N_7773,N_8693);
xnor U12131 (N_12131,N_9076,N_8707);
nand U12132 (N_12132,N_7514,N_7917);
nand U12133 (N_12133,N_6806,N_6666);
xor U12134 (N_12134,N_5084,N_5252);
and U12135 (N_12135,N_9630,N_7341);
and U12136 (N_12136,N_9742,N_5691);
nand U12137 (N_12137,N_9456,N_7970);
xnor U12138 (N_12138,N_9177,N_5018);
nor U12139 (N_12139,N_7647,N_9235);
nand U12140 (N_12140,N_8783,N_7185);
nand U12141 (N_12141,N_6240,N_8628);
and U12142 (N_12142,N_5530,N_6607);
xnor U12143 (N_12143,N_5145,N_9259);
xnor U12144 (N_12144,N_8159,N_5382);
nand U12145 (N_12145,N_6288,N_8708);
nor U12146 (N_12146,N_5734,N_8090);
and U12147 (N_12147,N_6332,N_5451);
and U12148 (N_12148,N_6830,N_9686);
or U12149 (N_12149,N_9121,N_5165);
nor U12150 (N_12150,N_5202,N_5008);
and U12151 (N_12151,N_6008,N_9483);
or U12152 (N_12152,N_9411,N_5534);
or U12153 (N_12153,N_8343,N_7208);
nor U12154 (N_12154,N_8740,N_8773);
or U12155 (N_12155,N_5375,N_8430);
and U12156 (N_12156,N_5875,N_9490);
nor U12157 (N_12157,N_9928,N_6718);
and U12158 (N_12158,N_5848,N_8880);
xor U12159 (N_12159,N_7885,N_5301);
xor U12160 (N_12160,N_7098,N_5641);
nor U12161 (N_12161,N_8258,N_8206);
and U12162 (N_12162,N_7681,N_7636);
xnor U12163 (N_12163,N_9085,N_5237);
and U12164 (N_12164,N_6178,N_7860);
xor U12165 (N_12165,N_8244,N_7687);
nor U12166 (N_12166,N_8588,N_9726);
nand U12167 (N_12167,N_8629,N_5394);
nand U12168 (N_12168,N_5810,N_7855);
nand U12169 (N_12169,N_7968,N_7685);
and U12170 (N_12170,N_8735,N_9518);
xor U12171 (N_12171,N_7124,N_7021);
or U12172 (N_12172,N_8951,N_8732);
and U12173 (N_12173,N_8179,N_5726);
and U12174 (N_12174,N_8657,N_6247);
nand U12175 (N_12175,N_9894,N_5561);
xor U12176 (N_12176,N_9093,N_8910);
nor U12177 (N_12177,N_6281,N_5573);
and U12178 (N_12178,N_6557,N_9433);
or U12179 (N_12179,N_7451,N_9161);
nor U12180 (N_12180,N_5802,N_8961);
or U12181 (N_12181,N_9029,N_6691);
xnor U12182 (N_12182,N_6326,N_8363);
nand U12183 (N_12183,N_8757,N_6974);
nor U12184 (N_12184,N_6193,N_9466);
xnor U12185 (N_12185,N_8694,N_7069);
or U12186 (N_12186,N_5525,N_7572);
xor U12187 (N_12187,N_8389,N_9687);
nand U12188 (N_12188,N_9838,N_6502);
nand U12189 (N_12189,N_5923,N_8314);
nand U12190 (N_12190,N_5967,N_9381);
and U12191 (N_12191,N_9900,N_6973);
or U12192 (N_12192,N_8627,N_8458);
nor U12193 (N_12193,N_5678,N_5819);
or U12194 (N_12194,N_7147,N_5899);
xnor U12195 (N_12195,N_7498,N_6507);
and U12196 (N_12196,N_8059,N_9795);
nand U12197 (N_12197,N_6149,N_5026);
nand U12198 (N_12198,N_8553,N_7414);
and U12199 (N_12199,N_8631,N_5529);
nor U12200 (N_12200,N_9662,N_8963);
nor U12201 (N_12201,N_9066,N_9295);
and U12202 (N_12202,N_7083,N_7713);
nand U12203 (N_12203,N_9583,N_5995);
and U12204 (N_12204,N_7234,N_6270);
xor U12205 (N_12205,N_6175,N_9975);
xnor U12206 (N_12206,N_5827,N_9370);
nor U12207 (N_12207,N_8421,N_7000);
nor U12208 (N_12208,N_7349,N_6138);
xnor U12209 (N_12209,N_6500,N_8274);
nand U12210 (N_12210,N_6180,N_8957);
nand U12211 (N_12211,N_5227,N_7455);
xnor U12212 (N_12212,N_6089,N_9476);
nor U12213 (N_12213,N_7507,N_6547);
and U12214 (N_12214,N_6278,N_5467);
nand U12215 (N_12215,N_6472,N_5234);
or U12216 (N_12216,N_6330,N_5208);
nand U12217 (N_12217,N_9347,N_6260);
nor U12218 (N_12218,N_9860,N_5116);
xnor U12219 (N_12219,N_5091,N_5442);
xor U12220 (N_12220,N_7186,N_7131);
nand U12221 (N_12221,N_9709,N_6743);
and U12222 (N_12222,N_7392,N_8316);
or U12223 (N_12223,N_6225,N_5682);
and U12224 (N_12224,N_5747,N_6369);
or U12225 (N_12225,N_7472,N_7427);
or U12226 (N_12226,N_5908,N_5080);
nand U12227 (N_12227,N_9083,N_6082);
nor U12228 (N_12228,N_8262,N_8736);
nand U12229 (N_12229,N_6854,N_7651);
nand U12230 (N_12230,N_7597,N_7887);
and U12231 (N_12231,N_7490,N_5191);
or U12232 (N_12232,N_5911,N_9106);
xnor U12233 (N_12233,N_7898,N_8606);
nor U12234 (N_12234,N_7637,N_5605);
xnor U12235 (N_12235,N_7984,N_5043);
nand U12236 (N_12236,N_5183,N_5454);
xnor U12237 (N_12237,N_9507,N_5347);
or U12238 (N_12238,N_9846,N_9097);
and U12239 (N_12239,N_9524,N_9681);
xnor U12240 (N_12240,N_9388,N_7799);
xor U12241 (N_12241,N_6581,N_9763);
nor U12242 (N_12242,N_9059,N_7189);
xnor U12243 (N_12243,N_6474,N_9803);
nor U12244 (N_12244,N_7100,N_6116);
nand U12245 (N_12245,N_6746,N_6426);
xnor U12246 (N_12246,N_6645,N_8287);
nand U12247 (N_12247,N_8512,N_6795);
nor U12248 (N_12248,N_6195,N_8415);
and U12249 (N_12249,N_9704,N_8191);
or U12250 (N_12250,N_5423,N_5049);
or U12251 (N_12251,N_8149,N_7928);
and U12252 (N_12252,N_9493,N_6465);
nor U12253 (N_12253,N_9854,N_9690);
xor U12254 (N_12254,N_9013,N_9651);
nand U12255 (N_12255,N_6084,N_6243);
and U12256 (N_12256,N_6459,N_9812);
and U12257 (N_12257,N_9326,N_9768);
or U12258 (N_12258,N_9873,N_5784);
and U12259 (N_12259,N_9231,N_7923);
or U12260 (N_12260,N_5134,N_5668);
or U12261 (N_12261,N_5371,N_5871);
or U12262 (N_12262,N_6464,N_7852);
or U12263 (N_12263,N_5782,N_6462);
nor U12264 (N_12264,N_5665,N_5215);
nor U12265 (N_12265,N_6501,N_8824);
and U12266 (N_12266,N_8878,N_8984);
nand U12267 (N_12267,N_7772,N_5024);
xor U12268 (N_12268,N_9659,N_5545);
nand U12269 (N_12269,N_7151,N_9604);
or U12270 (N_12270,N_9974,N_6119);
xnor U12271 (N_12271,N_5153,N_6072);
and U12272 (N_12272,N_6055,N_7216);
or U12273 (N_12273,N_8696,N_7273);
xor U12274 (N_12274,N_6659,N_8366);
or U12275 (N_12275,N_6267,N_7593);
nand U12276 (N_12276,N_6961,N_7740);
or U12277 (N_12277,N_7664,N_6914);
nand U12278 (N_12278,N_5857,N_5401);
and U12279 (N_12279,N_9440,N_5164);
or U12280 (N_12280,N_7207,N_9213);
and U12281 (N_12281,N_5696,N_6789);
nor U12282 (N_12282,N_6728,N_8765);
or U12283 (N_12283,N_8875,N_9984);
xnor U12284 (N_12284,N_5151,N_8602);
or U12285 (N_12285,N_9549,N_7366);
and U12286 (N_12286,N_6922,N_5162);
and U12287 (N_12287,N_6637,N_8803);
nand U12288 (N_12288,N_7260,N_8249);
xor U12289 (N_12289,N_5392,N_5412);
nand U12290 (N_12290,N_5809,N_9398);
nand U12291 (N_12291,N_9732,N_6923);
and U12292 (N_12292,N_5072,N_8977);
nor U12293 (N_12293,N_6256,N_8482);
nor U12294 (N_12294,N_8811,N_5278);
and U12295 (N_12295,N_8322,N_8084);
nand U12296 (N_12296,N_9441,N_6562);
xnor U12297 (N_12297,N_8645,N_9358);
or U12298 (N_12298,N_8554,N_9463);
or U12299 (N_12299,N_5892,N_5003);
xnor U12300 (N_12300,N_8438,N_5332);
or U12301 (N_12301,N_8243,N_9674);
nand U12302 (N_12302,N_5948,N_6561);
nor U12303 (N_12303,N_6176,N_6827);
xnor U12304 (N_12304,N_9915,N_8766);
xor U12305 (N_12305,N_5541,N_8771);
nor U12306 (N_12306,N_7442,N_7589);
or U12307 (N_12307,N_6358,N_5127);
and U12308 (N_12308,N_8467,N_5607);
and U12309 (N_12309,N_5128,N_5637);
or U12310 (N_12310,N_9730,N_7599);
nor U12311 (N_12311,N_5798,N_6259);
xor U12312 (N_12312,N_7237,N_7055);
nor U12313 (N_12313,N_8177,N_9926);
nand U12314 (N_12314,N_5624,N_6518);
and U12315 (N_12315,N_9723,N_8721);
nand U12316 (N_12316,N_9731,N_5299);
nand U12317 (N_12317,N_9351,N_6492);
and U12318 (N_12318,N_6906,N_8340);
or U12319 (N_12319,N_7489,N_9880);
nor U12320 (N_12320,N_5508,N_7196);
and U12321 (N_12321,N_7563,N_9496);
nor U12322 (N_12322,N_5720,N_8737);
nand U12323 (N_12323,N_5689,N_6183);
and U12324 (N_12324,N_6948,N_6756);
or U12325 (N_12325,N_6147,N_8223);
xnor U12326 (N_12326,N_7806,N_8747);
nand U12327 (N_12327,N_6210,N_9605);
and U12328 (N_12328,N_7158,N_5060);
xor U12329 (N_12329,N_5492,N_6466);
or U12330 (N_12330,N_8848,N_6739);
and U12331 (N_12331,N_7634,N_8662);
nor U12332 (N_12332,N_8789,N_5035);
nand U12333 (N_12333,N_8510,N_9044);
nor U12334 (N_12334,N_5193,N_6441);
nor U12335 (N_12335,N_6493,N_9939);
nand U12336 (N_12336,N_6952,N_5599);
or U12337 (N_12337,N_8265,N_9799);
xor U12338 (N_12338,N_9714,N_6376);
nor U12339 (N_12339,N_5225,N_5646);
xnor U12340 (N_12340,N_8255,N_5452);
nor U12341 (N_12341,N_8335,N_5814);
or U12342 (N_12342,N_6601,N_6614);
or U12343 (N_12343,N_5586,N_6976);
and U12344 (N_12344,N_7172,N_6971);
nor U12345 (N_12345,N_8120,N_9172);
or U12346 (N_12346,N_9807,N_9316);
or U12347 (N_12347,N_9751,N_9914);
nor U12348 (N_12348,N_5473,N_5219);
nor U12349 (N_12349,N_7085,N_5704);
xnor U12350 (N_12350,N_9017,N_6457);
nand U12351 (N_12351,N_9535,N_9970);
and U12352 (N_12352,N_6658,N_7046);
or U12353 (N_12353,N_5146,N_5389);
nand U12354 (N_12354,N_7696,N_9519);
nor U12355 (N_12355,N_5648,N_8560);
nand U12356 (N_12356,N_8454,N_5028);
xor U12357 (N_12357,N_9364,N_9879);
nand U12358 (N_12358,N_6010,N_5089);
nand U12359 (N_12359,N_8626,N_9040);
or U12360 (N_12360,N_5416,N_9156);
nor U12361 (N_12361,N_9434,N_7666);
nor U12362 (N_12362,N_8999,N_9305);
or U12363 (N_12363,N_8798,N_5951);
and U12364 (N_12364,N_8758,N_5837);
xor U12365 (N_12365,N_7670,N_6312);
nor U12366 (N_12366,N_5226,N_7892);
or U12367 (N_12367,N_7429,N_6965);
xor U12368 (N_12368,N_6184,N_7556);
nand U12369 (N_12369,N_8805,N_5283);
nand U12370 (N_12370,N_8371,N_6498);
nor U12371 (N_12371,N_9628,N_7523);
xnor U12372 (N_12372,N_9228,N_5500);
nor U12373 (N_12373,N_6413,N_5900);
nor U12374 (N_12374,N_9517,N_8125);
or U12375 (N_12375,N_8665,N_9998);
nor U12376 (N_12376,N_9292,N_7425);
or U12377 (N_12377,N_6804,N_6813);
xor U12378 (N_12378,N_5753,N_6998);
or U12379 (N_12379,N_9167,N_5653);
or U12380 (N_12380,N_6148,N_6941);
nor U12381 (N_12381,N_5103,N_6738);
xnor U12382 (N_12382,N_9342,N_9652);
and U12383 (N_12383,N_5635,N_5938);
nor U12384 (N_12384,N_5601,N_7316);
xor U12385 (N_12385,N_6171,N_9412);
nor U12386 (N_12386,N_7765,N_8015);
nand U12387 (N_12387,N_7364,N_5803);
or U12388 (N_12388,N_8099,N_9073);
and U12389 (N_12389,N_5520,N_8124);
or U12390 (N_12390,N_7691,N_6167);
and U12391 (N_12391,N_9427,N_9921);
xor U12392 (N_12392,N_5869,N_5942);
and U12393 (N_12393,N_7642,N_7295);
xor U12394 (N_12394,N_9022,N_9871);
or U12395 (N_12395,N_6157,N_7701);
and U12396 (N_12396,N_7146,N_9973);
nand U12397 (N_12397,N_5897,N_6077);
or U12398 (N_12398,N_9376,N_9010);
xnor U12399 (N_12399,N_7190,N_8684);
and U12400 (N_12400,N_8062,N_6947);
nor U12401 (N_12401,N_8136,N_9368);
and U12402 (N_12402,N_6404,N_6101);
nand U12403 (N_12403,N_8151,N_6698);
or U12404 (N_12404,N_6400,N_7454);
or U12405 (N_12405,N_6043,N_7070);
xor U12406 (N_12406,N_7989,N_9135);
and U12407 (N_12407,N_8359,N_5455);
xor U12408 (N_12408,N_8674,N_7746);
xor U12409 (N_12409,N_8028,N_9432);
or U12410 (N_12410,N_6764,N_9856);
nand U12411 (N_12411,N_5497,N_7441);
nor U12412 (N_12412,N_9875,N_9808);
or U12413 (N_12413,N_5918,N_9195);
and U12414 (N_12414,N_5768,N_7900);
nand U12415 (N_12415,N_9287,N_8330);
nand U12416 (N_12416,N_7232,N_5117);
or U12417 (N_12417,N_8632,N_6447);
xnor U12418 (N_12418,N_5514,N_5036);
xnor U12419 (N_12419,N_6891,N_8767);
or U12420 (N_12420,N_5673,N_7797);
nand U12421 (N_12421,N_8633,N_7646);
or U12422 (N_12422,N_7671,N_6519);
or U12423 (N_12423,N_5217,N_6328);
nor U12424 (N_12424,N_7838,N_6838);
nand U12425 (N_12425,N_8441,N_9408);
nand U12426 (N_12426,N_9204,N_9559);
xor U12427 (N_12427,N_8321,N_9356);
nor U12428 (N_12428,N_6366,N_5715);
nand U12429 (N_12429,N_9067,N_9500);
nor U12430 (N_12430,N_9623,N_8549);
and U12431 (N_12431,N_8853,N_5851);
xor U12432 (N_12432,N_9971,N_5883);
or U12433 (N_12433,N_8567,N_8100);
and U12434 (N_12434,N_9372,N_5289);
xor U12435 (N_12435,N_6003,N_5194);
nor U12436 (N_12436,N_7418,N_5391);
or U12437 (N_12437,N_9979,N_7356);
or U12438 (N_12438,N_9306,N_7850);
xnor U12439 (N_12439,N_9969,N_6133);
nor U12440 (N_12440,N_7434,N_9766);
nand U12441 (N_12441,N_8477,N_5531);
nand U12442 (N_12442,N_5478,N_7086);
or U12443 (N_12443,N_5204,N_6144);
and U12444 (N_12444,N_7375,N_7402);
or U12445 (N_12445,N_8292,N_8116);
and U12446 (N_12446,N_8904,N_7087);
xnor U12447 (N_12447,N_5038,N_8837);
or U12448 (N_12448,N_6690,N_6661);
nor U12449 (N_12449,N_9948,N_9512);
and U12450 (N_12450,N_8106,N_5387);
nand U12451 (N_12451,N_8667,N_8836);
or U12452 (N_12452,N_8040,N_9311);
nor U12453 (N_12453,N_8212,N_8382);
xor U12454 (N_12454,N_7805,N_8911);
nor U12455 (N_12455,N_9396,N_6253);
nor U12456 (N_12456,N_5047,N_7856);
and U12457 (N_12457,N_6300,N_9284);
or U12458 (N_12458,N_7843,N_6740);
or U12459 (N_12459,N_7584,N_5622);
nand U12460 (N_12460,N_7844,N_8066);
or U12461 (N_12461,N_8461,N_8480);
nor U12462 (N_12462,N_6910,N_7577);
and U12463 (N_12463,N_5463,N_6734);
nor U12464 (N_12464,N_7420,N_9713);
or U12465 (N_12465,N_7783,N_7978);
and U12466 (N_12466,N_9824,N_7360);
nand U12467 (N_12467,N_6234,N_5974);
or U12468 (N_12468,N_5730,N_5916);
xor U12469 (N_12469,N_6383,N_9771);
xor U12470 (N_12470,N_8862,N_6880);
nor U12471 (N_12471,N_5655,N_9353);
nor U12472 (N_12472,N_6411,N_5940);
xnor U12473 (N_12473,N_8456,N_9477);
nor U12474 (N_12474,N_6486,N_5729);
or U12475 (N_12475,N_5595,N_6235);
and U12476 (N_12476,N_5559,N_8261);
nand U12477 (N_12477,N_8075,N_9850);
nand U12478 (N_12478,N_5764,N_9074);
and U12479 (N_12479,N_5385,N_6761);
and U12480 (N_12480,N_7568,N_6602);
xor U12481 (N_12481,N_8916,N_6421);
and U12482 (N_12482,N_9157,N_8204);
and U12483 (N_12483,N_7362,N_5618);
and U12484 (N_12484,N_8964,N_6274);
nor U12485 (N_12485,N_7655,N_5121);
nand U12486 (N_12486,N_5081,N_5280);
nor U12487 (N_12487,N_7702,N_8563);
and U12488 (N_12488,N_5889,N_8272);
nand U12489 (N_12489,N_7045,N_8756);
nor U12490 (N_12490,N_6532,N_9787);
nor U12491 (N_12491,N_6015,N_9557);
nor U12492 (N_12492,N_7497,N_5355);
xor U12493 (N_12493,N_7211,N_8088);
or U12494 (N_12494,N_8038,N_6410);
or U12495 (N_12495,N_7096,N_6704);
and U12496 (N_12496,N_9443,N_5143);
nand U12497 (N_12497,N_6399,N_7798);
or U12498 (N_12498,N_8337,N_5638);
or U12499 (N_12499,N_5832,N_7380);
or U12500 (N_12500,N_9774,N_7785);
nand U12501 (N_12501,N_7486,N_8981);
and U12502 (N_12502,N_5343,N_5400);
and U12503 (N_12503,N_7274,N_6409);
nor U12504 (N_12504,N_7008,N_5166);
nand U12505 (N_12505,N_6111,N_9047);
nor U12506 (N_12506,N_6559,N_8772);
nand U12507 (N_12507,N_5621,N_8526);
and U12508 (N_12508,N_5266,N_9514);
nand U12509 (N_12509,N_7052,N_6725);
or U12510 (N_12510,N_8295,N_8325);
nand U12511 (N_12511,N_9937,N_6673);
nand U12512 (N_12512,N_8368,N_5825);
nor U12513 (N_12513,N_8540,N_5016);
and U12514 (N_12514,N_6644,N_8946);
nand U12515 (N_12515,N_9571,N_9697);
or U12516 (N_12516,N_8026,N_9845);
or U12517 (N_12517,N_8973,N_9122);
nor U12518 (N_12518,N_8550,N_8224);
xnor U12519 (N_12519,N_7184,N_5601);
or U12520 (N_12520,N_9899,N_9965);
xor U12521 (N_12521,N_9820,N_9535);
nand U12522 (N_12522,N_9799,N_6863);
xor U12523 (N_12523,N_8544,N_8752);
or U12524 (N_12524,N_9466,N_9710);
nor U12525 (N_12525,N_9410,N_8659);
or U12526 (N_12526,N_6587,N_7331);
nand U12527 (N_12527,N_9484,N_9838);
or U12528 (N_12528,N_6587,N_9634);
and U12529 (N_12529,N_7067,N_8935);
xnor U12530 (N_12530,N_8175,N_9020);
or U12531 (N_12531,N_7391,N_9899);
nor U12532 (N_12532,N_5266,N_7549);
and U12533 (N_12533,N_5555,N_6134);
xnor U12534 (N_12534,N_6842,N_8351);
xnor U12535 (N_12535,N_6793,N_8755);
xnor U12536 (N_12536,N_9665,N_8581);
or U12537 (N_12537,N_9039,N_8494);
xor U12538 (N_12538,N_8650,N_5984);
and U12539 (N_12539,N_6970,N_6749);
and U12540 (N_12540,N_6153,N_6564);
nand U12541 (N_12541,N_7183,N_7982);
or U12542 (N_12542,N_5012,N_8356);
nor U12543 (N_12543,N_8433,N_8055);
nor U12544 (N_12544,N_7805,N_6373);
or U12545 (N_12545,N_9085,N_5117);
or U12546 (N_12546,N_8928,N_9651);
and U12547 (N_12547,N_7314,N_9322);
nor U12548 (N_12548,N_8093,N_9249);
and U12549 (N_12549,N_9859,N_7389);
xor U12550 (N_12550,N_5414,N_5043);
nor U12551 (N_12551,N_8862,N_6540);
and U12552 (N_12552,N_6496,N_9560);
nand U12553 (N_12553,N_8237,N_9119);
xor U12554 (N_12554,N_8656,N_8600);
xor U12555 (N_12555,N_9286,N_7919);
nand U12556 (N_12556,N_5058,N_8971);
xnor U12557 (N_12557,N_9484,N_9495);
nand U12558 (N_12558,N_9466,N_8915);
xnor U12559 (N_12559,N_6723,N_8162);
nand U12560 (N_12560,N_8150,N_9049);
nor U12561 (N_12561,N_7727,N_8355);
xor U12562 (N_12562,N_5247,N_5664);
nor U12563 (N_12563,N_5812,N_7041);
or U12564 (N_12564,N_7342,N_8553);
and U12565 (N_12565,N_5234,N_5149);
xor U12566 (N_12566,N_7838,N_5686);
and U12567 (N_12567,N_7317,N_6067);
or U12568 (N_12568,N_9316,N_5822);
and U12569 (N_12569,N_7101,N_5510);
or U12570 (N_12570,N_9454,N_6095);
nor U12571 (N_12571,N_7584,N_8599);
nor U12572 (N_12572,N_8347,N_9208);
nand U12573 (N_12573,N_9021,N_8254);
or U12574 (N_12574,N_9469,N_9043);
nand U12575 (N_12575,N_5644,N_9927);
nor U12576 (N_12576,N_5813,N_8048);
nand U12577 (N_12577,N_5858,N_5159);
or U12578 (N_12578,N_5625,N_8939);
xnor U12579 (N_12579,N_5492,N_6276);
and U12580 (N_12580,N_9233,N_6020);
nor U12581 (N_12581,N_6827,N_6436);
nor U12582 (N_12582,N_5050,N_7386);
nor U12583 (N_12583,N_9281,N_9818);
nand U12584 (N_12584,N_7205,N_9563);
xnor U12585 (N_12585,N_9358,N_7581);
or U12586 (N_12586,N_5022,N_9710);
or U12587 (N_12587,N_6945,N_6064);
nand U12588 (N_12588,N_6567,N_6759);
and U12589 (N_12589,N_5939,N_8415);
nor U12590 (N_12590,N_9731,N_8375);
or U12591 (N_12591,N_9238,N_8042);
nand U12592 (N_12592,N_8717,N_5813);
and U12593 (N_12593,N_8521,N_9460);
nor U12594 (N_12594,N_5227,N_6644);
nor U12595 (N_12595,N_5213,N_9274);
or U12596 (N_12596,N_8901,N_5091);
or U12597 (N_12597,N_6494,N_5497);
xor U12598 (N_12598,N_9384,N_6165);
nor U12599 (N_12599,N_5995,N_9039);
nor U12600 (N_12600,N_6116,N_8859);
and U12601 (N_12601,N_5845,N_5570);
nand U12602 (N_12602,N_8912,N_7873);
nor U12603 (N_12603,N_9207,N_8451);
and U12604 (N_12604,N_8343,N_9687);
and U12605 (N_12605,N_9219,N_8941);
or U12606 (N_12606,N_5458,N_6858);
nor U12607 (N_12607,N_9002,N_9402);
xor U12608 (N_12608,N_6511,N_9588);
and U12609 (N_12609,N_5145,N_8693);
and U12610 (N_12610,N_8693,N_7873);
nand U12611 (N_12611,N_8467,N_8907);
or U12612 (N_12612,N_7508,N_9436);
xnor U12613 (N_12613,N_9561,N_6841);
xnor U12614 (N_12614,N_8895,N_8560);
xor U12615 (N_12615,N_6855,N_5791);
nor U12616 (N_12616,N_8581,N_8751);
xnor U12617 (N_12617,N_6257,N_6618);
xnor U12618 (N_12618,N_7718,N_6011);
and U12619 (N_12619,N_5331,N_7510);
nand U12620 (N_12620,N_8055,N_9469);
or U12621 (N_12621,N_6189,N_8474);
nor U12622 (N_12622,N_8691,N_6839);
or U12623 (N_12623,N_6455,N_8683);
nand U12624 (N_12624,N_6348,N_9032);
nor U12625 (N_12625,N_8756,N_5555);
nor U12626 (N_12626,N_9227,N_7190);
xnor U12627 (N_12627,N_8089,N_8489);
or U12628 (N_12628,N_7553,N_5504);
and U12629 (N_12629,N_8441,N_5702);
or U12630 (N_12630,N_6858,N_9619);
nand U12631 (N_12631,N_8834,N_9842);
nor U12632 (N_12632,N_6921,N_8222);
and U12633 (N_12633,N_6771,N_7772);
and U12634 (N_12634,N_6384,N_5500);
nor U12635 (N_12635,N_7136,N_9676);
nand U12636 (N_12636,N_8217,N_5254);
or U12637 (N_12637,N_9264,N_9328);
xor U12638 (N_12638,N_8752,N_8910);
nor U12639 (N_12639,N_5483,N_7556);
or U12640 (N_12640,N_9048,N_7821);
and U12641 (N_12641,N_6162,N_7883);
and U12642 (N_12642,N_8037,N_9970);
nand U12643 (N_12643,N_8312,N_6746);
xor U12644 (N_12644,N_8850,N_5119);
xnor U12645 (N_12645,N_7300,N_7647);
nor U12646 (N_12646,N_5714,N_9461);
and U12647 (N_12647,N_8751,N_5135);
or U12648 (N_12648,N_7107,N_7847);
xor U12649 (N_12649,N_5384,N_5689);
xnor U12650 (N_12650,N_6733,N_8592);
nand U12651 (N_12651,N_8944,N_7101);
or U12652 (N_12652,N_7310,N_5060);
and U12653 (N_12653,N_9317,N_9167);
nand U12654 (N_12654,N_5316,N_8467);
or U12655 (N_12655,N_9196,N_9162);
and U12656 (N_12656,N_6343,N_6474);
and U12657 (N_12657,N_6619,N_9920);
and U12658 (N_12658,N_5433,N_7695);
and U12659 (N_12659,N_5205,N_5499);
xnor U12660 (N_12660,N_5057,N_8092);
or U12661 (N_12661,N_5703,N_8106);
or U12662 (N_12662,N_9792,N_9878);
and U12663 (N_12663,N_9529,N_5387);
xor U12664 (N_12664,N_9078,N_6613);
and U12665 (N_12665,N_8589,N_7604);
nor U12666 (N_12666,N_7689,N_6334);
nor U12667 (N_12667,N_8619,N_5156);
and U12668 (N_12668,N_8321,N_7523);
xor U12669 (N_12669,N_6180,N_5412);
or U12670 (N_12670,N_9173,N_5074);
and U12671 (N_12671,N_7405,N_6154);
nor U12672 (N_12672,N_8050,N_7147);
or U12673 (N_12673,N_7327,N_8231);
and U12674 (N_12674,N_8734,N_8196);
or U12675 (N_12675,N_9883,N_8365);
xor U12676 (N_12676,N_9196,N_9010);
or U12677 (N_12677,N_6665,N_5794);
nand U12678 (N_12678,N_9695,N_5647);
nor U12679 (N_12679,N_8701,N_8197);
and U12680 (N_12680,N_6633,N_6341);
xnor U12681 (N_12681,N_7962,N_9989);
xor U12682 (N_12682,N_9165,N_7719);
and U12683 (N_12683,N_6887,N_6548);
nor U12684 (N_12684,N_9940,N_7226);
nor U12685 (N_12685,N_8805,N_6526);
xor U12686 (N_12686,N_8517,N_5937);
and U12687 (N_12687,N_8708,N_5182);
nor U12688 (N_12688,N_8182,N_5042);
or U12689 (N_12689,N_6575,N_7450);
or U12690 (N_12690,N_8712,N_5521);
nand U12691 (N_12691,N_6077,N_9758);
nor U12692 (N_12692,N_6469,N_9909);
nor U12693 (N_12693,N_5780,N_6311);
or U12694 (N_12694,N_8959,N_5197);
nor U12695 (N_12695,N_5386,N_6031);
nor U12696 (N_12696,N_8486,N_7512);
nand U12697 (N_12697,N_7107,N_6236);
nand U12698 (N_12698,N_8971,N_9677);
xnor U12699 (N_12699,N_5321,N_8853);
xnor U12700 (N_12700,N_8217,N_6966);
xnor U12701 (N_12701,N_5768,N_9065);
and U12702 (N_12702,N_6341,N_7899);
xor U12703 (N_12703,N_5123,N_8936);
and U12704 (N_12704,N_5632,N_8709);
nor U12705 (N_12705,N_5218,N_5106);
or U12706 (N_12706,N_7590,N_6207);
nor U12707 (N_12707,N_6105,N_6489);
xor U12708 (N_12708,N_5375,N_5274);
and U12709 (N_12709,N_5645,N_6441);
nand U12710 (N_12710,N_6190,N_5401);
and U12711 (N_12711,N_8483,N_8077);
xor U12712 (N_12712,N_7710,N_9267);
nor U12713 (N_12713,N_8451,N_5687);
nand U12714 (N_12714,N_5287,N_7100);
nand U12715 (N_12715,N_8515,N_6960);
or U12716 (N_12716,N_6359,N_8392);
nand U12717 (N_12717,N_9339,N_9175);
xnor U12718 (N_12718,N_7108,N_8322);
nand U12719 (N_12719,N_8060,N_8131);
or U12720 (N_12720,N_6753,N_9293);
nor U12721 (N_12721,N_9475,N_5438);
or U12722 (N_12722,N_8643,N_5063);
nor U12723 (N_12723,N_9016,N_7676);
and U12724 (N_12724,N_5082,N_6523);
nor U12725 (N_12725,N_7067,N_9233);
nor U12726 (N_12726,N_8396,N_5984);
nor U12727 (N_12727,N_7323,N_6524);
nand U12728 (N_12728,N_8117,N_7903);
or U12729 (N_12729,N_5586,N_9252);
and U12730 (N_12730,N_5423,N_8263);
xor U12731 (N_12731,N_8411,N_9035);
xnor U12732 (N_12732,N_6622,N_5466);
and U12733 (N_12733,N_6176,N_6725);
nand U12734 (N_12734,N_5943,N_7495);
nor U12735 (N_12735,N_9106,N_5398);
xnor U12736 (N_12736,N_6119,N_9666);
and U12737 (N_12737,N_7543,N_8563);
and U12738 (N_12738,N_7784,N_5491);
and U12739 (N_12739,N_7042,N_5431);
nor U12740 (N_12740,N_6659,N_6572);
and U12741 (N_12741,N_5482,N_6939);
xnor U12742 (N_12742,N_5122,N_8386);
and U12743 (N_12743,N_5222,N_8044);
xor U12744 (N_12744,N_7741,N_9334);
and U12745 (N_12745,N_8211,N_6575);
or U12746 (N_12746,N_6625,N_9935);
and U12747 (N_12747,N_5068,N_9247);
nor U12748 (N_12748,N_8839,N_5932);
nand U12749 (N_12749,N_9289,N_9462);
nor U12750 (N_12750,N_5189,N_8962);
and U12751 (N_12751,N_6903,N_6008);
nor U12752 (N_12752,N_5828,N_9857);
and U12753 (N_12753,N_7117,N_6824);
nor U12754 (N_12754,N_9019,N_5685);
and U12755 (N_12755,N_7587,N_9919);
and U12756 (N_12756,N_6649,N_8467);
xnor U12757 (N_12757,N_5798,N_9572);
nand U12758 (N_12758,N_5281,N_6979);
nand U12759 (N_12759,N_9975,N_7384);
xor U12760 (N_12760,N_7624,N_7256);
and U12761 (N_12761,N_7014,N_7479);
and U12762 (N_12762,N_6788,N_8938);
nand U12763 (N_12763,N_9897,N_6684);
and U12764 (N_12764,N_6756,N_5167);
xnor U12765 (N_12765,N_6143,N_6528);
nor U12766 (N_12766,N_6214,N_9849);
xor U12767 (N_12767,N_5580,N_8031);
and U12768 (N_12768,N_9662,N_9819);
and U12769 (N_12769,N_9592,N_9123);
nor U12770 (N_12770,N_8062,N_7761);
or U12771 (N_12771,N_6559,N_8012);
nand U12772 (N_12772,N_9562,N_9795);
or U12773 (N_12773,N_6455,N_5037);
nand U12774 (N_12774,N_9523,N_6248);
or U12775 (N_12775,N_8225,N_6472);
nand U12776 (N_12776,N_6759,N_5718);
or U12777 (N_12777,N_6781,N_9737);
and U12778 (N_12778,N_7261,N_6864);
or U12779 (N_12779,N_9689,N_8312);
and U12780 (N_12780,N_7690,N_5572);
nand U12781 (N_12781,N_5208,N_8002);
and U12782 (N_12782,N_7075,N_9120);
nor U12783 (N_12783,N_5309,N_7404);
and U12784 (N_12784,N_8424,N_8233);
or U12785 (N_12785,N_7148,N_8799);
and U12786 (N_12786,N_9106,N_9865);
and U12787 (N_12787,N_9362,N_7554);
nor U12788 (N_12788,N_6939,N_5727);
or U12789 (N_12789,N_7532,N_5630);
nand U12790 (N_12790,N_9786,N_6785);
and U12791 (N_12791,N_7843,N_6053);
nand U12792 (N_12792,N_8206,N_6697);
and U12793 (N_12793,N_9822,N_9983);
xor U12794 (N_12794,N_5693,N_5912);
nor U12795 (N_12795,N_5935,N_5051);
nor U12796 (N_12796,N_6725,N_5273);
or U12797 (N_12797,N_9092,N_8753);
nor U12798 (N_12798,N_6706,N_5119);
nand U12799 (N_12799,N_7484,N_6032);
nor U12800 (N_12800,N_8622,N_9436);
and U12801 (N_12801,N_8085,N_8748);
xor U12802 (N_12802,N_5685,N_7250);
or U12803 (N_12803,N_9202,N_6130);
nor U12804 (N_12804,N_8996,N_6195);
or U12805 (N_12805,N_7640,N_6999);
nor U12806 (N_12806,N_9853,N_6544);
or U12807 (N_12807,N_8817,N_5458);
nor U12808 (N_12808,N_6316,N_8794);
nor U12809 (N_12809,N_6583,N_7001);
nor U12810 (N_12810,N_8946,N_6815);
and U12811 (N_12811,N_7437,N_5045);
xor U12812 (N_12812,N_9353,N_8152);
nand U12813 (N_12813,N_8213,N_6393);
or U12814 (N_12814,N_8196,N_8804);
xnor U12815 (N_12815,N_6220,N_5945);
xor U12816 (N_12816,N_7015,N_9834);
nand U12817 (N_12817,N_7941,N_9811);
or U12818 (N_12818,N_5538,N_6564);
nand U12819 (N_12819,N_6181,N_9810);
nor U12820 (N_12820,N_9930,N_6494);
xor U12821 (N_12821,N_7021,N_9872);
nand U12822 (N_12822,N_6847,N_8698);
and U12823 (N_12823,N_7954,N_8756);
or U12824 (N_12824,N_6074,N_8702);
nand U12825 (N_12825,N_9410,N_7071);
nand U12826 (N_12826,N_7784,N_9070);
and U12827 (N_12827,N_6657,N_7685);
xor U12828 (N_12828,N_6885,N_6653);
nor U12829 (N_12829,N_8610,N_9894);
xor U12830 (N_12830,N_7516,N_5044);
or U12831 (N_12831,N_8429,N_8123);
and U12832 (N_12832,N_5176,N_9247);
nor U12833 (N_12833,N_6135,N_8945);
nor U12834 (N_12834,N_9148,N_8571);
and U12835 (N_12835,N_5990,N_9643);
nor U12836 (N_12836,N_9756,N_6762);
and U12837 (N_12837,N_5892,N_8044);
or U12838 (N_12838,N_9912,N_8478);
or U12839 (N_12839,N_9461,N_9265);
nand U12840 (N_12840,N_5445,N_5253);
and U12841 (N_12841,N_8468,N_7743);
nor U12842 (N_12842,N_8195,N_9725);
nor U12843 (N_12843,N_8294,N_6472);
or U12844 (N_12844,N_9181,N_6159);
or U12845 (N_12845,N_6490,N_9854);
or U12846 (N_12846,N_7330,N_8825);
xor U12847 (N_12847,N_5302,N_9694);
and U12848 (N_12848,N_6860,N_8297);
or U12849 (N_12849,N_9125,N_9416);
nor U12850 (N_12850,N_6648,N_6249);
nor U12851 (N_12851,N_8961,N_9476);
xnor U12852 (N_12852,N_7203,N_9020);
xnor U12853 (N_12853,N_9079,N_9779);
nor U12854 (N_12854,N_8766,N_7811);
nor U12855 (N_12855,N_9238,N_5974);
nand U12856 (N_12856,N_5175,N_9881);
or U12857 (N_12857,N_5859,N_6539);
and U12858 (N_12858,N_8468,N_6971);
nand U12859 (N_12859,N_7253,N_5544);
nor U12860 (N_12860,N_9166,N_6669);
or U12861 (N_12861,N_7071,N_9086);
nand U12862 (N_12862,N_9648,N_9339);
xor U12863 (N_12863,N_8982,N_6792);
nand U12864 (N_12864,N_5970,N_6983);
or U12865 (N_12865,N_5059,N_9985);
xor U12866 (N_12866,N_5916,N_7184);
nand U12867 (N_12867,N_9304,N_8987);
xnor U12868 (N_12868,N_6540,N_5449);
or U12869 (N_12869,N_7276,N_7386);
nand U12870 (N_12870,N_6944,N_9452);
or U12871 (N_12871,N_9241,N_9143);
xnor U12872 (N_12872,N_6039,N_5573);
xnor U12873 (N_12873,N_9939,N_9271);
or U12874 (N_12874,N_7683,N_5788);
and U12875 (N_12875,N_8933,N_8223);
and U12876 (N_12876,N_7682,N_9419);
or U12877 (N_12877,N_6605,N_5841);
or U12878 (N_12878,N_7718,N_6391);
nor U12879 (N_12879,N_9063,N_7027);
nor U12880 (N_12880,N_6745,N_6073);
xor U12881 (N_12881,N_8263,N_6273);
nor U12882 (N_12882,N_5154,N_8274);
nor U12883 (N_12883,N_8938,N_9577);
xnor U12884 (N_12884,N_9607,N_9403);
nor U12885 (N_12885,N_5475,N_9298);
xor U12886 (N_12886,N_7051,N_6089);
nor U12887 (N_12887,N_7254,N_7853);
xor U12888 (N_12888,N_9736,N_9934);
nand U12889 (N_12889,N_6517,N_8686);
nand U12890 (N_12890,N_5054,N_8274);
or U12891 (N_12891,N_5460,N_6806);
or U12892 (N_12892,N_7355,N_5906);
nand U12893 (N_12893,N_5552,N_7924);
nor U12894 (N_12894,N_6039,N_5497);
and U12895 (N_12895,N_8774,N_8075);
xor U12896 (N_12896,N_6241,N_8624);
and U12897 (N_12897,N_9144,N_6688);
xor U12898 (N_12898,N_8510,N_7054);
and U12899 (N_12899,N_9765,N_5276);
xor U12900 (N_12900,N_9487,N_7517);
nor U12901 (N_12901,N_9301,N_7731);
and U12902 (N_12902,N_9812,N_8335);
and U12903 (N_12903,N_6855,N_6024);
and U12904 (N_12904,N_9477,N_5887);
nor U12905 (N_12905,N_8196,N_8523);
nor U12906 (N_12906,N_7039,N_6657);
nand U12907 (N_12907,N_7972,N_8952);
nand U12908 (N_12908,N_5818,N_7165);
nand U12909 (N_12909,N_6475,N_6269);
nand U12910 (N_12910,N_6998,N_7308);
nand U12911 (N_12911,N_6520,N_5070);
nor U12912 (N_12912,N_9029,N_8259);
or U12913 (N_12913,N_8887,N_6404);
or U12914 (N_12914,N_5071,N_7729);
or U12915 (N_12915,N_8475,N_9473);
and U12916 (N_12916,N_5546,N_6429);
nand U12917 (N_12917,N_7627,N_8339);
xnor U12918 (N_12918,N_6705,N_5452);
xor U12919 (N_12919,N_9648,N_8907);
nand U12920 (N_12920,N_6590,N_9599);
and U12921 (N_12921,N_9455,N_5374);
nand U12922 (N_12922,N_6743,N_8068);
or U12923 (N_12923,N_8113,N_7738);
or U12924 (N_12924,N_8720,N_7223);
nand U12925 (N_12925,N_5293,N_7384);
and U12926 (N_12926,N_7411,N_9113);
nor U12927 (N_12927,N_8690,N_6410);
nand U12928 (N_12928,N_6447,N_9941);
or U12929 (N_12929,N_5090,N_9775);
xor U12930 (N_12930,N_9050,N_5495);
and U12931 (N_12931,N_6453,N_8069);
xor U12932 (N_12932,N_5065,N_7497);
and U12933 (N_12933,N_6213,N_9929);
nand U12934 (N_12934,N_8466,N_5694);
xor U12935 (N_12935,N_9670,N_9035);
or U12936 (N_12936,N_8972,N_6348);
or U12937 (N_12937,N_5709,N_5133);
nor U12938 (N_12938,N_7964,N_9568);
nand U12939 (N_12939,N_6636,N_9189);
nand U12940 (N_12940,N_8133,N_7649);
and U12941 (N_12941,N_5065,N_8205);
or U12942 (N_12942,N_7272,N_8961);
and U12943 (N_12943,N_8163,N_8858);
or U12944 (N_12944,N_5722,N_7631);
nor U12945 (N_12945,N_5157,N_6500);
nor U12946 (N_12946,N_9332,N_9952);
nand U12947 (N_12947,N_6131,N_5879);
and U12948 (N_12948,N_5457,N_9940);
and U12949 (N_12949,N_6885,N_5912);
nand U12950 (N_12950,N_8153,N_6037);
nor U12951 (N_12951,N_5308,N_8914);
nand U12952 (N_12952,N_9996,N_6817);
nor U12953 (N_12953,N_8020,N_7753);
xor U12954 (N_12954,N_9815,N_5797);
nand U12955 (N_12955,N_5342,N_9402);
or U12956 (N_12956,N_6123,N_7093);
xnor U12957 (N_12957,N_6755,N_8089);
nand U12958 (N_12958,N_5533,N_8824);
nor U12959 (N_12959,N_5039,N_8722);
and U12960 (N_12960,N_9545,N_6294);
and U12961 (N_12961,N_5639,N_5276);
nand U12962 (N_12962,N_8221,N_9602);
nor U12963 (N_12963,N_8523,N_5878);
xnor U12964 (N_12964,N_9398,N_6523);
nand U12965 (N_12965,N_9472,N_8914);
and U12966 (N_12966,N_7967,N_7547);
xor U12967 (N_12967,N_7771,N_9346);
nor U12968 (N_12968,N_9639,N_5608);
or U12969 (N_12969,N_7727,N_7801);
or U12970 (N_12970,N_6439,N_5060);
and U12971 (N_12971,N_7824,N_7766);
nor U12972 (N_12972,N_8940,N_7612);
nand U12973 (N_12973,N_6191,N_7184);
nor U12974 (N_12974,N_5073,N_5626);
xor U12975 (N_12975,N_7215,N_6595);
nand U12976 (N_12976,N_9144,N_5266);
xnor U12977 (N_12977,N_7859,N_6078);
and U12978 (N_12978,N_6396,N_7994);
nor U12979 (N_12979,N_8552,N_6089);
nand U12980 (N_12980,N_6274,N_6509);
nand U12981 (N_12981,N_9192,N_8831);
xor U12982 (N_12982,N_7218,N_6861);
nand U12983 (N_12983,N_5140,N_6265);
or U12984 (N_12984,N_8170,N_6856);
nor U12985 (N_12985,N_9797,N_6338);
or U12986 (N_12986,N_7393,N_7988);
and U12987 (N_12987,N_6766,N_6632);
or U12988 (N_12988,N_6387,N_5138);
xor U12989 (N_12989,N_9986,N_7678);
nor U12990 (N_12990,N_5239,N_8508);
nand U12991 (N_12991,N_5287,N_8721);
and U12992 (N_12992,N_5943,N_7799);
or U12993 (N_12993,N_9147,N_8992);
nand U12994 (N_12994,N_6681,N_5243);
and U12995 (N_12995,N_8718,N_5170);
or U12996 (N_12996,N_5856,N_8587);
nor U12997 (N_12997,N_5799,N_8328);
nand U12998 (N_12998,N_7023,N_5407);
nand U12999 (N_12999,N_6454,N_6908);
nand U13000 (N_13000,N_8343,N_6651);
and U13001 (N_13001,N_6763,N_6799);
xor U13002 (N_13002,N_9349,N_8038);
xnor U13003 (N_13003,N_7860,N_5591);
and U13004 (N_13004,N_7503,N_7907);
nand U13005 (N_13005,N_7105,N_9407);
nand U13006 (N_13006,N_8737,N_5144);
nor U13007 (N_13007,N_8685,N_8417);
and U13008 (N_13008,N_9113,N_6142);
or U13009 (N_13009,N_7056,N_8082);
xnor U13010 (N_13010,N_8816,N_5609);
nor U13011 (N_13011,N_8860,N_9337);
xnor U13012 (N_13012,N_6667,N_7605);
nand U13013 (N_13013,N_6583,N_9106);
xor U13014 (N_13014,N_6181,N_8011);
xnor U13015 (N_13015,N_7870,N_5737);
and U13016 (N_13016,N_8857,N_6859);
or U13017 (N_13017,N_5986,N_8239);
or U13018 (N_13018,N_9185,N_5654);
xor U13019 (N_13019,N_7573,N_6057);
nor U13020 (N_13020,N_6547,N_5252);
nand U13021 (N_13021,N_9007,N_9204);
and U13022 (N_13022,N_6465,N_9026);
and U13023 (N_13023,N_5310,N_9235);
nand U13024 (N_13024,N_6028,N_8722);
nand U13025 (N_13025,N_9487,N_9650);
nor U13026 (N_13026,N_7757,N_5337);
xor U13027 (N_13027,N_7766,N_8973);
or U13028 (N_13028,N_6420,N_7156);
xor U13029 (N_13029,N_9870,N_6854);
nor U13030 (N_13030,N_8216,N_8114);
or U13031 (N_13031,N_9577,N_8216);
or U13032 (N_13032,N_6592,N_6387);
nand U13033 (N_13033,N_8148,N_9627);
nor U13034 (N_13034,N_5852,N_9039);
nand U13035 (N_13035,N_5904,N_9832);
xor U13036 (N_13036,N_5526,N_8445);
xnor U13037 (N_13037,N_9655,N_7217);
nand U13038 (N_13038,N_8129,N_8270);
and U13039 (N_13039,N_5500,N_8574);
and U13040 (N_13040,N_6844,N_8848);
xnor U13041 (N_13041,N_9597,N_7676);
nor U13042 (N_13042,N_8461,N_7939);
or U13043 (N_13043,N_6888,N_5779);
nand U13044 (N_13044,N_6692,N_9919);
xor U13045 (N_13045,N_8481,N_7008);
nand U13046 (N_13046,N_7815,N_8562);
nor U13047 (N_13047,N_5091,N_7790);
nor U13048 (N_13048,N_5370,N_5867);
nor U13049 (N_13049,N_5475,N_7694);
nand U13050 (N_13050,N_9657,N_6007);
xnor U13051 (N_13051,N_6245,N_7871);
xnor U13052 (N_13052,N_8322,N_9288);
nor U13053 (N_13053,N_8928,N_7734);
or U13054 (N_13054,N_9550,N_9818);
nor U13055 (N_13055,N_8410,N_6420);
nor U13056 (N_13056,N_8634,N_6644);
nor U13057 (N_13057,N_5501,N_7943);
xor U13058 (N_13058,N_5360,N_9068);
nand U13059 (N_13059,N_9235,N_8775);
xnor U13060 (N_13060,N_6667,N_9244);
or U13061 (N_13061,N_5731,N_7752);
and U13062 (N_13062,N_5077,N_7025);
or U13063 (N_13063,N_5692,N_9315);
nand U13064 (N_13064,N_5877,N_6940);
or U13065 (N_13065,N_6451,N_6281);
xnor U13066 (N_13066,N_5415,N_9544);
nor U13067 (N_13067,N_7567,N_9673);
nor U13068 (N_13068,N_5930,N_9271);
and U13069 (N_13069,N_9134,N_9695);
or U13070 (N_13070,N_5310,N_7627);
or U13071 (N_13071,N_8218,N_9165);
and U13072 (N_13072,N_6826,N_6549);
nor U13073 (N_13073,N_5750,N_6899);
xor U13074 (N_13074,N_9199,N_9159);
and U13075 (N_13075,N_5267,N_5066);
and U13076 (N_13076,N_6927,N_9701);
or U13077 (N_13077,N_9510,N_9783);
nor U13078 (N_13078,N_7766,N_9073);
or U13079 (N_13079,N_7007,N_9952);
nand U13080 (N_13080,N_5760,N_5123);
or U13081 (N_13081,N_6254,N_5062);
nand U13082 (N_13082,N_5685,N_7430);
and U13083 (N_13083,N_9335,N_6709);
and U13084 (N_13084,N_7098,N_7970);
and U13085 (N_13085,N_5344,N_5272);
nand U13086 (N_13086,N_6052,N_5340);
xor U13087 (N_13087,N_6378,N_5854);
nor U13088 (N_13088,N_9395,N_9989);
xor U13089 (N_13089,N_7010,N_9875);
or U13090 (N_13090,N_7227,N_7318);
or U13091 (N_13091,N_9849,N_8390);
nor U13092 (N_13092,N_6382,N_9423);
xor U13093 (N_13093,N_5957,N_5310);
nand U13094 (N_13094,N_6139,N_8414);
nor U13095 (N_13095,N_9750,N_7687);
and U13096 (N_13096,N_9630,N_8147);
xor U13097 (N_13097,N_6715,N_6918);
xor U13098 (N_13098,N_7636,N_7784);
and U13099 (N_13099,N_6213,N_5533);
xnor U13100 (N_13100,N_9420,N_7032);
nand U13101 (N_13101,N_5250,N_8160);
nand U13102 (N_13102,N_5919,N_5351);
or U13103 (N_13103,N_9595,N_7704);
nor U13104 (N_13104,N_7538,N_5191);
nand U13105 (N_13105,N_8475,N_8474);
or U13106 (N_13106,N_7442,N_9551);
and U13107 (N_13107,N_7141,N_5173);
nand U13108 (N_13108,N_8545,N_9870);
xor U13109 (N_13109,N_9918,N_8578);
nand U13110 (N_13110,N_5448,N_9003);
nand U13111 (N_13111,N_6214,N_5261);
xnor U13112 (N_13112,N_8741,N_7419);
and U13113 (N_13113,N_8550,N_5990);
nand U13114 (N_13114,N_6930,N_6497);
nand U13115 (N_13115,N_7753,N_6045);
xor U13116 (N_13116,N_6436,N_8087);
and U13117 (N_13117,N_5930,N_5145);
xor U13118 (N_13118,N_8515,N_7078);
nor U13119 (N_13119,N_8717,N_5713);
nor U13120 (N_13120,N_7807,N_9792);
and U13121 (N_13121,N_6575,N_5396);
nor U13122 (N_13122,N_9702,N_9934);
nand U13123 (N_13123,N_9641,N_7661);
nand U13124 (N_13124,N_5938,N_6181);
or U13125 (N_13125,N_7782,N_6064);
and U13126 (N_13126,N_9803,N_7317);
and U13127 (N_13127,N_7643,N_9150);
nand U13128 (N_13128,N_7910,N_6785);
nand U13129 (N_13129,N_6267,N_9763);
and U13130 (N_13130,N_7374,N_7207);
or U13131 (N_13131,N_7185,N_5096);
xor U13132 (N_13132,N_6334,N_8971);
and U13133 (N_13133,N_9706,N_7571);
or U13134 (N_13134,N_9386,N_8685);
and U13135 (N_13135,N_7658,N_9857);
nor U13136 (N_13136,N_5336,N_9006);
xor U13137 (N_13137,N_9298,N_8843);
and U13138 (N_13138,N_6667,N_6181);
nor U13139 (N_13139,N_9170,N_7118);
nor U13140 (N_13140,N_6930,N_8986);
and U13141 (N_13141,N_6929,N_7614);
xor U13142 (N_13142,N_5084,N_5419);
nor U13143 (N_13143,N_9889,N_7349);
xor U13144 (N_13144,N_5418,N_7253);
nor U13145 (N_13145,N_5339,N_8699);
xnor U13146 (N_13146,N_7080,N_8567);
and U13147 (N_13147,N_8973,N_9579);
nand U13148 (N_13148,N_5282,N_9266);
or U13149 (N_13149,N_7020,N_9881);
nor U13150 (N_13150,N_8283,N_9658);
or U13151 (N_13151,N_6549,N_9982);
and U13152 (N_13152,N_9600,N_7020);
xor U13153 (N_13153,N_6888,N_8222);
nor U13154 (N_13154,N_9785,N_5252);
or U13155 (N_13155,N_7047,N_7626);
nor U13156 (N_13156,N_9919,N_6328);
or U13157 (N_13157,N_5861,N_9456);
nor U13158 (N_13158,N_7210,N_7264);
nand U13159 (N_13159,N_7230,N_7200);
or U13160 (N_13160,N_6526,N_7944);
and U13161 (N_13161,N_7663,N_5656);
or U13162 (N_13162,N_9061,N_7216);
xor U13163 (N_13163,N_7176,N_9738);
and U13164 (N_13164,N_9882,N_7309);
and U13165 (N_13165,N_7217,N_7733);
or U13166 (N_13166,N_5670,N_9438);
xnor U13167 (N_13167,N_9222,N_8229);
or U13168 (N_13168,N_5612,N_8588);
xnor U13169 (N_13169,N_5043,N_9522);
or U13170 (N_13170,N_9871,N_8718);
and U13171 (N_13171,N_9825,N_7846);
xor U13172 (N_13172,N_7721,N_6349);
or U13173 (N_13173,N_9998,N_7629);
nand U13174 (N_13174,N_7063,N_7227);
nand U13175 (N_13175,N_8208,N_7706);
or U13176 (N_13176,N_5900,N_5192);
nor U13177 (N_13177,N_5554,N_5348);
and U13178 (N_13178,N_9820,N_8731);
nand U13179 (N_13179,N_8067,N_8258);
and U13180 (N_13180,N_6274,N_7298);
nor U13181 (N_13181,N_6926,N_6627);
nand U13182 (N_13182,N_8796,N_9042);
or U13183 (N_13183,N_8588,N_7455);
or U13184 (N_13184,N_6861,N_9321);
or U13185 (N_13185,N_7020,N_7880);
nand U13186 (N_13186,N_8776,N_8502);
or U13187 (N_13187,N_5979,N_7042);
nor U13188 (N_13188,N_9025,N_6243);
xor U13189 (N_13189,N_8253,N_7664);
or U13190 (N_13190,N_6426,N_6792);
xnor U13191 (N_13191,N_6376,N_8984);
nor U13192 (N_13192,N_8018,N_5998);
and U13193 (N_13193,N_5984,N_8015);
or U13194 (N_13194,N_8433,N_7695);
or U13195 (N_13195,N_5606,N_8690);
nand U13196 (N_13196,N_6758,N_9392);
and U13197 (N_13197,N_9325,N_8302);
nand U13198 (N_13198,N_8761,N_8360);
nand U13199 (N_13199,N_8038,N_7172);
or U13200 (N_13200,N_5629,N_6876);
xor U13201 (N_13201,N_5490,N_5856);
nor U13202 (N_13202,N_8931,N_6274);
or U13203 (N_13203,N_9325,N_7599);
xnor U13204 (N_13204,N_9975,N_6790);
and U13205 (N_13205,N_8674,N_6264);
or U13206 (N_13206,N_9367,N_8230);
or U13207 (N_13207,N_8885,N_5960);
nand U13208 (N_13208,N_6260,N_7036);
or U13209 (N_13209,N_6735,N_8056);
nor U13210 (N_13210,N_8226,N_9028);
nor U13211 (N_13211,N_7005,N_5777);
nand U13212 (N_13212,N_6934,N_7856);
nand U13213 (N_13213,N_9493,N_7031);
or U13214 (N_13214,N_5973,N_7829);
nand U13215 (N_13215,N_7214,N_9628);
nand U13216 (N_13216,N_8289,N_5248);
and U13217 (N_13217,N_5910,N_5594);
nand U13218 (N_13218,N_9469,N_6854);
and U13219 (N_13219,N_5611,N_9803);
and U13220 (N_13220,N_6258,N_9304);
nor U13221 (N_13221,N_8996,N_9460);
nand U13222 (N_13222,N_6046,N_9153);
nor U13223 (N_13223,N_9704,N_7599);
nor U13224 (N_13224,N_9927,N_6142);
or U13225 (N_13225,N_7676,N_6590);
or U13226 (N_13226,N_7444,N_6064);
xnor U13227 (N_13227,N_9272,N_5811);
xnor U13228 (N_13228,N_9859,N_7568);
or U13229 (N_13229,N_7216,N_7313);
and U13230 (N_13230,N_5887,N_6806);
nand U13231 (N_13231,N_7522,N_8137);
xnor U13232 (N_13232,N_5637,N_8734);
xor U13233 (N_13233,N_7690,N_8774);
xnor U13234 (N_13234,N_8187,N_9397);
or U13235 (N_13235,N_9751,N_7121);
nand U13236 (N_13236,N_5683,N_8360);
or U13237 (N_13237,N_8237,N_5018);
or U13238 (N_13238,N_9438,N_9543);
xor U13239 (N_13239,N_8488,N_6666);
and U13240 (N_13240,N_7289,N_9422);
nand U13241 (N_13241,N_8230,N_7066);
nor U13242 (N_13242,N_6576,N_6019);
and U13243 (N_13243,N_8378,N_7712);
and U13244 (N_13244,N_6826,N_6752);
nor U13245 (N_13245,N_9143,N_6284);
or U13246 (N_13246,N_5353,N_8177);
or U13247 (N_13247,N_6464,N_5643);
or U13248 (N_13248,N_9179,N_9187);
nor U13249 (N_13249,N_5621,N_9429);
nand U13250 (N_13250,N_6575,N_7817);
nor U13251 (N_13251,N_6249,N_5498);
nand U13252 (N_13252,N_7082,N_6180);
nor U13253 (N_13253,N_6268,N_8543);
nor U13254 (N_13254,N_6974,N_8611);
xnor U13255 (N_13255,N_6728,N_9400);
nand U13256 (N_13256,N_6416,N_7467);
xor U13257 (N_13257,N_5636,N_6200);
nand U13258 (N_13258,N_7973,N_6142);
xor U13259 (N_13259,N_7672,N_7528);
and U13260 (N_13260,N_6298,N_9570);
and U13261 (N_13261,N_8616,N_6490);
nand U13262 (N_13262,N_8686,N_9240);
xnor U13263 (N_13263,N_5365,N_8992);
and U13264 (N_13264,N_6495,N_7406);
nand U13265 (N_13265,N_9111,N_5185);
or U13266 (N_13266,N_5039,N_5168);
xnor U13267 (N_13267,N_5854,N_9231);
nor U13268 (N_13268,N_5103,N_7706);
or U13269 (N_13269,N_6111,N_6345);
nor U13270 (N_13270,N_6542,N_5510);
xnor U13271 (N_13271,N_6706,N_7531);
xnor U13272 (N_13272,N_5623,N_8338);
or U13273 (N_13273,N_5997,N_8588);
nor U13274 (N_13274,N_7051,N_7596);
or U13275 (N_13275,N_5844,N_7861);
nand U13276 (N_13276,N_6076,N_9978);
or U13277 (N_13277,N_9199,N_9347);
or U13278 (N_13278,N_8906,N_5954);
nand U13279 (N_13279,N_8563,N_5107);
nor U13280 (N_13280,N_9029,N_9788);
xor U13281 (N_13281,N_8251,N_6073);
nand U13282 (N_13282,N_8418,N_5727);
or U13283 (N_13283,N_7090,N_5377);
nor U13284 (N_13284,N_7210,N_6205);
xnor U13285 (N_13285,N_6726,N_8870);
and U13286 (N_13286,N_5799,N_8009);
and U13287 (N_13287,N_6702,N_6925);
and U13288 (N_13288,N_5386,N_6321);
or U13289 (N_13289,N_9591,N_6156);
nor U13290 (N_13290,N_6643,N_5553);
nor U13291 (N_13291,N_6813,N_5293);
nor U13292 (N_13292,N_5512,N_6726);
and U13293 (N_13293,N_6273,N_5445);
nand U13294 (N_13294,N_5309,N_6459);
xnor U13295 (N_13295,N_5063,N_5653);
nor U13296 (N_13296,N_7609,N_7662);
or U13297 (N_13297,N_6043,N_7976);
and U13298 (N_13298,N_7499,N_5378);
and U13299 (N_13299,N_5992,N_9452);
nand U13300 (N_13300,N_7013,N_5067);
xor U13301 (N_13301,N_8154,N_7942);
nor U13302 (N_13302,N_7701,N_8371);
nor U13303 (N_13303,N_7472,N_9545);
nand U13304 (N_13304,N_8384,N_5283);
nand U13305 (N_13305,N_7326,N_5456);
or U13306 (N_13306,N_7437,N_6026);
nand U13307 (N_13307,N_9866,N_7112);
or U13308 (N_13308,N_8186,N_6782);
nand U13309 (N_13309,N_8795,N_7341);
or U13310 (N_13310,N_9298,N_9870);
and U13311 (N_13311,N_8803,N_7132);
and U13312 (N_13312,N_9893,N_7529);
nand U13313 (N_13313,N_8852,N_7596);
and U13314 (N_13314,N_9791,N_9377);
and U13315 (N_13315,N_7365,N_7008);
and U13316 (N_13316,N_8199,N_5086);
and U13317 (N_13317,N_6883,N_8489);
nor U13318 (N_13318,N_6228,N_5493);
and U13319 (N_13319,N_5206,N_9299);
nor U13320 (N_13320,N_7703,N_6357);
nor U13321 (N_13321,N_7546,N_6813);
or U13322 (N_13322,N_9844,N_9313);
nand U13323 (N_13323,N_8832,N_7866);
nor U13324 (N_13324,N_8105,N_9491);
xor U13325 (N_13325,N_6231,N_8463);
and U13326 (N_13326,N_9150,N_5760);
and U13327 (N_13327,N_8862,N_7924);
nor U13328 (N_13328,N_9299,N_8877);
or U13329 (N_13329,N_7804,N_8916);
nand U13330 (N_13330,N_6053,N_8994);
nand U13331 (N_13331,N_8931,N_6347);
and U13332 (N_13332,N_7251,N_8128);
nand U13333 (N_13333,N_5279,N_8223);
or U13334 (N_13334,N_9156,N_5143);
or U13335 (N_13335,N_9466,N_7556);
xor U13336 (N_13336,N_8170,N_6181);
xor U13337 (N_13337,N_5904,N_6063);
nand U13338 (N_13338,N_8185,N_8788);
nand U13339 (N_13339,N_6392,N_9373);
or U13340 (N_13340,N_8811,N_9902);
or U13341 (N_13341,N_6254,N_6472);
or U13342 (N_13342,N_7605,N_5909);
or U13343 (N_13343,N_9220,N_5769);
or U13344 (N_13344,N_8824,N_7991);
nand U13345 (N_13345,N_7598,N_5913);
and U13346 (N_13346,N_5383,N_5587);
or U13347 (N_13347,N_5337,N_6974);
and U13348 (N_13348,N_5545,N_8485);
nor U13349 (N_13349,N_6522,N_6031);
and U13350 (N_13350,N_5105,N_5926);
nor U13351 (N_13351,N_5398,N_7720);
nand U13352 (N_13352,N_6779,N_9746);
and U13353 (N_13353,N_8796,N_8300);
or U13354 (N_13354,N_5404,N_9157);
nor U13355 (N_13355,N_9975,N_6548);
and U13356 (N_13356,N_7436,N_7080);
or U13357 (N_13357,N_9474,N_7655);
xnor U13358 (N_13358,N_8580,N_7012);
or U13359 (N_13359,N_6766,N_8284);
xnor U13360 (N_13360,N_6443,N_5340);
nand U13361 (N_13361,N_9366,N_9050);
nor U13362 (N_13362,N_7526,N_9833);
nand U13363 (N_13363,N_8605,N_7028);
nand U13364 (N_13364,N_8627,N_9571);
nand U13365 (N_13365,N_8776,N_7731);
or U13366 (N_13366,N_9056,N_5384);
and U13367 (N_13367,N_5180,N_6032);
and U13368 (N_13368,N_8980,N_7218);
xnor U13369 (N_13369,N_9335,N_5400);
xnor U13370 (N_13370,N_7249,N_5837);
nand U13371 (N_13371,N_8457,N_7810);
nor U13372 (N_13372,N_7317,N_7985);
xnor U13373 (N_13373,N_6713,N_6689);
xor U13374 (N_13374,N_6328,N_7964);
or U13375 (N_13375,N_8590,N_8872);
nand U13376 (N_13376,N_5256,N_5245);
xor U13377 (N_13377,N_8970,N_5995);
or U13378 (N_13378,N_6022,N_9803);
or U13379 (N_13379,N_9130,N_7395);
or U13380 (N_13380,N_6160,N_9546);
nor U13381 (N_13381,N_8005,N_5765);
nor U13382 (N_13382,N_5979,N_5684);
nor U13383 (N_13383,N_9592,N_7428);
and U13384 (N_13384,N_9743,N_7271);
nor U13385 (N_13385,N_9480,N_8892);
and U13386 (N_13386,N_8446,N_9227);
nor U13387 (N_13387,N_7540,N_6095);
or U13388 (N_13388,N_5064,N_7293);
nor U13389 (N_13389,N_7113,N_8140);
xnor U13390 (N_13390,N_8686,N_6199);
nand U13391 (N_13391,N_7240,N_6004);
nor U13392 (N_13392,N_9369,N_9598);
or U13393 (N_13393,N_6565,N_6236);
and U13394 (N_13394,N_8209,N_9663);
and U13395 (N_13395,N_9231,N_6176);
xor U13396 (N_13396,N_6058,N_9428);
xor U13397 (N_13397,N_9447,N_8949);
nand U13398 (N_13398,N_7915,N_7757);
xor U13399 (N_13399,N_7194,N_9219);
and U13400 (N_13400,N_8901,N_8977);
nor U13401 (N_13401,N_8336,N_8598);
xnor U13402 (N_13402,N_6738,N_9588);
and U13403 (N_13403,N_8983,N_9172);
or U13404 (N_13404,N_5186,N_9433);
xor U13405 (N_13405,N_5453,N_8433);
nor U13406 (N_13406,N_6413,N_6643);
nor U13407 (N_13407,N_7548,N_9450);
and U13408 (N_13408,N_8943,N_7311);
and U13409 (N_13409,N_7049,N_9020);
or U13410 (N_13410,N_8590,N_7449);
nor U13411 (N_13411,N_9224,N_8022);
xor U13412 (N_13412,N_6975,N_7173);
nor U13413 (N_13413,N_6313,N_5024);
and U13414 (N_13414,N_8895,N_9183);
nor U13415 (N_13415,N_8437,N_7182);
nand U13416 (N_13416,N_8267,N_5598);
nand U13417 (N_13417,N_5786,N_7592);
and U13418 (N_13418,N_5921,N_9167);
nor U13419 (N_13419,N_7478,N_9593);
xnor U13420 (N_13420,N_9359,N_7559);
or U13421 (N_13421,N_8039,N_6057);
nor U13422 (N_13422,N_7931,N_6987);
nand U13423 (N_13423,N_7352,N_6080);
nand U13424 (N_13424,N_8306,N_9349);
nand U13425 (N_13425,N_6526,N_5315);
and U13426 (N_13426,N_9822,N_8189);
xnor U13427 (N_13427,N_7862,N_9548);
nand U13428 (N_13428,N_6089,N_9966);
and U13429 (N_13429,N_8256,N_7668);
nor U13430 (N_13430,N_6594,N_7381);
and U13431 (N_13431,N_6789,N_9917);
or U13432 (N_13432,N_6938,N_6771);
nor U13433 (N_13433,N_8026,N_5192);
nand U13434 (N_13434,N_6862,N_8228);
or U13435 (N_13435,N_6220,N_5302);
xnor U13436 (N_13436,N_5465,N_5607);
or U13437 (N_13437,N_5522,N_5465);
xor U13438 (N_13438,N_6903,N_8827);
nor U13439 (N_13439,N_6673,N_5407);
nand U13440 (N_13440,N_7960,N_9308);
or U13441 (N_13441,N_8755,N_7190);
nor U13442 (N_13442,N_7271,N_8536);
xnor U13443 (N_13443,N_7462,N_6119);
and U13444 (N_13444,N_7902,N_5681);
nand U13445 (N_13445,N_8575,N_6873);
or U13446 (N_13446,N_8488,N_7914);
nand U13447 (N_13447,N_6027,N_9340);
and U13448 (N_13448,N_5530,N_6540);
and U13449 (N_13449,N_8242,N_7264);
and U13450 (N_13450,N_6133,N_8619);
nand U13451 (N_13451,N_8501,N_9889);
xor U13452 (N_13452,N_9607,N_7080);
nand U13453 (N_13453,N_8997,N_6232);
and U13454 (N_13454,N_7180,N_6408);
xnor U13455 (N_13455,N_7739,N_9441);
and U13456 (N_13456,N_5211,N_5652);
nand U13457 (N_13457,N_5631,N_5092);
xor U13458 (N_13458,N_8984,N_8010);
xnor U13459 (N_13459,N_7350,N_7464);
and U13460 (N_13460,N_8393,N_7449);
xnor U13461 (N_13461,N_7932,N_7128);
and U13462 (N_13462,N_8463,N_7642);
or U13463 (N_13463,N_8675,N_9779);
or U13464 (N_13464,N_8140,N_8389);
or U13465 (N_13465,N_6382,N_6129);
and U13466 (N_13466,N_6161,N_8976);
nand U13467 (N_13467,N_9989,N_5614);
nand U13468 (N_13468,N_7863,N_9525);
nand U13469 (N_13469,N_5548,N_6270);
nor U13470 (N_13470,N_6796,N_9001);
or U13471 (N_13471,N_8654,N_5136);
and U13472 (N_13472,N_9075,N_6404);
nor U13473 (N_13473,N_6999,N_9287);
nand U13474 (N_13474,N_6564,N_7579);
nor U13475 (N_13475,N_5200,N_6722);
and U13476 (N_13476,N_9726,N_7776);
nand U13477 (N_13477,N_8832,N_5092);
or U13478 (N_13478,N_8139,N_9556);
xor U13479 (N_13479,N_6780,N_9898);
or U13480 (N_13480,N_8243,N_8703);
and U13481 (N_13481,N_7646,N_8942);
nor U13482 (N_13482,N_8918,N_8944);
nand U13483 (N_13483,N_7248,N_9770);
nor U13484 (N_13484,N_8458,N_6233);
nand U13485 (N_13485,N_5175,N_8868);
nor U13486 (N_13486,N_7195,N_6432);
or U13487 (N_13487,N_5927,N_9001);
and U13488 (N_13488,N_7639,N_8134);
nand U13489 (N_13489,N_7187,N_7343);
nor U13490 (N_13490,N_7663,N_9258);
or U13491 (N_13491,N_6490,N_8318);
nor U13492 (N_13492,N_5424,N_9688);
xnor U13493 (N_13493,N_5781,N_9567);
nand U13494 (N_13494,N_8810,N_7473);
and U13495 (N_13495,N_7823,N_8533);
xnor U13496 (N_13496,N_9254,N_6153);
and U13497 (N_13497,N_7889,N_6180);
nor U13498 (N_13498,N_8148,N_7783);
nor U13499 (N_13499,N_6020,N_7584);
nor U13500 (N_13500,N_6499,N_9282);
and U13501 (N_13501,N_6680,N_9700);
or U13502 (N_13502,N_5131,N_7822);
and U13503 (N_13503,N_5766,N_5229);
or U13504 (N_13504,N_8767,N_5002);
xnor U13505 (N_13505,N_6561,N_6269);
and U13506 (N_13506,N_5245,N_7822);
nand U13507 (N_13507,N_6610,N_6303);
xnor U13508 (N_13508,N_8068,N_7104);
and U13509 (N_13509,N_7343,N_9383);
xnor U13510 (N_13510,N_7280,N_9656);
xor U13511 (N_13511,N_7075,N_5234);
and U13512 (N_13512,N_5352,N_5278);
or U13513 (N_13513,N_7702,N_9652);
xnor U13514 (N_13514,N_6834,N_6805);
nor U13515 (N_13515,N_9813,N_9768);
nor U13516 (N_13516,N_7260,N_7342);
xor U13517 (N_13517,N_9660,N_9980);
and U13518 (N_13518,N_9567,N_9157);
or U13519 (N_13519,N_9710,N_7949);
and U13520 (N_13520,N_7262,N_5882);
nand U13521 (N_13521,N_7855,N_9070);
or U13522 (N_13522,N_8588,N_8599);
nor U13523 (N_13523,N_9404,N_9313);
and U13524 (N_13524,N_7211,N_9032);
xnor U13525 (N_13525,N_8106,N_7931);
or U13526 (N_13526,N_8134,N_6698);
nand U13527 (N_13527,N_7185,N_5253);
or U13528 (N_13528,N_5426,N_7138);
nand U13529 (N_13529,N_6970,N_9168);
nor U13530 (N_13530,N_8475,N_7458);
nand U13531 (N_13531,N_5958,N_7336);
nand U13532 (N_13532,N_8342,N_9236);
and U13533 (N_13533,N_5988,N_7524);
nor U13534 (N_13534,N_8191,N_9013);
nand U13535 (N_13535,N_8437,N_7990);
nor U13536 (N_13536,N_8723,N_9294);
and U13537 (N_13537,N_7894,N_5971);
nand U13538 (N_13538,N_5106,N_6659);
nand U13539 (N_13539,N_9680,N_6020);
nand U13540 (N_13540,N_5410,N_7946);
or U13541 (N_13541,N_6062,N_5872);
xnor U13542 (N_13542,N_5678,N_8522);
and U13543 (N_13543,N_7002,N_7783);
or U13544 (N_13544,N_7224,N_8204);
xor U13545 (N_13545,N_8568,N_9373);
or U13546 (N_13546,N_7124,N_5838);
or U13547 (N_13547,N_6243,N_8764);
nor U13548 (N_13548,N_5293,N_7374);
nor U13549 (N_13549,N_8114,N_8981);
nand U13550 (N_13550,N_6961,N_6512);
nor U13551 (N_13551,N_8216,N_9797);
nor U13552 (N_13552,N_8218,N_8600);
xor U13553 (N_13553,N_5689,N_9531);
nand U13554 (N_13554,N_6879,N_5911);
or U13555 (N_13555,N_7019,N_5246);
and U13556 (N_13556,N_7263,N_8888);
xnor U13557 (N_13557,N_8219,N_8163);
and U13558 (N_13558,N_9713,N_8374);
and U13559 (N_13559,N_9814,N_9387);
or U13560 (N_13560,N_8232,N_9701);
nand U13561 (N_13561,N_5868,N_8977);
or U13562 (N_13562,N_9071,N_7469);
nor U13563 (N_13563,N_8553,N_8617);
nand U13564 (N_13564,N_6838,N_8204);
nand U13565 (N_13565,N_7365,N_6062);
or U13566 (N_13566,N_8260,N_6015);
nand U13567 (N_13567,N_9932,N_5877);
and U13568 (N_13568,N_6807,N_6534);
nor U13569 (N_13569,N_6169,N_8180);
nand U13570 (N_13570,N_5859,N_5594);
and U13571 (N_13571,N_8446,N_6759);
nand U13572 (N_13572,N_6932,N_7480);
and U13573 (N_13573,N_5540,N_8732);
nand U13574 (N_13574,N_6015,N_6989);
or U13575 (N_13575,N_6650,N_7832);
and U13576 (N_13576,N_7650,N_9859);
or U13577 (N_13577,N_7944,N_9127);
or U13578 (N_13578,N_8246,N_6403);
and U13579 (N_13579,N_5885,N_9842);
or U13580 (N_13580,N_6398,N_6219);
or U13581 (N_13581,N_8102,N_6406);
xor U13582 (N_13582,N_6930,N_8809);
xnor U13583 (N_13583,N_6985,N_6473);
or U13584 (N_13584,N_9661,N_9769);
nor U13585 (N_13585,N_6854,N_8510);
xor U13586 (N_13586,N_8173,N_6472);
nand U13587 (N_13587,N_7099,N_6847);
and U13588 (N_13588,N_7478,N_8162);
and U13589 (N_13589,N_9803,N_6961);
and U13590 (N_13590,N_7022,N_7241);
nand U13591 (N_13591,N_5356,N_7673);
nor U13592 (N_13592,N_8811,N_6537);
or U13593 (N_13593,N_5418,N_8942);
and U13594 (N_13594,N_6883,N_5483);
nand U13595 (N_13595,N_9638,N_5860);
and U13596 (N_13596,N_9431,N_8281);
nor U13597 (N_13597,N_7756,N_5037);
nor U13598 (N_13598,N_9799,N_6359);
or U13599 (N_13599,N_8142,N_6095);
nor U13600 (N_13600,N_7829,N_8133);
nor U13601 (N_13601,N_9104,N_6316);
or U13602 (N_13602,N_9759,N_9039);
and U13603 (N_13603,N_9285,N_5280);
xnor U13604 (N_13604,N_5392,N_9499);
or U13605 (N_13605,N_7116,N_8032);
and U13606 (N_13606,N_5307,N_6816);
xor U13607 (N_13607,N_7341,N_5928);
and U13608 (N_13608,N_8411,N_9621);
or U13609 (N_13609,N_5885,N_7143);
nand U13610 (N_13610,N_8768,N_9363);
xnor U13611 (N_13611,N_6763,N_6776);
xnor U13612 (N_13612,N_7923,N_7657);
xnor U13613 (N_13613,N_9001,N_7028);
and U13614 (N_13614,N_7105,N_8158);
nor U13615 (N_13615,N_5578,N_6379);
or U13616 (N_13616,N_8095,N_6579);
and U13617 (N_13617,N_5698,N_8411);
nor U13618 (N_13618,N_5288,N_8054);
xnor U13619 (N_13619,N_7913,N_7223);
and U13620 (N_13620,N_9194,N_7498);
xnor U13621 (N_13621,N_9848,N_8380);
or U13622 (N_13622,N_8930,N_8737);
nor U13623 (N_13623,N_9804,N_6557);
nand U13624 (N_13624,N_6342,N_8905);
and U13625 (N_13625,N_8994,N_8960);
or U13626 (N_13626,N_6507,N_9428);
nand U13627 (N_13627,N_5866,N_7704);
and U13628 (N_13628,N_7125,N_6311);
or U13629 (N_13629,N_5872,N_8998);
or U13630 (N_13630,N_9087,N_6640);
or U13631 (N_13631,N_8852,N_5920);
nor U13632 (N_13632,N_5871,N_8809);
or U13633 (N_13633,N_9039,N_9449);
and U13634 (N_13634,N_5893,N_7730);
xnor U13635 (N_13635,N_5068,N_5931);
or U13636 (N_13636,N_6791,N_8337);
or U13637 (N_13637,N_6908,N_8454);
xor U13638 (N_13638,N_8391,N_7704);
xnor U13639 (N_13639,N_7282,N_8197);
nand U13640 (N_13640,N_5456,N_8636);
nand U13641 (N_13641,N_9700,N_5243);
or U13642 (N_13642,N_8172,N_8908);
and U13643 (N_13643,N_9200,N_9783);
nand U13644 (N_13644,N_6544,N_6849);
nand U13645 (N_13645,N_7468,N_9611);
and U13646 (N_13646,N_5281,N_9598);
and U13647 (N_13647,N_8182,N_6642);
xnor U13648 (N_13648,N_7065,N_8638);
or U13649 (N_13649,N_5951,N_7944);
nor U13650 (N_13650,N_7179,N_7727);
nand U13651 (N_13651,N_8437,N_6555);
nand U13652 (N_13652,N_5993,N_8384);
and U13653 (N_13653,N_5800,N_8518);
xor U13654 (N_13654,N_9232,N_7956);
nor U13655 (N_13655,N_9402,N_5764);
nand U13656 (N_13656,N_5786,N_5959);
and U13657 (N_13657,N_5683,N_5851);
xor U13658 (N_13658,N_8217,N_9213);
nor U13659 (N_13659,N_9577,N_5136);
nor U13660 (N_13660,N_7493,N_8056);
xnor U13661 (N_13661,N_7342,N_8273);
nand U13662 (N_13662,N_7305,N_7459);
nor U13663 (N_13663,N_7216,N_9376);
or U13664 (N_13664,N_9294,N_5235);
and U13665 (N_13665,N_5482,N_6631);
nor U13666 (N_13666,N_7667,N_8158);
and U13667 (N_13667,N_9940,N_8242);
and U13668 (N_13668,N_8542,N_8263);
xor U13669 (N_13669,N_5111,N_5914);
xor U13670 (N_13670,N_8053,N_6829);
nand U13671 (N_13671,N_5341,N_5096);
xnor U13672 (N_13672,N_8874,N_9313);
xor U13673 (N_13673,N_8320,N_7941);
nor U13674 (N_13674,N_6156,N_7371);
and U13675 (N_13675,N_8420,N_6241);
nor U13676 (N_13676,N_5999,N_5670);
xor U13677 (N_13677,N_8104,N_7568);
or U13678 (N_13678,N_6570,N_5579);
or U13679 (N_13679,N_7141,N_8542);
or U13680 (N_13680,N_8179,N_6354);
nand U13681 (N_13681,N_9297,N_9458);
or U13682 (N_13682,N_6184,N_8191);
nand U13683 (N_13683,N_5939,N_7726);
and U13684 (N_13684,N_6118,N_6908);
xor U13685 (N_13685,N_7765,N_6856);
or U13686 (N_13686,N_5775,N_6474);
or U13687 (N_13687,N_9027,N_7890);
xnor U13688 (N_13688,N_8927,N_5822);
nor U13689 (N_13689,N_9066,N_8083);
nor U13690 (N_13690,N_9531,N_5446);
or U13691 (N_13691,N_5561,N_9972);
nor U13692 (N_13692,N_8590,N_8920);
nand U13693 (N_13693,N_6634,N_6774);
or U13694 (N_13694,N_6323,N_6865);
nor U13695 (N_13695,N_5349,N_8046);
xnor U13696 (N_13696,N_8006,N_6356);
nor U13697 (N_13697,N_7355,N_7994);
nor U13698 (N_13698,N_6868,N_8661);
and U13699 (N_13699,N_8370,N_9458);
nand U13700 (N_13700,N_6942,N_8516);
nor U13701 (N_13701,N_7371,N_6402);
nor U13702 (N_13702,N_7022,N_7361);
xnor U13703 (N_13703,N_6034,N_8744);
nor U13704 (N_13704,N_7077,N_8249);
xor U13705 (N_13705,N_6205,N_6477);
and U13706 (N_13706,N_7164,N_8272);
and U13707 (N_13707,N_9263,N_8437);
nand U13708 (N_13708,N_7683,N_9113);
nand U13709 (N_13709,N_5636,N_5149);
or U13710 (N_13710,N_5663,N_6871);
xor U13711 (N_13711,N_6452,N_8766);
xor U13712 (N_13712,N_9486,N_9169);
xor U13713 (N_13713,N_5305,N_6517);
and U13714 (N_13714,N_6931,N_7303);
xor U13715 (N_13715,N_9613,N_9295);
or U13716 (N_13716,N_5084,N_6996);
or U13717 (N_13717,N_6938,N_9467);
xor U13718 (N_13718,N_6774,N_7105);
and U13719 (N_13719,N_6239,N_7040);
nor U13720 (N_13720,N_5342,N_8881);
nand U13721 (N_13721,N_9110,N_7615);
xor U13722 (N_13722,N_9708,N_9373);
and U13723 (N_13723,N_6774,N_7660);
nor U13724 (N_13724,N_5257,N_6598);
nand U13725 (N_13725,N_9127,N_7778);
nand U13726 (N_13726,N_8169,N_7540);
and U13727 (N_13727,N_6459,N_5592);
nand U13728 (N_13728,N_9048,N_7726);
nor U13729 (N_13729,N_7639,N_6839);
nor U13730 (N_13730,N_9695,N_9502);
or U13731 (N_13731,N_7802,N_8384);
and U13732 (N_13732,N_8017,N_7799);
and U13733 (N_13733,N_9576,N_6921);
nand U13734 (N_13734,N_5184,N_6367);
xnor U13735 (N_13735,N_6099,N_5477);
xnor U13736 (N_13736,N_5220,N_6744);
xnor U13737 (N_13737,N_9277,N_7905);
nand U13738 (N_13738,N_8813,N_5830);
nand U13739 (N_13739,N_5822,N_6583);
nor U13740 (N_13740,N_9239,N_7183);
or U13741 (N_13741,N_5147,N_5694);
xnor U13742 (N_13742,N_7077,N_6713);
xor U13743 (N_13743,N_5334,N_8645);
and U13744 (N_13744,N_9832,N_9263);
xor U13745 (N_13745,N_7319,N_8587);
nand U13746 (N_13746,N_6686,N_6315);
nand U13747 (N_13747,N_5260,N_8931);
and U13748 (N_13748,N_7476,N_6771);
or U13749 (N_13749,N_8013,N_7928);
xnor U13750 (N_13750,N_6185,N_5661);
xor U13751 (N_13751,N_6661,N_6015);
nand U13752 (N_13752,N_7229,N_7894);
or U13753 (N_13753,N_7054,N_8033);
xnor U13754 (N_13754,N_8048,N_8487);
xor U13755 (N_13755,N_9694,N_6369);
and U13756 (N_13756,N_8873,N_7781);
xnor U13757 (N_13757,N_8441,N_7836);
and U13758 (N_13758,N_8306,N_5644);
and U13759 (N_13759,N_8851,N_7048);
or U13760 (N_13760,N_8540,N_7062);
nand U13761 (N_13761,N_9648,N_6093);
xnor U13762 (N_13762,N_8988,N_8252);
nor U13763 (N_13763,N_8530,N_9058);
nor U13764 (N_13764,N_5433,N_8368);
nor U13765 (N_13765,N_8572,N_6332);
nor U13766 (N_13766,N_7308,N_6856);
nor U13767 (N_13767,N_5578,N_6493);
and U13768 (N_13768,N_9898,N_6891);
nand U13769 (N_13769,N_8093,N_5571);
or U13770 (N_13770,N_9274,N_9820);
and U13771 (N_13771,N_8357,N_8068);
nor U13772 (N_13772,N_9618,N_8697);
nor U13773 (N_13773,N_5318,N_6547);
nor U13774 (N_13774,N_6516,N_6355);
or U13775 (N_13775,N_8656,N_7528);
or U13776 (N_13776,N_8498,N_7227);
nor U13777 (N_13777,N_6499,N_6773);
and U13778 (N_13778,N_6022,N_9278);
and U13779 (N_13779,N_5686,N_5079);
and U13780 (N_13780,N_6137,N_6455);
nor U13781 (N_13781,N_5797,N_8227);
nor U13782 (N_13782,N_8950,N_9865);
and U13783 (N_13783,N_7433,N_5270);
or U13784 (N_13784,N_6465,N_6499);
nand U13785 (N_13785,N_7053,N_7149);
and U13786 (N_13786,N_6929,N_5488);
or U13787 (N_13787,N_8050,N_9937);
or U13788 (N_13788,N_6598,N_5565);
xor U13789 (N_13789,N_5580,N_6386);
nor U13790 (N_13790,N_5299,N_8026);
and U13791 (N_13791,N_6512,N_5106);
nand U13792 (N_13792,N_6339,N_8233);
nand U13793 (N_13793,N_9247,N_8749);
and U13794 (N_13794,N_7361,N_7954);
or U13795 (N_13795,N_9823,N_8780);
and U13796 (N_13796,N_6288,N_9129);
or U13797 (N_13797,N_7389,N_8515);
nor U13798 (N_13798,N_5020,N_9988);
and U13799 (N_13799,N_6140,N_8396);
xor U13800 (N_13800,N_7796,N_6672);
and U13801 (N_13801,N_9899,N_5480);
and U13802 (N_13802,N_9082,N_8788);
nand U13803 (N_13803,N_5283,N_5396);
or U13804 (N_13804,N_8302,N_5992);
or U13805 (N_13805,N_7761,N_7489);
and U13806 (N_13806,N_8881,N_7431);
or U13807 (N_13807,N_6192,N_9178);
and U13808 (N_13808,N_8794,N_6639);
and U13809 (N_13809,N_8278,N_7303);
or U13810 (N_13810,N_5665,N_6523);
or U13811 (N_13811,N_8063,N_8227);
nand U13812 (N_13812,N_8563,N_7773);
nand U13813 (N_13813,N_7319,N_5657);
or U13814 (N_13814,N_6325,N_7598);
or U13815 (N_13815,N_9875,N_7604);
nand U13816 (N_13816,N_5726,N_8406);
and U13817 (N_13817,N_9760,N_6954);
xor U13818 (N_13818,N_6251,N_6574);
nor U13819 (N_13819,N_6627,N_7474);
nand U13820 (N_13820,N_8802,N_7492);
nor U13821 (N_13821,N_7691,N_6944);
nor U13822 (N_13822,N_5393,N_8333);
nand U13823 (N_13823,N_9039,N_5094);
xnor U13824 (N_13824,N_9386,N_8445);
or U13825 (N_13825,N_8562,N_6841);
xor U13826 (N_13826,N_8059,N_8393);
nand U13827 (N_13827,N_5921,N_7150);
xor U13828 (N_13828,N_8503,N_8081);
or U13829 (N_13829,N_8336,N_7751);
and U13830 (N_13830,N_6177,N_7802);
and U13831 (N_13831,N_9275,N_7490);
nand U13832 (N_13832,N_5664,N_6626);
nor U13833 (N_13833,N_9984,N_8614);
xor U13834 (N_13834,N_7783,N_6461);
xor U13835 (N_13835,N_8882,N_9432);
xnor U13836 (N_13836,N_8353,N_6959);
nand U13837 (N_13837,N_5964,N_7203);
or U13838 (N_13838,N_6673,N_8123);
and U13839 (N_13839,N_7597,N_6249);
xnor U13840 (N_13840,N_6693,N_6280);
xnor U13841 (N_13841,N_9006,N_6222);
or U13842 (N_13842,N_5030,N_8321);
xnor U13843 (N_13843,N_8560,N_6056);
and U13844 (N_13844,N_9473,N_6739);
and U13845 (N_13845,N_9575,N_8894);
nand U13846 (N_13846,N_9724,N_5409);
nand U13847 (N_13847,N_6055,N_6581);
nor U13848 (N_13848,N_7021,N_6330);
nand U13849 (N_13849,N_6161,N_7564);
and U13850 (N_13850,N_7236,N_7938);
nand U13851 (N_13851,N_9605,N_6331);
nor U13852 (N_13852,N_5608,N_6168);
xnor U13853 (N_13853,N_8075,N_9838);
or U13854 (N_13854,N_8661,N_9331);
xor U13855 (N_13855,N_5708,N_9996);
nand U13856 (N_13856,N_8857,N_9132);
nor U13857 (N_13857,N_7656,N_7257);
xnor U13858 (N_13858,N_9235,N_6278);
nand U13859 (N_13859,N_7735,N_6881);
or U13860 (N_13860,N_6212,N_5526);
nand U13861 (N_13861,N_9701,N_5795);
nor U13862 (N_13862,N_8860,N_7956);
nor U13863 (N_13863,N_5289,N_8428);
xnor U13864 (N_13864,N_7637,N_7418);
xor U13865 (N_13865,N_6474,N_9561);
and U13866 (N_13866,N_6828,N_5166);
or U13867 (N_13867,N_9530,N_8787);
or U13868 (N_13868,N_6434,N_5374);
nand U13869 (N_13869,N_8654,N_5168);
nand U13870 (N_13870,N_7399,N_5227);
nor U13871 (N_13871,N_5410,N_8245);
nand U13872 (N_13872,N_9292,N_9772);
xor U13873 (N_13873,N_7739,N_8732);
nand U13874 (N_13874,N_7585,N_5033);
and U13875 (N_13875,N_7088,N_9591);
nand U13876 (N_13876,N_5426,N_5548);
nor U13877 (N_13877,N_5054,N_5778);
xor U13878 (N_13878,N_5018,N_7404);
and U13879 (N_13879,N_7179,N_9738);
xor U13880 (N_13880,N_5961,N_7854);
or U13881 (N_13881,N_6406,N_8217);
nand U13882 (N_13882,N_5421,N_8887);
nand U13883 (N_13883,N_9278,N_9753);
xor U13884 (N_13884,N_8331,N_9558);
or U13885 (N_13885,N_5881,N_5336);
xnor U13886 (N_13886,N_6291,N_8333);
or U13887 (N_13887,N_8911,N_8147);
and U13888 (N_13888,N_6756,N_8685);
nor U13889 (N_13889,N_7588,N_8934);
nand U13890 (N_13890,N_8368,N_7968);
nand U13891 (N_13891,N_8114,N_7999);
or U13892 (N_13892,N_9433,N_5074);
nand U13893 (N_13893,N_9208,N_8118);
nand U13894 (N_13894,N_8434,N_7468);
xor U13895 (N_13895,N_8006,N_9584);
and U13896 (N_13896,N_5453,N_8691);
xnor U13897 (N_13897,N_8665,N_6616);
nor U13898 (N_13898,N_5775,N_7189);
nor U13899 (N_13899,N_9349,N_6312);
nand U13900 (N_13900,N_9327,N_5912);
nand U13901 (N_13901,N_6564,N_7598);
xnor U13902 (N_13902,N_9683,N_8199);
or U13903 (N_13903,N_7497,N_9924);
nand U13904 (N_13904,N_5636,N_9781);
nor U13905 (N_13905,N_5943,N_6719);
or U13906 (N_13906,N_9733,N_8868);
nor U13907 (N_13907,N_6261,N_9752);
nor U13908 (N_13908,N_8348,N_7534);
or U13909 (N_13909,N_7149,N_8497);
xnor U13910 (N_13910,N_8214,N_6395);
and U13911 (N_13911,N_9741,N_8884);
or U13912 (N_13912,N_5668,N_6919);
nor U13913 (N_13913,N_9310,N_9295);
xnor U13914 (N_13914,N_8775,N_8540);
xor U13915 (N_13915,N_6358,N_5395);
nand U13916 (N_13916,N_9204,N_8142);
nand U13917 (N_13917,N_8176,N_6490);
and U13918 (N_13918,N_6063,N_7314);
and U13919 (N_13919,N_5435,N_6625);
nand U13920 (N_13920,N_6717,N_9776);
nand U13921 (N_13921,N_7397,N_5246);
or U13922 (N_13922,N_6774,N_7722);
and U13923 (N_13923,N_5250,N_5975);
xnor U13924 (N_13924,N_8169,N_9808);
nand U13925 (N_13925,N_7369,N_9249);
or U13926 (N_13926,N_5948,N_8712);
and U13927 (N_13927,N_8974,N_9241);
nor U13928 (N_13928,N_9197,N_5826);
xor U13929 (N_13929,N_6848,N_7212);
xor U13930 (N_13930,N_8570,N_5360);
or U13931 (N_13931,N_5125,N_5492);
and U13932 (N_13932,N_9889,N_5242);
nor U13933 (N_13933,N_9487,N_6459);
nand U13934 (N_13934,N_8092,N_7502);
nand U13935 (N_13935,N_6202,N_5078);
nand U13936 (N_13936,N_9098,N_5987);
or U13937 (N_13937,N_5638,N_7170);
nand U13938 (N_13938,N_6569,N_8902);
or U13939 (N_13939,N_8009,N_6412);
nand U13940 (N_13940,N_7556,N_5620);
xnor U13941 (N_13941,N_6136,N_9283);
and U13942 (N_13942,N_7030,N_9547);
xnor U13943 (N_13943,N_5342,N_8529);
nor U13944 (N_13944,N_8769,N_5377);
and U13945 (N_13945,N_7610,N_9812);
nand U13946 (N_13946,N_9227,N_9969);
or U13947 (N_13947,N_7941,N_7168);
or U13948 (N_13948,N_7626,N_5433);
and U13949 (N_13949,N_7412,N_6838);
xnor U13950 (N_13950,N_5571,N_7461);
nor U13951 (N_13951,N_6585,N_7696);
xnor U13952 (N_13952,N_8542,N_9776);
nor U13953 (N_13953,N_6283,N_6785);
xnor U13954 (N_13954,N_9748,N_8824);
or U13955 (N_13955,N_9558,N_9602);
and U13956 (N_13956,N_9118,N_6282);
nor U13957 (N_13957,N_7416,N_7812);
nand U13958 (N_13958,N_6874,N_9258);
nand U13959 (N_13959,N_5086,N_6119);
nor U13960 (N_13960,N_8620,N_6818);
or U13961 (N_13961,N_6576,N_8379);
nor U13962 (N_13962,N_9981,N_8414);
or U13963 (N_13963,N_6866,N_9065);
or U13964 (N_13964,N_9272,N_9228);
nor U13965 (N_13965,N_9988,N_5060);
nor U13966 (N_13966,N_6444,N_7316);
nand U13967 (N_13967,N_5357,N_9078);
nand U13968 (N_13968,N_6741,N_6037);
nand U13969 (N_13969,N_9822,N_5197);
or U13970 (N_13970,N_5058,N_9745);
nor U13971 (N_13971,N_5153,N_6107);
or U13972 (N_13972,N_5393,N_5874);
xor U13973 (N_13973,N_5089,N_8090);
or U13974 (N_13974,N_5904,N_8416);
and U13975 (N_13975,N_9884,N_8434);
xnor U13976 (N_13976,N_7650,N_7021);
xor U13977 (N_13977,N_6339,N_9199);
nand U13978 (N_13978,N_9635,N_6421);
nand U13979 (N_13979,N_9025,N_9212);
or U13980 (N_13980,N_8329,N_7289);
nor U13981 (N_13981,N_8981,N_5615);
nand U13982 (N_13982,N_6844,N_9509);
nor U13983 (N_13983,N_5414,N_9791);
or U13984 (N_13984,N_9161,N_8889);
and U13985 (N_13985,N_6055,N_5703);
xnor U13986 (N_13986,N_6264,N_5027);
xnor U13987 (N_13987,N_8821,N_6577);
nand U13988 (N_13988,N_8145,N_9789);
nor U13989 (N_13989,N_8128,N_9841);
nor U13990 (N_13990,N_6262,N_5317);
xnor U13991 (N_13991,N_9646,N_7639);
xor U13992 (N_13992,N_9293,N_7236);
xnor U13993 (N_13993,N_5237,N_5611);
xnor U13994 (N_13994,N_9240,N_5257);
or U13995 (N_13995,N_5092,N_8433);
xnor U13996 (N_13996,N_7473,N_9373);
nor U13997 (N_13997,N_8007,N_8541);
nor U13998 (N_13998,N_6841,N_9115);
nor U13999 (N_13999,N_6093,N_5523);
and U14000 (N_14000,N_5703,N_5066);
xnor U14001 (N_14001,N_8870,N_5145);
xnor U14002 (N_14002,N_6350,N_5593);
xor U14003 (N_14003,N_6854,N_6387);
nor U14004 (N_14004,N_5129,N_7669);
xor U14005 (N_14005,N_7179,N_5531);
nand U14006 (N_14006,N_7759,N_9215);
nand U14007 (N_14007,N_6904,N_5761);
nand U14008 (N_14008,N_7327,N_8306);
or U14009 (N_14009,N_6015,N_9042);
xnor U14010 (N_14010,N_8448,N_7748);
or U14011 (N_14011,N_9649,N_9352);
or U14012 (N_14012,N_7066,N_5357);
or U14013 (N_14013,N_9299,N_5621);
xor U14014 (N_14014,N_6258,N_5910);
nor U14015 (N_14015,N_5786,N_5299);
nor U14016 (N_14016,N_6788,N_5058);
and U14017 (N_14017,N_6148,N_6278);
xor U14018 (N_14018,N_7634,N_8936);
and U14019 (N_14019,N_9930,N_7861);
nand U14020 (N_14020,N_6779,N_8457);
or U14021 (N_14021,N_9748,N_7745);
and U14022 (N_14022,N_9543,N_9294);
nor U14023 (N_14023,N_7843,N_8197);
nor U14024 (N_14024,N_5183,N_8886);
and U14025 (N_14025,N_5160,N_7760);
nor U14026 (N_14026,N_6583,N_5815);
xnor U14027 (N_14027,N_5631,N_9801);
xor U14028 (N_14028,N_7953,N_5539);
xnor U14029 (N_14029,N_7989,N_6983);
and U14030 (N_14030,N_5837,N_5120);
or U14031 (N_14031,N_6045,N_9685);
and U14032 (N_14032,N_5987,N_5763);
nor U14033 (N_14033,N_8183,N_9258);
nand U14034 (N_14034,N_9579,N_8038);
and U14035 (N_14035,N_6080,N_9965);
or U14036 (N_14036,N_9366,N_7673);
nor U14037 (N_14037,N_6717,N_5650);
nor U14038 (N_14038,N_7616,N_9089);
nand U14039 (N_14039,N_7550,N_7363);
nor U14040 (N_14040,N_9366,N_9627);
nor U14041 (N_14041,N_5599,N_9727);
nor U14042 (N_14042,N_6565,N_8081);
xnor U14043 (N_14043,N_7413,N_7902);
nand U14044 (N_14044,N_6164,N_9200);
nand U14045 (N_14045,N_5137,N_7528);
nor U14046 (N_14046,N_7678,N_5941);
and U14047 (N_14047,N_6860,N_5902);
nor U14048 (N_14048,N_9129,N_7738);
and U14049 (N_14049,N_5637,N_9330);
or U14050 (N_14050,N_6196,N_9438);
nand U14051 (N_14051,N_9111,N_7119);
nor U14052 (N_14052,N_7747,N_9820);
xor U14053 (N_14053,N_9027,N_5662);
nor U14054 (N_14054,N_5949,N_5795);
nand U14055 (N_14055,N_8112,N_7983);
or U14056 (N_14056,N_9752,N_8554);
nor U14057 (N_14057,N_7573,N_6636);
and U14058 (N_14058,N_6110,N_8645);
or U14059 (N_14059,N_5492,N_9239);
xor U14060 (N_14060,N_8001,N_7086);
nor U14061 (N_14061,N_7784,N_6441);
nand U14062 (N_14062,N_6761,N_6284);
or U14063 (N_14063,N_6531,N_8769);
or U14064 (N_14064,N_6755,N_6249);
nand U14065 (N_14065,N_5909,N_5461);
nand U14066 (N_14066,N_8000,N_7963);
nor U14067 (N_14067,N_6937,N_6843);
nand U14068 (N_14068,N_5370,N_7787);
nor U14069 (N_14069,N_5895,N_5401);
xnor U14070 (N_14070,N_7822,N_7960);
nor U14071 (N_14071,N_5340,N_6395);
nor U14072 (N_14072,N_5899,N_9664);
nor U14073 (N_14073,N_9318,N_6423);
or U14074 (N_14074,N_5883,N_5067);
or U14075 (N_14075,N_7310,N_8809);
and U14076 (N_14076,N_5021,N_6779);
nand U14077 (N_14077,N_7957,N_5687);
xor U14078 (N_14078,N_8989,N_8225);
xnor U14079 (N_14079,N_5123,N_6309);
nand U14080 (N_14080,N_5566,N_5332);
nand U14081 (N_14081,N_8176,N_8462);
nand U14082 (N_14082,N_5954,N_5879);
and U14083 (N_14083,N_9937,N_7346);
and U14084 (N_14084,N_6046,N_9858);
nand U14085 (N_14085,N_8383,N_8321);
or U14086 (N_14086,N_8520,N_7689);
xnor U14087 (N_14087,N_5817,N_6913);
xnor U14088 (N_14088,N_9790,N_8871);
or U14089 (N_14089,N_8351,N_9729);
or U14090 (N_14090,N_6687,N_6994);
and U14091 (N_14091,N_7129,N_6356);
nor U14092 (N_14092,N_8341,N_9416);
xnor U14093 (N_14093,N_7831,N_7463);
and U14094 (N_14094,N_7498,N_6129);
nand U14095 (N_14095,N_6704,N_6470);
or U14096 (N_14096,N_8709,N_9473);
nand U14097 (N_14097,N_5806,N_7500);
nor U14098 (N_14098,N_6441,N_9126);
nand U14099 (N_14099,N_8951,N_5646);
nor U14100 (N_14100,N_9411,N_7600);
xor U14101 (N_14101,N_5831,N_7130);
xnor U14102 (N_14102,N_9588,N_6874);
nand U14103 (N_14103,N_9211,N_6252);
nor U14104 (N_14104,N_5993,N_6307);
nor U14105 (N_14105,N_9493,N_9587);
xnor U14106 (N_14106,N_7276,N_5508);
xnor U14107 (N_14107,N_6820,N_8433);
and U14108 (N_14108,N_8699,N_6157);
xor U14109 (N_14109,N_6650,N_9382);
or U14110 (N_14110,N_6336,N_6390);
nand U14111 (N_14111,N_6809,N_7234);
nor U14112 (N_14112,N_6962,N_6435);
nor U14113 (N_14113,N_9737,N_5966);
nand U14114 (N_14114,N_6095,N_6248);
nand U14115 (N_14115,N_7377,N_8217);
xor U14116 (N_14116,N_6540,N_6072);
nand U14117 (N_14117,N_5067,N_9783);
nor U14118 (N_14118,N_5359,N_9770);
xor U14119 (N_14119,N_7002,N_5725);
and U14120 (N_14120,N_6193,N_7733);
and U14121 (N_14121,N_7806,N_7539);
xnor U14122 (N_14122,N_7517,N_8331);
and U14123 (N_14123,N_6410,N_7002);
nor U14124 (N_14124,N_9142,N_6663);
or U14125 (N_14125,N_5859,N_8174);
and U14126 (N_14126,N_6749,N_8784);
nand U14127 (N_14127,N_8164,N_9230);
nand U14128 (N_14128,N_8061,N_6263);
nand U14129 (N_14129,N_6904,N_8388);
nor U14130 (N_14130,N_6380,N_9673);
nor U14131 (N_14131,N_5625,N_5991);
nor U14132 (N_14132,N_7935,N_7814);
nor U14133 (N_14133,N_7967,N_8799);
and U14134 (N_14134,N_7327,N_8181);
and U14135 (N_14135,N_9411,N_8520);
xnor U14136 (N_14136,N_7303,N_7848);
nand U14137 (N_14137,N_5369,N_6173);
or U14138 (N_14138,N_5787,N_5181);
xnor U14139 (N_14139,N_9303,N_7402);
and U14140 (N_14140,N_7673,N_8420);
or U14141 (N_14141,N_6736,N_8665);
nand U14142 (N_14142,N_6861,N_5411);
and U14143 (N_14143,N_8019,N_9773);
nand U14144 (N_14144,N_5165,N_9158);
nor U14145 (N_14145,N_8587,N_7799);
nor U14146 (N_14146,N_8016,N_9134);
nor U14147 (N_14147,N_6367,N_6563);
nand U14148 (N_14148,N_7523,N_8952);
xnor U14149 (N_14149,N_6572,N_8975);
xor U14150 (N_14150,N_6871,N_6839);
nor U14151 (N_14151,N_5485,N_6588);
nor U14152 (N_14152,N_9370,N_8578);
nand U14153 (N_14153,N_8812,N_6363);
and U14154 (N_14154,N_8930,N_9159);
nor U14155 (N_14155,N_8966,N_7058);
and U14156 (N_14156,N_7702,N_7498);
nor U14157 (N_14157,N_5220,N_9457);
and U14158 (N_14158,N_7984,N_7633);
nor U14159 (N_14159,N_9077,N_9237);
nand U14160 (N_14160,N_9181,N_5540);
xnor U14161 (N_14161,N_9355,N_8741);
nor U14162 (N_14162,N_7743,N_6541);
or U14163 (N_14163,N_6245,N_6049);
xnor U14164 (N_14164,N_6205,N_7718);
or U14165 (N_14165,N_7080,N_7452);
nor U14166 (N_14166,N_7470,N_6483);
xor U14167 (N_14167,N_8501,N_9104);
or U14168 (N_14168,N_8563,N_7285);
nor U14169 (N_14169,N_6495,N_8284);
or U14170 (N_14170,N_5847,N_7573);
xnor U14171 (N_14171,N_9620,N_8147);
nand U14172 (N_14172,N_5238,N_7436);
nor U14173 (N_14173,N_6144,N_8755);
and U14174 (N_14174,N_5961,N_5611);
and U14175 (N_14175,N_6799,N_8746);
and U14176 (N_14176,N_9415,N_6768);
or U14177 (N_14177,N_9715,N_5263);
nand U14178 (N_14178,N_5934,N_9280);
xnor U14179 (N_14179,N_8313,N_7530);
and U14180 (N_14180,N_6268,N_6798);
xnor U14181 (N_14181,N_6631,N_5617);
or U14182 (N_14182,N_7373,N_9065);
xnor U14183 (N_14183,N_6080,N_9909);
and U14184 (N_14184,N_5495,N_7201);
xor U14185 (N_14185,N_5227,N_6078);
nor U14186 (N_14186,N_8327,N_8869);
nor U14187 (N_14187,N_5480,N_6309);
nand U14188 (N_14188,N_7944,N_9073);
and U14189 (N_14189,N_9583,N_9862);
nand U14190 (N_14190,N_7986,N_7700);
nand U14191 (N_14191,N_5869,N_5148);
nand U14192 (N_14192,N_8123,N_5812);
and U14193 (N_14193,N_9919,N_8146);
nor U14194 (N_14194,N_9678,N_5473);
and U14195 (N_14195,N_9494,N_5989);
or U14196 (N_14196,N_8250,N_7887);
nand U14197 (N_14197,N_7087,N_9510);
xor U14198 (N_14198,N_7797,N_7227);
or U14199 (N_14199,N_6522,N_9413);
nor U14200 (N_14200,N_6101,N_5111);
nor U14201 (N_14201,N_8592,N_9546);
or U14202 (N_14202,N_9609,N_5519);
nand U14203 (N_14203,N_9542,N_7068);
nor U14204 (N_14204,N_9446,N_6937);
nand U14205 (N_14205,N_6408,N_6640);
and U14206 (N_14206,N_9632,N_6812);
or U14207 (N_14207,N_8794,N_7125);
and U14208 (N_14208,N_9993,N_9194);
nor U14209 (N_14209,N_5202,N_5856);
xnor U14210 (N_14210,N_5490,N_6945);
and U14211 (N_14211,N_6577,N_7996);
xnor U14212 (N_14212,N_9869,N_9158);
and U14213 (N_14213,N_6243,N_5968);
nand U14214 (N_14214,N_9922,N_5353);
and U14215 (N_14215,N_5109,N_9535);
xor U14216 (N_14216,N_5741,N_7814);
nand U14217 (N_14217,N_9647,N_6890);
nor U14218 (N_14218,N_6752,N_8998);
and U14219 (N_14219,N_6517,N_9767);
nand U14220 (N_14220,N_9671,N_6426);
or U14221 (N_14221,N_5550,N_8813);
nor U14222 (N_14222,N_5108,N_5052);
xor U14223 (N_14223,N_7082,N_6682);
nor U14224 (N_14224,N_6730,N_5811);
nand U14225 (N_14225,N_6611,N_6947);
or U14226 (N_14226,N_8203,N_8250);
nor U14227 (N_14227,N_8040,N_8124);
or U14228 (N_14228,N_7918,N_9450);
or U14229 (N_14229,N_8869,N_8220);
or U14230 (N_14230,N_8200,N_7466);
or U14231 (N_14231,N_7918,N_6186);
nor U14232 (N_14232,N_5385,N_9343);
xor U14233 (N_14233,N_9688,N_7443);
nor U14234 (N_14234,N_9687,N_9271);
nand U14235 (N_14235,N_7516,N_7800);
and U14236 (N_14236,N_6070,N_9348);
or U14237 (N_14237,N_6673,N_6960);
nor U14238 (N_14238,N_5214,N_5206);
nand U14239 (N_14239,N_7469,N_5617);
xnor U14240 (N_14240,N_8493,N_6013);
and U14241 (N_14241,N_9993,N_7477);
or U14242 (N_14242,N_5195,N_5568);
nor U14243 (N_14243,N_7920,N_9331);
or U14244 (N_14244,N_6024,N_9074);
and U14245 (N_14245,N_7399,N_5638);
xor U14246 (N_14246,N_8139,N_5014);
or U14247 (N_14247,N_8147,N_9279);
xor U14248 (N_14248,N_7609,N_7086);
xor U14249 (N_14249,N_7283,N_7525);
nand U14250 (N_14250,N_5663,N_5597);
or U14251 (N_14251,N_6599,N_5095);
nand U14252 (N_14252,N_5634,N_6243);
xor U14253 (N_14253,N_9742,N_7989);
nor U14254 (N_14254,N_9255,N_5479);
nor U14255 (N_14255,N_6988,N_7399);
nor U14256 (N_14256,N_5475,N_9517);
nand U14257 (N_14257,N_6970,N_8205);
and U14258 (N_14258,N_9014,N_5079);
xor U14259 (N_14259,N_9122,N_5937);
and U14260 (N_14260,N_7216,N_9656);
nand U14261 (N_14261,N_9036,N_5515);
or U14262 (N_14262,N_5519,N_7155);
nand U14263 (N_14263,N_6114,N_6236);
or U14264 (N_14264,N_7740,N_8087);
xnor U14265 (N_14265,N_6826,N_8165);
nor U14266 (N_14266,N_9466,N_9986);
and U14267 (N_14267,N_7193,N_6495);
nor U14268 (N_14268,N_5200,N_5133);
nor U14269 (N_14269,N_5345,N_5680);
nand U14270 (N_14270,N_7424,N_8680);
and U14271 (N_14271,N_6257,N_5149);
nor U14272 (N_14272,N_7730,N_5333);
and U14273 (N_14273,N_7648,N_8041);
nor U14274 (N_14274,N_5927,N_7795);
nor U14275 (N_14275,N_8824,N_7804);
nand U14276 (N_14276,N_7250,N_9834);
nand U14277 (N_14277,N_8008,N_5426);
nand U14278 (N_14278,N_9344,N_9351);
and U14279 (N_14279,N_5504,N_9992);
nor U14280 (N_14280,N_8812,N_7963);
nand U14281 (N_14281,N_7170,N_8402);
nor U14282 (N_14282,N_7299,N_6633);
and U14283 (N_14283,N_6852,N_8529);
nand U14284 (N_14284,N_6383,N_6658);
nor U14285 (N_14285,N_7896,N_7419);
or U14286 (N_14286,N_7328,N_5978);
and U14287 (N_14287,N_9034,N_8126);
xnor U14288 (N_14288,N_7887,N_7583);
nand U14289 (N_14289,N_8259,N_5664);
nor U14290 (N_14290,N_8413,N_9125);
or U14291 (N_14291,N_9559,N_9890);
xnor U14292 (N_14292,N_9126,N_9849);
and U14293 (N_14293,N_6645,N_7208);
nand U14294 (N_14294,N_9653,N_8698);
and U14295 (N_14295,N_5580,N_5433);
nand U14296 (N_14296,N_6402,N_7785);
and U14297 (N_14297,N_7086,N_5151);
nor U14298 (N_14298,N_6181,N_9395);
or U14299 (N_14299,N_7986,N_5455);
nor U14300 (N_14300,N_7518,N_9287);
and U14301 (N_14301,N_9689,N_5135);
xnor U14302 (N_14302,N_9724,N_9296);
nor U14303 (N_14303,N_7997,N_8163);
nor U14304 (N_14304,N_8535,N_8010);
or U14305 (N_14305,N_9206,N_8960);
or U14306 (N_14306,N_8339,N_8894);
and U14307 (N_14307,N_5728,N_9824);
nand U14308 (N_14308,N_7776,N_6263);
xor U14309 (N_14309,N_7751,N_8291);
xor U14310 (N_14310,N_9582,N_5535);
xor U14311 (N_14311,N_8893,N_5301);
nor U14312 (N_14312,N_9493,N_7219);
or U14313 (N_14313,N_7906,N_5717);
nand U14314 (N_14314,N_8364,N_6721);
and U14315 (N_14315,N_6347,N_7201);
nor U14316 (N_14316,N_9809,N_5247);
nor U14317 (N_14317,N_9974,N_8432);
and U14318 (N_14318,N_9450,N_9494);
and U14319 (N_14319,N_7140,N_7381);
nor U14320 (N_14320,N_7268,N_5399);
and U14321 (N_14321,N_7617,N_8961);
and U14322 (N_14322,N_5891,N_7780);
nand U14323 (N_14323,N_9975,N_9468);
and U14324 (N_14324,N_8441,N_9697);
nor U14325 (N_14325,N_7648,N_8008);
or U14326 (N_14326,N_7614,N_9848);
nand U14327 (N_14327,N_7613,N_7380);
and U14328 (N_14328,N_9683,N_6567);
and U14329 (N_14329,N_9089,N_8023);
nand U14330 (N_14330,N_7528,N_9713);
nor U14331 (N_14331,N_7866,N_7910);
or U14332 (N_14332,N_5665,N_6434);
and U14333 (N_14333,N_6094,N_7514);
xor U14334 (N_14334,N_5128,N_6540);
nand U14335 (N_14335,N_7469,N_9282);
or U14336 (N_14336,N_9767,N_9926);
xnor U14337 (N_14337,N_5111,N_8811);
nor U14338 (N_14338,N_7283,N_8716);
or U14339 (N_14339,N_8484,N_7150);
xnor U14340 (N_14340,N_5172,N_6691);
nor U14341 (N_14341,N_6613,N_8502);
nor U14342 (N_14342,N_7429,N_8290);
and U14343 (N_14343,N_8124,N_6394);
xnor U14344 (N_14344,N_5804,N_7444);
and U14345 (N_14345,N_6047,N_9819);
xor U14346 (N_14346,N_6436,N_5704);
nand U14347 (N_14347,N_7296,N_8247);
xor U14348 (N_14348,N_8463,N_6175);
and U14349 (N_14349,N_8498,N_8348);
nand U14350 (N_14350,N_6629,N_7428);
nor U14351 (N_14351,N_9525,N_8121);
or U14352 (N_14352,N_9413,N_7830);
xor U14353 (N_14353,N_5507,N_8896);
and U14354 (N_14354,N_8806,N_8850);
nand U14355 (N_14355,N_9869,N_6946);
or U14356 (N_14356,N_6214,N_6525);
or U14357 (N_14357,N_9361,N_9226);
and U14358 (N_14358,N_6198,N_7694);
or U14359 (N_14359,N_9664,N_9370);
and U14360 (N_14360,N_8174,N_6078);
and U14361 (N_14361,N_8639,N_8387);
nand U14362 (N_14362,N_8989,N_7386);
and U14363 (N_14363,N_7468,N_5782);
xor U14364 (N_14364,N_8263,N_5032);
nand U14365 (N_14365,N_9985,N_7549);
xor U14366 (N_14366,N_7845,N_7144);
xor U14367 (N_14367,N_7347,N_9160);
xnor U14368 (N_14368,N_8361,N_6208);
nand U14369 (N_14369,N_5542,N_6055);
and U14370 (N_14370,N_8699,N_7051);
or U14371 (N_14371,N_5315,N_5210);
nand U14372 (N_14372,N_7118,N_7998);
nand U14373 (N_14373,N_9374,N_5430);
and U14374 (N_14374,N_7351,N_6710);
nand U14375 (N_14375,N_9469,N_7052);
and U14376 (N_14376,N_9554,N_6025);
nand U14377 (N_14377,N_9151,N_9422);
nor U14378 (N_14378,N_5647,N_8833);
nor U14379 (N_14379,N_9813,N_7647);
nand U14380 (N_14380,N_6137,N_6568);
nand U14381 (N_14381,N_7804,N_8718);
nand U14382 (N_14382,N_8842,N_5545);
nor U14383 (N_14383,N_9459,N_9914);
and U14384 (N_14384,N_6284,N_7416);
xnor U14385 (N_14385,N_8602,N_6048);
nand U14386 (N_14386,N_7216,N_5002);
xor U14387 (N_14387,N_9080,N_8572);
xor U14388 (N_14388,N_7335,N_9631);
and U14389 (N_14389,N_8697,N_6258);
and U14390 (N_14390,N_8195,N_7326);
nor U14391 (N_14391,N_7145,N_6542);
xor U14392 (N_14392,N_5949,N_7191);
xor U14393 (N_14393,N_9585,N_5149);
and U14394 (N_14394,N_5200,N_6998);
nand U14395 (N_14395,N_7959,N_6629);
nor U14396 (N_14396,N_5741,N_7983);
nand U14397 (N_14397,N_7989,N_8034);
and U14398 (N_14398,N_6907,N_7761);
xor U14399 (N_14399,N_6964,N_5885);
and U14400 (N_14400,N_7785,N_7738);
and U14401 (N_14401,N_8734,N_8411);
and U14402 (N_14402,N_5679,N_6140);
and U14403 (N_14403,N_8701,N_6163);
xor U14404 (N_14404,N_5512,N_9066);
or U14405 (N_14405,N_7929,N_5077);
or U14406 (N_14406,N_6103,N_9435);
xnor U14407 (N_14407,N_7068,N_8462);
nand U14408 (N_14408,N_7661,N_6778);
or U14409 (N_14409,N_8037,N_7200);
and U14410 (N_14410,N_9652,N_5424);
and U14411 (N_14411,N_7018,N_7077);
nor U14412 (N_14412,N_7751,N_6085);
xnor U14413 (N_14413,N_6288,N_8625);
or U14414 (N_14414,N_9821,N_5026);
nand U14415 (N_14415,N_6065,N_8618);
and U14416 (N_14416,N_7076,N_6228);
nand U14417 (N_14417,N_9249,N_5401);
or U14418 (N_14418,N_7425,N_8022);
and U14419 (N_14419,N_9228,N_5465);
xnor U14420 (N_14420,N_6773,N_8757);
nand U14421 (N_14421,N_5823,N_9843);
or U14422 (N_14422,N_7277,N_7511);
and U14423 (N_14423,N_6837,N_5795);
or U14424 (N_14424,N_9922,N_7588);
xnor U14425 (N_14425,N_5376,N_7068);
xnor U14426 (N_14426,N_8819,N_5408);
or U14427 (N_14427,N_9394,N_9366);
nor U14428 (N_14428,N_8223,N_9302);
xor U14429 (N_14429,N_8949,N_5292);
nand U14430 (N_14430,N_8216,N_9005);
or U14431 (N_14431,N_9898,N_5931);
xor U14432 (N_14432,N_8879,N_7132);
or U14433 (N_14433,N_8290,N_8550);
nand U14434 (N_14434,N_5926,N_5743);
nor U14435 (N_14435,N_7265,N_7326);
nor U14436 (N_14436,N_7651,N_5133);
nand U14437 (N_14437,N_9693,N_6167);
nand U14438 (N_14438,N_8312,N_9589);
or U14439 (N_14439,N_6337,N_6832);
or U14440 (N_14440,N_7177,N_9288);
xor U14441 (N_14441,N_6510,N_5700);
and U14442 (N_14442,N_6157,N_5530);
and U14443 (N_14443,N_9695,N_5440);
or U14444 (N_14444,N_5124,N_7527);
nand U14445 (N_14445,N_8560,N_5170);
and U14446 (N_14446,N_7258,N_6872);
or U14447 (N_14447,N_7365,N_5977);
or U14448 (N_14448,N_9799,N_9922);
xor U14449 (N_14449,N_7869,N_9724);
or U14450 (N_14450,N_9902,N_7368);
xnor U14451 (N_14451,N_6641,N_9709);
nand U14452 (N_14452,N_8205,N_9481);
and U14453 (N_14453,N_8047,N_6507);
and U14454 (N_14454,N_6393,N_5576);
xnor U14455 (N_14455,N_6712,N_5126);
xor U14456 (N_14456,N_6449,N_5326);
or U14457 (N_14457,N_6404,N_6367);
nand U14458 (N_14458,N_8933,N_9625);
nor U14459 (N_14459,N_6794,N_6074);
and U14460 (N_14460,N_5099,N_6201);
and U14461 (N_14461,N_8191,N_8013);
nand U14462 (N_14462,N_7257,N_8116);
xnor U14463 (N_14463,N_8067,N_9393);
xnor U14464 (N_14464,N_7151,N_5494);
nor U14465 (N_14465,N_9230,N_5573);
nor U14466 (N_14466,N_9177,N_8433);
and U14467 (N_14467,N_9152,N_5262);
or U14468 (N_14468,N_7151,N_5194);
xnor U14469 (N_14469,N_6634,N_9770);
nand U14470 (N_14470,N_6192,N_8448);
and U14471 (N_14471,N_9871,N_5536);
xnor U14472 (N_14472,N_6420,N_7504);
nor U14473 (N_14473,N_5386,N_5934);
xor U14474 (N_14474,N_7746,N_6130);
and U14475 (N_14475,N_8999,N_9858);
or U14476 (N_14476,N_7113,N_9659);
xor U14477 (N_14477,N_5832,N_6636);
xnor U14478 (N_14478,N_6098,N_9836);
nand U14479 (N_14479,N_5749,N_9704);
nand U14480 (N_14480,N_8632,N_8563);
nor U14481 (N_14481,N_7454,N_8579);
and U14482 (N_14482,N_9286,N_9593);
and U14483 (N_14483,N_9370,N_8008);
and U14484 (N_14484,N_8424,N_8296);
xor U14485 (N_14485,N_9680,N_8143);
nand U14486 (N_14486,N_5935,N_6338);
nor U14487 (N_14487,N_9665,N_9378);
xnor U14488 (N_14488,N_8038,N_5659);
or U14489 (N_14489,N_7935,N_6634);
nand U14490 (N_14490,N_6080,N_6583);
xor U14491 (N_14491,N_7969,N_8968);
or U14492 (N_14492,N_9271,N_9390);
nor U14493 (N_14493,N_6977,N_5220);
and U14494 (N_14494,N_9849,N_5428);
and U14495 (N_14495,N_5691,N_8735);
nor U14496 (N_14496,N_6730,N_9673);
and U14497 (N_14497,N_9629,N_7324);
nand U14498 (N_14498,N_9997,N_5464);
xor U14499 (N_14499,N_7300,N_5261);
and U14500 (N_14500,N_5201,N_6199);
and U14501 (N_14501,N_9491,N_5779);
or U14502 (N_14502,N_9156,N_8390);
or U14503 (N_14503,N_6238,N_8759);
xnor U14504 (N_14504,N_7940,N_9811);
or U14505 (N_14505,N_9309,N_9916);
nor U14506 (N_14506,N_5151,N_9410);
nand U14507 (N_14507,N_8633,N_6135);
nor U14508 (N_14508,N_8599,N_7866);
nand U14509 (N_14509,N_8850,N_9191);
nand U14510 (N_14510,N_7098,N_9972);
or U14511 (N_14511,N_9442,N_7536);
or U14512 (N_14512,N_8411,N_8994);
and U14513 (N_14513,N_6591,N_8417);
and U14514 (N_14514,N_6087,N_9939);
nand U14515 (N_14515,N_7428,N_8041);
or U14516 (N_14516,N_9976,N_5774);
or U14517 (N_14517,N_7650,N_5899);
and U14518 (N_14518,N_7215,N_9172);
nand U14519 (N_14519,N_6389,N_9826);
xor U14520 (N_14520,N_5842,N_6000);
nand U14521 (N_14521,N_5075,N_8013);
nand U14522 (N_14522,N_8825,N_8752);
nand U14523 (N_14523,N_6988,N_5862);
nor U14524 (N_14524,N_5575,N_7217);
and U14525 (N_14525,N_5961,N_9711);
nand U14526 (N_14526,N_6874,N_7446);
and U14527 (N_14527,N_6811,N_8172);
nor U14528 (N_14528,N_7650,N_7361);
xnor U14529 (N_14529,N_8145,N_6237);
xor U14530 (N_14530,N_6555,N_9635);
nand U14531 (N_14531,N_8438,N_8981);
nand U14532 (N_14532,N_8345,N_9209);
xnor U14533 (N_14533,N_7950,N_7422);
nand U14534 (N_14534,N_9520,N_5296);
and U14535 (N_14535,N_9966,N_6362);
or U14536 (N_14536,N_7932,N_7121);
nor U14537 (N_14537,N_9058,N_6125);
nor U14538 (N_14538,N_9551,N_5299);
or U14539 (N_14539,N_7397,N_9986);
and U14540 (N_14540,N_8183,N_5165);
or U14541 (N_14541,N_7872,N_5946);
and U14542 (N_14542,N_6810,N_6389);
and U14543 (N_14543,N_7302,N_7165);
or U14544 (N_14544,N_5868,N_9700);
xnor U14545 (N_14545,N_8327,N_5196);
nand U14546 (N_14546,N_7765,N_8656);
and U14547 (N_14547,N_9554,N_9531);
or U14548 (N_14548,N_8088,N_7762);
and U14549 (N_14549,N_8732,N_6776);
and U14550 (N_14550,N_8786,N_6407);
or U14551 (N_14551,N_5330,N_6745);
xor U14552 (N_14552,N_8148,N_9500);
and U14553 (N_14553,N_7347,N_5790);
or U14554 (N_14554,N_6370,N_8622);
nand U14555 (N_14555,N_5087,N_8770);
nand U14556 (N_14556,N_9358,N_6142);
or U14557 (N_14557,N_8624,N_6112);
and U14558 (N_14558,N_8857,N_9849);
nand U14559 (N_14559,N_6633,N_7595);
or U14560 (N_14560,N_5651,N_6932);
xor U14561 (N_14561,N_7109,N_6572);
xnor U14562 (N_14562,N_8992,N_9283);
xnor U14563 (N_14563,N_7962,N_9452);
nand U14564 (N_14564,N_9077,N_8750);
and U14565 (N_14565,N_8252,N_5047);
xnor U14566 (N_14566,N_6151,N_5047);
nand U14567 (N_14567,N_7550,N_9718);
nand U14568 (N_14568,N_7522,N_6748);
nand U14569 (N_14569,N_6949,N_8250);
or U14570 (N_14570,N_5782,N_5147);
and U14571 (N_14571,N_7679,N_7854);
nand U14572 (N_14572,N_9568,N_7244);
and U14573 (N_14573,N_9525,N_7887);
nor U14574 (N_14574,N_5076,N_9755);
and U14575 (N_14575,N_5644,N_8105);
xnor U14576 (N_14576,N_7414,N_5665);
xor U14577 (N_14577,N_8698,N_6154);
and U14578 (N_14578,N_9393,N_6405);
or U14579 (N_14579,N_9132,N_9894);
and U14580 (N_14580,N_9313,N_9067);
xor U14581 (N_14581,N_8735,N_6031);
xnor U14582 (N_14582,N_8456,N_7240);
xnor U14583 (N_14583,N_7359,N_9957);
nand U14584 (N_14584,N_6474,N_7454);
nand U14585 (N_14585,N_6294,N_9017);
nand U14586 (N_14586,N_9406,N_7889);
nor U14587 (N_14587,N_9265,N_9904);
or U14588 (N_14588,N_5144,N_5603);
or U14589 (N_14589,N_9084,N_9096);
nor U14590 (N_14590,N_7128,N_8777);
nand U14591 (N_14591,N_7762,N_9286);
or U14592 (N_14592,N_9867,N_9706);
nand U14593 (N_14593,N_6924,N_5453);
and U14594 (N_14594,N_5010,N_9534);
xnor U14595 (N_14595,N_9884,N_5834);
xnor U14596 (N_14596,N_5371,N_6764);
nand U14597 (N_14597,N_5904,N_9895);
nand U14598 (N_14598,N_7857,N_5338);
nand U14599 (N_14599,N_5802,N_8428);
xnor U14600 (N_14600,N_7024,N_5327);
and U14601 (N_14601,N_9639,N_8572);
or U14602 (N_14602,N_5604,N_5378);
and U14603 (N_14603,N_6386,N_8581);
or U14604 (N_14604,N_6803,N_6012);
xnor U14605 (N_14605,N_9248,N_9432);
xor U14606 (N_14606,N_9030,N_6258);
nor U14607 (N_14607,N_8977,N_7780);
and U14608 (N_14608,N_7808,N_5075);
nand U14609 (N_14609,N_6998,N_9474);
nor U14610 (N_14610,N_5098,N_8938);
and U14611 (N_14611,N_8858,N_6335);
xor U14612 (N_14612,N_5342,N_9592);
nand U14613 (N_14613,N_5178,N_8163);
xor U14614 (N_14614,N_7373,N_5089);
and U14615 (N_14615,N_9929,N_6077);
xnor U14616 (N_14616,N_6033,N_7771);
and U14617 (N_14617,N_5879,N_9312);
or U14618 (N_14618,N_8682,N_5097);
or U14619 (N_14619,N_7672,N_6855);
xnor U14620 (N_14620,N_8383,N_5988);
or U14621 (N_14621,N_8324,N_6976);
or U14622 (N_14622,N_5926,N_9435);
nor U14623 (N_14623,N_5477,N_9883);
or U14624 (N_14624,N_6873,N_6908);
or U14625 (N_14625,N_7411,N_6466);
and U14626 (N_14626,N_5860,N_5997);
nor U14627 (N_14627,N_5528,N_8161);
nand U14628 (N_14628,N_8249,N_6753);
and U14629 (N_14629,N_8415,N_6642);
nor U14630 (N_14630,N_8654,N_7805);
or U14631 (N_14631,N_7966,N_9373);
nand U14632 (N_14632,N_9601,N_6086);
and U14633 (N_14633,N_7056,N_6396);
nor U14634 (N_14634,N_9927,N_9433);
nor U14635 (N_14635,N_7035,N_8275);
or U14636 (N_14636,N_7618,N_5309);
nand U14637 (N_14637,N_6443,N_7062);
or U14638 (N_14638,N_5316,N_6996);
or U14639 (N_14639,N_8761,N_5765);
or U14640 (N_14640,N_8268,N_9307);
nor U14641 (N_14641,N_9167,N_5723);
and U14642 (N_14642,N_9092,N_8904);
xor U14643 (N_14643,N_7506,N_6883);
nand U14644 (N_14644,N_7154,N_7596);
xor U14645 (N_14645,N_6265,N_7583);
nor U14646 (N_14646,N_6718,N_7882);
or U14647 (N_14647,N_6464,N_5014);
nand U14648 (N_14648,N_7575,N_5200);
or U14649 (N_14649,N_9227,N_5005);
nor U14650 (N_14650,N_6625,N_8025);
and U14651 (N_14651,N_7977,N_7233);
xnor U14652 (N_14652,N_7679,N_5320);
xor U14653 (N_14653,N_6686,N_7535);
nor U14654 (N_14654,N_9295,N_8207);
nor U14655 (N_14655,N_7156,N_5182);
nor U14656 (N_14656,N_5568,N_9630);
nor U14657 (N_14657,N_7403,N_8597);
or U14658 (N_14658,N_5660,N_7531);
xor U14659 (N_14659,N_7986,N_7046);
nor U14660 (N_14660,N_8060,N_8985);
xnor U14661 (N_14661,N_7952,N_5987);
and U14662 (N_14662,N_8171,N_9355);
or U14663 (N_14663,N_6963,N_5207);
nor U14664 (N_14664,N_7248,N_8748);
and U14665 (N_14665,N_9477,N_5148);
and U14666 (N_14666,N_5535,N_5387);
or U14667 (N_14667,N_8448,N_9769);
nand U14668 (N_14668,N_8424,N_5914);
or U14669 (N_14669,N_9473,N_7338);
and U14670 (N_14670,N_7215,N_5650);
nand U14671 (N_14671,N_9034,N_7756);
xnor U14672 (N_14672,N_5445,N_8751);
nand U14673 (N_14673,N_9137,N_7656);
or U14674 (N_14674,N_9930,N_6616);
or U14675 (N_14675,N_6816,N_7676);
nand U14676 (N_14676,N_5668,N_5154);
nand U14677 (N_14677,N_9765,N_8931);
xor U14678 (N_14678,N_6866,N_9901);
nor U14679 (N_14679,N_5911,N_9173);
and U14680 (N_14680,N_9429,N_9029);
nor U14681 (N_14681,N_6839,N_7927);
and U14682 (N_14682,N_7733,N_5533);
nor U14683 (N_14683,N_6567,N_8383);
and U14684 (N_14684,N_7507,N_8779);
or U14685 (N_14685,N_5510,N_9127);
xor U14686 (N_14686,N_7942,N_7361);
and U14687 (N_14687,N_6267,N_6432);
nand U14688 (N_14688,N_8182,N_7141);
nor U14689 (N_14689,N_7657,N_7866);
xnor U14690 (N_14690,N_9136,N_6915);
nor U14691 (N_14691,N_7582,N_5316);
nand U14692 (N_14692,N_9627,N_8074);
nor U14693 (N_14693,N_9238,N_8223);
xnor U14694 (N_14694,N_8435,N_7700);
nor U14695 (N_14695,N_8624,N_7744);
and U14696 (N_14696,N_6536,N_7026);
and U14697 (N_14697,N_6596,N_9092);
or U14698 (N_14698,N_7568,N_6672);
and U14699 (N_14699,N_5436,N_9737);
and U14700 (N_14700,N_6473,N_7180);
nand U14701 (N_14701,N_9645,N_8192);
or U14702 (N_14702,N_7564,N_5704);
or U14703 (N_14703,N_8593,N_6561);
xor U14704 (N_14704,N_8624,N_9768);
nor U14705 (N_14705,N_9320,N_5199);
xor U14706 (N_14706,N_8510,N_8957);
nand U14707 (N_14707,N_9395,N_8009);
xor U14708 (N_14708,N_9070,N_6221);
and U14709 (N_14709,N_6035,N_9200);
and U14710 (N_14710,N_8010,N_9608);
xor U14711 (N_14711,N_8381,N_7729);
nor U14712 (N_14712,N_7005,N_8486);
or U14713 (N_14713,N_9427,N_9915);
nand U14714 (N_14714,N_6308,N_8434);
nand U14715 (N_14715,N_6689,N_6913);
or U14716 (N_14716,N_8109,N_5203);
or U14717 (N_14717,N_5625,N_7032);
and U14718 (N_14718,N_7738,N_7002);
and U14719 (N_14719,N_8299,N_8836);
nand U14720 (N_14720,N_8991,N_9953);
and U14721 (N_14721,N_8861,N_9146);
or U14722 (N_14722,N_8877,N_8850);
xor U14723 (N_14723,N_6880,N_5690);
xor U14724 (N_14724,N_7241,N_6111);
xor U14725 (N_14725,N_9762,N_6707);
nand U14726 (N_14726,N_6815,N_5449);
nand U14727 (N_14727,N_9582,N_5046);
nor U14728 (N_14728,N_6018,N_9186);
or U14729 (N_14729,N_7946,N_5942);
nand U14730 (N_14730,N_5136,N_9816);
nor U14731 (N_14731,N_6272,N_9160);
or U14732 (N_14732,N_9499,N_7990);
xor U14733 (N_14733,N_6715,N_9894);
xnor U14734 (N_14734,N_5604,N_5882);
nor U14735 (N_14735,N_9164,N_6526);
nor U14736 (N_14736,N_6803,N_9417);
nor U14737 (N_14737,N_6787,N_6858);
nor U14738 (N_14738,N_8239,N_8223);
or U14739 (N_14739,N_8047,N_7233);
and U14740 (N_14740,N_6585,N_7634);
nand U14741 (N_14741,N_8536,N_8540);
xnor U14742 (N_14742,N_8686,N_5183);
and U14743 (N_14743,N_8903,N_8879);
or U14744 (N_14744,N_5691,N_5561);
xnor U14745 (N_14745,N_7870,N_8864);
nand U14746 (N_14746,N_9029,N_9828);
and U14747 (N_14747,N_8213,N_7405);
or U14748 (N_14748,N_6407,N_9551);
and U14749 (N_14749,N_9477,N_5714);
or U14750 (N_14750,N_6855,N_9865);
nand U14751 (N_14751,N_6891,N_6780);
nor U14752 (N_14752,N_5277,N_7735);
nand U14753 (N_14753,N_5222,N_9360);
xnor U14754 (N_14754,N_6829,N_7057);
xnor U14755 (N_14755,N_9850,N_5590);
and U14756 (N_14756,N_6057,N_9858);
nand U14757 (N_14757,N_6606,N_8010);
xor U14758 (N_14758,N_7790,N_6456);
nand U14759 (N_14759,N_7498,N_6494);
xor U14760 (N_14760,N_8147,N_8656);
nand U14761 (N_14761,N_9313,N_9328);
and U14762 (N_14762,N_8090,N_8533);
and U14763 (N_14763,N_5443,N_5441);
nor U14764 (N_14764,N_7934,N_6170);
xnor U14765 (N_14765,N_9200,N_9143);
xor U14766 (N_14766,N_7639,N_6451);
or U14767 (N_14767,N_7827,N_7343);
nand U14768 (N_14768,N_5584,N_5995);
xnor U14769 (N_14769,N_6711,N_9909);
or U14770 (N_14770,N_6081,N_5124);
xnor U14771 (N_14771,N_7164,N_8330);
and U14772 (N_14772,N_9371,N_7305);
nand U14773 (N_14773,N_9355,N_7837);
and U14774 (N_14774,N_8026,N_8389);
or U14775 (N_14775,N_7451,N_7298);
nand U14776 (N_14776,N_7303,N_8152);
and U14777 (N_14777,N_8673,N_8004);
nand U14778 (N_14778,N_9176,N_8431);
nand U14779 (N_14779,N_7325,N_7122);
nor U14780 (N_14780,N_6793,N_5047);
xor U14781 (N_14781,N_7214,N_9076);
nand U14782 (N_14782,N_7992,N_8391);
xnor U14783 (N_14783,N_8177,N_6358);
nor U14784 (N_14784,N_7622,N_9940);
or U14785 (N_14785,N_9286,N_8839);
nor U14786 (N_14786,N_8751,N_7127);
nor U14787 (N_14787,N_6210,N_5966);
or U14788 (N_14788,N_5488,N_7911);
nand U14789 (N_14789,N_6013,N_6570);
nor U14790 (N_14790,N_8476,N_5022);
xnor U14791 (N_14791,N_6648,N_5705);
nand U14792 (N_14792,N_8213,N_6594);
nor U14793 (N_14793,N_8447,N_8712);
nor U14794 (N_14794,N_6948,N_9376);
or U14795 (N_14795,N_5314,N_7396);
and U14796 (N_14796,N_7516,N_6947);
nand U14797 (N_14797,N_8620,N_8885);
nand U14798 (N_14798,N_9484,N_9768);
or U14799 (N_14799,N_9105,N_9797);
or U14800 (N_14800,N_7453,N_8919);
nand U14801 (N_14801,N_9820,N_6687);
nor U14802 (N_14802,N_5969,N_6363);
nor U14803 (N_14803,N_5214,N_5140);
xor U14804 (N_14804,N_9725,N_7593);
and U14805 (N_14805,N_7633,N_7690);
xnor U14806 (N_14806,N_7298,N_8204);
and U14807 (N_14807,N_6659,N_8690);
or U14808 (N_14808,N_6628,N_5835);
or U14809 (N_14809,N_6783,N_8055);
and U14810 (N_14810,N_9645,N_7488);
xnor U14811 (N_14811,N_9809,N_7311);
or U14812 (N_14812,N_8941,N_5346);
and U14813 (N_14813,N_8922,N_9481);
xor U14814 (N_14814,N_9563,N_7224);
nor U14815 (N_14815,N_8877,N_6391);
or U14816 (N_14816,N_7202,N_7321);
nand U14817 (N_14817,N_9983,N_8426);
nand U14818 (N_14818,N_8103,N_7457);
xor U14819 (N_14819,N_5231,N_6405);
and U14820 (N_14820,N_8408,N_6442);
and U14821 (N_14821,N_7218,N_5668);
xor U14822 (N_14822,N_7620,N_8844);
or U14823 (N_14823,N_9265,N_9727);
or U14824 (N_14824,N_7599,N_9519);
and U14825 (N_14825,N_6193,N_9142);
and U14826 (N_14826,N_5080,N_5820);
nor U14827 (N_14827,N_9725,N_9727);
or U14828 (N_14828,N_8871,N_6010);
nor U14829 (N_14829,N_9411,N_7714);
xor U14830 (N_14830,N_9662,N_5310);
xnor U14831 (N_14831,N_5726,N_6454);
nand U14832 (N_14832,N_5057,N_8365);
xor U14833 (N_14833,N_8314,N_7235);
or U14834 (N_14834,N_9709,N_7058);
nor U14835 (N_14835,N_5077,N_8446);
nor U14836 (N_14836,N_9306,N_6520);
nor U14837 (N_14837,N_7697,N_9711);
or U14838 (N_14838,N_7102,N_5353);
or U14839 (N_14839,N_6025,N_5021);
nand U14840 (N_14840,N_6799,N_8304);
xor U14841 (N_14841,N_9089,N_5546);
nand U14842 (N_14842,N_7449,N_5614);
nor U14843 (N_14843,N_8516,N_8914);
or U14844 (N_14844,N_7651,N_5483);
nor U14845 (N_14845,N_8998,N_8018);
nor U14846 (N_14846,N_9123,N_9435);
or U14847 (N_14847,N_9221,N_5038);
and U14848 (N_14848,N_8561,N_5858);
nor U14849 (N_14849,N_8684,N_9186);
nand U14850 (N_14850,N_7610,N_7433);
or U14851 (N_14851,N_5070,N_8285);
nand U14852 (N_14852,N_5675,N_9652);
nand U14853 (N_14853,N_6744,N_6115);
or U14854 (N_14854,N_8903,N_5435);
nor U14855 (N_14855,N_6157,N_7568);
or U14856 (N_14856,N_8291,N_6249);
nand U14857 (N_14857,N_6275,N_5786);
and U14858 (N_14858,N_8688,N_6560);
xor U14859 (N_14859,N_6894,N_8790);
and U14860 (N_14860,N_5449,N_5974);
and U14861 (N_14861,N_5571,N_5971);
or U14862 (N_14862,N_7715,N_6436);
and U14863 (N_14863,N_8061,N_5203);
xnor U14864 (N_14864,N_6280,N_9797);
and U14865 (N_14865,N_8996,N_5199);
or U14866 (N_14866,N_9787,N_9484);
nand U14867 (N_14867,N_6372,N_5487);
nand U14868 (N_14868,N_9789,N_7903);
or U14869 (N_14869,N_9783,N_9057);
xnor U14870 (N_14870,N_7778,N_5880);
xor U14871 (N_14871,N_7585,N_5295);
nor U14872 (N_14872,N_5995,N_7270);
or U14873 (N_14873,N_9924,N_6268);
or U14874 (N_14874,N_9164,N_9407);
xnor U14875 (N_14875,N_9046,N_6254);
nor U14876 (N_14876,N_7135,N_8068);
nor U14877 (N_14877,N_7125,N_5489);
xnor U14878 (N_14878,N_7299,N_9464);
nand U14879 (N_14879,N_7544,N_8498);
and U14880 (N_14880,N_7544,N_9163);
nand U14881 (N_14881,N_7914,N_5520);
and U14882 (N_14882,N_8667,N_5914);
nor U14883 (N_14883,N_9751,N_6592);
and U14884 (N_14884,N_5784,N_8229);
nor U14885 (N_14885,N_6230,N_6432);
xnor U14886 (N_14886,N_6893,N_8872);
nor U14887 (N_14887,N_6426,N_7979);
and U14888 (N_14888,N_5887,N_8036);
or U14889 (N_14889,N_7522,N_6279);
or U14890 (N_14890,N_9453,N_8537);
or U14891 (N_14891,N_8069,N_7123);
nor U14892 (N_14892,N_5406,N_5782);
nor U14893 (N_14893,N_6585,N_9186);
xor U14894 (N_14894,N_9351,N_9714);
and U14895 (N_14895,N_5903,N_8794);
xnor U14896 (N_14896,N_9398,N_5427);
and U14897 (N_14897,N_6505,N_5356);
and U14898 (N_14898,N_8540,N_7876);
and U14899 (N_14899,N_5121,N_6530);
nor U14900 (N_14900,N_6304,N_5298);
and U14901 (N_14901,N_6813,N_8139);
nor U14902 (N_14902,N_7919,N_5026);
nor U14903 (N_14903,N_5078,N_7027);
and U14904 (N_14904,N_8712,N_5447);
nand U14905 (N_14905,N_5628,N_6240);
nor U14906 (N_14906,N_6163,N_8127);
nand U14907 (N_14907,N_7355,N_9996);
or U14908 (N_14908,N_9364,N_9433);
nand U14909 (N_14909,N_5560,N_5007);
nand U14910 (N_14910,N_7809,N_8237);
nor U14911 (N_14911,N_7890,N_6387);
or U14912 (N_14912,N_5405,N_8842);
xnor U14913 (N_14913,N_8302,N_8238);
or U14914 (N_14914,N_5320,N_5433);
nand U14915 (N_14915,N_7658,N_9435);
nor U14916 (N_14916,N_8346,N_6287);
nor U14917 (N_14917,N_9195,N_9166);
nor U14918 (N_14918,N_8209,N_9932);
or U14919 (N_14919,N_6284,N_7477);
nand U14920 (N_14920,N_9940,N_6252);
and U14921 (N_14921,N_8429,N_7064);
nand U14922 (N_14922,N_9309,N_8990);
and U14923 (N_14923,N_9636,N_9327);
and U14924 (N_14924,N_7495,N_5669);
or U14925 (N_14925,N_6075,N_9999);
xnor U14926 (N_14926,N_5511,N_8616);
nand U14927 (N_14927,N_7818,N_7244);
and U14928 (N_14928,N_6067,N_7240);
nand U14929 (N_14929,N_5728,N_5720);
xnor U14930 (N_14930,N_5988,N_9107);
and U14931 (N_14931,N_7532,N_7561);
nor U14932 (N_14932,N_9350,N_7968);
xnor U14933 (N_14933,N_6576,N_9396);
xnor U14934 (N_14934,N_7748,N_8700);
nor U14935 (N_14935,N_8330,N_9859);
and U14936 (N_14936,N_7390,N_7640);
and U14937 (N_14937,N_6310,N_6366);
and U14938 (N_14938,N_8064,N_7561);
and U14939 (N_14939,N_6258,N_8932);
nand U14940 (N_14940,N_6375,N_5329);
xnor U14941 (N_14941,N_5317,N_8521);
nand U14942 (N_14942,N_7415,N_8091);
and U14943 (N_14943,N_5961,N_7443);
and U14944 (N_14944,N_5211,N_5461);
nor U14945 (N_14945,N_7967,N_7309);
and U14946 (N_14946,N_5377,N_9689);
nor U14947 (N_14947,N_5996,N_5754);
or U14948 (N_14948,N_8494,N_8357);
or U14949 (N_14949,N_8619,N_5901);
or U14950 (N_14950,N_9009,N_9390);
nand U14951 (N_14951,N_9478,N_7284);
nor U14952 (N_14952,N_6784,N_9627);
nor U14953 (N_14953,N_9267,N_9148);
and U14954 (N_14954,N_7232,N_6213);
nand U14955 (N_14955,N_7837,N_5975);
and U14956 (N_14956,N_8733,N_5674);
nor U14957 (N_14957,N_8095,N_5600);
and U14958 (N_14958,N_9787,N_9346);
or U14959 (N_14959,N_9103,N_6107);
or U14960 (N_14960,N_7242,N_5286);
or U14961 (N_14961,N_9790,N_6802);
and U14962 (N_14962,N_8651,N_5338);
nor U14963 (N_14963,N_8624,N_9248);
and U14964 (N_14964,N_6048,N_8515);
and U14965 (N_14965,N_8009,N_7561);
or U14966 (N_14966,N_5472,N_9584);
nor U14967 (N_14967,N_9052,N_8012);
and U14968 (N_14968,N_7004,N_5489);
nor U14969 (N_14969,N_9643,N_7589);
and U14970 (N_14970,N_5231,N_7629);
nand U14971 (N_14971,N_7791,N_6125);
nor U14972 (N_14972,N_7496,N_9739);
or U14973 (N_14973,N_8346,N_6127);
nand U14974 (N_14974,N_9592,N_9593);
or U14975 (N_14975,N_5847,N_6214);
and U14976 (N_14976,N_5195,N_6298);
nor U14977 (N_14977,N_5789,N_8343);
or U14978 (N_14978,N_9520,N_9081);
nor U14979 (N_14979,N_5543,N_6603);
xor U14980 (N_14980,N_9949,N_5406);
xor U14981 (N_14981,N_9120,N_7674);
and U14982 (N_14982,N_6382,N_8182);
xor U14983 (N_14983,N_8565,N_5955);
nor U14984 (N_14984,N_6642,N_5211);
nor U14985 (N_14985,N_8960,N_6034);
xnor U14986 (N_14986,N_6149,N_8366);
nand U14987 (N_14987,N_7954,N_8157);
and U14988 (N_14988,N_6411,N_5105);
or U14989 (N_14989,N_9221,N_6870);
or U14990 (N_14990,N_9503,N_8591);
and U14991 (N_14991,N_8212,N_8508);
xnor U14992 (N_14992,N_5982,N_5302);
and U14993 (N_14993,N_9493,N_6822);
xor U14994 (N_14994,N_8774,N_7163);
nand U14995 (N_14995,N_8314,N_9446);
xnor U14996 (N_14996,N_7433,N_9733);
and U14997 (N_14997,N_6695,N_5633);
nand U14998 (N_14998,N_8966,N_5506);
and U14999 (N_14999,N_6612,N_5603);
and U15000 (N_15000,N_12013,N_13684);
nand U15001 (N_15001,N_14873,N_12344);
and U15002 (N_15002,N_14224,N_11843);
nor U15003 (N_15003,N_13104,N_11120);
nand U15004 (N_15004,N_10425,N_11516);
nand U15005 (N_15005,N_10084,N_14513);
and U15006 (N_15006,N_13616,N_13846);
nand U15007 (N_15007,N_13119,N_11114);
or U15008 (N_15008,N_11102,N_14280);
nand U15009 (N_15009,N_13754,N_10810);
xor U15010 (N_15010,N_13664,N_11395);
nand U15011 (N_15011,N_14727,N_12882);
or U15012 (N_15012,N_12726,N_14980);
xnor U15013 (N_15013,N_11530,N_11468);
or U15014 (N_15014,N_12914,N_11913);
nor U15015 (N_15015,N_13940,N_11064);
and U15016 (N_15016,N_11668,N_14834);
nand U15017 (N_15017,N_13831,N_11579);
xnor U15018 (N_15018,N_12850,N_14916);
xor U15019 (N_15019,N_11664,N_11452);
and U15020 (N_15020,N_13612,N_11893);
nor U15021 (N_15021,N_14248,N_11820);
nand U15022 (N_15022,N_13400,N_10107);
nand U15023 (N_15023,N_13303,N_10748);
or U15024 (N_15024,N_11405,N_14522);
nand U15025 (N_15025,N_11385,N_11968);
nor U15026 (N_15026,N_14386,N_12301);
xnor U15027 (N_15027,N_13880,N_13385);
nand U15028 (N_15028,N_12753,N_10462);
nor U15029 (N_15029,N_12091,N_12052);
and U15030 (N_15030,N_13062,N_10141);
nor U15031 (N_15031,N_13339,N_11137);
xor U15032 (N_15032,N_14935,N_12967);
nor U15033 (N_15033,N_14125,N_11854);
or U15034 (N_15034,N_12051,N_10782);
xor U15035 (N_15035,N_12075,N_11510);
and U15036 (N_15036,N_12266,N_13023);
xnor U15037 (N_15037,N_10880,N_14880);
or U15038 (N_15038,N_11979,N_10453);
and U15039 (N_15039,N_13561,N_10696);
nand U15040 (N_15040,N_11814,N_14237);
or U15041 (N_15041,N_13092,N_13558);
or U15042 (N_15042,N_10223,N_10972);
nor U15043 (N_15043,N_13437,N_10088);
xnor U15044 (N_15044,N_14221,N_11790);
and U15045 (N_15045,N_10280,N_13990);
xor U15046 (N_15046,N_14740,N_11315);
nand U15047 (N_15047,N_10564,N_14694);
nand U15048 (N_15048,N_10197,N_12021);
xnor U15049 (N_15049,N_13228,N_14745);
nor U15050 (N_15050,N_14913,N_14432);
or U15051 (N_15051,N_10275,N_14380);
and U15052 (N_15052,N_14064,N_10302);
nand U15053 (N_15053,N_12233,N_11836);
xor U15054 (N_15054,N_13607,N_12763);
nor U15055 (N_15055,N_11795,N_10298);
nand U15056 (N_15056,N_12062,N_12210);
nor U15057 (N_15057,N_10733,N_11063);
and U15058 (N_15058,N_13251,N_12035);
and U15059 (N_15059,N_12134,N_12137);
xnor U15060 (N_15060,N_13703,N_10850);
and U15061 (N_15061,N_10556,N_14708);
nand U15062 (N_15062,N_11911,N_11841);
nor U15063 (N_15063,N_11691,N_14832);
xor U15064 (N_15064,N_11016,N_13806);
nor U15065 (N_15065,N_12949,N_14648);
nand U15066 (N_15066,N_11475,N_13589);
xor U15067 (N_15067,N_14074,N_12450);
nand U15068 (N_15068,N_11927,N_13999);
and U15069 (N_15069,N_12620,N_10473);
xor U15070 (N_15070,N_10747,N_13924);
nand U15071 (N_15071,N_14228,N_12343);
nand U15072 (N_15072,N_13549,N_11950);
xor U15073 (N_15073,N_10798,N_12001);
xor U15074 (N_15074,N_10382,N_13243);
xnor U15075 (N_15075,N_14122,N_13903);
nand U15076 (N_15076,N_13959,N_14545);
and U15077 (N_15077,N_12599,N_14375);
and U15078 (N_15078,N_12800,N_10918);
xnor U15079 (N_15079,N_13048,N_10185);
nand U15080 (N_15080,N_12182,N_13888);
nand U15081 (N_15081,N_14863,N_13256);
nor U15082 (N_15082,N_13517,N_10418);
nor U15083 (N_15083,N_13227,N_11878);
and U15084 (N_15084,N_11073,N_14210);
nor U15085 (N_15085,N_10091,N_12398);
nand U15086 (N_15086,N_11986,N_10006);
nand U15087 (N_15087,N_14554,N_10270);
xor U15088 (N_15088,N_10492,N_13186);
or U15089 (N_15089,N_13816,N_12567);
nand U15090 (N_15090,N_14267,N_14958);
nor U15091 (N_15091,N_10593,N_11519);
xor U15092 (N_15092,N_11630,N_13596);
and U15093 (N_15093,N_12140,N_11084);
nand U15094 (N_15094,N_14635,N_10947);
xnor U15095 (N_15095,N_11596,N_13440);
nor U15096 (N_15096,N_10834,N_14525);
xor U15097 (N_15097,N_10524,N_14529);
and U15098 (N_15098,N_11187,N_10236);
and U15099 (N_15099,N_11989,N_13151);
nand U15100 (N_15100,N_10176,N_12899);
xor U15101 (N_15101,N_12465,N_14550);
xor U15102 (N_15102,N_11767,N_10681);
nand U15103 (N_15103,N_10594,N_10714);
nand U15104 (N_15104,N_10755,N_13205);
or U15105 (N_15105,N_13380,N_10806);
or U15106 (N_15106,N_10826,N_11326);
xor U15107 (N_15107,N_13764,N_11258);
nand U15108 (N_15108,N_12965,N_13295);
and U15109 (N_15109,N_11148,N_14683);
or U15110 (N_15110,N_10884,N_13506);
and U15111 (N_15111,N_11141,N_10960);
xnor U15112 (N_15112,N_12177,N_11789);
or U15113 (N_15113,N_10741,N_12100);
xor U15114 (N_15114,N_11431,N_10590);
xnor U15115 (N_15115,N_13746,N_12770);
or U15116 (N_15116,N_13732,N_14706);
nor U15117 (N_15117,N_13886,N_14284);
and U15118 (N_15118,N_14911,N_14809);
nor U15119 (N_15119,N_10076,N_12889);
or U15120 (N_15120,N_11041,N_12616);
nand U15121 (N_15121,N_10893,N_12032);
nor U15122 (N_15122,N_13312,N_10397);
or U15123 (N_15123,N_10090,N_10175);
xnor U15124 (N_15124,N_12263,N_13969);
nand U15125 (N_15125,N_13139,N_10083);
nor U15126 (N_15126,N_11039,N_14742);
and U15127 (N_15127,N_11451,N_11866);
or U15128 (N_15128,N_10359,N_13722);
xnor U15129 (N_15129,N_10005,N_12783);
or U15130 (N_15130,N_11388,N_12797);
or U15131 (N_15131,N_14205,N_10668);
nand U15132 (N_15132,N_10670,N_10293);
or U15133 (N_15133,N_14507,N_13426);
and U15134 (N_15134,N_10173,N_10487);
nand U15135 (N_15135,N_12217,N_10892);
xnor U15136 (N_15136,N_11085,N_11639);
and U15137 (N_15137,N_10829,N_10046);
nand U15138 (N_15138,N_13237,N_13171);
nand U15139 (N_15139,N_10658,N_11822);
or U15140 (N_15140,N_13985,N_13190);
xnor U15141 (N_15141,N_14700,N_11711);
xnor U15142 (N_15142,N_14487,N_13065);
and U15143 (N_15143,N_14342,N_11233);
nor U15144 (N_15144,N_13707,N_11819);
or U15145 (N_15145,N_11648,N_13518);
or U15146 (N_15146,N_14548,N_12677);
nand U15147 (N_15147,N_10978,N_14352);
nand U15148 (N_15148,N_12084,N_13832);
and U15149 (N_15149,N_12861,N_12966);
xnor U15150 (N_15150,N_12578,N_13257);
nor U15151 (N_15151,N_14590,N_12820);
xor U15152 (N_15152,N_10125,N_10995);
and U15153 (N_15153,N_12817,N_10848);
or U15154 (N_15154,N_14308,N_14778);
or U15155 (N_15155,N_11474,N_11908);
nor U15156 (N_15156,N_13197,N_13284);
nand U15157 (N_15157,N_13821,N_10466);
nor U15158 (N_15158,N_10925,N_14844);
xnor U15159 (N_15159,N_11160,N_14572);
nor U15160 (N_15160,N_13322,N_14828);
or U15161 (N_15161,N_11192,N_14969);
nand U15162 (N_15162,N_12553,N_14830);
nand U15163 (N_15163,N_13807,N_11601);
or U15164 (N_15164,N_10011,N_13650);
nor U15165 (N_15165,N_11808,N_14769);
or U15166 (N_15166,N_12653,N_10503);
and U15167 (N_15167,N_12893,N_13855);
nand U15168 (N_15168,N_11353,N_10457);
and U15169 (N_15169,N_12980,N_13641);
nor U15170 (N_15170,N_13261,N_11533);
nor U15171 (N_15171,N_12467,N_11123);
xnor U15172 (N_15172,N_11965,N_12655);
nand U15173 (N_15173,N_14142,N_12179);
nand U15174 (N_15174,N_10423,N_13781);
or U15175 (N_15175,N_12088,N_13753);
or U15176 (N_15176,N_12365,N_11944);
or U15177 (N_15177,N_10991,N_13054);
nor U15178 (N_15178,N_13666,N_14362);
nand U15179 (N_15179,N_10786,N_10760);
nand U15180 (N_15180,N_11247,N_10445);
and U15181 (N_15181,N_10817,N_12373);
and U15182 (N_15182,N_14884,N_10534);
or U15183 (N_15183,N_14743,N_13763);
nand U15184 (N_15184,N_12998,N_13852);
xnor U15185 (N_15185,N_12552,N_10531);
nand U15186 (N_15186,N_11592,N_10544);
and U15187 (N_15187,N_14392,N_14758);
nor U15188 (N_15188,N_10586,N_10002);
nor U15189 (N_15189,N_11277,N_12443);
nand U15190 (N_15190,N_10429,N_13510);
nor U15191 (N_15191,N_10945,N_14685);
xor U15192 (N_15192,N_14629,N_12441);
nand U15193 (N_15193,N_11723,N_13498);
or U15194 (N_15194,N_10879,N_14597);
or U15195 (N_15195,N_10351,N_14804);
and U15196 (N_15196,N_13774,N_13696);
nand U15197 (N_15197,N_10142,N_13957);
and U15198 (N_15198,N_10229,N_11065);
nor U15199 (N_15199,N_10881,N_11453);
and U15200 (N_15200,N_12095,N_10761);
xor U15201 (N_15201,N_12057,N_12375);
nor U15202 (N_15202,N_14756,N_11858);
and U15203 (N_15203,N_12951,N_12496);
nand U15204 (N_15204,N_12534,N_10775);
or U15205 (N_15205,N_10491,N_13108);
nand U15206 (N_15206,N_10562,N_11086);
and U15207 (N_15207,N_12781,N_10154);
xor U15208 (N_15208,N_13912,N_13663);
nand U15209 (N_15209,N_11917,N_10456);
nor U15210 (N_15210,N_11645,N_11319);
nor U15211 (N_15211,N_10204,N_12413);
or U15212 (N_15212,N_14319,N_12658);
and U15213 (N_15213,N_11028,N_13509);
or U15214 (N_15214,N_12922,N_10105);
or U15215 (N_15215,N_10630,N_10227);
or U15216 (N_15216,N_10550,N_13210);
nor U15217 (N_15217,N_13093,N_13994);
xor U15218 (N_15218,N_14945,N_12792);
nor U15219 (N_15219,N_10546,N_13928);
or U15220 (N_15220,N_14455,N_10097);
and U15221 (N_15221,N_11118,N_14510);
nor U15222 (N_15222,N_13405,N_11887);
nor U15223 (N_15223,N_11752,N_12320);
xor U15224 (N_15224,N_10944,N_12941);
nor U15225 (N_15225,N_14164,N_13789);
nor U15226 (N_15226,N_13822,N_13038);
or U15227 (N_15227,N_12767,N_11071);
or U15228 (N_15228,N_12041,N_10948);
or U15229 (N_15229,N_13921,N_13505);
nand U15230 (N_15230,N_14094,N_14595);
nand U15231 (N_15231,N_14009,N_12937);
nor U15232 (N_15232,N_14070,N_10941);
nor U15233 (N_15233,N_10690,N_12045);
or U15234 (N_15234,N_11070,N_10067);
or U15235 (N_15235,N_12707,N_13291);
nor U15236 (N_15236,N_10647,N_12457);
or U15237 (N_15237,N_13450,N_14732);
or U15238 (N_15238,N_12419,N_13477);
xor U15239 (N_15239,N_11305,N_13591);
nand U15240 (N_15240,N_12948,N_12935);
xor U15241 (N_15241,N_12393,N_12777);
nand U15242 (N_15242,N_12485,N_12909);
nand U15243 (N_15243,N_12785,N_13189);
and U15244 (N_15244,N_11392,N_11484);
nand U15245 (N_15245,N_11881,N_13032);
and U15246 (N_15246,N_13468,N_13338);
xnor U15247 (N_15247,N_13608,N_12016);
and U15248 (N_15248,N_12651,N_11582);
nor U15249 (N_15249,N_12765,N_10009);
nor U15250 (N_15250,N_12348,N_13619);
nor U15251 (N_15251,N_12122,N_11417);
or U15252 (N_15252,N_11838,N_11750);
and U15253 (N_15253,N_13803,N_10752);
nand U15254 (N_15254,N_13164,N_12096);
and U15255 (N_15255,N_14903,N_12059);
and U15256 (N_15256,N_10923,N_10910);
xor U15257 (N_15257,N_12141,N_10527);
or U15258 (N_15258,N_11543,N_10132);
nand U15259 (N_15259,N_11244,N_13611);
and U15260 (N_15260,N_14617,N_12382);
or U15261 (N_15261,N_13947,N_13441);
nand U15262 (N_15262,N_10171,N_13422);
and U15263 (N_15263,N_13758,N_13528);
or U15264 (N_15264,N_10643,N_10042);
and U15265 (N_15265,N_10363,N_11505);
nor U15266 (N_15266,N_14602,N_13290);
nand U15267 (N_15267,N_12281,N_10857);
and U15268 (N_15268,N_14366,N_13337);
nand U15269 (N_15269,N_12440,N_11884);
and U15270 (N_15270,N_12157,N_14310);
xor U15271 (N_15271,N_12241,N_14148);
and U15272 (N_15272,N_14027,N_14393);
xor U15273 (N_15273,N_13165,N_11737);
xor U15274 (N_15274,N_11130,N_11446);
or U15275 (N_15275,N_14435,N_11285);
xor U15276 (N_15276,N_10169,N_14011);
nand U15277 (N_15277,N_12302,N_13709);
or U15278 (N_15278,N_13278,N_12019);
nor U15279 (N_15279,N_11501,N_13553);
and U15280 (N_15280,N_11355,N_10867);
and U15281 (N_15281,N_11939,N_10819);
or U15282 (N_15282,N_10207,N_12407);
xnor U15283 (N_15283,N_11536,N_10949);
nand U15284 (N_15284,N_13143,N_12492);
or U15285 (N_15285,N_14569,N_11865);
and U15286 (N_15286,N_10688,N_11310);
xor U15287 (N_15287,N_11846,N_13817);
nand U15288 (N_15288,N_10577,N_13315);
nand U15289 (N_15289,N_12869,N_10460);
xor U15290 (N_15290,N_14309,N_10767);
and U15291 (N_15291,N_14662,N_13386);
and U15292 (N_15292,N_11853,N_13979);
and U15293 (N_15293,N_11557,N_10386);
and U15294 (N_15294,N_11573,N_11801);
or U15295 (N_15295,N_13632,N_13540);
nand U15296 (N_15296,N_11807,N_12018);
or U15297 (N_15297,N_14212,N_14503);
xor U15298 (N_15298,N_14796,N_13909);
or U15299 (N_15299,N_10231,N_13798);
xnor U15300 (N_15300,N_11667,N_13705);
nor U15301 (N_15301,N_10324,N_10876);
nor U15302 (N_15302,N_13159,N_13094);
xor U15303 (N_15303,N_14437,N_13603);
nand U15304 (N_15304,N_13245,N_12895);
and U15305 (N_15305,N_12230,N_13593);
xnor U15306 (N_15306,N_10049,N_12451);
and U15307 (N_15307,N_12597,N_12417);
nor U15308 (N_15308,N_13293,N_11919);
or U15309 (N_15309,N_14047,N_11393);
xnor U15310 (N_15310,N_11239,N_13948);
and U15311 (N_15311,N_13355,N_12652);
nor U15312 (N_15312,N_11229,N_11649);
nor U15313 (N_15313,N_11830,N_14171);
nand U15314 (N_15314,N_12894,N_12181);
nor U15315 (N_15315,N_11428,N_10813);
nand U15316 (N_15316,N_14141,N_10264);
nor U15317 (N_15317,N_12357,N_14052);
nand U15318 (N_15318,N_12113,N_10238);
or U15319 (N_15319,N_14589,N_12974);
or U15320 (N_15320,N_12752,N_10045);
nand U15321 (N_15321,N_14560,N_11781);
or U15322 (N_15322,N_11299,N_10555);
nor U15323 (N_15323,N_10415,N_14851);
xor U15324 (N_15324,N_12943,N_13714);
or U15325 (N_15325,N_11738,N_10917);
nor U15326 (N_15326,N_14820,N_11554);
xor U15327 (N_15327,N_12338,N_10321);
xor U15328 (N_15328,N_13790,N_10058);
nor U15329 (N_15329,N_14591,N_14120);
or U15330 (N_15330,N_13066,N_14961);
nor U15331 (N_15331,N_14311,N_11816);
xor U15332 (N_15332,N_10277,N_11811);
xor U15333 (N_15333,N_12549,N_11054);
nand U15334 (N_15334,N_14644,N_12510);
and U15335 (N_15335,N_13799,N_10106);
xnor U15336 (N_15336,N_10950,N_10612);
or U15337 (N_15337,N_13728,N_11373);
and U15338 (N_15338,N_11741,N_14219);
xnor U15339 (N_15339,N_12730,N_13359);
or U15340 (N_15340,N_14842,N_10652);
xor U15341 (N_15341,N_11223,N_12685);
xnor U15342 (N_15342,N_13004,N_11707);
nor U15343 (N_15343,N_10519,N_14243);
nor U15344 (N_15344,N_12953,N_11414);
and U15345 (N_15345,N_13114,N_11276);
nand U15346 (N_15346,N_10729,N_13367);
xnor U15347 (N_15347,N_11013,N_14029);
and U15348 (N_15348,N_11313,N_14017);
nand U15349 (N_15349,N_11218,N_10254);
and U15350 (N_15350,N_10400,N_13242);
nor U15351 (N_15351,N_11851,N_12545);
or U15352 (N_15352,N_12854,N_14335);
nor U15353 (N_15353,N_12164,N_10913);
nand U15354 (N_15354,N_12316,N_10832);
and U15355 (N_15355,N_14316,N_13267);
nand U15356 (N_15356,N_11742,N_10003);
nor U15357 (N_15357,N_13701,N_14542);
and U15358 (N_15358,N_11524,N_14547);
xor U15359 (N_15359,N_12809,N_12630);
xnor U15360 (N_15360,N_11910,N_12003);
nand U15361 (N_15361,N_10345,N_12372);
or U15362 (N_15362,N_12853,N_12615);
xor U15363 (N_15363,N_11467,N_13453);
nor U15364 (N_15364,N_10816,N_13668);
xor U15365 (N_15365,N_11023,N_12170);
or U15366 (N_15366,N_14937,N_14091);
xnor U15367 (N_15367,N_14175,N_13811);
or U15368 (N_15368,N_14041,N_13212);
and U15369 (N_15369,N_13111,N_11418);
nand U15370 (N_15370,N_10568,N_14901);
or U15371 (N_15371,N_13455,N_14481);
or U15372 (N_15372,N_12619,N_13835);
or U15373 (N_15373,N_10517,N_10294);
or U15374 (N_15374,N_10256,N_11925);
nand U15375 (N_15375,N_12462,N_11762);
xnor U15376 (N_15376,N_10645,N_11976);
and U15377 (N_15377,N_14520,N_11672);
nand U15378 (N_15378,N_13334,N_14860);
nand U15379 (N_15379,N_14735,N_11034);
and U15380 (N_15380,N_13669,N_10967);
or U15381 (N_15381,N_14779,N_10358);
or U15382 (N_15382,N_14643,N_10977);
and U15383 (N_15383,N_13636,N_13025);
xor U15384 (N_15384,N_11796,N_14665);
nor U15385 (N_15385,N_11620,N_12144);
nor U15386 (N_15386,N_12336,N_10897);
xnor U15387 (N_15387,N_14431,N_14653);
or U15388 (N_15388,N_11714,N_10442);
or U15389 (N_15389,N_14677,N_10166);
xnor U15390 (N_15390,N_12605,N_12547);
xor U15391 (N_15391,N_14297,N_10575);
xor U15392 (N_15392,N_14124,N_13160);
and U15393 (N_15393,N_14921,N_14979);
and U15394 (N_15394,N_11547,N_14693);
xnor U15395 (N_15395,N_12400,N_11320);
or U15396 (N_15396,N_10904,N_11687);
xor U15397 (N_15397,N_13610,N_12845);
and U15398 (N_15398,N_10488,N_11942);
and U15399 (N_15399,N_11861,N_14268);
and U15400 (N_15400,N_10150,N_14535);
xor U15401 (N_15401,N_13890,N_10583);
nand U15402 (N_15402,N_11967,N_13706);
nand U15403 (N_15403,N_12565,N_13829);
nand U15404 (N_15404,N_10542,N_12818);
nand U15405 (N_15405,N_13269,N_11539);
or U15406 (N_15406,N_10420,N_11799);
and U15407 (N_15407,N_13604,N_12322);
and U15408 (N_15408,N_12863,N_12712);
nand U15409 (N_15409,N_12406,N_10489);
nor U15410 (N_15410,N_10102,N_10730);
or U15411 (N_15411,N_10720,N_11692);
and U15412 (N_15412,N_11528,N_12643);
and U15413 (N_15413,N_11981,N_11608);
nor U15414 (N_15414,N_12906,N_11551);
nor U15415 (N_15415,N_13460,N_10984);
nand U15416 (N_15416,N_11295,N_10168);
nor U15417 (N_15417,N_10452,N_10669);
and U15418 (N_15418,N_11609,N_12819);
xor U15419 (N_15419,N_11765,N_11008);
or U15420 (N_15420,N_10877,N_13230);
xor U15421 (N_15421,N_12986,N_14391);
nor U15422 (N_15422,N_13949,N_13439);
nor U15423 (N_15423,N_12060,N_13225);
or U15424 (N_15424,N_11088,N_10538);
or U15425 (N_15425,N_14600,N_12624);
nor U15426 (N_15426,N_12370,N_13067);
xnor U15427 (N_15427,N_13894,N_10287);
and U15428 (N_15428,N_14050,N_13218);
xnor U15429 (N_15429,N_10258,N_11659);
nor U15430 (N_15430,N_13856,N_11012);
or U15431 (N_15431,N_10056,N_13578);
and U15432 (N_15432,N_14849,N_11104);
nor U15433 (N_15433,N_12275,N_10261);
or U15434 (N_15434,N_12970,N_11507);
nor U15435 (N_15435,N_13953,N_10290);
nor U15436 (N_15436,N_14870,N_11232);
nand U15437 (N_15437,N_11751,N_13087);
and U15438 (N_15438,N_12146,N_13531);
nor U15439 (N_15439,N_12644,N_14229);
and U15440 (N_15440,N_11045,N_13466);
or U15441 (N_15441,N_12904,N_14028);
nand U15442 (N_15442,N_13541,N_10980);
and U15443 (N_15443,N_12416,N_14610);
and U15444 (N_15444,N_11756,N_13676);
xor U15445 (N_15445,N_12627,N_11931);
xor U15446 (N_15446,N_13292,N_12232);
nand U15447 (N_15447,N_14014,N_10387);
and U15448 (N_15448,N_11905,N_14003);
nand U15449 (N_15449,N_11203,N_10717);
nor U15450 (N_15450,N_14493,N_12831);
or U15451 (N_15451,N_11384,N_11671);
nand U15452 (N_15452,N_10776,N_13156);
nand U15453 (N_15453,N_10121,N_10123);
or U15454 (N_15454,N_11768,N_12234);
and U15455 (N_15455,N_12764,N_12477);
xor U15456 (N_15456,N_12721,N_13998);
nor U15457 (N_15457,N_10447,N_10651);
xnor U15458 (N_15458,N_11934,N_11760);
or U15459 (N_15459,N_10522,N_14815);
or U15460 (N_15460,N_11732,N_14876);
or U15461 (N_15461,N_14526,N_13661);
or U15462 (N_15462,N_11613,N_11496);
nor U15463 (N_15463,N_11426,N_14523);
and U15464 (N_15464,N_13830,N_13018);
and U15465 (N_15465,N_13582,N_12706);
and U15466 (N_15466,N_10026,N_11912);
nor U15467 (N_15467,N_12648,N_14954);
and U15468 (N_15468,N_11726,N_11537);
xnor U15469 (N_15469,N_13936,N_13741);
or U15470 (N_15470,N_14775,N_10312);
or U15471 (N_15471,N_13298,N_10780);
nand U15472 (N_15472,N_12086,N_12256);
or U15473 (N_15473,N_12504,N_11398);
xnor U15474 (N_15474,N_10288,N_13394);
or U15475 (N_15475,N_11655,N_12608);
nand U15476 (N_15476,N_14465,N_11334);
nand U15477 (N_15477,N_12229,N_13778);
and U15478 (N_15478,N_10310,N_12881);
nand U15479 (N_15479,N_12436,N_13609);
or U15480 (N_15480,N_11993,N_14462);
nand U15481 (N_15481,N_11302,N_14084);
nor U15482 (N_15482,N_10769,N_14430);
nand U15483 (N_15483,N_14150,N_12471);
xnor U15484 (N_15484,N_14934,N_14145);
nor U15485 (N_15485,N_13050,N_14755);
nor U15486 (N_15486,N_12246,N_11587);
or U15487 (N_15487,N_12249,N_14428);
xor U15488 (N_15488,N_11217,N_12154);
and U15489 (N_15489,N_10909,N_12053);
nor U15490 (N_15490,N_12657,N_11863);
or U15491 (N_15491,N_12807,N_14917);
xnor U15492 (N_15492,N_13929,N_14146);
nand U15493 (N_15493,N_10554,N_11055);
or U15494 (N_15494,N_10887,N_11440);
nand U15495 (N_15495,N_13028,N_14261);
or U15496 (N_15496,N_12046,N_12039);
xor U15497 (N_15497,N_12927,N_12991);
and U15498 (N_15498,N_12388,N_13224);
nor U15499 (N_15499,N_14461,N_14555);
nor U15500 (N_15500,N_11325,N_11403);
and U15501 (N_15501,N_13715,N_12544);
xor U15502 (N_15502,N_10833,N_10269);
nor U15503 (N_15503,N_12642,N_10308);
and U15504 (N_15504,N_12033,N_13991);
and U15505 (N_15505,N_11840,N_14867);
nor U15506 (N_15506,N_10214,N_13074);
nor U15507 (N_15507,N_12508,N_10621);
or U15508 (N_15508,N_12579,N_13417);
nor U15509 (N_15509,N_12743,N_10565);
and U15510 (N_15510,N_10147,N_10140);
xor U15511 (N_15511,N_10676,N_14208);
and U15512 (N_15512,N_11698,N_14875);
or U15513 (N_15513,N_11643,N_13071);
or U15514 (N_15514,N_14115,N_13524);
nor U15515 (N_15515,N_13956,N_14689);
xnor U15516 (N_15516,N_14165,N_14826);
nand U15517 (N_15517,N_11832,N_13571);
or U15518 (N_15518,N_12649,N_10533);
or U15519 (N_15519,N_14398,N_11745);
nor U15520 (N_15520,N_14975,N_12097);
xnor U15521 (N_15521,N_10915,N_12360);
xnor U15522 (N_15522,N_11438,N_14187);
and U15523 (N_15523,N_10186,N_12833);
xnor U15524 (N_15524,N_11590,N_11270);
and U15525 (N_15525,N_11996,N_10854);
and U15526 (N_15526,N_10161,N_14127);
xor U15527 (N_15527,N_13679,N_14783);
or U15528 (N_15528,N_13321,N_12815);
or U15529 (N_15529,N_14587,N_10235);
or U15530 (N_15530,N_14885,N_11198);
xnor U15531 (N_15531,N_12222,N_10475);
xnor U15532 (N_15532,N_13934,N_13736);
nor U15533 (N_15533,N_14456,N_14962);
and U15534 (N_15534,N_11694,N_13503);
nand U15535 (N_15535,N_14073,N_14519);
or U15536 (N_15536,N_10362,N_11769);
and U15537 (N_15537,N_14822,N_13565);
nand U15538 (N_15538,N_11242,N_14236);
and U15539 (N_15539,N_13459,N_10641);
nor U15540 (N_15540,N_13195,N_10044);
and U15541 (N_15541,N_13031,N_12150);
and U15542 (N_15542,N_14785,N_13299);
nor U15543 (N_15543,N_13389,N_10886);
nand U15544 (N_15544,N_11140,N_13564);
and U15545 (N_15545,N_10632,N_13688);
xor U15546 (N_15546,N_12747,N_10458);
xor U15547 (N_15547,N_10032,N_13390);
nor U15548 (N_15548,N_10799,N_12623);
nand U15549 (N_15549,N_13738,N_14479);
nand U15550 (N_15550,N_12802,N_11346);
nor U15551 (N_15551,N_11317,N_11240);
xnor U15552 (N_15552,N_12589,N_14898);
and U15553 (N_15553,N_13384,N_13136);
or U15554 (N_15554,N_10112,N_11735);
nor U15555 (N_15555,N_10388,N_12933);
nand U15556 (N_15556,N_10289,N_10642);
and U15557 (N_15557,N_10124,N_12453);
xor U15558 (N_15558,N_12849,N_14172);
nand U15559 (N_15559,N_11015,N_14544);
and U15560 (N_15560,N_11206,N_11509);
nor U15561 (N_15561,N_14744,N_14304);
nor U15562 (N_15562,N_14757,N_10136);
or U15563 (N_15563,N_11215,N_13347);
xnor U15564 (N_15564,N_10329,N_12358);
or U15565 (N_15565,N_10649,N_12618);
or U15566 (N_15566,N_10841,N_14388);
nor U15567 (N_15567,N_10571,N_10367);
and U15568 (N_15568,N_10405,N_11518);
and U15569 (N_15569,N_14337,N_12840);
and U15570 (N_15570,N_10859,N_13145);
and U15571 (N_15571,N_11169,N_12020);
and U15572 (N_15572,N_10956,N_11115);
xor U15573 (N_15573,N_13249,N_10201);
nand U15574 (N_15574,N_10240,N_11162);
nor U15575 (N_15575,N_10153,N_10521);
xnor U15576 (N_15576,N_12221,N_10114);
xnor U15577 (N_15577,N_11684,N_14372);
nand U15578 (N_15578,N_10812,N_13134);
xor U15579 (N_15579,N_13276,N_12520);
nand U15580 (N_15580,N_12541,N_12334);
and U15581 (N_15581,N_11152,N_13056);
or U15582 (N_15582,N_14241,N_13035);
or U15583 (N_15583,N_13351,N_14320);
nand U15584 (N_15584,N_14666,N_10520);
and U15585 (N_15585,N_10932,N_13131);
nand U15586 (N_15586,N_12201,N_13326);
xnor U15587 (N_15587,N_10566,N_10530);
and U15588 (N_15588,N_10273,N_10041);
and U15589 (N_15589,N_13533,N_13393);
nand U15590 (N_15590,N_13470,N_13857);
or U15591 (N_15591,N_12717,N_12784);
and U15592 (N_15592,N_13946,N_14982);
nand U15593 (N_15593,N_14104,N_11214);
nand U15594 (N_15594,N_13493,N_12913);
xor U15595 (N_15595,N_14797,N_10198);
nand U15596 (N_15596,N_13353,N_14043);
nand U15597 (N_15597,N_12077,N_13375);
or U15598 (N_15598,N_11076,N_10536);
or U15599 (N_15599,N_10424,N_11686);
nand U15600 (N_15600,N_10875,N_13834);
nand U15601 (N_15601,N_12128,N_12061);
or U15602 (N_15602,N_10784,N_12566);
or U15603 (N_15603,N_12573,N_14209);
nand U15604 (N_15604,N_11455,N_13487);
and U15605 (N_15605,N_12464,N_14607);
xor U15606 (N_15606,N_10305,N_10485);
xor U15607 (N_15607,N_13550,N_13319);
nor U15608 (N_15608,N_14577,N_12110);
or U15609 (N_15609,N_10148,N_12257);
nand U15610 (N_15610,N_11847,N_13323);
xor U15611 (N_15611,N_11108,N_13984);
and U15612 (N_15612,N_10771,N_11193);
xnor U15613 (N_15613,N_14579,N_12040);
xnor U15614 (N_15614,N_14782,N_12524);
xor U15615 (N_15615,N_12826,N_12696);
xor U15616 (N_15616,N_11183,N_13902);
nor U15617 (N_15617,N_12151,N_10844);
xnor U15618 (N_15618,N_11143,N_11977);
nand U15619 (N_15619,N_10557,N_12447);
nand U15620 (N_15620,N_12848,N_11042);
xor U15621 (N_15621,N_11324,N_11158);
xnor U15622 (N_15622,N_13447,N_13708);
xor U15623 (N_15623,N_14925,N_12847);
xor U15624 (N_15624,N_11379,N_11443);
and U15625 (N_15625,N_13495,N_11932);
and U15626 (N_15626,N_13140,N_13235);
nand U15627 (N_15627,N_10985,N_10347);
or U15628 (N_15628,N_10545,N_14847);
or U15629 (N_15629,N_13486,N_11771);
and U15630 (N_15630,N_11298,N_10732);
xnor U15631 (N_15631,N_11599,N_11424);
xor U15632 (N_15632,N_13827,N_14825);
and U15633 (N_15633,N_11534,N_13568);
or U15634 (N_15634,N_12228,N_12478);
or U15635 (N_15635,N_14508,N_14791);
or U15636 (N_15636,N_13154,N_13277);
nand U15637 (N_15637,N_14259,N_13011);
and U15638 (N_15638,N_12102,N_12507);
nor U15639 (N_15639,N_13120,N_10507);
nand U15640 (N_15640,N_14060,N_13200);
nor U15641 (N_15641,N_11168,N_13760);
or U15642 (N_15642,N_14298,N_14680);
nor U15643 (N_15643,N_14896,N_14609);
nand U15644 (N_15644,N_11382,N_14696);
xor U15645 (N_15645,N_10976,N_11363);
xnor U15646 (N_15646,N_11278,N_13499);
xor U15647 (N_15647,N_12920,N_13395);
nand U15648 (N_15648,N_13874,N_11960);
or U15649 (N_15649,N_12694,N_12202);
and U15650 (N_15650,N_14562,N_11958);
or U15651 (N_15651,N_11571,N_14299);
nor U15652 (N_15652,N_11647,N_11150);
xnor U15653 (N_15653,N_13027,N_11813);
or U15654 (N_15654,N_10131,N_13192);
and U15655 (N_15655,N_14275,N_10212);
nand U15656 (N_15656,N_14703,N_10682);
or U15657 (N_15657,N_14927,N_14657);
nor U15658 (N_15658,N_14088,N_11920);
or U15659 (N_15659,N_11935,N_13718);
xor U15660 (N_15660,N_14394,N_12183);
xnor U15661 (N_15661,N_11241,N_10737);
nand U15662 (N_15662,N_10074,N_10143);
or U15663 (N_15663,N_10080,N_10523);
and U15664 (N_15664,N_13115,N_10831);
nand U15665 (N_15665,N_11564,N_12917);
or U15666 (N_15666,N_14090,N_12647);
and U15667 (N_15667,N_12514,N_14929);
and U15668 (N_15668,N_14225,N_14707);
and U15669 (N_15669,N_14850,N_10390);
nand U15670 (N_15670,N_10811,N_12168);
or U15671 (N_15671,N_11867,N_14664);
nor U15672 (N_15672,N_10818,N_11998);
or U15673 (N_15673,N_13881,N_10033);
nand U15674 (N_15674,N_14904,N_11730);
xor U15675 (N_15675,N_12437,N_13808);
or U15676 (N_15676,N_12127,N_14367);
xor U15677 (N_15677,N_14458,N_14232);
nor U15678 (N_15678,N_12445,N_11089);
and U15679 (N_15679,N_13329,N_12198);
nand U15680 (N_15680,N_11641,N_12130);
nor U15681 (N_15681,N_11629,N_14192);
xnor U15682 (N_15682,N_12460,N_13244);
or U15683 (N_15683,N_11480,N_10281);
and U15684 (N_15684,N_12409,N_11352);
nor U15685 (N_15685,N_10407,N_14681);
nand U15686 (N_15686,N_14258,N_12292);
xor U15687 (N_15687,N_10990,N_10317);
or U15688 (N_15688,N_11350,N_12570);
nand U15689 (N_15689,N_11117,N_11555);
nor U15690 (N_15690,N_13449,N_13859);
xor U15691 (N_15691,N_11764,N_14780);
xnor U15692 (N_15692,N_11784,N_13916);
nand U15693 (N_15693,N_10419,N_12650);
nor U15694 (N_15694,N_13411,N_13254);
nor U15695 (N_15695,N_11237,N_11900);
nor U15696 (N_15696,N_11275,N_13026);
nor U15697 (N_15697,N_14000,N_14266);
xnor U15698 (N_15698,N_11415,N_11461);
or U15699 (N_15699,N_10861,N_12213);
and U15700 (N_15700,N_11876,N_14245);
and U15701 (N_15701,N_13461,N_12262);
or U15702 (N_15702,N_14618,N_13073);
xor U15703 (N_15703,N_13838,N_13365);
xnor U15704 (N_15704,N_10210,N_13231);
nor U15705 (N_15705,N_10380,N_10560);
xnor U15706 (N_15706,N_13118,N_14425);
xor U15707 (N_15707,N_14036,N_14346);
or U15708 (N_15708,N_11212,N_12219);
nand U15709 (N_15709,N_10582,N_10241);
nor U15710 (N_15710,N_12352,N_10278);
or U15711 (N_15711,N_12924,N_14322);
and U15712 (N_15712,N_11857,N_14719);
and U15713 (N_15713,N_14906,N_10872);
nand U15714 (N_15714,N_12092,N_10246);
and U15715 (N_15715,N_11653,N_14692);
xor U15716 (N_15716,N_13907,N_10567);
and U15717 (N_15717,N_10398,N_10216);
or U15718 (N_15718,N_14810,N_14857);
xor U15719 (N_15719,N_12969,N_13711);
or U15720 (N_15720,N_13085,N_13864);
nor U15721 (N_15721,N_11109,N_10408);
nand U15722 (N_15722,N_12311,N_12719);
and U15723 (N_15723,N_10493,N_10993);
and U15724 (N_15724,N_13335,N_11387);
nand U15725 (N_15725,N_14816,N_12024);
nor U15726 (N_15726,N_12601,N_12192);
nor U15727 (N_15727,N_10078,N_12429);
or U15728 (N_15728,N_13640,N_10332);
and U15729 (N_15729,N_10842,N_11003);
or U15730 (N_15730,N_10624,N_13240);
xor U15731 (N_15731,N_11713,N_13465);
nor U15732 (N_15732,N_14512,N_12121);
nand U15733 (N_15733,N_10878,N_14784);
nand U15734 (N_15734,N_13662,N_13173);
or U15735 (N_15735,N_10973,N_14712);
and U15736 (N_15736,N_14673,N_12962);
nand U15737 (N_15737,N_13656,N_14058);
and U15738 (N_15738,N_13622,N_10064);
nand U15739 (N_15739,N_12314,N_11591);
xnor U15740 (N_15740,N_10365,N_13950);
nor U15741 (N_15741,N_14289,N_14698);
nand U15742 (N_15742,N_10709,N_14423);
and U15743 (N_15743,N_13316,N_13364);
nand U15744 (N_15744,N_11002,N_11422);
xor U15745 (N_15745,N_13016,N_10890);
nand U15746 (N_15746,N_11378,N_10862);
xor U15747 (N_15747,N_13939,N_10942);
nand U15748 (N_15748,N_11744,N_13587);
or U15749 (N_15749,N_10292,N_10639);
and U15750 (N_15750,N_11116,N_12581);
nor U15751 (N_15751,N_11222,N_10417);
and U15752 (N_15752,N_10025,N_12963);
nor U15753 (N_15753,N_12759,N_13635);
and U15754 (N_15754,N_12979,N_11262);
and U15755 (N_15755,N_13340,N_12633);
nand U15756 (N_15756,N_11069,N_11204);
and U15757 (N_15757,N_13148,N_14651);
nor U15758 (N_15758,N_14099,N_13552);
nor U15759 (N_15759,N_10039,N_14747);
nor U15760 (N_15760,N_12555,N_10206);
nand U15761 (N_15761,N_12226,N_11151);
and U15762 (N_15762,N_14966,N_14184);
nor U15763 (N_15763,N_14216,N_12775);
or U15764 (N_15764,N_12683,N_11017);
nand U15765 (N_15765,N_14965,N_11487);
nand U15766 (N_15766,N_11062,N_11068);
or U15767 (N_15767,N_10659,N_13017);
or U15768 (N_15768,N_14957,N_12596);
xnor U15769 (N_15769,N_11777,N_12461);
xor U15770 (N_15770,N_11036,N_10739);
or U15771 (N_15771,N_13402,N_14524);
xnor U15772 (N_15772,N_13201,N_13986);
and U15773 (N_15773,N_13421,N_11096);
or U15774 (N_15774,N_11043,N_12082);
and U15775 (N_15775,N_11618,N_13586);
xnor U15776 (N_15776,N_14718,N_13149);
nand U15777 (N_15777,N_10103,N_13793);
nor U15778 (N_15778,N_12813,N_13861);
nand U15779 (N_15779,N_14194,N_13058);
nor U15780 (N_15780,N_14095,N_11673);
nor U15781 (N_15781,N_14688,N_10774);
or U15782 (N_15782,N_13842,N_12295);
nand U15783 (N_15783,N_10779,N_12982);
or U15784 (N_15784,N_13845,N_12528);
nor U15785 (N_15785,N_13869,N_10971);
and U15786 (N_15786,N_11485,N_13762);
nor U15787 (N_15787,N_14072,N_14994);
and U15788 (N_15788,N_10803,N_13501);
nand U15789 (N_15789,N_10181,N_14402);
nor U15790 (N_15790,N_13490,N_11025);
nor U15791 (N_15791,N_11472,N_14573);
nand U15792 (N_15792,N_13141,N_14533);
or U15793 (N_15793,N_11250,N_14470);
and U15794 (N_15794,N_12031,N_13765);
or U15795 (N_15795,N_11888,N_10694);
and U15796 (N_15796,N_11314,N_14601);
and U15797 (N_15797,N_13301,N_10071);
nand U15798 (N_15798,N_10836,N_12816);
nand U15799 (N_15799,N_14663,N_13860);
xnor U15800 (N_15800,N_12007,N_12286);
xnor U15801 (N_15801,N_10128,N_14494);
or U15802 (N_15802,N_10242,N_13314);
or U15803 (N_15803,N_10605,N_12328);
or U15804 (N_15804,N_12656,N_14615);
nor U15805 (N_15805,N_14155,N_11891);
nor U15806 (N_15806,N_14789,N_12108);
and U15807 (N_15807,N_11770,N_13853);
and U15808 (N_15808,N_10558,N_14326);
xor U15809 (N_15809,N_10706,N_12563);
and U15810 (N_15810,N_14119,N_10448);
nand U15811 (N_15811,N_13188,N_10922);
and U15812 (N_15812,N_11909,N_13502);
nor U15813 (N_15813,N_12109,N_12498);
xnor U15814 (N_15814,N_13489,N_13229);
or U15815 (N_15815,N_12794,N_10361);
nor U15816 (N_15816,N_12810,N_11594);
xor U15817 (N_15817,N_14946,N_14034);
or U15818 (N_15818,N_12855,N_11962);
xor U15819 (N_15819,N_13818,N_10552);
nand U15820 (N_15820,N_10664,N_13534);
nand U15821 (N_15821,N_10072,N_13125);
or U15822 (N_15822,N_14650,N_13922);
nand U15823 (N_15823,N_10611,N_10034);
or U15824 (N_15824,N_11127,N_14625);
or U15825 (N_15825,N_13788,N_11282);
and U15826 (N_15826,N_14988,N_13751);
nand U15827 (N_15827,N_10268,N_14720);
nand U15828 (N_15828,N_12587,N_12766);
nand U15829 (N_15829,N_10030,N_10335);
and U15830 (N_15830,N_10959,N_12125);
xnor U15831 (N_15831,N_11430,N_10412);
xor U15832 (N_15832,N_11005,N_13216);
and U15833 (N_15833,N_12004,N_13147);
and U15834 (N_15834,N_11105,N_13471);
xor U15835 (N_15835,N_12635,N_12945);
xnor U15836 (N_15836,N_12558,N_12512);
or U15837 (N_15837,N_11227,N_14353);
and U15838 (N_15838,N_14158,N_12483);
and U15839 (N_15839,N_12174,N_12376);
and U15840 (N_15840,N_13246,N_10433);
or U15841 (N_15841,N_14619,N_11356);
or U15842 (N_15842,N_13575,N_12148);
nor U15843 (N_15843,N_11914,N_10193);
or U15844 (N_15844,N_12364,N_10855);
nand U15845 (N_15845,N_11907,N_13002);
and U15846 (N_15846,N_12708,N_13937);
nand U15847 (N_15847,N_12463,N_10213);
xnor U15848 (N_15848,N_13423,N_12374);
xnor U15849 (N_15849,N_12715,N_13360);
nand U15850 (N_15850,N_14262,N_13629);
or U15851 (N_15851,N_12890,N_13884);
xor U15852 (N_15852,N_13012,N_10661);
or U15853 (N_15853,N_12636,N_10969);
nand U15854 (N_15854,N_10916,N_14515);
and U15855 (N_15855,N_14325,N_14549);
or U15856 (N_15856,N_13882,N_12442);
xor U15857 (N_15857,N_14675,N_13265);
nand U15858 (N_15858,N_13126,N_13475);
nand U15859 (N_15859,N_10699,N_13734);
nand U15860 (N_15860,N_14705,N_11690);
or U15861 (N_15861,N_12359,N_11883);
xnor U15862 (N_15862,N_13849,N_10253);
and U15863 (N_15863,N_14837,N_12337);
xnor U15864 (N_15864,N_11292,N_13387);
nand U15865 (N_15865,N_13841,N_13088);
or U15866 (N_15866,N_12333,N_14998);
nor U15867 (N_15867,N_13651,N_13770);
xnor U15868 (N_15868,N_11321,N_11139);
or U15869 (N_15869,N_14476,N_11066);
or U15870 (N_15870,N_11077,N_14217);
nand U15871 (N_15871,N_13454,N_12378);
and U15872 (N_15872,N_12695,N_13976);
xor U15873 (N_15873,N_13698,N_11007);
xnor U15874 (N_15874,N_11234,N_10497);
nand U15875 (N_15875,N_10736,N_11153);
xor U15876 (N_15876,N_14269,N_10465);
or U15877 (N_15877,N_14713,N_13989);
and U15878 (N_15878,N_12835,N_10768);
nor U15879 (N_15879,N_10928,N_10144);
nor U15880 (N_15880,N_12204,N_12165);
or U15881 (N_15881,N_12868,N_13434);
xnor U15882 (N_15882,N_10087,N_11688);
nor U15883 (N_15883,N_12896,N_12106);
nor U15884 (N_15884,N_10727,N_14963);
nor U15885 (N_15885,N_10529,N_12300);
or U15886 (N_15886,N_13511,N_11231);
and U15887 (N_15887,N_13621,N_14944);
nor U15888 (N_15888,N_10435,N_13076);
nand U15889 (N_15889,N_10471,N_10964);
xor U15890 (N_15890,N_13369,N_13392);
and U15891 (N_15891,N_12509,N_12803);
or U15892 (N_15892,N_11999,N_11580);
xnor U15893 (N_15893,N_12583,N_12131);
xor U15894 (N_15894,N_11155,N_11506);
and U15895 (N_15895,N_11458,N_13382);
nor U15896 (N_15896,N_10099,N_12038);
and U15897 (N_15897,N_12988,N_11380);
nor U15898 (N_15898,N_14583,N_11021);
xor U15899 (N_15899,N_12641,N_10975);
nor U15900 (N_15900,N_13399,N_10498);
and U15901 (N_15901,N_11703,N_10259);
or U15902 (N_15902,N_14471,N_14598);
nand U15903 (N_15903,N_12325,N_11291);
and U15904 (N_15904,N_12119,N_13556);
and U15905 (N_15905,N_13563,N_14883);
or U15906 (N_15906,N_10628,N_13700);
and U15907 (N_15907,N_10540,N_10958);
nand U15908 (N_15908,N_10200,N_12722);
or U15909 (N_15909,N_14191,N_13286);
nand U15910 (N_15910,N_12242,N_14948);
nor U15911 (N_15911,N_11323,N_13530);
and U15912 (N_15912,N_11251,N_14450);
and U15913 (N_15913,N_13878,N_11040);
nand U15914 (N_15914,N_14459,N_12960);
nand U15915 (N_15915,N_14363,N_12836);
xnor U15916 (N_15916,N_12678,N_14136);
and U15917 (N_15917,N_13819,N_12480);
nor U15918 (N_15918,N_11486,N_10219);
nand U15919 (N_15919,N_12446,N_10476);
xnor U15920 (N_15920,N_12540,N_11588);
xor U15921 (N_15921,N_10146,N_14347);
and U15922 (N_15922,N_13920,N_12026);
nor U15923 (N_15923,N_12315,N_14078);
and U15924 (N_15924,N_13693,N_14420);
xnor U15925 (N_15925,N_10589,N_10587);
and U15926 (N_15926,N_13311,N_10888);
and U15927 (N_15927,N_13226,N_14176);
nand U15928 (N_15928,N_12875,N_11558);
and U15929 (N_15929,N_13414,N_12782);
or U15930 (N_15930,N_12897,N_12976);
nor U15931 (N_15931,N_14005,N_11793);
nor U15932 (N_15932,N_12622,N_12698);
nand U15933 (N_15933,N_10745,N_10172);
nand U15934 (N_15934,N_12274,N_10203);
nand U15935 (N_15935,N_10341,N_13252);
xor U15936 (N_15936,N_10244,N_11953);
xnor U15937 (N_15937,N_13796,N_13208);
or U15938 (N_15938,N_11774,N_13597);
xor U15939 (N_15939,N_14731,N_10673);
nor U15940 (N_15940,N_12501,N_11103);
and U15941 (N_15941,N_10883,N_11101);
or U15942 (N_15942,N_14226,N_13469);
xnor U15943 (N_15943,N_14403,N_10701);
nand U15944 (N_15944,N_14126,N_14761);
nor U15945 (N_15945,N_13480,N_11831);
nand U15946 (N_15946,N_13580,N_14286);
xnor U15947 (N_15947,N_12385,N_13342);
or U15948 (N_15948,N_13199,N_14077);
or U15949 (N_15949,N_12700,N_13072);
nand U15950 (N_15950,N_11705,N_11522);
nor U15951 (N_15951,N_14287,N_12871);
or U15952 (N_15952,N_11179,N_10177);
or U15953 (N_15953,N_12529,N_12392);
or U15954 (N_15954,N_14624,N_13452);
and U15955 (N_15955,N_13546,N_10635);
nor U15956 (N_15956,N_12796,N_10982);
or U15957 (N_15957,N_12548,N_14636);
xnor U15958 (N_15958,N_10384,N_14318);
or U15959 (N_15959,N_10392,N_13771);
nor U15960 (N_15960,N_13341,N_11207);
or U15961 (N_15961,N_11182,N_13627);
xor U15962 (N_15962,N_11491,N_13101);
nor U15963 (N_15963,N_10297,N_14485);
or U15964 (N_15964,N_14912,N_13645);
nor U15965 (N_15965,N_12735,N_10657);
nand U15966 (N_15966,N_14632,N_11136);
and U15967 (N_15967,N_10785,N_12438);
or U15968 (N_15968,N_10416,N_13097);
nand U15969 (N_15969,N_14888,N_14025);
nand U15970 (N_15970,N_14278,N_13483);
or U15971 (N_15971,N_14411,N_14446);
nand U15972 (N_15972,N_14853,N_11868);
or U15973 (N_15973,N_10232,N_11757);
or U15974 (N_15974,N_14670,N_12332);
nand U15975 (N_15975,N_13420,N_12617);
and U15976 (N_15976,N_11180,N_12702);
xnor U15977 (N_15977,N_13833,N_11860);
nand U15978 (N_15978,N_11748,N_11340);
and U15979 (N_15979,N_10098,N_10981);
and U15980 (N_15980,N_14652,N_13776);
and U15981 (N_15981,N_10350,N_13307);
nor U15982 (N_15982,N_11376,N_12449);
or U15983 (N_15983,N_12469,N_12245);
nand U15984 (N_15984,N_13581,N_13572);
and U15985 (N_15985,N_10095,N_11681);
xnor U15986 (N_15986,N_11817,N_13997);
xor U15987 (N_15987,N_14385,N_12395);
or U15988 (N_15988,N_14575,N_14559);
nor U15989 (N_15989,N_12162,N_12741);
or U15990 (N_15990,N_11556,N_13983);
nand U15991 (N_15991,N_12877,N_11004);
or U15992 (N_15992,N_13919,N_11272);
and U15993 (N_15993,N_11733,N_12386);
or U15994 (N_15994,N_14737,N_12044);
nand U15995 (N_15995,N_11584,N_10506);
and U15996 (N_15996,N_11095,N_14121);
nor U15997 (N_15997,N_13982,N_13378);
or U15998 (N_15998,N_12898,N_10120);
nand U15999 (N_15999,N_11142,N_14329);
and U16000 (N_16000,N_10414,N_12142);
xor U16001 (N_16001,N_11010,N_14442);
or U16002 (N_16002,N_14408,N_14593);
nor U16003 (N_16003,N_12664,N_10644);
xor U16004 (N_16004,N_12176,N_10743);
nand U16005 (N_16005,N_14214,N_14447);
nor U16006 (N_16006,N_13488,N_14613);
and U16007 (N_16007,N_14818,N_11281);
and U16008 (N_16008,N_12701,N_11172);
or U16009 (N_16009,N_11416,N_13317);
nand U16010 (N_16010,N_11006,N_10697);
nand U16011 (N_16011,N_13409,N_14833);
nand U16012 (N_16012,N_13634,N_13613);
nand U16013 (N_16013,N_14943,N_11951);
nand U16014 (N_16014,N_12123,N_10898);
or U16015 (N_16015,N_12236,N_13313);
or U16016 (N_16016,N_13041,N_10252);
xor U16017 (N_16017,N_12002,N_10631);
xor U16018 (N_16018,N_10048,N_13516);
or U16019 (N_16019,N_14829,N_14736);
nor U16020 (N_16020,N_11146,N_12472);
nor U16021 (N_16021,N_14709,N_12104);
nor U16022 (N_16022,N_12269,N_12037);
xor U16023 (N_16023,N_11330,N_11651);
or U16024 (N_16024,N_13117,N_13992);
and U16025 (N_16025,N_14062,N_13719);
xnor U16026 (N_16026,N_12883,N_11449);
or U16027 (N_16027,N_14467,N_11870);
or U16028 (N_16028,N_12418,N_13900);
xnor U16029 (N_16029,N_10063,N_10082);
and U16030 (N_16030,N_14357,N_14321);
or U16031 (N_16031,N_14019,N_11982);
nand U16032 (N_16032,N_14701,N_12267);
nor U16033 (N_16033,N_13617,N_14405);
or U16034 (N_16034,N_12659,N_12277);
nor U16035 (N_16035,N_12342,N_13304);
nand U16036 (N_16036,N_14371,N_14879);
nand U16037 (N_16037,N_11423,N_14251);
xnor U16038 (N_16038,N_14990,N_14100);
or U16039 (N_16039,N_12139,N_10401);
and U16040 (N_16040,N_13980,N_13828);
nand U16041 (N_16041,N_13464,N_14861);
xor U16042 (N_16042,N_12543,N_13336);
and U16043 (N_16043,N_11997,N_14546);
nand U16044 (N_16044,N_13010,N_11924);
nand U16045 (N_16045,N_13047,N_12614);
nor U16046 (N_16046,N_14383,N_10986);
nor U16047 (N_16047,N_10031,N_10116);
and U16048 (N_16048,N_14033,N_13383);
nor U16049 (N_16049,N_14543,N_10914);
xnor U16050 (N_16050,N_10924,N_14180);
nor U16051 (N_16051,N_11540,N_13373);
or U16052 (N_16052,N_14631,N_14163);
nand U16053 (N_16053,N_13966,N_11181);
xor U16054 (N_16054,N_14203,N_10344);
xor U16055 (N_16055,N_12261,N_11778);
or U16056 (N_16056,N_10225,N_11531);
nand U16057 (N_16057,N_11877,N_11624);
xnor U16058 (N_16058,N_14273,N_14160);
and U16059 (N_16059,N_14586,N_12830);
nor U16060 (N_16060,N_14324,N_12905);
nor U16061 (N_16061,N_12065,N_13648);
nand U16062 (N_16062,N_12194,N_12805);
nor U16063 (N_16063,N_13194,N_11918);
xnor U16064 (N_16064,N_11632,N_12431);
nand U16065 (N_16065,N_11368,N_14928);
xnor U16066 (N_16066,N_10393,N_14117);
nand U16067 (N_16067,N_10505,N_14162);
and U16068 (N_16068,N_13630,N_14397);
nor U16069 (N_16069,N_11057,N_14055);
nor U16070 (N_16070,N_10998,N_13787);
nand U16071 (N_16071,N_14083,N_11826);
and U16072 (N_16072,N_14933,N_13467);
xor U16073 (N_16073,N_12779,N_14862);
or U16074 (N_16074,N_12220,N_13238);
or U16075 (N_16075,N_13723,N_13743);
nor U16076 (N_16076,N_10679,N_11701);
nor U16077 (N_16077,N_13960,N_13812);
xnor U16078 (N_16078,N_12903,N_10163);
or U16079 (N_16079,N_14596,N_10762);
or U16080 (N_16080,N_13491,N_11454);
or U16081 (N_16081,N_10866,N_12070);
nor U16082 (N_16082,N_11676,N_11797);
xor U16083 (N_16083,N_13448,N_14959);
nand U16084 (N_16084,N_11409,N_13963);
xor U16085 (N_16085,N_11704,N_13926);
or U16086 (N_16086,N_12312,N_10921);
or U16087 (N_16087,N_11776,N_10614);
and U16088 (N_16088,N_13320,N_11047);
or U16089 (N_16089,N_10160,N_10968);
nand U16090 (N_16090,N_14452,N_11773);
or U16091 (N_16091,N_12774,N_10135);
xnor U16092 (N_16092,N_14079,N_14722);
nand U16093 (N_16093,N_11923,N_10316);
or U16094 (N_16094,N_14039,N_12838);
nand U16095 (N_16095,N_10957,N_11607);
nor U16096 (N_16096,N_14093,N_10221);
nand U16097 (N_16097,N_12280,N_12101);
nand U16098 (N_16098,N_10581,N_10765);
or U16099 (N_16099,N_11175,N_14684);
and U16100 (N_16100,N_12756,N_10366);
nand U16101 (N_16101,N_11048,N_10629);
and U16102 (N_16102,N_13485,N_12012);
nor U16103 (N_16103,N_13748,N_14290);
or U16104 (N_16104,N_11009,N_13318);
nor U16105 (N_16105,N_10856,N_11695);
xor U16106 (N_16106,N_13851,N_13070);
nor U16107 (N_16107,N_13773,N_11447);
and U16108 (N_16108,N_12746,N_13435);
or U16109 (N_16109,N_14007,N_14497);
nor U16110 (N_16110,N_10864,N_10260);
nand U16111 (N_16111,N_11921,N_13752);
or U16112 (N_16112,N_11210,N_10778);
nand U16113 (N_16113,N_10413,N_14532);
or U16114 (N_16114,N_14606,N_14801);
nor U16115 (N_16115,N_11755,N_10858);
or U16116 (N_16116,N_13539,N_10022);
nor U16117 (N_16117,N_13105,N_12564);
xnor U16118 (N_16118,N_14864,N_11190);
nor U16119 (N_16119,N_13951,N_12769);
xor U16120 (N_16120,N_13416,N_13779);
nor U16121 (N_16121,N_13562,N_12427);
nand U16122 (N_16122,N_12910,N_12184);
nand U16123 (N_16123,N_12640,N_14981);
xor U16124 (N_16124,N_10263,N_12932);
xor U16125 (N_16125,N_12159,N_10051);
nand U16126 (N_16126,N_11366,N_14960);
and U16127 (N_16127,N_10797,N_12105);
and U16128 (N_16128,N_10174,N_11815);
and U16129 (N_16129,N_14473,N_10920);
or U16130 (N_16130,N_13600,N_11844);
and U16131 (N_16131,N_13241,N_12401);
and U16132 (N_16132,N_11538,N_11280);
nor U16133 (N_16133,N_13014,N_12433);
or U16134 (N_16134,N_14189,N_13925);
nor U16135 (N_16135,N_13196,N_12594);
xnor U16136 (N_16136,N_14201,N_13941);
nand U16137 (N_16137,N_14418,N_10908);
nor U16138 (N_16138,N_12632,N_11898);
and U16139 (N_16139,N_11216,N_14854);
nor U16140 (N_16140,N_11563,N_11099);
and U16141 (N_16141,N_12676,N_10796);
nor U16142 (N_16142,N_14739,N_14292);
xnor U16143 (N_16143,N_12203,N_12056);
xnor U16144 (N_16144,N_13783,N_14293);
xnor U16145 (N_16145,N_10459,N_12864);
or U16146 (N_16146,N_12742,N_13425);
xor U16147 (N_16147,N_14477,N_11938);
or U16148 (N_16148,N_12660,N_12476);
xnor U16149 (N_16149,N_10307,N_10600);
or U16150 (N_16150,N_13690,N_14419);
or U16151 (N_16151,N_14553,N_14331);
or U16152 (N_16152,N_12673,N_13178);
nand U16153 (N_16153,N_11915,N_13850);
or U16154 (N_16154,N_12568,N_14422);
or U16155 (N_16155,N_14107,N_13713);
xor U16156 (N_16156,N_13476,N_12490);
nand U16157 (N_16157,N_11051,N_10127);
nor U16158 (N_16158,N_11544,N_11377);
nand U16159 (N_16159,N_12984,N_13167);
nor U16160 (N_16160,N_13560,N_11902);
and U16161 (N_16161,N_14843,N_14947);
or U16162 (N_16162,N_13875,N_10478);
nand U16163 (N_16163,N_13305,N_12430);
and U16164 (N_16164,N_11364,N_13935);
nand U16165 (N_16165,N_11886,N_12539);
and U16166 (N_16166,N_12149,N_13374);
or U16167 (N_16167,N_11248,N_10588);
nand U16168 (N_16168,N_14006,N_14628);
nor U16169 (N_16169,N_13692,N_10903);
nand U16170 (N_16170,N_12180,N_12475);
xnor U16171 (N_16171,N_10075,N_11656);
or U16172 (N_16172,N_11621,N_10027);
xnor U16173 (N_16173,N_11297,N_13772);
nand U16174 (N_16174,N_10821,N_10115);
and U16175 (N_16175,N_14604,N_12087);
xnor U16176 (N_16176,N_14626,N_11895);
and U16177 (N_16177,N_14865,N_14741);
nor U16178 (N_16178,N_14620,N_12874);
and U16179 (N_16179,N_10421,N_11132);
nor U16180 (N_16180,N_14206,N_13583);
and U16181 (N_16181,N_13775,N_13174);
nand U16182 (N_16182,N_13602,N_12738);
or U16183 (N_16183,N_12574,N_14765);
and U16184 (N_16184,N_10667,N_10962);
nor U16185 (N_16185,N_14993,N_11772);
xnor U16186 (N_16186,N_10262,N_12919);
or U16187 (N_16187,N_11164,N_13354);
nand U16188 (N_16188,N_13843,N_12952);
xor U16189 (N_16189,N_12027,N_13747);
and U16190 (N_16190,N_12533,N_14469);
or U16191 (N_16191,N_14018,N_12929);
and U16192 (N_16192,N_10710,N_10060);
or U16193 (N_16193,N_13906,N_14215);
xnor U16194 (N_16194,N_14240,N_12598);
xor U16195 (N_16195,N_11633,N_14764);
nand U16196 (N_16196,N_13784,N_14151);
or U16197 (N_16197,N_10756,N_14188);
nor U16198 (N_16198,N_14725,N_14491);
and U16199 (N_16199,N_13036,N_13804);
xor U16200 (N_16200,N_10983,N_13044);
nor U16201 (N_16201,N_13155,N_11661);
and U16202 (N_16202,N_12050,N_14972);
nand U16203 (N_16203,N_12055,N_11787);
and U16204 (N_16204,N_12290,N_10479);
nor U16205 (N_16205,N_12347,N_14389);
nand U16206 (N_16206,N_12638,N_14436);
or U16207 (N_16207,N_11683,N_14915);
and U16208 (N_16208,N_14807,N_13368);
or U16209 (N_16209,N_10970,N_14111);
xnor U16210 (N_16210,N_13847,N_14866);
and U16211 (N_16211,N_10808,N_11189);
or U16212 (N_16212,N_14300,N_12591);
and U16213 (N_16213,N_13146,N_10579);
or U16214 (N_16214,N_14582,N_12839);
or U16215 (N_16215,N_14859,N_12155);
and U16216 (N_16216,N_13977,N_14530);
nor U16217 (N_16217,N_13129,N_11075);
or U16218 (N_16218,N_10961,N_14616);
xor U16219 (N_16219,N_12788,N_13331);
nor U16220 (N_16220,N_12212,N_10019);
or U16221 (N_16221,N_11469,N_13068);
nor U16222 (N_16222,N_12580,N_12585);
or U16223 (N_16223,N_14106,N_10623);
xnor U16224 (N_16224,N_11129,N_12349);
and U16225 (N_16225,N_11837,N_11429);
nor U16226 (N_16226,N_11058,N_11312);
xor U16227 (N_16227,N_14271,N_14679);
nand U16228 (N_16228,N_12479,N_10410);
xnor U16229 (N_16229,N_10597,N_10130);
nor U16230 (N_16230,N_13082,N_14336);
and U16231 (N_16231,N_10770,N_14667);
nor U16232 (N_16232,N_12603,N_13442);
xor U16233 (N_16233,N_14894,N_12852);
or U16234 (N_16234,N_11957,N_14728);
xor U16235 (N_16235,N_13777,N_11859);
nand U16236 (N_16236,N_12542,N_14584);
xnor U16237 (N_16237,N_10191,N_14277);
or U16238 (N_16238,N_13737,N_10300);
nor U16239 (N_16239,N_13107,N_12879);
nand U16240 (N_16240,N_11791,N_11476);
or U16241 (N_16241,N_13532,N_11508);
xnor U16242 (N_16242,N_12902,N_13809);
and U16243 (N_16243,N_13854,N_11548);
and U16244 (N_16244,N_13494,N_10627);
and U16245 (N_16245,N_10724,N_11027);
nor U16246 (N_16246,N_12167,N_11369);
or U16247 (N_16247,N_13638,N_11637);
nand U16248 (N_16248,N_12218,N_14611);
or U16249 (N_16249,N_14770,N_10655);
or U16250 (N_16250,N_13381,N_11456);
nand U16251 (N_16251,N_13497,N_10687);
nor U16252 (N_16252,N_11565,N_11593);
xnor U16253 (N_16253,N_12550,N_14976);
nand U16254 (N_16254,N_14200,N_11082);
nand U16255 (N_16255,N_14365,N_14762);
nand U16256 (N_16256,N_13133,N_11666);
nand U16257 (N_16257,N_11731,N_14647);
and U16258 (N_16258,N_12843,N_14812);
xor U16259 (N_16259,N_12734,N_12994);
xnor U16260 (N_16260,N_10444,N_10477);
nand U16261 (N_16261,N_12631,N_14968);
nor U16262 (N_16262,N_14198,N_10700);
or U16263 (N_16263,N_10195,N_11125);
or U16264 (N_16264,N_12138,N_11389);
nand U16265 (N_16265,N_10274,N_13204);
xnor U16266 (N_16266,N_12169,N_12190);
nand U16267 (N_16267,N_12858,N_12456);
xnor U16268 (N_16268,N_10101,N_12957);
nor U16269 (N_16269,N_14531,N_12748);
xnor U16270 (N_16270,N_12186,N_10315);
and U16271 (N_16271,N_10373,N_10874);
xnor U16272 (N_16272,N_14379,N_10901);
or U16273 (N_16273,N_10192,N_11083);
nand U16274 (N_16274,N_11603,N_12891);
xnor U16275 (N_16275,N_11402,N_12389);
nor U16276 (N_16276,N_12205,N_13180);
and U16277 (N_16277,N_13332,N_12248);
nor U16278 (N_16278,N_10402,N_14874);
or U16279 (N_16279,N_11460,N_12613);
xor U16280 (N_16280,N_14895,N_12670);
nor U16281 (N_16281,N_14247,N_10744);
nor U16282 (N_16282,N_13514,N_11038);
nor U16283 (N_16283,N_14478,N_12405);
or U16284 (N_16284,N_14835,N_12728);
and U16285 (N_16285,N_12946,N_14114);
nor U16286 (N_16286,N_12054,N_14265);
xor U16287 (N_16287,N_13297,N_11973);
nor U16288 (N_16288,N_12637,N_11246);
nor U16289 (N_16289,N_10299,N_13735);
xor U16290 (N_16290,N_10772,N_13345);
xor U16291 (N_16291,N_11626,N_10070);
xnor U16292 (N_16292,N_10368,N_13325);
xor U16293 (N_16293,N_13211,N_13625);
nor U16294 (N_16294,N_10211,N_14930);
xor U16295 (N_16295,N_13264,N_13478);
or U16296 (N_16296,N_12327,N_12196);
nand U16297 (N_16297,N_10551,N_10868);
nand U16298 (N_16298,N_12718,N_13914);
nor U16299 (N_16299,N_13513,N_14031);
or U16300 (N_16300,N_11074,N_12771);
and U16301 (N_16301,N_12276,N_11948);
nand U16302 (N_16302,N_14166,N_14900);
nor U16303 (N_16303,N_12278,N_11087);
nand U16304 (N_16304,N_12798,N_13671);
nand U16305 (N_16305,N_11408,N_11185);
and U16306 (N_16306,N_10480,N_13930);
or U16307 (N_16307,N_10054,N_10754);
and U16308 (N_16308,N_11602,N_13428);
nand U16309 (N_16309,N_11032,N_11161);
and U16310 (N_16310,N_13233,N_10118);
and U16311 (N_16311,N_10486,N_14138);
and U16312 (N_16312,N_14686,N_12313);
and U16313 (N_16313,N_14848,N_12317);
xnor U16314 (N_16314,N_14678,N_10722);
xor U16315 (N_16315,N_14040,N_13911);
and U16316 (N_16316,N_10468,N_13069);
and U16317 (N_16317,N_13844,N_14541);
xnor U16318 (N_16318,N_10483,N_14410);
nor U16319 (N_16319,N_12834,N_10654);
nand U16320 (N_16320,N_12519,N_11254);
and U16321 (N_16321,N_12353,N_14227);
and U16322 (N_16322,N_11583,N_14087);
or U16323 (N_16323,N_13137,N_11677);
or U16324 (N_16324,N_11188,N_11080);
xnor U16325 (N_16325,N_12661,N_11482);
and U16326 (N_16326,N_13344,N_11788);
nor U16327 (N_16327,N_14939,N_10113);
xor U16328 (N_16328,N_13896,N_10539);
and U16329 (N_16329,N_13507,N_12363);
nand U16330 (N_16330,N_13554,N_12844);
xor U16331 (N_16331,N_10239,N_11990);
or U16332 (N_16332,N_14985,N_14089);
nand U16333 (N_16333,N_10499,N_10689);
or U16334 (N_16334,N_12575,N_13521);
nor U16335 (N_16335,N_13266,N_11037);
or U16336 (N_16336,N_11421,N_11894);
xor U16337 (N_16337,N_10122,N_14222);
nor U16338 (N_16338,N_13122,N_13750);
nor U16339 (N_16339,N_11810,N_11381);
and U16340 (N_16340,N_14204,N_12029);
xor U16341 (N_16341,N_13725,N_12408);
or U16342 (N_16342,N_13699,N_13280);
nor U16343 (N_16343,N_12699,N_10357);
nor U16344 (N_16344,N_14551,N_11994);
xnor U16345 (N_16345,N_14839,N_11174);
or U16346 (N_16346,N_12915,N_10721);
nand U16347 (N_16347,N_10648,N_14348);
nor U16348 (N_16348,N_14838,N_14788);
nand U16349 (N_16349,N_10481,N_10441);
or U16350 (N_16350,N_11562,N_12209);
xnor U16351 (N_16351,N_10451,N_12287);
or U16352 (N_16352,N_14622,N_13474);
xnor U16353 (N_16353,N_11802,N_14082);
or U16354 (N_16354,N_13191,N_11194);
or U16355 (N_16355,N_13545,N_11749);
nand U16356 (N_16356,N_12537,N_11171);
nand U16357 (N_16357,N_11874,N_10513);
or U16358 (N_16358,N_12466,N_11243);
nor U16359 (N_16359,N_11351,N_12094);
and U16360 (N_16360,N_13837,N_14537);
xnor U16361 (N_16361,N_14986,N_11715);
or U16362 (N_16362,N_13710,N_13084);
or U16363 (N_16363,N_12208,N_12118);
xnor U16364 (N_16364,N_11483,N_11823);
nor U16365 (N_16365,N_12977,N_12921);
nand U16366 (N_16366,N_11875,N_14012);
xnor U16367 (N_16367,N_13863,N_10598);
and U16368 (N_16368,N_11941,N_10422);
or U16369 (N_16369,N_10622,N_12755);
nor U16370 (N_16370,N_12132,N_11343);
and U16371 (N_16371,N_14474,N_11586);
xnor U16372 (N_16372,N_12188,N_14185);
nand U16373 (N_16373,N_12487,N_12856);
nand U16374 (N_16374,N_13096,N_10750);
xnor U16375 (N_16375,N_13481,N_11899);
xnor U16376 (N_16376,N_11780,N_12704);
xnor U16377 (N_16377,N_12971,N_13971);
nand U16378 (N_16378,N_12538,N_10230);
nor U16379 (N_16379,N_14674,N_12247);
xor U16380 (N_16380,N_13150,N_14159);
nor U16381 (N_16381,N_10646,N_14852);
xor U16382 (N_16382,N_10528,N_10802);
nand U16383 (N_16383,N_11566,N_12939);
nand U16384 (N_16384,N_11678,N_14910);
nor U16385 (N_16385,N_13363,N_10548);
nor U16386 (N_16386,N_13862,N_11611);
nor U16387 (N_16387,N_12955,N_13579);
nand U16388 (N_16388,N_14563,N_13893);
and U16389 (N_16389,N_13310,N_13757);
nand U16390 (N_16390,N_13644,N_14890);
nand U16391 (N_16391,N_11265,N_10911);
and U16392 (N_16392,N_14932,N_10847);
nand U16393 (N_16393,N_12595,N_11479);
nand U16394 (N_16394,N_14951,N_11856);
or U16395 (N_16395,N_13239,N_12892);
and U16396 (N_16396,N_13013,N_11407);
and U16397 (N_16397,N_12993,N_12074);
and U16398 (N_16398,N_11561,N_12488);
nor U16399 (N_16399,N_14974,N_12944);
nand U16400 (N_16400,N_11892,N_13288);
and U16401 (N_16401,N_14135,N_12954);
xnor U16402 (N_16402,N_11514,N_12873);
xnor U16403 (N_16403,N_13161,N_14133);
nand U16404 (N_16404,N_11995,N_14167);
or U16405 (N_16405,N_10763,N_14153);
xnor U16406 (N_16406,N_12522,N_12403);
or U16407 (N_16407,N_14302,N_11019);
nor U16408 (N_16408,N_10638,N_12114);
nor U16409 (N_16409,N_10023,N_14502);
nand U16410 (N_16410,N_11974,N_14506);
nor U16411 (N_16411,N_13064,N_11457);
xnor U16412 (N_16412,N_11842,N_11249);
nor U16413 (N_16413,N_12662,N_10871);
nor U16414 (N_16414,N_13599,N_11956);
or U16415 (N_16415,N_12577,N_11663);
xnor U16416 (N_16416,N_13079,N_12505);
nor U16417 (N_16417,N_12224,N_10715);
or U16418 (N_16418,N_11311,N_13877);
nand U16419 (N_16419,N_10430,N_13769);
nor U16420 (N_16420,N_12532,N_10712);
nor U16421 (N_16421,N_11286,N_10591);
nand U16422 (N_16422,N_14416,N_13704);
and U16423 (N_16423,N_10311,N_12610);
and U16424 (N_16424,N_11783,N_14658);
xnor U16425 (N_16425,N_14578,N_14908);
nor U16426 (N_16426,N_14174,N_11804);
or U16427 (N_16427,N_14101,N_14108);
nand U16428 (N_16428,N_13258,N_13153);
and U16429 (N_16429,N_11674,N_13889);
xor U16430 (N_16430,N_14881,N_14811);
nor U16431 (N_16431,N_13250,N_12525);
xor U16432 (N_16432,N_12448,N_13767);
and U16433 (N_16433,N_10381,N_10085);
and U16434 (N_16434,N_10374,N_13388);
nand U16435 (N_16435,N_12681,N_14374);
and U16436 (N_16436,N_10515,N_12938);
or U16437 (N_16437,N_12366,N_11978);
nand U16438 (N_16438,N_11669,N_13975);
nand U16439 (N_16439,N_14585,N_13883);
and U16440 (N_16440,N_11308,N_13198);
and U16441 (N_16441,N_11303,N_14926);
xor U16442 (N_16442,N_11371,N_11014);
nand U16443 (N_16443,N_12870,N_12017);
nand U16444 (N_16444,N_10753,N_11113);
nor U16445 (N_16445,N_10825,N_11236);
and U16446 (N_16446,N_10987,N_14332);
or U16447 (N_16447,N_13512,N_14433);
or U16448 (N_16448,N_14396,N_14333);
nor U16449 (N_16449,N_11177,N_11775);
xnor U16450 (N_16450,N_13972,N_14472);
and U16451 (N_16451,N_11644,N_13268);
xor U16452 (N_16452,N_11434,N_10194);
xnor U16453 (N_16453,N_11359,N_13116);
xnor U16454 (N_16454,N_14605,N_10822);
or U16455 (N_16455,N_12160,N_10360);
xnor U16456 (N_16456,N_12454,N_13868);
nand U16457 (N_16457,N_12171,N_10369);
or U16458 (N_16458,N_13910,N_10134);
and U16459 (N_16459,N_10640,N_11225);
nor U16460 (N_16460,N_11259,N_11512);
and U16461 (N_16461,N_11338,N_12305);
and U16462 (N_16462,N_11570,N_10929);
or U16463 (N_16463,N_12380,N_13300);
nand U16464 (N_16464,N_14518,N_10839);
and U16465 (N_16465,N_12298,N_14914);
nand U16466 (N_16466,N_14889,N_12412);
nand U16467 (N_16467,N_13247,N_11610);
or U16468 (N_16468,N_10149,N_14378);
nor U16469 (N_16469,N_13407,N_10553);
or U16470 (N_16470,N_13203,N_13045);
xor U16471 (N_16471,N_14024,N_12014);
nand U16472 (N_16472,N_12072,N_14406);
or U16473 (N_16473,N_10438,N_11606);
or U16474 (N_16474,N_11662,N_10618);
xor U16475 (N_16475,N_11432,N_13965);
xnor U16476 (N_16476,N_13234,N_11943);
or U16477 (N_16477,N_12368,N_12686);
xnor U16478 (N_16478,N_14250,N_12452);
xor U16479 (N_16479,N_10339,N_14887);
nor U16480 (N_16480,N_13932,N_14669);
or U16481 (N_16481,N_11585,N_11205);
nor U16482 (N_16482,N_13712,N_14656);
or U16483 (N_16483,N_14130,N_10974);
nand U16484 (N_16484,N_14781,N_12536);
nor U16485 (N_16485,N_12592,N_12264);
or U16486 (N_16486,N_10024,N_12251);
or U16487 (N_16487,N_14110,N_11614);
or U16488 (N_16488,N_14642,N_14897);
nand U16489 (N_16489,N_13248,N_11855);
and U16490 (N_16490,N_10279,N_11110);
xnor U16491 (N_16491,N_12908,N_10482);
or U16492 (N_16492,N_11575,N_13281);
xor U16493 (N_16493,N_11226,N_11022);
nand U16494 (N_16494,N_10758,N_13207);
nand U16495 (N_16495,N_14360,N_12424);
or U16496 (N_16496,N_11033,N_10965);
and U16497 (N_16497,N_13592,N_14754);
and U16498 (N_16498,N_14242,N_13273);
xnor U16499 (N_16499,N_11937,N_13049);
or U16500 (N_16500,N_14235,N_14368);
xnor U16501 (N_16501,N_11372,N_11156);
nand U16502 (N_16502,N_13098,N_11631);
xnor U16503 (N_16503,N_13152,N_13020);
and U16504 (N_16504,N_12432,N_10885);
and U16505 (N_16505,N_13639,N_13158);
nor U16506 (N_16506,N_13255,N_13768);
xor U16507 (N_16507,N_11178,N_11309);
nor U16508 (N_16508,N_13901,N_11331);
xor U16509 (N_16509,N_11078,N_11612);
xnor U16510 (N_16510,N_11195,N_14305);
or U16511 (N_16511,N_14239,N_14909);
xor U16512 (N_16512,N_10543,N_10138);
xor U16513 (N_16513,N_14427,N_12762);
xor U16514 (N_16514,N_10606,N_10001);
and U16515 (N_16515,N_11274,N_11464);
or U16516 (N_16516,N_10052,N_12390);
nor U16517 (N_16517,N_14264,N_11052);
xnor U16518 (N_16518,N_10718,N_14521);
nand U16519 (N_16519,N_12812,N_10894);
xnor U16520 (N_16520,N_12885,N_14749);
nor U16521 (N_16521,N_11107,N_11511);
or U16522 (N_16522,N_11200,N_10265);
xor U16523 (N_16523,N_10702,N_12513);
or U16524 (N_16524,N_11394,N_13749);
nor U16525 (N_16525,N_11439,N_13657);
nand U16526 (N_16526,N_11734,N_12047);
xor U16527 (N_16527,N_11035,N_12030);
and U16528 (N_16528,N_12790,N_12768);
and U16529 (N_16529,N_10208,N_11365);
nor U16530 (N_16530,N_10930,N_10617);
nand U16531 (N_16531,N_13970,N_11329);
xnor U16532 (N_16532,N_11636,N_11521);
or U16533 (N_16533,N_11720,N_12489);
and U16534 (N_16534,N_12444,N_12772);
and U16535 (N_16535,N_13408,N_12063);
or U16536 (N_16536,N_11922,N_11597);
or U16537 (N_16537,N_14877,N_13647);
xor U16538 (N_16538,N_12593,N_11399);
nand U16539 (N_16539,N_10953,N_10572);
xor U16540 (N_16540,N_12503,N_10869);
and U16541 (N_16541,N_10336,N_10018);
or U16542 (N_16542,N_10364,N_10711);
xor U16543 (N_16543,N_11442,N_10788);
and U16544 (N_16544,N_12482,N_10757);
nand U16545 (N_16545,N_14919,N_13660);
nor U16546 (N_16546,N_12355,N_14823);
xor U16547 (N_16547,N_13606,N_14112);
nand U16548 (N_16548,N_14260,N_13780);
nand U16549 (N_16549,N_11517,N_14500);
or U16550 (N_16550,N_13995,N_14661);
nor U16551 (N_16551,N_11201,N_11642);
nand U16552 (N_16552,N_11880,N_12126);
nand U16553 (N_16553,N_14878,N_13130);
nor U16554 (N_16554,N_12822,N_12085);
or U16555 (N_16555,N_11709,N_12629);
nor U16556 (N_16556,N_12474,N_12502);
nand U16557 (N_16557,N_14069,N_14552);
nor U16558 (N_16558,N_13427,N_11834);
or U16559 (N_16559,N_12497,N_10807);
xor U16560 (N_16560,N_14891,N_14147);
and U16561 (N_16561,N_14841,N_10992);
or U16562 (N_16562,N_12689,N_12625);
nor U16563 (N_16563,N_13726,N_13302);
or U16564 (N_16564,N_11628,N_13655);
nor U16565 (N_16565,N_14931,N_10057);
and U16566 (N_16566,N_13905,N_12720);
nor U16567 (N_16567,N_12521,N_13601);
xnor U16568 (N_16568,N_13555,N_13458);
or U16569 (N_16569,N_10707,N_10406);
nor U16570 (N_16570,N_12925,N_14053);
nand U16571 (N_16571,N_12120,N_12166);
and U16572 (N_16572,N_13052,N_14869);
and U16573 (N_16573,N_10291,N_14177);
nor U16574 (N_16574,N_13162,N_11494);
nor U16575 (N_16575,N_14109,N_14803);
nor U16576 (N_16576,N_10454,N_14413);
nor U16577 (N_16577,N_12857,N_11747);
and U16578 (N_16578,N_12733,N_13015);
xor U16579 (N_16579,N_13357,N_13981);
nand U16580 (N_16580,N_11053,N_11616);
or U16581 (N_16581,N_14444,N_11413);
nor U16582 (N_16582,N_13618,N_10343);
nand U16583 (N_16583,N_14746,N_10284);
and U16584 (N_16584,N_11576,N_10532);
and U16585 (N_16585,N_13672,N_10852);
nor U16586 (N_16586,N_10704,N_10996);
or U16587 (N_16587,N_10352,N_12259);
or U16588 (N_16588,N_12028,N_13624);
xor U16589 (N_16589,N_10703,N_12985);
or U16590 (N_16590,N_14460,N_13456);
and U16591 (N_16591,N_14254,N_12999);
xnor U16592 (N_16592,N_14480,N_14808);
xnor U16593 (N_16593,N_13529,N_11839);
nand U16594 (N_16594,N_11357,N_11318);
nand U16595 (N_16595,N_14920,N_10066);
and U16596 (N_16596,N_10164,N_10470);
or U16597 (N_16597,N_10394,N_12043);
nor U16598 (N_16598,N_12590,N_12888);
nor U16599 (N_16599,N_12115,N_13952);
xnor U16600 (N_16600,N_14338,N_10111);
and U16601 (N_16601,N_10226,N_14358);
or U16602 (N_16602,N_10403,N_12340);
nor U16603 (N_16603,N_11940,N_10726);
nor U16604 (N_16604,N_12083,N_14008);
nor U16605 (N_16605,N_12411,N_14496);
nand U16606 (N_16606,N_12710,N_12291);
nand U16607 (N_16607,N_10376,N_14068);
xnor U16608 (N_16608,N_14439,N_13030);
nor U16609 (N_16609,N_12711,N_11882);
nand U16610 (N_16610,N_11970,N_13282);
nand U16611 (N_16611,N_11293,N_13206);
or U16612 (N_16612,N_11134,N_14813);
xor U16613 (N_16613,N_14483,N_14565);
nand U16614 (N_16614,N_12143,N_12586);
nor U16615 (N_16615,N_12776,N_10338);
and U16616 (N_16616,N_13683,N_10330);
xor U16617 (N_16617,N_13538,N_14395);
and U16618 (N_16618,N_10109,N_14345);
nor U16619 (N_16619,N_12240,N_12928);
xor U16620 (N_16620,N_12107,N_13942);
nor U16621 (N_16621,N_11862,N_13681);
or U16622 (N_16622,N_11167,N_12646);
xnor U16623 (N_16623,N_11577,N_12740);
xor U16624 (N_16624,N_13631,N_13484);
xnor U16625 (N_16625,N_12258,N_11386);
and U16626 (N_16626,N_13436,N_11779);
or U16627 (N_16627,N_13598,N_11336);
nor U16628 (N_16628,N_10151,N_10931);
or U16629 (N_16629,N_14953,N_14384);
or U16630 (N_16630,N_10303,N_14768);
nor U16631 (N_16631,N_12042,N_10156);
and U16632 (N_16632,N_13742,N_11969);
or U16633 (N_16633,N_13927,N_12806);
xor U16634 (N_16634,N_12557,N_10792);
and U16635 (N_16635,N_11252,N_11685);
and U16636 (N_16636,N_10653,N_13005);
nand U16637 (N_16637,N_10610,N_10110);
nor U16638 (N_16638,N_12112,N_10671);
or U16639 (N_16639,N_12950,N_10008);
xnor U16640 (N_16640,N_11879,N_11952);
xor U16641 (N_16641,N_10725,N_13135);
nand U16642 (N_16642,N_11307,N_11196);
and U16643 (N_16643,N_10396,N_11322);
nor U16644 (N_16644,N_11348,N_13132);
and U16645 (N_16645,N_11955,N_14772);
nand U16646 (N_16646,N_14645,N_11044);
and U16647 (N_16647,N_14558,N_10267);
or U16648 (N_16648,N_11419,N_11235);
or U16649 (N_16649,N_14257,N_11300);
xnor U16650 (N_16650,N_10014,N_14370);
xnor U16651 (N_16651,N_12303,N_12404);
or U16652 (N_16652,N_13110,N_14464);
nand U16653 (N_16653,N_10749,N_12535);
or U16654 (N_16654,N_12067,N_11871);
nor U16655 (N_16655,N_14760,N_11809);
and U16656 (N_16656,N_12022,N_12350);
nor U16657 (N_16657,N_10137,N_12609);
nand U16658 (N_16658,N_13039,N_11682);
xnor U16659 (N_16659,N_13665,N_10951);
xor U16660 (N_16660,N_11526,N_10674);
xnor U16661 (N_16661,N_10625,N_14168);
nor U16662 (N_16662,N_11213,N_13406);
or U16663 (N_16663,N_10666,N_14924);
and U16664 (N_16664,N_10318,N_11850);
xor U16665 (N_16665,N_12273,N_12147);
nand U16666 (N_16666,N_12331,N_13620);
and U16667 (N_16667,N_10899,N_11157);
nor U16668 (N_16668,N_10891,N_14787);
and U16669 (N_16669,N_14170,N_12716);
xor U16670 (N_16670,N_10549,N_12760);
xnor U16671 (N_16671,N_14899,N_14997);
nand U16672 (N_16672,N_13202,N_14538);
nor U16673 (N_16673,N_12884,N_12866);
nor U16674 (N_16674,N_12069,N_11092);
and U16675 (N_16675,N_11821,N_12296);
nand U16676 (N_16676,N_11697,N_10428);
xnor U16677 (N_16677,N_12600,N_12152);
nand U16678 (N_16678,N_14995,N_11046);
xor U16679 (N_16679,N_13962,N_11983);
nand U16680 (N_16680,N_11341,N_10355);
xnor U16681 (N_16681,N_13724,N_14182);
or U16682 (N_16682,N_13283,N_10801);
xnor U16683 (N_16683,N_13413,N_14790);
xnor U16684 (N_16684,N_11724,N_11503);
nor U16685 (N_16685,N_11165,N_13327);
or U16686 (N_16686,N_14445,N_13100);
and U16687 (N_16687,N_13873,N_10604);
and U16688 (N_16688,N_10595,N_12823);
or U16689 (N_16689,N_10895,N_12426);
nand U16690 (N_16690,N_14294,N_11425);
nand U16691 (N_16691,N_14400,N_11401);
nand U16692 (N_16692,N_13308,N_13628);
xnor U16693 (N_16693,N_10182,N_13170);
xnor U16694 (N_16694,N_13106,N_12865);
nor U16695 (N_16695,N_13978,N_10015);
nor U16696 (N_16696,N_14517,N_12829);
nand U16697 (N_16697,N_10205,N_14315);
and U16698 (N_16698,N_12008,N_11301);
nor U16699 (N_16699,N_12500,N_13795);
nor U16700 (N_16700,N_12399,N_10738);
nand U16701 (N_16701,N_13674,N_11361);
or U16702 (N_16702,N_10043,N_11197);
and U16703 (N_16703,N_14567,N_12079);
or U16704 (N_16704,N_13000,N_14030);
or U16705 (N_16705,N_12422,N_12397);
or U16706 (N_16706,N_13519,N_14627);
or U16707 (N_16707,N_14774,N_14872);
xnor U16708 (N_16708,N_12758,N_12081);
or U16709 (N_16709,N_10940,N_10255);
nand U16710 (N_16710,N_14283,N_10079);
or U16711 (N_16711,N_11090,N_10547);
or U16712 (N_16712,N_13166,N_12330);
nor U16713 (N_16713,N_13260,N_14814);
and U16714 (N_16714,N_11018,N_10047);
xor U16715 (N_16715,N_14716,N_13785);
xnor U16716 (N_16716,N_12959,N_11933);
or U16717 (N_16717,N_11256,N_13275);
nor U16718 (N_16718,N_14103,N_11445);
or U16719 (N_16719,N_12339,N_11056);
or U16720 (N_16720,N_10865,N_13691);
nor U16721 (N_16721,N_13522,N_14724);
nand U16722 (N_16722,N_10461,N_14952);
or U16723 (N_16723,N_11572,N_10165);
xor U16724 (N_16724,N_10129,N_10824);
nand U16725 (N_16725,N_10133,N_10119);
and U16726 (N_16726,N_13432,N_12626);
xor U16727 (N_16727,N_10375,N_12238);
nor U16728 (N_16728,N_14075,N_11758);
xnor U16729 (N_16729,N_10592,N_10237);
and U16730 (N_16730,N_12714,N_14417);
or U16731 (N_16731,N_10789,N_13815);
xor U16732 (N_16732,N_14081,N_12973);
and U16733 (N_16733,N_11094,N_14092);
nor U16734 (N_16734,N_12420,N_13127);
nand U16735 (N_16735,N_12153,N_10705);
nor U16736 (N_16736,N_14536,N_11335);
or U16737 (N_16737,N_13123,N_12787);
or U16738 (N_16738,N_11574,N_10728);
or U16739 (N_16739,N_14154,N_12724);
xnor U16740 (N_16740,N_14295,N_10809);
nor U16741 (N_16741,N_14249,N_11370);
and U16742 (N_16742,N_14691,N_11725);
xnor U16743 (N_16743,N_13217,N_12279);
and U16744 (N_16744,N_14682,N_12987);
or U16745 (N_16745,N_12978,N_12034);
nor U16746 (N_16746,N_12193,N_13537);
xnor U16747 (N_16747,N_14800,N_11050);
nor U16748 (N_16748,N_14361,N_11897);
xnor U16749 (N_16749,N_10434,N_13330);
or U16750 (N_16750,N_14571,N_11568);
xnor U16751 (N_16751,N_11546,N_11347);
nor U16752 (N_16752,N_14051,N_11798);
nor U16753 (N_16753,N_13791,N_13396);
nand U16754 (N_16754,N_12918,N_12992);
and U16755 (N_16755,N_14984,N_12414);
nor U16756 (N_16756,N_13309,N_14149);
or U16757 (N_16757,N_12697,N_10158);
and U16758 (N_16758,N_10860,N_10170);
nor U16759 (N_16759,N_12191,N_14918);
and U16760 (N_16760,N_11545,N_14639);
and U16761 (N_16761,N_13961,N_14054);
nor U16762 (N_16762,N_10504,N_10636);
and U16763 (N_16763,N_10372,N_13397);
or U16764 (N_16764,N_10184,N_14845);
xor U16765 (N_16765,N_11947,N_12556);
nand U16766 (N_16766,N_10999,N_10516);
or U16767 (N_16767,N_13043,N_11138);
xnor U16768 (N_16768,N_12859,N_10734);
and U16769 (N_16769,N_11706,N_14369);
or U16770 (N_16770,N_10838,N_10016);
nand U16771 (N_16771,N_13687,N_11535);
or U16772 (N_16772,N_10439,N_11283);
nand U16773 (N_16773,N_13733,N_12253);
nor U16774 (N_16774,N_10089,N_14817);
xnor U16775 (N_16775,N_12791,N_13836);
nor U16776 (N_16776,N_12199,N_12569);
xor U16777 (N_16777,N_12048,N_13654);
or U16778 (N_16778,N_10245,N_13053);
nand U16779 (N_16779,N_12351,N_10314);
or U16780 (N_16780,N_10882,N_13653);
and U16781 (N_16781,N_10708,N_11000);
nor U16782 (N_16782,N_14941,N_10740);
nand U16783 (N_16783,N_13358,N_13716);
xor U16784 (N_16784,N_12073,N_10849);
nor U16785 (N_16785,N_14113,N_12470);
nor U16786 (N_16786,N_13103,N_12814);
xnor U16787 (N_16787,N_14759,N_14197);
or U16788 (N_16788,N_11946,N_10677);
nor U16789 (N_16789,N_14016,N_12223);
nand U16790 (N_16790,N_10840,N_10573);
xor U16791 (N_16791,N_14105,N_12481);
nand U16792 (N_16792,N_13673,N_12271);
xnor U16793 (N_16793,N_10286,N_12808);
and U16794 (N_16794,N_10020,N_14488);
or U16795 (N_16795,N_10851,N_10919);
and U16796 (N_16796,N_14231,N_14858);
nand U16797 (N_16797,N_12304,N_13262);
nor U16798 (N_16798,N_13745,N_11930);
nor U16799 (N_16799,N_13333,N_11623);
nor U16800 (N_16800,N_11221,N_11696);
and U16801 (N_16801,N_11245,N_10295);
nor U16802 (N_16802,N_14426,N_12916);
or U16803 (N_16803,N_12294,N_14046);
nand U16804 (N_16804,N_10501,N_12133);
nand U16805 (N_16805,N_14276,N_13424);
or U16806 (N_16806,N_12005,N_13187);
nand U16807 (N_16807,N_10304,N_13055);
xnor U16808 (N_16808,N_10059,N_12956);
or U16809 (N_16809,N_13051,N_14714);
nand U16810 (N_16810,N_11238,N_12588);
nor U16811 (N_16811,N_11288,N_13075);
or U16812 (N_16812,N_14312,N_14161);
and U16813 (N_16813,N_11459,N_12239);
xnor U16814 (N_16814,N_14751,N_14646);
nor U16815 (N_16815,N_10805,N_11390);
or U16816 (N_16816,N_10202,N_12754);
xnor U16817 (N_16817,N_13086,N_14038);
xnor U16818 (N_16818,N_14967,N_12136);
and U16819 (N_16819,N_10900,N_13179);
and U16820 (N_16820,N_10257,N_14306);
or U16821 (N_16821,N_10250,N_13685);
or U16822 (N_16822,N_14144,N_10742);
nand U16823 (N_16823,N_14255,N_13090);
nor U16824 (N_16824,N_11906,N_12324);
nand U16825 (N_16825,N_11383,N_11079);
nor U16826 (N_16826,N_10510,N_13175);
or U16827 (N_16827,N_11658,N_14612);
nor U16828 (N_16828,N_12318,N_10665);
or U16829 (N_16829,N_12669,N_12402);
nand U16830 (N_16830,N_12527,N_10698);
and U16831 (N_16831,N_12703,N_10370);
xor U16832 (N_16832,N_12972,N_12000);
nor U16833 (N_16833,N_13945,N_13642);
xor U16834 (N_16834,N_13430,N_13376);
nand U16835 (N_16835,N_14059,N_10938);
and U16836 (N_16836,N_14527,N_14451);
xnor U16837 (N_16837,N_14355,N_12421);
nand U16838 (N_16838,N_13042,N_14274);
or U16839 (N_16839,N_11753,N_13915);
and U16840 (N_16840,N_13457,N_12793);
xnor U16841 (N_16841,N_11966,N_11680);
and U16842 (N_16842,N_14350,N_10518);
nand U16843 (N_16843,N_14218,N_12439);
or U16844 (N_16844,N_11220,N_13694);
nand U16845 (N_16845,N_11718,N_14086);
or U16846 (N_16846,N_12757,N_14211);
nor U16847 (N_16847,N_11264,N_10889);
nor U16848 (N_16848,N_10152,N_10325);
nor U16849 (N_16849,N_13352,N_11059);
and U16850 (N_16850,N_10389,N_10271);
nand U16851 (N_16851,N_13759,N_10399);
nor U16852 (N_16852,N_11358,N_13897);
xnor U16853 (N_16853,N_14344,N_11581);
nand U16854 (N_16854,N_13270,N_12841);
or U16855 (N_16855,N_12321,N_13800);
xor U16856 (N_16856,N_12582,N_11872);
xnor U16857 (N_16857,N_10835,N_13968);
or U16858 (N_16858,N_12821,N_11097);
xor U16859 (N_16859,N_10870,N_13181);
or U16860 (N_16860,N_11253,N_10248);
nor U16861 (N_16861,N_14750,N_11163);
nor U16862 (N_16862,N_13987,N_12940);
xor U16863 (N_16863,N_10000,N_14288);
nor U16864 (N_16864,N_13801,N_11916);
nand U16865 (N_16865,N_11255,N_14238);
nand U16866 (N_16866,N_14621,N_13938);
or U16867 (N_16867,N_12872,N_11619);
and U16868 (N_16868,N_14637,N_14449);
xor U16869 (N_16869,N_13221,N_11766);
xor U16870 (N_16870,N_14183,N_13078);
and U16871 (N_16871,N_12435,N_14726);
xnor U16872 (N_16872,N_14021,N_14570);
and U16873 (N_16873,N_14404,N_10685);
nor U16874 (N_16874,N_13944,N_14263);
nor U16875 (N_16875,N_14840,N_13346);
and U16876 (N_16876,N_12231,N_14207);
or U16877 (N_16877,N_12674,N_11654);
nand U16878 (N_16878,N_12778,N_10563);
xor U16879 (N_16879,N_12428,N_10791);
and U16880 (N_16880,N_14010,N_14490);
and U16881 (N_16881,N_12499,N_11736);
or U16882 (N_16882,N_13418,N_11011);
nor U16883 (N_16883,N_13670,N_14443);
or U16884 (N_16884,N_10678,N_14399);
and U16885 (N_16885,N_14763,N_13786);
nand U16886 (N_16886,N_13060,N_12930);
xnor U16887 (N_16887,N_10450,N_11404);
and U16888 (N_16888,N_14285,N_11848);
nor U16889 (N_16889,N_14169,N_13964);
xnor U16890 (N_16890,N_10218,N_12867);
nand U16891 (N_16891,N_11595,N_14035);
and U16892 (N_16892,N_13429,N_14137);
and U16893 (N_16893,N_14753,N_14132);
nor U16894 (N_16894,N_13285,N_14373);
nand U16895 (N_16895,N_13520,N_10764);
nand U16896 (N_16896,N_13077,N_14581);
nor U16897 (N_16897,N_12049,N_14557);
nand U16898 (N_16898,N_12394,N_11743);
xnor U16899 (N_16899,N_14734,N_14733);
or U16900 (N_16900,N_13887,N_12308);
nor U16901 (N_16901,N_11061,N_11615);
nand U16902 (N_16902,N_12495,N_10320);
and U16903 (N_16903,N_14085,N_12161);
and U16904 (N_16904,N_10672,N_11746);
nand U16905 (N_16905,N_13525,N_11625);
nor U16906 (N_16906,N_12387,N_11261);
and U16907 (N_16907,N_12285,N_11176);
nand U16908 (N_16908,N_11444,N_13659);
xnor U16909 (N_16909,N_14798,N_10234);
nand U16910 (N_16910,N_14989,N_11761);
nor U16911 (N_16911,N_11569,N_10222);
and U16912 (N_16912,N_12111,N_11436);
nand U16913 (N_16913,N_13438,N_12878);
nand U16914 (N_16914,N_10603,N_10596);
nand U16915 (N_16915,N_14498,N_12103);
and U16916 (N_16916,N_12491,N_11441);
nand U16917 (N_16917,N_12837,N_10828);
and U16918 (N_16918,N_13089,N_14766);
or U16919 (N_16919,N_13823,N_10077);
nand U16920 (N_16920,N_13566,N_13169);
xnor U16921 (N_16921,N_12145,N_12628);
xor U16922 (N_16922,N_14634,N_12207);
nor U16923 (N_16923,N_11984,N_13001);
nor U16924 (N_16924,N_10061,N_14831);
nand U16925 (N_16925,N_10946,N_13236);
nand U16926 (N_16926,N_14950,N_11471);
nand U16927 (N_16927,N_11604,N_10065);
xnor U16928 (N_16928,N_13904,N_13523);
nand U16929 (N_16929,N_13348,N_13865);
nand U16930 (N_16930,N_10494,N_10793);
nor U16931 (N_16931,N_13729,N_13996);
nor U16932 (N_16932,N_14179,N_10155);
nor U16933 (N_16933,N_10180,N_13755);
nand U16934 (N_16934,N_12745,N_14630);
or U16935 (N_16935,N_12584,N_11971);
nor U16936 (N_16936,N_10490,N_10187);
nor U16937 (N_16937,N_13955,N_13727);
nand U16938 (N_16938,N_12323,N_11650);
or U16939 (N_16939,N_13404,N_12078);
nor U16940 (N_16940,N_10409,N_10837);
or U16941 (N_16941,N_10794,N_10994);
nor U16942 (N_16942,N_11354,N_10615);
and U16943 (N_16943,N_13825,N_10952);
and U16944 (N_16944,N_14711,N_14307);
xnor U16945 (N_16945,N_12667,N_13542);
nor U16946 (N_16946,N_10773,N_10228);
nand U16947 (N_16947,N_12562,N_10449);
and U16948 (N_16948,N_10391,N_10937);
and U16949 (N_16949,N_14729,N_14364);
nand U16950 (N_16950,N_12486,N_13993);
nor U16951 (N_16951,N_11945,N_10934);
nand U16952 (N_16952,N_13091,N_11362);
or U16953 (N_16953,N_13024,N_14343);
nor U16954 (N_16954,N_13569,N_10036);
and U16955 (N_16955,N_12602,N_11477);
and U16956 (N_16956,N_12227,N_10266);
or U16957 (N_16957,N_13034,N_12058);
nor U16958 (N_16958,N_10686,N_12842);
nand U16959 (N_16959,N_12214,N_11144);
or U16960 (N_16960,N_10979,N_12254);
or U16961 (N_16961,N_13372,N_10282);
nor U16962 (N_16962,N_12709,N_12611);
nor U16963 (N_16963,N_12178,N_11122);
nor U16964 (N_16964,N_10104,N_12023);
or U16965 (N_16965,N_10073,N_14821);
and U16966 (N_16966,N_13756,N_13259);
xor U16967 (N_16967,N_11928,N_14723);
and U16968 (N_16968,N_11170,N_14991);
nor U16969 (N_16969,N_13958,N_11473);
xnor U16970 (N_16970,N_10609,N_11638);
xor U16971 (N_16971,N_13652,N_11640);
nand U16972 (N_16972,N_12459,N_11700);
and U16973 (N_16973,N_12506,N_10607);
or U16974 (N_16974,N_13037,N_10342);
and U16975 (N_16975,N_11124,N_12561);
xnor U16976 (N_16976,N_10766,N_12684);
and U16977 (N_16977,N_11803,N_13021);
or U16978 (N_16978,N_10989,N_14882);
and U16979 (N_16979,N_11499,N_11693);
nand U16980 (N_16980,N_12068,N_11410);
nor U16981 (N_16981,N_13839,N_14492);
nand U16982 (N_16982,N_13840,N_12828);
or U16983 (N_16983,N_11154,N_10017);
and U16984 (N_16984,N_11634,N_12326);
or U16985 (N_16985,N_13232,N_13398);
or U16986 (N_16986,N_11490,N_11500);
nor U16987 (N_16987,N_12309,N_12036);
nor U16988 (N_16988,N_12572,N_11228);
nor U16989 (N_16989,N_11800,N_12691);
or U16990 (N_16990,N_14412,N_13720);
xor U16991 (N_16991,N_14234,N_12384);
and U16992 (N_16992,N_10814,N_14660);
xnor U16993 (N_16993,N_12926,N_10069);
and U16994 (N_16994,N_14061,N_12377);
nand U16995 (N_16995,N_12346,N_12912);
or U16996 (N_16996,N_14004,N_14970);
xnor U16997 (N_16997,N_13184,N_14767);
xor U16998 (N_16998,N_14128,N_13895);
nor U16999 (N_16999,N_14339,N_10660);
nor U17000 (N_17000,N_10139,N_14334);
nand U17001 (N_17001,N_14576,N_11328);
nor U17002 (N_17002,N_14202,N_10525);
and U17003 (N_17003,N_11833,N_14341);
xor U17004 (N_17004,N_10013,N_14697);
or U17005 (N_17005,N_14793,N_12727);
xor U17006 (N_17006,N_10731,N_10301);
xor U17007 (N_17007,N_13667,N_14907);
xnor U17008 (N_17008,N_11337,N_10035);
and U17009 (N_17009,N_11289,N_10680);
xnor U17010 (N_17010,N_12379,N_13379);
xor U17011 (N_17011,N_13142,N_13451);
and U17012 (N_17012,N_12679,N_14499);
xnor U17013 (N_17013,N_13879,N_12299);
or U17014 (N_17014,N_14441,N_10693);
or U17015 (N_17015,N_10055,N_12455);
or U17016 (N_17016,N_12484,N_11287);
and U17017 (N_17017,N_13637,N_11835);
nor U17018 (N_17018,N_10695,N_12526);
and U17019 (N_17019,N_14871,N_12010);
nand U17020 (N_17020,N_14973,N_14045);
xnor U17021 (N_17021,N_10787,N_11098);
xnor U17022 (N_17022,N_13415,N_14390);
nor U17023 (N_17023,N_14475,N_13677);
nand U17024 (N_17024,N_14220,N_13740);
and U17025 (N_17025,N_13813,N_11466);
xor U17026 (N_17026,N_14824,N_13099);
nand U17027 (N_17027,N_13007,N_14695);
or U17028 (N_17028,N_10815,N_14638);
or U17029 (N_17029,N_14580,N_13033);
nor U17030 (N_17030,N_14654,N_12975);
xnor U17031 (N_17031,N_11100,N_14902);
nand U17032 (N_17032,N_12270,N_14608);
nor U17033 (N_17033,N_11391,N_10500);
nor U17034 (N_17034,N_12687,N_13473);
nand U17035 (N_17035,N_12851,N_12076);
nand U17036 (N_17036,N_11567,N_14421);
or U17037 (N_17037,N_12801,N_11901);
nand U17038 (N_17038,N_10179,N_11437);
and U17039 (N_17039,N_14486,N_11549);
nand U17040 (N_17040,N_13577,N_14922);
nand U17041 (N_17041,N_14349,N_14655);
xor U17042 (N_17042,N_13866,N_11294);
or U17043 (N_17043,N_12391,N_13633);
nand U17044 (N_17044,N_13614,N_11794);
or U17045 (N_17045,N_13279,N_13766);
and U17046 (N_17046,N_10243,N_14588);
nand U17047 (N_17047,N_11091,N_10029);
xnor U17048 (N_17048,N_13820,N_14317);
xor U17049 (N_17049,N_13401,N_10010);
and U17050 (N_17050,N_13029,N_14296);
and U17051 (N_17051,N_14827,N_14381);
xor U17052 (N_17052,N_10777,N_12931);
nor U17053 (N_17053,N_14438,N_13294);
nor U17054 (N_17054,N_11145,N_10804);
and U17055 (N_17055,N_11578,N_12795);
or U17056 (N_17056,N_10283,N_12071);
xnor U17057 (N_17057,N_11622,N_11093);
or U17058 (N_17058,N_10637,N_10220);
xor U17059 (N_17059,N_10322,N_11260);
nor U17060 (N_17060,N_10827,N_11985);
nand U17061 (N_17061,N_12255,N_10038);
and U17062 (N_17062,N_10395,N_14978);
xnor U17063 (N_17063,N_11689,N_11759);
and U17064 (N_17064,N_13433,N_11131);
or U17065 (N_17065,N_11553,N_13462);
nor U17066 (N_17066,N_12997,N_14434);
and U17067 (N_17067,N_14279,N_13899);
or U17068 (N_17068,N_11827,N_11520);
xor U17069 (N_17069,N_11936,N_12639);
or U17070 (N_17070,N_14129,N_14328);
nor U17071 (N_17071,N_14893,N_14414);
and U17072 (N_17072,N_13003,N_13391);
or U17073 (N_17073,N_14710,N_13931);
xor U17074 (N_17074,N_10663,N_14152);
xnor U17075 (N_17075,N_14892,N_14614);
nand U17076 (N_17076,N_13891,N_14999);
xor U17077 (N_17077,N_10309,N_14792);
xnor U17078 (N_17078,N_11269,N_14992);
xor U17079 (N_17079,N_11652,N_10830);
nor U17080 (N_17080,N_10455,N_11829);
nand U17081 (N_17081,N_14291,N_11559);
and U17082 (N_17082,N_10126,N_11708);
nor U17083 (N_17083,N_10484,N_14199);
and U17084 (N_17084,N_13588,N_12098);
or U17085 (N_17085,N_12173,N_13623);
xnor U17086 (N_17086,N_10100,N_12989);
nand U17087 (N_17087,N_14178,N_10662);
xor U17088 (N_17088,N_11903,N_12356);
or U17089 (N_17089,N_14511,N_11702);
or U17090 (N_17090,N_12362,N_10379);
xnor U17091 (N_17091,N_10719,N_14173);
or U17092 (N_17092,N_12668,N_14942);
nor U17093 (N_17093,N_10905,N_12135);
nor U17094 (N_17094,N_13876,N_12607);
or U17095 (N_17095,N_10313,N_11975);
and U17096 (N_17096,N_12025,N_14504);
nand U17097 (N_17097,N_13761,N_11679);
nor U17098 (N_17098,N_10502,N_12901);
xnor U17099 (N_17099,N_10939,N_11029);
and U17100 (N_17100,N_10907,N_14281);
nand U17101 (N_17101,N_10511,N_11627);
nand U17102 (N_17102,N_11332,N_11670);
nor U17103 (N_17103,N_14301,N_12172);
or U17104 (N_17104,N_14057,N_13172);
nor U17105 (N_17105,N_10012,N_11740);
xnor U17106 (N_17106,N_10021,N_14463);
nand U17107 (N_17107,N_14056,N_12690);
and U17108 (N_17108,N_13403,N_13057);
nor U17109 (N_17109,N_12739,N_10713);
xor U17110 (N_17110,N_13274,N_14599);
or U17111 (N_17111,N_11845,N_10569);
nor U17112 (N_17112,N_12983,N_11339);
nor U17113 (N_17113,N_13933,N_12252);
nor U17114 (N_17114,N_11306,N_11929);
or U17115 (N_17115,N_11184,N_14065);
or U17116 (N_17116,N_10578,N_10249);
xor U17117 (N_17117,N_12124,N_12282);
nand U17118 (N_17118,N_11722,N_11665);
or U17119 (N_17119,N_14794,N_13083);
and U17120 (N_17120,N_11208,N_10613);
or U17121 (N_17121,N_10650,N_13527);
nand U17122 (N_17122,N_10037,N_13272);
nor U17123 (N_17123,N_13526,N_10936);
nand U17124 (N_17124,N_11792,N_13658);
or U17125 (N_17125,N_11159,N_14097);
or U17126 (N_17126,N_13744,N_10178);
or U17127 (N_17127,N_10108,N_14001);
xor U17128 (N_17128,N_11135,N_11478);
or U17129 (N_17129,N_12345,N_11600);
xor U17130 (N_17130,N_13954,N_14633);
and U17131 (N_17131,N_10846,N_12737);
nor U17132 (N_17132,N_14564,N_11067);
nand U17133 (N_17133,N_14272,N_10233);
or U17134 (N_17134,N_14253,N_14282);
nor U17135 (N_17135,N_10691,N_10616);
or U17136 (N_17136,N_14574,N_14592);
or U17137 (N_17137,N_13324,N_12064);
or U17138 (N_17138,N_11504,N_10117);
and U17139 (N_17139,N_14964,N_14048);
nor U17140 (N_17140,N_13371,N_13689);
or U17141 (N_17141,N_11498,N_10094);
xnor U17142 (N_17142,N_12225,N_10306);
and U17143 (N_17143,N_14354,N_12473);
nor U17144 (N_17144,N_13377,N_12682);
nand U17145 (N_17145,N_14181,N_12571);
nor U17146 (N_17146,N_10326,N_11739);
and U17147 (N_17147,N_14071,N_11552);
nor U17148 (N_17148,N_13009,N_14594);
nor U17149 (N_17149,N_10927,N_12260);
nand U17150 (N_17150,N_13543,N_11873);
nand U17151 (N_17151,N_11304,N_10188);
nor U17152 (N_17152,N_12511,N_12235);
or U17153 (N_17153,N_14454,N_11550);
nand U17154 (N_17154,N_11375,N_13917);
or U17155 (N_17155,N_10656,N_14699);
nand U17156 (N_17156,N_12015,N_13515);
xor U17157 (N_17157,N_11542,N_10467);
nand U17158 (N_17158,N_11316,N_11890);
xnor U17159 (N_17159,N_11991,N_13102);
nand U17160 (N_17160,N_11926,N_14802);
nor U17161 (N_17161,N_10385,N_10162);
or U17162 (N_17162,N_14156,N_13585);
and U17163 (N_17163,N_11488,N_10348);
nor U17164 (N_17164,N_13215,N_14856);
xnor U17165 (N_17165,N_10323,N_12080);
and U17166 (N_17166,N_14096,N_11710);
and U17167 (N_17167,N_11489,N_13739);
nor U17168 (N_17168,N_14799,N_12268);
xnor U17169 (N_17169,N_13157,N_12116);
nor U17170 (N_17170,N_11828,N_11818);
and U17171 (N_17171,N_14453,N_14022);
and U17172 (N_17172,N_14886,N_13605);
xor U17173 (N_17173,N_12517,N_12306);
and U17174 (N_17174,N_12671,N_10272);
or U17175 (N_17175,N_11825,N_12250);
or U17176 (N_17176,N_13168,N_10004);
and U17177 (N_17177,N_12723,N_12750);
nor U17178 (N_17178,N_11266,N_11400);
and U17179 (N_17179,N_13022,N_14987);
and U17180 (N_17180,N_13913,N_14313);
nand U17181 (N_17181,N_13504,N_11128);
and U17182 (N_17182,N_13343,N_13697);
nor U17183 (N_17183,N_12621,N_11721);
or U17184 (N_17184,N_14687,N_11660);
nand U17185 (N_17185,N_13943,N_14819);
nand U17186 (N_17186,N_14116,N_13496);
xor U17187 (N_17187,N_14776,N_12947);
nor U17188 (N_17188,N_11527,N_14923);
and U17189 (N_17189,N_11949,N_13479);
nor U17190 (N_17190,N_13695,N_12680);
nand U17191 (N_17191,N_14868,N_14495);
or U17192 (N_17192,N_11617,N_13213);
and U17193 (N_17193,N_11972,N_13109);
or U17194 (N_17194,N_11719,N_14717);
nor U17195 (N_17195,N_14123,N_12876);
xor U17196 (N_17196,N_10692,N_14977);
and U17197 (N_17197,N_13967,N_12297);
or U17198 (N_17198,N_11954,N_14327);
or U17199 (N_17199,N_11349,N_10716);
nand U17200 (N_17200,N_10371,N_14623);
nand U17201 (N_17201,N_13361,N_14157);
and U17202 (N_17202,N_13548,N_11224);
xor U17203 (N_17203,N_13222,N_11515);
nand U17204 (N_17204,N_10040,N_11727);
nand U17205 (N_17205,N_11806,N_13567);
nor U17206 (N_17206,N_12516,N_11525);
nor U17207 (N_17207,N_11284,N_13584);
nor U17208 (N_17208,N_12011,N_11433);
nand U17209 (N_17209,N_13219,N_14246);
nor U17210 (N_17210,N_10331,N_13508);
or U17211 (N_17211,N_12996,N_10602);
or U17212 (N_17212,N_13576,N_12961);
xor U17213 (N_17213,N_12786,N_12185);
nor U17214 (N_17214,N_10508,N_12434);
nor U17215 (N_17215,N_14516,N_10570);
and U17216 (N_17216,N_10783,N_13797);
xor U17217 (N_17217,N_13124,N_12175);
nor U17218 (N_17218,N_10251,N_13419);
or U17219 (N_17219,N_14539,N_10823);
or U17220 (N_17220,N_13121,N_11869);
xor U17221 (N_17221,N_14377,N_11199);
xnor U17222 (N_17222,N_13615,N_11729);
or U17223 (N_17223,N_14505,N_13356);
and U17224 (N_17224,N_14063,N_12341);
or U17225 (N_17225,N_13595,N_13482);
or U17226 (N_17226,N_14659,N_13923);
or U17227 (N_17227,N_10902,N_13061);
and U17228 (N_17228,N_13802,N_13443);
or U17229 (N_17229,N_12634,N_12284);
xor U17230 (N_17230,N_12688,N_13551);
nand U17231 (N_17231,N_14440,N_11111);
and U17232 (N_17232,N_13731,N_12900);
and U17233 (N_17233,N_10746,N_10599);
nand U17234 (N_17234,N_14971,N_14509);
xnor U17235 (N_17235,N_10050,N_12862);
or U17236 (N_17236,N_12725,N_14501);
or U17237 (N_17237,N_13463,N_11904);
nor U17238 (N_17238,N_13848,N_13287);
or U17239 (N_17239,N_14140,N_13649);
nor U17240 (N_17240,N_14407,N_12523);
nand U17241 (N_17241,N_13350,N_11988);
or U17242 (N_17242,N_11279,N_12211);
xor U17243 (N_17243,N_13885,N_13792);
and U17244 (N_17244,N_13500,N_11646);
nor U17245 (N_17245,N_14855,N_14566);
nand U17246 (N_17246,N_11360,N_12934);
nand U17247 (N_17247,N_10353,N_14196);
nand U17248 (N_17248,N_11992,N_11230);
nand U17249 (N_17249,N_12361,N_11782);
or U17250 (N_17250,N_10584,N_12066);
xnor U17251 (N_17251,N_13858,N_12158);
xor U17252 (N_17252,N_13144,N_10328);
and U17253 (N_17253,N_11406,N_12518);
xor U17254 (N_17254,N_14323,N_13289);
nand U17255 (N_17255,N_10935,N_14032);
nand U17256 (N_17256,N_11020,N_10781);
or U17257 (N_17257,N_12761,N_11495);
or U17258 (N_17258,N_11049,N_13063);
and U17259 (N_17259,N_14482,N_11296);
and U17260 (N_17260,N_11889,N_12156);
xor U17261 (N_17261,N_14466,N_10167);
or U17262 (N_17262,N_12968,N_11397);
nor U17263 (N_17263,N_12751,N_10926);
or U17264 (N_17264,N_10843,N_12530);
or U17265 (N_17265,N_10626,N_13590);
and U17266 (N_17266,N_13081,N_14690);
and U17267 (N_17267,N_13446,N_10496);
and U17268 (N_17268,N_10845,N_14002);
or U17269 (N_17269,N_13040,N_12990);
nor U17270 (N_17270,N_14401,N_13824);
and U17271 (N_17271,N_10159,N_11290);
xnor U17272 (N_17272,N_12093,N_13138);
nor U17273 (N_17273,N_13492,N_11211);
nor U17274 (N_17274,N_13431,N_13080);
and U17275 (N_17275,N_13445,N_12117);
xnor U17276 (N_17276,N_10795,N_10954);
nand U17277 (N_17277,N_13872,N_12880);
xor U17278 (N_17278,N_10675,N_12006);
nand U17279 (N_17279,N_10247,N_12832);
xor U17280 (N_17280,N_10955,N_10472);
nand U17281 (N_17281,N_12515,N_11026);
nand U17282 (N_17282,N_12329,N_10541);
nor U17283 (N_17283,N_11812,N_10377);
nand U17284 (N_17284,N_12713,N_10906);
nor U17285 (N_17285,N_10683,N_10189);
or U17286 (N_17286,N_11268,N_14786);
and U17287 (N_17287,N_10463,N_13973);
or U17288 (N_17288,N_10096,N_14244);
and U17289 (N_17289,N_11030,N_11961);
xnor U17290 (N_17290,N_13412,N_13296);
xor U17291 (N_17291,N_12272,N_10585);
nand U17292 (N_17292,N_11885,N_14996);
or U17293 (N_17293,N_10443,N_12307);
nor U17294 (N_17294,N_14738,N_13682);
xor U17295 (N_17295,N_10912,N_13721);
nor U17296 (N_17296,N_14730,N_10081);
xor U17297 (N_17297,N_12383,N_11173);
and U17298 (N_17298,N_14468,N_12749);
nand U17299 (N_17299,N_11465,N_14983);
and U17300 (N_17300,N_11374,N_14640);
xor U17301 (N_17301,N_13646,N_13209);
xor U17302 (N_17302,N_10800,N_13163);
nand U17303 (N_17303,N_12860,N_11717);
and U17304 (N_17304,N_13730,N_13535);
or U17305 (N_17305,N_11560,N_12824);
nand U17306 (N_17306,N_11427,N_10512);
and U17307 (N_17307,N_10863,N_12371);
xor U17308 (N_17308,N_14102,N_12493);
nand U17309 (N_17309,N_13680,N_10209);
or U17310 (N_17310,N_10068,N_11716);
nor U17311 (N_17311,N_10053,N_14139);
xor U17312 (N_17312,N_11333,N_12665);
nor U17313 (N_17313,N_13113,N_10190);
and U17314 (N_17314,N_12789,N_13046);
nor U17315 (N_17315,N_10093,N_10157);
or U17316 (N_17316,N_13717,N_14230);
or U17317 (N_17317,N_11523,N_12732);
and U17318 (N_17318,N_12468,N_13892);
xor U17319 (N_17319,N_13686,N_11106);
nor U17320 (N_17320,N_12675,N_14256);
nand U17321 (N_17321,N_14351,N_14641);
xnor U17322 (N_17322,N_13974,N_10535);
nand U17323 (N_17323,N_14649,N_14026);
and U17324 (N_17324,N_14568,N_13223);
and U17325 (N_17325,N_11987,N_11112);
or U17326 (N_17326,N_10346,N_11327);
nor U17327 (N_17327,N_13006,N_12396);
nor U17328 (N_17328,N_14704,N_13306);
or U17329 (N_17329,N_12293,N_10349);
nand U17330 (N_17330,N_11541,N_12604);
nor U17331 (N_17331,N_13362,N_14448);
nor U17332 (N_17332,N_12425,N_10759);
xor U17333 (N_17333,N_12187,N_11824);
xnor U17334 (N_17334,N_12215,N_13177);
nor U17335 (N_17335,N_10469,N_14376);
or U17336 (N_17336,N_10896,N_10684);
and U17337 (N_17337,N_10790,N_14186);
and U17338 (N_17338,N_13702,N_12729);
nor U17339 (N_17339,N_12244,N_13871);
or U17340 (N_17340,N_12692,N_12551);
xnor U17341 (N_17341,N_14721,N_10145);
and U17342 (N_17342,N_11149,N_14409);
xor U17343 (N_17343,N_12089,N_13794);
xnor U17344 (N_17344,N_10354,N_14015);
nor U17345 (N_17345,N_12958,N_14936);
and U17346 (N_17346,N_10319,N_14949);
and U17347 (N_17347,N_11345,N_10735);
xnor U17348 (N_17348,N_10062,N_12825);
or U17349 (N_17349,N_11849,N_13678);
and U17350 (N_17350,N_11785,N_10853);
nand U17351 (N_17351,N_13918,N_10963);
xnor U17352 (N_17352,N_11257,N_11060);
nand U17353 (N_17353,N_12423,N_10196);
xor U17354 (N_17354,N_10561,N_14415);
nor U17355 (N_17355,N_14042,N_14940);
or U17356 (N_17356,N_13573,N_13626);
or U17357 (N_17357,N_11031,N_14514);
or U17358 (N_17358,N_13574,N_14270);
nand U17359 (N_17359,N_10411,N_14044);
nand U17360 (N_17360,N_12319,N_10092);
nand U17361 (N_17361,N_12369,N_11209);
xor U17362 (N_17362,N_12811,N_12163);
or U17363 (N_17363,N_11513,N_12288);
nand U17364 (N_17364,N_11470,N_14905);
nor U17365 (N_17365,N_13176,N_11133);
or U17366 (N_17366,N_11589,N_14846);
nor U17367 (N_17367,N_12129,N_12206);
nand U17368 (N_17368,N_13444,N_12606);
nand U17369 (N_17369,N_12560,N_12216);
nand U17370 (N_17370,N_14131,N_12846);
or U17371 (N_17371,N_13193,N_13271);
nor U17372 (N_17372,N_14748,N_14080);
and U17373 (N_17373,N_14534,N_14252);
xor U17374 (N_17374,N_13112,N_10723);
xnor U17375 (N_17375,N_10285,N_11492);
xor U17376 (N_17376,N_13349,N_14752);
xor U17377 (N_17377,N_10276,N_12886);
xnor U17378 (N_17378,N_11605,N_14429);
nand U17379 (N_17379,N_13366,N_12410);
xnor U17380 (N_17380,N_13988,N_12335);
nand U17381 (N_17381,N_10966,N_10580);
xor U17382 (N_17382,N_12458,N_11493);
or U17383 (N_17383,N_14777,N_12663);
and U17384 (N_17384,N_12827,N_12705);
or U17385 (N_17385,N_10495,N_12654);
nand U17386 (N_17386,N_10559,N_11420);
xnor U17387 (N_17387,N_14098,N_11191);
and U17388 (N_17388,N_10427,N_11367);
nor U17389 (N_17389,N_10601,N_11411);
nor U17390 (N_17390,N_11786,N_10296);
xor U17391 (N_17391,N_10327,N_11763);
and U17392 (N_17392,N_12099,N_13410);
nor U17393 (N_17393,N_12243,N_12265);
xor U17394 (N_17394,N_11963,N_12936);
or U17395 (N_17395,N_14484,N_14013);
nand U17396 (N_17396,N_10333,N_14049);
or U17397 (N_17397,N_14340,N_14561);
or U17398 (N_17398,N_13867,N_12090);
nand U17399 (N_17399,N_14195,N_11412);
nand U17400 (N_17400,N_11502,N_14134);
nand U17401 (N_17401,N_11166,N_10215);
or U17402 (N_17402,N_10432,N_10820);
or U17403 (N_17403,N_12576,N_12494);
xnor U17404 (N_17404,N_14118,N_14672);
nand U17405 (N_17405,N_10576,N_12195);
or U17406 (N_17406,N_10217,N_12237);
nand U17407 (N_17407,N_14956,N_13214);
or U17408 (N_17408,N_13182,N_12645);
xor U17409 (N_17409,N_14806,N_10464);
nor U17410 (N_17410,N_14067,N_12310);
nor U17411 (N_17411,N_14076,N_14556);
and U17412 (N_17412,N_11267,N_14773);
or U17413 (N_17413,N_14805,N_14795);
xor U17414 (N_17414,N_10634,N_14489);
nor U17415 (N_17415,N_13544,N_11396);
nand U17416 (N_17416,N_11081,N_11450);
or U17417 (N_17417,N_10873,N_11121);
nand U17418 (N_17418,N_12200,N_10619);
or U17419 (N_17419,N_14314,N_11712);
nand U17420 (N_17420,N_11532,N_11072);
and U17421 (N_17421,N_10404,N_10337);
nor U17422 (N_17422,N_14771,N_10378);
or U17423 (N_17423,N_13826,N_11481);
or U17424 (N_17424,N_14359,N_11271);
xor U17425 (N_17425,N_12780,N_11448);
nor U17426 (N_17426,N_10086,N_11186);
nand U17427 (N_17427,N_11754,N_13220);
nand U17428 (N_17428,N_14702,N_11529);
and U17429 (N_17429,N_12546,N_14020);
xor U17430 (N_17430,N_10356,N_11497);
nor U17431 (N_17431,N_14193,N_10440);
xnor U17432 (N_17432,N_11657,N_11896);
xnor U17433 (N_17433,N_11462,N_10474);
nor U17434 (N_17434,N_13805,N_13185);
or U17435 (N_17435,N_12559,N_14023);
and U17436 (N_17436,N_14938,N_13536);
or U17437 (N_17437,N_10509,N_14233);
nor U17438 (N_17438,N_12744,N_10340);
nor U17439 (N_17439,N_10383,N_11147);
xor U17440 (N_17440,N_14066,N_13472);
xor U17441 (N_17441,N_13675,N_12942);
nand U17442 (N_17442,N_13570,N_12804);
nor U17443 (N_17443,N_13059,N_11344);
nand U17444 (N_17444,N_12731,N_14424);
nor U17445 (N_17445,N_10537,N_13814);
nand U17446 (N_17446,N_11728,N_12612);
nor U17447 (N_17447,N_13898,N_10199);
and U17448 (N_17448,N_11001,N_13547);
or U17449 (N_17449,N_14143,N_14223);
and U17450 (N_17450,N_12887,N_11219);
nand U17451 (N_17451,N_11980,N_12189);
xnor U17452 (N_17452,N_12354,N_14671);
nor U17453 (N_17453,N_11024,N_14603);
xnor U17454 (N_17454,N_12981,N_14836);
nand U17455 (N_17455,N_11805,N_13128);
nand U17456 (N_17456,N_10431,N_10436);
xnor U17457 (N_17457,N_14303,N_10751);
xor U17458 (N_17458,N_10997,N_10633);
and U17459 (N_17459,N_13559,N_14387);
nor U17460 (N_17460,N_12289,N_13870);
and U17461 (N_17461,N_10007,N_13557);
and U17462 (N_17462,N_11598,N_10943);
nand U17463 (N_17463,N_11635,N_14668);
or U17464 (N_17464,N_10334,N_12197);
and U17465 (N_17465,N_12964,N_13782);
or U17466 (N_17466,N_14715,N_12554);
and U17467 (N_17467,N_13908,N_10514);
nor U17468 (N_17468,N_10224,N_11675);
nand U17469 (N_17469,N_11964,N_12531);
xor U17470 (N_17470,N_14190,N_14356);
or U17471 (N_17471,N_11273,N_14037);
or U17472 (N_17472,N_11435,N_11342);
nor U17473 (N_17473,N_12907,N_11852);
or U17474 (N_17474,N_10426,N_12693);
xor U17475 (N_17475,N_14330,N_13263);
nand U17476 (N_17476,N_10933,N_11126);
or U17477 (N_17477,N_10620,N_14676);
xor U17478 (N_17478,N_13370,N_12995);
and U17479 (N_17479,N_12367,N_12923);
xor U17480 (N_17480,N_12736,N_13810);
nor U17481 (N_17481,N_13095,N_11202);
or U17482 (N_17482,N_12911,N_12799);
xor U17483 (N_17483,N_14213,N_12415);
xor U17484 (N_17484,N_13019,N_12672);
or U17485 (N_17485,N_13183,N_12773);
and U17486 (N_17486,N_10526,N_11699);
and U17487 (N_17487,N_14955,N_14457);
or U17488 (N_17488,N_12283,N_10446);
nand U17489 (N_17489,N_10608,N_11959);
xnor U17490 (N_17490,N_11119,N_14540);
or U17491 (N_17491,N_10574,N_12666);
or U17492 (N_17492,N_13253,N_13643);
or U17493 (N_17493,N_12381,N_10028);
nor U17494 (N_17494,N_10183,N_13328);
nor U17495 (N_17495,N_11463,N_13594);
nand U17496 (N_17496,N_11263,N_11864);
and U17497 (N_17497,N_14382,N_14528);
xor U17498 (N_17498,N_13008,N_10988);
xor U17499 (N_17499,N_12009,N_10437);
xnor U17500 (N_17500,N_14989,N_14855);
nand U17501 (N_17501,N_14177,N_13423);
xnor U17502 (N_17502,N_14439,N_14381);
and U17503 (N_17503,N_10164,N_11641);
nor U17504 (N_17504,N_10381,N_10821);
nand U17505 (N_17505,N_14710,N_14037);
or U17506 (N_17506,N_14504,N_10168);
and U17507 (N_17507,N_14255,N_13623);
xor U17508 (N_17508,N_11645,N_13610);
and U17509 (N_17509,N_11673,N_12767);
and U17510 (N_17510,N_13521,N_11755);
nor U17511 (N_17511,N_10599,N_12671);
nor U17512 (N_17512,N_11372,N_11231);
nor U17513 (N_17513,N_13023,N_13076);
nor U17514 (N_17514,N_13386,N_11282);
nor U17515 (N_17515,N_12931,N_11732);
nand U17516 (N_17516,N_11511,N_10117);
and U17517 (N_17517,N_10215,N_14501);
nand U17518 (N_17518,N_12084,N_13090);
and U17519 (N_17519,N_11829,N_14253);
nand U17520 (N_17520,N_10827,N_14923);
nand U17521 (N_17521,N_14470,N_11490);
or U17522 (N_17522,N_13874,N_11978);
or U17523 (N_17523,N_10445,N_14525);
nand U17524 (N_17524,N_10675,N_11773);
xor U17525 (N_17525,N_14937,N_14319);
or U17526 (N_17526,N_12132,N_14908);
nand U17527 (N_17527,N_12762,N_11715);
or U17528 (N_17528,N_10985,N_10809);
nand U17529 (N_17529,N_12571,N_13698);
nand U17530 (N_17530,N_12245,N_12861);
nand U17531 (N_17531,N_13229,N_13633);
and U17532 (N_17532,N_10246,N_13342);
and U17533 (N_17533,N_12824,N_13414);
nor U17534 (N_17534,N_10912,N_13253);
or U17535 (N_17535,N_12538,N_11156);
nor U17536 (N_17536,N_14655,N_11956);
or U17537 (N_17537,N_11154,N_11790);
nor U17538 (N_17538,N_10698,N_10141);
nand U17539 (N_17539,N_12104,N_12373);
nand U17540 (N_17540,N_12173,N_12957);
xnor U17541 (N_17541,N_11209,N_10988);
or U17542 (N_17542,N_14847,N_12800);
and U17543 (N_17543,N_14862,N_14483);
or U17544 (N_17544,N_10775,N_11352);
nor U17545 (N_17545,N_13494,N_13903);
nor U17546 (N_17546,N_13578,N_10037);
or U17547 (N_17547,N_12549,N_11647);
nand U17548 (N_17548,N_12336,N_12770);
xor U17549 (N_17549,N_14362,N_12187);
xor U17550 (N_17550,N_13423,N_10610);
or U17551 (N_17551,N_12732,N_14429);
nand U17552 (N_17552,N_10913,N_12616);
and U17553 (N_17553,N_11837,N_13466);
xor U17554 (N_17554,N_10387,N_13541);
or U17555 (N_17555,N_12766,N_14022);
xnor U17556 (N_17556,N_14679,N_10589);
xnor U17557 (N_17557,N_10249,N_11596);
nand U17558 (N_17558,N_13843,N_13334);
and U17559 (N_17559,N_12143,N_12505);
or U17560 (N_17560,N_12412,N_10549);
nor U17561 (N_17561,N_11725,N_14047);
nand U17562 (N_17562,N_14972,N_12929);
or U17563 (N_17563,N_11045,N_10601);
nor U17564 (N_17564,N_10090,N_14862);
xnor U17565 (N_17565,N_12001,N_14054);
and U17566 (N_17566,N_11276,N_10906);
or U17567 (N_17567,N_10935,N_10544);
nand U17568 (N_17568,N_10127,N_13872);
and U17569 (N_17569,N_13527,N_13390);
and U17570 (N_17570,N_10733,N_10022);
nand U17571 (N_17571,N_10341,N_14563);
nand U17572 (N_17572,N_14293,N_10679);
nand U17573 (N_17573,N_13877,N_12131);
nand U17574 (N_17574,N_14332,N_12473);
nand U17575 (N_17575,N_10233,N_11502);
and U17576 (N_17576,N_11872,N_12688);
nor U17577 (N_17577,N_12150,N_12157);
nand U17578 (N_17578,N_13150,N_14249);
nor U17579 (N_17579,N_12231,N_12010);
nand U17580 (N_17580,N_13326,N_10578);
nand U17581 (N_17581,N_10989,N_13437);
nor U17582 (N_17582,N_11430,N_12839);
xor U17583 (N_17583,N_13092,N_10515);
or U17584 (N_17584,N_13219,N_12989);
and U17585 (N_17585,N_11184,N_12762);
xor U17586 (N_17586,N_10123,N_12644);
nand U17587 (N_17587,N_14122,N_13820);
nor U17588 (N_17588,N_14365,N_13279);
xnor U17589 (N_17589,N_11182,N_13623);
nor U17590 (N_17590,N_12895,N_11734);
xor U17591 (N_17591,N_12839,N_14275);
and U17592 (N_17592,N_10503,N_13154);
or U17593 (N_17593,N_11626,N_14103);
nor U17594 (N_17594,N_14365,N_10597);
or U17595 (N_17595,N_14746,N_11694);
xnor U17596 (N_17596,N_10067,N_10848);
or U17597 (N_17597,N_13509,N_12515);
nand U17598 (N_17598,N_12976,N_10907);
or U17599 (N_17599,N_11619,N_14657);
nand U17600 (N_17600,N_12891,N_10752);
nand U17601 (N_17601,N_14256,N_12248);
nor U17602 (N_17602,N_14109,N_10627);
or U17603 (N_17603,N_10348,N_11188);
nor U17604 (N_17604,N_11545,N_11360);
or U17605 (N_17605,N_12732,N_14912);
and U17606 (N_17606,N_12281,N_13658);
and U17607 (N_17607,N_11106,N_13380);
and U17608 (N_17608,N_10441,N_14977);
xor U17609 (N_17609,N_13599,N_12191);
xor U17610 (N_17610,N_14418,N_13848);
xor U17611 (N_17611,N_10902,N_10883);
xnor U17612 (N_17612,N_14468,N_12737);
and U17613 (N_17613,N_12797,N_13860);
or U17614 (N_17614,N_12109,N_14289);
or U17615 (N_17615,N_10490,N_12107);
or U17616 (N_17616,N_13922,N_11223);
nand U17617 (N_17617,N_14968,N_11670);
and U17618 (N_17618,N_14862,N_14188);
or U17619 (N_17619,N_10923,N_10397);
xnor U17620 (N_17620,N_12268,N_11494);
and U17621 (N_17621,N_12161,N_11378);
and U17622 (N_17622,N_13424,N_14211);
xor U17623 (N_17623,N_13511,N_10295);
nand U17624 (N_17624,N_10138,N_10205);
xor U17625 (N_17625,N_13408,N_13748);
nand U17626 (N_17626,N_11096,N_14578);
nor U17627 (N_17627,N_10834,N_13797);
xor U17628 (N_17628,N_11554,N_12778);
nor U17629 (N_17629,N_10500,N_10060);
nand U17630 (N_17630,N_13297,N_11471);
nand U17631 (N_17631,N_12862,N_14399);
xnor U17632 (N_17632,N_11647,N_14469);
nand U17633 (N_17633,N_14241,N_10031);
nor U17634 (N_17634,N_12162,N_10053);
xnor U17635 (N_17635,N_12106,N_14252);
xnor U17636 (N_17636,N_12085,N_13401);
and U17637 (N_17637,N_10947,N_12666);
xnor U17638 (N_17638,N_13555,N_10319);
nor U17639 (N_17639,N_10098,N_14159);
nor U17640 (N_17640,N_12827,N_13022);
or U17641 (N_17641,N_14205,N_13177);
or U17642 (N_17642,N_10361,N_14373);
nand U17643 (N_17643,N_11057,N_14493);
and U17644 (N_17644,N_11745,N_13551);
xnor U17645 (N_17645,N_11632,N_14191);
nor U17646 (N_17646,N_14871,N_14068);
and U17647 (N_17647,N_11665,N_14130);
xnor U17648 (N_17648,N_14767,N_13319);
and U17649 (N_17649,N_10415,N_10699);
nor U17650 (N_17650,N_14876,N_12853);
nor U17651 (N_17651,N_14534,N_12990);
xor U17652 (N_17652,N_14216,N_10996);
and U17653 (N_17653,N_10134,N_13904);
xnor U17654 (N_17654,N_10339,N_14711);
and U17655 (N_17655,N_10831,N_12905);
nor U17656 (N_17656,N_14896,N_14887);
nand U17657 (N_17657,N_13525,N_14228);
nor U17658 (N_17658,N_10531,N_12337);
and U17659 (N_17659,N_14564,N_10591);
nand U17660 (N_17660,N_11769,N_14744);
and U17661 (N_17661,N_14739,N_10877);
or U17662 (N_17662,N_11408,N_12511);
nand U17663 (N_17663,N_14118,N_14762);
nand U17664 (N_17664,N_12975,N_12600);
nand U17665 (N_17665,N_11263,N_13375);
xnor U17666 (N_17666,N_11421,N_13412);
nand U17667 (N_17667,N_10510,N_10464);
nor U17668 (N_17668,N_13542,N_13444);
nand U17669 (N_17669,N_10443,N_13232);
or U17670 (N_17670,N_10856,N_11809);
and U17671 (N_17671,N_11043,N_14701);
nor U17672 (N_17672,N_12364,N_11804);
nor U17673 (N_17673,N_10003,N_14385);
xor U17674 (N_17674,N_13778,N_13398);
nor U17675 (N_17675,N_10334,N_11537);
or U17676 (N_17676,N_12747,N_10598);
nor U17677 (N_17677,N_14409,N_11059);
or U17678 (N_17678,N_12528,N_11562);
nor U17679 (N_17679,N_12102,N_14308);
nor U17680 (N_17680,N_11626,N_13926);
nand U17681 (N_17681,N_10401,N_11290);
xnor U17682 (N_17682,N_12661,N_10287);
or U17683 (N_17683,N_12182,N_11756);
xnor U17684 (N_17684,N_13732,N_14930);
and U17685 (N_17685,N_10091,N_10811);
and U17686 (N_17686,N_11983,N_12796);
and U17687 (N_17687,N_14651,N_11352);
and U17688 (N_17688,N_14632,N_11645);
nor U17689 (N_17689,N_10993,N_11119);
and U17690 (N_17690,N_13299,N_14378);
nand U17691 (N_17691,N_10172,N_10188);
nor U17692 (N_17692,N_11566,N_14434);
or U17693 (N_17693,N_11741,N_12110);
nor U17694 (N_17694,N_14247,N_14552);
and U17695 (N_17695,N_13094,N_14492);
or U17696 (N_17696,N_11274,N_12570);
or U17697 (N_17697,N_14649,N_11114);
and U17698 (N_17698,N_14298,N_12939);
nand U17699 (N_17699,N_13429,N_13148);
nand U17700 (N_17700,N_13064,N_14321);
or U17701 (N_17701,N_10784,N_11212);
nand U17702 (N_17702,N_11733,N_13547);
nor U17703 (N_17703,N_14982,N_13235);
nor U17704 (N_17704,N_14600,N_14964);
or U17705 (N_17705,N_14405,N_12263);
or U17706 (N_17706,N_10956,N_12487);
nor U17707 (N_17707,N_12653,N_13162);
nand U17708 (N_17708,N_13290,N_11273);
nand U17709 (N_17709,N_11619,N_11603);
nand U17710 (N_17710,N_12974,N_13559);
and U17711 (N_17711,N_10252,N_13289);
nor U17712 (N_17712,N_11593,N_11205);
or U17713 (N_17713,N_12288,N_14884);
and U17714 (N_17714,N_13069,N_13252);
or U17715 (N_17715,N_14973,N_14135);
xnor U17716 (N_17716,N_13071,N_12092);
nor U17717 (N_17717,N_14501,N_14113);
nand U17718 (N_17718,N_12916,N_11964);
and U17719 (N_17719,N_13608,N_14565);
and U17720 (N_17720,N_14425,N_12694);
nor U17721 (N_17721,N_10221,N_13711);
nor U17722 (N_17722,N_12004,N_12081);
and U17723 (N_17723,N_11279,N_14989);
or U17724 (N_17724,N_10442,N_13010);
or U17725 (N_17725,N_10368,N_12777);
and U17726 (N_17726,N_11437,N_12902);
or U17727 (N_17727,N_13860,N_11308);
or U17728 (N_17728,N_11679,N_12616);
xnor U17729 (N_17729,N_10336,N_14822);
and U17730 (N_17730,N_14198,N_10778);
or U17731 (N_17731,N_10317,N_10863);
or U17732 (N_17732,N_11663,N_11765);
nor U17733 (N_17733,N_11007,N_11168);
nand U17734 (N_17734,N_11191,N_14707);
xor U17735 (N_17735,N_11775,N_14617);
or U17736 (N_17736,N_11424,N_10273);
or U17737 (N_17737,N_14040,N_12894);
nor U17738 (N_17738,N_10565,N_14680);
nor U17739 (N_17739,N_13522,N_12179);
nor U17740 (N_17740,N_12104,N_10979);
xor U17741 (N_17741,N_13810,N_10256);
and U17742 (N_17742,N_11268,N_14847);
nand U17743 (N_17743,N_10544,N_14846);
nor U17744 (N_17744,N_12539,N_10244);
nand U17745 (N_17745,N_10894,N_13819);
xnor U17746 (N_17746,N_11764,N_10148);
and U17747 (N_17747,N_13162,N_12333);
or U17748 (N_17748,N_13419,N_11714);
nor U17749 (N_17749,N_10721,N_12666);
nand U17750 (N_17750,N_14488,N_11171);
nand U17751 (N_17751,N_12041,N_11512);
and U17752 (N_17752,N_13383,N_14560);
or U17753 (N_17753,N_11303,N_13624);
xnor U17754 (N_17754,N_10067,N_13706);
xor U17755 (N_17755,N_10055,N_11404);
nor U17756 (N_17756,N_13800,N_14555);
xnor U17757 (N_17757,N_12099,N_13982);
or U17758 (N_17758,N_12930,N_11899);
nand U17759 (N_17759,N_12593,N_12863);
nand U17760 (N_17760,N_12809,N_10192);
xor U17761 (N_17761,N_10991,N_13090);
and U17762 (N_17762,N_13351,N_12758);
or U17763 (N_17763,N_11455,N_11443);
or U17764 (N_17764,N_11048,N_12897);
and U17765 (N_17765,N_13702,N_14083);
xor U17766 (N_17766,N_10104,N_13282);
and U17767 (N_17767,N_13275,N_13088);
nor U17768 (N_17768,N_12346,N_11275);
and U17769 (N_17769,N_10090,N_13781);
nand U17770 (N_17770,N_13999,N_14917);
or U17771 (N_17771,N_14825,N_14325);
nor U17772 (N_17772,N_14905,N_14798);
nor U17773 (N_17773,N_14054,N_13557);
nand U17774 (N_17774,N_13961,N_11256);
nor U17775 (N_17775,N_14606,N_12805);
and U17776 (N_17776,N_10621,N_13532);
nand U17777 (N_17777,N_12752,N_11870);
nor U17778 (N_17778,N_10335,N_13571);
xor U17779 (N_17779,N_13287,N_10896);
nand U17780 (N_17780,N_13576,N_14331);
nor U17781 (N_17781,N_13427,N_13407);
or U17782 (N_17782,N_11320,N_13812);
nor U17783 (N_17783,N_13952,N_13237);
nor U17784 (N_17784,N_12494,N_10266);
nor U17785 (N_17785,N_12665,N_14772);
nand U17786 (N_17786,N_10357,N_13286);
and U17787 (N_17787,N_13309,N_11961);
nand U17788 (N_17788,N_13099,N_13185);
and U17789 (N_17789,N_10411,N_10356);
and U17790 (N_17790,N_13408,N_10870);
nand U17791 (N_17791,N_13316,N_11804);
nor U17792 (N_17792,N_13904,N_10336);
and U17793 (N_17793,N_13506,N_11218);
xor U17794 (N_17794,N_14632,N_14584);
or U17795 (N_17795,N_12427,N_14247);
xnor U17796 (N_17796,N_11857,N_11555);
and U17797 (N_17797,N_14361,N_11554);
nor U17798 (N_17798,N_10429,N_14576);
xnor U17799 (N_17799,N_13974,N_10711);
and U17800 (N_17800,N_11677,N_13525);
xor U17801 (N_17801,N_14052,N_12676);
nor U17802 (N_17802,N_11736,N_14875);
nor U17803 (N_17803,N_14402,N_10627);
nor U17804 (N_17804,N_10904,N_10699);
nor U17805 (N_17805,N_10947,N_14570);
and U17806 (N_17806,N_10584,N_11975);
and U17807 (N_17807,N_14911,N_10946);
nor U17808 (N_17808,N_12501,N_10379);
and U17809 (N_17809,N_13647,N_14588);
nand U17810 (N_17810,N_11464,N_14806);
nand U17811 (N_17811,N_10104,N_11666);
nand U17812 (N_17812,N_13888,N_10480);
and U17813 (N_17813,N_14897,N_14601);
and U17814 (N_17814,N_14288,N_12328);
xor U17815 (N_17815,N_13012,N_12393);
or U17816 (N_17816,N_12525,N_10658);
xnor U17817 (N_17817,N_10974,N_13705);
nand U17818 (N_17818,N_13068,N_12496);
nor U17819 (N_17819,N_12011,N_13171);
nor U17820 (N_17820,N_13977,N_14603);
nand U17821 (N_17821,N_13332,N_12635);
nor U17822 (N_17822,N_10226,N_10124);
and U17823 (N_17823,N_12541,N_13267);
xnor U17824 (N_17824,N_13867,N_14509);
xor U17825 (N_17825,N_13794,N_13693);
or U17826 (N_17826,N_10779,N_11981);
nor U17827 (N_17827,N_12021,N_10557);
nand U17828 (N_17828,N_10228,N_14678);
or U17829 (N_17829,N_13434,N_13499);
xnor U17830 (N_17830,N_12049,N_10308);
nand U17831 (N_17831,N_10596,N_11699);
nor U17832 (N_17832,N_11592,N_10181);
xor U17833 (N_17833,N_12166,N_13253);
xnor U17834 (N_17834,N_13251,N_14294);
nand U17835 (N_17835,N_12012,N_10983);
and U17836 (N_17836,N_13897,N_11719);
xor U17837 (N_17837,N_10800,N_13238);
nand U17838 (N_17838,N_13996,N_12175);
nand U17839 (N_17839,N_13496,N_10992);
xor U17840 (N_17840,N_14417,N_13249);
and U17841 (N_17841,N_13190,N_11050);
nor U17842 (N_17842,N_14594,N_14719);
nor U17843 (N_17843,N_11983,N_11492);
nor U17844 (N_17844,N_11614,N_13039);
nor U17845 (N_17845,N_14406,N_12020);
and U17846 (N_17846,N_10049,N_11221);
nor U17847 (N_17847,N_11209,N_11021);
nor U17848 (N_17848,N_14171,N_11037);
and U17849 (N_17849,N_12911,N_10463);
and U17850 (N_17850,N_13328,N_14656);
nand U17851 (N_17851,N_14349,N_12351);
or U17852 (N_17852,N_13982,N_13383);
and U17853 (N_17853,N_11644,N_11673);
nor U17854 (N_17854,N_13105,N_12448);
and U17855 (N_17855,N_10807,N_14733);
nand U17856 (N_17856,N_10999,N_11190);
and U17857 (N_17857,N_10545,N_10025);
and U17858 (N_17858,N_14874,N_11637);
or U17859 (N_17859,N_11161,N_13905);
nand U17860 (N_17860,N_10596,N_14352);
nand U17861 (N_17861,N_14468,N_14692);
xor U17862 (N_17862,N_11624,N_14733);
and U17863 (N_17863,N_10788,N_10281);
and U17864 (N_17864,N_10352,N_13111);
xor U17865 (N_17865,N_13406,N_10716);
and U17866 (N_17866,N_12759,N_10647);
or U17867 (N_17867,N_14584,N_14427);
and U17868 (N_17868,N_10525,N_11373);
xor U17869 (N_17869,N_10909,N_10220);
or U17870 (N_17870,N_13468,N_11882);
nand U17871 (N_17871,N_11541,N_11630);
xnor U17872 (N_17872,N_10836,N_12532);
nand U17873 (N_17873,N_12173,N_11315);
nor U17874 (N_17874,N_13588,N_10449);
or U17875 (N_17875,N_11395,N_13890);
and U17876 (N_17876,N_12204,N_12685);
or U17877 (N_17877,N_14873,N_13248);
xor U17878 (N_17878,N_11383,N_14965);
or U17879 (N_17879,N_10786,N_13345);
nand U17880 (N_17880,N_14221,N_10957);
xor U17881 (N_17881,N_11317,N_11561);
xnor U17882 (N_17882,N_12498,N_10020);
nor U17883 (N_17883,N_13022,N_12471);
xnor U17884 (N_17884,N_10989,N_13573);
nand U17885 (N_17885,N_14041,N_10310);
or U17886 (N_17886,N_13903,N_12910);
xnor U17887 (N_17887,N_13773,N_10151);
xnor U17888 (N_17888,N_11041,N_11443);
and U17889 (N_17889,N_11491,N_11811);
and U17890 (N_17890,N_14092,N_11617);
nand U17891 (N_17891,N_13260,N_10877);
or U17892 (N_17892,N_11394,N_12787);
or U17893 (N_17893,N_11467,N_12699);
and U17894 (N_17894,N_13868,N_14923);
or U17895 (N_17895,N_13012,N_11069);
nand U17896 (N_17896,N_10481,N_13574);
xor U17897 (N_17897,N_13551,N_13329);
xnor U17898 (N_17898,N_10745,N_11173);
nand U17899 (N_17899,N_14634,N_13003);
and U17900 (N_17900,N_11731,N_14895);
nor U17901 (N_17901,N_12365,N_14634);
nand U17902 (N_17902,N_12102,N_14901);
xor U17903 (N_17903,N_13789,N_13921);
or U17904 (N_17904,N_12236,N_12906);
or U17905 (N_17905,N_11527,N_13341);
xor U17906 (N_17906,N_10561,N_14016);
nor U17907 (N_17907,N_13887,N_11276);
and U17908 (N_17908,N_12136,N_14889);
and U17909 (N_17909,N_10860,N_14064);
nand U17910 (N_17910,N_12610,N_13915);
xor U17911 (N_17911,N_10276,N_10081);
and U17912 (N_17912,N_13261,N_14006);
nor U17913 (N_17913,N_13911,N_10891);
nor U17914 (N_17914,N_11002,N_13881);
nand U17915 (N_17915,N_11287,N_10389);
nor U17916 (N_17916,N_13102,N_14277);
or U17917 (N_17917,N_10842,N_10013);
and U17918 (N_17918,N_10080,N_14849);
nor U17919 (N_17919,N_10204,N_13139);
xnor U17920 (N_17920,N_12534,N_13374);
nor U17921 (N_17921,N_10849,N_11931);
nor U17922 (N_17922,N_11221,N_11583);
nand U17923 (N_17923,N_14575,N_11831);
nand U17924 (N_17924,N_13030,N_11109);
and U17925 (N_17925,N_13421,N_11495);
nand U17926 (N_17926,N_10551,N_10699);
nand U17927 (N_17927,N_11034,N_12869);
or U17928 (N_17928,N_13543,N_13580);
xor U17929 (N_17929,N_14457,N_12206);
nand U17930 (N_17930,N_12337,N_12575);
nor U17931 (N_17931,N_11480,N_11802);
xor U17932 (N_17932,N_11213,N_12942);
nand U17933 (N_17933,N_10966,N_12519);
nand U17934 (N_17934,N_11432,N_10341);
or U17935 (N_17935,N_14804,N_13790);
or U17936 (N_17936,N_10795,N_13230);
nor U17937 (N_17937,N_12623,N_11804);
and U17938 (N_17938,N_12661,N_13120);
or U17939 (N_17939,N_14761,N_14024);
xnor U17940 (N_17940,N_10157,N_11737);
nor U17941 (N_17941,N_10853,N_14971);
nand U17942 (N_17942,N_14629,N_12093);
nor U17943 (N_17943,N_12552,N_13645);
or U17944 (N_17944,N_10301,N_10421);
and U17945 (N_17945,N_12433,N_10402);
nand U17946 (N_17946,N_13923,N_11662);
nor U17947 (N_17947,N_13807,N_14655);
and U17948 (N_17948,N_13773,N_14501);
nor U17949 (N_17949,N_12754,N_12863);
nand U17950 (N_17950,N_14014,N_12182);
or U17951 (N_17951,N_11300,N_12704);
nor U17952 (N_17952,N_11705,N_13073);
or U17953 (N_17953,N_10948,N_10117);
nor U17954 (N_17954,N_14390,N_14812);
and U17955 (N_17955,N_10296,N_13072);
xnor U17956 (N_17956,N_10811,N_11201);
xor U17957 (N_17957,N_12754,N_11630);
and U17958 (N_17958,N_14372,N_13895);
nor U17959 (N_17959,N_11555,N_13340);
nand U17960 (N_17960,N_11587,N_14173);
nor U17961 (N_17961,N_14583,N_14638);
nand U17962 (N_17962,N_11311,N_13334);
nor U17963 (N_17963,N_14491,N_10377);
xor U17964 (N_17964,N_12088,N_13505);
nand U17965 (N_17965,N_12943,N_11671);
nand U17966 (N_17966,N_13554,N_12414);
or U17967 (N_17967,N_14464,N_10714);
xor U17968 (N_17968,N_14733,N_11133);
and U17969 (N_17969,N_13937,N_11372);
nor U17970 (N_17970,N_11511,N_12837);
or U17971 (N_17971,N_10773,N_11550);
or U17972 (N_17972,N_13649,N_14343);
nand U17973 (N_17973,N_13488,N_11230);
and U17974 (N_17974,N_11284,N_14078);
xor U17975 (N_17975,N_10816,N_13409);
nor U17976 (N_17976,N_14307,N_12135);
nand U17977 (N_17977,N_10037,N_11112);
or U17978 (N_17978,N_10987,N_11305);
or U17979 (N_17979,N_10435,N_11968);
nand U17980 (N_17980,N_10104,N_14327);
nand U17981 (N_17981,N_10101,N_10788);
nand U17982 (N_17982,N_13601,N_11918);
xor U17983 (N_17983,N_10531,N_10455);
nor U17984 (N_17984,N_14687,N_10655);
nand U17985 (N_17985,N_12418,N_13417);
and U17986 (N_17986,N_12655,N_14698);
nand U17987 (N_17987,N_14511,N_14058);
nor U17988 (N_17988,N_13932,N_11604);
xnor U17989 (N_17989,N_14296,N_13755);
xor U17990 (N_17990,N_14177,N_14514);
nand U17991 (N_17991,N_11766,N_13375);
nor U17992 (N_17992,N_11084,N_11359);
and U17993 (N_17993,N_14002,N_14799);
nand U17994 (N_17994,N_12545,N_11433);
xnor U17995 (N_17995,N_11890,N_13126);
nand U17996 (N_17996,N_12839,N_10104);
nor U17997 (N_17997,N_10056,N_14391);
xnor U17998 (N_17998,N_14683,N_14225);
and U17999 (N_17999,N_10990,N_11791);
nand U18000 (N_18000,N_13412,N_12720);
xor U18001 (N_18001,N_11507,N_13577);
and U18002 (N_18002,N_10975,N_12372);
and U18003 (N_18003,N_12964,N_11527);
or U18004 (N_18004,N_10846,N_13782);
and U18005 (N_18005,N_14889,N_13711);
nor U18006 (N_18006,N_14373,N_10831);
xor U18007 (N_18007,N_11233,N_10525);
or U18008 (N_18008,N_10265,N_11191);
xnor U18009 (N_18009,N_11595,N_12306);
nand U18010 (N_18010,N_12035,N_12581);
nor U18011 (N_18011,N_14265,N_14380);
nand U18012 (N_18012,N_12139,N_11377);
or U18013 (N_18013,N_10134,N_11143);
and U18014 (N_18014,N_13993,N_10493);
xnor U18015 (N_18015,N_11068,N_14207);
nor U18016 (N_18016,N_13633,N_10481);
xnor U18017 (N_18017,N_12551,N_13000);
and U18018 (N_18018,N_11020,N_13553);
or U18019 (N_18019,N_10993,N_13678);
or U18020 (N_18020,N_11208,N_14968);
nand U18021 (N_18021,N_13754,N_10877);
and U18022 (N_18022,N_12993,N_10716);
or U18023 (N_18023,N_12480,N_14514);
nand U18024 (N_18024,N_11765,N_13375);
xor U18025 (N_18025,N_14559,N_14033);
and U18026 (N_18026,N_10970,N_13380);
xor U18027 (N_18027,N_14460,N_11588);
and U18028 (N_18028,N_10013,N_10230);
and U18029 (N_18029,N_12931,N_12828);
nand U18030 (N_18030,N_12451,N_13145);
and U18031 (N_18031,N_14117,N_10643);
and U18032 (N_18032,N_14756,N_12327);
xor U18033 (N_18033,N_12709,N_11658);
and U18034 (N_18034,N_11062,N_13297);
nand U18035 (N_18035,N_11407,N_14425);
xnor U18036 (N_18036,N_11367,N_14076);
xnor U18037 (N_18037,N_10996,N_10229);
and U18038 (N_18038,N_11229,N_11288);
and U18039 (N_18039,N_13317,N_14930);
and U18040 (N_18040,N_14573,N_10323);
xnor U18041 (N_18041,N_12816,N_11505);
nor U18042 (N_18042,N_10302,N_14226);
xnor U18043 (N_18043,N_10046,N_13006);
nand U18044 (N_18044,N_13537,N_13743);
xor U18045 (N_18045,N_10066,N_11520);
nor U18046 (N_18046,N_10227,N_11409);
xor U18047 (N_18047,N_13316,N_14676);
nor U18048 (N_18048,N_11393,N_12302);
or U18049 (N_18049,N_13897,N_12320);
xor U18050 (N_18050,N_11068,N_13053);
nor U18051 (N_18051,N_12135,N_10558);
and U18052 (N_18052,N_11217,N_10073);
nand U18053 (N_18053,N_11002,N_11217);
and U18054 (N_18054,N_13394,N_10794);
or U18055 (N_18055,N_11712,N_13762);
or U18056 (N_18056,N_10039,N_12243);
nor U18057 (N_18057,N_14772,N_10548);
nand U18058 (N_18058,N_12960,N_13551);
nand U18059 (N_18059,N_12055,N_11173);
and U18060 (N_18060,N_11367,N_11712);
or U18061 (N_18061,N_12881,N_12583);
and U18062 (N_18062,N_11515,N_14112);
and U18063 (N_18063,N_14646,N_13717);
and U18064 (N_18064,N_14968,N_13439);
nand U18065 (N_18065,N_13355,N_14251);
nand U18066 (N_18066,N_14201,N_10577);
nor U18067 (N_18067,N_12227,N_11023);
xor U18068 (N_18068,N_11044,N_12807);
and U18069 (N_18069,N_10365,N_14123);
nand U18070 (N_18070,N_14761,N_11991);
xor U18071 (N_18071,N_11384,N_14090);
nor U18072 (N_18072,N_10222,N_13680);
xor U18073 (N_18073,N_11617,N_11085);
nor U18074 (N_18074,N_10131,N_12274);
or U18075 (N_18075,N_10354,N_10086);
xor U18076 (N_18076,N_13182,N_13484);
xnor U18077 (N_18077,N_11467,N_10524);
xor U18078 (N_18078,N_12461,N_11532);
or U18079 (N_18079,N_14444,N_10577);
nand U18080 (N_18080,N_14250,N_12684);
nand U18081 (N_18081,N_11058,N_12555);
and U18082 (N_18082,N_14412,N_13399);
xor U18083 (N_18083,N_14579,N_14210);
and U18084 (N_18084,N_10146,N_14167);
and U18085 (N_18085,N_10843,N_11561);
and U18086 (N_18086,N_11245,N_11044);
xnor U18087 (N_18087,N_12228,N_13629);
nand U18088 (N_18088,N_10219,N_11693);
or U18089 (N_18089,N_11423,N_10252);
nor U18090 (N_18090,N_10070,N_10901);
xor U18091 (N_18091,N_12867,N_11322);
or U18092 (N_18092,N_12087,N_10269);
nor U18093 (N_18093,N_14426,N_13126);
and U18094 (N_18094,N_11001,N_10111);
nor U18095 (N_18095,N_10643,N_12709);
and U18096 (N_18096,N_12375,N_13652);
xnor U18097 (N_18097,N_12094,N_14259);
or U18098 (N_18098,N_14765,N_10588);
nand U18099 (N_18099,N_11904,N_11119);
or U18100 (N_18100,N_12658,N_14290);
nor U18101 (N_18101,N_10830,N_10722);
or U18102 (N_18102,N_11443,N_11852);
nand U18103 (N_18103,N_11813,N_11069);
or U18104 (N_18104,N_13816,N_14447);
or U18105 (N_18105,N_10596,N_11583);
and U18106 (N_18106,N_10401,N_11057);
xnor U18107 (N_18107,N_13115,N_13569);
or U18108 (N_18108,N_14319,N_11439);
nor U18109 (N_18109,N_11229,N_14677);
nand U18110 (N_18110,N_11187,N_13806);
and U18111 (N_18111,N_14237,N_11374);
and U18112 (N_18112,N_14715,N_12514);
and U18113 (N_18113,N_12940,N_14599);
nand U18114 (N_18114,N_11707,N_11377);
or U18115 (N_18115,N_12031,N_12672);
nand U18116 (N_18116,N_11468,N_10220);
and U18117 (N_18117,N_14961,N_11624);
and U18118 (N_18118,N_11290,N_12260);
xor U18119 (N_18119,N_10883,N_13156);
and U18120 (N_18120,N_11439,N_12232);
xnor U18121 (N_18121,N_14855,N_13183);
nand U18122 (N_18122,N_11970,N_10826);
and U18123 (N_18123,N_13382,N_10020);
xor U18124 (N_18124,N_11127,N_14247);
or U18125 (N_18125,N_10796,N_14675);
xor U18126 (N_18126,N_13308,N_10527);
and U18127 (N_18127,N_13598,N_13514);
and U18128 (N_18128,N_12157,N_12769);
and U18129 (N_18129,N_10709,N_12614);
and U18130 (N_18130,N_12546,N_10055);
and U18131 (N_18131,N_13494,N_10129);
nand U18132 (N_18132,N_12158,N_14951);
nand U18133 (N_18133,N_10543,N_14488);
and U18134 (N_18134,N_12714,N_10016);
xnor U18135 (N_18135,N_10549,N_12700);
or U18136 (N_18136,N_12270,N_14307);
xor U18137 (N_18137,N_10532,N_13087);
or U18138 (N_18138,N_13088,N_10848);
or U18139 (N_18139,N_10397,N_12626);
and U18140 (N_18140,N_11923,N_10688);
or U18141 (N_18141,N_13014,N_13480);
or U18142 (N_18142,N_11256,N_12921);
xor U18143 (N_18143,N_11944,N_11865);
nor U18144 (N_18144,N_12259,N_11191);
nand U18145 (N_18145,N_13124,N_11273);
xor U18146 (N_18146,N_11813,N_12751);
xnor U18147 (N_18147,N_14496,N_13286);
nor U18148 (N_18148,N_10902,N_10672);
nor U18149 (N_18149,N_12588,N_12884);
nor U18150 (N_18150,N_10880,N_11356);
nand U18151 (N_18151,N_10123,N_10086);
nand U18152 (N_18152,N_13080,N_12567);
nand U18153 (N_18153,N_10163,N_10459);
nand U18154 (N_18154,N_14950,N_13060);
nor U18155 (N_18155,N_10175,N_12467);
xnor U18156 (N_18156,N_13183,N_12606);
nor U18157 (N_18157,N_10885,N_12951);
xor U18158 (N_18158,N_12236,N_10882);
nand U18159 (N_18159,N_14760,N_14117);
and U18160 (N_18160,N_14197,N_13082);
xnor U18161 (N_18161,N_13595,N_11267);
or U18162 (N_18162,N_12406,N_11711);
nor U18163 (N_18163,N_11615,N_11339);
and U18164 (N_18164,N_13984,N_14245);
xor U18165 (N_18165,N_14938,N_13739);
and U18166 (N_18166,N_10493,N_12528);
nand U18167 (N_18167,N_10660,N_14334);
nor U18168 (N_18168,N_12184,N_12862);
nor U18169 (N_18169,N_14098,N_11106);
and U18170 (N_18170,N_13043,N_11562);
nor U18171 (N_18171,N_11857,N_10097);
nor U18172 (N_18172,N_12286,N_14189);
xor U18173 (N_18173,N_12609,N_14368);
xnor U18174 (N_18174,N_14415,N_13242);
or U18175 (N_18175,N_13901,N_13092);
nand U18176 (N_18176,N_11779,N_10466);
nor U18177 (N_18177,N_10866,N_11746);
nand U18178 (N_18178,N_11929,N_14752);
nor U18179 (N_18179,N_11447,N_11092);
or U18180 (N_18180,N_10689,N_13442);
xnor U18181 (N_18181,N_13160,N_14499);
xor U18182 (N_18182,N_12104,N_14523);
xor U18183 (N_18183,N_12672,N_13951);
xnor U18184 (N_18184,N_10821,N_14692);
nor U18185 (N_18185,N_14670,N_11910);
or U18186 (N_18186,N_12438,N_12412);
nor U18187 (N_18187,N_11085,N_14087);
or U18188 (N_18188,N_11694,N_11096);
nand U18189 (N_18189,N_12212,N_14679);
nor U18190 (N_18190,N_13962,N_14709);
and U18191 (N_18191,N_13328,N_14231);
or U18192 (N_18192,N_13487,N_13781);
xnor U18193 (N_18193,N_13811,N_10658);
and U18194 (N_18194,N_10613,N_12648);
nand U18195 (N_18195,N_11200,N_12148);
xnor U18196 (N_18196,N_13019,N_11011);
or U18197 (N_18197,N_12918,N_10899);
nor U18198 (N_18198,N_12921,N_11136);
nor U18199 (N_18199,N_11141,N_11897);
xnor U18200 (N_18200,N_13452,N_12236);
xor U18201 (N_18201,N_11628,N_11150);
nor U18202 (N_18202,N_14708,N_13441);
and U18203 (N_18203,N_14822,N_10973);
xnor U18204 (N_18204,N_10599,N_12516);
and U18205 (N_18205,N_10961,N_10828);
xnor U18206 (N_18206,N_11009,N_11906);
nor U18207 (N_18207,N_11055,N_13469);
nor U18208 (N_18208,N_10599,N_12186);
nand U18209 (N_18209,N_12132,N_11225);
nor U18210 (N_18210,N_10326,N_12538);
nand U18211 (N_18211,N_12237,N_13799);
xor U18212 (N_18212,N_11107,N_14766);
nand U18213 (N_18213,N_11068,N_10178);
nor U18214 (N_18214,N_14734,N_10520);
nand U18215 (N_18215,N_11802,N_11407);
or U18216 (N_18216,N_12618,N_12785);
nor U18217 (N_18217,N_10133,N_13369);
nand U18218 (N_18218,N_10838,N_13062);
nand U18219 (N_18219,N_10161,N_13236);
or U18220 (N_18220,N_11661,N_13978);
nor U18221 (N_18221,N_14660,N_12107);
nand U18222 (N_18222,N_12924,N_11055);
xnor U18223 (N_18223,N_13133,N_10860);
nor U18224 (N_18224,N_14715,N_11030);
and U18225 (N_18225,N_10897,N_13920);
and U18226 (N_18226,N_10446,N_12027);
or U18227 (N_18227,N_11353,N_12607);
and U18228 (N_18228,N_14976,N_12353);
xor U18229 (N_18229,N_10114,N_13995);
nand U18230 (N_18230,N_10170,N_12543);
or U18231 (N_18231,N_13601,N_10186);
nand U18232 (N_18232,N_14790,N_10569);
nor U18233 (N_18233,N_14553,N_12897);
nor U18234 (N_18234,N_12740,N_12023);
or U18235 (N_18235,N_14214,N_14399);
or U18236 (N_18236,N_13422,N_10940);
nor U18237 (N_18237,N_11365,N_14446);
nand U18238 (N_18238,N_10796,N_14928);
xor U18239 (N_18239,N_10883,N_12342);
xor U18240 (N_18240,N_10207,N_12282);
nand U18241 (N_18241,N_10147,N_13614);
xor U18242 (N_18242,N_13536,N_10208);
or U18243 (N_18243,N_14137,N_13409);
and U18244 (N_18244,N_14990,N_11991);
xnor U18245 (N_18245,N_12989,N_10134);
xor U18246 (N_18246,N_11527,N_14060);
nor U18247 (N_18247,N_13166,N_13044);
and U18248 (N_18248,N_11026,N_12208);
nand U18249 (N_18249,N_12056,N_13527);
nand U18250 (N_18250,N_11683,N_13048);
and U18251 (N_18251,N_11932,N_12983);
or U18252 (N_18252,N_10819,N_11277);
nand U18253 (N_18253,N_13680,N_10730);
and U18254 (N_18254,N_14001,N_14482);
nor U18255 (N_18255,N_13445,N_10431);
nand U18256 (N_18256,N_14920,N_10653);
and U18257 (N_18257,N_13393,N_13061);
xnor U18258 (N_18258,N_13091,N_10740);
nand U18259 (N_18259,N_10614,N_14347);
or U18260 (N_18260,N_10655,N_12124);
nor U18261 (N_18261,N_10017,N_13600);
xor U18262 (N_18262,N_10646,N_14409);
nor U18263 (N_18263,N_14596,N_13504);
or U18264 (N_18264,N_13805,N_14370);
nand U18265 (N_18265,N_14754,N_12511);
nor U18266 (N_18266,N_13488,N_10067);
and U18267 (N_18267,N_14298,N_14459);
or U18268 (N_18268,N_12303,N_11687);
nand U18269 (N_18269,N_14802,N_12446);
and U18270 (N_18270,N_14353,N_12204);
nand U18271 (N_18271,N_14185,N_11267);
and U18272 (N_18272,N_10506,N_12762);
xor U18273 (N_18273,N_10030,N_10878);
xor U18274 (N_18274,N_11082,N_14157);
nor U18275 (N_18275,N_12631,N_13762);
nand U18276 (N_18276,N_14328,N_12253);
xnor U18277 (N_18277,N_12117,N_12192);
and U18278 (N_18278,N_13849,N_11492);
or U18279 (N_18279,N_11329,N_11232);
nand U18280 (N_18280,N_12925,N_13586);
and U18281 (N_18281,N_12900,N_11479);
or U18282 (N_18282,N_12266,N_12497);
nor U18283 (N_18283,N_13776,N_12191);
xor U18284 (N_18284,N_14242,N_12889);
xnor U18285 (N_18285,N_14674,N_14499);
nor U18286 (N_18286,N_11010,N_14764);
xor U18287 (N_18287,N_12907,N_13847);
or U18288 (N_18288,N_11098,N_10427);
xor U18289 (N_18289,N_11895,N_10731);
and U18290 (N_18290,N_14589,N_14196);
and U18291 (N_18291,N_12050,N_12463);
nor U18292 (N_18292,N_12993,N_12519);
and U18293 (N_18293,N_14443,N_12388);
or U18294 (N_18294,N_10676,N_13378);
xnor U18295 (N_18295,N_11013,N_11635);
and U18296 (N_18296,N_10248,N_10088);
xor U18297 (N_18297,N_13792,N_14379);
xnor U18298 (N_18298,N_12125,N_10786);
or U18299 (N_18299,N_13959,N_11690);
or U18300 (N_18300,N_11317,N_10540);
nor U18301 (N_18301,N_11542,N_10167);
or U18302 (N_18302,N_10272,N_13039);
or U18303 (N_18303,N_13108,N_12362);
xor U18304 (N_18304,N_12256,N_13404);
xor U18305 (N_18305,N_11292,N_14292);
and U18306 (N_18306,N_13924,N_13136);
nand U18307 (N_18307,N_12756,N_14312);
nand U18308 (N_18308,N_14431,N_12026);
or U18309 (N_18309,N_14552,N_13446);
nor U18310 (N_18310,N_11147,N_13907);
nor U18311 (N_18311,N_11063,N_10017);
or U18312 (N_18312,N_12851,N_13993);
nor U18313 (N_18313,N_11834,N_10391);
and U18314 (N_18314,N_11369,N_13194);
xnor U18315 (N_18315,N_12611,N_11597);
nor U18316 (N_18316,N_12417,N_14066);
and U18317 (N_18317,N_11820,N_14917);
xnor U18318 (N_18318,N_13920,N_13179);
or U18319 (N_18319,N_10108,N_13608);
nand U18320 (N_18320,N_14463,N_12950);
and U18321 (N_18321,N_13537,N_11590);
or U18322 (N_18322,N_12074,N_10186);
or U18323 (N_18323,N_13703,N_12169);
nand U18324 (N_18324,N_14776,N_10611);
and U18325 (N_18325,N_12718,N_12091);
nor U18326 (N_18326,N_13432,N_11270);
or U18327 (N_18327,N_14293,N_10913);
nor U18328 (N_18328,N_11506,N_14215);
nor U18329 (N_18329,N_13996,N_10045);
xor U18330 (N_18330,N_14978,N_10601);
or U18331 (N_18331,N_11999,N_14832);
or U18332 (N_18332,N_10677,N_10235);
nor U18333 (N_18333,N_13269,N_14875);
and U18334 (N_18334,N_12475,N_12375);
nand U18335 (N_18335,N_13287,N_12775);
xnor U18336 (N_18336,N_14584,N_10728);
nor U18337 (N_18337,N_11814,N_10234);
nand U18338 (N_18338,N_12080,N_12722);
nand U18339 (N_18339,N_12292,N_10455);
nor U18340 (N_18340,N_14761,N_13382);
and U18341 (N_18341,N_14886,N_12723);
nand U18342 (N_18342,N_14368,N_11388);
nor U18343 (N_18343,N_13420,N_13214);
xnor U18344 (N_18344,N_12820,N_10029);
or U18345 (N_18345,N_11051,N_10576);
and U18346 (N_18346,N_12069,N_12600);
nor U18347 (N_18347,N_14153,N_13046);
or U18348 (N_18348,N_13149,N_11517);
nand U18349 (N_18349,N_10420,N_14546);
and U18350 (N_18350,N_10779,N_11138);
nand U18351 (N_18351,N_13847,N_13125);
xor U18352 (N_18352,N_11368,N_13598);
nand U18353 (N_18353,N_11115,N_11487);
nand U18354 (N_18354,N_12899,N_11207);
nor U18355 (N_18355,N_11103,N_10535);
xnor U18356 (N_18356,N_12450,N_14570);
and U18357 (N_18357,N_14523,N_14339);
nor U18358 (N_18358,N_12813,N_11902);
nor U18359 (N_18359,N_12370,N_10037);
and U18360 (N_18360,N_11542,N_11923);
or U18361 (N_18361,N_13344,N_11616);
nor U18362 (N_18362,N_12704,N_12487);
xnor U18363 (N_18363,N_12252,N_10147);
nand U18364 (N_18364,N_10378,N_10820);
nand U18365 (N_18365,N_11370,N_12836);
xnor U18366 (N_18366,N_14607,N_14684);
nor U18367 (N_18367,N_13758,N_11374);
nor U18368 (N_18368,N_11274,N_12189);
or U18369 (N_18369,N_10759,N_12978);
nor U18370 (N_18370,N_14150,N_11277);
xor U18371 (N_18371,N_12197,N_13277);
nand U18372 (N_18372,N_13681,N_10182);
and U18373 (N_18373,N_11057,N_13276);
or U18374 (N_18374,N_12768,N_13194);
nor U18375 (N_18375,N_12713,N_14039);
nand U18376 (N_18376,N_13183,N_14624);
or U18377 (N_18377,N_14667,N_14590);
nor U18378 (N_18378,N_14541,N_13536);
or U18379 (N_18379,N_11270,N_11423);
xor U18380 (N_18380,N_14275,N_14495);
or U18381 (N_18381,N_11000,N_12193);
nor U18382 (N_18382,N_12921,N_10010);
and U18383 (N_18383,N_13800,N_11111);
or U18384 (N_18384,N_13241,N_11872);
nand U18385 (N_18385,N_10311,N_14705);
nand U18386 (N_18386,N_14520,N_14271);
xor U18387 (N_18387,N_10201,N_12267);
nand U18388 (N_18388,N_10243,N_14387);
xor U18389 (N_18389,N_13206,N_11138);
nand U18390 (N_18390,N_13975,N_10863);
nand U18391 (N_18391,N_12445,N_10778);
and U18392 (N_18392,N_13170,N_14982);
xnor U18393 (N_18393,N_10474,N_12456);
nor U18394 (N_18394,N_12812,N_14806);
xor U18395 (N_18395,N_11592,N_11570);
nand U18396 (N_18396,N_14957,N_13259);
or U18397 (N_18397,N_11475,N_10203);
nand U18398 (N_18398,N_14100,N_10389);
nor U18399 (N_18399,N_14392,N_10956);
and U18400 (N_18400,N_12229,N_14976);
nor U18401 (N_18401,N_12282,N_12654);
or U18402 (N_18402,N_12638,N_14929);
nor U18403 (N_18403,N_11811,N_13195);
or U18404 (N_18404,N_14244,N_14327);
and U18405 (N_18405,N_11256,N_13594);
nand U18406 (N_18406,N_11666,N_12759);
nor U18407 (N_18407,N_11247,N_14125);
xor U18408 (N_18408,N_11013,N_13571);
xor U18409 (N_18409,N_14632,N_14653);
and U18410 (N_18410,N_13321,N_11958);
and U18411 (N_18411,N_10413,N_10639);
and U18412 (N_18412,N_12080,N_11487);
xnor U18413 (N_18413,N_10933,N_13854);
nor U18414 (N_18414,N_13754,N_13368);
nand U18415 (N_18415,N_12072,N_14150);
nor U18416 (N_18416,N_11138,N_11368);
or U18417 (N_18417,N_14938,N_11835);
xnor U18418 (N_18418,N_14776,N_12507);
nand U18419 (N_18419,N_11776,N_10766);
or U18420 (N_18420,N_14725,N_12139);
or U18421 (N_18421,N_12050,N_14441);
nand U18422 (N_18422,N_10930,N_13077);
or U18423 (N_18423,N_11189,N_13461);
nand U18424 (N_18424,N_10413,N_14750);
nand U18425 (N_18425,N_10916,N_10339);
xnor U18426 (N_18426,N_10676,N_12554);
xnor U18427 (N_18427,N_11665,N_11407);
nand U18428 (N_18428,N_13292,N_12387);
and U18429 (N_18429,N_10374,N_12181);
xnor U18430 (N_18430,N_11131,N_11351);
or U18431 (N_18431,N_12813,N_10306);
and U18432 (N_18432,N_11438,N_13336);
xor U18433 (N_18433,N_12708,N_11765);
nand U18434 (N_18434,N_14828,N_11607);
and U18435 (N_18435,N_11233,N_10690);
or U18436 (N_18436,N_11690,N_12213);
nand U18437 (N_18437,N_11064,N_10617);
or U18438 (N_18438,N_10287,N_11473);
nor U18439 (N_18439,N_11978,N_11416);
and U18440 (N_18440,N_12865,N_11648);
xnor U18441 (N_18441,N_11271,N_10166);
and U18442 (N_18442,N_12669,N_14823);
nor U18443 (N_18443,N_12393,N_11102);
nand U18444 (N_18444,N_14851,N_11039);
xor U18445 (N_18445,N_13256,N_13130);
nand U18446 (N_18446,N_10670,N_10965);
or U18447 (N_18447,N_10644,N_12702);
or U18448 (N_18448,N_12974,N_14300);
xor U18449 (N_18449,N_11626,N_12714);
or U18450 (N_18450,N_11944,N_13295);
nor U18451 (N_18451,N_12046,N_14279);
or U18452 (N_18452,N_10727,N_10597);
xor U18453 (N_18453,N_11058,N_12209);
and U18454 (N_18454,N_13508,N_10550);
or U18455 (N_18455,N_12546,N_10743);
xor U18456 (N_18456,N_14692,N_14032);
nor U18457 (N_18457,N_14871,N_12842);
or U18458 (N_18458,N_14666,N_12559);
nand U18459 (N_18459,N_12172,N_10952);
xor U18460 (N_18460,N_12756,N_11692);
nand U18461 (N_18461,N_14436,N_10627);
and U18462 (N_18462,N_12586,N_12695);
and U18463 (N_18463,N_12592,N_14746);
or U18464 (N_18464,N_10641,N_14130);
and U18465 (N_18465,N_14608,N_14019);
or U18466 (N_18466,N_10349,N_10678);
or U18467 (N_18467,N_10544,N_13065);
and U18468 (N_18468,N_11106,N_12964);
xnor U18469 (N_18469,N_12502,N_13275);
nand U18470 (N_18470,N_11815,N_11124);
and U18471 (N_18471,N_10283,N_10539);
or U18472 (N_18472,N_11086,N_14895);
nor U18473 (N_18473,N_14548,N_12958);
nor U18474 (N_18474,N_12816,N_14155);
nor U18475 (N_18475,N_10810,N_12058);
xor U18476 (N_18476,N_10101,N_12268);
nor U18477 (N_18477,N_13667,N_12217);
nand U18478 (N_18478,N_11256,N_12843);
and U18479 (N_18479,N_14609,N_13759);
xnor U18480 (N_18480,N_13271,N_11704);
xor U18481 (N_18481,N_12824,N_10099);
and U18482 (N_18482,N_12215,N_13415);
nor U18483 (N_18483,N_12823,N_11625);
nand U18484 (N_18484,N_10713,N_11475);
or U18485 (N_18485,N_12856,N_10046);
xor U18486 (N_18486,N_10198,N_12927);
or U18487 (N_18487,N_11801,N_12936);
and U18488 (N_18488,N_11596,N_14162);
xnor U18489 (N_18489,N_13292,N_10135);
and U18490 (N_18490,N_11953,N_11018);
and U18491 (N_18491,N_11587,N_12026);
and U18492 (N_18492,N_12071,N_14641);
and U18493 (N_18493,N_11212,N_14930);
xor U18494 (N_18494,N_11155,N_12456);
xor U18495 (N_18495,N_13272,N_10265);
and U18496 (N_18496,N_11435,N_14540);
and U18497 (N_18497,N_14992,N_13109);
nand U18498 (N_18498,N_10319,N_10799);
and U18499 (N_18499,N_13323,N_12899);
nand U18500 (N_18500,N_11969,N_13992);
or U18501 (N_18501,N_13669,N_12093);
or U18502 (N_18502,N_11475,N_11570);
or U18503 (N_18503,N_11682,N_10684);
xnor U18504 (N_18504,N_12450,N_14295);
and U18505 (N_18505,N_11430,N_14442);
nand U18506 (N_18506,N_11162,N_11595);
or U18507 (N_18507,N_14294,N_14042);
and U18508 (N_18508,N_13610,N_14881);
xor U18509 (N_18509,N_11335,N_13420);
nand U18510 (N_18510,N_14571,N_11173);
nor U18511 (N_18511,N_13130,N_14762);
and U18512 (N_18512,N_11245,N_12312);
nor U18513 (N_18513,N_11976,N_14595);
or U18514 (N_18514,N_12143,N_11946);
and U18515 (N_18515,N_13332,N_10197);
nand U18516 (N_18516,N_13427,N_12741);
and U18517 (N_18517,N_10861,N_14350);
and U18518 (N_18518,N_12666,N_11072);
xnor U18519 (N_18519,N_14892,N_13869);
nor U18520 (N_18520,N_10015,N_14984);
nor U18521 (N_18521,N_14274,N_12437);
nor U18522 (N_18522,N_12064,N_12695);
and U18523 (N_18523,N_13027,N_11681);
and U18524 (N_18524,N_11768,N_10323);
nand U18525 (N_18525,N_12839,N_14465);
and U18526 (N_18526,N_10921,N_11337);
nor U18527 (N_18527,N_13548,N_11568);
nand U18528 (N_18528,N_10418,N_13247);
and U18529 (N_18529,N_14111,N_13831);
xnor U18530 (N_18530,N_13001,N_11461);
and U18531 (N_18531,N_14238,N_14652);
xor U18532 (N_18532,N_13722,N_12104);
nor U18533 (N_18533,N_13894,N_10540);
xnor U18534 (N_18534,N_11434,N_11480);
and U18535 (N_18535,N_14282,N_11689);
xor U18536 (N_18536,N_11783,N_11023);
xor U18537 (N_18537,N_10438,N_12666);
or U18538 (N_18538,N_11912,N_11678);
xnor U18539 (N_18539,N_13523,N_10180);
nor U18540 (N_18540,N_10763,N_13150);
nor U18541 (N_18541,N_12428,N_13929);
xor U18542 (N_18542,N_14387,N_14304);
xor U18543 (N_18543,N_11339,N_14870);
nand U18544 (N_18544,N_10333,N_10016);
or U18545 (N_18545,N_10393,N_13337);
xnor U18546 (N_18546,N_12652,N_12779);
nand U18547 (N_18547,N_12470,N_12028);
xor U18548 (N_18548,N_11891,N_14350);
or U18549 (N_18549,N_13780,N_10999);
and U18550 (N_18550,N_12933,N_14873);
and U18551 (N_18551,N_11334,N_14170);
and U18552 (N_18552,N_13464,N_10150);
nor U18553 (N_18553,N_14781,N_13589);
nor U18554 (N_18554,N_14099,N_11078);
and U18555 (N_18555,N_12186,N_13951);
xor U18556 (N_18556,N_11813,N_12863);
nor U18557 (N_18557,N_13518,N_10069);
and U18558 (N_18558,N_10009,N_12817);
nor U18559 (N_18559,N_12342,N_14467);
nor U18560 (N_18560,N_14127,N_12089);
or U18561 (N_18561,N_14285,N_12519);
and U18562 (N_18562,N_11687,N_13735);
and U18563 (N_18563,N_12597,N_10132);
nand U18564 (N_18564,N_11547,N_14660);
xnor U18565 (N_18565,N_11893,N_10881);
nor U18566 (N_18566,N_13289,N_11220);
nand U18567 (N_18567,N_10495,N_14262);
nand U18568 (N_18568,N_14303,N_10986);
or U18569 (N_18569,N_10754,N_12576);
xnor U18570 (N_18570,N_13781,N_13768);
and U18571 (N_18571,N_14177,N_11442);
xnor U18572 (N_18572,N_14993,N_11584);
nand U18573 (N_18573,N_14542,N_14010);
and U18574 (N_18574,N_14777,N_14389);
or U18575 (N_18575,N_10835,N_13778);
or U18576 (N_18576,N_12647,N_11384);
or U18577 (N_18577,N_12859,N_10464);
xnor U18578 (N_18578,N_13388,N_13730);
nor U18579 (N_18579,N_14819,N_11788);
nand U18580 (N_18580,N_11483,N_10681);
and U18581 (N_18581,N_12785,N_11649);
nand U18582 (N_18582,N_12835,N_12484);
or U18583 (N_18583,N_14511,N_13298);
nand U18584 (N_18584,N_12942,N_10623);
or U18585 (N_18585,N_12566,N_13786);
nand U18586 (N_18586,N_11574,N_10078);
xnor U18587 (N_18587,N_11719,N_13754);
xor U18588 (N_18588,N_14200,N_10241);
nor U18589 (N_18589,N_13446,N_11624);
nor U18590 (N_18590,N_13250,N_14806);
xnor U18591 (N_18591,N_12075,N_14600);
or U18592 (N_18592,N_14808,N_10550);
or U18593 (N_18593,N_11323,N_14560);
xor U18594 (N_18594,N_14355,N_11845);
nor U18595 (N_18595,N_14652,N_14721);
nor U18596 (N_18596,N_13185,N_13737);
or U18597 (N_18597,N_14786,N_10746);
or U18598 (N_18598,N_10893,N_13153);
xnor U18599 (N_18599,N_14838,N_10154);
nor U18600 (N_18600,N_13353,N_11647);
nor U18601 (N_18601,N_12241,N_14123);
or U18602 (N_18602,N_11336,N_11560);
nor U18603 (N_18603,N_13069,N_14664);
nor U18604 (N_18604,N_11306,N_10189);
or U18605 (N_18605,N_10316,N_10443);
nor U18606 (N_18606,N_10115,N_13451);
or U18607 (N_18607,N_12512,N_11274);
xnor U18608 (N_18608,N_11143,N_14090);
and U18609 (N_18609,N_11962,N_10475);
or U18610 (N_18610,N_10011,N_11794);
and U18611 (N_18611,N_11588,N_13045);
nand U18612 (N_18612,N_13080,N_14076);
nand U18613 (N_18613,N_12470,N_11678);
nand U18614 (N_18614,N_10676,N_11791);
and U18615 (N_18615,N_14777,N_10141);
nand U18616 (N_18616,N_12558,N_12857);
nor U18617 (N_18617,N_14894,N_10256);
and U18618 (N_18618,N_12134,N_12273);
xor U18619 (N_18619,N_10079,N_14168);
xnor U18620 (N_18620,N_13912,N_11828);
or U18621 (N_18621,N_13829,N_12922);
xor U18622 (N_18622,N_10851,N_14279);
and U18623 (N_18623,N_11861,N_10024);
and U18624 (N_18624,N_14054,N_14056);
nand U18625 (N_18625,N_11393,N_13457);
nor U18626 (N_18626,N_11732,N_14342);
nand U18627 (N_18627,N_10275,N_14718);
and U18628 (N_18628,N_11828,N_13866);
nand U18629 (N_18629,N_12617,N_13714);
or U18630 (N_18630,N_11826,N_11788);
nand U18631 (N_18631,N_12257,N_12503);
and U18632 (N_18632,N_10202,N_13068);
and U18633 (N_18633,N_10982,N_11865);
nor U18634 (N_18634,N_13796,N_11620);
xor U18635 (N_18635,N_10093,N_13140);
xor U18636 (N_18636,N_13840,N_11256);
xor U18637 (N_18637,N_11752,N_13156);
or U18638 (N_18638,N_13960,N_10054);
nor U18639 (N_18639,N_10956,N_10636);
xnor U18640 (N_18640,N_14108,N_12340);
xnor U18641 (N_18641,N_12444,N_11703);
nand U18642 (N_18642,N_11960,N_12578);
nand U18643 (N_18643,N_10179,N_10385);
nor U18644 (N_18644,N_10294,N_12755);
or U18645 (N_18645,N_13958,N_14443);
nand U18646 (N_18646,N_14834,N_13183);
and U18647 (N_18647,N_11962,N_14710);
and U18648 (N_18648,N_10851,N_13045);
and U18649 (N_18649,N_10547,N_10484);
xnor U18650 (N_18650,N_13692,N_10056);
xnor U18651 (N_18651,N_13389,N_12916);
xnor U18652 (N_18652,N_11724,N_10450);
nand U18653 (N_18653,N_13439,N_13803);
xnor U18654 (N_18654,N_13814,N_14089);
or U18655 (N_18655,N_10641,N_10836);
or U18656 (N_18656,N_12358,N_10630);
xnor U18657 (N_18657,N_10504,N_12079);
xor U18658 (N_18658,N_11746,N_12072);
nor U18659 (N_18659,N_10073,N_11656);
nor U18660 (N_18660,N_12803,N_13629);
or U18661 (N_18661,N_14925,N_10645);
or U18662 (N_18662,N_10151,N_10096);
nand U18663 (N_18663,N_14416,N_10495);
nand U18664 (N_18664,N_14477,N_14771);
xor U18665 (N_18665,N_12317,N_10400);
nor U18666 (N_18666,N_13218,N_10283);
or U18667 (N_18667,N_10892,N_11620);
or U18668 (N_18668,N_14487,N_10239);
and U18669 (N_18669,N_14684,N_12253);
nor U18670 (N_18670,N_13750,N_12004);
or U18671 (N_18671,N_14782,N_10633);
nor U18672 (N_18672,N_11402,N_12031);
nand U18673 (N_18673,N_13436,N_10208);
and U18674 (N_18674,N_13246,N_13245);
and U18675 (N_18675,N_13050,N_12842);
nor U18676 (N_18676,N_12176,N_13927);
nor U18677 (N_18677,N_10001,N_13989);
or U18678 (N_18678,N_11241,N_14890);
nand U18679 (N_18679,N_13797,N_10168);
nor U18680 (N_18680,N_10025,N_14919);
or U18681 (N_18681,N_13957,N_13346);
nand U18682 (N_18682,N_12290,N_13962);
and U18683 (N_18683,N_14497,N_13945);
or U18684 (N_18684,N_10881,N_11617);
or U18685 (N_18685,N_11451,N_11120);
xor U18686 (N_18686,N_10814,N_10424);
and U18687 (N_18687,N_13937,N_10974);
and U18688 (N_18688,N_10748,N_11239);
or U18689 (N_18689,N_14918,N_11041);
nor U18690 (N_18690,N_12933,N_12825);
nand U18691 (N_18691,N_13123,N_10670);
xnor U18692 (N_18692,N_12225,N_13473);
and U18693 (N_18693,N_10258,N_10595);
nand U18694 (N_18694,N_11682,N_14876);
nand U18695 (N_18695,N_11826,N_10809);
nand U18696 (N_18696,N_13244,N_14859);
and U18697 (N_18697,N_11776,N_12073);
xor U18698 (N_18698,N_10692,N_11478);
and U18699 (N_18699,N_12697,N_12400);
xnor U18700 (N_18700,N_12018,N_12980);
nor U18701 (N_18701,N_12394,N_10363);
nor U18702 (N_18702,N_12495,N_14429);
xor U18703 (N_18703,N_14862,N_10666);
xnor U18704 (N_18704,N_14549,N_11479);
or U18705 (N_18705,N_12917,N_13712);
xnor U18706 (N_18706,N_12672,N_14008);
and U18707 (N_18707,N_13306,N_10437);
or U18708 (N_18708,N_13696,N_14737);
nor U18709 (N_18709,N_12551,N_10138);
or U18710 (N_18710,N_14192,N_11015);
and U18711 (N_18711,N_12978,N_10050);
or U18712 (N_18712,N_10684,N_13543);
and U18713 (N_18713,N_14247,N_11331);
nand U18714 (N_18714,N_12583,N_10592);
nor U18715 (N_18715,N_13919,N_11370);
xnor U18716 (N_18716,N_14182,N_14363);
and U18717 (N_18717,N_11960,N_14800);
nand U18718 (N_18718,N_10124,N_13828);
nand U18719 (N_18719,N_14546,N_12448);
nor U18720 (N_18720,N_12906,N_14720);
and U18721 (N_18721,N_10180,N_11980);
xor U18722 (N_18722,N_13753,N_13672);
or U18723 (N_18723,N_13369,N_12327);
or U18724 (N_18724,N_11905,N_12491);
nand U18725 (N_18725,N_13117,N_14131);
and U18726 (N_18726,N_12901,N_12221);
nor U18727 (N_18727,N_10166,N_14618);
nand U18728 (N_18728,N_11987,N_11520);
nand U18729 (N_18729,N_12510,N_12500);
nand U18730 (N_18730,N_14271,N_11946);
or U18731 (N_18731,N_11024,N_14693);
and U18732 (N_18732,N_13761,N_10112);
and U18733 (N_18733,N_13617,N_10768);
or U18734 (N_18734,N_13945,N_11684);
xor U18735 (N_18735,N_14473,N_14972);
nand U18736 (N_18736,N_12833,N_13989);
xnor U18737 (N_18737,N_10016,N_12579);
and U18738 (N_18738,N_10782,N_11975);
nand U18739 (N_18739,N_13363,N_14207);
nor U18740 (N_18740,N_11201,N_12577);
or U18741 (N_18741,N_14298,N_14718);
nor U18742 (N_18742,N_12351,N_13109);
and U18743 (N_18743,N_10162,N_10923);
xnor U18744 (N_18744,N_13808,N_14799);
and U18745 (N_18745,N_14636,N_14299);
nand U18746 (N_18746,N_11978,N_11320);
and U18747 (N_18747,N_12084,N_13112);
nand U18748 (N_18748,N_10057,N_12581);
and U18749 (N_18749,N_11035,N_10380);
nor U18750 (N_18750,N_14246,N_13108);
or U18751 (N_18751,N_11438,N_13415);
nor U18752 (N_18752,N_12421,N_13511);
or U18753 (N_18753,N_12013,N_10884);
xnor U18754 (N_18754,N_10548,N_10165);
nor U18755 (N_18755,N_11265,N_11327);
or U18756 (N_18756,N_14518,N_10041);
and U18757 (N_18757,N_11642,N_13294);
nor U18758 (N_18758,N_10791,N_12261);
xnor U18759 (N_18759,N_10857,N_12060);
nor U18760 (N_18760,N_10634,N_13701);
nand U18761 (N_18761,N_12486,N_12984);
xor U18762 (N_18762,N_14923,N_14537);
or U18763 (N_18763,N_14436,N_12744);
or U18764 (N_18764,N_12624,N_13954);
xor U18765 (N_18765,N_11018,N_13270);
nor U18766 (N_18766,N_10148,N_10353);
and U18767 (N_18767,N_14241,N_13042);
or U18768 (N_18768,N_13510,N_13880);
and U18769 (N_18769,N_12677,N_13949);
nor U18770 (N_18770,N_12854,N_10554);
and U18771 (N_18771,N_13852,N_12924);
nor U18772 (N_18772,N_14340,N_13993);
or U18773 (N_18773,N_10026,N_14622);
nor U18774 (N_18774,N_12505,N_10856);
xnor U18775 (N_18775,N_11846,N_13858);
and U18776 (N_18776,N_10417,N_10696);
nor U18777 (N_18777,N_13001,N_14664);
xor U18778 (N_18778,N_10753,N_14240);
and U18779 (N_18779,N_13047,N_11896);
nand U18780 (N_18780,N_13391,N_12204);
nand U18781 (N_18781,N_14727,N_12915);
nor U18782 (N_18782,N_12578,N_10454);
xor U18783 (N_18783,N_11412,N_14537);
nand U18784 (N_18784,N_12646,N_12639);
and U18785 (N_18785,N_13446,N_13616);
or U18786 (N_18786,N_11890,N_14039);
nor U18787 (N_18787,N_14037,N_10150);
xnor U18788 (N_18788,N_12793,N_13785);
nor U18789 (N_18789,N_10884,N_14233);
nor U18790 (N_18790,N_13078,N_10389);
nand U18791 (N_18791,N_14062,N_14822);
xor U18792 (N_18792,N_13856,N_11391);
and U18793 (N_18793,N_13062,N_11772);
nor U18794 (N_18794,N_12883,N_12611);
nor U18795 (N_18795,N_13024,N_12383);
nand U18796 (N_18796,N_14055,N_12916);
or U18797 (N_18797,N_10480,N_11780);
nor U18798 (N_18798,N_12161,N_10393);
xnor U18799 (N_18799,N_13450,N_13957);
xnor U18800 (N_18800,N_13044,N_11492);
nand U18801 (N_18801,N_14552,N_13379);
nor U18802 (N_18802,N_11844,N_11316);
nand U18803 (N_18803,N_10261,N_13353);
xnor U18804 (N_18804,N_10284,N_14774);
nor U18805 (N_18805,N_13044,N_11535);
nor U18806 (N_18806,N_11988,N_12122);
and U18807 (N_18807,N_12862,N_14779);
and U18808 (N_18808,N_14610,N_10867);
xnor U18809 (N_18809,N_11109,N_12195);
nor U18810 (N_18810,N_14480,N_10573);
xnor U18811 (N_18811,N_12191,N_12261);
nand U18812 (N_18812,N_13386,N_12171);
nand U18813 (N_18813,N_14390,N_14001);
nand U18814 (N_18814,N_13341,N_11171);
xnor U18815 (N_18815,N_13000,N_10517);
or U18816 (N_18816,N_10250,N_11947);
and U18817 (N_18817,N_11437,N_12771);
nand U18818 (N_18818,N_13955,N_13443);
and U18819 (N_18819,N_10529,N_14019);
nand U18820 (N_18820,N_14642,N_13131);
or U18821 (N_18821,N_11848,N_10378);
or U18822 (N_18822,N_10505,N_11175);
or U18823 (N_18823,N_11985,N_11957);
and U18824 (N_18824,N_14785,N_11770);
and U18825 (N_18825,N_11943,N_12990);
xor U18826 (N_18826,N_14319,N_10953);
nand U18827 (N_18827,N_11062,N_12192);
nor U18828 (N_18828,N_11178,N_14034);
xnor U18829 (N_18829,N_13966,N_14677);
or U18830 (N_18830,N_13024,N_11570);
and U18831 (N_18831,N_14220,N_14661);
nor U18832 (N_18832,N_14135,N_10760);
xnor U18833 (N_18833,N_12863,N_10324);
or U18834 (N_18834,N_14952,N_14092);
and U18835 (N_18835,N_12258,N_11698);
nand U18836 (N_18836,N_14035,N_14570);
or U18837 (N_18837,N_14592,N_10426);
nor U18838 (N_18838,N_12592,N_13198);
nor U18839 (N_18839,N_11720,N_14785);
nor U18840 (N_18840,N_13945,N_13313);
xor U18841 (N_18841,N_11272,N_14621);
nor U18842 (N_18842,N_11338,N_14990);
nand U18843 (N_18843,N_11305,N_13316);
xor U18844 (N_18844,N_11884,N_12318);
and U18845 (N_18845,N_14099,N_12565);
nand U18846 (N_18846,N_12639,N_12014);
nor U18847 (N_18847,N_10422,N_12281);
nor U18848 (N_18848,N_13585,N_11916);
xor U18849 (N_18849,N_14102,N_12474);
and U18850 (N_18850,N_11797,N_12632);
and U18851 (N_18851,N_14410,N_11489);
xor U18852 (N_18852,N_12854,N_11164);
or U18853 (N_18853,N_14500,N_14857);
nand U18854 (N_18854,N_10823,N_11995);
and U18855 (N_18855,N_11837,N_12473);
nand U18856 (N_18856,N_12491,N_13497);
and U18857 (N_18857,N_11882,N_11950);
xnor U18858 (N_18858,N_10249,N_11634);
nor U18859 (N_18859,N_11097,N_10612);
nand U18860 (N_18860,N_11276,N_14705);
xor U18861 (N_18861,N_11947,N_13894);
and U18862 (N_18862,N_13862,N_13193);
nand U18863 (N_18863,N_12715,N_14915);
nand U18864 (N_18864,N_13805,N_12418);
nand U18865 (N_18865,N_11125,N_11758);
nand U18866 (N_18866,N_12193,N_12878);
or U18867 (N_18867,N_10770,N_11825);
nand U18868 (N_18868,N_12285,N_11726);
nor U18869 (N_18869,N_10566,N_13580);
or U18870 (N_18870,N_10403,N_13630);
and U18871 (N_18871,N_10992,N_12398);
nand U18872 (N_18872,N_12146,N_14594);
nor U18873 (N_18873,N_14894,N_13306);
or U18874 (N_18874,N_12177,N_12735);
xnor U18875 (N_18875,N_13999,N_10991);
nor U18876 (N_18876,N_10770,N_10091);
xor U18877 (N_18877,N_14359,N_14650);
and U18878 (N_18878,N_13684,N_10684);
xor U18879 (N_18879,N_14009,N_13551);
nand U18880 (N_18880,N_12668,N_13318);
xor U18881 (N_18881,N_11686,N_12786);
nand U18882 (N_18882,N_10032,N_11936);
and U18883 (N_18883,N_10415,N_13305);
or U18884 (N_18884,N_14398,N_13443);
or U18885 (N_18885,N_13691,N_14454);
nand U18886 (N_18886,N_11283,N_10165);
xnor U18887 (N_18887,N_10513,N_14463);
nand U18888 (N_18888,N_10889,N_13952);
nor U18889 (N_18889,N_13495,N_10495);
nand U18890 (N_18890,N_14058,N_14931);
nor U18891 (N_18891,N_10306,N_11502);
and U18892 (N_18892,N_14137,N_10082);
nand U18893 (N_18893,N_11753,N_11165);
nand U18894 (N_18894,N_12076,N_13963);
or U18895 (N_18895,N_12498,N_13297);
or U18896 (N_18896,N_12167,N_10588);
and U18897 (N_18897,N_12226,N_14473);
nand U18898 (N_18898,N_14975,N_12393);
and U18899 (N_18899,N_11629,N_14178);
and U18900 (N_18900,N_10297,N_13652);
or U18901 (N_18901,N_12695,N_14782);
nand U18902 (N_18902,N_14740,N_13740);
and U18903 (N_18903,N_13498,N_14239);
and U18904 (N_18904,N_10736,N_12617);
and U18905 (N_18905,N_10239,N_12826);
and U18906 (N_18906,N_10957,N_13887);
xor U18907 (N_18907,N_10052,N_10663);
and U18908 (N_18908,N_13828,N_12114);
xor U18909 (N_18909,N_12295,N_14232);
nand U18910 (N_18910,N_10723,N_13023);
nor U18911 (N_18911,N_14181,N_11961);
and U18912 (N_18912,N_12272,N_14424);
nand U18913 (N_18913,N_13438,N_14510);
xnor U18914 (N_18914,N_11514,N_11302);
and U18915 (N_18915,N_11958,N_14792);
nor U18916 (N_18916,N_12566,N_11805);
and U18917 (N_18917,N_10037,N_11779);
nor U18918 (N_18918,N_14609,N_14000);
and U18919 (N_18919,N_13707,N_10123);
nor U18920 (N_18920,N_12088,N_13681);
or U18921 (N_18921,N_13549,N_14073);
xor U18922 (N_18922,N_13472,N_12276);
nand U18923 (N_18923,N_11347,N_10947);
and U18924 (N_18924,N_10158,N_12198);
xnor U18925 (N_18925,N_11040,N_14420);
nor U18926 (N_18926,N_13754,N_11052);
nor U18927 (N_18927,N_10203,N_10969);
or U18928 (N_18928,N_14172,N_10452);
and U18929 (N_18929,N_13009,N_13820);
xnor U18930 (N_18930,N_10376,N_14643);
or U18931 (N_18931,N_14517,N_12291);
nand U18932 (N_18932,N_11880,N_11680);
xnor U18933 (N_18933,N_12839,N_12588);
nand U18934 (N_18934,N_11893,N_10588);
nand U18935 (N_18935,N_10527,N_11376);
and U18936 (N_18936,N_13613,N_12486);
xnor U18937 (N_18937,N_10970,N_13710);
and U18938 (N_18938,N_12641,N_12357);
xor U18939 (N_18939,N_13412,N_11303);
and U18940 (N_18940,N_13273,N_12549);
and U18941 (N_18941,N_14555,N_14748);
xor U18942 (N_18942,N_10102,N_14294);
and U18943 (N_18943,N_12941,N_12949);
nor U18944 (N_18944,N_14202,N_13244);
and U18945 (N_18945,N_10741,N_11900);
nor U18946 (N_18946,N_11416,N_13600);
nand U18947 (N_18947,N_13126,N_11223);
nor U18948 (N_18948,N_12630,N_10900);
and U18949 (N_18949,N_13476,N_12497);
and U18950 (N_18950,N_10530,N_10860);
or U18951 (N_18951,N_11854,N_12897);
nor U18952 (N_18952,N_13582,N_11789);
or U18953 (N_18953,N_13765,N_12895);
nand U18954 (N_18954,N_12146,N_11247);
nand U18955 (N_18955,N_12079,N_13232);
xor U18956 (N_18956,N_13472,N_14765);
nor U18957 (N_18957,N_14746,N_12751);
or U18958 (N_18958,N_11326,N_14174);
xor U18959 (N_18959,N_10904,N_14929);
xnor U18960 (N_18960,N_14525,N_13037);
nand U18961 (N_18961,N_10278,N_11704);
or U18962 (N_18962,N_13262,N_13304);
or U18963 (N_18963,N_13513,N_12064);
or U18964 (N_18964,N_12279,N_10875);
or U18965 (N_18965,N_13921,N_10924);
or U18966 (N_18966,N_10433,N_13037);
and U18967 (N_18967,N_10513,N_13300);
or U18968 (N_18968,N_10773,N_14548);
or U18969 (N_18969,N_13884,N_13285);
and U18970 (N_18970,N_11542,N_14914);
and U18971 (N_18971,N_13423,N_12783);
xnor U18972 (N_18972,N_11782,N_13802);
and U18973 (N_18973,N_14452,N_14363);
nor U18974 (N_18974,N_11662,N_10686);
xnor U18975 (N_18975,N_13883,N_13495);
xor U18976 (N_18976,N_10949,N_13737);
xor U18977 (N_18977,N_11191,N_10650);
nor U18978 (N_18978,N_14829,N_11932);
xnor U18979 (N_18979,N_13197,N_10178);
nor U18980 (N_18980,N_11568,N_10735);
nor U18981 (N_18981,N_10288,N_12714);
or U18982 (N_18982,N_13015,N_12463);
or U18983 (N_18983,N_11599,N_14982);
nand U18984 (N_18984,N_12771,N_11337);
xnor U18985 (N_18985,N_13049,N_10197);
or U18986 (N_18986,N_11475,N_10632);
or U18987 (N_18987,N_13669,N_13573);
nor U18988 (N_18988,N_12046,N_13222);
and U18989 (N_18989,N_13634,N_11875);
xnor U18990 (N_18990,N_11968,N_14099);
and U18991 (N_18991,N_11931,N_13277);
nand U18992 (N_18992,N_14659,N_11253);
xnor U18993 (N_18993,N_11855,N_10599);
or U18994 (N_18994,N_11463,N_14259);
nand U18995 (N_18995,N_11241,N_13470);
and U18996 (N_18996,N_13090,N_12012);
nand U18997 (N_18997,N_13309,N_10042);
nor U18998 (N_18998,N_10689,N_10128);
or U18999 (N_18999,N_11070,N_10747);
xnor U19000 (N_19000,N_14408,N_12220);
xor U19001 (N_19001,N_13439,N_11192);
nand U19002 (N_19002,N_11844,N_10303);
and U19003 (N_19003,N_11412,N_13339);
or U19004 (N_19004,N_12538,N_14108);
or U19005 (N_19005,N_13458,N_14142);
or U19006 (N_19006,N_14504,N_13672);
nor U19007 (N_19007,N_10097,N_12278);
nand U19008 (N_19008,N_14310,N_10348);
nand U19009 (N_19009,N_12381,N_14713);
or U19010 (N_19010,N_13719,N_12838);
nand U19011 (N_19011,N_12661,N_11831);
or U19012 (N_19012,N_12349,N_13868);
nor U19013 (N_19013,N_12602,N_14195);
and U19014 (N_19014,N_11259,N_12949);
nand U19015 (N_19015,N_10653,N_14090);
or U19016 (N_19016,N_11435,N_11290);
and U19017 (N_19017,N_11828,N_11886);
xnor U19018 (N_19018,N_10327,N_13750);
xnor U19019 (N_19019,N_14846,N_10638);
or U19020 (N_19020,N_11744,N_14003);
nor U19021 (N_19021,N_12602,N_13750);
xor U19022 (N_19022,N_14562,N_13713);
and U19023 (N_19023,N_14107,N_12926);
nor U19024 (N_19024,N_11755,N_12772);
nand U19025 (N_19025,N_10151,N_13454);
and U19026 (N_19026,N_13746,N_14905);
nand U19027 (N_19027,N_12738,N_12756);
xor U19028 (N_19028,N_10083,N_10339);
xnor U19029 (N_19029,N_12211,N_11827);
nand U19030 (N_19030,N_14399,N_13963);
nor U19031 (N_19031,N_13063,N_12832);
nor U19032 (N_19032,N_11856,N_10497);
nor U19033 (N_19033,N_10855,N_14946);
nand U19034 (N_19034,N_12347,N_12403);
and U19035 (N_19035,N_13880,N_12566);
and U19036 (N_19036,N_10168,N_12682);
nand U19037 (N_19037,N_10145,N_11304);
and U19038 (N_19038,N_13820,N_13674);
and U19039 (N_19039,N_14862,N_10588);
nand U19040 (N_19040,N_10712,N_11534);
nand U19041 (N_19041,N_10349,N_10464);
nor U19042 (N_19042,N_12227,N_10220);
and U19043 (N_19043,N_12709,N_10541);
nor U19044 (N_19044,N_10304,N_11806);
xnor U19045 (N_19045,N_11953,N_14000);
nor U19046 (N_19046,N_10284,N_12337);
nor U19047 (N_19047,N_13835,N_12080);
and U19048 (N_19048,N_13197,N_10487);
or U19049 (N_19049,N_14549,N_10236);
xor U19050 (N_19050,N_11419,N_13538);
or U19051 (N_19051,N_14625,N_10667);
xor U19052 (N_19052,N_13445,N_14637);
and U19053 (N_19053,N_12765,N_14633);
nor U19054 (N_19054,N_12832,N_14488);
or U19055 (N_19055,N_10336,N_14371);
nor U19056 (N_19056,N_13635,N_12571);
nand U19057 (N_19057,N_12740,N_10918);
and U19058 (N_19058,N_11273,N_11784);
or U19059 (N_19059,N_11566,N_10913);
and U19060 (N_19060,N_10367,N_12958);
nor U19061 (N_19061,N_10266,N_10689);
xor U19062 (N_19062,N_14542,N_13632);
nor U19063 (N_19063,N_14775,N_14470);
xor U19064 (N_19064,N_14384,N_14487);
or U19065 (N_19065,N_13319,N_14511);
nand U19066 (N_19066,N_14483,N_12273);
or U19067 (N_19067,N_14067,N_14409);
nor U19068 (N_19068,N_14374,N_12946);
nor U19069 (N_19069,N_10734,N_10692);
or U19070 (N_19070,N_10415,N_10353);
nand U19071 (N_19071,N_10305,N_11480);
or U19072 (N_19072,N_13133,N_14373);
nand U19073 (N_19073,N_13783,N_13284);
or U19074 (N_19074,N_13194,N_10142);
nor U19075 (N_19075,N_11567,N_13329);
xnor U19076 (N_19076,N_12720,N_14931);
nor U19077 (N_19077,N_13777,N_12029);
nor U19078 (N_19078,N_10858,N_11026);
or U19079 (N_19079,N_11878,N_11000);
and U19080 (N_19080,N_14450,N_11853);
nand U19081 (N_19081,N_13139,N_14774);
nand U19082 (N_19082,N_12312,N_12416);
nor U19083 (N_19083,N_14052,N_13894);
nor U19084 (N_19084,N_12733,N_12867);
nor U19085 (N_19085,N_12813,N_11225);
or U19086 (N_19086,N_10518,N_14346);
nand U19087 (N_19087,N_12662,N_10865);
xnor U19088 (N_19088,N_11364,N_11549);
nor U19089 (N_19089,N_12906,N_13603);
nor U19090 (N_19090,N_10919,N_12537);
nor U19091 (N_19091,N_10387,N_11273);
nand U19092 (N_19092,N_12912,N_12842);
xor U19093 (N_19093,N_10872,N_10046);
nor U19094 (N_19094,N_10131,N_13222);
and U19095 (N_19095,N_12009,N_10993);
nor U19096 (N_19096,N_11184,N_12283);
and U19097 (N_19097,N_10047,N_11031);
nor U19098 (N_19098,N_12325,N_11150);
xnor U19099 (N_19099,N_13703,N_14543);
nor U19100 (N_19100,N_13338,N_11648);
and U19101 (N_19101,N_14573,N_11315);
xnor U19102 (N_19102,N_12960,N_13053);
xor U19103 (N_19103,N_11293,N_13264);
and U19104 (N_19104,N_10677,N_11846);
nor U19105 (N_19105,N_12379,N_10758);
nor U19106 (N_19106,N_13919,N_12830);
and U19107 (N_19107,N_10543,N_11347);
and U19108 (N_19108,N_13499,N_10142);
nand U19109 (N_19109,N_14909,N_11899);
nor U19110 (N_19110,N_13309,N_14289);
or U19111 (N_19111,N_10641,N_11195);
nand U19112 (N_19112,N_12014,N_12706);
xnor U19113 (N_19113,N_13999,N_12727);
nand U19114 (N_19114,N_13925,N_11589);
nand U19115 (N_19115,N_12513,N_11969);
nor U19116 (N_19116,N_13410,N_12913);
xor U19117 (N_19117,N_11904,N_14667);
and U19118 (N_19118,N_12255,N_10193);
or U19119 (N_19119,N_11264,N_12591);
or U19120 (N_19120,N_11746,N_13989);
and U19121 (N_19121,N_11433,N_10736);
and U19122 (N_19122,N_12116,N_14143);
and U19123 (N_19123,N_11763,N_11364);
and U19124 (N_19124,N_10575,N_10406);
and U19125 (N_19125,N_11683,N_12202);
nor U19126 (N_19126,N_10593,N_13669);
or U19127 (N_19127,N_10967,N_12839);
nand U19128 (N_19128,N_12073,N_14752);
nand U19129 (N_19129,N_10654,N_10824);
and U19130 (N_19130,N_11554,N_14810);
or U19131 (N_19131,N_14898,N_10392);
or U19132 (N_19132,N_10023,N_14268);
and U19133 (N_19133,N_10387,N_14435);
or U19134 (N_19134,N_11955,N_13552);
or U19135 (N_19135,N_13091,N_11574);
nand U19136 (N_19136,N_10550,N_14013);
or U19137 (N_19137,N_13546,N_11510);
or U19138 (N_19138,N_13440,N_13229);
xnor U19139 (N_19139,N_13427,N_11157);
and U19140 (N_19140,N_11010,N_11936);
and U19141 (N_19141,N_11595,N_14744);
nor U19142 (N_19142,N_13115,N_11560);
nand U19143 (N_19143,N_11962,N_10306);
xnor U19144 (N_19144,N_13494,N_12295);
nand U19145 (N_19145,N_10376,N_10991);
and U19146 (N_19146,N_14819,N_12311);
and U19147 (N_19147,N_14624,N_13112);
or U19148 (N_19148,N_11974,N_10304);
or U19149 (N_19149,N_13499,N_14379);
nand U19150 (N_19150,N_14689,N_10952);
and U19151 (N_19151,N_13098,N_13028);
nand U19152 (N_19152,N_13580,N_12689);
nand U19153 (N_19153,N_12435,N_11290);
and U19154 (N_19154,N_12432,N_10032);
nor U19155 (N_19155,N_14138,N_14501);
nor U19156 (N_19156,N_12229,N_14839);
nand U19157 (N_19157,N_12851,N_12557);
or U19158 (N_19158,N_12277,N_14872);
or U19159 (N_19159,N_11425,N_10971);
or U19160 (N_19160,N_13933,N_11098);
nand U19161 (N_19161,N_11323,N_12946);
nand U19162 (N_19162,N_10149,N_10085);
nor U19163 (N_19163,N_10138,N_14118);
xnor U19164 (N_19164,N_12364,N_12026);
and U19165 (N_19165,N_10501,N_13229);
and U19166 (N_19166,N_13800,N_12844);
nand U19167 (N_19167,N_12563,N_11517);
nand U19168 (N_19168,N_11053,N_10558);
xor U19169 (N_19169,N_14164,N_13976);
xnor U19170 (N_19170,N_14899,N_11686);
and U19171 (N_19171,N_12935,N_14066);
and U19172 (N_19172,N_14984,N_14264);
or U19173 (N_19173,N_14002,N_13567);
nor U19174 (N_19174,N_12060,N_13714);
xnor U19175 (N_19175,N_12582,N_11717);
or U19176 (N_19176,N_10334,N_12391);
nor U19177 (N_19177,N_10894,N_13845);
nand U19178 (N_19178,N_11923,N_10711);
xor U19179 (N_19179,N_11873,N_14369);
and U19180 (N_19180,N_13915,N_14832);
or U19181 (N_19181,N_13825,N_13299);
or U19182 (N_19182,N_13202,N_10567);
nor U19183 (N_19183,N_14232,N_11206);
and U19184 (N_19184,N_14519,N_11077);
nor U19185 (N_19185,N_13920,N_11472);
or U19186 (N_19186,N_10476,N_14629);
or U19187 (N_19187,N_10442,N_10900);
nor U19188 (N_19188,N_13649,N_13984);
and U19189 (N_19189,N_11034,N_14483);
nor U19190 (N_19190,N_10260,N_11220);
or U19191 (N_19191,N_14484,N_13036);
and U19192 (N_19192,N_13431,N_10064);
and U19193 (N_19193,N_11815,N_11689);
and U19194 (N_19194,N_12775,N_12590);
nand U19195 (N_19195,N_12895,N_13946);
xnor U19196 (N_19196,N_10389,N_14639);
xor U19197 (N_19197,N_13510,N_14502);
nor U19198 (N_19198,N_10387,N_11537);
nor U19199 (N_19199,N_10930,N_11484);
xnor U19200 (N_19200,N_13713,N_10117);
nor U19201 (N_19201,N_13784,N_14673);
xor U19202 (N_19202,N_10675,N_14310);
or U19203 (N_19203,N_13777,N_13181);
nor U19204 (N_19204,N_13225,N_12193);
nor U19205 (N_19205,N_11546,N_11872);
and U19206 (N_19206,N_11614,N_10425);
xnor U19207 (N_19207,N_10399,N_14227);
xor U19208 (N_19208,N_13244,N_10401);
nor U19209 (N_19209,N_13382,N_10357);
nand U19210 (N_19210,N_11176,N_11688);
xor U19211 (N_19211,N_10417,N_12105);
or U19212 (N_19212,N_12275,N_12174);
nand U19213 (N_19213,N_14585,N_12395);
or U19214 (N_19214,N_13960,N_11265);
nand U19215 (N_19215,N_14534,N_10890);
nand U19216 (N_19216,N_12057,N_12126);
nor U19217 (N_19217,N_12758,N_11809);
nand U19218 (N_19218,N_13224,N_14465);
xnor U19219 (N_19219,N_13995,N_14588);
or U19220 (N_19220,N_12766,N_11656);
xor U19221 (N_19221,N_11502,N_13478);
nand U19222 (N_19222,N_13719,N_13495);
nor U19223 (N_19223,N_10745,N_14624);
nand U19224 (N_19224,N_10679,N_10267);
xor U19225 (N_19225,N_11540,N_10751);
nand U19226 (N_19226,N_14139,N_12384);
nand U19227 (N_19227,N_12859,N_10975);
nand U19228 (N_19228,N_13726,N_11328);
or U19229 (N_19229,N_13293,N_11652);
nand U19230 (N_19230,N_10937,N_10457);
nand U19231 (N_19231,N_10962,N_12941);
nand U19232 (N_19232,N_12716,N_14462);
or U19233 (N_19233,N_11576,N_11568);
or U19234 (N_19234,N_14298,N_14163);
nand U19235 (N_19235,N_14712,N_14219);
and U19236 (N_19236,N_11251,N_12536);
nand U19237 (N_19237,N_10868,N_10049);
nand U19238 (N_19238,N_10663,N_12316);
nand U19239 (N_19239,N_14026,N_11295);
and U19240 (N_19240,N_14024,N_11830);
nor U19241 (N_19241,N_14306,N_11456);
nor U19242 (N_19242,N_10105,N_11652);
or U19243 (N_19243,N_14314,N_12287);
xor U19244 (N_19244,N_14951,N_14634);
or U19245 (N_19245,N_14771,N_10548);
or U19246 (N_19246,N_10545,N_12828);
xnor U19247 (N_19247,N_13812,N_13167);
and U19248 (N_19248,N_14902,N_14686);
and U19249 (N_19249,N_11081,N_10655);
or U19250 (N_19250,N_10489,N_12126);
nand U19251 (N_19251,N_10179,N_12226);
and U19252 (N_19252,N_10653,N_13752);
xnor U19253 (N_19253,N_12111,N_13308);
or U19254 (N_19254,N_12646,N_13109);
and U19255 (N_19255,N_14078,N_11393);
nor U19256 (N_19256,N_11908,N_10137);
nor U19257 (N_19257,N_13912,N_10325);
and U19258 (N_19258,N_14260,N_12075);
xor U19259 (N_19259,N_14196,N_14989);
xnor U19260 (N_19260,N_10046,N_12866);
nand U19261 (N_19261,N_12402,N_13919);
nand U19262 (N_19262,N_10656,N_12786);
nor U19263 (N_19263,N_12115,N_12881);
or U19264 (N_19264,N_12322,N_12332);
nand U19265 (N_19265,N_10840,N_14645);
or U19266 (N_19266,N_12175,N_12576);
nor U19267 (N_19267,N_12665,N_12965);
and U19268 (N_19268,N_10965,N_10078);
or U19269 (N_19269,N_14093,N_12221);
or U19270 (N_19270,N_11170,N_11104);
and U19271 (N_19271,N_11229,N_12244);
and U19272 (N_19272,N_14970,N_11693);
xor U19273 (N_19273,N_11019,N_12945);
or U19274 (N_19274,N_13920,N_12434);
or U19275 (N_19275,N_13715,N_13766);
and U19276 (N_19276,N_14924,N_11777);
nor U19277 (N_19277,N_13762,N_12915);
and U19278 (N_19278,N_13465,N_13696);
nand U19279 (N_19279,N_13465,N_14119);
xor U19280 (N_19280,N_11361,N_14883);
or U19281 (N_19281,N_14345,N_11676);
nand U19282 (N_19282,N_14176,N_11772);
and U19283 (N_19283,N_11326,N_14567);
nor U19284 (N_19284,N_12823,N_12724);
nand U19285 (N_19285,N_14406,N_10456);
or U19286 (N_19286,N_14137,N_12749);
xor U19287 (N_19287,N_10379,N_14745);
and U19288 (N_19288,N_10117,N_11018);
or U19289 (N_19289,N_14358,N_10235);
nor U19290 (N_19290,N_10625,N_10857);
nor U19291 (N_19291,N_10565,N_14696);
or U19292 (N_19292,N_11912,N_11148);
nand U19293 (N_19293,N_13535,N_10529);
nor U19294 (N_19294,N_14007,N_13040);
nand U19295 (N_19295,N_11352,N_13532);
xor U19296 (N_19296,N_12147,N_11833);
nor U19297 (N_19297,N_11215,N_12579);
and U19298 (N_19298,N_14581,N_11727);
or U19299 (N_19299,N_11855,N_10637);
or U19300 (N_19300,N_11510,N_10378);
or U19301 (N_19301,N_11635,N_12803);
and U19302 (N_19302,N_13701,N_12341);
xor U19303 (N_19303,N_12249,N_13394);
nand U19304 (N_19304,N_12520,N_10627);
xnor U19305 (N_19305,N_10378,N_13740);
nand U19306 (N_19306,N_10049,N_13155);
nand U19307 (N_19307,N_12064,N_13765);
and U19308 (N_19308,N_10134,N_12196);
and U19309 (N_19309,N_10118,N_10014);
or U19310 (N_19310,N_13507,N_10624);
nor U19311 (N_19311,N_13682,N_12251);
nand U19312 (N_19312,N_10922,N_14750);
xor U19313 (N_19313,N_14812,N_11964);
xor U19314 (N_19314,N_12202,N_13875);
xor U19315 (N_19315,N_10647,N_11974);
nor U19316 (N_19316,N_12157,N_10423);
nor U19317 (N_19317,N_11360,N_13389);
nand U19318 (N_19318,N_13516,N_13609);
xnor U19319 (N_19319,N_12738,N_11126);
nand U19320 (N_19320,N_10807,N_10703);
xnor U19321 (N_19321,N_12239,N_14773);
nand U19322 (N_19322,N_10168,N_10894);
xor U19323 (N_19323,N_11363,N_11292);
xor U19324 (N_19324,N_14624,N_11309);
or U19325 (N_19325,N_12134,N_14054);
and U19326 (N_19326,N_13833,N_11146);
or U19327 (N_19327,N_12877,N_13921);
nand U19328 (N_19328,N_14557,N_11278);
or U19329 (N_19329,N_12014,N_12576);
nand U19330 (N_19330,N_10506,N_13638);
nor U19331 (N_19331,N_13663,N_14181);
nor U19332 (N_19332,N_12117,N_10041);
nor U19333 (N_19333,N_14052,N_13760);
xnor U19334 (N_19334,N_14502,N_14208);
xor U19335 (N_19335,N_13507,N_13337);
nor U19336 (N_19336,N_10409,N_11202);
nor U19337 (N_19337,N_11109,N_13335);
nor U19338 (N_19338,N_14106,N_14267);
nand U19339 (N_19339,N_10576,N_10186);
nor U19340 (N_19340,N_10285,N_11539);
nor U19341 (N_19341,N_13686,N_13913);
nor U19342 (N_19342,N_14945,N_13844);
nand U19343 (N_19343,N_10109,N_13095);
nor U19344 (N_19344,N_10493,N_11353);
or U19345 (N_19345,N_11360,N_13325);
xnor U19346 (N_19346,N_12066,N_14538);
nor U19347 (N_19347,N_12133,N_12598);
or U19348 (N_19348,N_14251,N_12347);
nor U19349 (N_19349,N_11058,N_14956);
and U19350 (N_19350,N_14345,N_10031);
and U19351 (N_19351,N_14953,N_11958);
nand U19352 (N_19352,N_14155,N_11518);
xnor U19353 (N_19353,N_12547,N_11382);
nand U19354 (N_19354,N_10927,N_14708);
and U19355 (N_19355,N_14813,N_13125);
and U19356 (N_19356,N_14951,N_12666);
xor U19357 (N_19357,N_12078,N_10662);
and U19358 (N_19358,N_11791,N_13111);
xnor U19359 (N_19359,N_13360,N_14519);
nand U19360 (N_19360,N_13812,N_11958);
nand U19361 (N_19361,N_14074,N_10981);
nand U19362 (N_19362,N_13524,N_12863);
nor U19363 (N_19363,N_12538,N_11208);
or U19364 (N_19364,N_14231,N_12207);
nand U19365 (N_19365,N_14982,N_13808);
or U19366 (N_19366,N_10890,N_10332);
and U19367 (N_19367,N_14976,N_14895);
nand U19368 (N_19368,N_14404,N_12817);
nor U19369 (N_19369,N_14257,N_10256);
and U19370 (N_19370,N_11702,N_14438);
or U19371 (N_19371,N_10528,N_14602);
nand U19372 (N_19372,N_14367,N_14844);
or U19373 (N_19373,N_13069,N_14678);
nor U19374 (N_19374,N_13173,N_13774);
nor U19375 (N_19375,N_13239,N_12564);
nand U19376 (N_19376,N_14084,N_11934);
or U19377 (N_19377,N_10528,N_14457);
or U19378 (N_19378,N_10860,N_13776);
nor U19379 (N_19379,N_10923,N_10961);
nor U19380 (N_19380,N_12682,N_12763);
nand U19381 (N_19381,N_10470,N_12236);
or U19382 (N_19382,N_12210,N_10806);
nand U19383 (N_19383,N_12394,N_13805);
nand U19384 (N_19384,N_10379,N_10023);
nand U19385 (N_19385,N_12766,N_11901);
nand U19386 (N_19386,N_10786,N_13458);
and U19387 (N_19387,N_12432,N_13130);
or U19388 (N_19388,N_13494,N_12177);
or U19389 (N_19389,N_14837,N_12530);
and U19390 (N_19390,N_10689,N_10682);
nor U19391 (N_19391,N_12968,N_13619);
xor U19392 (N_19392,N_11254,N_10835);
nor U19393 (N_19393,N_11544,N_13597);
nand U19394 (N_19394,N_13373,N_10994);
nand U19395 (N_19395,N_10451,N_12853);
nor U19396 (N_19396,N_13786,N_11811);
or U19397 (N_19397,N_12533,N_13394);
nand U19398 (N_19398,N_12590,N_13086);
xnor U19399 (N_19399,N_10236,N_10196);
or U19400 (N_19400,N_12668,N_13488);
nand U19401 (N_19401,N_11728,N_13701);
xnor U19402 (N_19402,N_14552,N_13211);
xnor U19403 (N_19403,N_11055,N_13188);
nor U19404 (N_19404,N_13652,N_10594);
and U19405 (N_19405,N_11198,N_12556);
and U19406 (N_19406,N_13331,N_10825);
nor U19407 (N_19407,N_13531,N_11828);
and U19408 (N_19408,N_10671,N_12511);
xnor U19409 (N_19409,N_14710,N_10781);
or U19410 (N_19410,N_12299,N_14579);
or U19411 (N_19411,N_13086,N_14072);
and U19412 (N_19412,N_10451,N_11073);
and U19413 (N_19413,N_12546,N_11520);
nand U19414 (N_19414,N_14941,N_11616);
or U19415 (N_19415,N_11823,N_12843);
and U19416 (N_19416,N_14357,N_14163);
xnor U19417 (N_19417,N_10172,N_10277);
or U19418 (N_19418,N_14753,N_12576);
xor U19419 (N_19419,N_11982,N_13827);
xnor U19420 (N_19420,N_11853,N_14166);
and U19421 (N_19421,N_13878,N_11429);
and U19422 (N_19422,N_14990,N_13801);
xor U19423 (N_19423,N_13416,N_12847);
xor U19424 (N_19424,N_12159,N_14125);
nor U19425 (N_19425,N_12959,N_11949);
nor U19426 (N_19426,N_12950,N_11682);
and U19427 (N_19427,N_10344,N_10436);
xor U19428 (N_19428,N_14647,N_12378);
xor U19429 (N_19429,N_13828,N_13793);
xnor U19430 (N_19430,N_11750,N_10942);
nand U19431 (N_19431,N_12018,N_11439);
nor U19432 (N_19432,N_14886,N_10849);
nand U19433 (N_19433,N_13231,N_11177);
and U19434 (N_19434,N_13712,N_13762);
xor U19435 (N_19435,N_14039,N_11815);
or U19436 (N_19436,N_14172,N_11342);
nor U19437 (N_19437,N_13974,N_12185);
xor U19438 (N_19438,N_11385,N_10231);
xor U19439 (N_19439,N_10369,N_12779);
xnor U19440 (N_19440,N_14864,N_13823);
and U19441 (N_19441,N_14911,N_10536);
xnor U19442 (N_19442,N_13899,N_10354);
or U19443 (N_19443,N_13949,N_12974);
and U19444 (N_19444,N_10161,N_13028);
xnor U19445 (N_19445,N_14082,N_14087);
and U19446 (N_19446,N_12771,N_14671);
or U19447 (N_19447,N_13860,N_14853);
and U19448 (N_19448,N_14833,N_14867);
and U19449 (N_19449,N_12940,N_13269);
and U19450 (N_19450,N_14435,N_11329);
and U19451 (N_19451,N_13397,N_14040);
nor U19452 (N_19452,N_10645,N_10363);
nor U19453 (N_19453,N_11047,N_10846);
xor U19454 (N_19454,N_13745,N_14604);
nor U19455 (N_19455,N_14245,N_12488);
nand U19456 (N_19456,N_12477,N_13951);
nand U19457 (N_19457,N_10460,N_14030);
or U19458 (N_19458,N_11151,N_12705);
and U19459 (N_19459,N_10460,N_14864);
nand U19460 (N_19460,N_10205,N_14824);
and U19461 (N_19461,N_13684,N_14453);
or U19462 (N_19462,N_11983,N_13514);
and U19463 (N_19463,N_11519,N_12611);
nor U19464 (N_19464,N_14378,N_14954);
and U19465 (N_19465,N_13557,N_11714);
xor U19466 (N_19466,N_10593,N_10476);
or U19467 (N_19467,N_11433,N_14626);
nor U19468 (N_19468,N_10665,N_11696);
xnor U19469 (N_19469,N_14748,N_11697);
xor U19470 (N_19470,N_11718,N_13118);
or U19471 (N_19471,N_13820,N_13373);
xnor U19472 (N_19472,N_11081,N_12754);
xnor U19473 (N_19473,N_13112,N_14678);
and U19474 (N_19474,N_11156,N_11107);
or U19475 (N_19475,N_14346,N_11857);
or U19476 (N_19476,N_12879,N_12545);
or U19477 (N_19477,N_10843,N_11131);
and U19478 (N_19478,N_13316,N_12152);
nand U19479 (N_19479,N_13315,N_13089);
nand U19480 (N_19480,N_11690,N_12366);
or U19481 (N_19481,N_10793,N_11771);
xor U19482 (N_19482,N_10523,N_11065);
and U19483 (N_19483,N_12354,N_10584);
nor U19484 (N_19484,N_11097,N_13258);
or U19485 (N_19485,N_13145,N_13376);
or U19486 (N_19486,N_13713,N_12730);
and U19487 (N_19487,N_10608,N_12521);
and U19488 (N_19488,N_12887,N_11640);
and U19489 (N_19489,N_10255,N_13501);
nor U19490 (N_19490,N_14708,N_12336);
or U19491 (N_19491,N_13552,N_13511);
nand U19492 (N_19492,N_13213,N_12958);
or U19493 (N_19493,N_14611,N_12764);
xor U19494 (N_19494,N_10261,N_13513);
nor U19495 (N_19495,N_10686,N_10164);
nand U19496 (N_19496,N_11249,N_13762);
nand U19497 (N_19497,N_11632,N_12729);
and U19498 (N_19498,N_10257,N_10596);
nor U19499 (N_19499,N_11471,N_14793);
and U19500 (N_19500,N_14088,N_10759);
nand U19501 (N_19501,N_13553,N_12835);
or U19502 (N_19502,N_14181,N_14445);
nand U19503 (N_19503,N_14427,N_12838);
or U19504 (N_19504,N_12995,N_12228);
or U19505 (N_19505,N_12209,N_10938);
or U19506 (N_19506,N_12238,N_11128);
xnor U19507 (N_19507,N_11197,N_13130);
xor U19508 (N_19508,N_10491,N_12295);
xor U19509 (N_19509,N_11369,N_13695);
nor U19510 (N_19510,N_12148,N_13327);
xor U19511 (N_19511,N_11802,N_12201);
nor U19512 (N_19512,N_10034,N_10566);
nand U19513 (N_19513,N_14062,N_10241);
and U19514 (N_19514,N_14370,N_13557);
nor U19515 (N_19515,N_14879,N_14393);
and U19516 (N_19516,N_10118,N_11745);
nand U19517 (N_19517,N_11668,N_12710);
nand U19518 (N_19518,N_14995,N_12838);
or U19519 (N_19519,N_14251,N_11066);
or U19520 (N_19520,N_14791,N_10032);
or U19521 (N_19521,N_14887,N_13505);
xnor U19522 (N_19522,N_13559,N_13410);
or U19523 (N_19523,N_11592,N_12524);
nand U19524 (N_19524,N_10626,N_13053);
xor U19525 (N_19525,N_10111,N_13633);
nand U19526 (N_19526,N_14793,N_14789);
nand U19527 (N_19527,N_11828,N_14392);
nor U19528 (N_19528,N_13301,N_10400);
nand U19529 (N_19529,N_11280,N_12454);
xnor U19530 (N_19530,N_11213,N_11028);
or U19531 (N_19531,N_12594,N_13229);
nand U19532 (N_19532,N_13685,N_14976);
and U19533 (N_19533,N_12717,N_10910);
nand U19534 (N_19534,N_11502,N_10912);
nand U19535 (N_19535,N_11824,N_13637);
nand U19536 (N_19536,N_11379,N_12773);
xor U19537 (N_19537,N_12039,N_11850);
and U19538 (N_19538,N_13279,N_13725);
and U19539 (N_19539,N_13758,N_13541);
xor U19540 (N_19540,N_11348,N_12851);
or U19541 (N_19541,N_10404,N_11536);
or U19542 (N_19542,N_12963,N_10680);
nor U19543 (N_19543,N_10789,N_12354);
or U19544 (N_19544,N_13003,N_14738);
or U19545 (N_19545,N_14355,N_14077);
nor U19546 (N_19546,N_13782,N_12972);
nand U19547 (N_19547,N_12882,N_13937);
nand U19548 (N_19548,N_13343,N_10409);
or U19549 (N_19549,N_11117,N_14977);
nor U19550 (N_19550,N_12827,N_14687);
or U19551 (N_19551,N_12402,N_13478);
nor U19552 (N_19552,N_12876,N_13591);
nor U19553 (N_19553,N_14626,N_10469);
nor U19554 (N_19554,N_12660,N_12305);
or U19555 (N_19555,N_11916,N_12614);
nand U19556 (N_19556,N_12280,N_12000);
xor U19557 (N_19557,N_14683,N_11170);
or U19558 (N_19558,N_13110,N_12138);
and U19559 (N_19559,N_10388,N_14039);
and U19560 (N_19560,N_11079,N_13648);
nor U19561 (N_19561,N_14321,N_12928);
xor U19562 (N_19562,N_11913,N_10128);
xnor U19563 (N_19563,N_10456,N_11125);
xnor U19564 (N_19564,N_11000,N_14974);
or U19565 (N_19565,N_13486,N_13075);
xnor U19566 (N_19566,N_14823,N_13833);
nor U19567 (N_19567,N_10625,N_12286);
or U19568 (N_19568,N_12953,N_12064);
nor U19569 (N_19569,N_13108,N_10483);
nor U19570 (N_19570,N_13206,N_13745);
and U19571 (N_19571,N_13680,N_12573);
nand U19572 (N_19572,N_13682,N_12176);
and U19573 (N_19573,N_12664,N_10228);
or U19574 (N_19574,N_12079,N_10435);
nand U19575 (N_19575,N_11331,N_11062);
xor U19576 (N_19576,N_13467,N_13245);
and U19577 (N_19577,N_13915,N_10577);
and U19578 (N_19578,N_13568,N_14359);
or U19579 (N_19579,N_14980,N_14070);
or U19580 (N_19580,N_10142,N_11465);
or U19581 (N_19581,N_14567,N_11432);
or U19582 (N_19582,N_13228,N_12988);
or U19583 (N_19583,N_14673,N_12881);
nor U19584 (N_19584,N_11574,N_11217);
and U19585 (N_19585,N_11415,N_13730);
nor U19586 (N_19586,N_14325,N_11827);
and U19587 (N_19587,N_10901,N_12550);
nand U19588 (N_19588,N_10068,N_13514);
nor U19589 (N_19589,N_13363,N_12509);
or U19590 (N_19590,N_13002,N_14951);
nand U19591 (N_19591,N_12878,N_12224);
nand U19592 (N_19592,N_12033,N_14595);
or U19593 (N_19593,N_11917,N_11900);
or U19594 (N_19594,N_12917,N_10152);
or U19595 (N_19595,N_10221,N_11978);
or U19596 (N_19596,N_14233,N_12167);
and U19597 (N_19597,N_12788,N_10099);
and U19598 (N_19598,N_12855,N_12159);
nor U19599 (N_19599,N_10218,N_14839);
nor U19600 (N_19600,N_10740,N_12311);
and U19601 (N_19601,N_13854,N_13624);
nor U19602 (N_19602,N_10890,N_11476);
or U19603 (N_19603,N_14600,N_12955);
and U19604 (N_19604,N_14085,N_14567);
or U19605 (N_19605,N_14054,N_13744);
and U19606 (N_19606,N_10792,N_10797);
and U19607 (N_19607,N_11057,N_14640);
or U19608 (N_19608,N_14306,N_11519);
and U19609 (N_19609,N_11128,N_10157);
or U19610 (N_19610,N_12472,N_11901);
nor U19611 (N_19611,N_13666,N_14059);
and U19612 (N_19612,N_14738,N_10804);
and U19613 (N_19613,N_11348,N_14129);
nor U19614 (N_19614,N_10791,N_11144);
and U19615 (N_19615,N_12137,N_14108);
or U19616 (N_19616,N_11284,N_13636);
nor U19617 (N_19617,N_14380,N_10673);
nor U19618 (N_19618,N_11944,N_13243);
nand U19619 (N_19619,N_13379,N_12616);
nor U19620 (N_19620,N_12940,N_12214);
nand U19621 (N_19621,N_12200,N_11958);
and U19622 (N_19622,N_11146,N_10805);
nand U19623 (N_19623,N_14125,N_10508);
or U19624 (N_19624,N_12668,N_10969);
nand U19625 (N_19625,N_12222,N_11561);
and U19626 (N_19626,N_11628,N_12712);
xnor U19627 (N_19627,N_10198,N_14177);
nand U19628 (N_19628,N_12010,N_12891);
nand U19629 (N_19629,N_13525,N_11361);
nor U19630 (N_19630,N_14254,N_10335);
and U19631 (N_19631,N_11522,N_11190);
xor U19632 (N_19632,N_10728,N_14100);
and U19633 (N_19633,N_13225,N_10799);
and U19634 (N_19634,N_14348,N_14114);
and U19635 (N_19635,N_13517,N_12954);
and U19636 (N_19636,N_13000,N_11334);
xnor U19637 (N_19637,N_13383,N_12996);
nor U19638 (N_19638,N_10999,N_10975);
and U19639 (N_19639,N_14196,N_11063);
nand U19640 (N_19640,N_10331,N_11129);
nand U19641 (N_19641,N_13085,N_13244);
or U19642 (N_19642,N_10474,N_11141);
nor U19643 (N_19643,N_11623,N_12312);
or U19644 (N_19644,N_13107,N_12336);
or U19645 (N_19645,N_11949,N_12585);
nor U19646 (N_19646,N_13533,N_12463);
and U19647 (N_19647,N_13047,N_14355);
nor U19648 (N_19648,N_14721,N_12099);
and U19649 (N_19649,N_14031,N_11875);
and U19650 (N_19650,N_11194,N_10046);
or U19651 (N_19651,N_12975,N_12711);
nand U19652 (N_19652,N_12897,N_11736);
xor U19653 (N_19653,N_12716,N_12892);
or U19654 (N_19654,N_13711,N_14619);
nand U19655 (N_19655,N_13420,N_13609);
or U19656 (N_19656,N_12783,N_13525);
and U19657 (N_19657,N_10549,N_12912);
nand U19658 (N_19658,N_11446,N_14763);
or U19659 (N_19659,N_12804,N_14532);
and U19660 (N_19660,N_14241,N_12706);
nand U19661 (N_19661,N_10471,N_10694);
or U19662 (N_19662,N_11706,N_10246);
or U19663 (N_19663,N_12582,N_10809);
nor U19664 (N_19664,N_11404,N_14808);
or U19665 (N_19665,N_14709,N_10469);
nor U19666 (N_19666,N_10245,N_14073);
nand U19667 (N_19667,N_11561,N_11900);
or U19668 (N_19668,N_14075,N_10760);
or U19669 (N_19669,N_11351,N_13592);
xnor U19670 (N_19670,N_12745,N_13368);
nand U19671 (N_19671,N_11867,N_14505);
nand U19672 (N_19672,N_11698,N_14934);
or U19673 (N_19673,N_13766,N_13323);
xor U19674 (N_19674,N_14833,N_12538);
nand U19675 (N_19675,N_14704,N_10207);
xor U19676 (N_19676,N_11613,N_10981);
or U19677 (N_19677,N_11631,N_11614);
nand U19678 (N_19678,N_13881,N_10674);
nand U19679 (N_19679,N_10601,N_10568);
nor U19680 (N_19680,N_14637,N_13708);
nor U19681 (N_19681,N_14560,N_13948);
and U19682 (N_19682,N_10795,N_10285);
and U19683 (N_19683,N_12376,N_11936);
nand U19684 (N_19684,N_10502,N_12349);
or U19685 (N_19685,N_14036,N_12738);
xor U19686 (N_19686,N_10356,N_12794);
or U19687 (N_19687,N_12416,N_12857);
nand U19688 (N_19688,N_10421,N_11188);
xor U19689 (N_19689,N_12458,N_11320);
xor U19690 (N_19690,N_13227,N_11058);
or U19691 (N_19691,N_11528,N_13748);
nor U19692 (N_19692,N_11985,N_11464);
nor U19693 (N_19693,N_14302,N_14559);
nor U19694 (N_19694,N_12743,N_11307);
and U19695 (N_19695,N_11629,N_10172);
or U19696 (N_19696,N_12636,N_13047);
nand U19697 (N_19697,N_14873,N_11200);
and U19698 (N_19698,N_12225,N_10463);
xnor U19699 (N_19699,N_12189,N_10303);
nor U19700 (N_19700,N_10646,N_10982);
and U19701 (N_19701,N_12451,N_13659);
nor U19702 (N_19702,N_11021,N_13356);
nand U19703 (N_19703,N_11380,N_11959);
nand U19704 (N_19704,N_13389,N_14006);
or U19705 (N_19705,N_14381,N_14364);
xor U19706 (N_19706,N_10091,N_11109);
and U19707 (N_19707,N_10609,N_12567);
nor U19708 (N_19708,N_14893,N_10971);
nand U19709 (N_19709,N_13958,N_12784);
or U19710 (N_19710,N_11570,N_10004);
and U19711 (N_19711,N_10791,N_12390);
or U19712 (N_19712,N_11049,N_12351);
nand U19713 (N_19713,N_13788,N_11536);
nand U19714 (N_19714,N_14397,N_13547);
and U19715 (N_19715,N_11695,N_10392);
nor U19716 (N_19716,N_13565,N_10595);
or U19717 (N_19717,N_11232,N_11753);
xnor U19718 (N_19718,N_10101,N_13007);
xnor U19719 (N_19719,N_14008,N_11828);
nor U19720 (N_19720,N_11326,N_11979);
nor U19721 (N_19721,N_10457,N_13131);
and U19722 (N_19722,N_11062,N_10626);
xor U19723 (N_19723,N_12916,N_13109);
and U19724 (N_19724,N_14482,N_12757);
and U19725 (N_19725,N_13617,N_12330);
or U19726 (N_19726,N_12751,N_13661);
and U19727 (N_19727,N_12362,N_10918);
and U19728 (N_19728,N_11653,N_13813);
nor U19729 (N_19729,N_14752,N_11944);
nor U19730 (N_19730,N_12433,N_11906);
or U19731 (N_19731,N_13609,N_14165);
nor U19732 (N_19732,N_12604,N_10052);
and U19733 (N_19733,N_10043,N_12897);
and U19734 (N_19734,N_14941,N_11763);
xor U19735 (N_19735,N_14265,N_14398);
xnor U19736 (N_19736,N_14071,N_12824);
and U19737 (N_19737,N_14431,N_14917);
and U19738 (N_19738,N_13649,N_10139);
xor U19739 (N_19739,N_13322,N_12238);
or U19740 (N_19740,N_14113,N_12991);
or U19741 (N_19741,N_13661,N_12615);
nor U19742 (N_19742,N_11478,N_12001);
and U19743 (N_19743,N_12536,N_14015);
or U19744 (N_19744,N_10688,N_12773);
nor U19745 (N_19745,N_12185,N_10090);
nand U19746 (N_19746,N_11058,N_13425);
nor U19747 (N_19747,N_14388,N_13546);
nand U19748 (N_19748,N_10199,N_12626);
nor U19749 (N_19749,N_13967,N_12467);
or U19750 (N_19750,N_14173,N_13504);
xor U19751 (N_19751,N_11496,N_14242);
or U19752 (N_19752,N_14537,N_14865);
nor U19753 (N_19753,N_11779,N_13776);
nand U19754 (N_19754,N_12751,N_14492);
or U19755 (N_19755,N_10973,N_13008);
and U19756 (N_19756,N_12398,N_13490);
or U19757 (N_19757,N_14325,N_11587);
xor U19758 (N_19758,N_14601,N_14312);
nor U19759 (N_19759,N_14889,N_11453);
and U19760 (N_19760,N_10189,N_12860);
nand U19761 (N_19761,N_11429,N_11367);
and U19762 (N_19762,N_13765,N_10683);
nand U19763 (N_19763,N_12184,N_13071);
nor U19764 (N_19764,N_11716,N_13901);
and U19765 (N_19765,N_10842,N_14420);
or U19766 (N_19766,N_11333,N_11725);
nor U19767 (N_19767,N_14722,N_11070);
and U19768 (N_19768,N_14018,N_11305);
and U19769 (N_19769,N_10094,N_14024);
or U19770 (N_19770,N_12543,N_10829);
and U19771 (N_19771,N_11445,N_10250);
or U19772 (N_19772,N_14606,N_13694);
nand U19773 (N_19773,N_14060,N_10439);
xor U19774 (N_19774,N_10486,N_12417);
nor U19775 (N_19775,N_14554,N_14859);
nand U19776 (N_19776,N_11924,N_10832);
nor U19777 (N_19777,N_12797,N_12184);
nor U19778 (N_19778,N_11290,N_14698);
and U19779 (N_19779,N_13053,N_11562);
nor U19780 (N_19780,N_13273,N_12392);
xnor U19781 (N_19781,N_10537,N_13600);
or U19782 (N_19782,N_12834,N_11166);
xnor U19783 (N_19783,N_12545,N_11210);
xor U19784 (N_19784,N_14820,N_11798);
nand U19785 (N_19785,N_13601,N_10877);
nand U19786 (N_19786,N_10309,N_11642);
xnor U19787 (N_19787,N_14434,N_14799);
nor U19788 (N_19788,N_13406,N_14821);
or U19789 (N_19789,N_14780,N_10038);
nor U19790 (N_19790,N_10163,N_10358);
or U19791 (N_19791,N_14734,N_11302);
xor U19792 (N_19792,N_10486,N_12244);
and U19793 (N_19793,N_13080,N_11725);
nand U19794 (N_19794,N_12283,N_13155);
and U19795 (N_19795,N_13891,N_12534);
xor U19796 (N_19796,N_13334,N_13196);
nand U19797 (N_19797,N_12122,N_11546);
and U19798 (N_19798,N_10223,N_12228);
nor U19799 (N_19799,N_12160,N_13094);
or U19800 (N_19800,N_11764,N_12385);
and U19801 (N_19801,N_13985,N_13589);
nor U19802 (N_19802,N_13863,N_10904);
nand U19803 (N_19803,N_11065,N_12471);
and U19804 (N_19804,N_11308,N_12364);
or U19805 (N_19805,N_13861,N_14100);
xnor U19806 (N_19806,N_14186,N_11249);
and U19807 (N_19807,N_14301,N_14040);
and U19808 (N_19808,N_13539,N_13506);
nand U19809 (N_19809,N_11316,N_12023);
nand U19810 (N_19810,N_12397,N_14193);
xor U19811 (N_19811,N_14516,N_11535);
nor U19812 (N_19812,N_11769,N_12106);
and U19813 (N_19813,N_14127,N_14674);
and U19814 (N_19814,N_13926,N_10391);
and U19815 (N_19815,N_10612,N_11798);
xor U19816 (N_19816,N_11511,N_12723);
and U19817 (N_19817,N_13254,N_13736);
and U19818 (N_19818,N_13695,N_11340);
or U19819 (N_19819,N_14088,N_10403);
and U19820 (N_19820,N_14156,N_14429);
nand U19821 (N_19821,N_13649,N_14417);
nor U19822 (N_19822,N_10058,N_14078);
nand U19823 (N_19823,N_10279,N_12355);
nand U19824 (N_19824,N_10763,N_11241);
nor U19825 (N_19825,N_10643,N_11359);
xor U19826 (N_19826,N_10391,N_13865);
nor U19827 (N_19827,N_11095,N_12418);
and U19828 (N_19828,N_13004,N_13990);
xor U19829 (N_19829,N_10503,N_14150);
or U19830 (N_19830,N_10354,N_10470);
and U19831 (N_19831,N_11614,N_14950);
or U19832 (N_19832,N_11945,N_12371);
nand U19833 (N_19833,N_14577,N_12090);
and U19834 (N_19834,N_12634,N_13374);
nand U19835 (N_19835,N_11884,N_10180);
nor U19836 (N_19836,N_13978,N_13512);
nor U19837 (N_19837,N_12967,N_12299);
nand U19838 (N_19838,N_12085,N_12551);
nor U19839 (N_19839,N_12475,N_14632);
and U19840 (N_19840,N_14577,N_10807);
nand U19841 (N_19841,N_11771,N_12023);
nor U19842 (N_19842,N_12872,N_10348);
or U19843 (N_19843,N_14000,N_13532);
xor U19844 (N_19844,N_13602,N_11550);
xnor U19845 (N_19845,N_14315,N_13030);
or U19846 (N_19846,N_11286,N_12269);
xor U19847 (N_19847,N_10128,N_14040);
nand U19848 (N_19848,N_10024,N_13413);
or U19849 (N_19849,N_12839,N_13160);
nand U19850 (N_19850,N_12612,N_14433);
or U19851 (N_19851,N_10540,N_11215);
and U19852 (N_19852,N_14717,N_12074);
and U19853 (N_19853,N_13076,N_10277);
or U19854 (N_19854,N_13575,N_13198);
and U19855 (N_19855,N_14588,N_10680);
and U19856 (N_19856,N_14570,N_13888);
or U19857 (N_19857,N_10495,N_12180);
nor U19858 (N_19858,N_14782,N_12289);
xor U19859 (N_19859,N_13289,N_14795);
or U19860 (N_19860,N_10514,N_12105);
nor U19861 (N_19861,N_11122,N_11169);
xnor U19862 (N_19862,N_10635,N_13853);
or U19863 (N_19863,N_10634,N_14926);
xor U19864 (N_19864,N_10014,N_11517);
and U19865 (N_19865,N_10393,N_10356);
nor U19866 (N_19866,N_13199,N_12368);
or U19867 (N_19867,N_14088,N_12800);
nand U19868 (N_19868,N_12181,N_14695);
nor U19869 (N_19869,N_10829,N_10108);
nor U19870 (N_19870,N_12411,N_13124);
nor U19871 (N_19871,N_14519,N_13810);
and U19872 (N_19872,N_13651,N_10942);
nand U19873 (N_19873,N_10845,N_12252);
xor U19874 (N_19874,N_14531,N_11751);
xor U19875 (N_19875,N_14173,N_14904);
xnor U19876 (N_19876,N_14573,N_10825);
xor U19877 (N_19877,N_11413,N_13373);
or U19878 (N_19878,N_12981,N_11806);
and U19879 (N_19879,N_14807,N_14126);
or U19880 (N_19880,N_13088,N_14347);
nand U19881 (N_19881,N_11964,N_13927);
and U19882 (N_19882,N_11064,N_11924);
nand U19883 (N_19883,N_13257,N_11041);
and U19884 (N_19884,N_10257,N_10813);
and U19885 (N_19885,N_10793,N_14693);
and U19886 (N_19886,N_13817,N_10323);
nand U19887 (N_19887,N_12764,N_11171);
nand U19888 (N_19888,N_10442,N_10297);
or U19889 (N_19889,N_14528,N_12175);
and U19890 (N_19890,N_11420,N_12836);
nand U19891 (N_19891,N_10628,N_10445);
and U19892 (N_19892,N_10223,N_14055);
nor U19893 (N_19893,N_13639,N_14033);
and U19894 (N_19894,N_11312,N_12048);
and U19895 (N_19895,N_14865,N_11188);
xor U19896 (N_19896,N_13559,N_10952);
nand U19897 (N_19897,N_13341,N_14157);
xor U19898 (N_19898,N_11404,N_10527);
nand U19899 (N_19899,N_12745,N_14933);
xor U19900 (N_19900,N_10449,N_10885);
xnor U19901 (N_19901,N_10704,N_11274);
nor U19902 (N_19902,N_12074,N_10223);
xor U19903 (N_19903,N_13937,N_14741);
xor U19904 (N_19904,N_10701,N_10014);
and U19905 (N_19905,N_11020,N_10471);
nand U19906 (N_19906,N_11146,N_13988);
nor U19907 (N_19907,N_10319,N_13480);
and U19908 (N_19908,N_11704,N_13709);
xnor U19909 (N_19909,N_13240,N_10386);
xnor U19910 (N_19910,N_14292,N_10908);
and U19911 (N_19911,N_10406,N_14837);
xnor U19912 (N_19912,N_12040,N_14596);
nand U19913 (N_19913,N_11411,N_10162);
or U19914 (N_19914,N_13466,N_12546);
or U19915 (N_19915,N_10609,N_10186);
nand U19916 (N_19916,N_10857,N_14771);
nand U19917 (N_19917,N_14317,N_10897);
xor U19918 (N_19918,N_14287,N_14524);
xnor U19919 (N_19919,N_10843,N_10833);
or U19920 (N_19920,N_13135,N_14461);
and U19921 (N_19921,N_13464,N_11641);
nand U19922 (N_19922,N_13687,N_11778);
and U19923 (N_19923,N_13580,N_11364);
nand U19924 (N_19924,N_13624,N_10253);
nor U19925 (N_19925,N_10581,N_10964);
or U19926 (N_19926,N_13003,N_13610);
nor U19927 (N_19927,N_13678,N_10053);
and U19928 (N_19928,N_12088,N_10886);
nand U19929 (N_19929,N_12461,N_11471);
nor U19930 (N_19930,N_13666,N_10277);
or U19931 (N_19931,N_14029,N_10546);
xor U19932 (N_19932,N_10906,N_13693);
xnor U19933 (N_19933,N_13844,N_13204);
or U19934 (N_19934,N_10023,N_11968);
nor U19935 (N_19935,N_10226,N_11230);
xnor U19936 (N_19936,N_12818,N_10854);
nor U19937 (N_19937,N_11181,N_11775);
nor U19938 (N_19938,N_11411,N_10399);
or U19939 (N_19939,N_11068,N_11870);
nor U19940 (N_19940,N_14760,N_12046);
nor U19941 (N_19941,N_14533,N_11873);
xor U19942 (N_19942,N_11458,N_13086);
or U19943 (N_19943,N_13770,N_14654);
or U19944 (N_19944,N_12413,N_12199);
or U19945 (N_19945,N_13680,N_14772);
nand U19946 (N_19946,N_13078,N_14324);
or U19947 (N_19947,N_12495,N_12873);
nand U19948 (N_19948,N_13444,N_11432);
xor U19949 (N_19949,N_12585,N_10361);
and U19950 (N_19950,N_14118,N_13769);
or U19951 (N_19951,N_12574,N_14669);
or U19952 (N_19952,N_11025,N_11022);
nor U19953 (N_19953,N_14394,N_13640);
nand U19954 (N_19954,N_14013,N_13968);
nand U19955 (N_19955,N_13857,N_11019);
nand U19956 (N_19956,N_12111,N_12480);
or U19957 (N_19957,N_12153,N_10038);
nand U19958 (N_19958,N_11806,N_10269);
nand U19959 (N_19959,N_11728,N_12730);
nor U19960 (N_19960,N_13781,N_11003);
and U19961 (N_19961,N_14321,N_11486);
xor U19962 (N_19962,N_14498,N_14178);
xor U19963 (N_19963,N_13154,N_14062);
xnor U19964 (N_19964,N_13338,N_10087);
or U19965 (N_19965,N_12052,N_11964);
nand U19966 (N_19966,N_10623,N_12324);
and U19967 (N_19967,N_13950,N_13237);
nand U19968 (N_19968,N_14005,N_10515);
and U19969 (N_19969,N_14840,N_11336);
or U19970 (N_19970,N_14011,N_13210);
nand U19971 (N_19971,N_12884,N_10530);
nand U19972 (N_19972,N_11758,N_11088);
nor U19973 (N_19973,N_10174,N_12901);
xor U19974 (N_19974,N_13775,N_13098);
nand U19975 (N_19975,N_12260,N_14330);
and U19976 (N_19976,N_14656,N_14010);
nor U19977 (N_19977,N_10436,N_12523);
xor U19978 (N_19978,N_10199,N_13033);
nand U19979 (N_19979,N_13904,N_12899);
and U19980 (N_19980,N_12477,N_10048);
nand U19981 (N_19981,N_13671,N_13384);
or U19982 (N_19982,N_11342,N_12841);
xor U19983 (N_19983,N_13554,N_10953);
nand U19984 (N_19984,N_14841,N_10614);
nor U19985 (N_19985,N_11840,N_10968);
xnor U19986 (N_19986,N_14704,N_12704);
or U19987 (N_19987,N_13509,N_13842);
and U19988 (N_19988,N_14712,N_13605);
or U19989 (N_19989,N_10075,N_12476);
or U19990 (N_19990,N_10882,N_13269);
and U19991 (N_19991,N_12261,N_10041);
nand U19992 (N_19992,N_13898,N_13650);
xor U19993 (N_19993,N_12259,N_11811);
and U19994 (N_19994,N_13853,N_11726);
nor U19995 (N_19995,N_13591,N_10473);
xnor U19996 (N_19996,N_13384,N_11594);
and U19997 (N_19997,N_14444,N_14716);
and U19998 (N_19998,N_10136,N_13101);
or U19999 (N_19999,N_10399,N_13604);
or U20000 (N_20000,N_17438,N_19332);
nor U20001 (N_20001,N_18395,N_15795);
nand U20002 (N_20002,N_18972,N_18575);
and U20003 (N_20003,N_15275,N_16220);
xor U20004 (N_20004,N_17072,N_15497);
and U20005 (N_20005,N_18125,N_16335);
nand U20006 (N_20006,N_16769,N_17393);
nand U20007 (N_20007,N_17725,N_15581);
nand U20008 (N_20008,N_17914,N_17480);
and U20009 (N_20009,N_16307,N_16849);
or U20010 (N_20010,N_19126,N_16576);
xnor U20011 (N_20011,N_16938,N_15096);
or U20012 (N_20012,N_17340,N_15819);
and U20013 (N_20013,N_15638,N_15250);
nor U20014 (N_20014,N_18362,N_18692);
and U20015 (N_20015,N_18416,N_15804);
and U20016 (N_20016,N_15435,N_19453);
nand U20017 (N_20017,N_17614,N_18374);
and U20018 (N_20018,N_16937,N_15583);
nor U20019 (N_20019,N_16908,N_19174);
nor U20020 (N_20020,N_18386,N_18223);
or U20021 (N_20021,N_16579,N_17530);
xor U20022 (N_20022,N_16582,N_15613);
xor U20023 (N_20023,N_17141,N_18045);
and U20024 (N_20024,N_17732,N_18502);
nor U20025 (N_20025,N_18244,N_17039);
xnor U20026 (N_20026,N_15454,N_15786);
nor U20027 (N_20027,N_15157,N_16763);
and U20028 (N_20028,N_17381,N_15646);
nand U20029 (N_20029,N_19208,N_19482);
nor U20030 (N_20030,N_16506,N_16987);
nor U20031 (N_20031,N_19399,N_16215);
nand U20032 (N_20032,N_18171,N_15494);
or U20033 (N_20033,N_17212,N_18151);
nand U20034 (N_20034,N_15088,N_18780);
and U20035 (N_20035,N_19913,N_18616);
xnor U20036 (N_20036,N_16600,N_15046);
nor U20037 (N_20037,N_17851,N_17207);
nor U20038 (N_20038,N_18352,N_16030);
nor U20039 (N_20039,N_19690,N_18378);
or U20040 (N_20040,N_19470,N_17360);
and U20041 (N_20041,N_17861,N_18375);
xor U20042 (N_20042,N_15008,N_18681);
and U20043 (N_20043,N_15632,N_16322);
xor U20044 (N_20044,N_16850,N_16507);
nor U20045 (N_20045,N_15016,N_18269);
xor U20046 (N_20046,N_16602,N_16489);
nor U20047 (N_20047,N_19286,N_16328);
nor U20048 (N_20048,N_17475,N_15884);
and U20049 (N_20049,N_15981,N_19378);
xnor U20050 (N_20050,N_17291,N_19737);
nor U20051 (N_20051,N_17929,N_17432);
nor U20052 (N_20052,N_16567,N_15263);
nor U20053 (N_20053,N_16263,N_18331);
and U20054 (N_20054,N_18825,N_18593);
nand U20055 (N_20055,N_17910,N_17037);
nand U20056 (N_20056,N_15160,N_18700);
or U20057 (N_20057,N_15099,N_17306);
or U20058 (N_20058,N_19140,N_17703);
or U20059 (N_20059,N_16390,N_19664);
nor U20060 (N_20060,N_15251,N_15711);
nand U20061 (N_20061,N_15586,N_19304);
and U20062 (N_20062,N_19112,N_17259);
nand U20063 (N_20063,N_16812,N_15402);
and U20064 (N_20064,N_19864,N_19924);
nand U20065 (N_20065,N_19518,N_19039);
or U20066 (N_20066,N_17024,N_17652);
nor U20067 (N_20067,N_15350,N_15489);
nor U20068 (N_20068,N_17499,N_19160);
nor U20069 (N_20069,N_19407,N_17382);
and U20070 (N_20070,N_17988,N_19083);
and U20071 (N_20071,N_16695,N_18007);
xnor U20072 (N_20072,N_15243,N_15375);
xor U20073 (N_20073,N_17778,N_19299);
xnor U20074 (N_20074,N_16749,N_19561);
or U20075 (N_20075,N_16327,N_18259);
xnor U20076 (N_20076,N_19629,N_17734);
or U20077 (N_20077,N_18071,N_16179);
nor U20078 (N_20078,N_16424,N_17656);
nand U20079 (N_20079,N_18577,N_17273);
and U20080 (N_20080,N_16197,N_17053);
xor U20081 (N_20081,N_16842,N_17045);
or U20082 (N_20082,N_18366,N_17794);
or U20083 (N_20083,N_17253,N_17644);
nor U20084 (N_20084,N_19461,N_15906);
xnor U20085 (N_20085,N_17846,N_15824);
nor U20086 (N_20086,N_19484,N_16133);
or U20087 (N_20087,N_16120,N_18511);
or U20088 (N_20088,N_17174,N_18434);
or U20089 (N_20089,N_17043,N_19581);
nor U20090 (N_20090,N_16866,N_17190);
nand U20091 (N_20091,N_16990,N_16451);
nor U20092 (N_20092,N_19632,N_16712);
xor U20093 (N_20093,N_15078,N_17814);
and U20094 (N_20094,N_15756,N_19305);
nand U20095 (N_20095,N_16187,N_19040);
or U20096 (N_20096,N_16248,N_18124);
nor U20097 (N_20097,N_17669,N_16679);
xor U20098 (N_20098,N_19566,N_18069);
or U20099 (N_20099,N_17631,N_15085);
nor U20100 (N_20100,N_19845,N_19687);
nand U20101 (N_20101,N_16747,N_15066);
nor U20102 (N_20102,N_18288,N_15943);
nor U20103 (N_20103,N_17471,N_15984);
nor U20104 (N_20104,N_16977,N_15641);
or U20105 (N_20105,N_18799,N_16472);
and U20106 (N_20106,N_15109,N_19075);
nor U20107 (N_20107,N_19852,N_19188);
nand U20108 (N_20108,N_15974,N_15865);
and U20109 (N_20109,N_17803,N_19285);
or U20110 (N_20110,N_15691,N_18327);
and U20111 (N_20111,N_15947,N_15635);
nor U20112 (N_20112,N_19171,N_17210);
and U20113 (N_20113,N_17399,N_18879);
or U20114 (N_20114,N_19398,N_17078);
and U20115 (N_20115,N_18443,N_15627);
and U20116 (N_20116,N_17158,N_19206);
nand U20117 (N_20117,N_19143,N_17551);
nand U20118 (N_20118,N_19142,N_19814);
xor U20119 (N_20119,N_17233,N_15098);
and U20120 (N_20120,N_17057,N_15812);
and U20121 (N_20121,N_15068,N_17153);
or U20122 (N_20122,N_16397,N_19015);
and U20123 (N_20123,N_19556,N_15833);
nand U20124 (N_20124,N_17465,N_18026);
nor U20125 (N_20125,N_18721,N_18785);
nand U20126 (N_20126,N_17646,N_16337);
nor U20127 (N_20127,N_16776,N_15619);
nor U20128 (N_20128,N_19485,N_18877);
nor U20129 (N_20129,N_15544,N_17904);
xnor U20130 (N_20130,N_17874,N_18465);
xor U20131 (N_20131,N_18190,N_18381);
nand U20132 (N_20132,N_15216,N_17596);
nor U20133 (N_20133,N_18008,N_17666);
nand U20134 (N_20134,N_15675,N_19988);
and U20135 (N_20135,N_15976,N_19109);
and U20136 (N_20136,N_17654,N_17731);
nor U20137 (N_20137,N_15000,N_15789);
and U20138 (N_20138,N_17785,N_19750);
and U20139 (N_20139,N_15942,N_15441);
and U20140 (N_20140,N_17815,N_16673);
xor U20141 (N_20141,N_18408,N_17941);
and U20142 (N_20142,N_19444,N_18301);
or U20143 (N_20143,N_15241,N_15877);
nand U20144 (N_20144,N_15736,N_16400);
nor U20145 (N_20145,N_17926,N_16874);
and U20146 (N_20146,N_15411,N_17080);
nand U20147 (N_20147,N_15870,N_16268);
xnor U20148 (N_20148,N_15885,N_15103);
xnor U20149 (N_20149,N_16002,N_17224);
and U20150 (N_20150,N_15737,N_16720);
xnor U20151 (N_20151,N_16855,N_19319);
or U20152 (N_20152,N_19134,N_16165);
and U20153 (N_20153,N_15591,N_17554);
nor U20154 (N_20154,N_19231,N_18064);
and U20155 (N_20155,N_17775,N_16562);
or U20156 (N_20156,N_19681,N_16453);
xor U20157 (N_20157,N_17795,N_15432);
nor U20158 (N_20158,N_15939,N_18931);
and U20159 (N_20159,N_17375,N_19094);
xnor U20160 (N_20160,N_19867,N_17012);
or U20161 (N_20161,N_16980,N_19607);
and U20162 (N_20162,N_19584,N_17034);
xnor U20163 (N_20163,N_16645,N_19092);
or U20164 (N_20164,N_17637,N_15805);
or U20165 (N_20165,N_16366,N_18439);
nor U20166 (N_20166,N_16604,N_17966);
nand U20167 (N_20167,N_19099,N_18657);
nor U20168 (N_20168,N_17274,N_19908);
xor U20169 (N_20169,N_19164,N_16707);
and U20170 (N_20170,N_17154,N_17305);
nand U20171 (N_20171,N_16456,N_19834);
xor U20172 (N_20172,N_16641,N_19048);
or U20173 (N_20173,N_15826,N_19106);
and U20174 (N_20174,N_18076,N_16341);
and U20175 (N_20175,N_16279,N_15968);
or U20176 (N_20176,N_18889,N_19595);
nand U20177 (N_20177,N_18903,N_19663);
and U20178 (N_20178,N_17527,N_16206);
and U20179 (N_20179,N_18454,N_15513);
nor U20180 (N_20180,N_16088,N_17925);
nand U20181 (N_20181,N_17780,N_16898);
nor U20182 (N_20182,N_15086,N_19795);
nand U20183 (N_20183,N_19655,N_15121);
or U20184 (N_20184,N_18000,N_17495);
and U20185 (N_20185,N_15816,N_17899);
nand U20186 (N_20186,N_19416,N_18299);
or U20187 (N_20187,N_18963,N_19131);
xor U20188 (N_20188,N_16224,N_18226);
xnor U20189 (N_20189,N_16753,N_19059);
nand U20190 (N_20190,N_18309,N_16156);
nand U20191 (N_20191,N_15470,N_19323);
or U20192 (N_20192,N_17246,N_15897);
and U20193 (N_20193,N_16670,N_19812);
and U20194 (N_20194,N_17576,N_18427);
and U20195 (N_20195,N_18444,N_18099);
and U20196 (N_20196,N_16996,N_15751);
xnor U20197 (N_20197,N_18858,N_17326);
or U20198 (N_20198,N_19382,N_19989);
and U20199 (N_20199,N_17159,N_18129);
nor U20200 (N_20200,N_16677,N_19159);
nor U20201 (N_20201,N_15861,N_19187);
and U20202 (N_20202,N_16967,N_15941);
nand U20203 (N_20203,N_19747,N_15881);
or U20204 (N_20204,N_18498,N_19042);
xnor U20205 (N_20205,N_19239,N_16796);
nor U20206 (N_20206,N_16176,N_16192);
or U20207 (N_20207,N_19771,N_18635);
nor U20208 (N_20208,N_16527,N_15418);
xor U20209 (N_20209,N_19506,N_18974);
nor U20210 (N_20210,N_19216,N_16942);
nor U20211 (N_20211,N_18642,N_16485);
xnor U20212 (N_20212,N_18709,N_16919);
and U20213 (N_20213,N_17130,N_15592);
nand U20214 (N_20214,N_15831,N_16291);
nor U20215 (N_20215,N_18756,N_16803);
and U20216 (N_20216,N_18899,N_18051);
nor U20217 (N_20217,N_17139,N_15719);
and U20218 (N_20218,N_18722,N_15959);
nor U20219 (N_20219,N_19331,N_16635);
or U20220 (N_20220,N_16974,N_17805);
nand U20221 (N_20221,N_19851,N_16563);
xor U20222 (N_20222,N_17423,N_18203);
nand U20223 (N_20223,N_16984,N_16080);
xor U20224 (N_20224,N_16049,N_17201);
and U20225 (N_20225,N_15252,N_18118);
nor U20226 (N_20226,N_18634,N_17738);
nor U20227 (N_20227,N_17541,N_18415);
and U20228 (N_20228,N_16564,N_16816);
xor U20229 (N_20229,N_18316,N_19635);
nor U20230 (N_20230,N_16345,N_16892);
or U20231 (N_20231,N_19272,N_19365);
or U20232 (N_20232,N_15571,N_15305);
and U20233 (N_20233,N_19610,N_16033);
and U20234 (N_20234,N_15873,N_17128);
or U20235 (N_20235,N_18038,N_18512);
nand U20236 (N_20236,N_17807,N_17221);
nor U20237 (N_20237,N_19643,N_18403);
nor U20238 (N_20238,N_15134,N_18941);
nor U20239 (N_20239,N_15945,N_16003);
nand U20240 (N_20240,N_18334,N_19302);
xor U20241 (N_20241,N_17332,N_18543);
xnor U20242 (N_20242,N_16696,N_16698);
nand U20243 (N_20243,N_16168,N_16237);
and U20244 (N_20244,N_17176,N_16151);
nand U20245 (N_20245,N_15633,N_15295);
nor U20246 (N_20246,N_15159,N_15230);
nor U20247 (N_20247,N_15425,N_18370);
and U20248 (N_20248,N_17871,N_15208);
nand U20249 (N_20249,N_15264,N_19978);
nor U20250 (N_20250,N_17492,N_19489);
and U20251 (N_20251,N_15353,N_16417);
xor U20252 (N_20252,N_16655,N_18531);
xnor U20253 (N_20253,N_19275,N_17006);
and U20254 (N_20254,N_18686,N_19904);
xnor U20255 (N_20255,N_19839,N_17730);
nor U20256 (N_20256,N_17044,N_16916);
xnor U20257 (N_20257,N_18246,N_18711);
nand U20258 (N_20258,N_15644,N_18341);
or U20259 (N_20259,N_16543,N_16784);
and U20260 (N_20260,N_17342,N_15142);
nor U20261 (N_20261,N_18845,N_16492);
xnor U20262 (N_20262,N_16123,N_16352);
xor U20263 (N_20263,N_19582,N_15330);
nor U20264 (N_20264,N_17206,N_15965);
nand U20265 (N_20265,N_18310,N_16734);
nand U20266 (N_20266,N_16349,N_16449);
nor U20267 (N_20267,N_15584,N_16137);
nand U20268 (N_20268,N_16947,N_19583);
nand U20269 (N_20269,N_15666,N_15368);
and U20270 (N_20270,N_16330,N_15137);
or U20271 (N_20271,N_15887,N_17869);
or U20272 (N_20272,N_18419,N_15024);
nor U20273 (N_20273,N_16909,N_16791);
and U20274 (N_20274,N_17630,N_15201);
and U20275 (N_20275,N_19500,N_15809);
and U20276 (N_20276,N_16011,N_17142);
nor U20277 (N_20277,N_17888,N_15900);
and U20278 (N_20278,N_15993,N_18535);
nand U20279 (N_20279,N_17515,N_15559);
and U20280 (N_20280,N_17521,N_19822);
xnor U20281 (N_20281,N_15090,N_17028);
xor U20282 (N_20282,N_15191,N_18983);
and U20283 (N_20283,N_18487,N_18919);
and U20284 (N_20284,N_18679,N_18075);
and U20285 (N_20285,N_15808,N_16369);
nand U20286 (N_20286,N_15572,N_15476);
nand U20287 (N_20287,N_18201,N_19574);
nand U20288 (N_20288,N_19598,N_16323);
or U20289 (N_20289,N_19809,N_18414);
xnor U20290 (N_20290,N_17443,N_15154);
nand U20291 (N_20291,N_18844,N_17106);
nor U20292 (N_20292,N_15079,N_17769);
xnor U20293 (N_20293,N_15912,N_18995);
or U20294 (N_20294,N_19009,N_18098);
nor U20295 (N_20295,N_15101,N_16319);
and U20296 (N_20296,N_19150,N_17696);
xnor U20297 (N_20297,N_16583,N_19120);
or U20298 (N_20298,N_17556,N_15317);
nor U20299 (N_20299,N_17565,N_15950);
nor U20300 (N_20300,N_16954,N_17082);
nor U20301 (N_20301,N_17767,N_19511);
and U20302 (N_20302,N_16629,N_15936);
nor U20303 (N_20303,N_16886,N_17557);
or U20304 (N_20304,N_18472,N_16353);
and U20305 (N_20305,N_19668,N_19316);
nand U20306 (N_20306,N_15240,N_19135);
and U20307 (N_20307,N_15962,N_16493);
and U20308 (N_20308,N_18985,N_17651);
or U20309 (N_20309,N_15662,N_17401);
or U20310 (N_20310,N_16797,N_15143);
or U20311 (N_20311,N_15612,N_16570);
or U20312 (N_20312,N_19127,N_16683);
and U20313 (N_20313,N_19800,N_16068);
or U20314 (N_20314,N_18939,N_16218);
nand U20315 (N_20315,N_16173,N_17096);
nor U20316 (N_20316,N_19027,N_18878);
and U20317 (N_20317,N_15025,N_17473);
xor U20318 (N_20318,N_19066,N_16839);
nor U20319 (N_20319,N_18032,N_16031);
or U20320 (N_20320,N_17107,N_19395);
xor U20321 (N_20321,N_17486,N_19569);
xnor U20322 (N_20322,N_19789,N_16672);
nor U20323 (N_20323,N_16304,N_18364);
nand U20324 (N_20324,N_16549,N_19963);
xor U20325 (N_20325,N_16025,N_18451);
xnor U20326 (N_20326,N_19955,N_19038);
and U20327 (N_20327,N_17531,N_15127);
xnor U20328 (N_20328,N_16568,N_16910);
xnor U20329 (N_20329,N_15339,N_18441);
and U20330 (N_20330,N_15080,N_15533);
and U20331 (N_20331,N_19758,N_16084);
and U20332 (N_20332,N_19707,N_16415);
nor U20333 (N_20333,N_15554,N_16962);
nand U20334 (N_20334,N_17774,N_17897);
and U20335 (N_20335,N_16281,N_18435);
nand U20336 (N_20336,N_15791,N_16768);
or U20337 (N_20337,N_15963,N_15729);
xnor U20338 (N_20338,N_15651,N_16950);
or U20339 (N_20339,N_17574,N_19163);
and U20340 (N_20340,N_16346,N_18705);
nand U20341 (N_20341,N_16101,N_18927);
and U20342 (N_20342,N_17365,N_16370);
and U20343 (N_20343,N_19090,N_15175);
xor U20344 (N_20344,N_17783,N_18815);
nor U20345 (N_20345,N_18908,N_18503);
xnor U20346 (N_20346,N_15714,N_15565);
or U20347 (N_20347,N_15184,N_16975);
and U20348 (N_20348,N_15899,N_18569);
nand U20349 (N_20349,N_19446,N_16789);
nor U20350 (N_20350,N_18034,N_17667);
or U20351 (N_20351,N_17972,N_15033);
xor U20352 (N_20352,N_18514,N_16100);
xor U20353 (N_20353,N_15130,N_17655);
xor U20354 (N_20354,N_16648,N_17507);
or U20355 (N_20355,N_17835,N_17996);
xor U20356 (N_20356,N_17995,N_15952);
nor U20357 (N_20357,N_16065,N_19105);
and U20358 (N_20358,N_19424,N_15862);
xnor U20359 (N_20359,N_18275,N_19937);
nor U20360 (N_20360,N_18023,N_18716);
xor U20361 (N_20361,N_16536,N_16627);
or U20362 (N_20362,N_15163,N_17884);
or U20363 (N_20363,N_15074,N_18518);
and U20364 (N_20364,N_18956,N_18238);
or U20365 (N_20365,N_19894,N_17035);
xor U20366 (N_20366,N_19145,N_16053);
or U20367 (N_20367,N_19890,N_16717);
nand U20368 (N_20368,N_15994,N_18563);
xor U20369 (N_20369,N_15469,N_17810);
xnor U20370 (N_20370,N_16300,N_15828);
and U20371 (N_20371,N_16716,N_16216);
nor U20372 (N_20372,N_16535,N_17601);
nor U20373 (N_20373,N_18971,N_17297);
nor U20374 (N_20374,N_18738,N_19396);
and U20375 (N_20375,N_19405,N_17817);
nand U20376 (N_20376,N_15466,N_15672);
nand U20377 (N_20377,N_17196,N_17101);
nand U20378 (N_20378,N_19880,N_15656);
xnor U20379 (N_20379,N_15563,N_15311);
xnor U20380 (N_20380,N_17674,N_16952);
and U20381 (N_20381,N_17735,N_18942);
nand U20382 (N_20382,N_16110,N_16588);
nor U20383 (N_20383,N_15189,N_19480);
nor U20384 (N_20384,N_15307,N_16209);
xor U20385 (N_20385,N_16982,N_15111);
or U20386 (N_20386,N_16409,N_19290);
xor U20387 (N_20387,N_19261,N_19197);
xor U20388 (N_20388,N_18794,N_15510);
nand U20389 (N_20389,N_19732,N_19225);
and U20390 (N_20390,N_17881,N_18804);
xor U20391 (N_20391,N_19454,N_17203);
nand U20392 (N_20392,N_16912,N_17061);
nand U20393 (N_20393,N_19706,N_19630);
and U20394 (N_20394,N_15539,N_15829);
nand U20395 (N_20395,N_19141,N_18774);
or U20396 (N_20396,N_15686,N_17093);
nor U20397 (N_20397,N_16070,N_16143);
nor U20398 (N_20398,N_19775,N_18533);
and U20399 (N_20399,N_15126,N_17388);
and U20400 (N_20400,N_18687,N_19226);
nor U20401 (N_20401,N_15723,N_19199);
nand U20402 (N_20402,N_15355,N_15859);
or U20403 (N_20403,N_19406,N_16112);
nor U20404 (N_20404,N_19786,N_15265);
and U20405 (N_20405,N_16085,N_19169);
and U20406 (N_20406,N_15601,N_17252);
xnor U20407 (N_20407,N_15215,N_19601);
and U20408 (N_20408,N_16907,N_16018);
xor U20409 (N_20409,N_16636,N_15938);
or U20410 (N_20410,N_17430,N_17310);
xnor U20411 (N_20411,N_19397,N_16838);
nor U20412 (N_20412,N_17880,N_17526);
nand U20413 (N_20413,N_15648,N_16766);
and U20414 (N_20414,N_16879,N_19847);
xor U20415 (N_20415,N_18207,N_18909);
and U20416 (N_20416,N_19223,N_15594);
and U20417 (N_20417,N_19350,N_16693);
nand U20418 (N_20418,N_17315,N_18752);
nor U20419 (N_20419,N_17325,N_16444);
or U20420 (N_20420,N_15058,N_16230);
nand U20421 (N_20421,N_18528,N_18139);
or U20422 (N_20422,N_19773,N_19958);
and U20423 (N_20423,N_19412,N_19028);
nand U20424 (N_20424,N_18240,N_19073);
nor U20425 (N_20425,N_19428,N_19389);
or U20426 (N_20426,N_19578,N_17192);
or U20427 (N_20427,N_15660,N_18052);
xnor U20428 (N_20428,N_19268,N_19976);
and U20429 (N_20429,N_15203,N_15561);
nand U20430 (N_20430,N_15420,N_16392);
and U20431 (N_20431,N_16212,N_17915);
xor U20432 (N_20432,N_17514,N_18406);
and U20433 (N_20433,N_18148,N_19493);
or U20434 (N_20434,N_16733,N_18729);
xnor U20435 (N_20435,N_19155,N_15763);
or U20436 (N_20436,N_15503,N_17434);
and U20437 (N_20437,N_19052,N_19183);
and U20438 (N_20438,N_18773,N_19486);
nor U20439 (N_20439,N_15610,N_16571);
xnor U20440 (N_20440,N_15212,N_18142);
and U20441 (N_20441,N_15224,N_19981);
nor U20442 (N_20442,N_19563,N_15290);
or U20443 (N_20443,N_18954,N_19759);
xor U20444 (N_20444,N_19118,N_19766);
nor U20445 (N_20445,N_18935,N_19280);
nand U20446 (N_20446,N_18306,N_16483);
nand U20447 (N_20447,N_15574,N_19861);
and U20448 (N_20448,N_18629,N_17249);
xnor U20449 (N_20449,N_18585,N_17793);
and U20450 (N_20450,N_19572,N_18957);
xor U20451 (N_20451,N_18996,N_15720);
nand U20452 (N_20452,N_19019,N_19338);
and U20453 (N_20453,N_19125,N_18473);
nor U20454 (N_20454,N_16280,N_15585);
nand U20455 (N_20455,N_17208,N_19430);
nand U20456 (N_20456,N_18633,N_15905);
and U20457 (N_20457,N_16804,N_16373);
nand U20458 (N_20458,N_19368,N_16959);
nor U20459 (N_20459,N_15433,N_19877);
xor U20460 (N_20460,N_16376,N_15374);
and U20461 (N_20461,N_17197,N_17209);
nand U20462 (N_20462,N_19097,N_19599);
nor U20463 (N_20463,N_16873,N_15760);
xnor U20464 (N_20464,N_17337,N_16930);
nand U20465 (N_20465,N_18311,N_18833);
nor U20466 (N_20466,N_16701,N_17427);
nand U20467 (N_20467,N_19673,N_19785);
nor U20468 (N_20468,N_18732,N_19128);
xnor U20469 (N_20469,N_16667,N_18183);
nor U20470 (N_20470,N_18222,N_16454);
and U20471 (N_20471,N_17503,N_19520);
or U20472 (N_20472,N_19311,N_19242);
nor U20473 (N_20473,N_17216,N_17917);
nor U20474 (N_20474,N_17765,N_15128);
xnor U20475 (N_20475,N_17855,N_18807);
nor U20476 (N_20476,N_15937,N_15615);
nor U20477 (N_20477,N_18425,N_19526);
or U20478 (N_20478,N_18191,N_18164);
nand U20479 (N_20479,N_15838,N_18614);
xor U20480 (N_20480,N_16458,N_17701);
xnor U20481 (N_20481,N_19529,N_15570);
xor U20482 (N_20482,N_16028,N_17419);
or U20483 (N_20483,N_17277,N_15582);
nor U20484 (N_20484,N_17322,N_16198);
xor U20485 (N_20485,N_16332,N_17251);
or U20486 (N_20486,N_16214,N_16069);
nor U20487 (N_20487,N_16964,N_17245);
xor U20488 (N_20488,N_16097,N_19494);
or U20489 (N_20489,N_19445,N_18644);
nor U20490 (N_20490,N_17281,N_17830);
nor U20491 (N_20491,N_19589,N_19096);
nor U20492 (N_20492,N_17369,N_17612);
xnor U20493 (N_20493,N_18035,N_19604);
nor U20494 (N_20494,N_18250,N_18955);
or U20495 (N_20495,N_16826,N_18280);
xor U20496 (N_20496,N_15269,N_15495);
nor U20497 (N_20497,N_15524,N_15314);
and U20498 (N_20498,N_19436,N_17955);
or U20499 (N_20499,N_17300,N_16587);
nand U20500 (N_20500,N_16978,N_15661);
or U20501 (N_20501,N_19342,N_15765);
nand U20502 (N_20502,N_15391,N_16480);
xnor U20503 (N_20503,N_19863,N_19693);
nor U20504 (N_20504,N_18856,N_19644);
and U20505 (N_20505,N_19247,N_16094);
or U20506 (N_20506,N_18237,N_16722);
or U20507 (N_20507,N_15966,N_17750);
xnor U20508 (N_20508,N_19548,N_19071);
nand U20509 (N_20509,N_17714,N_18335);
nor U20510 (N_20510,N_18278,N_18631);
nor U20511 (N_20511,N_16945,N_18611);
xnor U20512 (N_20512,N_18279,N_16546);
or U20513 (N_20513,N_15842,N_16460);
nor U20514 (N_20514,N_16994,N_17927);
or U20515 (N_20515,N_15455,N_15929);
nor U20516 (N_20516,N_16482,N_15580);
nand U20517 (N_20517,N_17125,N_16131);
xnor U20518 (N_20518,N_16043,N_17126);
xor U20519 (N_20519,N_17566,N_19296);
or U20520 (N_20520,N_19712,N_15461);
and U20521 (N_20521,N_16423,N_16277);
xor U20522 (N_20522,N_18430,N_16552);
or U20523 (N_20523,N_18161,N_18177);
xnor U20524 (N_20524,N_19472,N_19119);
nor U20525 (N_20525,N_17813,N_16073);
xor U20526 (N_20526,N_15507,N_16022);
nor U20527 (N_20527,N_16762,N_15268);
nor U20528 (N_20528,N_18477,N_19661);
xor U20529 (N_20529,N_17356,N_19914);
xnor U20530 (N_20530,N_17877,N_18276);
nand U20531 (N_20531,N_17677,N_17323);
xor U20532 (N_20532,N_15379,N_15071);
xor U20533 (N_20533,N_17602,N_19537);
and U20534 (N_20534,N_16985,N_19952);
xor U20535 (N_20535,N_16751,N_18938);
or U20536 (N_20536,N_18663,N_19440);
nand U20537 (N_20537,N_15598,N_15110);
xnor U20538 (N_20538,N_18777,N_19373);
and U20539 (N_20539,N_17095,N_15850);
or U20540 (N_20540,N_16878,N_18329);
and U20541 (N_20541,N_19815,N_15112);
or U20542 (N_20542,N_16194,N_15185);
or U20543 (N_20543,N_17230,N_19767);
and U20544 (N_20544,N_15035,N_15548);
or U20545 (N_20545,N_19209,N_16888);
xor U20546 (N_20546,N_17071,N_18597);
nand U20547 (N_20547,N_16809,N_16481);
nand U20548 (N_20548,N_15386,N_19306);
nand U20549 (N_20549,N_19091,N_18049);
or U20550 (N_20550,N_17736,N_17358);
nand U20551 (N_20551,N_15405,N_18840);
and U20552 (N_20552,N_19917,N_18336);
and U20553 (N_20553,N_19799,N_19002);
xor U20554 (N_20554,N_18819,N_19794);
xnor U20555 (N_20555,N_15915,N_19315);
nor U20556 (N_20556,N_16282,N_19699);
nand U20557 (N_20557,N_18524,N_18295);
nand U20558 (N_20558,N_19464,N_19902);
nand U20559 (N_20559,N_19431,N_19927);
xor U20560 (N_20560,N_19999,N_19069);
nor U20561 (N_20561,N_16316,N_18656);
and U20562 (N_20562,N_17762,N_19666);
nor U20563 (N_20563,N_16226,N_16617);
nand U20564 (N_20564,N_16724,N_18229);
nor U20565 (N_20565,N_18688,N_19692);
and U20566 (N_20566,N_17011,N_19512);
nor U20567 (N_20567,N_15556,N_15650);
or U20568 (N_20568,N_19817,N_19269);
xor U20569 (N_20569,N_15879,N_19628);
or U20570 (N_20570,N_16664,N_19915);
nand U20571 (N_20571,N_15534,N_18233);
nand U20572 (N_20572,N_18489,N_15464);
xor U20573 (N_20573,N_15682,N_15499);
nor U20574 (N_20574,N_19603,N_15232);
or U20575 (N_20575,N_18483,N_19103);
nand U20576 (N_20576,N_15320,N_15274);
xnor U20577 (N_20577,N_19483,N_17218);
and U20578 (N_20578,N_15562,N_18652);
nor U20579 (N_20579,N_16616,N_19920);
nor U20580 (N_20580,N_15385,N_16391);
and U20581 (N_20581,N_16668,N_16737);
nor U20582 (N_20582,N_17699,N_17478);
nor U20583 (N_20583,N_18736,N_19035);
nor U20584 (N_20584,N_18286,N_17550);
or U20585 (N_20585,N_19810,N_19860);
nor U20586 (N_20586,N_18485,N_18422);
or U20587 (N_20587,N_15589,N_15625);
or U20588 (N_20588,N_18172,N_18636);
xnor U20589 (N_20589,N_19818,N_15056);
nor U20590 (N_20590,N_16380,N_19029);
nand U20591 (N_20591,N_19702,N_17103);
or U20592 (N_20592,N_18554,N_19393);
or U20593 (N_20593,N_15748,N_17491);
and U20594 (N_20594,N_16399,N_16278);
nand U20595 (N_20595,N_18852,N_18116);
or U20596 (N_20596,N_18429,N_18730);
and U20597 (N_20597,N_18361,N_17352);
or U20598 (N_20598,N_16502,N_18496);
or U20599 (N_20599,N_17711,N_16265);
and U20600 (N_20600,N_15673,N_17826);
and U20601 (N_20601,N_19391,N_17608);
xnor U20602 (N_20602,N_15182,N_17016);
and U20603 (N_20603,N_19068,N_18011);
nand U20604 (N_20604,N_16993,N_16694);
or U20605 (N_20605,N_18220,N_18111);
and U20606 (N_20606,N_18015,N_16711);
nor U20607 (N_20607,N_17758,N_16862);
or U20608 (N_20608,N_18432,N_16815);
or U20609 (N_20609,N_17618,N_15902);
and U20610 (N_20610,N_18495,N_16859);
nor U20611 (N_20611,N_19195,N_16473);
or U20612 (N_20612,N_17148,N_17999);
or U20613 (N_20613,N_19297,N_16231);
xnor U20614 (N_20614,N_15634,N_19662);
or U20615 (N_20615,N_16183,N_16933);
and U20616 (N_20616,N_16594,N_15542);
xnor U20617 (N_20617,N_15444,N_16633);
xnor U20618 (N_20618,N_15106,N_16609);
and U20619 (N_20619,N_16150,N_16295);
nor U20620 (N_20620,N_15172,N_16246);
nand U20621 (N_20621,N_18167,N_15985);
and U20622 (N_20622,N_16525,N_15220);
and U20623 (N_20623,N_16624,N_18864);
nor U20624 (N_20624,N_18902,N_18070);
nand U20625 (N_20625,N_17700,N_18493);
xnor U20626 (N_20626,N_19997,N_16271);
xnor U20627 (N_20627,N_15063,N_18224);
and U20628 (N_20628,N_16309,N_17119);
nand U20629 (N_20629,N_17578,N_17470);
and U20630 (N_20630,N_18086,N_19022);
xnor U20631 (N_20631,N_15266,N_18211);
or U20632 (N_20632,N_18270,N_19570);
nand U20633 (N_20633,N_18782,N_18816);
nand U20634 (N_20634,N_15349,N_18480);
xor U20635 (N_20635,N_15999,N_19946);
nor U20636 (N_20636,N_18789,N_17193);
xnor U20637 (N_20637,N_18580,N_18952);
nor U20638 (N_20638,N_17607,N_15055);
and U20639 (N_20639,N_16389,N_19432);
xor U20640 (N_20640,N_16310,N_16432);
nor U20641 (N_20641,N_16596,N_17050);
nor U20642 (N_20642,N_18982,N_16394);
and U20643 (N_20643,N_17435,N_15827);
nor U20644 (N_20644,N_18453,N_15926);
and U20645 (N_20645,N_15231,N_17186);
nor U20646 (N_20646,N_18841,N_16652);
or U20647 (N_20647,N_16505,N_18558);
or U20648 (N_20648,N_16169,N_16963);
nor U20649 (N_20649,N_15930,N_15097);
xnor U20650 (N_20650,N_16026,N_18993);
nand U20651 (N_20651,N_19542,N_16038);
nor U20652 (N_20652,N_19985,N_19949);
nand U20653 (N_20653,N_19696,N_15649);
or U20654 (N_20654,N_17553,N_16443);
nor U20655 (N_20655,N_15597,N_16190);
and U20656 (N_20656,N_16884,N_17820);
nand U20657 (N_20657,N_17353,N_19728);
nor U20658 (N_20658,N_16808,N_15132);
xor U20659 (N_20659,N_16852,N_15023);
xnor U20660 (N_20660,N_15781,N_16960);
xnor U20661 (N_20661,N_19326,N_19243);
nand U20662 (N_20662,N_17560,N_17916);
and U20663 (N_20663,N_17453,N_18192);
and U20664 (N_20664,N_15752,N_19961);
nand U20665 (N_20665,N_16051,N_15034);
nand U20666 (N_20666,N_18714,N_18765);
or U20667 (N_20667,N_18043,N_16755);
nand U20668 (N_20668,N_18591,N_19552);
or U20669 (N_20669,N_18751,N_19611);
xnor U20670 (N_20670,N_18258,N_16378);
xnor U20671 (N_20671,N_16740,N_18849);
or U20672 (N_20672,N_17009,N_15095);
nor U20673 (N_20673,N_16440,N_19654);
xor U20674 (N_20674,N_15690,N_18987);
or U20675 (N_20675,N_15329,N_16523);
or U20676 (N_20676,N_18622,N_17963);
xor U20677 (N_20677,N_15693,N_17001);
nand U20678 (N_20678,N_19364,N_17304);
or U20679 (N_20679,N_15479,N_19928);
and U20680 (N_20680,N_18552,N_17373);
or U20681 (N_20681,N_19051,N_17284);
xnor U20682 (N_20682,N_18886,N_15529);
or U20683 (N_20683,N_15310,N_18085);
and U20684 (N_20684,N_19376,N_16007);
xor U20685 (N_20685,N_19683,N_15322);
xnor U20686 (N_20686,N_18638,N_18459);
nor U20687 (N_20687,N_17739,N_16621);
and U20688 (N_20688,N_15958,N_19234);
nand U20689 (N_20689,N_16853,N_15049);
xnor U20690 (N_20690,N_15011,N_16467);
xnor U20691 (N_20691,N_17286,N_16188);
xor U20692 (N_20692,N_17876,N_15249);
nor U20693 (N_20693,N_18605,N_19903);
xor U20694 (N_20694,N_19176,N_15400);
and U20695 (N_20695,N_17879,N_19760);
or U20696 (N_20696,N_17385,N_17529);
and U20697 (N_20697,N_19554,N_18028);
and U20698 (N_20698,N_15370,N_15626);
or U20699 (N_20699,N_16461,N_16625);
or U20700 (N_20700,N_17087,N_17671);
or U20701 (N_20701,N_19944,N_15478);
or U20702 (N_20702,N_17688,N_15136);
xor U20703 (N_20703,N_19442,N_15467);
and U20704 (N_20704,N_16508,N_18092);
or U20705 (N_20705,N_16012,N_17609);
nor U20706 (N_20706,N_18741,N_19749);
xnor U20707 (N_20707,N_18670,N_18097);
or U20708 (N_20708,N_15849,N_18596);
and U20709 (N_20709,N_15787,N_15335);
or U20710 (N_20710,N_19855,N_19597);
xor U20711 (N_20711,N_18242,N_19361);
or U20712 (N_20712,N_15807,N_19005);
nor U20713 (N_20713,N_18468,N_16250);
xnor U20714 (N_20714,N_19129,N_18448);
nand U20715 (N_20715,N_15170,N_15694);
or U20716 (N_20716,N_15778,N_15652);
and U20717 (N_20717,N_15239,N_19729);
and U20718 (N_20718,N_18389,N_15659);
nand U20719 (N_20719,N_15026,N_19359);
nand U20720 (N_20720,N_17363,N_19330);
nand U20721 (N_20721,N_17479,N_16294);
nand U20722 (N_20722,N_16869,N_19152);
nor U20723 (N_20723,N_18517,N_16306);
nand U20724 (N_20724,N_18134,N_17663);
xnor U20725 (N_20725,N_18297,N_19682);
nor U20726 (N_20726,N_19372,N_15917);
nand U20727 (N_20727,N_15642,N_16243);
nor U20728 (N_20728,N_16713,N_18959);
and U20729 (N_20729,N_19856,N_16802);
xor U20730 (N_20730,N_18317,N_17720);
nand U20731 (N_20731,N_18355,N_16560);
nand U20732 (N_20732,N_18411,N_19166);
xnor U20733 (N_20733,N_17098,N_15039);
or U20734 (N_20734,N_19335,N_17535);
xor U20735 (N_20735,N_19259,N_15568);
xnor U20736 (N_20736,N_17328,N_16781);
and U20737 (N_20737,N_18981,N_18772);
and U20738 (N_20738,N_18992,N_18904);
nand U20739 (N_20739,N_17127,N_18146);
nand U20740 (N_20740,N_17187,N_17600);
nor U20741 (N_20741,N_17394,N_19726);
nand U20742 (N_20742,N_19633,N_18968);
or U20743 (N_20743,N_17500,N_15604);
nor U20744 (N_20744,N_17215,N_18961);
and U20745 (N_20745,N_18775,N_19782);
nand U20746 (N_20746,N_19363,N_15797);
nand U20747 (N_20747,N_18475,N_19990);
or U20748 (N_20748,N_16767,N_18321);
nor U20749 (N_20749,N_17684,N_15587);
xor U20750 (N_20750,N_17288,N_15458);
xor U20751 (N_20751,N_18186,N_18758);
or U20752 (N_20752,N_15131,N_16222);
or U20753 (N_20753,N_16611,N_18156);
and U20754 (N_20754,N_16058,N_15194);
nor U20755 (N_20755,N_16684,N_18771);
or U20756 (N_20756,N_18025,N_15472);
and U20757 (N_20757,N_17073,N_15259);
nand U20758 (N_20758,N_18354,N_16210);
nor U20759 (N_20759,N_19993,N_19972);
nand U20760 (N_20760,N_15308,N_16160);
nor U20761 (N_20761,N_17463,N_17374);
nand U20762 (N_20762,N_16372,N_16067);
nand U20763 (N_20763,N_18109,N_16810);
xnor U20764 (N_20764,N_15342,N_16072);
xnor U20765 (N_20765,N_16823,N_19032);
or U20766 (N_20766,N_19341,N_17886);
nand U20767 (N_20767,N_15073,N_18147);
nor U20768 (N_20768,N_19776,N_19701);
nor U20769 (N_20769,N_15417,N_16266);
nor U20770 (N_20770,N_16213,N_17635);
or U20771 (N_20771,N_19355,N_15825);
nor U20772 (N_20772,N_19254,N_19139);
nor U20773 (N_20773,N_19317,N_15173);
nor U20774 (N_20774,N_18655,N_18728);
or U20775 (N_20775,N_17267,N_17355);
or U20776 (N_20776,N_18128,N_18353);
or U20777 (N_20777,N_18458,N_17719);
and U20778 (N_20778,N_19474,N_18544);
or U20779 (N_20779,N_18140,N_15683);
xnor U20780 (N_20780,N_17474,N_19201);
or U20781 (N_20781,N_18157,N_19218);
nand U20782 (N_20782,N_16728,N_15798);
and U20783 (N_20783,N_18205,N_15818);
nand U20784 (N_20784,N_18505,N_16413);
or U20785 (N_20785,N_16557,N_15313);
or U20786 (N_20786,N_16702,N_17439);
and U20787 (N_20787,N_18087,N_17942);
nor U20788 (N_20788,N_18304,N_17512);
or U20789 (N_20789,N_18977,N_15438);
xor U20790 (N_20790,N_18784,N_17235);
and U20791 (N_20791,N_15631,N_16398);
or U20792 (N_20792,N_19891,N_18407);
or U20793 (N_20793,N_19813,N_19715);
xnor U20794 (N_20794,N_18615,N_17990);
nor U20795 (N_20795,N_18463,N_16495);
and U20796 (N_20796,N_17962,N_19402);
nand U20797 (N_20797,N_16738,N_16175);
and U20798 (N_20798,N_15223,N_17658);
nor U20799 (N_20799,N_18519,N_17105);
nand U20800 (N_20800,N_16688,N_19536);
xor U20801 (N_20801,N_15210,N_17403);
nand U20802 (N_20802,N_19354,N_19148);
xnor U20803 (N_20803,N_19144,N_16761);
nand U20804 (N_20804,N_18060,N_18783);
and U20805 (N_20805,N_18870,N_18625);
nor U20806 (N_20806,N_16537,N_18228);
nor U20807 (N_20807,N_18821,N_16887);
nor U20808 (N_20808,N_18742,N_17308);
nand U20809 (N_20809,N_16127,N_17488);
nor U20810 (N_20810,N_16860,N_19034);
nor U20811 (N_20811,N_16401,N_15316);
xor U20812 (N_20812,N_16500,N_15813);
nand U20813 (N_20813,N_18236,N_17983);
xnor U20814 (N_20814,N_19467,N_15640);
or U20815 (N_20815,N_15995,N_17961);
nand U20816 (N_20816,N_18057,N_18294);
or U20817 (N_20817,N_18433,N_17448);
nor U20818 (N_20818,N_15853,N_17561);
nand U20819 (N_20819,N_18997,N_19806);
nand U20820 (N_20820,N_19044,N_15176);
xor U20821 (N_20821,N_19862,N_19865);
nor U20822 (N_20822,N_18491,N_17889);
and U20823 (N_20823,N_15409,N_16178);
and U20824 (N_20824,N_19527,N_17449);
xnor U20825 (N_20825,N_17653,N_17191);
nor U20826 (N_20826,N_17108,N_18159);
or U20827 (N_20827,N_15536,N_19672);
or U20828 (N_20828,N_18578,N_18267);
xor U20829 (N_20829,N_19616,N_15480);
or U20830 (N_20830,N_19264,N_18947);
or U20831 (N_20831,N_17636,N_15992);
xor U20832 (N_20832,N_18016,N_15260);
nor U20833 (N_20833,N_16119,N_16682);
or U20834 (N_20834,N_15091,N_15286);
nor U20835 (N_20835,N_16538,N_16727);
nand U20836 (N_20836,N_19626,N_16877);
xor U20837 (N_20837,N_16425,N_18174);
and U20838 (N_20838,N_19846,N_17268);
nand U20839 (N_20839,N_16772,N_19240);
and U20840 (N_20840,N_16921,N_18813);
nor U20841 (N_20841,N_17086,N_18302);
xnor U20842 (N_20842,N_19764,N_19752);
or U20843 (N_20843,N_17241,N_16819);
or U20844 (N_20844,N_17865,N_19130);
xnor U20845 (N_20845,N_19115,N_16584);
nor U20846 (N_20846,N_16699,N_17217);
nor U20847 (N_20847,N_19433,N_15371);
nand U20848 (N_20848,N_17490,N_17939);
and U20849 (N_20849,N_17791,N_19213);
or U20850 (N_20850,N_15141,N_18937);
and U20851 (N_20851,N_16238,N_17264);
and U20852 (N_20852,N_16411,N_19191);
and U20853 (N_20853,N_17664,N_17951);
and U20854 (N_20854,N_19777,N_16039);
nor U20855 (N_20855,N_18102,N_15758);
nor U20856 (N_20856,N_17675,N_18488);
and U20857 (N_20857,N_15306,N_19741);
xnor U20858 (N_20858,N_18456,N_15990);
xor U20859 (N_20859,N_18628,N_15738);
nor U20860 (N_20860,N_18158,N_15713);
xnor U20861 (N_20861,N_15543,N_18504);
and U20862 (N_20862,N_19910,N_15338);
nand U20863 (N_20863,N_18497,N_15971);
or U20864 (N_20864,N_15204,N_16090);
and U20865 (N_20865,N_17661,N_17633);
and U20866 (N_20866,N_16968,N_16329);
and U20867 (N_20867,N_19057,N_18573);
xnor U20868 (N_20868,N_15779,N_19455);
and U20869 (N_20869,N_16419,N_15357);
and U20870 (N_20870,N_19441,N_16628);
nand U20871 (N_20871,N_19892,N_17766);
and U20872 (N_20872,N_19838,N_17694);
and U20873 (N_20873,N_15334,N_17166);
nand U20874 (N_20874,N_17276,N_15717);
nor U20875 (N_20875,N_18936,N_15505);
or U20876 (N_20876,N_15679,N_16517);
nand U20877 (N_20877,N_15312,N_18464);
and U20878 (N_20878,N_15727,N_15567);
nand U20879 (N_20879,N_19992,N_19205);
xnor U20880 (N_20880,N_17704,N_15578);
xor U20881 (N_20881,N_18138,N_16359);
nor U20882 (N_20882,N_17184,N_19987);
nor U20883 (N_20883,N_17524,N_15983);
or U20884 (N_20884,N_15007,N_19000);
xnor U20885 (N_20885,N_19642,N_18770);
xnor U20886 (N_20886,N_15732,N_15323);
nand U20887 (N_20887,N_17338,N_15235);
and U20888 (N_20888,N_18719,N_16714);
nand U20889 (N_20889,N_17200,N_18617);
xnor U20890 (N_20890,N_17248,N_16060);
nor U20891 (N_20891,N_15219,N_18632);
and U20892 (N_20892,N_19836,N_19550);
and U20893 (N_20893,N_17414,N_18713);
or U20894 (N_20894,N_16433,N_15407);
or U20895 (N_20895,N_19640,N_16124);
nor U20896 (N_20896,N_15383,N_19866);
and U20897 (N_20897,N_16554,N_18896);
xor U20898 (N_20898,N_18307,N_16706);
nand U20899 (N_20899,N_16245,N_18749);
nor U20900 (N_20900,N_15852,N_18602);
or U20901 (N_20901,N_19893,N_19070);
and U20902 (N_20902,N_18893,N_18506);
xnor U20903 (N_20903,N_16903,N_18666);
and U20904 (N_20904,N_16368,N_15643);
and U20905 (N_20905,N_16745,N_19021);
nor U20906 (N_20906,N_15378,N_17952);
or U20907 (N_20907,N_18900,N_18053);
and U20908 (N_20908,N_18283,N_18873);
nand U20909 (N_20909,N_15856,N_16340);
nand U20910 (N_20910,N_19101,N_19887);
or U20911 (N_20911,N_19637,N_15577);
and U20912 (N_20912,N_17898,N_16997);
and U20913 (N_20913,N_15015,N_17377);
and U20914 (N_20914,N_17429,N_19658);
and U20915 (N_20915,N_16759,N_16824);
nand U20916 (N_20916,N_17536,N_15940);
or U20917 (N_20917,N_19524,N_15115);
nand U20918 (N_20918,N_18476,N_16800);
nor U20919 (N_20919,N_17025,N_19279);
and U20920 (N_20920,N_16649,N_18723);
or U20921 (N_20921,N_18779,N_17506);
nor U20922 (N_20922,N_15924,N_18894);
or U20923 (N_20923,N_19532,N_19568);
xnor U20924 (N_20924,N_19965,N_16788);
xnor U20925 (N_20925,N_19964,N_18200);
nand U20926 (N_20926,N_18871,N_17017);
nor U20927 (N_20927,N_18412,N_17513);
or U20928 (N_20928,N_15273,N_19671);
nor U20929 (N_20929,N_16741,N_18746);
xor U20930 (N_20930,N_18926,N_16420);
or U20931 (N_20931,N_19170,N_17391);
or U20932 (N_20932,N_16431,N_18262);
xnor U20933 (N_20933,N_16820,N_19872);
nor U20934 (N_20934,N_18958,N_19688);
xnor U20935 (N_20935,N_19623,N_16503);
xor U20936 (N_20936,N_17483,N_19345);
or U20937 (N_20937,N_19189,N_18768);
nor U20938 (N_20938,N_17542,N_19745);
nor U20939 (N_20939,N_16793,N_16157);
or U20940 (N_20940,N_17572,N_19956);
nand U20941 (N_20941,N_17319,N_17969);
nor U20942 (N_20942,N_17410,N_18834);
and U20943 (N_20943,N_17998,N_15309);
nand U20944 (N_20944,N_15869,N_17872);
or U20945 (N_20945,N_19606,N_17645);
xnor U20946 (N_20946,N_17058,N_17975);
or U20947 (N_20947,N_16144,N_18546);
nor U20948 (N_20948,N_16555,N_17121);
and U20949 (N_20949,N_17749,N_16988);
xor U20950 (N_20950,N_19652,N_19074);
xnor U20951 (N_20951,N_17912,N_16843);
nor U20952 (N_20952,N_18347,N_19995);
nor U20953 (N_20953,N_19418,N_16556);
nand U20954 (N_20954,N_19896,N_17875);
and U20955 (N_20955,N_18315,N_19023);
nand U20956 (N_20956,N_19923,N_16105);
nand U20957 (N_20957,N_16317,N_19411);
nor U20958 (N_20958,N_16474,N_19953);
nor U20959 (N_20959,N_15944,N_15550);
nor U20960 (N_20960,N_19576,N_15848);
and U20961 (N_20961,N_16936,N_19933);
and U20962 (N_20962,N_16868,N_18469);
xnor U20963 (N_20963,N_18912,N_15721);
nand U20964 (N_20964,N_19780,N_17136);
or U20965 (N_20965,N_16412,N_18081);
xor U20966 (N_20966,N_17177,N_17420);
or U20967 (N_20967,N_17953,N_16047);
nor U20968 (N_20968,N_15302,N_18221);
nor U20969 (N_20969,N_16093,N_15796);
or U20970 (N_20970,N_18839,N_18951);
or U20971 (N_20971,N_18725,N_19255);
or U20972 (N_20972,N_18404,N_16760);
nand U20973 (N_20973,N_18303,N_16447);
and U20974 (N_20974,N_19375,N_19844);
and U20975 (N_20975,N_18039,N_16783);
and U20976 (N_20976,N_17721,N_15255);
or U20977 (N_20977,N_19694,N_15680);
and U20978 (N_20978,N_19172,N_17339);
or U20979 (N_20979,N_16331,N_18103);
and U20980 (N_20980,N_18019,N_17974);
nor U20981 (N_20981,N_17102,N_19849);
nor U20982 (N_20982,N_17978,N_17175);
and U20983 (N_20983,N_15428,N_19543);
xor U20984 (N_20984,N_19492,N_18486);
nand U20985 (N_20985,N_19107,N_18054);
xnor U20986 (N_20986,N_19986,N_17831);
nor U20987 (N_20987,N_16619,N_15573);
nand U20988 (N_20988,N_17819,N_18918);
and U20989 (N_20989,N_17351,N_17318);
nand U20990 (N_20990,N_19819,N_17051);
nor U20991 (N_20991,N_15922,N_19738);
xnor U20992 (N_20992,N_19717,N_15525);
nor U20993 (N_20993,N_17079,N_17046);
and U20994 (N_20994,N_15281,N_15667);
nand U20995 (N_20995,N_17022,N_15171);
and U20996 (N_20996,N_19698,N_16172);
and U20997 (N_20997,N_17114,N_18536);
nor U20998 (N_20998,N_17816,N_16995);
or U20999 (N_20999,N_18388,N_16643);
xnor U21000 (N_21000,N_19173,N_18661);
or U21001 (N_21001,N_17182,N_18913);
nand U21002 (N_21002,N_17173,N_18197);
nor U21003 (N_21003,N_19013,N_19667);
xor U21004 (N_21004,N_19804,N_16509);
or U21005 (N_21005,N_18678,N_19224);
nand U21006 (N_21006,N_18254,N_18291);
nor U21007 (N_21007,N_19263,N_17818);
nor U21008 (N_21008,N_15836,N_17844);
nor U21009 (N_21009,N_19387,N_19564);
xor U21010 (N_21010,N_19344,N_18175);
nor U21011 (N_21011,N_16669,N_16050);
nor U21012 (N_21012,N_18832,N_18349);
or U21013 (N_21013,N_17920,N_15380);
nor U21014 (N_21014,N_17687,N_18822);
xnor U21015 (N_21015,N_19328,N_15397);
xor U21016 (N_21016,N_19515,N_17347);
and U21017 (N_21017,N_18757,N_15287);
and U21018 (N_21018,N_16662,N_19041);
nor U21019 (N_21019,N_18787,N_16487);
nor U21020 (N_21020,N_16139,N_18037);
nand U21021 (N_21021,N_17662,N_15081);
nor U21022 (N_21022,N_16466,N_18450);
nor U21023 (N_21023,N_16189,N_16710);
and U21024 (N_21024,N_16911,N_17188);
or U21025 (N_21025,N_15670,N_19579);
or U21026 (N_21026,N_15792,N_18020);
xnor U21027 (N_21027,N_15989,N_15072);
nand U21028 (N_21028,N_17343,N_17258);
xor U21029 (N_21029,N_16742,N_18319);
nor U21030 (N_21030,N_19384,N_18170);
xnor U21031 (N_21031,N_15412,N_17755);
xnor U21032 (N_21032,N_15655,N_18484);
nand U21033 (N_21033,N_15366,N_17583);
nand U21034 (N_21034,N_16836,N_18022);
xor U21035 (N_21035,N_17751,N_15916);
nand U21036 (N_21036,N_16148,N_16697);
or U21037 (N_21037,N_16632,N_15414);
xnor U21038 (N_21038,N_19098,N_15535);
nor U21039 (N_21039,N_17269,N_15764);
nor U21040 (N_21040,N_18627,N_17219);
xnor U21041 (N_21041,N_16360,N_17074);
nor U21042 (N_21042,N_19415,N_17647);
nor U21043 (N_21043,N_18861,N_17852);
or U21044 (N_21044,N_18541,N_15674);
nand U21045 (N_21045,N_19049,N_18239);
nand U21046 (N_21046,N_19462,N_16739);
nand U21047 (N_21047,N_19111,N_15957);
nand U21048 (N_21048,N_15164,N_15401);
nand U21049 (N_21049,N_17321,N_17562);
or U21050 (N_21050,N_18119,N_16109);
xor U21051 (N_21051,N_17540,N_17183);
nor U21052 (N_21052,N_19756,N_18290);
nor U21053 (N_21053,N_17683,N_18710);
nor U21054 (N_21054,N_16872,N_19733);
or U21055 (N_21055,N_16801,N_19390);
nand U21056 (N_21056,N_16145,N_18574);
nor U21057 (N_21057,N_17244,N_15045);
or U21058 (N_21058,N_19605,N_19840);
or U21059 (N_21059,N_16106,N_15579);
or U21060 (N_21060,N_18482,N_18726);
or U21061 (N_21061,N_18764,N_15388);
xor U21062 (N_21062,N_16056,N_18731);
or U21063 (N_21063,N_17092,N_18874);
nor U21064 (N_21064,N_16159,N_15837);
nand U21065 (N_21065,N_19909,N_16914);
and U21066 (N_21066,N_19221,N_15595);
or U21067 (N_21067,N_17026,N_16931);
nor U21068 (N_21068,N_19796,N_17055);
or U21069 (N_21069,N_19530,N_15703);
nor U21070 (N_21070,N_19289,N_16757);
nor U21071 (N_21071,N_18313,N_15076);
xnor U21072 (N_21072,N_17729,N_19843);
nor U21073 (N_21073,N_18885,N_17497);
nor U21074 (N_21074,N_18013,N_15234);
nand U21075 (N_21075,N_15715,N_18582);
or U21076 (N_21076,N_17690,N_17133);
nor U21077 (N_21077,N_19830,N_15814);
nor U21078 (N_21078,N_15611,N_17295);
nor U21079 (N_21079,N_17402,N_15948);
or U21080 (N_21080,N_17744,N_19380);
and U21081 (N_21081,N_15546,N_18922);
xnor U21082 (N_21082,N_19488,N_18798);
and U21083 (N_21083,N_15463,N_17389);
xnor U21084 (N_21084,N_19905,N_16074);
or U21085 (N_21085,N_17610,N_17538);
and U21086 (N_21086,N_16725,N_19580);
xnor U21087 (N_21087,N_16395,N_18198);
or U21088 (N_21088,N_18106,N_18179);
nor U21089 (N_21089,N_15389,N_16138);
or U21090 (N_21090,N_17189,N_18557);
nand U21091 (N_21091,N_16009,N_15282);
or U21092 (N_21092,N_19653,N_17670);
nor U21093 (N_21093,N_17296,N_18810);
or U21094 (N_21094,N_15704,N_17812);
nor U21095 (N_21095,N_17376,N_15277);
xnor U21096 (N_21096,N_19011,N_16147);
nand U21097 (N_21097,N_18795,N_19967);
nor U21098 (N_21098,N_15381,N_18376);
nor U21099 (N_21099,N_18762,N_15782);
or U21100 (N_21100,N_15617,N_18357);
or U21101 (N_21101,N_19627,N_17997);
nand U21102 (N_21102,N_19394,N_15628);
and U21103 (N_21103,N_17263,N_17317);
xor U21104 (N_21104,N_16292,N_19510);
nor U21105 (N_21105,N_15028,N_18289);
nor U21106 (N_21106,N_16448,N_15986);
nand U21107 (N_21107,N_17109,N_19854);
xor U21108 (N_21108,N_15700,N_17407);
xor U21109 (N_21109,N_15188,N_16686);
xor U21110 (N_21110,N_15845,N_16152);
or U21111 (N_21111,N_16992,N_17959);
nand U21112 (N_21112,N_16488,N_19744);
nor U21113 (N_21113,N_18800,N_17908);
xnor U21114 (N_21114,N_18113,N_19451);
nand U21115 (N_21115,N_15500,N_18143);
nor U21116 (N_21116,N_15996,N_15304);
or U21117 (N_21117,N_19823,N_17029);
xor U21118 (N_21118,N_16199,N_18027);
and U21119 (N_21119,N_15197,N_17331);
nand U21120 (N_21120,N_19740,N_17064);
xnor U21121 (N_21121,N_17031,N_15707);
xnor U21122 (N_21122,N_17532,N_16848);
nand U21123 (N_21123,N_17302,N_19680);
xor U21124 (N_21124,N_16153,N_19313);
or U21125 (N_21125,N_15771,N_19596);
nand U21126 (N_21126,N_16180,N_15354);
xor U21127 (N_21127,N_18630,N_17413);
or U21128 (N_21128,N_15767,N_18830);
xnor U21129 (N_21129,N_18715,N_17821);
nor U21130 (N_21130,N_16864,N_19631);
and U21131 (N_21131,N_17214,N_17918);
nor U21132 (N_21132,N_17181,N_15858);
nor U21133 (N_21133,N_16284,N_17824);
nand U21134 (N_21134,N_15123,N_19293);
xor U21135 (N_21135,N_19063,N_15436);
nor U21136 (N_21136,N_19553,N_15695);
or U21137 (N_21137,N_17946,N_17528);
xor U21138 (N_21138,N_17168,N_16958);
nor U21139 (N_21139,N_15139,N_18875);
xor U21140 (N_21140,N_15289,N_17070);
nand U21141 (N_21141,N_17907,N_16610);
or U21142 (N_21142,N_17756,N_16091);
and U21143 (N_21143,N_17796,N_15490);
xnor U21144 (N_21144,N_16748,N_16613);
xor U21145 (N_21145,N_15083,N_16846);
and U21146 (N_21146,N_18127,N_15783);
or U21147 (N_21147,N_18865,N_17924);
and U21148 (N_21148,N_18108,N_18168);
nor U21149 (N_21149,N_17712,N_17944);
nor U21150 (N_21150,N_16255,N_18598);
xor U21151 (N_21151,N_18348,N_19056);
or U21152 (N_21152,N_17619,N_16121);
xnor U21153 (N_21153,N_15705,N_19190);
xor U21154 (N_21154,N_17657,N_15785);
xnor U21155 (N_21155,N_19460,N_18809);
nand U21156 (N_21156,N_17104,N_19882);
nor U21157 (N_21157,N_16362,N_17964);
nand U21158 (N_21158,N_15253,N_18668);
nor U21159 (N_21159,N_18872,N_18743);
nand U21160 (N_21160,N_19132,N_18869);
and U21161 (N_21161,N_19138,N_15030);
xnor U21162 (N_21162,N_16223,N_17091);
or U21163 (N_21163,N_17786,N_19571);
nand U21164 (N_21164,N_16283,N_19158);
and U21165 (N_21165,N_19587,N_18589);
xor U21166 (N_21166,N_15753,N_17621);
or U21167 (N_21167,N_17937,N_17426);
or U21168 (N_21168,N_17679,N_16302);
and U21169 (N_21169,N_18863,N_19168);
and U21170 (N_21170,N_19837,N_16000);
nor U21171 (N_21171,N_15914,N_17116);
or U21172 (N_21172,N_16377,N_16078);
xor U21173 (N_21173,N_19641,N_17702);
nand U21174 (N_21174,N_17099,N_15969);
and U21175 (N_21175,N_15291,N_19320);
nand U21176 (N_21176,N_16253,N_19720);
nor U21177 (N_21177,N_19868,N_17698);
and U21178 (N_21178,N_15151,N_16045);
nor U21179 (N_21179,N_16128,N_15806);
xnor U21180 (N_21180,N_17194,N_15337);
or U21181 (N_21181,N_18145,N_18232);
xnor U21182 (N_21182,N_17066,N_16177);
and U21183 (N_21183,N_19757,N_18187);
xor U21184 (N_21184,N_18921,N_16765);
nand U21185 (N_21185,N_17002,N_15978);
and U21186 (N_21186,N_18978,N_15757);
and U21187 (N_21187,N_16468,N_16989);
nor U21188 (N_21188,N_18428,N_18314);
xor U21189 (N_21189,N_15657,N_15776);
nor U21190 (N_21190,N_16671,N_18658);
xnor U21191 (N_21191,N_17477,N_15222);
nor U21192 (N_21192,N_18745,N_18182);
xor U21193 (N_21193,N_18501,N_18284);
and U21194 (N_21194,N_18363,N_15689);
or U21195 (N_21195,N_17444,N_16743);
or U21196 (N_21196,N_19309,N_17094);
or U21197 (N_21197,N_15445,N_19826);
and U21198 (N_21198,N_15822,N_15488);
or U21199 (N_21199,N_18235,N_15485);
xor U21200 (N_21200,N_16615,N_17019);
and U21201 (N_21201,N_16515,N_17980);
and U21202 (N_21202,N_16347,N_15328);
nand U21203 (N_21203,N_17771,N_18105);
or U21204 (N_21204,N_16817,N_19951);
or U21205 (N_21205,N_17706,N_18216);
or U21206 (N_21206,N_18033,N_18160);
nor U21207 (N_21207,N_16690,N_15802);
or U21208 (N_21208,N_18964,N_18928);
xnor U21209 (N_21209,N_16744,N_18231);
nor U21210 (N_21210,N_16861,N_17973);
xor U21211 (N_21211,N_19123,N_18583);
xor U21212 (N_21212,N_15895,N_16103);
nand U21213 (N_21213,N_17629,N_19452);
nand U21214 (N_21214,N_17827,N_17431);
nand U21215 (N_21215,N_17003,N_17487);
nand U21216 (N_21216,N_17828,N_19291);
or U21217 (N_21217,N_18761,N_16544);
xor U21218 (N_21218,N_19998,N_19685);
nand U21219 (N_21219,N_19165,N_19353);
nor U21220 (N_21220,N_16320,N_16393);
xor U21221 (N_21221,N_17994,N_15346);
nand U21222 (N_21222,N_19030,N_19634);
nand U21223 (N_21223,N_15523,N_19736);
and U21224 (N_21224,N_18607,N_17842);
nand U21225 (N_21225,N_18516,N_18648);
or U21226 (N_21226,N_17893,N_18640);
nand U21227 (N_21227,N_19651,N_16269);
or U21228 (N_21228,N_15815,N_15344);
or U21229 (N_21229,N_19931,N_15775);
and U21230 (N_21230,N_15238,N_18532);
or U21231 (N_21231,N_16863,N_15347);
or U21232 (N_21232,N_18265,N_15624);
nand U21233 (N_21233,N_17027,N_18066);
or U21234 (N_21234,N_17668,N_19458);
and U21235 (N_21235,N_19783,N_16841);
xnor U21236 (N_21236,N_16099,N_19533);
nand U21237 (N_21237,N_17577,N_16086);
nor U21238 (N_21238,N_18551,N_16719);
or U21239 (N_21239,N_19062,N_17349);
nor U21240 (N_21240,N_16036,N_18801);
or U21241 (N_21241,N_16371,N_18209);
or U21242 (N_21242,N_19104,N_17509);
xor U21243 (N_21243,N_16939,N_16638);
nand U21244 (N_21244,N_15794,N_16118);
nor U21245 (N_21245,N_16314,N_16098);
xnor U21246 (N_21246,N_19608,N_18547);
nor U21247 (N_21247,N_17227,N_19657);
or U21248 (N_21248,N_18788,N_17255);
and U21249 (N_21249,N_17036,N_15933);
or U21250 (N_21250,N_15245,N_16986);
or U21251 (N_21251,N_17151,N_15516);
nor U21252 (N_21252,N_18359,N_18933);
and U21253 (N_21253,N_18300,N_16574);
and U21254 (N_21254,N_18462,N_17977);
nand U21255 (N_21255,N_19842,N_16251);
or U21256 (N_21256,N_15886,N_15484);
or U21257 (N_21257,N_16599,N_16902);
nand U21258 (N_21258,N_18778,N_18587);
nand U21259 (N_21259,N_17242,N_18112);
nor U21260 (N_21260,N_15158,N_17864);
or U21261 (N_21261,N_15262,N_17545);
xor U21262 (N_21262,N_17623,N_18522);
or U21263 (N_21263,N_16678,N_17333);
or U21264 (N_21264,N_15919,N_17015);
nor U21265 (N_21265,N_18887,N_19055);
nand U21266 (N_21266,N_15630,N_16894);
and U21267 (N_21267,N_18608,N_19932);
nand U21268 (N_21268,N_16416,N_17563);
nand U21269 (N_21269,N_15766,N_19401);
and U21270 (N_21270,N_17330,N_16149);
nand U21271 (N_21271,N_19016,N_19721);
or U21272 (N_21272,N_19859,N_16408);
xor U21273 (N_21273,N_15153,N_15671);
and U21274 (N_21274,N_18820,N_19110);
nand U21275 (N_21275,N_16015,N_17534);
or U21276 (N_21276,N_18181,N_17505);
or U21277 (N_21277,N_19377,N_15772);
xor U21278 (N_21278,N_16244,N_17458);
or U21279 (N_21279,N_16129,N_18860);
and U21280 (N_21280,N_16275,N_16795);
nand U21281 (N_21281,N_18384,N_19645);
xnor U21282 (N_21282,N_18653,N_19768);
xor U21283 (N_21283,N_15725,N_18760);
xor U21284 (N_21284,N_15512,N_16414);
or U21285 (N_21285,N_16272,N_17841);
xor U21286 (N_21286,N_16476,N_19077);
and U21287 (N_21287,N_19695,N_18689);
or U21288 (N_21288,N_15193,N_18371);
nor U21289 (N_21289,N_15450,N_15509);
nor U21290 (N_21290,N_16356,N_16020);
and U21291 (N_21291,N_15421,N_19490);
nor U21292 (N_21292,N_16233,N_17344);
nand U21293 (N_21293,N_19318,N_19471);
and U21294 (N_21294,N_19018,N_16623);
or U21295 (N_21295,N_17262,N_17616);
and U21296 (N_21296,N_18368,N_16847);
nor U21297 (N_21297,N_16891,N_15237);
nand U21298 (N_21298,N_16607,N_18296);
or U21299 (N_21299,N_15761,N_16708);
and U21300 (N_21300,N_19833,N_18990);
nand U21301 (N_21301,N_18048,N_16361);
nor U21302 (N_21302,N_18096,N_15152);
or U21303 (N_21303,N_19793,N_18382);
nand U21304 (N_21304,N_16577,N_16249);
nor U21305 (N_21305,N_15552,N_19502);
or U21306 (N_21306,N_16239,N_18130);
and U21307 (N_21307,N_17293,N_17366);
nand U21308 (N_21308,N_15773,N_15688);
xnor U21309 (N_21309,N_16550,N_17134);
nand U21310 (N_21310,N_19459,N_16510);
or U21311 (N_21311,N_17226,N_19080);
nor U21312 (N_21312,N_18115,N_18492);
nand U21313 (N_21313,N_16062,N_16054);
nand U21314 (N_21314,N_18014,N_18230);
nand U21315 (N_21315,N_15367,N_19060);
and U21316 (N_21316,N_19966,N_17836);
or U21317 (N_21317,N_19043,N_17620);
nor U21318 (N_21318,N_15468,N_17649);
and U21319 (N_21319,N_17839,N_19014);
nand U21320 (N_21320,N_16354,N_15551);
nand U21321 (N_21321,N_18612,N_15521);
nand U21322 (N_21322,N_15053,N_15424);
or U21323 (N_21323,N_18455,N_17260);
nor U21324 (N_21324,N_16905,N_18478);
nor U21325 (N_21325,N_15221,N_16104);
xnor U21326 (N_21326,N_15607,N_17782);
nand U21327 (N_21327,N_17498,N_17862);
xor U21328 (N_21328,N_15616,N_15698);
nor U21329 (N_21329,N_16606,N_18274);
nand U21330 (N_21330,N_17501,N_15423);
nor U21331 (N_21331,N_16972,N_18603);
nor U21332 (N_21332,N_15005,N_17543);
xor U21333 (N_21333,N_18623,N_16422);
nand U21334 (N_21334,N_15687,N_16844);
or U21335 (N_21335,N_16676,N_19274);
and U21336 (N_21336,N_15967,N_19249);
xnor U21337 (N_21337,N_19322,N_18010);
xor U21338 (N_21338,N_18494,N_19260);
or U21339 (N_21339,N_18350,N_18252);
nor U21340 (N_21340,N_15530,N_18855);
nand U21341 (N_21341,N_18717,N_16313);
and U21342 (N_21342,N_19541,N_17728);
nand U21343 (N_21343,N_19417,N_16016);
nand U21344 (N_21344,N_18424,N_17135);
or U21345 (N_21345,N_17949,N_17425);
xnor U21346 (N_21346,N_16082,N_16450);
or U21347 (N_21347,N_17412,N_19012);
xnor U21348 (N_21348,N_17059,N_15871);
or U21349 (N_21349,N_19936,N_18499);
and U21350 (N_21350,N_15393,N_16856);
and U21351 (N_21351,N_16818,N_18916);
and U21352 (N_21352,N_15599,N_16498);
nand U21353 (N_21353,N_19093,N_19739);
or U21354 (N_21354,N_17856,N_17747);
or U21355 (N_21355,N_16287,N_17165);
or U21356 (N_21356,N_15745,N_17062);
nand U21357 (N_21357,N_18827,N_16654);
xnor U21358 (N_21358,N_17991,N_17523);
nand U21359 (N_21359,N_17613,N_19710);
nand U21360 (N_21360,N_15032,N_16746);
nor U21361 (N_21361,N_15280,N_16464);
and U21362 (N_21362,N_19157,N_18836);
nor U21363 (N_21363,N_18698,N_19938);
and U21364 (N_21364,N_18649,N_18797);
nor U21365 (N_21365,N_18180,N_15840);
or U21366 (N_21366,N_18217,N_17727);
xnor U21367 (N_21367,N_17587,N_15834);
nand U21368 (N_21368,N_16651,N_15522);
and U21369 (N_21369,N_17829,N_19456);
nand U21370 (N_21370,N_16573,N_18817);
or U21371 (N_21371,N_18586,N_19122);
or U21372 (N_21372,N_15910,N_15196);
or U21373 (N_21373,N_16396,N_16539);
and U21374 (N_21374,N_17965,N_19114);
nor U21375 (N_21375,N_16512,N_18040);
or U21376 (N_21376,N_17680,N_18581);
nor U21377 (N_21377,N_19565,N_19646);
xor U21378 (N_21378,N_16463,N_19617);
nand U21379 (N_21379,N_17150,N_18338);
or U21380 (N_21380,N_18467,N_17948);
and U21381 (N_21381,N_18271,N_15664);
nand U21382 (N_21382,N_15718,N_16927);
nand U21383 (N_21383,N_17143,N_18576);
and U21384 (N_21384,N_17447,N_19930);
or U21385 (N_21385,N_15629,N_19674);
xnor U21386 (N_21386,N_15605,N_17316);
nand U21387 (N_21387,N_18204,N_19774);
and U21388 (N_21388,N_17894,N_15874);
or U21389 (N_21389,N_18268,N_19487);
nor U21390 (N_21390,N_16917,N_15864);
nor U21391 (N_21391,N_19185,N_19562);
xnor U21392 (N_21392,N_18396,N_17834);
or U21393 (N_21393,N_16991,N_17254);
and U21394 (N_21394,N_18708,N_17537);
nor U21395 (N_21395,N_16333,N_16981);
or U21396 (N_21396,N_19256,N_19434);
nand U21397 (N_21397,N_17076,N_19250);
xor U21398 (N_21398,N_18104,N_17773);
nand U21399 (N_21399,N_16729,N_15603);
or U21400 (N_21400,N_17247,N_15384);
nor U21401 (N_21401,N_18421,N_19481);
or U21402 (N_21402,N_17167,N_16754);
nand U21403 (N_21403,N_17569,N_16504);
and U21404 (N_21404,N_16944,N_16775);
and U21405 (N_21405,N_15722,N_18943);
nor U21406 (N_21406,N_18895,N_16731);
xnor U21407 (N_21407,N_16174,N_17354);
nand U21408 (N_21408,N_15150,N_17581);
nand U21409 (N_21409,N_15810,N_16915);
or U21410 (N_21410,N_15042,N_19602);
or U21411 (N_21411,N_16024,N_17672);
xnor U21412 (N_21412,N_18791,N_18227);
and U21413 (N_21413,N_19875,N_19301);
xor U21414 (N_21414,N_15351,N_18802);
xnor U21415 (N_21415,N_18521,N_16955);
nand U21416 (N_21416,N_15471,N_16170);
xor U21417 (N_21417,N_18471,N_18684);
xnor U21418 (N_21418,N_19534,N_15860);
xnor U21419 (N_21419,N_15129,N_18529);
nor U21420 (N_21420,N_17887,N_19876);
xnor U21421 (N_21421,N_15457,N_15883);
xor U21422 (N_21422,N_19947,N_15678);
nand U21423 (N_21423,N_18846,N_15360);
nor U21424 (N_21424,N_15206,N_17640);
xnor U21425 (N_21425,N_19575,N_17032);
nand U21426 (N_21426,N_18392,N_17590);
xnor U21427 (N_21427,N_17232,N_18136);
or U21428 (N_21428,N_19468,N_17164);
nand U21429 (N_21429,N_18988,N_19210);
xor U21430 (N_21430,N_18405,N_15538);
and U21431 (N_21431,N_17090,N_15031);
or U21432 (N_21432,N_16113,N_16008);
or U21433 (N_21433,N_16477,N_17900);
xnor U21434 (N_21434,N_18555,N_17013);
or U21435 (N_21435,N_19647,N_17896);
nand U21436 (N_21436,N_16875,N_15953);
nand U21437 (N_21437,N_18702,N_15602);
xnor U21438 (N_21438,N_19421,N_16167);
and U21439 (N_21439,N_19689,N_19507);
or U21440 (N_21440,N_18332,N_16225);
nor U21441 (N_21441,N_18744,N_19095);
or U21442 (N_21442,N_17740,N_16857);
or U21443 (N_21443,N_17724,N_17052);
and U21444 (N_21444,N_15755,N_15395);
nor U21445 (N_21445,N_17938,N_17837);
xnor U21446 (N_21446,N_16455,N_15964);
and U21447 (N_21447,N_17660,N_19941);
and U21448 (N_21448,N_18553,N_17776);
and U21449 (N_21449,N_17909,N_19622);
or U21450 (N_21450,N_18055,N_16374);
nor U21451 (N_21451,N_18413,N_17278);
and U21452 (N_21452,N_16897,N_19942);
xnor U21453 (N_21453,N_15178,N_19665);
and U21454 (N_21454,N_18385,N_17313);
xor U21455 (N_21455,N_18967,N_17709);
nor U21456 (N_21456,N_19636,N_16837);
nor U21457 (N_21457,N_15165,N_19252);
xor U21458 (N_21458,N_17777,N_17840);
and U21459 (N_21459,N_18975,N_15658);
and U21460 (N_21460,N_19010,N_16089);
nand U21461 (N_21461,N_15821,N_19266);
and U21462 (N_21462,N_16704,N_16365);
or U21463 (N_21463,N_18042,N_16591);
nor U21464 (N_21464,N_19713,N_18892);
nand U21465 (N_21465,N_19991,N_19790);
nor U21466 (N_21466,N_18540,N_16096);
nor U21467 (N_21467,N_16771,N_17710);
xnor U21468 (N_21468,N_19620,N_18423);
and U21469 (N_21469,N_16572,N_19121);
and U21470 (N_21470,N_18154,N_15403);
or U21471 (N_21471,N_15207,N_18859);
and U21472 (N_21472,N_19560,N_15070);
xor U21473 (N_21473,N_16608,N_19079);
and U21474 (N_21474,N_19241,N_17508);
nand U21475 (N_21475,N_16141,N_18805);
or U21476 (N_21476,N_17144,N_17883);
xor U21477 (N_21477,N_19358,N_19146);
xor U21478 (N_21478,N_18883,N_16079);
nor U21479 (N_21479,N_19245,N_16021);
xnor U21480 (N_21480,N_18293,N_16524);
xor U21481 (N_21481,N_18383,N_17695);
xor U21482 (N_21482,N_19883,N_19153);
nor U21483 (N_21483,N_19509,N_19886);
nor U21484 (N_21484,N_18056,N_19926);
and U21485 (N_21485,N_17152,N_18166);
nor U21486 (N_21486,N_16185,N_19778);
nor U21487 (N_21487,N_18447,N_15392);
nor U21488 (N_21488,N_16723,N_18330);
and U21489 (N_21489,N_15118,N_19948);
or U21490 (N_21490,N_17626,N_17752);
nand U21491 (N_21491,N_19222,N_16924);
and U21492 (N_21492,N_19498,N_15896);
or U21493 (N_21493,N_19957,N_15988);
nor U21494 (N_21494,N_19974,N_16247);
nand U21495 (N_21495,N_16870,N_17665);
and U21496 (N_21496,N_17510,N_15211);
and U21497 (N_21497,N_19528,N_19265);
xor U21498 (N_21498,N_19900,N_19615);
and U21499 (N_21499,N_16896,N_15456);
nand U21500 (N_21500,N_16943,N_16348);
nor U21501 (N_21501,N_18944,N_19508);
or U21502 (N_21502,N_19828,N_18621);
nor U21503 (N_21503,N_15365,N_19984);
nand U21504 (N_21504,N_17772,N_17822);
xnor U21505 (N_21505,N_16620,N_16042);
nor U21506 (N_21506,N_15973,N_16234);
xnor U21507 (N_21507,N_16779,N_18680);
xnor U21508 (N_21508,N_16680,N_16114);
and U21509 (N_21509,N_19334,N_19426);
xor U21510 (N_21510,N_17606,N_19853);
nor U21511 (N_21511,N_18568,N_16405);
or U21512 (N_21512,N_15588,N_16262);
nor U21513 (N_21513,N_18953,N_15069);
nand U21514 (N_21514,N_15909,N_17584);
nor U21515 (N_21515,N_16973,N_18107);
nor U21516 (N_21516,N_15555,N_17987);
nand U21517 (N_21517,N_17113,N_18906);
and U21518 (N_21518,N_18141,N_17863);
xor U21519 (N_21519,N_19088,N_17742);
nor U21520 (N_21520,N_15769,N_17257);
xor U21521 (N_21521,N_17364,N_15318);
or U21522 (N_21522,N_18660,N_15749);
nand U21523 (N_21523,N_15526,N_16004);
nand U21524 (N_21524,N_17442,N_17689);
and U21525 (N_21525,N_15590,N_18089);
nand U21526 (N_21526,N_18460,N_19465);
or U21527 (N_21527,N_19929,N_18991);
nand U21528 (N_21528,N_17359,N_16640);
and U21529 (N_21529,N_15187,N_18090);
nand U21530 (N_21530,N_19339,N_18911);
nor U21531 (N_21531,N_15326,N_19386);
nor U21532 (N_21532,N_18135,N_18002);
or U21533 (N_21533,N_16430,N_15054);
xnor U21534 (N_21534,N_19202,N_18212);
nor U21535 (N_21535,N_16075,N_17068);
and U21536 (N_21536,N_16647,N_19705);
nor U21537 (N_21537,N_18654,N_17309);
nand U21538 (N_21538,N_15663,N_15774);
nand U21539 (N_21539,N_19873,N_17789);
nand U21540 (N_21540,N_19503,N_19117);
or U21541 (N_21541,N_18358,N_18969);
xor U21542 (N_21542,N_17549,N_16027);
nor U21543 (N_21543,N_16286,N_16900);
xor U21544 (N_21544,N_18564,N_19161);
nor U21545 (N_21545,N_16081,N_16134);
nor U21546 (N_21546,N_18351,N_15040);
or U21547 (N_21547,N_17390,N_15133);
xor U21548 (N_21548,N_16595,N_18344);
nor U21549 (N_21549,N_17482,N_15434);
and U21550 (N_21550,N_18263,N_18989);
nand U21551 (N_21551,N_16315,N_16490);
xor U21552 (N_21552,N_16949,N_19539);
nand U21553 (N_21553,N_16881,N_16459);
nand U21554 (N_21554,N_18523,N_19277);
and U21555 (N_21555,N_19945,N_17625);
nand U21556 (N_21556,N_18114,N_19513);
nand U21557 (N_21557,N_17692,N_18442);
or U21558 (N_21558,N_17005,N_18562);
nand U21559 (N_21559,N_19884,N_15746);
nor U21560 (N_21560,N_16922,N_17272);
or U21561 (N_21561,N_18047,N_19592);
or U21562 (N_21562,N_15894,N_16559);
xnor U21563 (N_21563,N_18980,N_19531);
nor U21564 (N_21564,N_17298,N_18452);
and U21565 (N_21565,N_19980,N_18901);
xnor U21566 (N_21566,N_18253,N_19102);
or U21567 (N_21567,N_19003,N_18976);
and U21568 (N_21568,N_16770,N_16561);
or U21569 (N_21569,N_19648,N_18470);
nor U21570 (N_21570,N_19343,N_17100);
xnor U21571 (N_21571,N_19447,N_16532);
and U21572 (N_21572,N_17599,N_19366);
nand U21573 (N_21573,N_18604,N_15501);
nor U21574 (N_21574,N_19787,N_19081);
nor U21575 (N_21575,N_19555,N_19282);
nor U21576 (N_21576,N_16592,N_16446);
nand U21577 (N_21577,N_15060,N_19977);
nor U21578 (N_21578,N_19204,N_17781);
nor U21579 (N_21579,N_17225,N_17934);
xor U21580 (N_21580,N_19497,N_19504);
nand U21581 (N_21581,N_17041,N_15645);
or U21582 (N_21582,N_19895,N_17546);
or U21583 (N_21583,N_15491,N_17441);
xnor U21584 (N_21584,N_17223,N_17042);
xor U21585 (N_21585,N_17229,N_17030);
nand U21586 (N_21586,N_17147,N_16475);
and U21587 (N_21587,N_16285,N_16469);
and U21588 (N_21588,N_17455,N_15882);
or U21589 (N_21589,N_17460,N_19085);
or U21590 (N_21590,N_15248,N_15903);
or U21591 (N_21591,N_17040,N_18340);
and U21592 (N_21592,N_19175,N_18606);
nand U21593 (N_21593,N_17459,N_18061);
and U21594 (N_21594,N_18298,N_18500);
and U21595 (N_21595,N_16799,N_16705);
and U21596 (N_21596,N_16794,N_16736);
and U21597 (N_21597,N_16547,N_17081);
nand U21598 (N_21598,N_18152,N_15668);
xor U21599 (N_21599,N_19940,N_19762);
and U21600 (N_21600,N_17792,N_17809);
or U21601 (N_21601,N_16195,N_18210);
and U21602 (N_21602,N_18639,N_18219);
nor U21603 (N_21603,N_17370,N_19594);
or U21604 (N_21604,N_15991,N_15013);
xor U21605 (N_21605,N_19477,N_15256);
xor U21606 (N_21606,N_18697,N_17715);
nand U21607 (N_21607,N_18342,N_19735);
xor U21608 (N_21608,N_18367,N_16044);
nor U21609 (N_21609,N_17084,N_17598);
and U21610 (N_21610,N_18095,N_18882);
xor U21611 (N_21611,N_17800,N_18824);
and U21612 (N_21612,N_18646,N_15292);
nand U21613 (N_21613,N_18009,N_19676);
or U21614 (N_21614,N_17157,N_15740);
nand U21615 (N_21615,N_15997,N_18693);
or U21616 (N_21616,N_18984,N_16427);
and U21617 (N_21617,N_19065,N_15528);
nand U21618 (N_21618,N_18509,N_16014);
nor U21619 (N_21619,N_18850,N_15018);
or U21620 (N_21620,N_16675,N_16829);
xor U21621 (N_21621,N_15217,N_19211);
xnor U21622 (N_21622,N_19797,N_18030);
nand U21623 (N_21623,N_18394,N_18556);
nor U21624 (N_21624,N_18786,N_18673);
and U21625 (N_21625,N_15359,N_15147);
and U21626 (N_21626,N_17593,N_15474);
or U21627 (N_21627,N_17400,N_17582);
nand U21628 (N_21628,N_18243,N_16382);
xor U21629 (N_21629,N_17868,N_17605);
nor U21630 (N_21630,N_17484,N_15564);
nand U21631 (N_21631,N_18044,N_16528);
or U21632 (N_21632,N_17717,N_19639);
and U21633 (N_21633,N_19679,N_19281);
and U21634 (N_21634,N_17960,N_15557);
nor U21635 (N_21635,N_16589,N_16321);
and U21636 (N_21636,N_17327,N_15108);
or U21637 (N_21637,N_17873,N_17161);
nor U21638 (N_21638,N_19333,N_17801);
nand U21639 (N_21639,N_18890,N_17947);
nor U21640 (N_21640,N_19207,N_17632);
nor U21641 (N_21641,N_15092,N_18753);
nand U21642 (N_21642,N_17905,N_16001);
nor U21643 (N_21643,N_16087,N_17559);
or U21644 (N_21644,N_17110,N_15540);
nor U21645 (N_21645,N_19577,N_16305);
xnor U21646 (N_21646,N_18707,N_19147);
nand U21647 (N_21647,N_15502,N_18932);
nand U21648 (N_21648,N_15006,N_18566);
nand U21649 (N_21649,N_15677,N_15114);
and U21650 (N_21650,N_18409,N_19108);
nor U21651 (N_21651,N_17416,N_15743);
and U21652 (N_21652,N_15593,N_16219);
xor U21653 (N_21653,N_17462,N_18041);
nand U21654 (N_21654,N_19409,N_17511);
nand U21655 (N_21655,N_18664,N_19959);
nand U21656 (N_21656,N_19381,N_15363);
xnor U21657 (N_21657,N_19237,N_15155);
and U21658 (N_21658,N_17446,N_19053);
xor U21659 (N_21659,N_19214,N_16575);
nand U21660 (N_21660,N_19906,N_17798);
xor U21661 (N_21661,N_16059,N_19294);
nand U21662 (N_21662,N_19523,N_16164);
nand U21663 (N_21663,N_16057,N_19613);
xor U21664 (N_21664,N_15100,N_15823);
xnor U21665 (N_21665,N_17676,N_19975);
nand U21666 (N_21666,N_15186,N_15923);
nand U21667 (N_21667,N_15770,N_15439);
xnor U21668 (N_21668,N_19278,N_18750);
or U21669 (N_21669,N_18754,N_17638);
nand U21670 (N_21670,N_15465,N_16363);
and U21671 (N_21671,N_19824,N_18923);
xnor U21672 (N_21672,N_17832,N_19435);
and U21673 (N_21673,N_18898,N_16406);
or U21674 (N_21674,N_15077,N_17014);
or U21675 (N_21675,N_18251,N_18137);
nor U21676 (N_21676,N_18417,N_18510);
xor U21677 (N_21677,N_16650,N_17118);
nor U21678 (N_21678,N_19593,N_15961);
nor U21679 (N_21679,N_16542,N_19479);
nand U21680 (N_21680,N_16445,N_15161);
xnor U21681 (N_21681,N_16404,N_16115);
or U21682 (N_21682,N_18739,N_17639);
xor U21683 (N_21683,N_19730,N_18811);
or U21684 (N_21684,N_18377,N_16130);
and U21685 (N_21685,N_16929,N_17642);
and U21686 (N_21686,N_18826,N_15430);
or U21687 (N_21687,N_16135,N_15174);
or U21688 (N_21688,N_16626,N_15998);
nor U21689 (N_21689,N_16326,N_19425);
nor U21690 (N_21690,N_15839,N_17589);
nand U21691 (N_21691,N_18399,N_17982);
and U21692 (N_21692,N_15437,N_19033);
nand U21693 (N_21693,N_17643,N_17571);
xnor U21694 (N_21694,N_17054,N_15733);
nand U21695 (N_21695,N_16786,N_17697);
or U21696 (N_21696,N_18973,N_19273);
nor U21697 (N_21697,N_15558,N_18074);
or U21698 (N_21698,N_18584,N_17129);
nand U21699 (N_21699,N_17768,N_17170);
xnor U21700 (N_21700,N_16041,N_16913);
and U21701 (N_21701,N_15742,N_15422);
or U21702 (N_21702,N_16518,N_15037);
xor U21703 (N_21703,N_19346,N_16037);
and U21704 (N_21704,N_16171,N_19609);
xnor U21705 (N_21705,N_19496,N_16565);
or U21706 (N_21706,N_19414,N_17878);
xnor U21707 (N_21707,N_15162,N_15800);
nor U21708 (N_21708,N_15167,N_17307);
or U21709 (N_21709,N_19614,N_15228);
or U21710 (N_21710,N_16946,N_19540);
nand U21711 (N_21711,N_18260,N_19919);
nand U21712 (N_21712,N_16311,N_16436);
nand U21713 (N_21713,N_17726,N_15288);
nor U21714 (N_21714,N_18812,N_18093);
nor U21715 (N_21715,N_15932,N_18436);
and U21716 (N_21716,N_16035,N_16979);
nand U21717 (N_21717,N_16585,N_17004);
nand U21718 (N_21718,N_16646,N_19879);
nand U21719 (N_21719,N_19007,N_16598);
xor U21720 (N_21720,N_19969,N_15777);
and U21721 (N_21721,N_16111,N_19624);
nand U21722 (N_21722,N_15880,N_16790);
nor U21723 (N_21723,N_17238,N_19874);
or U21724 (N_21724,N_16205,N_16835);
or U21725 (N_21725,N_17838,N_18853);
nor U21726 (N_21726,N_15296,N_16833);
xor U21727 (N_21727,N_19934,N_15637);
nand U21728 (N_21728,N_17585,N_18176);
or U21729 (N_21729,N_19292,N_19954);
nand U21730 (N_21730,N_16983,N_15229);
and U21731 (N_21731,N_17705,N_16040);
and U21732 (N_21732,N_17956,N_16484);
xor U21733 (N_21733,N_18410,N_16013);
nor U21734 (N_21734,N_19983,N_17361);
nand U21735 (N_21735,N_17334,N_18398);
and U21736 (N_21736,N_19889,N_19588);
nor U21737 (N_21737,N_15038,N_19357);
or U21738 (N_21738,N_18379,N_19136);
xnor U21739 (N_21739,N_19638,N_19870);
nand U21740 (N_21740,N_16241,N_16548);
nor U21741 (N_21741,N_15257,N_15841);
nor U21742 (N_21742,N_15475,N_17163);
nand U21743 (N_21743,N_18507,N_19669);
and U21744 (N_21744,N_18910,N_15790);
or U21745 (N_21745,N_18402,N_18393);
nor U21746 (N_21746,N_19538,N_18326);
or U21747 (N_21747,N_15065,N_17930);
nor U21748 (N_21748,N_16976,N_19351);
nand U21749 (N_21749,N_15285,N_16948);
nor U21750 (N_21750,N_16252,N_15951);
or U21751 (N_21751,N_17069,N_17409);
nand U21752 (N_21752,N_19525,N_17371);
xor U21753 (N_21753,N_15954,N_15925);
or U21754 (N_21754,N_16336,N_16227);
and U21755 (N_21755,N_19348,N_19916);
xnor U21756 (N_21756,N_15913,N_19788);
and U21757 (N_21757,N_17833,N_15911);
xnor U21758 (N_21758,N_17745,N_15741);
xor U21759 (N_21759,N_18960,N_16095);
and U21760 (N_21760,N_16956,N_15872);
xnor U21761 (N_21761,N_17989,N_17850);
nand U21762 (N_21762,N_18082,N_16261);
xnor U21763 (N_21763,N_19037,N_15541);
and U21764 (N_21764,N_16957,N_18920);
and U21765 (N_21765,N_16514,N_15893);
or U21766 (N_21766,N_17202,N_16644);
nand U21767 (N_21767,N_17075,N_17033);
and U21768 (N_21768,N_15654,N_17943);
or U21769 (N_21769,N_17748,N_19036);
xor U21770 (N_21770,N_15888,N_18004);
and U21771 (N_21771,N_15029,N_15041);
and U21772 (N_21772,N_17378,N_19196);
and U21773 (N_21773,N_17060,N_15192);
xor U21774 (N_21774,N_15547,N_17088);
xor U21775 (N_21775,N_15803,N_19996);
or U21776 (N_21776,N_15728,N_19374);
or U21777 (N_21777,N_16832,N_15442);
nor U21778 (N_21778,N_17799,N_15048);
xnor U21779 (N_21779,N_18005,N_17685);
nand U21780 (N_21780,N_19251,N_16264);
nand U21781 (N_21781,N_19558,N_16941);
xor U21782 (N_21782,N_19761,N_15844);
xor U21783 (N_21783,N_19659,N_17398);
or U21784 (N_21784,N_15453,N_16052);
nand U21785 (N_21785,N_18880,N_18662);
and U21786 (N_21786,N_16274,N_15270);
and U21787 (N_21787,N_17172,N_19026);
and U21788 (N_21788,N_17048,N_19899);
or U21789 (N_21789,N_19307,N_19349);
nand U21790 (N_21790,N_17693,N_18962);
xnor U21791 (N_21791,N_17825,N_18273);
nand U21792 (N_21792,N_16019,N_16254);
and U21793 (N_21793,N_16155,N_15125);
and U21794 (N_21794,N_16410,N_19370);
nor U21795 (N_21795,N_19180,N_17279);
nand U21796 (N_21796,N_16586,N_17266);
nand U21797 (N_21797,N_18072,N_18572);
or U21798 (N_21798,N_16017,N_17784);
nand U21799 (N_21799,N_15685,N_18831);
xnor U21800 (N_21800,N_18346,N_15730);
xnor U21801 (N_21801,N_15473,N_17362);
or U21802 (N_21802,N_15181,N_17418);
nor U21803 (N_21803,N_15443,N_19067);
xor U21804 (N_21804,N_16462,N_19618);
or U21805 (N_21805,N_17971,N_15051);
nor U21806 (N_21806,N_19050,N_15920);
or U21807 (N_21807,N_15987,N_15177);
nand U21808 (N_21808,N_19922,N_18063);
nand U21809 (N_21809,N_19257,N_16308);
nand U21810 (N_21810,N_19288,N_16970);
xor U21811 (N_21811,N_18257,N_17759);
nand U21812 (N_21812,N_15498,N_17552);
and U21813 (N_21813,N_16140,N_17650);
and U21814 (N_21814,N_17627,N_18948);
nand U21815 (N_21815,N_19379,N_15710);
nor U21816 (N_21816,N_15084,N_15140);
nand U21817 (N_21817,N_17452,N_16782);
nand U21818 (N_21818,N_16730,N_16674);
and U21819 (N_21819,N_17312,N_16478);
xnor U21820 (N_21820,N_18884,N_17870);
nand U21821 (N_21821,N_16756,N_17882);
nor U21822 (N_21822,N_19064,N_17020);
nand U21823 (N_21823,N_17858,N_17283);
nand U21824 (N_21824,N_18234,N_16046);
xor U21825 (N_21825,N_19621,N_16893);
nor U21826 (N_21826,N_16203,N_17903);
and U21827 (N_21827,N_16055,N_18537);
or U21828 (N_21828,N_19422,N_16499);
nand U21829 (N_21829,N_17659,N_17913);
and U21830 (N_21830,N_17617,N_16063);
xnor U21831 (N_21831,N_15708,N_18854);
and U21832 (N_21832,N_18155,N_16534);
and U21833 (N_21833,N_17761,N_19547);
and U21834 (N_21834,N_16318,N_19848);
and U21835 (N_21835,N_15319,N_15702);
and U21836 (N_21836,N_17179,N_19805);
and U21837 (N_21837,N_16969,N_16181);
xor U21838 (N_21838,N_18998,N_18285);
nor U21839 (N_21839,N_19082,N_19167);
or U21840 (N_21840,N_18248,N_15875);
or U21841 (N_21841,N_19670,N_17733);
xor U21842 (N_21842,N_17213,N_15213);
and U21843 (N_21843,N_19427,N_17845);
xnor U21844 (N_21844,N_18165,N_19270);
nand U21845 (N_21845,N_17236,N_15890);
and U21846 (N_21846,N_18185,N_19360);
nand U21847 (N_21847,N_15062,N_16653);
nand U21848 (N_21848,N_15596,N_15750);
xnor U21849 (N_21849,N_19557,N_15854);
and U21850 (N_21850,N_15107,N_19076);
nand U21851 (N_21851,N_19356,N_16511);
and U21852 (N_21852,N_19742,N_19765);
or U21853 (N_21853,N_15198,N_19546);
nand U21854 (N_21854,N_15614,N_18538);
and U21855 (N_21855,N_17010,N_18567);
xor U21856 (N_21856,N_18131,N_18088);
and U21857 (N_21857,N_16774,N_19388);
xnor U21858 (N_21858,N_19649,N_17885);
xor U21859 (N_21859,N_18247,N_18373);
xor U21860 (N_21860,N_16901,N_16858);
or U21861 (N_21861,N_17597,N_19429);
nand U21862 (N_21862,N_18189,N_16479);
nand U21863 (N_21863,N_15094,N_15768);
nand U21864 (N_21864,N_19369,N_19514);
nand U21865 (N_21865,N_18891,N_16657);
or U21866 (N_21866,N_16407,N_16940);
nor U21867 (N_21867,N_16665,N_18121);
nor U21868 (N_21868,N_16999,N_19807);
nor U21869 (N_21869,N_19825,N_15706);
nor U21870 (N_21870,N_17387,N_17940);
nor U21871 (N_21871,N_15348,N_18202);
nor U21872 (N_21872,N_15331,N_15093);
nor U21873 (N_21873,N_16297,N_18445);
xnor U21874 (N_21874,N_17008,N_17341);
and U21875 (N_21875,N_19943,N_16867);
xnor U21876 (N_21876,N_19232,N_15975);
or U21877 (N_21877,N_18626,N_19516);
and U21878 (N_21878,N_19960,N_15908);
nand U21879 (N_21879,N_16605,N_17290);
nor U21880 (N_21880,N_17007,N_18907);
nand U21881 (N_21881,N_18194,N_17544);
or U21882 (N_21882,N_16034,N_18390);
xor U21883 (N_21883,N_16208,N_18305);
xor U21884 (N_21884,N_18461,N_16418);
nor U21885 (N_21885,N_16437,N_16496);
xor U21886 (N_21886,N_18387,N_18438);
and U21887 (N_21887,N_15027,N_18677);
nor U21888 (N_21888,N_15168,N_18755);
nor U21889 (N_21889,N_16202,N_17922);
or U21890 (N_21890,N_18669,N_18851);
or U21891 (N_21891,N_17615,N_16465);
and U21892 (N_21892,N_18847,N_19801);
and U21893 (N_21893,N_16364,N_16966);
nor U21894 (N_21894,N_18790,N_16290);
xor U21895 (N_21895,N_18592,N_16117);
nor U21896 (N_21896,N_16692,N_16721);
nor U21897 (N_21897,N_17350,N_17860);
and U21898 (N_21898,N_15517,N_16529);
and U21899 (N_21899,N_18083,N_18618);
nor U21900 (N_21900,N_19229,N_16814);
xor U21901 (N_21901,N_19832,N_16876);
nand U21902 (N_21902,N_17682,N_16792);
or U21903 (N_21903,N_15931,N_19763);
and U21904 (N_21904,N_15209,N_17445);
nand U21905 (N_21905,N_16752,N_19755);
nand U21906 (N_21906,N_17968,N_19179);
and U21907 (N_21907,N_17421,N_18866);
xor U21908 (N_21908,N_17461,N_15117);
and U21909 (N_21909,N_15226,N_15149);
or U21910 (N_21910,N_19781,N_15195);
or U21911 (N_21911,N_16381,N_19325);
nand U21912 (N_21912,N_16928,N_18545);
nor U21913 (N_21913,N_16240,N_16923);
nor U21914 (N_21914,N_15712,N_18837);
nand U21915 (N_21915,N_15431,N_15608);
nor U21916 (N_21916,N_15956,N_19718);
or U21917 (N_21917,N_19723,N_18718);
and U21918 (N_21918,N_16083,N_19408);
xor U21919 (N_21919,N_18117,N_19367);
and U21920 (N_21920,N_17386,N_16553);
xnor U21921 (N_21921,N_15399,N_18925);
xnor U21922 (N_21922,N_17928,N_18966);
nor U21923 (N_21923,N_15333,N_18073);
and U21924 (N_21924,N_18740,N_15014);
nand U21925 (N_21925,N_15519,N_16403);
or U21926 (N_21926,N_19457,N_18637);
or U21927 (N_21927,N_16355,N_19897);
xor U21928 (N_21928,N_15970,N_17472);
or U21929 (N_21929,N_19001,N_18345);
nand U21930 (N_21930,N_16603,N_17588);
or U21931 (N_21931,N_18080,N_18867);
nor U21932 (N_21932,N_18018,N_17417);
xor U21933 (N_21933,N_19925,N_17848);
nor U21934 (N_21934,N_16601,N_16798);
and U21935 (N_21935,N_17854,N_18776);
or U21936 (N_21936,N_18525,N_15972);
nor U21937 (N_21937,N_19186,N_15560);
xor U21938 (N_21938,N_17902,N_19820);
and U21939 (N_21939,N_16232,N_16343);
nand U21940 (N_21940,N_18324,N_16196);
nor U21941 (N_21941,N_19235,N_19133);
and U21942 (N_21942,N_15227,N_17145);
nor U21943 (N_21943,N_16342,N_17282);
or U21944 (N_21944,N_19327,N_15148);
xor U21945 (N_21945,N_15293,N_16971);
and U21946 (N_21946,N_18163,N_16344);
nor U21947 (N_21947,N_16161,N_15246);
nor U21948 (N_21948,N_16703,N_18695);
or U21949 (N_21949,N_15297,N_16260);
or U21950 (N_21950,N_19156,N_16387);
or U21951 (N_21951,N_15398,N_17519);
or U21952 (N_21952,N_16383,N_18012);
xor U21953 (N_21953,N_16637,N_18372);
nor U21954 (N_21954,N_17681,N_18474);
xnor U21955 (N_21955,N_17380,N_17089);
or U21956 (N_21956,N_19177,N_19734);
xor U21957 (N_21957,N_15927,N_15341);
xnor U21958 (N_21958,N_19352,N_17467);
and U21959 (N_21959,N_15321,N_15276);
nand U21960 (N_21960,N_16048,N_16324);
and U21961 (N_21961,N_16358,N_16787);
xor U21962 (N_21962,N_19625,N_15146);
nor U21963 (N_21963,N_19025,N_15892);
nor U21964 (N_21964,N_18667,N_19869);
and U21965 (N_21965,N_15448,N_15180);
or U21966 (N_21966,N_18682,N_15452);
or U21967 (N_21967,N_15653,N_15921);
nor U21968 (N_21968,N_17415,N_19802);
nand U21969 (N_21969,N_16806,N_15343);
nand U21970 (N_21970,N_16618,N_19858);
nand U21971 (N_21971,N_17496,N_18193);
xnor U21972 (N_21972,N_19835,N_19463);
and U21973 (N_21973,N_16357,N_16351);
nor U21974 (N_21974,N_19008,N_18036);
nor U21975 (N_21975,N_17294,N_19267);
and U21976 (N_21976,N_19545,N_18024);
nor U21977 (N_21977,N_17804,N_15218);
nor U21978 (N_21978,N_18766,N_15009);
xor U21979 (N_21979,N_18594,N_18767);
nand U21980 (N_21980,N_19192,N_18225);
nand U21981 (N_21981,N_17797,N_15681);
nand U21982 (N_21982,N_15233,N_17146);
xor U21983 (N_21983,N_15482,N_19779);
xnor U21984 (N_21984,N_18466,N_15537);
nor U21985 (N_21985,N_16831,N_16865);
and U21986 (N_21986,N_15271,N_19162);
xor U21987 (N_21987,N_17456,N_18318);
nor U21988 (N_21988,N_15665,N_17932);
nand U21989 (N_21989,N_18068,N_16184);
xnor U21990 (N_21990,N_17077,N_16526);
and U21991 (N_21991,N_15278,N_18256);
xnor U21992 (N_21992,N_17123,N_16126);
and U21993 (N_21993,N_17155,N_16221);
or U21994 (N_21994,N_18059,N_17494);
or U21995 (N_21995,N_18735,N_16519);
and U21996 (N_21996,N_17757,N_18659);
or U21997 (N_21997,N_19310,N_17866);
and U21998 (N_21998,N_15169,N_16551);
nor U21999 (N_21999,N_19058,N_19312);
or U22000 (N_22000,N_16758,N_18843);
nand U22001 (N_22001,N_18624,N_16166);
and U22002 (N_22002,N_15481,N_15325);
and U22003 (N_22003,N_19753,N_15669);
xor U22004 (N_22004,N_15303,N_19700);
and U22005 (N_22005,N_19124,N_18829);
and U22006 (N_22006,N_15549,N_15477);
and U22007 (N_22007,N_17580,N_15036);
or U22008 (N_22008,N_15784,N_15918);
nand U22009 (N_22009,N_19677,N_15258);
xnor U22010 (N_22010,N_17788,N_18703);
nand U22011 (N_22011,N_19831,N_19935);
nor U22012 (N_22012,N_17811,N_15527);
or U22013 (N_22013,N_16885,N_16435);
nor U22014 (N_22014,N_16325,N_15061);
nand U22015 (N_22015,N_18914,N_15462);
xnor U22016 (N_22016,N_16566,N_16732);
nor U22017 (N_22017,N_17132,N_18940);
xor U22018 (N_22018,N_17450,N_16597);
nand U22019 (N_22019,N_15021,N_16421);
nand U22020 (N_22020,N_16207,N_18748);
xnor U22021 (N_22021,N_19784,N_19054);
or U22022 (N_22022,N_18986,N_19725);
nand U22023 (N_22023,N_19276,N_17250);
nand U22024 (N_22024,N_18133,N_15225);
nand U22025 (N_22025,N_17787,N_17454);
or U22026 (N_22026,N_17314,N_19982);
or U22027 (N_22027,N_17504,N_16895);
nand U22028 (N_22028,N_15267,N_15851);
and U22029 (N_22029,N_19519,N_17906);
or U22030 (N_22030,N_19650,N_15801);
or U22031 (N_22031,N_18930,N_18534);
or U22032 (N_22032,N_19888,N_15647);
nor U22033 (N_22033,N_17853,N_19450);
xor U22034 (N_22034,N_18737,N_16661);
xor U22035 (N_22035,N_19184,N_16715);
xnor U22036 (N_22036,N_18905,N_17708);
or U22037 (N_22037,N_18249,N_15003);
nor U22038 (N_22038,N_15352,N_18255);
nor U22039 (N_22039,N_16204,N_16614);
nand U22040 (N_22040,N_18208,N_15960);
and U22041 (N_22041,N_15369,N_15242);
xnor U22042 (N_22042,N_15701,N_15606);
nor U22043 (N_22043,N_18343,N_15780);
nor U22044 (N_22044,N_18699,N_18665);
nor U22045 (N_22045,N_17754,N_18218);
or U22046 (N_22046,N_17292,N_16541);
nand U22047 (N_22047,N_16828,N_17149);
or U22048 (N_22048,N_18588,N_16709);
or U22049 (N_22049,N_18292,N_15618);
xor U22050 (N_22050,N_16951,N_15866);
and U22051 (N_22051,N_19087,N_15447);
or U22052 (N_22052,N_18862,N_17867);
xnor U22053 (N_22053,N_18734,N_17823);
or U22054 (N_22054,N_19675,N_16825);
and U22055 (N_22055,N_17384,N_19727);
nor U22056 (N_22056,N_19113,N_15935);
and U22057 (N_22057,N_19708,N_19284);
or U22058 (N_22058,N_15891,N_19994);
and U22059 (N_22059,N_17594,N_19228);
or U22060 (N_22060,N_19420,N_19045);
xnor U22061 (N_22061,N_17573,N_17628);
nand U22062 (N_22062,N_18876,N_15410);
nor U22063 (N_22063,N_17950,N_18641);
or U22064 (N_22064,N_18312,N_17406);
and U22065 (N_22065,N_19612,N_19912);
and U22066 (N_22066,N_17335,N_15620);
nand U22067 (N_22067,N_17502,N_18949);
nor U22068 (N_22068,N_18701,N_19691);
nand U22069 (N_22069,N_19178,N_16273);
and U22070 (N_22070,N_19586,N_17641);
xor U22071 (N_22071,N_18706,N_18613);
nand U22072 (N_22072,N_19324,N_15356);
xnor U22073 (N_22073,N_18599,N_15394);
nand U22074 (N_22074,N_18001,N_19973);
nand U22075 (N_22075,N_16700,N_17802);
and U22076 (N_22076,N_16656,N_16071);
nor U22077 (N_22077,N_18513,N_15362);
nand U22078 (N_22078,N_18793,N_15064);
or U22079 (N_22079,N_16780,N_15057);
and U22080 (N_22080,N_15982,N_16639);
nor U22081 (N_22081,N_15735,N_16545);
and U22082 (N_22082,N_19505,N_19151);
nor U22083 (N_22083,N_15759,N_17112);
xnor U22084 (N_22084,N_17555,N_19478);
or U22085 (N_22085,N_19438,N_16434);
and U22086 (N_22086,N_18643,N_15376);
nor U22087 (N_22087,N_17716,N_16312);
nor U22088 (N_22088,N_15408,N_18720);
or U22089 (N_22089,N_19911,N_16270);
nand U22090 (N_22090,N_16882,N_17979);
nand U22091 (N_22091,N_16681,N_16851);
nor U22092 (N_22092,N_18759,N_16822);
and U22093 (N_22093,N_16961,N_17843);
and U22094 (N_22094,N_19501,N_17228);
or U22095 (N_22095,N_15697,N_18418);
nand U22096 (N_22096,N_15284,N_17859);
nor U22097 (N_22097,N_17464,N_17021);
xor U22098 (N_22098,N_17117,N_19816);
nand U22099 (N_22099,N_18084,N_16350);
or U22100 (N_22100,N_16154,N_18724);
and U22101 (N_22101,N_17220,N_18747);
nor U22102 (N_22102,N_15105,N_17243);
nor U22103 (N_22103,N_16076,N_17023);
xnor U22104 (N_22104,N_16660,N_15022);
nand U22105 (N_22105,N_16522,N_19600);
nor U22106 (N_22106,N_18062,N_18620);
nor U22107 (N_22107,N_17433,N_18333);
and U22108 (N_22108,N_19217,N_17517);
nor U22109 (N_22109,N_15744,N_19203);
or U22110 (N_22110,N_16486,N_15446);
nor U22111 (N_22111,N_19885,N_19499);
nor U22112 (N_22112,N_18929,N_18123);
nand U22113 (N_22113,N_18685,N_18595);
xnor U22114 (N_22114,N_16899,N_17320);
and U22115 (N_22115,N_17301,N_16880);
and U22116 (N_22116,N_17764,N_15300);
and U22117 (N_22117,N_17691,N_18337);
or U22118 (N_22118,N_18100,N_17408);
and U22119 (N_22119,N_19466,N_16298);
or U22120 (N_22120,N_19544,N_15396);
nor U22121 (N_22121,N_15413,N_19017);
xor U22122 (N_22122,N_17440,N_15835);
nor U22123 (N_22123,N_18651,N_15205);
and U22124 (N_22124,N_18542,N_17085);
or U22125 (N_22125,N_19968,N_15044);
nor U22126 (N_22126,N_16642,N_19340);
nand U22127 (N_22127,N_15855,N_19769);
and U22128 (N_22128,N_16883,N_16735);
or U22129 (N_22129,N_17324,N_15336);
and U22130 (N_22130,N_15120,N_18391);
and U22131 (N_22131,N_19898,N_19970);
nor U22132 (N_22132,N_18065,N_15955);
or U22133 (N_22133,N_16491,N_16228);
nor U22134 (N_22134,N_17204,N_17558);
xnor U22135 (N_22135,N_19230,N_18565);
xnor U22136 (N_22136,N_16229,N_18199);
or U22137 (N_22137,N_16630,N_15934);
nor U22138 (N_22138,N_17476,N_18356);
nand U22139 (N_22139,N_19573,N_15575);
nand U22140 (N_22140,N_16146,N_17169);
nand U22141 (N_22141,N_19078,N_19182);
nor U22142 (N_22142,N_15531,N_16906);
nand U22143 (N_22143,N_15949,N_15709);
xnor U22144 (N_22144,N_17137,N_18029);
xnor U22145 (N_22145,N_19149,N_19298);
and U22146 (N_22146,N_16267,N_17180);
nand U22147 (N_22147,N_18814,N_19714);
xnor U22148 (N_22148,N_19559,N_16666);
or U22149 (N_22149,N_16061,N_16441);
xnor U22150 (N_22150,N_18094,N_17405);
nor U22151 (N_22151,N_18178,N_17622);
xnor U22152 (N_22152,N_17603,N_17211);
and U22153 (N_22153,N_16612,N_16200);
or U22154 (N_22154,N_17857,N_18792);
and U22155 (N_22155,N_16494,N_16805);
xnor U22156 (N_22156,N_19193,N_15052);
and U22157 (N_22157,N_17162,N_18440);
and U22158 (N_22158,N_17984,N_16920);
and U22159 (N_22159,N_19495,N_15419);
and U22160 (N_22160,N_19100,N_18214);
nor U22161 (N_22161,N_17522,N_18150);
nand U22162 (N_22162,N_15361,N_15202);
or U22163 (N_22163,N_17936,N_19400);
and U22164 (N_22164,N_15059,N_18449);
xnor U22165 (N_22165,N_17849,N_17411);
nand U22166 (N_22166,N_18188,N_16687);
xor U22167 (N_22167,N_15511,N_16520);
or U22168 (N_22168,N_17673,N_19901);
xnor U22169 (N_22169,N_16116,N_19551);
and U22170 (N_22170,N_15907,N_17743);
nor U22171 (N_22171,N_17518,N_18808);
nor U22172 (N_22172,N_19798,N_19881);
xnor U22173 (N_22173,N_17568,N_15373);
nor U22174 (N_22174,N_17586,N_18609);
and U22175 (N_22175,N_18674,N_16211);
and U22176 (N_22176,N_15082,N_15200);
and U22177 (N_22177,N_19212,N_15980);
xnor U22178 (N_22178,N_19347,N_15144);
nand U22179 (N_22179,N_15876,N_15600);
or U22180 (N_22180,N_19950,N_15623);
xnor U22181 (N_22181,N_17428,N_16242);
nor U22182 (N_22182,N_19549,N_16293);
and U22183 (N_22183,N_18196,N_19535);
or U22184 (N_22184,N_18245,N_18515);
or U22185 (N_22185,N_15122,N_18122);
nor U22186 (N_22186,N_18579,N_18550);
and U22187 (N_22187,N_15002,N_15486);
nor U22188 (N_22188,N_18241,N_17808);
xor U22189 (N_22189,N_19410,N_19215);
and U22190 (N_22190,N_16773,N_15138);
xor U22191 (N_22191,N_18490,N_19031);
and U22192 (N_22192,N_16064,N_15820);
or U22193 (N_22193,N_17790,N_19089);
or U22194 (N_22194,N_18272,N_15004);
nor U22195 (N_22195,N_16256,N_16622);
or U22196 (N_22196,N_15487,N_17345);
and U22197 (N_22197,N_16032,N_16925);
or U22198 (N_22198,N_18479,N_16193);
nand U22199 (N_22199,N_16142,N_16934);
nand U22200 (N_22200,N_16689,N_18835);
and U22201 (N_22201,N_17539,N_16777);
xor U22202 (N_22202,N_19476,N_15492);
nand U22203 (N_22203,N_18322,N_15504);
and U22204 (N_22204,N_16429,N_15199);
and U22205 (N_22205,N_18675,N_18527);
nor U22206 (N_22206,N_19403,N_18610);
and U22207 (N_22207,N_19962,N_16807);
xnor U22208 (N_22208,N_17185,N_17992);
nand U22209 (N_22209,N_19258,N_17469);
nor U22210 (N_22210,N_17579,N_17000);
or U22211 (N_22211,N_17237,N_16122);
nor U22212 (N_22212,N_15214,N_17124);
nor U22213 (N_22213,N_15377,N_16186);
nor U22214 (N_22214,N_17437,N_16691);
and U22215 (N_22215,N_17120,N_15817);
nand U22216 (N_22216,N_17424,N_16935);
nand U22217 (N_22217,N_18888,N_15857);
or U22218 (N_22218,N_16578,N_19792);
nand U22219 (N_22219,N_17280,N_15047);
nor U22220 (N_22220,N_17122,N_19770);
and U22221 (N_22221,N_17231,N_15788);
nand U22222 (N_22222,N_16531,N_18400);
xnor U22223 (N_22223,N_16926,N_15087);
and U22224 (N_22224,N_19006,N_17923);
or U22225 (N_22225,N_19061,N_17138);
nand U22226 (N_22226,N_17049,N_18881);
nor U22227 (N_22227,N_19238,N_18266);
or U22228 (N_22228,N_17993,N_16108);
and U22229 (N_22229,N_16580,N_15116);
nand U22230 (N_22230,N_15089,N_15294);
nand U22231 (N_22231,N_17140,N_18559);
and U22232 (N_22232,N_16136,N_15358);
nor U22233 (N_22233,N_18763,N_19181);
nand U22234 (N_22234,N_17547,N_16367);
and U22235 (N_22235,N_16581,N_17891);
nor U22236 (N_22236,N_15867,N_17285);
or U22237 (N_22237,N_16513,N_19439);
nor U22238 (N_22238,N_18530,N_15012);
xnor U22239 (N_22239,N_18287,N_17516);
xor U22240 (N_22240,N_17567,N_18144);
xor U22241 (N_22241,N_19703,N_17595);
or U22242 (N_22242,N_19491,N_15236);
nor U22243 (N_22243,N_18046,N_17933);
nand U22244 (N_22244,N_15050,N_18184);
nand U22245 (N_22245,N_17760,N_16497);
or U22246 (N_22246,N_18868,N_15532);
and U22247 (N_22247,N_16659,N_19449);
nor U22248 (N_22248,N_16162,N_17240);
xnor U22249 (N_22249,N_18945,N_18676);
and U22250 (N_22250,N_19200,N_15416);
and U22251 (N_22251,N_17624,N_19253);
and U22252 (N_22252,N_15390,N_17199);
nand U22253 (N_22253,N_16764,N_19448);
nand U22254 (N_22254,N_18277,N_19746);
xor U22255 (N_22255,N_15518,N_15979);
nand U22256 (N_22256,N_16426,N_17265);
or U22257 (N_22257,N_18828,N_18549);
or U22258 (N_22258,N_17957,N_17741);
xor U22259 (N_22259,N_18571,N_17847);
nor U22260 (N_22260,N_19751,N_15696);
xnor U22261 (N_22261,N_19754,N_18365);
nand U22262 (N_22262,N_15459,N_18781);
xnor U22263 (N_22263,N_17404,N_17275);
nor U22264 (N_22264,N_15508,N_18601);
and U22265 (N_22265,N_17678,N_17489);
nor U22266 (N_22266,N_15493,N_15327);
and U22267 (N_22267,N_15946,N_15102);
xor U22268 (N_22268,N_16558,N_15382);
nor U22269 (N_22269,N_19590,N_17967);
or U22270 (N_22270,N_17981,N_15261);
or U22271 (N_22271,N_18003,N_16182);
and U22272 (N_22272,N_17770,N_19517);
or U22273 (N_22273,N_18126,N_18691);
and U22274 (N_22274,N_16217,N_17018);
or U22275 (N_22275,N_18308,N_18727);
or U22276 (N_22276,N_18526,N_16077);
or U22277 (N_22277,N_15684,N_18173);
or U22278 (N_22278,N_19660,N_16375);
nand U22279 (N_22279,N_18647,N_15145);
nor U22280 (N_22280,N_16235,N_16685);
or U22281 (N_22281,N_18206,N_17919);
or U22282 (N_22282,N_15372,N_19619);
nor U22283 (N_22283,N_15754,N_17945);
xnor U22284 (N_22284,N_17564,N_17958);
nor U22285 (N_22285,N_19821,N_19383);
or U22286 (N_22286,N_17686,N_19678);
nor U22287 (N_22287,N_15811,N_16540);
nor U22288 (N_22288,N_18561,N_17311);
or U22289 (N_22289,N_17570,N_16530);
xnor U22290 (N_22290,N_17806,N_16726);
nand U22291 (N_22291,N_15846,N_18078);
or U22292 (N_22292,N_16236,N_19227);
and U22293 (N_22293,N_17063,N_16918);
and U22294 (N_22294,N_19731,N_19748);
nor U22295 (N_22295,N_18590,N_15569);
or U22296 (N_22296,N_17372,N_16569);
nand U22297 (N_22297,N_15340,N_17097);
and U22298 (N_22298,N_18570,N_17396);
xor U22299 (N_22299,N_16658,N_15622);
and U22300 (N_22300,N_19591,N_16158);
nor U22301 (N_22301,N_19827,N_19803);
nor U22302 (N_22302,N_17611,N_15724);
xor U22303 (N_22303,N_15460,N_18077);
and U22304 (N_22304,N_17779,N_15726);
or U22305 (N_22305,N_18481,N_15017);
xor U22306 (N_22306,N_17115,N_18360);
nand U22307 (N_22307,N_19329,N_15166);
xnor U22308 (N_22308,N_15406,N_16871);
nor U22309 (N_22309,N_19719,N_16778);
and U22310 (N_22310,N_19437,N_17485);
and U22311 (N_22311,N_17056,N_17195);
xor U22312 (N_22312,N_19236,N_19423);
xor U22313 (N_22313,N_15119,N_16845);
nor U22314 (N_22314,N_15449,N_16439);
nor U22315 (N_22315,N_16288,N_17270);
and U22316 (N_22316,N_17379,N_19047);
xor U22317 (N_22317,N_16830,N_19137);
nand U22318 (N_22318,N_15247,N_15020);
xor U22319 (N_22319,N_19808,N_15387);
nand U22320 (N_22320,N_18457,N_15576);
nand U22321 (N_22321,N_19287,N_19303);
nor U22322 (N_22322,N_17336,N_19262);
and U22323 (N_22323,N_19475,N_17481);
and U22324 (N_22324,N_17239,N_15832);
nor U22325 (N_22325,N_17592,N_19878);
xnor U22326 (N_22326,N_15315,N_16299);
xor U22327 (N_22327,N_18696,N_16593);
nor U22328 (N_22328,N_18325,N_18823);
nor U22329 (N_22329,N_18965,N_15977);
or U22330 (N_22330,N_19392,N_16163);
nor U22331 (N_22331,N_15043,N_16840);
nand U22332 (N_22332,N_18694,N_16276);
nor U22333 (N_22333,N_17397,N_17533);
xnor U22334 (N_22334,N_18671,N_15699);
and U22335 (N_22335,N_18769,N_16821);
nor U22336 (N_22336,N_17892,N_16006);
nand U22337 (N_22337,N_19295,N_16259);
xor U22338 (N_22338,N_17901,N_18934);
or U22339 (N_22339,N_16442,N_15747);
nor U22340 (N_22340,N_17395,N_17986);
nand U22341 (N_22341,N_17548,N_15001);
or U22342 (N_22342,N_19443,N_18520);
nand U22343 (N_22343,N_15183,N_19194);
nor U22344 (N_22344,N_16634,N_19046);
nand U22345 (N_22345,N_15609,N_15863);
nand U22346 (N_22346,N_19473,N_19469);
and U22347 (N_22347,N_19246,N_16501);
nor U22348 (N_22348,N_18067,N_17436);
nor U22349 (N_22349,N_16889,N_16904);
or U22350 (N_22350,N_19684,N_15878);
or U22351 (N_22351,N_17457,N_17111);
and U22352 (N_22352,N_19724,N_16010);
nor U22353 (N_22353,N_18924,N_15244);
nor U22354 (N_22354,N_19314,N_16827);
nand U22355 (N_22355,N_19697,N_19791);
or U22356 (N_22356,N_17575,N_17329);
xor U22357 (N_22357,N_19024,N_18320);
nor U22358 (N_22358,N_17198,N_19004);
and U22359 (N_22359,N_17287,N_18369);
and U22360 (N_22360,N_18213,N_18380);
or U22361 (N_22361,N_19419,N_18264);
nand U22362 (N_22362,N_16388,N_15928);
or U22363 (N_22363,N_17921,N_18796);
xnor U22364 (N_22364,N_18848,N_18842);
nor U22365 (N_22365,N_16457,N_17890);
nand U22366 (N_22366,N_18915,N_15426);
nand U22367 (N_22367,N_18857,N_19921);
and U22368 (N_22368,N_15124,N_18110);
or U22369 (N_22369,N_19283,N_18683);
xnor U22370 (N_22370,N_15739,N_16890);
or U22371 (N_22371,N_18323,N_17493);
nand U22372 (N_22372,N_18153,N_16521);
and U22373 (N_22373,N_16191,N_19198);
nor U22374 (N_22374,N_15345,N_15440);
nand U22375 (N_22375,N_16029,N_18619);
or U22376 (N_22376,N_18994,N_16834);
nand U22377 (N_22377,N_19567,N_19244);
nand U22378 (N_22378,N_17367,N_18917);
nor U22379 (N_22379,N_15156,N_15639);
and U22380 (N_22380,N_16296,N_15451);
nand U22381 (N_22381,N_15847,N_16631);
and U22382 (N_22382,N_19362,N_19686);
or U22383 (N_22383,N_16201,N_18397);
and U22384 (N_22384,N_18838,N_17911);
and U22385 (N_22385,N_17038,N_15889);
xnor U22386 (N_22386,N_18437,N_15415);
or U22387 (N_22387,N_16107,N_16750);
xor U22388 (N_22388,N_17422,N_18979);
xor U22389 (N_22389,N_17525,N_16965);
and U22390 (N_22390,N_15692,N_19829);
and U22391 (N_22391,N_15179,N_19084);
or U22392 (N_22392,N_17737,N_18600);
nor U22393 (N_22393,N_19220,N_17895);
nand U22394 (N_22394,N_17713,N_15135);
and U22395 (N_22395,N_15113,N_16533);
nand U22396 (N_22396,N_19321,N_16813);
or U22397 (N_22397,N_16590,N_18712);
xor U22398 (N_22398,N_16516,N_15283);
nand U22399 (N_22399,N_19219,N_17160);
nand U22400 (N_22400,N_18431,N_16932);
and U22401 (N_22401,N_15734,N_18733);
nand U22402 (N_22402,N_17346,N_16470);
or U22403 (N_22403,N_16102,N_19404);
and U22404 (N_22404,N_15520,N_15716);
nor U22405 (N_22405,N_18101,N_18261);
xor U22406 (N_22406,N_17763,N_18508);
nand U22407 (N_22407,N_15010,N_19772);
nor U22408 (N_22408,N_17392,N_17083);
nand U22409 (N_22409,N_17707,N_18050);
or U22410 (N_22410,N_17722,N_16132);
nand U22411 (N_22411,N_17931,N_19711);
or U22412 (N_22412,N_16718,N_18446);
and U22413 (N_22413,N_17065,N_16257);
and U22414 (N_22414,N_15324,N_16379);
nor U22415 (N_22415,N_17451,N_15279);
nor U22416 (N_22416,N_16334,N_16438);
and U22417 (N_22417,N_18120,N_17954);
xnor U22418 (N_22418,N_19116,N_18162);
xnor U22419 (N_22419,N_19907,N_19857);
and U22420 (N_22420,N_17234,N_18058);
or U22421 (N_22421,N_18946,N_15636);
or U22422 (N_22422,N_17348,N_17222);
nand U22423 (N_22423,N_19918,N_18645);
nand U22424 (N_22424,N_16854,N_16386);
nand U22425 (N_22425,N_16338,N_17131);
nand U22426 (N_22426,N_17303,N_17723);
or U22427 (N_22427,N_19979,N_19709);
xor U22428 (N_22428,N_19971,N_15429);
or U22429 (N_22429,N_18999,N_19154);
and U22430 (N_22430,N_15104,N_17753);
nor U22431 (N_22431,N_16125,N_15067);
nor U22432 (N_22432,N_16023,N_15483);
nor U22433 (N_22433,N_18328,N_18017);
nand U22434 (N_22434,N_18950,N_15830);
or U22435 (N_22435,N_15506,N_19385);
xor U22436 (N_22436,N_15799,N_15545);
and U22437 (N_22437,N_18690,N_15553);
nor U22438 (N_22438,N_17746,N_15566);
or U22439 (N_22439,N_15496,N_18169);
and U22440 (N_22440,N_18401,N_17171);
and U22441 (N_22441,N_18031,N_15621);
nand U22442 (N_22442,N_17289,N_17205);
nor U22443 (N_22443,N_15731,N_15190);
nor U22444 (N_22444,N_18704,N_15901);
nor U22445 (N_22445,N_15272,N_16385);
xor U22446 (N_22446,N_19871,N_19271);
or U22447 (N_22447,N_19939,N_17178);
or U22448 (N_22448,N_19248,N_18339);
xnor U22449 (N_22449,N_17634,N_15298);
and U22450 (N_22450,N_19337,N_16303);
xnor U22451 (N_22451,N_17256,N_15898);
nor U22452 (N_22452,N_19841,N_16066);
xnor U22453 (N_22453,N_18021,N_19716);
or U22454 (N_22454,N_19521,N_16785);
and U22455 (N_22455,N_15514,N_15075);
nand U22456 (N_22456,N_17468,N_17985);
xnor U22457 (N_22457,N_15904,N_17648);
nor U22458 (N_22458,N_16471,N_16258);
and U22459 (N_22459,N_16663,N_16289);
nor U22460 (N_22460,N_15254,N_18006);
or U22461 (N_22461,N_17299,N_16301);
and U22462 (N_22462,N_18897,N_15364);
nor U22463 (N_22463,N_17466,N_15762);
and U22464 (N_22464,N_15843,N_19371);
or U22465 (N_22465,N_18548,N_16384);
nor U22466 (N_22466,N_17067,N_16998);
and U22467 (N_22467,N_17520,N_17271);
nor U22468 (N_22468,N_19072,N_18539);
and U22469 (N_22469,N_19522,N_19850);
and U22470 (N_22470,N_17383,N_16339);
nor U22471 (N_22471,N_17261,N_17357);
nor U22472 (N_22472,N_15301,N_18281);
nand U22473 (N_22473,N_17156,N_19086);
nand U22474 (N_22474,N_19300,N_19722);
xor U22475 (N_22475,N_15427,N_16953);
xnor U22476 (N_22476,N_18650,N_18672);
and U22477 (N_22477,N_17976,N_18132);
nand U22478 (N_22478,N_18970,N_19020);
or U22479 (N_22479,N_17718,N_18215);
nand U22480 (N_22480,N_19656,N_17935);
nand U22481 (N_22481,N_15868,N_18149);
nand U22482 (N_22482,N_19413,N_16092);
or U22483 (N_22483,N_19704,N_18803);
nor U22484 (N_22484,N_19308,N_15676);
or U22485 (N_22485,N_18818,N_17591);
and U22486 (N_22486,N_16811,N_15299);
and U22487 (N_22487,N_17970,N_15019);
nand U22488 (N_22488,N_15404,N_16005);
nand U22489 (N_22489,N_18420,N_15332);
or U22490 (N_22490,N_17368,N_18282);
nand U22491 (N_22491,N_17047,N_16452);
nand U22492 (N_22492,N_19336,N_18426);
xor U22493 (N_22493,N_17604,N_16428);
xor U22494 (N_22494,N_18079,N_16402);
nor U22495 (N_22495,N_18195,N_18091);
and U22496 (N_22496,N_19811,N_19585);
or U22497 (N_22497,N_15515,N_19743);
nor U22498 (N_22498,N_15793,N_18806);
and U22499 (N_22499,N_18560,N_19233);
xnor U22500 (N_22500,N_18106,N_19073);
or U22501 (N_22501,N_17774,N_19654);
or U22502 (N_22502,N_15505,N_19525);
and U22503 (N_22503,N_15396,N_18021);
and U22504 (N_22504,N_17337,N_18327);
xor U22505 (N_22505,N_15281,N_18482);
nor U22506 (N_22506,N_19533,N_19142);
and U22507 (N_22507,N_15762,N_16139);
nand U22508 (N_22508,N_16910,N_17487);
or U22509 (N_22509,N_17106,N_15628);
and U22510 (N_22510,N_15968,N_17489);
nor U22511 (N_22511,N_17583,N_19487);
or U22512 (N_22512,N_19909,N_19624);
nand U22513 (N_22513,N_19952,N_17033);
or U22514 (N_22514,N_19068,N_18680);
nor U22515 (N_22515,N_17022,N_19858);
nor U22516 (N_22516,N_16834,N_17093);
or U22517 (N_22517,N_18858,N_17085);
xor U22518 (N_22518,N_16889,N_15105);
xnor U22519 (N_22519,N_19711,N_17888);
nor U22520 (N_22520,N_19859,N_16258);
nand U22521 (N_22521,N_19613,N_18854);
or U22522 (N_22522,N_18744,N_18978);
or U22523 (N_22523,N_17441,N_17264);
xor U22524 (N_22524,N_15354,N_17850);
or U22525 (N_22525,N_16084,N_19542);
nor U22526 (N_22526,N_19481,N_18760);
nor U22527 (N_22527,N_15479,N_16515);
or U22528 (N_22528,N_17429,N_16205);
nand U22529 (N_22529,N_18498,N_16355);
nor U22530 (N_22530,N_17101,N_15964);
nand U22531 (N_22531,N_17569,N_15133);
nor U22532 (N_22532,N_18221,N_16604);
and U22533 (N_22533,N_16659,N_18547);
or U22534 (N_22534,N_15788,N_16208);
nor U22535 (N_22535,N_19241,N_15208);
nor U22536 (N_22536,N_17359,N_18716);
nand U22537 (N_22537,N_15571,N_18997);
nand U22538 (N_22538,N_19963,N_15198);
or U22539 (N_22539,N_15700,N_19508);
and U22540 (N_22540,N_19609,N_17880);
xor U22541 (N_22541,N_17704,N_15776);
nand U22542 (N_22542,N_18834,N_16600);
nand U22543 (N_22543,N_16074,N_15661);
or U22544 (N_22544,N_18024,N_15853);
or U22545 (N_22545,N_15872,N_16299);
nor U22546 (N_22546,N_18748,N_19100);
or U22547 (N_22547,N_16032,N_17106);
nor U22548 (N_22548,N_15113,N_18014);
or U22549 (N_22549,N_16708,N_18632);
and U22550 (N_22550,N_19151,N_16872);
or U22551 (N_22551,N_18792,N_16312);
nor U22552 (N_22552,N_19774,N_16168);
nand U22553 (N_22553,N_19383,N_17563);
or U22554 (N_22554,N_18943,N_18444);
and U22555 (N_22555,N_18732,N_18842);
xor U22556 (N_22556,N_19367,N_19194);
nor U22557 (N_22557,N_16314,N_18965);
nor U22558 (N_22558,N_16665,N_15229);
xnor U22559 (N_22559,N_19575,N_15533);
nand U22560 (N_22560,N_18573,N_19253);
xor U22561 (N_22561,N_18073,N_16458);
nand U22562 (N_22562,N_15801,N_16059);
nand U22563 (N_22563,N_17608,N_17516);
and U22564 (N_22564,N_17303,N_18116);
xor U22565 (N_22565,N_17263,N_15689);
or U22566 (N_22566,N_15469,N_15547);
xor U22567 (N_22567,N_18381,N_16198);
or U22568 (N_22568,N_18948,N_19031);
nand U22569 (N_22569,N_18019,N_17115);
and U22570 (N_22570,N_16308,N_18550);
nand U22571 (N_22571,N_16371,N_15501);
and U22572 (N_22572,N_15842,N_15264);
xnor U22573 (N_22573,N_16401,N_18474);
xor U22574 (N_22574,N_18364,N_17148);
nand U22575 (N_22575,N_19901,N_15504);
or U22576 (N_22576,N_16241,N_17435);
and U22577 (N_22577,N_15501,N_15351);
nor U22578 (N_22578,N_15023,N_15237);
and U22579 (N_22579,N_19423,N_19726);
nand U22580 (N_22580,N_16302,N_18736);
and U22581 (N_22581,N_18955,N_17506);
nand U22582 (N_22582,N_19207,N_19290);
or U22583 (N_22583,N_17647,N_17481);
nand U22584 (N_22584,N_19029,N_17823);
xor U22585 (N_22585,N_17235,N_16823);
xor U22586 (N_22586,N_17587,N_16056);
or U22587 (N_22587,N_16588,N_16479);
or U22588 (N_22588,N_16135,N_17360);
nor U22589 (N_22589,N_18549,N_17937);
xnor U22590 (N_22590,N_18081,N_18825);
nand U22591 (N_22591,N_16670,N_15767);
or U22592 (N_22592,N_16583,N_19348);
or U22593 (N_22593,N_18054,N_17795);
nand U22594 (N_22594,N_16416,N_15013);
or U22595 (N_22595,N_18523,N_18660);
nor U22596 (N_22596,N_19246,N_15930);
and U22597 (N_22597,N_19982,N_15789);
xor U22598 (N_22598,N_16227,N_19861);
nor U22599 (N_22599,N_15596,N_17248);
nor U22600 (N_22600,N_15441,N_17024);
or U22601 (N_22601,N_19252,N_17061);
nor U22602 (N_22602,N_17045,N_17968);
xnor U22603 (N_22603,N_18556,N_16916);
nand U22604 (N_22604,N_17202,N_17121);
xnor U22605 (N_22605,N_19550,N_19830);
xor U22606 (N_22606,N_18156,N_18394);
and U22607 (N_22607,N_15428,N_17764);
and U22608 (N_22608,N_16118,N_16824);
nand U22609 (N_22609,N_16865,N_15438);
nor U22610 (N_22610,N_18237,N_18440);
nor U22611 (N_22611,N_15474,N_19815);
xor U22612 (N_22612,N_19925,N_19616);
xor U22613 (N_22613,N_16725,N_17990);
or U22614 (N_22614,N_17329,N_16668);
or U22615 (N_22615,N_19535,N_18456);
nand U22616 (N_22616,N_17107,N_15231);
nor U22617 (N_22617,N_15545,N_15176);
nor U22618 (N_22618,N_15524,N_18385);
xnor U22619 (N_22619,N_16243,N_18183);
nand U22620 (N_22620,N_17770,N_19557);
nor U22621 (N_22621,N_16030,N_16273);
and U22622 (N_22622,N_16887,N_15330);
or U22623 (N_22623,N_17752,N_17506);
nor U22624 (N_22624,N_15599,N_18042);
nand U22625 (N_22625,N_18303,N_19785);
xor U22626 (N_22626,N_18763,N_16708);
or U22627 (N_22627,N_16173,N_18231);
nand U22628 (N_22628,N_19335,N_19295);
xor U22629 (N_22629,N_19495,N_17070);
nand U22630 (N_22630,N_16128,N_19821);
and U22631 (N_22631,N_17679,N_19076);
nor U22632 (N_22632,N_17124,N_15281);
and U22633 (N_22633,N_15838,N_17987);
nor U22634 (N_22634,N_17623,N_19360);
nand U22635 (N_22635,N_15372,N_16681);
and U22636 (N_22636,N_18818,N_19310);
nand U22637 (N_22637,N_18572,N_16531);
and U22638 (N_22638,N_16699,N_15466);
nor U22639 (N_22639,N_15933,N_16077);
nand U22640 (N_22640,N_17863,N_17339);
nand U22641 (N_22641,N_15064,N_18320);
and U22642 (N_22642,N_19989,N_17864);
nor U22643 (N_22643,N_18075,N_17205);
xnor U22644 (N_22644,N_19111,N_16939);
or U22645 (N_22645,N_15655,N_16520);
nand U22646 (N_22646,N_16897,N_17131);
nor U22647 (N_22647,N_16619,N_19920);
nor U22648 (N_22648,N_18580,N_19368);
nand U22649 (N_22649,N_19500,N_17826);
or U22650 (N_22650,N_16787,N_15140);
nand U22651 (N_22651,N_15862,N_15130);
nor U22652 (N_22652,N_19488,N_16065);
xnor U22653 (N_22653,N_15047,N_17216);
and U22654 (N_22654,N_17413,N_16991);
nand U22655 (N_22655,N_17881,N_17030);
nand U22656 (N_22656,N_19584,N_19197);
nand U22657 (N_22657,N_18159,N_19327);
nand U22658 (N_22658,N_15887,N_17547);
and U22659 (N_22659,N_17921,N_19067);
xnor U22660 (N_22660,N_16104,N_19269);
and U22661 (N_22661,N_19673,N_19031);
nand U22662 (N_22662,N_15030,N_19091);
nand U22663 (N_22663,N_17783,N_17313);
xor U22664 (N_22664,N_16855,N_19090);
xnor U22665 (N_22665,N_15793,N_18515);
or U22666 (N_22666,N_17539,N_19461);
or U22667 (N_22667,N_19881,N_16884);
nor U22668 (N_22668,N_17866,N_16722);
nor U22669 (N_22669,N_19259,N_19897);
nor U22670 (N_22670,N_19266,N_18623);
nand U22671 (N_22671,N_17522,N_19857);
xor U22672 (N_22672,N_15819,N_18012);
or U22673 (N_22673,N_17072,N_17667);
xor U22674 (N_22674,N_19816,N_17723);
nor U22675 (N_22675,N_16859,N_18859);
nand U22676 (N_22676,N_19141,N_16666);
nor U22677 (N_22677,N_15879,N_19447);
nor U22678 (N_22678,N_19302,N_16587);
xnor U22679 (N_22679,N_15487,N_19532);
nor U22680 (N_22680,N_18003,N_19504);
xor U22681 (N_22681,N_18342,N_17765);
nor U22682 (N_22682,N_19202,N_18159);
nor U22683 (N_22683,N_18812,N_18579);
xor U22684 (N_22684,N_17620,N_19303);
nor U22685 (N_22685,N_16053,N_19261);
nand U22686 (N_22686,N_15622,N_18639);
nand U22687 (N_22687,N_17898,N_15883);
or U22688 (N_22688,N_17575,N_15054);
nand U22689 (N_22689,N_17263,N_18030);
or U22690 (N_22690,N_15020,N_17106);
and U22691 (N_22691,N_19455,N_18864);
xor U22692 (N_22692,N_18500,N_17562);
xor U22693 (N_22693,N_16398,N_19333);
and U22694 (N_22694,N_19926,N_19837);
or U22695 (N_22695,N_17088,N_19090);
or U22696 (N_22696,N_17272,N_16294);
xnor U22697 (N_22697,N_15557,N_15910);
xnor U22698 (N_22698,N_19103,N_18728);
and U22699 (N_22699,N_18709,N_15058);
nand U22700 (N_22700,N_17729,N_19039);
or U22701 (N_22701,N_18695,N_16732);
and U22702 (N_22702,N_15746,N_16083);
nor U22703 (N_22703,N_15172,N_18579);
nor U22704 (N_22704,N_16021,N_16563);
or U22705 (N_22705,N_15696,N_16016);
nand U22706 (N_22706,N_18484,N_19936);
nand U22707 (N_22707,N_19702,N_17813);
and U22708 (N_22708,N_19588,N_17717);
xor U22709 (N_22709,N_16684,N_18712);
xnor U22710 (N_22710,N_16486,N_17024);
and U22711 (N_22711,N_16328,N_15416);
or U22712 (N_22712,N_18352,N_17181);
and U22713 (N_22713,N_15489,N_16713);
and U22714 (N_22714,N_16807,N_19591);
or U22715 (N_22715,N_19289,N_18490);
nor U22716 (N_22716,N_18421,N_18854);
or U22717 (N_22717,N_17067,N_15146);
and U22718 (N_22718,N_15414,N_17779);
or U22719 (N_22719,N_16734,N_18201);
or U22720 (N_22720,N_17241,N_16867);
nand U22721 (N_22721,N_15502,N_15053);
or U22722 (N_22722,N_15225,N_17147);
nor U22723 (N_22723,N_15512,N_17429);
or U22724 (N_22724,N_15355,N_18196);
nor U22725 (N_22725,N_16419,N_16560);
nand U22726 (N_22726,N_15628,N_19044);
nand U22727 (N_22727,N_17346,N_18494);
or U22728 (N_22728,N_18431,N_16973);
or U22729 (N_22729,N_19443,N_18788);
xnor U22730 (N_22730,N_17094,N_19401);
or U22731 (N_22731,N_18594,N_19060);
and U22732 (N_22732,N_18533,N_15590);
xnor U22733 (N_22733,N_19361,N_16911);
nand U22734 (N_22734,N_16048,N_19556);
nor U22735 (N_22735,N_18050,N_18864);
nor U22736 (N_22736,N_19885,N_19626);
nand U22737 (N_22737,N_15197,N_15771);
nor U22738 (N_22738,N_15206,N_16232);
or U22739 (N_22739,N_15345,N_16367);
nand U22740 (N_22740,N_19523,N_18014);
nor U22741 (N_22741,N_19942,N_15805);
nand U22742 (N_22742,N_16065,N_16020);
nand U22743 (N_22743,N_15755,N_19726);
nand U22744 (N_22744,N_19512,N_15003);
nor U22745 (N_22745,N_16653,N_19156);
xnor U22746 (N_22746,N_17142,N_15249);
and U22747 (N_22747,N_18306,N_19714);
and U22748 (N_22748,N_18051,N_17247);
nand U22749 (N_22749,N_16816,N_18474);
and U22750 (N_22750,N_16725,N_16059);
and U22751 (N_22751,N_16340,N_15332);
and U22752 (N_22752,N_18024,N_19010);
or U22753 (N_22753,N_18765,N_18435);
nand U22754 (N_22754,N_16725,N_18019);
xnor U22755 (N_22755,N_19481,N_19239);
nand U22756 (N_22756,N_17216,N_18770);
and U22757 (N_22757,N_18617,N_16334);
nor U22758 (N_22758,N_17007,N_16916);
nand U22759 (N_22759,N_18095,N_16967);
xnor U22760 (N_22760,N_18916,N_19235);
nor U22761 (N_22761,N_15643,N_19852);
or U22762 (N_22762,N_15252,N_16109);
xor U22763 (N_22763,N_16234,N_19991);
nand U22764 (N_22764,N_19323,N_16662);
nand U22765 (N_22765,N_18124,N_15576);
nor U22766 (N_22766,N_16163,N_19555);
and U22767 (N_22767,N_19294,N_17286);
xnor U22768 (N_22768,N_17253,N_19563);
nand U22769 (N_22769,N_15103,N_18609);
and U22770 (N_22770,N_18961,N_18037);
or U22771 (N_22771,N_17430,N_15642);
and U22772 (N_22772,N_19854,N_19493);
and U22773 (N_22773,N_15635,N_19119);
nor U22774 (N_22774,N_17317,N_16781);
or U22775 (N_22775,N_16369,N_16506);
nand U22776 (N_22776,N_17891,N_16788);
nand U22777 (N_22777,N_19354,N_17760);
nand U22778 (N_22778,N_16154,N_15785);
nand U22779 (N_22779,N_19067,N_18148);
or U22780 (N_22780,N_17843,N_18181);
xnor U22781 (N_22781,N_18892,N_18684);
xor U22782 (N_22782,N_17922,N_17935);
nand U22783 (N_22783,N_19128,N_17988);
nor U22784 (N_22784,N_16247,N_15797);
or U22785 (N_22785,N_18209,N_17536);
xor U22786 (N_22786,N_15604,N_19440);
nand U22787 (N_22787,N_19165,N_18682);
nand U22788 (N_22788,N_15088,N_15907);
nor U22789 (N_22789,N_16983,N_17141);
nand U22790 (N_22790,N_18880,N_19372);
or U22791 (N_22791,N_16046,N_18711);
or U22792 (N_22792,N_16843,N_15806);
and U22793 (N_22793,N_18734,N_18685);
or U22794 (N_22794,N_16424,N_19255);
xnor U22795 (N_22795,N_16790,N_18981);
or U22796 (N_22796,N_19608,N_16118);
nor U22797 (N_22797,N_19145,N_18790);
xor U22798 (N_22798,N_15249,N_16216);
nand U22799 (N_22799,N_16665,N_19033);
nor U22800 (N_22800,N_17513,N_18497);
nor U22801 (N_22801,N_16806,N_16292);
and U22802 (N_22802,N_18073,N_15051);
or U22803 (N_22803,N_15755,N_18508);
nor U22804 (N_22804,N_18046,N_16684);
xor U22805 (N_22805,N_17151,N_15965);
and U22806 (N_22806,N_17201,N_17012);
nor U22807 (N_22807,N_19373,N_18069);
or U22808 (N_22808,N_18660,N_18693);
nor U22809 (N_22809,N_16017,N_15727);
nand U22810 (N_22810,N_18168,N_18432);
or U22811 (N_22811,N_17409,N_15773);
nor U22812 (N_22812,N_17404,N_16539);
or U22813 (N_22813,N_15108,N_19097);
xor U22814 (N_22814,N_15970,N_18910);
nand U22815 (N_22815,N_17749,N_19446);
and U22816 (N_22816,N_17476,N_18717);
nor U22817 (N_22817,N_18362,N_15602);
or U22818 (N_22818,N_16781,N_19541);
and U22819 (N_22819,N_16884,N_17437);
xor U22820 (N_22820,N_16870,N_15361);
and U22821 (N_22821,N_17255,N_18594);
or U22822 (N_22822,N_17583,N_15495);
xor U22823 (N_22823,N_15949,N_18567);
xor U22824 (N_22824,N_16974,N_15392);
nand U22825 (N_22825,N_17322,N_17158);
or U22826 (N_22826,N_18517,N_19182);
xnor U22827 (N_22827,N_19397,N_19157);
nor U22828 (N_22828,N_19013,N_17982);
and U22829 (N_22829,N_16360,N_19508);
nand U22830 (N_22830,N_16118,N_16659);
nor U22831 (N_22831,N_17690,N_18607);
and U22832 (N_22832,N_19840,N_18211);
nor U22833 (N_22833,N_15558,N_18824);
xor U22834 (N_22834,N_16919,N_16243);
or U22835 (N_22835,N_15070,N_16051);
nand U22836 (N_22836,N_17689,N_17981);
nand U22837 (N_22837,N_15857,N_18100);
xor U22838 (N_22838,N_17917,N_17498);
nor U22839 (N_22839,N_18930,N_17624);
or U22840 (N_22840,N_15863,N_17021);
or U22841 (N_22841,N_18503,N_19323);
nand U22842 (N_22842,N_17633,N_16024);
nand U22843 (N_22843,N_15622,N_15271);
nand U22844 (N_22844,N_18471,N_19689);
and U22845 (N_22845,N_17349,N_15622);
nand U22846 (N_22846,N_18688,N_15453);
xnor U22847 (N_22847,N_19807,N_15669);
and U22848 (N_22848,N_19586,N_17206);
nand U22849 (N_22849,N_17604,N_16065);
xor U22850 (N_22850,N_17425,N_15948);
xnor U22851 (N_22851,N_16178,N_17623);
nand U22852 (N_22852,N_15005,N_15633);
xor U22853 (N_22853,N_15765,N_17449);
xnor U22854 (N_22854,N_17513,N_18285);
nand U22855 (N_22855,N_17124,N_15683);
and U22856 (N_22856,N_17091,N_16559);
and U22857 (N_22857,N_19639,N_17511);
and U22858 (N_22858,N_16933,N_16573);
nor U22859 (N_22859,N_16254,N_17972);
xnor U22860 (N_22860,N_18375,N_17374);
nor U22861 (N_22861,N_16594,N_17689);
or U22862 (N_22862,N_19808,N_15256);
and U22863 (N_22863,N_17522,N_17676);
nand U22864 (N_22864,N_15977,N_16927);
and U22865 (N_22865,N_16119,N_18486);
or U22866 (N_22866,N_17075,N_18790);
and U22867 (N_22867,N_17634,N_18632);
and U22868 (N_22868,N_17303,N_17610);
nor U22869 (N_22869,N_15565,N_19661);
nand U22870 (N_22870,N_18877,N_17262);
or U22871 (N_22871,N_19331,N_16841);
and U22872 (N_22872,N_16242,N_19536);
xor U22873 (N_22873,N_15882,N_19850);
or U22874 (N_22874,N_19321,N_15494);
and U22875 (N_22875,N_17280,N_15340);
xor U22876 (N_22876,N_18378,N_15518);
or U22877 (N_22877,N_17877,N_17727);
or U22878 (N_22878,N_16885,N_15259);
nand U22879 (N_22879,N_17581,N_19516);
or U22880 (N_22880,N_19171,N_17392);
and U22881 (N_22881,N_17162,N_16397);
xnor U22882 (N_22882,N_19065,N_16249);
nand U22883 (N_22883,N_16320,N_16531);
or U22884 (N_22884,N_19728,N_18691);
nor U22885 (N_22885,N_16723,N_19331);
nand U22886 (N_22886,N_17335,N_19218);
xor U22887 (N_22887,N_16729,N_16087);
nor U22888 (N_22888,N_19804,N_15300);
nand U22889 (N_22889,N_16619,N_16512);
and U22890 (N_22890,N_18225,N_16698);
and U22891 (N_22891,N_15417,N_17532);
and U22892 (N_22892,N_17371,N_15633);
nand U22893 (N_22893,N_19250,N_18197);
nor U22894 (N_22894,N_19741,N_19032);
or U22895 (N_22895,N_16922,N_17411);
nand U22896 (N_22896,N_18017,N_17101);
or U22897 (N_22897,N_19488,N_17712);
and U22898 (N_22898,N_17848,N_16278);
and U22899 (N_22899,N_18271,N_16439);
nor U22900 (N_22900,N_15386,N_16078);
nand U22901 (N_22901,N_16660,N_18029);
nor U22902 (N_22902,N_18100,N_19532);
nand U22903 (N_22903,N_15972,N_15303);
nand U22904 (N_22904,N_16556,N_16452);
xor U22905 (N_22905,N_19990,N_15106);
xor U22906 (N_22906,N_16465,N_15188);
nand U22907 (N_22907,N_18702,N_16047);
nand U22908 (N_22908,N_17296,N_17284);
nor U22909 (N_22909,N_19297,N_15338);
nand U22910 (N_22910,N_17019,N_15216);
nor U22911 (N_22911,N_16874,N_19479);
xor U22912 (N_22912,N_19790,N_18811);
xor U22913 (N_22913,N_18441,N_18772);
nor U22914 (N_22914,N_18117,N_17425);
nand U22915 (N_22915,N_18298,N_17492);
and U22916 (N_22916,N_19105,N_15648);
nand U22917 (N_22917,N_19288,N_17471);
or U22918 (N_22918,N_19285,N_19708);
nor U22919 (N_22919,N_15482,N_15337);
xnor U22920 (N_22920,N_19221,N_19410);
and U22921 (N_22921,N_15392,N_18877);
and U22922 (N_22922,N_17892,N_15852);
nand U22923 (N_22923,N_16582,N_17649);
nand U22924 (N_22924,N_18212,N_16475);
and U22925 (N_22925,N_19944,N_19860);
nor U22926 (N_22926,N_16149,N_19253);
and U22927 (N_22927,N_19849,N_16294);
nand U22928 (N_22928,N_15323,N_15033);
xnor U22929 (N_22929,N_15383,N_15875);
xnor U22930 (N_22930,N_19272,N_18075);
or U22931 (N_22931,N_17223,N_17414);
xor U22932 (N_22932,N_19790,N_15856);
and U22933 (N_22933,N_18810,N_15229);
or U22934 (N_22934,N_17926,N_17218);
xor U22935 (N_22935,N_16494,N_19254);
or U22936 (N_22936,N_19962,N_15472);
or U22937 (N_22937,N_17531,N_19612);
nor U22938 (N_22938,N_17521,N_15646);
nor U22939 (N_22939,N_18641,N_16625);
nor U22940 (N_22940,N_16038,N_19728);
or U22941 (N_22941,N_17910,N_16269);
or U22942 (N_22942,N_19949,N_19293);
nor U22943 (N_22943,N_17682,N_15846);
xnor U22944 (N_22944,N_15326,N_15091);
nand U22945 (N_22945,N_17925,N_18475);
and U22946 (N_22946,N_19387,N_18088);
nor U22947 (N_22947,N_15247,N_18624);
nor U22948 (N_22948,N_16708,N_19870);
nor U22949 (N_22949,N_18399,N_18329);
or U22950 (N_22950,N_18686,N_19087);
xnor U22951 (N_22951,N_18062,N_16828);
nor U22952 (N_22952,N_16429,N_16376);
or U22953 (N_22953,N_17352,N_19682);
nor U22954 (N_22954,N_15680,N_19278);
xnor U22955 (N_22955,N_18476,N_18859);
or U22956 (N_22956,N_19030,N_19124);
and U22957 (N_22957,N_15378,N_19514);
or U22958 (N_22958,N_17207,N_15115);
and U22959 (N_22959,N_16466,N_19312);
xor U22960 (N_22960,N_18069,N_17565);
xnor U22961 (N_22961,N_15287,N_17358);
or U22962 (N_22962,N_16741,N_19328);
nand U22963 (N_22963,N_16070,N_18249);
nor U22964 (N_22964,N_19054,N_18429);
nand U22965 (N_22965,N_19394,N_15932);
and U22966 (N_22966,N_15328,N_16022);
nor U22967 (N_22967,N_19468,N_19777);
and U22968 (N_22968,N_17021,N_15834);
and U22969 (N_22969,N_19391,N_19777);
nand U22970 (N_22970,N_17636,N_19611);
and U22971 (N_22971,N_18435,N_17690);
nand U22972 (N_22972,N_15816,N_16132);
nand U22973 (N_22973,N_16659,N_19910);
or U22974 (N_22974,N_16748,N_15711);
or U22975 (N_22975,N_19370,N_18679);
and U22976 (N_22976,N_17269,N_18277);
nand U22977 (N_22977,N_15462,N_18067);
xnor U22978 (N_22978,N_16525,N_16234);
and U22979 (N_22979,N_19742,N_16942);
nand U22980 (N_22980,N_16620,N_18420);
or U22981 (N_22981,N_17095,N_16452);
or U22982 (N_22982,N_16901,N_17591);
nand U22983 (N_22983,N_17876,N_17984);
or U22984 (N_22984,N_19354,N_19345);
or U22985 (N_22985,N_16069,N_19997);
and U22986 (N_22986,N_17269,N_19911);
and U22987 (N_22987,N_15677,N_18641);
or U22988 (N_22988,N_15401,N_15422);
or U22989 (N_22989,N_16679,N_16823);
nand U22990 (N_22990,N_15646,N_17310);
or U22991 (N_22991,N_17153,N_19599);
or U22992 (N_22992,N_18530,N_19854);
and U22993 (N_22993,N_18845,N_16339);
or U22994 (N_22994,N_19740,N_19410);
and U22995 (N_22995,N_16179,N_16965);
and U22996 (N_22996,N_17292,N_16798);
xor U22997 (N_22997,N_15756,N_19026);
and U22998 (N_22998,N_19507,N_19723);
xor U22999 (N_22999,N_15337,N_18563);
nand U23000 (N_23000,N_16952,N_16607);
and U23001 (N_23001,N_16691,N_19450);
or U23002 (N_23002,N_18787,N_16322);
and U23003 (N_23003,N_15053,N_17584);
or U23004 (N_23004,N_18603,N_17166);
nand U23005 (N_23005,N_15487,N_17805);
nand U23006 (N_23006,N_16909,N_19209);
or U23007 (N_23007,N_19255,N_18248);
and U23008 (N_23008,N_19542,N_18939);
nor U23009 (N_23009,N_17056,N_18941);
xnor U23010 (N_23010,N_17633,N_19337);
nor U23011 (N_23011,N_16988,N_19203);
and U23012 (N_23012,N_16056,N_19661);
or U23013 (N_23013,N_16980,N_16101);
or U23014 (N_23014,N_19822,N_16910);
nand U23015 (N_23015,N_15038,N_17182);
nor U23016 (N_23016,N_15780,N_19531);
xnor U23017 (N_23017,N_18654,N_16743);
or U23018 (N_23018,N_18993,N_17692);
or U23019 (N_23019,N_19316,N_15570);
nor U23020 (N_23020,N_18701,N_19093);
nand U23021 (N_23021,N_17984,N_15433);
or U23022 (N_23022,N_18228,N_19218);
xor U23023 (N_23023,N_15684,N_15101);
or U23024 (N_23024,N_18064,N_16943);
xnor U23025 (N_23025,N_18738,N_17131);
or U23026 (N_23026,N_17590,N_18909);
nand U23027 (N_23027,N_16445,N_18617);
nor U23028 (N_23028,N_16049,N_19727);
xnor U23029 (N_23029,N_16242,N_16445);
or U23030 (N_23030,N_19001,N_18218);
and U23031 (N_23031,N_15137,N_17297);
xor U23032 (N_23032,N_19105,N_16184);
nand U23033 (N_23033,N_19422,N_17840);
xnor U23034 (N_23034,N_17467,N_19583);
nand U23035 (N_23035,N_19929,N_17401);
or U23036 (N_23036,N_17199,N_18068);
xnor U23037 (N_23037,N_15865,N_16630);
nor U23038 (N_23038,N_19496,N_18078);
and U23039 (N_23039,N_19270,N_17725);
xnor U23040 (N_23040,N_16769,N_19349);
and U23041 (N_23041,N_18390,N_19201);
nand U23042 (N_23042,N_16732,N_19949);
nor U23043 (N_23043,N_18184,N_15285);
nand U23044 (N_23044,N_18285,N_16591);
or U23045 (N_23045,N_19927,N_16428);
and U23046 (N_23046,N_18123,N_15065);
nor U23047 (N_23047,N_19199,N_19586);
xnor U23048 (N_23048,N_19921,N_19905);
xnor U23049 (N_23049,N_17083,N_19420);
xor U23050 (N_23050,N_16826,N_16491);
nand U23051 (N_23051,N_17439,N_15708);
nor U23052 (N_23052,N_19340,N_19816);
nor U23053 (N_23053,N_17391,N_16259);
nor U23054 (N_23054,N_15831,N_15481);
xor U23055 (N_23055,N_17643,N_17125);
nor U23056 (N_23056,N_18932,N_17658);
nor U23057 (N_23057,N_15233,N_16672);
nor U23058 (N_23058,N_15690,N_16896);
nand U23059 (N_23059,N_17157,N_19210);
nor U23060 (N_23060,N_19772,N_16038);
or U23061 (N_23061,N_19066,N_15705);
and U23062 (N_23062,N_18324,N_17294);
and U23063 (N_23063,N_15585,N_16996);
xnor U23064 (N_23064,N_18400,N_17853);
nand U23065 (N_23065,N_15704,N_17539);
and U23066 (N_23066,N_18289,N_18090);
xnor U23067 (N_23067,N_19718,N_18039);
or U23068 (N_23068,N_15160,N_19170);
and U23069 (N_23069,N_19883,N_19565);
or U23070 (N_23070,N_18323,N_17364);
and U23071 (N_23071,N_18474,N_17999);
or U23072 (N_23072,N_16609,N_15391);
nor U23073 (N_23073,N_18354,N_15793);
and U23074 (N_23074,N_16375,N_18524);
nor U23075 (N_23075,N_18318,N_19769);
nor U23076 (N_23076,N_17235,N_16551);
nand U23077 (N_23077,N_15659,N_17271);
and U23078 (N_23078,N_16629,N_17327);
xnor U23079 (N_23079,N_19067,N_16715);
xnor U23080 (N_23080,N_19453,N_17428);
or U23081 (N_23081,N_17042,N_18523);
xnor U23082 (N_23082,N_15497,N_16614);
and U23083 (N_23083,N_17233,N_18788);
nor U23084 (N_23084,N_15752,N_17127);
xnor U23085 (N_23085,N_15399,N_18695);
nor U23086 (N_23086,N_19175,N_18134);
nor U23087 (N_23087,N_15653,N_16703);
and U23088 (N_23088,N_19478,N_15958);
nand U23089 (N_23089,N_18327,N_19020);
xor U23090 (N_23090,N_17993,N_19325);
and U23091 (N_23091,N_19633,N_19567);
nand U23092 (N_23092,N_18612,N_18778);
nand U23093 (N_23093,N_15095,N_16669);
xnor U23094 (N_23094,N_19405,N_17657);
xor U23095 (N_23095,N_15137,N_17905);
and U23096 (N_23096,N_16017,N_17375);
nor U23097 (N_23097,N_17979,N_17236);
nor U23098 (N_23098,N_17681,N_15281);
or U23099 (N_23099,N_16026,N_19998);
nand U23100 (N_23100,N_17853,N_18613);
and U23101 (N_23101,N_18039,N_18687);
nand U23102 (N_23102,N_17034,N_15071);
nand U23103 (N_23103,N_19134,N_18930);
nand U23104 (N_23104,N_19333,N_16531);
nor U23105 (N_23105,N_18234,N_16311);
xnor U23106 (N_23106,N_16154,N_17155);
xnor U23107 (N_23107,N_19548,N_16285);
nor U23108 (N_23108,N_16583,N_19001);
or U23109 (N_23109,N_17244,N_15127);
or U23110 (N_23110,N_19614,N_16693);
and U23111 (N_23111,N_15949,N_16899);
xor U23112 (N_23112,N_17794,N_19377);
or U23113 (N_23113,N_16808,N_17155);
nand U23114 (N_23114,N_17243,N_18666);
nor U23115 (N_23115,N_17165,N_17052);
nand U23116 (N_23116,N_18797,N_15835);
nor U23117 (N_23117,N_16355,N_17663);
xnor U23118 (N_23118,N_17092,N_17475);
xor U23119 (N_23119,N_19190,N_19231);
xnor U23120 (N_23120,N_16332,N_18191);
nand U23121 (N_23121,N_18319,N_18219);
nor U23122 (N_23122,N_17240,N_16544);
or U23123 (N_23123,N_19912,N_17939);
or U23124 (N_23124,N_16990,N_17583);
or U23125 (N_23125,N_19853,N_17770);
nand U23126 (N_23126,N_18985,N_18865);
xor U23127 (N_23127,N_17326,N_17429);
or U23128 (N_23128,N_18837,N_16747);
or U23129 (N_23129,N_15874,N_16693);
nand U23130 (N_23130,N_19239,N_17790);
xor U23131 (N_23131,N_15553,N_17960);
nor U23132 (N_23132,N_17429,N_17317);
or U23133 (N_23133,N_18076,N_18266);
nor U23134 (N_23134,N_17814,N_17052);
xnor U23135 (N_23135,N_18417,N_15893);
nor U23136 (N_23136,N_15193,N_18966);
nor U23137 (N_23137,N_19855,N_17081);
nand U23138 (N_23138,N_19114,N_18835);
nor U23139 (N_23139,N_18812,N_15743);
xnor U23140 (N_23140,N_16785,N_15334);
nand U23141 (N_23141,N_16927,N_16217);
and U23142 (N_23142,N_19443,N_16260);
or U23143 (N_23143,N_16444,N_17219);
or U23144 (N_23144,N_16010,N_17728);
nand U23145 (N_23145,N_17472,N_15452);
and U23146 (N_23146,N_19965,N_16767);
or U23147 (N_23147,N_17567,N_19903);
nor U23148 (N_23148,N_19372,N_18727);
nand U23149 (N_23149,N_19550,N_18602);
nor U23150 (N_23150,N_19946,N_15524);
xor U23151 (N_23151,N_18687,N_16857);
nand U23152 (N_23152,N_19275,N_16661);
nor U23153 (N_23153,N_19503,N_16609);
xnor U23154 (N_23154,N_19078,N_18959);
or U23155 (N_23155,N_19728,N_19531);
and U23156 (N_23156,N_15287,N_19563);
nor U23157 (N_23157,N_19679,N_19779);
nand U23158 (N_23158,N_18652,N_17348);
nor U23159 (N_23159,N_19547,N_16285);
or U23160 (N_23160,N_19249,N_18540);
and U23161 (N_23161,N_17486,N_16393);
and U23162 (N_23162,N_15511,N_16076);
nor U23163 (N_23163,N_16327,N_17946);
and U23164 (N_23164,N_17127,N_16609);
xnor U23165 (N_23165,N_15672,N_15356);
or U23166 (N_23166,N_16748,N_17402);
or U23167 (N_23167,N_17908,N_18570);
xor U23168 (N_23168,N_18568,N_17675);
xor U23169 (N_23169,N_19775,N_17542);
xor U23170 (N_23170,N_17549,N_17820);
xor U23171 (N_23171,N_18009,N_17811);
xor U23172 (N_23172,N_18661,N_15683);
nand U23173 (N_23173,N_17894,N_17455);
nand U23174 (N_23174,N_16013,N_16947);
or U23175 (N_23175,N_15727,N_19644);
nand U23176 (N_23176,N_17576,N_19573);
and U23177 (N_23177,N_19017,N_16678);
or U23178 (N_23178,N_16657,N_18802);
or U23179 (N_23179,N_16840,N_19397);
xor U23180 (N_23180,N_15744,N_18093);
xnor U23181 (N_23181,N_18038,N_16380);
nand U23182 (N_23182,N_18430,N_16426);
and U23183 (N_23183,N_17017,N_15371);
nand U23184 (N_23184,N_15184,N_17704);
and U23185 (N_23185,N_15548,N_18881);
xnor U23186 (N_23186,N_15062,N_15813);
and U23187 (N_23187,N_15148,N_16977);
or U23188 (N_23188,N_17648,N_16101);
or U23189 (N_23189,N_17526,N_18940);
nor U23190 (N_23190,N_17564,N_19007);
or U23191 (N_23191,N_16220,N_17490);
xor U23192 (N_23192,N_16337,N_19442);
xnor U23193 (N_23193,N_15791,N_19669);
or U23194 (N_23194,N_18857,N_19700);
or U23195 (N_23195,N_16069,N_16862);
and U23196 (N_23196,N_16494,N_15374);
nor U23197 (N_23197,N_16470,N_17758);
xnor U23198 (N_23198,N_16801,N_15467);
nor U23199 (N_23199,N_16443,N_17266);
or U23200 (N_23200,N_18051,N_17633);
xor U23201 (N_23201,N_18704,N_19782);
and U23202 (N_23202,N_15343,N_19929);
and U23203 (N_23203,N_17426,N_15331);
xnor U23204 (N_23204,N_19345,N_18923);
nor U23205 (N_23205,N_16070,N_16358);
nor U23206 (N_23206,N_16911,N_15033);
and U23207 (N_23207,N_16544,N_18374);
and U23208 (N_23208,N_16882,N_19275);
nand U23209 (N_23209,N_15202,N_18598);
nor U23210 (N_23210,N_16245,N_19153);
nor U23211 (N_23211,N_17565,N_17359);
nand U23212 (N_23212,N_18879,N_17137);
nand U23213 (N_23213,N_15098,N_15331);
and U23214 (N_23214,N_18712,N_15211);
xnor U23215 (N_23215,N_15079,N_19530);
xnor U23216 (N_23216,N_18337,N_15275);
xor U23217 (N_23217,N_17063,N_17294);
and U23218 (N_23218,N_18352,N_15861);
and U23219 (N_23219,N_17674,N_19097);
nor U23220 (N_23220,N_15101,N_16010);
or U23221 (N_23221,N_15546,N_16333);
and U23222 (N_23222,N_18969,N_15482);
nor U23223 (N_23223,N_16579,N_17435);
and U23224 (N_23224,N_15901,N_18598);
nand U23225 (N_23225,N_16341,N_16862);
xor U23226 (N_23226,N_15709,N_15041);
and U23227 (N_23227,N_17416,N_16269);
and U23228 (N_23228,N_19317,N_15517);
nor U23229 (N_23229,N_16339,N_15240);
or U23230 (N_23230,N_16882,N_17844);
nor U23231 (N_23231,N_18183,N_19996);
and U23232 (N_23232,N_15836,N_16597);
xor U23233 (N_23233,N_15069,N_18278);
xor U23234 (N_23234,N_16012,N_15914);
xor U23235 (N_23235,N_18071,N_18183);
nor U23236 (N_23236,N_19456,N_16241);
nand U23237 (N_23237,N_18539,N_16543);
nor U23238 (N_23238,N_18447,N_18344);
xor U23239 (N_23239,N_17101,N_19784);
xor U23240 (N_23240,N_19206,N_17319);
nand U23241 (N_23241,N_15140,N_15981);
nand U23242 (N_23242,N_19845,N_15868);
nand U23243 (N_23243,N_19672,N_18561);
and U23244 (N_23244,N_17273,N_18164);
and U23245 (N_23245,N_15504,N_17310);
xnor U23246 (N_23246,N_19464,N_18027);
nor U23247 (N_23247,N_19600,N_18732);
xor U23248 (N_23248,N_17455,N_18397);
or U23249 (N_23249,N_15645,N_17016);
nor U23250 (N_23250,N_15227,N_15193);
nor U23251 (N_23251,N_17325,N_19050);
xor U23252 (N_23252,N_19786,N_19197);
xnor U23253 (N_23253,N_17313,N_18920);
nor U23254 (N_23254,N_19737,N_17340);
and U23255 (N_23255,N_17491,N_15523);
and U23256 (N_23256,N_19574,N_16104);
nand U23257 (N_23257,N_17277,N_15866);
nand U23258 (N_23258,N_15442,N_17019);
or U23259 (N_23259,N_16832,N_15277);
nor U23260 (N_23260,N_15350,N_16861);
and U23261 (N_23261,N_18159,N_16830);
xor U23262 (N_23262,N_18727,N_16792);
nor U23263 (N_23263,N_19296,N_19200);
nor U23264 (N_23264,N_15461,N_19228);
and U23265 (N_23265,N_15540,N_18353);
nand U23266 (N_23266,N_19739,N_17079);
and U23267 (N_23267,N_15965,N_17740);
and U23268 (N_23268,N_19162,N_17516);
xor U23269 (N_23269,N_19172,N_16123);
xor U23270 (N_23270,N_15181,N_16567);
or U23271 (N_23271,N_18691,N_17181);
nor U23272 (N_23272,N_19769,N_15488);
xnor U23273 (N_23273,N_19409,N_18370);
nand U23274 (N_23274,N_17006,N_16148);
and U23275 (N_23275,N_17014,N_17207);
xor U23276 (N_23276,N_17158,N_19235);
nor U23277 (N_23277,N_18000,N_18382);
or U23278 (N_23278,N_15828,N_19211);
nand U23279 (N_23279,N_17251,N_16703);
xnor U23280 (N_23280,N_19404,N_19804);
or U23281 (N_23281,N_15754,N_19157);
nand U23282 (N_23282,N_19929,N_15043);
xor U23283 (N_23283,N_16206,N_15775);
and U23284 (N_23284,N_19265,N_19232);
nor U23285 (N_23285,N_19422,N_19296);
or U23286 (N_23286,N_18103,N_17810);
and U23287 (N_23287,N_16247,N_18762);
nand U23288 (N_23288,N_15042,N_19472);
xnor U23289 (N_23289,N_17284,N_15069);
or U23290 (N_23290,N_16361,N_17306);
nand U23291 (N_23291,N_19901,N_18854);
nand U23292 (N_23292,N_15154,N_19686);
xor U23293 (N_23293,N_16575,N_17975);
and U23294 (N_23294,N_15101,N_17921);
xor U23295 (N_23295,N_16742,N_16290);
nand U23296 (N_23296,N_16330,N_15212);
xnor U23297 (N_23297,N_16935,N_19219);
xor U23298 (N_23298,N_16915,N_15282);
and U23299 (N_23299,N_15715,N_15293);
and U23300 (N_23300,N_18168,N_18123);
nor U23301 (N_23301,N_15426,N_15095);
nor U23302 (N_23302,N_15928,N_15100);
nand U23303 (N_23303,N_15848,N_18167);
nand U23304 (N_23304,N_19952,N_19628);
and U23305 (N_23305,N_18155,N_16384);
nor U23306 (N_23306,N_15712,N_18963);
and U23307 (N_23307,N_16726,N_19584);
and U23308 (N_23308,N_19352,N_15707);
or U23309 (N_23309,N_18885,N_15762);
nand U23310 (N_23310,N_19304,N_17092);
or U23311 (N_23311,N_16623,N_18299);
and U23312 (N_23312,N_15183,N_18421);
nand U23313 (N_23313,N_16230,N_19482);
or U23314 (N_23314,N_16051,N_15560);
xor U23315 (N_23315,N_15704,N_16186);
xnor U23316 (N_23316,N_17137,N_15696);
or U23317 (N_23317,N_17137,N_16616);
and U23318 (N_23318,N_19606,N_17958);
or U23319 (N_23319,N_15594,N_17496);
or U23320 (N_23320,N_15877,N_17185);
nand U23321 (N_23321,N_19975,N_16928);
xor U23322 (N_23322,N_18300,N_19998);
xnor U23323 (N_23323,N_17221,N_19406);
nand U23324 (N_23324,N_18746,N_17384);
and U23325 (N_23325,N_19143,N_18577);
and U23326 (N_23326,N_16713,N_16613);
or U23327 (N_23327,N_19812,N_16710);
and U23328 (N_23328,N_17866,N_19213);
or U23329 (N_23329,N_19279,N_17065);
and U23330 (N_23330,N_19242,N_15737);
and U23331 (N_23331,N_19064,N_18097);
nor U23332 (N_23332,N_15777,N_18268);
or U23333 (N_23333,N_15999,N_18592);
nand U23334 (N_23334,N_16360,N_16782);
nor U23335 (N_23335,N_18211,N_16647);
nor U23336 (N_23336,N_16217,N_15728);
and U23337 (N_23337,N_18110,N_16416);
xnor U23338 (N_23338,N_19727,N_16086);
nand U23339 (N_23339,N_18588,N_16392);
nor U23340 (N_23340,N_18990,N_16524);
and U23341 (N_23341,N_15324,N_17250);
nor U23342 (N_23342,N_17328,N_17044);
nand U23343 (N_23343,N_16372,N_19498);
nor U23344 (N_23344,N_16561,N_16741);
xnor U23345 (N_23345,N_16847,N_18959);
xnor U23346 (N_23346,N_16167,N_16919);
and U23347 (N_23347,N_18702,N_17404);
xor U23348 (N_23348,N_19870,N_17275);
nor U23349 (N_23349,N_19732,N_19144);
nor U23350 (N_23350,N_18719,N_16359);
or U23351 (N_23351,N_19127,N_19628);
or U23352 (N_23352,N_15461,N_19425);
nand U23353 (N_23353,N_18241,N_19468);
and U23354 (N_23354,N_17356,N_18483);
and U23355 (N_23355,N_18830,N_16349);
xnor U23356 (N_23356,N_16124,N_15821);
or U23357 (N_23357,N_16708,N_19748);
nand U23358 (N_23358,N_19741,N_15074);
xor U23359 (N_23359,N_17109,N_15779);
or U23360 (N_23360,N_16013,N_18114);
nor U23361 (N_23361,N_16334,N_19429);
xnor U23362 (N_23362,N_17792,N_18129);
or U23363 (N_23363,N_19138,N_17011);
nand U23364 (N_23364,N_15191,N_18566);
and U23365 (N_23365,N_16428,N_15909);
nor U23366 (N_23366,N_16912,N_16024);
or U23367 (N_23367,N_18283,N_18234);
xnor U23368 (N_23368,N_16557,N_18823);
and U23369 (N_23369,N_18867,N_17953);
and U23370 (N_23370,N_15956,N_16740);
nor U23371 (N_23371,N_15465,N_15576);
and U23372 (N_23372,N_16054,N_17722);
nor U23373 (N_23373,N_18844,N_17137);
xor U23374 (N_23374,N_15525,N_15683);
and U23375 (N_23375,N_19575,N_19174);
nand U23376 (N_23376,N_17836,N_16679);
xor U23377 (N_23377,N_19793,N_18426);
and U23378 (N_23378,N_18326,N_17978);
nor U23379 (N_23379,N_18395,N_16679);
nand U23380 (N_23380,N_17164,N_19438);
or U23381 (N_23381,N_18348,N_18829);
and U23382 (N_23382,N_19244,N_16266);
or U23383 (N_23383,N_16617,N_15613);
nand U23384 (N_23384,N_15509,N_18410);
and U23385 (N_23385,N_19429,N_15927);
nand U23386 (N_23386,N_15540,N_17418);
and U23387 (N_23387,N_15496,N_15864);
and U23388 (N_23388,N_18124,N_17316);
nor U23389 (N_23389,N_17049,N_17484);
xnor U23390 (N_23390,N_15773,N_18688);
xnor U23391 (N_23391,N_18808,N_15841);
xor U23392 (N_23392,N_19283,N_16976);
or U23393 (N_23393,N_16360,N_19502);
or U23394 (N_23394,N_19922,N_17742);
or U23395 (N_23395,N_15906,N_19562);
xnor U23396 (N_23396,N_18096,N_16891);
nand U23397 (N_23397,N_19165,N_15673);
nand U23398 (N_23398,N_15629,N_15059);
xnor U23399 (N_23399,N_16323,N_19831);
nor U23400 (N_23400,N_18682,N_16284);
nand U23401 (N_23401,N_17881,N_17738);
and U23402 (N_23402,N_17568,N_19138);
or U23403 (N_23403,N_17686,N_19883);
nand U23404 (N_23404,N_16504,N_16670);
and U23405 (N_23405,N_15252,N_17872);
nand U23406 (N_23406,N_18840,N_19550);
or U23407 (N_23407,N_18620,N_18070);
xnor U23408 (N_23408,N_15410,N_18125);
xor U23409 (N_23409,N_17792,N_19536);
or U23410 (N_23410,N_19686,N_15265);
or U23411 (N_23411,N_17942,N_19420);
nand U23412 (N_23412,N_16218,N_16416);
or U23413 (N_23413,N_15245,N_15042);
nor U23414 (N_23414,N_16266,N_16155);
and U23415 (N_23415,N_18043,N_15141);
nand U23416 (N_23416,N_19047,N_19096);
nor U23417 (N_23417,N_15239,N_18963);
and U23418 (N_23418,N_18631,N_18658);
nand U23419 (N_23419,N_16730,N_15339);
nor U23420 (N_23420,N_18152,N_19374);
or U23421 (N_23421,N_15457,N_17572);
or U23422 (N_23422,N_16632,N_16447);
nand U23423 (N_23423,N_17946,N_15707);
nand U23424 (N_23424,N_15827,N_19374);
and U23425 (N_23425,N_17647,N_15461);
and U23426 (N_23426,N_16552,N_19091);
xnor U23427 (N_23427,N_17566,N_17999);
and U23428 (N_23428,N_17780,N_19086);
xor U23429 (N_23429,N_15484,N_16300);
nor U23430 (N_23430,N_17803,N_17060);
xor U23431 (N_23431,N_19645,N_19814);
xnor U23432 (N_23432,N_16026,N_15023);
and U23433 (N_23433,N_17885,N_17350);
nor U23434 (N_23434,N_15457,N_19325);
xor U23435 (N_23435,N_16754,N_18366);
and U23436 (N_23436,N_16460,N_19662);
nand U23437 (N_23437,N_19079,N_16541);
xnor U23438 (N_23438,N_18221,N_15183);
nor U23439 (N_23439,N_18442,N_17112);
or U23440 (N_23440,N_15693,N_16344);
xnor U23441 (N_23441,N_18120,N_17060);
nand U23442 (N_23442,N_19440,N_18825);
nand U23443 (N_23443,N_16924,N_18524);
or U23444 (N_23444,N_18382,N_18995);
xor U23445 (N_23445,N_17071,N_17210);
nor U23446 (N_23446,N_17682,N_19367);
xnor U23447 (N_23447,N_19462,N_17332);
nor U23448 (N_23448,N_16564,N_18643);
nand U23449 (N_23449,N_19945,N_18989);
and U23450 (N_23450,N_17915,N_19410);
or U23451 (N_23451,N_15999,N_17278);
and U23452 (N_23452,N_15541,N_15090);
xor U23453 (N_23453,N_16088,N_17223);
and U23454 (N_23454,N_16654,N_18426);
xnor U23455 (N_23455,N_15003,N_19669);
and U23456 (N_23456,N_18593,N_17136);
nor U23457 (N_23457,N_15437,N_15883);
or U23458 (N_23458,N_16502,N_16527);
nor U23459 (N_23459,N_19423,N_16268);
nor U23460 (N_23460,N_18609,N_18354);
or U23461 (N_23461,N_15606,N_18527);
or U23462 (N_23462,N_19493,N_18740);
and U23463 (N_23463,N_16036,N_17871);
nor U23464 (N_23464,N_19870,N_19029);
and U23465 (N_23465,N_19197,N_16040);
or U23466 (N_23466,N_17391,N_18364);
nor U23467 (N_23467,N_18701,N_19532);
nor U23468 (N_23468,N_16596,N_15795);
nor U23469 (N_23469,N_17020,N_16014);
or U23470 (N_23470,N_15343,N_16513);
and U23471 (N_23471,N_17670,N_19005);
nand U23472 (N_23472,N_19096,N_19387);
or U23473 (N_23473,N_15368,N_15809);
and U23474 (N_23474,N_17058,N_15288);
nand U23475 (N_23475,N_15266,N_17095);
nand U23476 (N_23476,N_15888,N_15402);
nand U23477 (N_23477,N_16094,N_19434);
or U23478 (N_23478,N_18300,N_18559);
xnor U23479 (N_23479,N_19476,N_19253);
xnor U23480 (N_23480,N_19213,N_18142);
and U23481 (N_23481,N_18702,N_17786);
or U23482 (N_23482,N_17291,N_15962);
and U23483 (N_23483,N_18852,N_18134);
nand U23484 (N_23484,N_16078,N_18023);
nand U23485 (N_23485,N_15046,N_15297);
xnor U23486 (N_23486,N_16519,N_19918);
or U23487 (N_23487,N_17601,N_18161);
or U23488 (N_23488,N_16423,N_15269);
or U23489 (N_23489,N_18156,N_15145);
nand U23490 (N_23490,N_18173,N_18780);
or U23491 (N_23491,N_19535,N_19043);
nand U23492 (N_23492,N_18157,N_17415);
or U23493 (N_23493,N_19049,N_15682);
nand U23494 (N_23494,N_17888,N_16396);
xnor U23495 (N_23495,N_16191,N_19089);
xnor U23496 (N_23496,N_15300,N_18711);
or U23497 (N_23497,N_18253,N_18109);
xnor U23498 (N_23498,N_19462,N_19884);
or U23499 (N_23499,N_18870,N_18638);
and U23500 (N_23500,N_17233,N_17754);
nor U23501 (N_23501,N_19011,N_19342);
and U23502 (N_23502,N_19875,N_17962);
or U23503 (N_23503,N_15233,N_17319);
or U23504 (N_23504,N_17437,N_16472);
and U23505 (N_23505,N_19777,N_18571);
xnor U23506 (N_23506,N_16304,N_17747);
and U23507 (N_23507,N_15938,N_15446);
or U23508 (N_23508,N_16121,N_16627);
and U23509 (N_23509,N_18245,N_18026);
nor U23510 (N_23510,N_16463,N_17215);
and U23511 (N_23511,N_18265,N_19346);
or U23512 (N_23512,N_15541,N_18858);
or U23513 (N_23513,N_18815,N_16158);
nor U23514 (N_23514,N_19442,N_15874);
and U23515 (N_23515,N_16484,N_19733);
nor U23516 (N_23516,N_19877,N_19237);
nand U23517 (N_23517,N_17129,N_18457);
xor U23518 (N_23518,N_18811,N_18551);
and U23519 (N_23519,N_15418,N_17033);
nand U23520 (N_23520,N_19598,N_16308);
xor U23521 (N_23521,N_18239,N_15345);
xnor U23522 (N_23522,N_16828,N_19155);
nand U23523 (N_23523,N_18787,N_17807);
xnor U23524 (N_23524,N_18192,N_16899);
xor U23525 (N_23525,N_17427,N_17730);
nand U23526 (N_23526,N_17288,N_18602);
and U23527 (N_23527,N_19287,N_15885);
or U23528 (N_23528,N_16526,N_17059);
nor U23529 (N_23529,N_16579,N_19276);
and U23530 (N_23530,N_19397,N_15794);
or U23531 (N_23531,N_18569,N_15729);
nand U23532 (N_23532,N_15316,N_16345);
xor U23533 (N_23533,N_16280,N_16709);
or U23534 (N_23534,N_19279,N_16304);
or U23535 (N_23535,N_16413,N_16185);
xor U23536 (N_23536,N_16233,N_16221);
and U23537 (N_23537,N_17698,N_16473);
or U23538 (N_23538,N_16279,N_15220);
and U23539 (N_23539,N_18336,N_16486);
nand U23540 (N_23540,N_19803,N_18206);
nor U23541 (N_23541,N_17333,N_19871);
and U23542 (N_23542,N_19088,N_15935);
and U23543 (N_23543,N_16307,N_17515);
nor U23544 (N_23544,N_16059,N_17923);
or U23545 (N_23545,N_18022,N_15035);
nand U23546 (N_23546,N_19429,N_16923);
nand U23547 (N_23547,N_15002,N_18118);
xnor U23548 (N_23548,N_15670,N_18723);
or U23549 (N_23549,N_15610,N_17893);
nand U23550 (N_23550,N_17490,N_19792);
nor U23551 (N_23551,N_18465,N_18150);
and U23552 (N_23552,N_18884,N_19793);
xor U23553 (N_23553,N_19005,N_17142);
nand U23554 (N_23554,N_18460,N_16481);
and U23555 (N_23555,N_16590,N_17196);
nand U23556 (N_23556,N_15165,N_17918);
xnor U23557 (N_23557,N_15391,N_17906);
nor U23558 (N_23558,N_18514,N_15026);
nor U23559 (N_23559,N_15052,N_15266);
and U23560 (N_23560,N_15914,N_18388);
or U23561 (N_23561,N_17302,N_19309);
nand U23562 (N_23562,N_17827,N_18662);
nor U23563 (N_23563,N_16727,N_18780);
nand U23564 (N_23564,N_17235,N_19135);
nand U23565 (N_23565,N_19855,N_19976);
nand U23566 (N_23566,N_16758,N_18974);
nand U23567 (N_23567,N_18648,N_17345);
xnor U23568 (N_23568,N_18863,N_16484);
and U23569 (N_23569,N_18458,N_15240);
xor U23570 (N_23570,N_19284,N_15337);
nand U23571 (N_23571,N_19080,N_19467);
or U23572 (N_23572,N_17842,N_15527);
xor U23573 (N_23573,N_19990,N_16621);
nand U23574 (N_23574,N_16755,N_17981);
or U23575 (N_23575,N_15227,N_19986);
nand U23576 (N_23576,N_17361,N_15104);
nor U23577 (N_23577,N_18321,N_15689);
and U23578 (N_23578,N_18020,N_17264);
nand U23579 (N_23579,N_16883,N_18096);
or U23580 (N_23580,N_18378,N_17958);
nor U23581 (N_23581,N_17738,N_16072);
or U23582 (N_23582,N_15534,N_18055);
nand U23583 (N_23583,N_19022,N_15692);
or U23584 (N_23584,N_17832,N_16300);
nand U23585 (N_23585,N_15501,N_17229);
nor U23586 (N_23586,N_18922,N_16933);
nand U23587 (N_23587,N_17798,N_16440);
or U23588 (N_23588,N_16465,N_16411);
nor U23589 (N_23589,N_18565,N_15788);
or U23590 (N_23590,N_18546,N_18974);
nor U23591 (N_23591,N_18575,N_19040);
or U23592 (N_23592,N_19962,N_17812);
xor U23593 (N_23593,N_17328,N_19864);
xnor U23594 (N_23594,N_18541,N_18472);
nand U23595 (N_23595,N_19717,N_17311);
nand U23596 (N_23596,N_15639,N_16892);
xnor U23597 (N_23597,N_16505,N_18958);
nor U23598 (N_23598,N_15064,N_19619);
or U23599 (N_23599,N_15325,N_19662);
nand U23600 (N_23600,N_19362,N_18430);
xnor U23601 (N_23601,N_15583,N_15180);
nand U23602 (N_23602,N_16683,N_15386);
xnor U23603 (N_23603,N_15668,N_15124);
nor U23604 (N_23604,N_19065,N_18664);
xnor U23605 (N_23605,N_15188,N_15676);
and U23606 (N_23606,N_18595,N_16887);
and U23607 (N_23607,N_15997,N_15183);
xor U23608 (N_23608,N_15840,N_15279);
and U23609 (N_23609,N_15893,N_17883);
xor U23610 (N_23610,N_16550,N_18285);
nor U23611 (N_23611,N_18708,N_17429);
and U23612 (N_23612,N_18348,N_19949);
nand U23613 (N_23613,N_15860,N_16392);
nor U23614 (N_23614,N_16336,N_18860);
and U23615 (N_23615,N_19238,N_15856);
or U23616 (N_23616,N_19188,N_17795);
and U23617 (N_23617,N_19600,N_18338);
and U23618 (N_23618,N_15845,N_18832);
xor U23619 (N_23619,N_15071,N_16943);
and U23620 (N_23620,N_17959,N_19199);
nand U23621 (N_23621,N_19535,N_16423);
nor U23622 (N_23622,N_19006,N_18807);
nor U23623 (N_23623,N_17088,N_16385);
and U23624 (N_23624,N_16968,N_17275);
or U23625 (N_23625,N_16773,N_16651);
nor U23626 (N_23626,N_17451,N_18192);
nand U23627 (N_23627,N_15255,N_18104);
or U23628 (N_23628,N_15597,N_15806);
nand U23629 (N_23629,N_16334,N_18316);
or U23630 (N_23630,N_19291,N_18679);
and U23631 (N_23631,N_19624,N_17109);
nand U23632 (N_23632,N_18515,N_17826);
nand U23633 (N_23633,N_17522,N_19809);
xnor U23634 (N_23634,N_15416,N_15058);
nand U23635 (N_23635,N_15836,N_16066);
or U23636 (N_23636,N_17511,N_19984);
nor U23637 (N_23637,N_18776,N_17737);
and U23638 (N_23638,N_15425,N_19926);
or U23639 (N_23639,N_15008,N_19520);
or U23640 (N_23640,N_15625,N_17072);
nor U23641 (N_23641,N_17612,N_17533);
nor U23642 (N_23642,N_17264,N_15799);
xor U23643 (N_23643,N_18232,N_18146);
or U23644 (N_23644,N_19709,N_17772);
and U23645 (N_23645,N_19781,N_17471);
and U23646 (N_23646,N_17089,N_16603);
and U23647 (N_23647,N_18181,N_18505);
nor U23648 (N_23648,N_19435,N_15691);
and U23649 (N_23649,N_18075,N_17915);
and U23650 (N_23650,N_19626,N_16229);
nand U23651 (N_23651,N_15533,N_15837);
xor U23652 (N_23652,N_17653,N_18779);
or U23653 (N_23653,N_17586,N_19286);
and U23654 (N_23654,N_17155,N_16428);
nor U23655 (N_23655,N_18836,N_18672);
xnor U23656 (N_23656,N_19838,N_18445);
and U23657 (N_23657,N_17020,N_16065);
nor U23658 (N_23658,N_16254,N_17494);
and U23659 (N_23659,N_17888,N_18614);
nor U23660 (N_23660,N_18111,N_19037);
xnor U23661 (N_23661,N_17106,N_17353);
xor U23662 (N_23662,N_17466,N_18380);
nand U23663 (N_23663,N_19995,N_17521);
or U23664 (N_23664,N_16740,N_15615);
or U23665 (N_23665,N_17041,N_16630);
and U23666 (N_23666,N_19926,N_17663);
nor U23667 (N_23667,N_15517,N_17623);
or U23668 (N_23668,N_17419,N_16114);
nand U23669 (N_23669,N_19168,N_18072);
and U23670 (N_23670,N_18442,N_16436);
and U23671 (N_23671,N_19061,N_18445);
or U23672 (N_23672,N_19310,N_19939);
nand U23673 (N_23673,N_18729,N_15706);
and U23674 (N_23674,N_19396,N_16339);
nor U23675 (N_23675,N_15612,N_15618);
or U23676 (N_23676,N_18980,N_18731);
xnor U23677 (N_23677,N_15834,N_15329);
nand U23678 (N_23678,N_18603,N_17373);
nand U23679 (N_23679,N_19921,N_16586);
nand U23680 (N_23680,N_18021,N_19125);
nand U23681 (N_23681,N_17762,N_18974);
nand U23682 (N_23682,N_19477,N_19711);
or U23683 (N_23683,N_17193,N_16731);
xor U23684 (N_23684,N_18643,N_18383);
and U23685 (N_23685,N_15585,N_18193);
nand U23686 (N_23686,N_16762,N_17978);
nor U23687 (N_23687,N_16607,N_18360);
and U23688 (N_23688,N_18895,N_15947);
and U23689 (N_23689,N_19860,N_18617);
or U23690 (N_23690,N_17446,N_18119);
or U23691 (N_23691,N_18785,N_16815);
nor U23692 (N_23692,N_16911,N_16421);
xnor U23693 (N_23693,N_19161,N_17479);
or U23694 (N_23694,N_15951,N_17271);
and U23695 (N_23695,N_17209,N_15174);
and U23696 (N_23696,N_15583,N_16686);
or U23697 (N_23697,N_16924,N_19810);
or U23698 (N_23698,N_16840,N_17511);
xnor U23699 (N_23699,N_15916,N_17141);
and U23700 (N_23700,N_18608,N_18302);
and U23701 (N_23701,N_17773,N_16680);
and U23702 (N_23702,N_15515,N_17783);
and U23703 (N_23703,N_15643,N_18630);
xor U23704 (N_23704,N_17833,N_16859);
xor U23705 (N_23705,N_16437,N_18066);
xor U23706 (N_23706,N_16867,N_15359);
or U23707 (N_23707,N_18709,N_16095);
or U23708 (N_23708,N_18825,N_19670);
xor U23709 (N_23709,N_19877,N_17781);
xor U23710 (N_23710,N_15619,N_15349);
and U23711 (N_23711,N_18693,N_16315);
nand U23712 (N_23712,N_18754,N_16771);
xnor U23713 (N_23713,N_16291,N_16121);
nor U23714 (N_23714,N_18614,N_16106);
nand U23715 (N_23715,N_16494,N_16498);
nand U23716 (N_23716,N_18908,N_19976);
xnor U23717 (N_23717,N_18190,N_18998);
xnor U23718 (N_23718,N_17628,N_19964);
or U23719 (N_23719,N_17275,N_16599);
nand U23720 (N_23720,N_15949,N_19391);
nor U23721 (N_23721,N_17784,N_17352);
and U23722 (N_23722,N_15260,N_15073);
nor U23723 (N_23723,N_19998,N_19960);
or U23724 (N_23724,N_16919,N_15522);
nand U23725 (N_23725,N_19543,N_16244);
xor U23726 (N_23726,N_16234,N_19757);
nand U23727 (N_23727,N_15351,N_17555);
nor U23728 (N_23728,N_15058,N_16448);
or U23729 (N_23729,N_19104,N_18169);
and U23730 (N_23730,N_15019,N_16783);
xnor U23731 (N_23731,N_15144,N_15774);
and U23732 (N_23732,N_17068,N_15282);
and U23733 (N_23733,N_19204,N_16830);
nand U23734 (N_23734,N_18215,N_18707);
or U23735 (N_23735,N_18685,N_16472);
or U23736 (N_23736,N_18610,N_18776);
and U23737 (N_23737,N_16635,N_16967);
xnor U23738 (N_23738,N_19243,N_17964);
or U23739 (N_23739,N_16615,N_16172);
nand U23740 (N_23740,N_15236,N_16587);
or U23741 (N_23741,N_15432,N_18087);
nand U23742 (N_23742,N_18787,N_18790);
nand U23743 (N_23743,N_18222,N_17403);
nand U23744 (N_23744,N_16414,N_16651);
nand U23745 (N_23745,N_19357,N_19047);
or U23746 (N_23746,N_18165,N_17261);
or U23747 (N_23747,N_16852,N_15212);
or U23748 (N_23748,N_18898,N_19647);
and U23749 (N_23749,N_19833,N_15994);
nor U23750 (N_23750,N_16804,N_16557);
nand U23751 (N_23751,N_18816,N_19743);
or U23752 (N_23752,N_15537,N_16149);
nand U23753 (N_23753,N_19090,N_18536);
nand U23754 (N_23754,N_16605,N_17104);
or U23755 (N_23755,N_18414,N_17856);
xor U23756 (N_23756,N_15482,N_16461);
xor U23757 (N_23757,N_19642,N_15315);
xnor U23758 (N_23758,N_15190,N_15872);
nor U23759 (N_23759,N_15571,N_19375);
xor U23760 (N_23760,N_15147,N_17587);
nor U23761 (N_23761,N_18604,N_18248);
and U23762 (N_23762,N_19553,N_17516);
nor U23763 (N_23763,N_17916,N_17523);
nor U23764 (N_23764,N_17834,N_18302);
nand U23765 (N_23765,N_15939,N_19064);
nor U23766 (N_23766,N_17313,N_18921);
and U23767 (N_23767,N_17763,N_15368);
and U23768 (N_23768,N_16187,N_15134);
and U23769 (N_23769,N_16962,N_16012);
or U23770 (N_23770,N_15258,N_15944);
xor U23771 (N_23771,N_19252,N_18489);
nand U23772 (N_23772,N_18918,N_15127);
nand U23773 (N_23773,N_16811,N_19434);
nand U23774 (N_23774,N_17396,N_18057);
nor U23775 (N_23775,N_17834,N_15260);
nor U23776 (N_23776,N_17677,N_15488);
or U23777 (N_23777,N_15614,N_18974);
or U23778 (N_23778,N_17350,N_18826);
and U23779 (N_23779,N_16619,N_17650);
nor U23780 (N_23780,N_15520,N_16186);
or U23781 (N_23781,N_15139,N_16736);
xor U23782 (N_23782,N_18326,N_19592);
or U23783 (N_23783,N_17673,N_17529);
or U23784 (N_23784,N_16215,N_18177);
and U23785 (N_23785,N_16620,N_15448);
and U23786 (N_23786,N_15523,N_17007);
xnor U23787 (N_23787,N_19154,N_15681);
xnor U23788 (N_23788,N_17321,N_17391);
or U23789 (N_23789,N_19178,N_16342);
or U23790 (N_23790,N_19167,N_17899);
nor U23791 (N_23791,N_17363,N_17635);
nor U23792 (N_23792,N_16734,N_16475);
or U23793 (N_23793,N_19544,N_18601);
or U23794 (N_23794,N_15478,N_16781);
xnor U23795 (N_23795,N_16480,N_18662);
nor U23796 (N_23796,N_19789,N_19040);
nand U23797 (N_23797,N_15840,N_15708);
or U23798 (N_23798,N_18281,N_15609);
xnor U23799 (N_23799,N_18105,N_19106);
nand U23800 (N_23800,N_16100,N_18761);
xnor U23801 (N_23801,N_16136,N_19715);
or U23802 (N_23802,N_16744,N_15699);
and U23803 (N_23803,N_15139,N_17036);
or U23804 (N_23804,N_17218,N_18240);
or U23805 (N_23805,N_16979,N_16227);
or U23806 (N_23806,N_18411,N_18813);
nand U23807 (N_23807,N_15010,N_15849);
nand U23808 (N_23808,N_17814,N_15656);
or U23809 (N_23809,N_19579,N_18303);
nand U23810 (N_23810,N_17237,N_17978);
and U23811 (N_23811,N_16201,N_16820);
or U23812 (N_23812,N_15791,N_15262);
and U23813 (N_23813,N_18153,N_15754);
xor U23814 (N_23814,N_16730,N_15267);
nand U23815 (N_23815,N_19915,N_18546);
nor U23816 (N_23816,N_16641,N_15369);
and U23817 (N_23817,N_17556,N_18912);
xor U23818 (N_23818,N_19211,N_19188);
nor U23819 (N_23819,N_15877,N_15198);
or U23820 (N_23820,N_15617,N_15606);
xor U23821 (N_23821,N_15992,N_15225);
and U23822 (N_23822,N_16472,N_15198);
or U23823 (N_23823,N_18623,N_16062);
and U23824 (N_23824,N_17160,N_17380);
and U23825 (N_23825,N_19982,N_19140);
or U23826 (N_23826,N_17717,N_18167);
and U23827 (N_23827,N_18112,N_19982);
xor U23828 (N_23828,N_15479,N_18200);
xor U23829 (N_23829,N_15756,N_18640);
xnor U23830 (N_23830,N_16592,N_16177);
xnor U23831 (N_23831,N_16439,N_19146);
nand U23832 (N_23832,N_16231,N_19123);
or U23833 (N_23833,N_15765,N_18337);
xor U23834 (N_23834,N_15404,N_17019);
or U23835 (N_23835,N_17457,N_16584);
xor U23836 (N_23836,N_19939,N_16735);
and U23837 (N_23837,N_18581,N_18161);
nor U23838 (N_23838,N_17882,N_18624);
nor U23839 (N_23839,N_18488,N_19035);
xor U23840 (N_23840,N_16678,N_16520);
or U23841 (N_23841,N_19016,N_18608);
and U23842 (N_23842,N_19714,N_18887);
nor U23843 (N_23843,N_15992,N_15354);
xnor U23844 (N_23844,N_17336,N_18139);
nor U23845 (N_23845,N_15693,N_19806);
and U23846 (N_23846,N_18447,N_15403);
or U23847 (N_23847,N_19348,N_17560);
xnor U23848 (N_23848,N_19437,N_15309);
nor U23849 (N_23849,N_19368,N_19262);
xnor U23850 (N_23850,N_17232,N_16881);
nand U23851 (N_23851,N_15899,N_19889);
nor U23852 (N_23852,N_15196,N_17677);
nor U23853 (N_23853,N_18821,N_15997);
and U23854 (N_23854,N_17565,N_19832);
nor U23855 (N_23855,N_19550,N_17896);
and U23856 (N_23856,N_19795,N_16032);
and U23857 (N_23857,N_15092,N_18169);
xor U23858 (N_23858,N_15693,N_17900);
xor U23859 (N_23859,N_18319,N_19930);
and U23860 (N_23860,N_19939,N_18777);
nor U23861 (N_23861,N_19607,N_17254);
or U23862 (N_23862,N_16814,N_18567);
nor U23863 (N_23863,N_16760,N_19192);
xnor U23864 (N_23864,N_19370,N_16975);
nor U23865 (N_23865,N_18666,N_16908);
xnor U23866 (N_23866,N_19289,N_17730);
or U23867 (N_23867,N_17062,N_18539);
nor U23868 (N_23868,N_15269,N_18269);
or U23869 (N_23869,N_19534,N_19911);
xor U23870 (N_23870,N_17903,N_15938);
nor U23871 (N_23871,N_19729,N_15518);
nand U23872 (N_23872,N_18327,N_16342);
xor U23873 (N_23873,N_16365,N_17470);
nor U23874 (N_23874,N_19235,N_18461);
or U23875 (N_23875,N_18964,N_17829);
and U23876 (N_23876,N_18277,N_18946);
nor U23877 (N_23877,N_17230,N_18910);
or U23878 (N_23878,N_19726,N_18300);
nand U23879 (N_23879,N_16789,N_19240);
xor U23880 (N_23880,N_17223,N_18524);
or U23881 (N_23881,N_17374,N_15428);
nor U23882 (N_23882,N_15351,N_18358);
nor U23883 (N_23883,N_17955,N_19244);
and U23884 (N_23884,N_19125,N_17435);
and U23885 (N_23885,N_16011,N_15908);
xnor U23886 (N_23886,N_17624,N_18388);
or U23887 (N_23887,N_15805,N_17636);
xor U23888 (N_23888,N_17643,N_17504);
or U23889 (N_23889,N_18072,N_16607);
nand U23890 (N_23890,N_18772,N_17739);
nand U23891 (N_23891,N_18807,N_19698);
nor U23892 (N_23892,N_18336,N_15727);
and U23893 (N_23893,N_17155,N_17335);
nor U23894 (N_23894,N_17862,N_19180);
nor U23895 (N_23895,N_15617,N_19794);
nand U23896 (N_23896,N_18308,N_19289);
and U23897 (N_23897,N_17415,N_16658);
xnor U23898 (N_23898,N_16445,N_19178);
or U23899 (N_23899,N_18834,N_16465);
nand U23900 (N_23900,N_15083,N_18297);
and U23901 (N_23901,N_19520,N_19875);
xnor U23902 (N_23902,N_17133,N_19868);
or U23903 (N_23903,N_15166,N_18588);
and U23904 (N_23904,N_16637,N_17183);
xor U23905 (N_23905,N_18052,N_15485);
and U23906 (N_23906,N_17197,N_19200);
nand U23907 (N_23907,N_15734,N_16046);
nand U23908 (N_23908,N_16421,N_17386);
and U23909 (N_23909,N_17915,N_15176);
and U23910 (N_23910,N_15446,N_19260);
or U23911 (N_23911,N_17540,N_18108);
xor U23912 (N_23912,N_19469,N_19600);
nor U23913 (N_23913,N_17596,N_16004);
or U23914 (N_23914,N_16310,N_18128);
nor U23915 (N_23915,N_18157,N_19737);
nand U23916 (N_23916,N_18546,N_16347);
xnor U23917 (N_23917,N_17310,N_15575);
nand U23918 (N_23918,N_17570,N_17685);
and U23919 (N_23919,N_16683,N_18467);
nor U23920 (N_23920,N_16086,N_17267);
and U23921 (N_23921,N_19457,N_18851);
nor U23922 (N_23922,N_18815,N_18239);
and U23923 (N_23923,N_18054,N_19673);
nand U23924 (N_23924,N_19762,N_17142);
nor U23925 (N_23925,N_18561,N_16029);
nand U23926 (N_23926,N_15227,N_19924);
xor U23927 (N_23927,N_19642,N_17713);
nor U23928 (N_23928,N_19277,N_17086);
nor U23929 (N_23929,N_18199,N_16903);
nand U23930 (N_23930,N_18220,N_15304);
and U23931 (N_23931,N_17024,N_19938);
xnor U23932 (N_23932,N_15695,N_19710);
nand U23933 (N_23933,N_15145,N_17236);
or U23934 (N_23934,N_16688,N_17861);
and U23935 (N_23935,N_17223,N_18912);
nand U23936 (N_23936,N_19877,N_18236);
nor U23937 (N_23937,N_17634,N_16021);
and U23938 (N_23938,N_17933,N_19182);
and U23939 (N_23939,N_15664,N_19066);
and U23940 (N_23940,N_19425,N_15839);
or U23941 (N_23941,N_15009,N_18379);
or U23942 (N_23942,N_15060,N_18109);
or U23943 (N_23943,N_19676,N_19033);
nor U23944 (N_23944,N_19907,N_16625);
xor U23945 (N_23945,N_19813,N_16507);
or U23946 (N_23946,N_18214,N_17280);
xnor U23947 (N_23947,N_15885,N_15112);
nor U23948 (N_23948,N_19334,N_18852);
and U23949 (N_23949,N_16879,N_18928);
nor U23950 (N_23950,N_18701,N_19948);
and U23951 (N_23951,N_16850,N_17581);
nor U23952 (N_23952,N_18909,N_16280);
or U23953 (N_23953,N_17043,N_16426);
nand U23954 (N_23954,N_15763,N_18353);
nor U23955 (N_23955,N_19734,N_19555);
xor U23956 (N_23956,N_19226,N_19095);
or U23957 (N_23957,N_18007,N_18104);
nor U23958 (N_23958,N_17017,N_18783);
nor U23959 (N_23959,N_17672,N_17629);
xnor U23960 (N_23960,N_15418,N_17092);
nor U23961 (N_23961,N_19241,N_18327);
nor U23962 (N_23962,N_15677,N_17795);
or U23963 (N_23963,N_19537,N_16566);
xnor U23964 (N_23964,N_15980,N_18079);
or U23965 (N_23965,N_15635,N_16711);
and U23966 (N_23966,N_17728,N_18868);
nor U23967 (N_23967,N_18168,N_16629);
or U23968 (N_23968,N_18847,N_18876);
nor U23969 (N_23969,N_19874,N_16401);
nand U23970 (N_23970,N_19349,N_16220);
xnor U23971 (N_23971,N_19549,N_16396);
nor U23972 (N_23972,N_16417,N_15445);
nand U23973 (N_23973,N_15601,N_19648);
and U23974 (N_23974,N_18853,N_17418);
nor U23975 (N_23975,N_16677,N_16605);
xor U23976 (N_23976,N_16173,N_16501);
xnor U23977 (N_23977,N_19815,N_19628);
nand U23978 (N_23978,N_18654,N_16023);
and U23979 (N_23979,N_17904,N_17425);
or U23980 (N_23980,N_16634,N_17922);
nor U23981 (N_23981,N_17568,N_19416);
nor U23982 (N_23982,N_18879,N_15949);
nor U23983 (N_23983,N_19583,N_16287);
or U23984 (N_23984,N_15448,N_15166);
or U23985 (N_23985,N_15200,N_17840);
xnor U23986 (N_23986,N_17560,N_19857);
nand U23987 (N_23987,N_17692,N_19985);
nand U23988 (N_23988,N_18765,N_16751);
xor U23989 (N_23989,N_16613,N_17859);
and U23990 (N_23990,N_18665,N_15381);
nor U23991 (N_23991,N_18818,N_15986);
nor U23992 (N_23992,N_16528,N_18530);
or U23993 (N_23993,N_15159,N_19625);
and U23994 (N_23994,N_19282,N_15820);
or U23995 (N_23995,N_16348,N_16686);
and U23996 (N_23996,N_17469,N_17026);
and U23997 (N_23997,N_15617,N_18771);
xor U23998 (N_23998,N_16974,N_18615);
or U23999 (N_23999,N_15480,N_18359);
nand U24000 (N_24000,N_17688,N_17361);
xor U24001 (N_24001,N_16071,N_16038);
or U24002 (N_24002,N_16049,N_16460);
and U24003 (N_24003,N_18511,N_17485);
and U24004 (N_24004,N_18306,N_19765);
nand U24005 (N_24005,N_19230,N_16494);
or U24006 (N_24006,N_18851,N_19154);
nor U24007 (N_24007,N_17948,N_19142);
xor U24008 (N_24008,N_18285,N_18273);
and U24009 (N_24009,N_18225,N_19349);
or U24010 (N_24010,N_15371,N_19657);
nor U24011 (N_24011,N_19905,N_16048);
nor U24012 (N_24012,N_18508,N_17688);
and U24013 (N_24013,N_18601,N_17254);
or U24014 (N_24014,N_16246,N_19123);
or U24015 (N_24015,N_16949,N_15948);
or U24016 (N_24016,N_17759,N_17437);
or U24017 (N_24017,N_17691,N_18873);
and U24018 (N_24018,N_16186,N_17635);
xnor U24019 (N_24019,N_16001,N_15638);
and U24020 (N_24020,N_18375,N_18372);
and U24021 (N_24021,N_17685,N_17609);
xor U24022 (N_24022,N_19125,N_19098);
xor U24023 (N_24023,N_16698,N_17065);
nor U24024 (N_24024,N_15939,N_19727);
nor U24025 (N_24025,N_15381,N_18882);
nor U24026 (N_24026,N_15556,N_17003);
nor U24027 (N_24027,N_19305,N_17670);
nor U24028 (N_24028,N_17274,N_19206);
nor U24029 (N_24029,N_16408,N_16189);
xnor U24030 (N_24030,N_16716,N_16023);
or U24031 (N_24031,N_19606,N_17394);
xor U24032 (N_24032,N_16928,N_17157);
xor U24033 (N_24033,N_16391,N_15005);
nor U24034 (N_24034,N_18955,N_16301);
and U24035 (N_24035,N_15226,N_17454);
or U24036 (N_24036,N_15291,N_16622);
nor U24037 (N_24037,N_15490,N_16776);
nand U24038 (N_24038,N_16104,N_17611);
nand U24039 (N_24039,N_17023,N_16216);
and U24040 (N_24040,N_17146,N_17944);
nand U24041 (N_24041,N_18310,N_15460);
nor U24042 (N_24042,N_15787,N_15511);
xnor U24043 (N_24043,N_16229,N_16705);
and U24044 (N_24044,N_17977,N_16773);
xor U24045 (N_24045,N_18225,N_18034);
xor U24046 (N_24046,N_17528,N_15590);
or U24047 (N_24047,N_18464,N_19496);
xor U24048 (N_24048,N_18463,N_19439);
nand U24049 (N_24049,N_18594,N_16452);
xnor U24050 (N_24050,N_16123,N_19609);
and U24051 (N_24051,N_15472,N_17560);
nand U24052 (N_24052,N_17515,N_17854);
nand U24053 (N_24053,N_19159,N_19125);
nor U24054 (N_24054,N_18045,N_17497);
nor U24055 (N_24055,N_17339,N_17731);
and U24056 (N_24056,N_17866,N_18150);
and U24057 (N_24057,N_19203,N_15556);
or U24058 (N_24058,N_15067,N_19218);
and U24059 (N_24059,N_18625,N_19174);
nand U24060 (N_24060,N_15510,N_19171);
and U24061 (N_24061,N_16872,N_19000);
or U24062 (N_24062,N_15255,N_19172);
xor U24063 (N_24063,N_17649,N_17427);
xor U24064 (N_24064,N_15849,N_15856);
nor U24065 (N_24065,N_15183,N_16726);
or U24066 (N_24066,N_18859,N_15699);
nand U24067 (N_24067,N_17850,N_19981);
nand U24068 (N_24068,N_16910,N_19439);
and U24069 (N_24069,N_16711,N_17363);
and U24070 (N_24070,N_15329,N_17713);
and U24071 (N_24071,N_17860,N_17954);
xor U24072 (N_24072,N_16264,N_17154);
or U24073 (N_24073,N_17387,N_17137);
xor U24074 (N_24074,N_19381,N_17099);
and U24075 (N_24075,N_15177,N_17304);
and U24076 (N_24076,N_19129,N_17997);
or U24077 (N_24077,N_19818,N_16029);
and U24078 (N_24078,N_19081,N_16221);
nand U24079 (N_24079,N_16285,N_19912);
xnor U24080 (N_24080,N_17210,N_16064);
or U24081 (N_24081,N_16271,N_19056);
nand U24082 (N_24082,N_15410,N_16684);
nor U24083 (N_24083,N_18696,N_16932);
and U24084 (N_24084,N_15446,N_19760);
nor U24085 (N_24085,N_19723,N_15293);
nand U24086 (N_24086,N_16918,N_16625);
and U24087 (N_24087,N_16651,N_16164);
or U24088 (N_24088,N_15231,N_16474);
and U24089 (N_24089,N_15181,N_16420);
nor U24090 (N_24090,N_19061,N_18041);
nand U24091 (N_24091,N_18270,N_15567);
nand U24092 (N_24092,N_19634,N_16368);
or U24093 (N_24093,N_15129,N_15184);
nand U24094 (N_24094,N_19416,N_18769);
and U24095 (N_24095,N_17560,N_19798);
xor U24096 (N_24096,N_17288,N_17363);
nor U24097 (N_24097,N_16852,N_18178);
xnor U24098 (N_24098,N_15902,N_15532);
xor U24099 (N_24099,N_15602,N_15952);
or U24100 (N_24100,N_16733,N_18721);
nand U24101 (N_24101,N_18021,N_19751);
nor U24102 (N_24102,N_16313,N_16176);
and U24103 (N_24103,N_16338,N_17167);
or U24104 (N_24104,N_15999,N_17946);
and U24105 (N_24105,N_19738,N_15307);
and U24106 (N_24106,N_16894,N_19423);
xnor U24107 (N_24107,N_16991,N_18872);
and U24108 (N_24108,N_17729,N_15151);
and U24109 (N_24109,N_17391,N_18935);
or U24110 (N_24110,N_18609,N_16816);
and U24111 (N_24111,N_18418,N_15905);
nor U24112 (N_24112,N_15543,N_15866);
or U24113 (N_24113,N_16886,N_19643);
nor U24114 (N_24114,N_15044,N_17916);
or U24115 (N_24115,N_17209,N_16427);
nor U24116 (N_24116,N_19425,N_19482);
or U24117 (N_24117,N_18267,N_15567);
or U24118 (N_24118,N_18155,N_16876);
xnor U24119 (N_24119,N_18752,N_19270);
or U24120 (N_24120,N_19197,N_17021);
and U24121 (N_24121,N_18644,N_18635);
and U24122 (N_24122,N_18098,N_19007);
and U24123 (N_24123,N_18760,N_18690);
or U24124 (N_24124,N_17317,N_16788);
and U24125 (N_24125,N_17122,N_19084);
xor U24126 (N_24126,N_16368,N_18622);
nor U24127 (N_24127,N_15441,N_19059);
nand U24128 (N_24128,N_17908,N_15333);
nor U24129 (N_24129,N_15820,N_17321);
or U24130 (N_24130,N_16991,N_15943);
xnor U24131 (N_24131,N_16367,N_19251);
nand U24132 (N_24132,N_17903,N_16104);
and U24133 (N_24133,N_18889,N_18175);
nor U24134 (N_24134,N_15793,N_19046);
or U24135 (N_24135,N_16747,N_18891);
nor U24136 (N_24136,N_18368,N_16608);
or U24137 (N_24137,N_15107,N_19351);
nand U24138 (N_24138,N_17182,N_16993);
or U24139 (N_24139,N_19578,N_16281);
nand U24140 (N_24140,N_19411,N_18310);
nor U24141 (N_24141,N_17681,N_17370);
xnor U24142 (N_24142,N_15883,N_16798);
or U24143 (N_24143,N_16366,N_19168);
nor U24144 (N_24144,N_15948,N_17447);
xnor U24145 (N_24145,N_16741,N_17114);
xnor U24146 (N_24146,N_19897,N_19378);
xnor U24147 (N_24147,N_18445,N_18705);
nor U24148 (N_24148,N_15260,N_19775);
xor U24149 (N_24149,N_17391,N_18459);
xor U24150 (N_24150,N_19992,N_18748);
or U24151 (N_24151,N_18882,N_16179);
or U24152 (N_24152,N_15540,N_18023);
and U24153 (N_24153,N_19409,N_15720);
xor U24154 (N_24154,N_16879,N_16609);
nor U24155 (N_24155,N_18126,N_16728);
nand U24156 (N_24156,N_15066,N_17016);
and U24157 (N_24157,N_19201,N_16276);
or U24158 (N_24158,N_16616,N_15699);
nand U24159 (N_24159,N_15017,N_15122);
or U24160 (N_24160,N_15728,N_19535);
and U24161 (N_24161,N_17572,N_18720);
xor U24162 (N_24162,N_16473,N_19380);
nand U24163 (N_24163,N_16029,N_16017);
xor U24164 (N_24164,N_15819,N_18571);
or U24165 (N_24165,N_16053,N_16510);
or U24166 (N_24166,N_15082,N_15822);
nor U24167 (N_24167,N_19244,N_16393);
or U24168 (N_24168,N_18312,N_15185);
or U24169 (N_24169,N_15412,N_18047);
nand U24170 (N_24170,N_19203,N_18294);
nor U24171 (N_24171,N_18280,N_16991);
or U24172 (N_24172,N_15395,N_18120);
nand U24173 (N_24173,N_16953,N_16803);
and U24174 (N_24174,N_17768,N_16648);
and U24175 (N_24175,N_17376,N_19131);
nand U24176 (N_24176,N_15776,N_18711);
or U24177 (N_24177,N_19259,N_18074);
xnor U24178 (N_24178,N_18356,N_19454);
or U24179 (N_24179,N_15167,N_17502);
or U24180 (N_24180,N_18892,N_19529);
nand U24181 (N_24181,N_16304,N_19320);
or U24182 (N_24182,N_15632,N_18373);
xor U24183 (N_24183,N_17611,N_19131);
xnor U24184 (N_24184,N_15378,N_16288);
and U24185 (N_24185,N_16632,N_15081);
nor U24186 (N_24186,N_16660,N_17309);
nor U24187 (N_24187,N_16292,N_18383);
xnor U24188 (N_24188,N_16308,N_19135);
nor U24189 (N_24189,N_16873,N_17146);
nor U24190 (N_24190,N_18754,N_17351);
nand U24191 (N_24191,N_19491,N_18058);
and U24192 (N_24192,N_19573,N_19409);
xor U24193 (N_24193,N_18580,N_15960);
and U24194 (N_24194,N_15352,N_16438);
nand U24195 (N_24195,N_18335,N_15640);
xnor U24196 (N_24196,N_17638,N_16897);
nor U24197 (N_24197,N_19279,N_19605);
nand U24198 (N_24198,N_19918,N_15245);
nor U24199 (N_24199,N_16070,N_19116);
nor U24200 (N_24200,N_19953,N_19448);
or U24201 (N_24201,N_18091,N_15174);
nand U24202 (N_24202,N_15578,N_19530);
and U24203 (N_24203,N_18631,N_15439);
and U24204 (N_24204,N_19663,N_19381);
and U24205 (N_24205,N_16666,N_19910);
xor U24206 (N_24206,N_18018,N_17181);
nor U24207 (N_24207,N_19558,N_17876);
or U24208 (N_24208,N_19851,N_17009);
or U24209 (N_24209,N_15982,N_16791);
nor U24210 (N_24210,N_17053,N_17774);
or U24211 (N_24211,N_17601,N_15217);
nand U24212 (N_24212,N_15502,N_15301);
nor U24213 (N_24213,N_17180,N_16828);
and U24214 (N_24214,N_19551,N_16362);
or U24215 (N_24215,N_17148,N_18477);
nand U24216 (N_24216,N_19756,N_16231);
xor U24217 (N_24217,N_17851,N_16564);
xor U24218 (N_24218,N_18105,N_19078);
or U24219 (N_24219,N_16206,N_19980);
nand U24220 (N_24220,N_19850,N_19559);
nand U24221 (N_24221,N_18100,N_16236);
or U24222 (N_24222,N_19505,N_19724);
nor U24223 (N_24223,N_16975,N_17718);
or U24224 (N_24224,N_19908,N_17129);
nand U24225 (N_24225,N_16806,N_15039);
nor U24226 (N_24226,N_19097,N_18781);
or U24227 (N_24227,N_19596,N_15618);
xor U24228 (N_24228,N_19351,N_15323);
nand U24229 (N_24229,N_19364,N_18227);
xor U24230 (N_24230,N_17309,N_17362);
and U24231 (N_24231,N_18171,N_15229);
xnor U24232 (N_24232,N_18660,N_18565);
nor U24233 (N_24233,N_18259,N_19230);
and U24234 (N_24234,N_16741,N_17231);
nand U24235 (N_24235,N_19000,N_15459);
and U24236 (N_24236,N_17529,N_18217);
nor U24237 (N_24237,N_18967,N_15064);
or U24238 (N_24238,N_17685,N_19741);
nor U24239 (N_24239,N_19349,N_18677);
xor U24240 (N_24240,N_15810,N_19428);
or U24241 (N_24241,N_16926,N_17564);
and U24242 (N_24242,N_17342,N_15568);
and U24243 (N_24243,N_19201,N_15777);
nor U24244 (N_24244,N_17595,N_18291);
nor U24245 (N_24245,N_17133,N_16867);
nand U24246 (N_24246,N_17220,N_15298);
xor U24247 (N_24247,N_16802,N_19298);
xnor U24248 (N_24248,N_18141,N_16040);
xnor U24249 (N_24249,N_18337,N_18973);
xor U24250 (N_24250,N_18993,N_17734);
xnor U24251 (N_24251,N_17729,N_15853);
nor U24252 (N_24252,N_18852,N_15448);
xnor U24253 (N_24253,N_17109,N_16117);
nor U24254 (N_24254,N_18861,N_18113);
xnor U24255 (N_24255,N_16015,N_16138);
or U24256 (N_24256,N_18218,N_18102);
xor U24257 (N_24257,N_19390,N_16819);
nand U24258 (N_24258,N_17598,N_19271);
or U24259 (N_24259,N_19331,N_18253);
and U24260 (N_24260,N_19316,N_18596);
or U24261 (N_24261,N_19124,N_16600);
nor U24262 (N_24262,N_16983,N_18956);
xnor U24263 (N_24263,N_15089,N_15287);
nor U24264 (N_24264,N_18478,N_16853);
and U24265 (N_24265,N_15491,N_15059);
nand U24266 (N_24266,N_15556,N_17941);
or U24267 (N_24267,N_16901,N_17559);
xor U24268 (N_24268,N_18248,N_18738);
nor U24269 (N_24269,N_16755,N_19915);
xnor U24270 (N_24270,N_15003,N_17583);
nand U24271 (N_24271,N_19307,N_18090);
nand U24272 (N_24272,N_15356,N_15825);
nor U24273 (N_24273,N_15596,N_16354);
nand U24274 (N_24274,N_15936,N_19089);
xor U24275 (N_24275,N_15214,N_19219);
xnor U24276 (N_24276,N_19233,N_16418);
nor U24277 (N_24277,N_15174,N_15799);
nand U24278 (N_24278,N_18274,N_16867);
xnor U24279 (N_24279,N_15548,N_16458);
or U24280 (N_24280,N_16784,N_18463);
or U24281 (N_24281,N_19203,N_18833);
and U24282 (N_24282,N_18869,N_18671);
nand U24283 (N_24283,N_18781,N_15605);
and U24284 (N_24284,N_17874,N_16352);
xnor U24285 (N_24285,N_17846,N_18294);
xnor U24286 (N_24286,N_16545,N_18739);
or U24287 (N_24287,N_16365,N_16571);
nor U24288 (N_24288,N_17430,N_17266);
nand U24289 (N_24289,N_17904,N_16627);
and U24290 (N_24290,N_18329,N_16885);
nor U24291 (N_24291,N_19264,N_15639);
nand U24292 (N_24292,N_17663,N_16677);
xnor U24293 (N_24293,N_19903,N_17938);
nand U24294 (N_24294,N_18701,N_17215);
nor U24295 (N_24295,N_15017,N_16368);
or U24296 (N_24296,N_17308,N_18391);
nor U24297 (N_24297,N_15423,N_15210);
nand U24298 (N_24298,N_19323,N_17606);
or U24299 (N_24299,N_17738,N_18107);
and U24300 (N_24300,N_19702,N_19974);
xnor U24301 (N_24301,N_15664,N_18169);
and U24302 (N_24302,N_19002,N_19152);
or U24303 (N_24303,N_17188,N_18815);
xor U24304 (N_24304,N_15841,N_18059);
and U24305 (N_24305,N_15965,N_16332);
xnor U24306 (N_24306,N_15676,N_17323);
and U24307 (N_24307,N_17542,N_17076);
and U24308 (N_24308,N_17164,N_19205);
nor U24309 (N_24309,N_18019,N_15873);
or U24310 (N_24310,N_19632,N_18400);
nor U24311 (N_24311,N_18019,N_18095);
nand U24312 (N_24312,N_17255,N_19146);
nand U24313 (N_24313,N_15964,N_18031);
or U24314 (N_24314,N_17994,N_17123);
xor U24315 (N_24315,N_16908,N_19253);
and U24316 (N_24316,N_17568,N_17726);
nor U24317 (N_24317,N_15748,N_15379);
or U24318 (N_24318,N_15702,N_17557);
and U24319 (N_24319,N_15586,N_15045);
or U24320 (N_24320,N_18966,N_16648);
and U24321 (N_24321,N_19369,N_15471);
or U24322 (N_24322,N_18611,N_17615);
xnor U24323 (N_24323,N_16431,N_18547);
xor U24324 (N_24324,N_15507,N_17607);
xor U24325 (N_24325,N_16191,N_19571);
nand U24326 (N_24326,N_19539,N_15244);
and U24327 (N_24327,N_18675,N_19801);
nor U24328 (N_24328,N_16858,N_19814);
nor U24329 (N_24329,N_18607,N_19648);
xor U24330 (N_24330,N_18092,N_16885);
nand U24331 (N_24331,N_16306,N_19642);
or U24332 (N_24332,N_15394,N_18244);
xnor U24333 (N_24333,N_15301,N_17546);
xnor U24334 (N_24334,N_18487,N_19649);
nand U24335 (N_24335,N_16558,N_18159);
and U24336 (N_24336,N_17431,N_16636);
or U24337 (N_24337,N_18580,N_19997);
and U24338 (N_24338,N_18838,N_17796);
nor U24339 (N_24339,N_16587,N_17873);
and U24340 (N_24340,N_16513,N_16540);
or U24341 (N_24341,N_19712,N_15591);
or U24342 (N_24342,N_17783,N_19358);
nand U24343 (N_24343,N_15523,N_18494);
or U24344 (N_24344,N_18926,N_17832);
xnor U24345 (N_24345,N_15725,N_18391);
and U24346 (N_24346,N_17185,N_19534);
nand U24347 (N_24347,N_19769,N_15394);
nor U24348 (N_24348,N_15068,N_18260);
and U24349 (N_24349,N_16152,N_19130);
nor U24350 (N_24350,N_15057,N_15295);
nand U24351 (N_24351,N_16917,N_16316);
nor U24352 (N_24352,N_17978,N_18066);
xor U24353 (N_24353,N_15057,N_19543);
xor U24354 (N_24354,N_15837,N_16033);
or U24355 (N_24355,N_16584,N_17530);
and U24356 (N_24356,N_15692,N_16659);
nor U24357 (N_24357,N_18764,N_19060);
and U24358 (N_24358,N_17993,N_18015);
nor U24359 (N_24359,N_19031,N_16944);
xnor U24360 (N_24360,N_18279,N_17804);
and U24361 (N_24361,N_16897,N_16423);
or U24362 (N_24362,N_18113,N_16581);
nor U24363 (N_24363,N_16195,N_18675);
nand U24364 (N_24364,N_18549,N_18798);
and U24365 (N_24365,N_17720,N_18502);
nand U24366 (N_24366,N_15897,N_19778);
and U24367 (N_24367,N_19017,N_16551);
nand U24368 (N_24368,N_16707,N_16016);
or U24369 (N_24369,N_19747,N_18125);
or U24370 (N_24370,N_16655,N_19053);
nor U24371 (N_24371,N_16033,N_16501);
or U24372 (N_24372,N_15691,N_18571);
or U24373 (N_24373,N_16860,N_19848);
xor U24374 (N_24374,N_16567,N_18292);
or U24375 (N_24375,N_18450,N_15661);
or U24376 (N_24376,N_18150,N_16679);
nand U24377 (N_24377,N_17847,N_15174);
xor U24378 (N_24378,N_18000,N_18251);
nor U24379 (N_24379,N_15278,N_19957);
nand U24380 (N_24380,N_19557,N_15874);
and U24381 (N_24381,N_17932,N_16348);
xnor U24382 (N_24382,N_17419,N_17520);
and U24383 (N_24383,N_18276,N_17274);
nor U24384 (N_24384,N_15618,N_15423);
or U24385 (N_24385,N_15643,N_17780);
nand U24386 (N_24386,N_15552,N_16469);
xnor U24387 (N_24387,N_19282,N_19753);
and U24388 (N_24388,N_15201,N_18047);
or U24389 (N_24389,N_19305,N_18543);
or U24390 (N_24390,N_15074,N_18730);
nand U24391 (N_24391,N_15176,N_17526);
or U24392 (N_24392,N_17181,N_17396);
nor U24393 (N_24393,N_17267,N_19845);
nor U24394 (N_24394,N_15914,N_15002);
or U24395 (N_24395,N_16712,N_19450);
and U24396 (N_24396,N_18951,N_16905);
xnor U24397 (N_24397,N_19234,N_15285);
or U24398 (N_24398,N_17962,N_15013);
nand U24399 (N_24399,N_18171,N_19862);
xnor U24400 (N_24400,N_19742,N_17884);
nor U24401 (N_24401,N_15457,N_19335);
nand U24402 (N_24402,N_15749,N_18043);
nand U24403 (N_24403,N_17257,N_18818);
or U24404 (N_24404,N_19010,N_15750);
nand U24405 (N_24405,N_16890,N_16058);
and U24406 (N_24406,N_18964,N_18795);
or U24407 (N_24407,N_18011,N_16774);
xnor U24408 (N_24408,N_16929,N_17072);
nor U24409 (N_24409,N_18294,N_16659);
nor U24410 (N_24410,N_18270,N_17917);
and U24411 (N_24411,N_16675,N_17828);
and U24412 (N_24412,N_19247,N_17860);
or U24413 (N_24413,N_17230,N_17079);
nor U24414 (N_24414,N_17336,N_15735);
nand U24415 (N_24415,N_19735,N_19402);
xor U24416 (N_24416,N_17262,N_15336);
nand U24417 (N_24417,N_18532,N_15921);
and U24418 (N_24418,N_17997,N_16222);
nand U24419 (N_24419,N_18906,N_16842);
xnor U24420 (N_24420,N_15559,N_19007);
and U24421 (N_24421,N_17815,N_18377);
nor U24422 (N_24422,N_15281,N_17424);
or U24423 (N_24423,N_16441,N_16078);
nand U24424 (N_24424,N_19856,N_16639);
and U24425 (N_24425,N_15072,N_18042);
nand U24426 (N_24426,N_19918,N_19144);
xor U24427 (N_24427,N_18269,N_16743);
xor U24428 (N_24428,N_19738,N_16043);
nand U24429 (N_24429,N_16467,N_18791);
xnor U24430 (N_24430,N_15641,N_15126);
nand U24431 (N_24431,N_18062,N_16696);
nor U24432 (N_24432,N_18425,N_17169);
nor U24433 (N_24433,N_15768,N_18095);
xor U24434 (N_24434,N_15853,N_17176);
nand U24435 (N_24435,N_16363,N_19057);
and U24436 (N_24436,N_18410,N_17690);
and U24437 (N_24437,N_16498,N_16234);
nand U24438 (N_24438,N_17929,N_15780);
nor U24439 (N_24439,N_19508,N_16361);
xnor U24440 (N_24440,N_18722,N_17081);
nand U24441 (N_24441,N_19677,N_18388);
xnor U24442 (N_24442,N_19962,N_17084);
nand U24443 (N_24443,N_19560,N_17035);
nor U24444 (N_24444,N_16792,N_15007);
and U24445 (N_24445,N_15995,N_17849);
and U24446 (N_24446,N_19878,N_15125);
and U24447 (N_24447,N_17448,N_19056);
nor U24448 (N_24448,N_19000,N_19661);
xnor U24449 (N_24449,N_15065,N_19152);
xor U24450 (N_24450,N_18532,N_18370);
xor U24451 (N_24451,N_19583,N_16090);
xor U24452 (N_24452,N_17202,N_19882);
xnor U24453 (N_24453,N_19693,N_18835);
nor U24454 (N_24454,N_19698,N_16258);
or U24455 (N_24455,N_18754,N_16130);
nor U24456 (N_24456,N_15841,N_16733);
or U24457 (N_24457,N_16952,N_19684);
nor U24458 (N_24458,N_15934,N_16280);
or U24459 (N_24459,N_18497,N_17351);
or U24460 (N_24460,N_18634,N_16168);
or U24461 (N_24461,N_18474,N_19782);
nand U24462 (N_24462,N_18015,N_19347);
or U24463 (N_24463,N_19880,N_15545);
or U24464 (N_24464,N_19262,N_17777);
or U24465 (N_24465,N_18883,N_18403);
nand U24466 (N_24466,N_18711,N_18297);
and U24467 (N_24467,N_17015,N_17947);
xor U24468 (N_24468,N_18968,N_15496);
or U24469 (N_24469,N_16706,N_15427);
nor U24470 (N_24470,N_18991,N_17126);
nand U24471 (N_24471,N_15089,N_19197);
or U24472 (N_24472,N_19330,N_18504);
or U24473 (N_24473,N_16363,N_19697);
nand U24474 (N_24474,N_19774,N_18771);
xnor U24475 (N_24475,N_15840,N_15575);
nand U24476 (N_24476,N_19487,N_15633);
and U24477 (N_24477,N_15787,N_19726);
or U24478 (N_24478,N_19618,N_19163);
or U24479 (N_24479,N_15610,N_15191);
xnor U24480 (N_24480,N_18083,N_15309);
or U24481 (N_24481,N_16569,N_15745);
nand U24482 (N_24482,N_16946,N_17837);
and U24483 (N_24483,N_19741,N_18681);
nand U24484 (N_24484,N_17698,N_17460);
nand U24485 (N_24485,N_17219,N_17385);
xor U24486 (N_24486,N_15603,N_16127);
or U24487 (N_24487,N_15585,N_15553);
and U24488 (N_24488,N_16060,N_15280);
nand U24489 (N_24489,N_19144,N_19207);
nor U24490 (N_24490,N_19628,N_16594);
xnor U24491 (N_24491,N_17546,N_16382);
or U24492 (N_24492,N_19744,N_15222);
nor U24493 (N_24493,N_19316,N_16140);
or U24494 (N_24494,N_15167,N_17858);
xor U24495 (N_24495,N_16668,N_15860);
and U24496 (N_24496,N_18704,N_19025);
xnor U24497 (N_24497,N_18827,N_18188);
and U24498 (N_24498,N_16605,N_18165);
nor U24499 (N_24499,N_18471,N_18784);
or U24500 (N_24500,N_16937,N_15403);
xor U24501 (N_24501,N_17662,N_18297);
nand U24502 (N_24502,N_17525,N_19440);
xnor U24503 (N_24503,N_18622,N_16922);
nor U24504 (N_24504,N_18612,N_18988);
nor U24505 (N_24505,N_16498,N_17199);
and U24506 (N_24506,N_19306,N_17213);
xnor U24507 (N_24507,N_15387,N_19955);
xnor U24508 (N_24508,N_18347,N_16458);
or U24509 (N_24509,N_19259,N_16366);
or U24510 (N_24510,N_18954,N_16037);
nand U24511 (N_24511,N_19675,N_17365);
and U24512 (N_24512,N_16445,N_17959);
nand U24513 (N_24513,N_18385,N_19677);
nor U24514 (N_24514,N_18561,N_19555);
nor U24515 (N_24515,N_18279,N_18793);
nand U24516 (N_24516,N_15498,N_19326);
xnor U24517 (N_24517,N_18830,N_15354);
and U24518 (N_24518,N_19078,N_16861);
nor U24519 (N_24519,N_15171,N_17102);
nand U24520 (N_24520,N_16286,N_15873);
nand U24521 (N_24521,N_15279,N_16450);
xor U24522 (N_24522,N_15551,N_19078);
or U24523 (N_24523,N_18736,N_15283);
nand U24524 (N_24524,N_17701,N_15038);
or U24525 (N_24525,N_16791,N_19537);
xor U24526 (N_24526,N_15846,N_15013);
nor U24527 (N_24527,N_19045,N_19957);
or U24528 (N_24528,N_18183,N_16620);
and U24529 (N_24529,N_18892,N_15465);
nor U24530 (N_24530,N_17104,N_17324);
xor U24531 (N_24531,N_19333,N_15935);
and U24532 (N_24532,N_16135,N_19919);
nand U24533 (N_24533,N_17663,N_17817);
or U24534 (N_24534,N_17885,N_17983);
xor U24535 (N_24535,N_17611,N_16287);
nand U24536 (N_24536,N_16940,N_15387);
nand U24537 (N_24537,N_15104,N_17226);
xor U24538 (N_24538,N_15334,N_16859);
or U24539 (N_24539,N_15205,N_15841);
nand U24540 (N_24540,N_16538,N_19664);
nor U24541 (N_24541,N_19714,N_17380);
nand U24542 (N_24542,N_17441,N_15315);
xor U24543 (N_24543,N_18156,N_15696);
nor U24544 (N_24544,N_18446,N_16862);
nor U24545 (N_24545,N_18367,N_19527);
xnor U24546 (N_24546,N_18166,N_15663);
nor U24547 (N_24547,N_15422,N_19473);
nand U24548 (N_24548,N_15042,N_18848);
and U24549 (N_24549,N_17014,N_15084);
or U24550 (N_24550,N_18590,N_17522);
nand U24551 (N_24551,N_18064,N_17270);
or U24552 (N_24552,N_15420,N_19773);
nand U24553 (N_24553,N_19876,N_15156);
xnor U24554 (N_24554,N_16774,N_19372);
nand U24555 (N_24555,N_17611,N_18993);
or U24556 (N_24556,N_18057,N_15689);
nand U24557 (N_24557,N_16437,N_15239);
or U24558 (N_24558,N_15822,N_18793);
and U24559 (N_24559,N_16842,N_17172);
nor U24560 (N_24560,N_19396,N_15143);
xnor U24561 (N_24561,N_16178,N_18858);
xor U24562 (N_24562,N_16582,N_16759);
xor U24563 (N_24563,N_15498,N_17759);
nor U24564 (N_24564,N_19581,N_15481);
xnor U24565 (N_24565,N_17568,N_15197);
xor U24566 (N_24566,N_16196,N_19200);
and U24567 (N_24567,N_16973,N_19825);
xnor U24568 (N_24568,N_16355,N_15442);
nand U24569 (N_24569,N_17186,N_19359);
or U24570 (N_24570,N_15879,N_15896);
nor U24571 (N_24571,N_15227,N_17726);
xnor U24572 (N_24572,N_17475,N_15301);
nor U24573 (N_24573,N_17173,N_19826);
and U24574 (N_24574,N_18029,N_16869);
and U24575 (N_24575,N_18374,N_19035);
xnor U24576 (N_24576,N_17319,N_16232);
xor U24577 (N_24577,N_15343,N_17433);
nor U24578 (N_24578,N_19704,N_19556);
nor U24579 (N_24579,N_19748,N_15568);
or U24580 (N_24580,N_19257,N_16134);
nor U24581 (N_24581,N_17442,N_18020);
nand U24582 (N_24582,N_15704,N_18723);
xnor U24583 (N_24583,N_17634,N_19845);
xor U24584 (N_24584,N_18446,N_17134);
xor U24585 (N_24585,N_15994,N_19917);
nand U24586 (N_24586,N_17168,N_15378);
nand U24587 (N_24587,N_18914,N_16499);
xnor U24588 (N_24588,N_18967,N_15710);
xor U24589 (N_24589,N_19668,N_16712);
xnor U24590 (N_24590,N_15438,N_16931);
nor U24591 (N_24591,N_19638,N_15204);
nor U24592 (N_24592,N_16452,N_17264);
nand U24593 (N_24593,N_17058,N_16547);
nand U24594 (N_24594,N_17153,N_19071);
and U24595 (N_24595,N_18287,N_15164);
nand U24596 (N_24596,N_17773,N_18731);
and U24597 (N_24597,N_18281,N_15273);
or U24598 (N_24598,N_17138,N_16682);
nand U24599 (N_24599,N_19335,N_18015);
and U24600 (N_24600,N_15319,N_19450);
xnor U24601 (N_24601,N_17898,N_17180);
and U24602 (N_24602,N_16179,N_15520);
xnor U24603 (N_24603,N_18733,N_19446);
nand U24604 (N_24604,N_15396,N_16769);
nor U24605 (N_24605,N_19146,N_15525);
nand U24606 (N_24606,N_15395,N_18822);
and U24607 (N_24607,N_17813,N_19595);
or U24608 (N_24608,N_19540,N_17176);
and U24609 (N_24609,N_19995,N_18953);
xor U24610 (N_24610,N_16939,N_16836);
xnor U24611 (N_24611,N_17695,N_18639);
nor U24612 (N_24612,N_17325,N_15216);
xor U24613 (N_24613,N_17881,N_15481);
nor U24614 (N_24614,N_15799,N_17002);
nand U24615 (N_24615,N_18077,N_15479);
or U24616 (N_24616,N_17081,N_17713);
xnor U24617 (N_24617,N_18700,N_19604);
nand U24618 (N_24618,N_15281,N_19313);
and U24619 (N_24619,N_16758,N_18916);
and U24620 (N_24620,N_17499,N_18420);
nand U24621 (N_24621,N_17742,N_19610);
nor U24622 (N_24622,N_18285,N_16272);
and U24623 (N_24623,N_19284,N_16966);
and U24624 (N_24624,N_15637,N_15737);
xor U24625 (N_24625,N_18750,N_15388);
nand U24626 (N_24626,N_19055,N_18576);
nor U24627 (N_24627,N_17646,N_17498);
nand U24628 (N_24628,N_15061,N_15741);
xor U24629 (N_24629,N_19789,N_18471);
or U24630 (N_24630,N_19043,N_18317);
and U24631 (N_24631,N_16239,N_19207);
nor U24632 (N_24632,N_16502,N_15234);
nand U24633 (N_24633,N_18873,N_18144);
nor U24634 (N_24634,N_19693,N_19305);
nand U24635 (N_24635,N_19446,N_17314);
or U24636 (N_24636,N_18670,N_16336);
nand U24637 (N_24637,N_17397,N_16741);
or U24638 (N_24638,N_18010,N_19394);
and U24639 (N_24639,N_18440,N_16200);
nand U24640 (N_24640,N_17602,N_17357);
nor U24641 (N_24641,N_18956,N_16644);
xnor U24642 (N_24642,N_15497,N_19808);
xnor U24643 (N_24643,N_16251,N_16726);
and U24644 (N_24644,N_16726,N_18220);
nand U24645 (N_24645,N_15171,N_16065);
xor U24646 (N_24646,N_19674,N_17102);
nand U24647 (N_24647,N_18145,N_15068);
nor U24648 (N_24648,N_16092,N_18939);
or U24649 (N_24649,N_17410,N_18848);
nand U24650 (N_24650,N_16229,N_17257);
nand U24651 (N_24651,N_16135,N_15058);
nand U24652 (N_24652,N_16454,N_19684);
or U24653 (N_24653,N_18270,N_15274);
nand U24654 (N_24654,N_15977,N_15809);
xnor U24655 (N_24655,N_16746,N_17814);
and U24656 (N_24656,N_17007,N_15342);
or U24657 (N_24657,N_17037,N_16098);
or U24658 (N_24658,N_19047,N_16071);
nand U24659 (N_24659,N_17640,N_15443);
nor U24660 (N_24660,N_16324,N_18025);
nor U24661 (N_24661,N_18699,N_16841);
xor U24662 (N_24662,N_16813,N_16664);
xnor U24663 (N_24663,N_15170,N_18672);
xor U24664 (N_24664,N_19075,N_18783);
and U24665 (N_24665,N_19009,N_16356);
nand U24666 (N_24666,N_18144,N_19553);
xor U24667 (N_24667,N_16238,N_16242);
and U24668 (N_24668,N_16215,N_19386);
xor U24669 (N_24669,N_16880,N_18573);
or U24670 (N_24670,N_18782,N_16737);
nor U24671 (N_24671,N_17479,N_17309);
or U24672 (N_24672,N_15663,N_19597);
and U24673 (N_24673,N_17857,N_18798);
xnor U24674 (N_24674,N_17540,N_18593);
xor U24675 (N_24675,N_17216,N_17343);
nor U24676 (N_24676,N_19220,N_18529);
xor U24677 (N_24677,N_15957,N_15419);
and U24678 (N_24678,N_17825,N_16209);
nand U24679 (N_24679,N_17640,N_15417);
nand U24680 (N_24680,N_18283,N_18657);
nor U24681 (N_24681,N_15235,N_18967);
or U24682 (N_24682,N_16837,N_18192);
nand U24683 (N_24683,N_18580,N_18230);
or U24684 (N_24684,N_17957,N_15077);
xnor U24685 (N_24685,N_19723,N_16894);
or U24686 (N_24686,N_18792,N_19143);
xor U24687 (N_24687,N_17736,N_15200);
or U24688 (N_24688,N_19792,N_18819);
and U24689 (N_24689,N_16367,N_16837);
nor U24690 (N_24690,N_16187,N_17618);
and U24691 (N_24691,N_18657,N_16418);
and U24692 (N_24692,N_16595,N_15648);
xor U24693 (N_24693,N_18518,N_15890);
xnor U24694 (N_24694,N_16611,N_16810);
nor U24695 (N_24695,N_15877,N_19794);
and U24696 (N_24696,N_19621,N_16848);
nand U24697 (N_24697,N_16353,N_18071);
and U24698 (N_24698,N_19501,N_15922);
xnor U24699 (N_24699,N_18206,N_17945);
nand U24700 (N_24700,N_19198,N_15369);
and U24701 (N_24701,N_17044,N_19452);
nor U24702 (N_24702,N_16437,N_18239);
and U24703 (N_24703,N_15884,N_19395);
or U24704 (N_24704,N_16800,N_15376);
and U24705 (N_24705,N_15636,N_15455);
xnor U24706 (N_24706,N_17385,N_17843);
or U24707 (N_24707,N_15835,N_19229);
nor U24708 (N_24708,N_15245,N_19411);
nand U24709 (N_24709,N_19977,N_19281);
nand U24710 (N_24710,N_17518,N_16292);
or U24711 (N_24711,N_18032,N_15821);
or U24712 (N_24712,N_18026,N_15765);
xor U24713 (N_24713,N_18813,N_18589);
nand U24714 (N_24714,N_15950,N_16701);
or U24715 (N_24715,N_15358,N_19335);
xor U24716 (N_24716,N_16075,N_18356);
nand U24717 (N_24717,N_17697,N_16617);
or U24718 (N_24718,N_16902,N_19996);
and U24719 (N_24719,N_16686,N_15092);
or U24720 (N_24720,N_19227,N_19111);
nor U24721 (N_24721,N_19346,N_15899);
xnor U24722 (N_24722,N_16584,N_19386);
nand U24723 (N_24723,N_15266,N_19878);
or U24724 (N_24724,N_18141,N_18666);
nor U24725 (N_24725,N_18131,N_18837);
and U24726 (N_24726,N_16031,N_16155);
nor U24727 (N_24727,N_17097,N_15338);
nand U24728 (N_24728,N_18199,N_17206);
xnor U24729 (N_24729,N_16481,N_18193);
xor U24730 (N_24730,N_19259,N_17130);
or U24731 (N_24731,N_18950,N_19349);
nor U24732 (N_24732,N_19242,N_18665);
nor U24733 (N_24733,N_17048,N_18563);
nand U24734 (N_24734,N_17372,N_15573);
nor U24735 (N_24735,N_19257,N_17141);
and U24736 (N_24736,N_19340,N_16305);
nor U24737 (N_24737,N_15631,N_16882);
and U24738 (N_24738,N_17832,N_18961);
and U24739 (N_24739,N_17776,N_17591);
nor U24740 (N_24740,N_19906,N_15526);
xor U24741 (N_24741,N_19553,N_16274);
nor U24742 (N_24742,N_17817,N_17131);
and U24743 (N_24743,N_16874,N_17450);
nor U24744 (N_24744,N_17628,N_18878);
or U24745 (N_24745,N_15944,N_16900);
and U24746 (N_24746,N_19000,N_16236);
nand U24747 (N_24747,N_15038,N_15721);
xnor U24748 (N_24748,N_17384,N_16279);
nand U24749 (N_24749,N_16699,N_18798);
nand U24750 (N_24750,N_19597,N_16642);
nand U24751 (N_24751,N_16984,N_15795);
nor U24752 (N_24752,N_17864,N_16391);
or U24753 (N_24753,N_19663,N_19817);
and U24754 (N_24754,N_16736,N_15616);
or U24755 (N_24755,N_15046,N_15820);
xnor U24756 (N_24756,N_18245,N_16485);
or U24757 (N_24757,N_15426,N_18753);
or U24758 (N_24758,N_15470,N_16599);
nand U24759 (N_24759,N_19987,N_17325);
or U24760 (N_24760,N_15871,N_19979);
xnor U24761 (N_24761,N_18207,N_19560);
xnor U24762 (N_24762,N_19086,N_16518);
xor U24763 (N_24763,N_17768,N_16759);
nand U24764 (N_24764,N_15634,N_15238);
and U24765 (N_24765,N_19351,N_15259);
xor U24766 (N_24766,N_16893,N_16013);
and U24767 (N_24767,N_15013,N_19184);
nor U24768 (N_24768,N_15378,N_16776);
nor U24769 (N_24769,N_16803,N_18502);
nand U24770 (N_24770,N_17591,N_15330);
nor U24771 (N_24771,N_16021,N_18387);
or U24772 (N_24772,N_15780,N_17158);
or U24773 (N_24773,N_17928,N_18288);
nor U24774 (N_24774,N_18224,N_16632);
and U24775 (N_24775,N_16421,N_19625);
nand U24776 (N_24776,N_19258,N_15856);
and U24777 (N_24777,N_18162,N_16317);
and U24778 (N_24778,N_15980,N_16068);
nor U24779 (N_24779,N_18911,N_18249);
nand U24780 (N_24780,N_19905,N_15121);
and U24781 (N_24781,N_19432,N_18635);
xor U24782 (N_24782,N_19613,N_15628);
and U24783 (N_24783,N_16142,N_18947);
nor U24784 (N_24784,N_16179,N_17173);
and U24785 (N_24785,N_19967,N_16392);
xnor U24786 (N_24786,N_16081,N_16758);
nand U24787 (N_24787,N_19976,N_15391);
and U24788 (N_24788,N_19766,N_18741);
nand U24789 (N_24789,N_15290,N_19556);
nor U24790 (N_24790,N_16347,N_18912);
and U24791 (N_24791,N_17065,N_19252);
xnor U24792 (N_24792,N_15267,N_18331);
and U24793 (N_24793,N_18793,N_15993);
xnor U24794 (N_24794,N_18350,N_15360);
nor U24795 (N_24795,N_19709,N_15926);
or U24796 (N_24796,N_18505,N_17653);
nand U24797 (N_24797,N_15232,N_18419);
and U24798 (N_24798,N_17952,N_16533);
nor U24799 (N_24799,N_17207,N_18116);
nand U24800 (N_24800,N_15449,N_17728);
or U24801 (N_24801,N_18674,N_17759);
or U24802 (N_24802,N_17340,N_17033);
nor U24803 (N_24803,N_19813,N_17625);
xnor U24804 (N_24804,N_19696,N_16092);
xnor U24805 (N_24805,N_17329,N_17409);
xor U24806 (N_24806,N_17320,N_16110);
nor U24807 (N_24807,N_17742,N_17459);
xor U24808 (N_24808,N_17247,N_18841);
xnor U24809 (N_24809,N_16830,N_18150);
or U24810 (N_24810,N_15137,N_15277);
xnor U24811 (N_24811,N_19026,N_15327);
nor U24812 (N_24812,N_16316,N_15378);
or U24813 (N_24813,N_17426,N_15557);
xor U24814 (N_24814,N_15235,N_18694);
or U24815 (N_24815,N_17815,N_17643);
or U24816 (N_24816,N_18027,N_19336);
nor U24817 (N_24817,N_16607,N_18960);
nand U24818 (N_24818,N_19830,N_15526);
nand U24819 (N_24819,N_18831,N_19918);
nand U24820 (N_24820,N_16056,N_17769);
nand U24821 (N_24821,N_19457,N_18653);
nor U24822 (N_24822,N_15087,N_16910);
xnor U24823 (N_24823,N_17961,N_18428);
nor U24824 (N_24824,N_18056,N_18978);
nor U24825 (N_24825,N_15550,N_16865);
nor U24826 (N_24826,N_17003,N_19470);
and U24827 (N_24827,N_19392,N_15531);
nand U24828 (N_24828,N_18558,N_16356);
nor U24829 (N_24829,N_16778,N_16115);
or U24830 (N_24830,N_15487,N_15678);
and U24831 (N_24831,N_16964,N_16777);
or U24832 (N_24832,N_19780,N_15612);
and U24833 (N_24833,N_16855,N_19438);
nor U24834 (N_24834,N_19797,N_15317);
or U24835 (N_24835,N_18306,N_16407);
or U24836 (N_24836,N_16567,N_19750);
and U24837 (N_24837,N_16639,N_15752);
nand U24838 (N_24838,N_19214,N_18851);
or U24839 (N_24839,N_17925,N_16680);
nor U24840 (N_24840,N_16458,N_17136);
and U24841 (N_24841,N_16371,N_18098);
or U24842 (N_24842,N_19637,N_16549);
and U24843 (N_24843,N_18230,N_16843);
xor U24844 (N_24844,N_18428,N_16962);
and U24845 (N_24845,N_17993,N_17697);
and U24846 (N_24846,N_15126,N_18019);
xnor U24847 (N_24847,N_18775,N_18499);
or U24848 (N_24848,N_19012,N_18347);
or U24849 (N_24849,N_19657,N_16653);
nor U24850 (N_24850,N_16312,N_18709);
nor U24851 (N_24851,N_15090,N_17809);
and U24852 (N_24852,N_18201,N_19771);
or U24853 (N_24853,N_19125,N_15793);
nand U24854 (N_24854,N_19075,N_16287);
and U24855 (N_24855,N_18348,N_16280);
nand U24856 (N_24856,N_16268,N_18030);
and U24857 (N_24857,N_19702,N_15352);
or U24858 (N_24858,N_17730,N_15532);
nand U24859 (N_24859,N_16019,N_18666);
nand U24860 (N_24860,N_19643,N_15172);
nand U24861 (N_24861,N_19706,N_15208);
and U24862 (N_24862,N_18294,N_15036);
nand U24863 (N_24863,N_15654,N_16527);
or U24864 (N_24864,N_18688,N_19345);
nand U24865 (N_24865,N_15037,N_16419);
and U24866 (N_24866,N_15089,N_17531);
nor U24867 (N_24867,N_17450,N_16763);
or U24868 (N_24868,N_17597,N_19554);
and U24869 (N_24869,N_17774,N_19699);
xor U24870 (N_24870,N_19753,N_18733);
or U24871 (N_24871,N_18384,N_19051);
nor U24872 (N_24872,N_19112,N_16325);
nand U24873 (N_24873,N_16270,N_16692);
nand U24874 (N_24874,N_16770,N_16211);
nand U24875 (N_24875,N_15890,N_17893);
nor U24876 (N_24876,N_16943,N_19538);
nor U24877 (N_24877,N_18867,N_17151);
nor U24878 (N_24878,N_15752,N_15511);
nor U24879 (N_24879,N_18722,N_18765);
xor U24880 (N_24880,N_15979,N_15059);
and U24881 (N_24881,N_19634,N_18425);
and U24882 (N_24882,N_18195,N_18727);
xnor U24883 (N_24883,N_18941,N_18299);
or U24884 (N_24884,N_15142,N_17624);
or U24885 (N_24885,N_16358,N_18396);
nand U24886 (N_24886,N_15151,N_18658);
nor U24887 (N_24887,N_16623,N_17431);
xnor U24888 (N_24888,N_16616,N_15111);
nand U24889 (N_24889,N_18175,N_19237);
nor U24890 (N_24890,N_18466,N_15310);
and U24891 (N_24891,N_19055,N_17581);
or U24892 (N_24892,N_16334,N_17559);
nor U24893 (N_24893,N_19527,N_17093);
nor U24894 (N_24894,N_16321,N_18335);
and U24895 (N_24895,N_17117,N_18308);
nand U24896 (N_24896,N_16608,N_16373);
and U24897 (N_24897,N_17326,N_16631);
nand U24898 (N_24898,N_15496,N_15466);
nand U24899 (N_24899,N_18297,N_19064);
or U24900 (N_24900,N_19795,N_19702);
xor U24901 (N_24901,N_16772,N_15959);
xnor U24902 (N_24902,N_17065,N_17497);
and U24903 (N_24903,N_17088,N_15298);
xor U24904 (N_24904,N_19546,N_18402);
nand U24905 (N_24905,N_18477,N_19794);
xor U24906 (N_24906,N_18055,N_16097);
xnor U24907 (N_24907,N_16225,N_19040);
xor U24908 (N_24908,N_16132,N_19682);
nor U24909 (N_24909,N_16498,N_16998);
nand U24910 (N_24910,N_19253,N_18404);
and U24911 (N_24911,N_15098,N_19416);
nand U24912 (N_24912,N_17237,N_15495);
nand U24913 (N_24913,N_17875,N_17824);
and U24914 (N_24914,N_18715,N_18138);
xnor U24915 (N_24915,N_15683,N_18219);
and U24916 (N_24916,N_19766,N_17713);
nor U24917 (N_24917,N_15246,N_19226);
nand U24918 (N_24918,N_15252,N_19770);
or U24919 (N_24919,N_18438,N_19347);
xor U24920 (N_24920,N_15269,N_18186);
xor U24921 (N_24921,N_19207,N_17112);
nor U24922 (N_24922,N_18159,N_19967);
nor U24923 (N_24923,N_19387,N_16406);
nor U24924 (N_24924,N_16741,N_17587);
nand U24925 (N_24925,N_15178,N_18999);
nor U24926 (N_24926,N_15699,N_16929);
and U24927 (N_24927,N_16718,N_16262);
xnor U24928 (N_24928,N_17326,N_18456);
xor U24929 (N_24929,N_18784,N_15959);
and U24930 (N_24930,N_16837,N_15861);
or U24931 (N_24931,N_19035,N_15401);
and U24932 (N_24932,N_19110,N_18390);
nor U24933 (N_24933,N_16911,N_19268);
nor U24934 (N_24934,N_18704,N_15175);
nand U24935 (N_24935,N_19728,N_18283);
xnor U24936 (N_24936,N_17947,N_18308);
or U24937 (N_24937,N_17257,N_18361);
or U24938 (N_24938,N_16616,N_18248);
xor U24939 (N_24939,N_18166,N_16860);
nand U24940 (N_24940,N_19869,N_15181);
or U24941 (N_24941,N_19944,N_15176);
xor U24942 (N_24942,N_16986,N_19497);
xnor U24943 (N_24943,N_17487,N_18644);
nor U24944 (N_24944,N_16805,N_19033);
nor U24945 (N_24945,N_15932,N_15076);
nor U24946 (N_24946,N_19048,N_19385);
nand U24947 (N_24947,N_16816,N_15343);
xor U24948 (N_24948,N_16200,N_19797);
and U24949 (N_24949,N_19332,N_15458);
nand U24950 (N_24950,N_17862,N_17843);
nor U24951 (N_24951,N_19745,N_17810);
nand U24952 (N_24952,N_17920,N_17401);
and U24953 (N_24953,N_16343,N_15215);
nand U24954 (N_24954,N_16969,N_19716);
nand U24955 (N_24955,N_18163,N_17195);
or U24956 (N_24956,N_15991,N_15192);
and U24957 (N_24957,N_16183,N_17408);
xor U24958 (N_24958,N_16201,N_15323);
or U24959 (N_24959,N_19005,N_17820);
nor U24960 (N_24960,N_17302,N_17943);
and U24961 (N_24961,N_17553,N_18697);
xnor U24962 (N_24962,N_15378,N_17463);
nor U24963 (N_24963,N_16900,N_18238);
or U24964 (N_24964,N_16476,N_15269);
or U24965 (N_24965,N_19106,N_18195);
and U24966 (N_24966,N_18057,N_17548);
and U24967 (N_24967,N_19631,N_18773);
and U24968 (N_24968,N_19095,N_17599);
xor U24969 (N_24969,N_16402,N_19341);
nor U24970 (N_24970,N_16692,N_17133);
nor U24971 (N_24971,N_18515,N_18024);
nand U24972 (N_24972,N_17971,N_17114);
nor U24973 (N_24973,N_17658,N_18093);
and U24974 (N_24974,N_16683,N_17666);
and U24975 (N_24975,N_16614,N_18353);
and U24976 (N_24976,N_17316,N_15197);
and U24977 (N_24977,N_18616,N_18857);
nand U24978 (N_24978,N_19494,N_18911);
or U24979 (N_24979,N_17722,N_17815);
nand U24980 (N_24980,N_15206,N_17917);
xnor U24981 (N_24981,N_17319,N_16445);
nand U24982 (N_24982,N_18472,N_18265);
nor U24983 (N_24983,N_15600,N_19296);
nand U24984 (N_24984,N_17021,N_17328);
or U24985 (N_24985,N_18566,N_15765);
xor U24986 (N_24986,N_16334,N_17783);
nor U24987 (N_24987,N_18748,N_16716);
xnor U24988 (N_24988,N_16818,N_15589);
and U24989 (N_24989,N_17689,N_18381);
xnor U24990 (N_24990,N_16784,N_15809);
or U24991 (N_24991,N_17591,N_18318);
or U24992 (N_24992,N_16721,N_16569);
nor U24993 (N_24993,N_18855,N_16355);
and U24994 (N_24994,N_18050,N_19930);
nor U24995 (N_24995,N_19500,N_15716);
or U24996 (N_24996,N_18908,N_16510);
or U24997 (N_24997,N_16464,N_19085);
nand U24998 (N_24998,N_17176,N_19978);
and U24999 (N_24999,N_16512,N_15808);
xnor U25000 (N_25000,N_23929,N_21176);
nand U25001 (N_25001,N_24087,N_22633);
xnor U25002 (N_25002,N_22098,N_23247);
and U25003 (N_25003,N_23939,N_24893);
nand U25004 (N_25004,N_23759,N_20522);
nor U25005 (N_25005,N_23249,N_22999);
xor U25006 (N_25006,N_22447,N_24405);
or U25007 (N_25007,N_22785,N_24657);
nand U25008 (N_25008,N_22599,N_22404);
or U25009 (N_25009,N_24293,N_21877);
and U25010 (N_25010,N_20744,N_20113);
or U25011 (N_25011,N_22317,N_23331);
xor U25012 (N_25012,N_21283,N_20394);
or U25013 (N_25013,N_23550,N_20712);
or U25014 (N_25014,N_22102,N_20550);
and U25015 (N_25015,N_20591,N_22957);
nand U25016 (N_25016,N_24027,N_20554);
and U25017 (N_25017,N_22901,N_23298);
xnor U25018 (N_25018,N_20290,N_22644);
nand U25019 (N_25019,N_24997,N_24151);
and U25020 (N_25020,N_20806,N_20029);
nor U25021 (N_25021,N_23506,N_20224);
xnor U25022 (N_25022,N_23885,N_22530);
nor U25023 (N_25023,N_22402,N_21145);
and U25024 (N_25024,N_23496,N_21686);
xnor U25025 (N_25025,N_24472,N_21815);
xnor U25026 (N_25026,N_21329,N_22139);
and U25027 (N_25027,N_22024,N_23756);
nand U25028 (N_25028,N_21761,N_20539);
or U25029 (N_25029,N_21494,N_20731);
xnor U25030 (N_25030,N_24306,N_21078);
nand U25031 (N_25031,N_20455,N_22258);
nor U25032 (N_25032,N_23605,N_21959);
nor U25033 (N_25033,N_20634,N_20015);
and U25034 (N_25034,N_20312,N_23351);
xnor U25035 (N_25035,N_24240,N_20851);
nor U25036 (N_25036,N_22089,N_24917);
nor U25037 (N_25037,N_21270,N_23902);
nor U25038 (N_25038,N_20748,N_20449);
nor U25039 (N_25039,N_21546,N_24009);
nor U25040 (N_25040,N_21440,N_24316);
nor U25041 (N_25041,N_22656,N_24442);
and U25042 (N_25042,N_22699,N_23014);
nor U25043 (N_25043,N_24611,N_21096);
or U25044 (N_25044,N_24006,N_21169);
nand U25045 (N_25045,N_23648,N_24628);
or U25046 (N_25046,N_21294,N_24677);
or U25047 (N_25047,N_23676,N_21420);
and U25048 (N_25048,N_24062,N_23522);
nand U25049 (N_25049,N_22483,N_24666);
nor U25050 (N_25050,N_22923,N_22053);
nor U25051 (N_25051,N_21062,N_22032);
nand U25052 (N_25052,N_20509,N_22013);
or U25053 (N_25053,N_22109,N_20733);
xor U25054 (N_25054,N_21056,N_24169);
and U25055 (N_25055,N_24230,N_21637);
nor U25056 (N_25056,N_21499,N_24681);
nor U25057 (N_25057,N_22927,N_20054);
xnor U25058 (N_25058,N_20175,N_22141);
xnor U25059 (N_25059,N_20708,N_20264);
xor U25060 (N_25060,N_24511,N_24645);
or U25061 (N_25061,N_23115,N_24323);
xor U25062 (N_25062,N_24703,N_21852);
xor U25063 (N_25063,N_23056,N_20258);
nor U25064 (N_25064,N_22010,N_20407);
or U25065 (N_25065,N_24848,N_20494);
nand U25066 (N_25066,N_22216,N_24491);
nand U25067 (N_25067,N_24918,N_22496);
or U25068 (N_25068,N_23089,N_22261);
or U25069 (N_25069,N_20027,N_20391);
and U25070 (N_25070,N_22097,N_20686);
xnor U25071 (N_25071,N_23141,N_23256);
or U25072 (N_25072,N_23575,N_24107);
and U25073 (N_25073,N_24079,N_23576);
and U25074 (N_25074,N_24127,N_21951);
nand U25075 (N_25075,N_20935,N_22197);
and U25076 (N_25076,N_24742,N_21010);
xor U25077 (N_25077,N_24845,N_21006);
or U25078 (N_25078,N_23457,N_21766);
and U25079 (N_25079,N_20414,N_21895);
or U25080 (N_25080,N_24739,N_24732);
nor U25081 (N_25081,N_22045,N_22409);
xor U25082 (N_25082,N_21927,N_23895);
and U25083 (N_25083,N_22533,N_21591);
xor U25084 (N_25084,N_23454,N_22889);
and U25085 (N_25085,N_21059,N_20021);
nor U25086 (N_25086,N_23438,N_24969);
or U25087 (N_25087,N_22275,N_20001);
nand U25088 (N_25088,N_21736,N_20133);
or U25089 (N_25089,N_24250,N_24595);
or U25090 (N_25090,N_20805,N_22674);
or U25091 (N_25091,N_21476,N_20062);
xor U25092 (N_25092,N_24584,N_21029);
or U25093 (N_25093,N_22913,N_22757);
or U25094 (N_25094,N_20913,N_23326);
xor U25095 (N_25095,N_24721,N_20716);
nand U25096 (N_25096,N_22048,N_21525);
xor U25097 (N_25097,N_24229,N_24541);
xnor U25098 (N_25098,N_24867,N_21965);
or U25099 (N_25099,N_20372,N_24887);
and U25100 (N_25100,N_20431,N_22738);
and U25101 (N_25101,N_21847,N_22398);
and U25102 (N_25102,N_21986,N_23119);
or U25103 (N_25103,N_21336,N_21475);
and U25104 (N_25104,N_21653,N_20227);
nor U25105 (N_25105,N_24847,N_23928);
xnor U25106 (N_25106,N_24691,N_24105);
nor U25107 (N_25107,N_20259,N_21880);
and U25108 (N_25108,N_21694,N_24274);
xor U25109 (N_25109,N_21011,N_20102);
nor U25110 (N_25110,N_23931,N_23707);
and U25111 (N_25111,N_23938,N_21536);
nand U25112 (N_25112,N_20613,N_24227);
and U25113 (N_25113,N_21627,N_23007);
nand U25114 (N_25114,N_22778,N_23603);
and U25115 (N_25115,N_24746,N_23975);
nor U25116 (N_25116,N_20226,N_24618);
nor U25117 (N_25117,N_23746,N_21495);
nor U25118 (N_25118,N_24520,N_23234);
nor U25119 (N_25119,N_21679,N_22017);
xnor U25120 (N_25120,N_22969,N_21256);
and U25121 (N_25121,N_22801,N_24297);
xor U25122 (N_25122,N_22371,N_23560);
or U25123 (N_25123,N_21372,N_21121);
and U25124 (N_25124,N_21991,N_22745);
nor U25125 (N_25125,N_21043,N_24366);
or U25126 (N_25126,N_23003,N_20840);
or U25127 (N_25127,N_21930,N_20364);
nand U25128 (N_25128,N_23835,N_24299);
nand U25129 (N_25129,N_23842,N_21133);
xor U25130 (N_25130,N_24514,N_21837);
and U25131 (N_25131,N_21397,N_22176);
xnor U25132 (N_25132,N_23330,N_21483);
xnor U25133 (N_25133,N_24008,N_21517);
nand U25134 (N_25134,N_22948,N_21949);
and U25135 (N_25135,N_22982,N_23568);
nand U25136 (N_25136,N_20230,N_22046);
nand U25137 (N_25137,N_24815,N_21758);
and U25138 (N_25138,N_23161,N_20888);
nor U25139 (N_25139,N_24148,N_20490);
nor U25140 (N_25140,N_21723,N_21109);
nor U25141 (N_25141,N_21819,N_20602);
nor U25142 (N_25142,N_24115,N_23742);
xor U25143 (N_25143,N_20982,N_22967);
or U25144 (N_25144,N_24673,N_23536);
nand U25145 (N_25145,N_23060,N_20432);
nand U25146 (N_25146,N_23961,N_22627);
xnor U25147 (N_25147,N_21273,N_22219);
xor U25148 (N_25148,N_24271,N_23787);
nand U25149 (N_25149,N_21400,N_24425);
or U25150 (N_25150,N_21441,N_23292);
xor U25151 (N_25151,N_20501,N_21768);
nor U25152 (N_25152,N_24290,N_20667);
nor U25153 (N_25153,N_21197,N_22993);
xnor U25154 (N_25154,N_24521,N_21333);
nand U25155 (N_25155,N_20082,N_22320);
xnor U25156 (N_25156,N_24621,N_24857);
and U25157 (N_25157,N_22457,N_21613);
xor U25158 (N_25158,N_20864,N_20108);
nor U25159 (N_25159,N_20083,N_23586);
nand U25160 (N_25160,N_21269,N_24486);
nand U25161 (N_25161,N_20053,N_23205);
or U25162 (N_25162,N_21276,N_20039);
nor U25163 (N_25163,N_22857,N_24423);
nor U25164 (N_25164,N_24529,N_22846);
or U25165 (N_25165,N_23230,N_23433);
xor U25166 (N_25166,N_21136,N_23659);
xnor U25167 (N_25167,N_24586,N_22008);
and U25168 (N_25168,N_24363,N_24633);
nor U25169 (N_25169,N_21363,N_22207);
nor U25170 (N_25170,N_24463,N_24600);
nand U25171 (N_25171,N_23054,N_20237);
nand U25172 (N_25172,N_21080,N_23017);
and U25173 (N_25173,N_20361,N_21426);
xnor U25174 (N_25174,N_20477,N_23967);
or U25175 (N_25175,N_24589,N_22907);
xor U25176 (N_25176,N_23724,N_23564);
and U25177 (N_25177,N_22583,N_24559);
or U25178 (N_25178,N_24455,N_23156);
xnor U25179 (N_25179,N_21647,N_23263);
nor U25180 (N_25180,N_22077,N_23406);
xnor U25181 (N_25181,N_22694,N_21886);
and U25182 (N_25182,N_22463,N_24412);
nand U25183 (N_25183,N_20420,N_23591);
nand U25184 (N_25184,N_20110,N_21921);
and U25185 (N_25185,N_24723,N_22569);
nand U25186 (N_25186,N_23511,N_23758);
xor U25187 (N_25187,N_23739,N_20019);
or U25188 (N_25188,N_24434,N_22980);
xor U25189 (N_25189,N_24563,N_22511);
or U25190 (N_25190,N_23892,N_21322);
or U25191 (N_25191,N_21353,N_22874);
or U25192 (N_25192,N_24970,N_23136);
nand U25193 (N_25193,N_20183,N_22775);
and U25194 (N_25194,N_21784,N_23543);
nor U25195 (N_25195,N_22677,N_23268);
nor U25196 (N_25196,N_24640,N_23203);
and U25197 (N_25197,N_21009,N_21057);
xor U25198 (N_25198,N_21289,N_24740);
and U25199 (N_25199,N_20441,N_23019);
xnor U25200 (N_25200,N_20630,N_21069);
nand U25201 (N_25201,N_22971,N_20445);
xnor U25202 (N_25202,N_21326,N_22137);
nand U25203 (N_25203,N_21541,N_20886);
nand U25204 (N_25204,N_20808,N_20974);
xnor U25205 (N_25205,N_23529,N_21602);
nor U25206 (N_25206,N_21459,N_23012);
or U25207 (N_25207,N_23872,N_24489);
or U25208 (N_25208,N_24116,N_24095);
or U25209 (N_25209,N_20486,N_20485);
xor U25210 (N_25210,N_23376,N_24838);
and U25211 (N_25211,N_24136,N_22099);
and U25212 (N_25212,N_22337,N_23647);
nor U25213 (N_25213,N_24038,N_23020);
xnor U25214 (N_25214,N_20474,N_21045);
or U25215 (N_25215,N_24987,N_23080);
or U25216 (N_25216,N_22940,N_24710);
xor U25217 (N_25217,N_24462,N_20067);
or U25218 (N_25218,N_21449,N_24468);
nor U25219 (N_25219,N_20997,N_22461);
and U25220 (N_25220,N_24764,N_23688);
xnor U25221 (N_25221,N_20696,N_23004);
nor U25222 (N_25222,N_22895,N_20355);
and U25223 (N_25223,N_23366,N_24971);
nor U25224 (N_25224,N_24243,N_23635);
and U25225 (N_25225,N_22189,N_20729);
nor U25226 (N_25226,N_20127,N_24558);
nand U25227 (N_25227,N_24490,N_21733);
and U25228 (N_25228,N_23195,N_24421);
and U25229 (N_25229,N_24817,N_24142);
nor U25230 (N_25230,N_22848,N_24149);
xor U25231 (N_25231,N_21091,N_21415);
nand U25232 (N_25232,N_20637,N_23152);
nand U25233 (N_25233,N_24004,N_24916);
nor U25234 (N_25234,N_21926,N_23436);
or U25235 (N_25235,N_20567,N_21649);
nand U25236 (N_25236,N_24736,N_23941);
nand U25237 (N_25237,N_24449,N_21047);
nand U25238 (N_25238,N_20827,N_21140);
and U25239 (N_25239,N_20625,N_23159);
nand U25240 (N_25240,N_24317,N_24818);
xor U25241 (N_25241,N_22288,N_22826);
or U25242 (N_25242,N_23548,N_20581);
and U25243 (N_25243,N_23915,N_20291);
and U25244 (N_25244,N_20471,N_22472);
nor U25245 (N_25245,N_23018,N_23657);
nor U25246 (N_25246,N_23927,N_23876);
or U25247 (N_25247,N_24076,N_24548);
nand U25248 (N_25248,N_24846,N_23969);
and U25249 (N_25249,N_20203,N_24292);
nor U25250 (N_25250,N_23949,N_23528);
xor U25251 (N_25251,N_22921,N_23907);
and U25252 (N_25252,N_21493,N_22213);
and U25253 (N_25253,N_22296,N_21755);
nor U25254 (N_25254,N_21938,N_23871);
and U25255 (N_25255,N_22661,N_20294);
or U25256 (N_25256,N_21302,N_24877);
nor U25257 (N_25257,N_21244,N_20106);
or U25258 (N_25258,N_21825,N_20908);
nand U25259 (N_25259,N_22366,N_20545);
or U25260 (N_25260,N_20919,N_21317);
nor U25261 (N_25261,N_23899,N_21143);
xor U25262 (N_25262,N_20762,N_21100);
or U25263 (N_25263,N_23840,N_23533);
or U25264 (N_25264,N_24033,N_23449);
xor U25265 (N_25265,N_24061,N_22196);
or U25266 (N_25266,N_24789,N_20159);
xnor U25267 (N_25267,N_22932,N_24480);
xnor U25268 (N_25268,N_24594,N_23180);
nor U25269 (N_25269,N_20723,N_22323);
nand U25270 (N_25270,N_20789,N_23801);
nand U25271 (N_25271,N_22349,N_22410);
nand U25272 (N_25272,N_21841,N_21490);
or U25273 (N_25273,N_20791,N_24536);
or U25274 (N_25274,N_22170,N_24193);
nand U25275 (N_25275,N_22458,N_24379);
and U25276 (N_25276,N_21498,N_24911);
and U25277 (N_25277,N_22985,N_20005);
nand U25278 (N_25278,N_24748,N_24530);
and U25279 (N_25279,N_23687,N_21559);
nor U25280 (N_25280,N_20998,N_22313);
nor U25281 (N_25281,N_21690,N_21416);
and U25282 (N_25282,N_20350,N_24289);
xnor U25283 (N_25283,N_22960,N_23715);
or U25284 (N_25284,N_20713,N_20426);
nor U25285 (N_25285,N_24200,N_23919);
or U25286 (N_25286,N_22844,N_24663);
nand U25287 (N_25287,N_24899,N_23191);
xor U25288 (N_25288,N_24864,N_20836);
or U25289 (N_25289,N_20629,N_23182);
nor U25290 (N_25290,N_24670,N_23118);
nor U25291 (N_25291,N_24053,N_21090);
and U25292 (N_25292,N_21263,N_24201);
or U25293 (N_25293,N_22153,N_23765);
nor U25294 (N_25294,N_24500,N_22289);
and U25295 (N_25295,N_22858,N_21696);
xnor U25296 (N_25296,N_23187,N_24927);
nand U25297 (N_25297,N_21829,N_23057);
or U25298 (N_25298,N_24475,N_24662);
xnor U25299 (N_25299,N_22678,N_21560);
and U25300 (N_25300,N_20680,N_24701);
nor U25301 (N_25301,N_22016,N_22491);
xor U25302 (N_25302,N_21668,N_24422);
nand U25303 (N_25303,N_23459,N_24459);
or U25304 (N_25304,N_21568,N_23750);
xor U25305 (N_25305,N_23743,N_23309);
and U25306 (N_25306,N_24859,N_22838);
nand U25307 (N_25307,N_21425,N_24411);
or U25308 (N_25308,N_22558,N_22735);
xor U25309 (N_25309,N_24938,N_22285);
and U25310 (N_25310,N_24623,N_22292);
xnor U25311 (N_25311,N_24144,N_22369);
and U25312 (N_25312,N_22345,N_24431);
nand U25313 (N_25313,N_24044,N_22783);
or U25314 (N_25314,N_21812,N_20472);
nand U25315 (N_25315,N_23149,N_20508);
xor U25316 (N_25316,N_21948,N_22361);
nand U25317 (N_25317,N_24156,N_21291);
and U25318 (N_25318,N_24767,N_23458);
nor U25319 (N_25319,N_23546,N_20790);
nand U25320 (N_25320,N_24183,N_23270);
xnor U25321 (N_25321,N_22332,N_22038);
or U25322 (N_25322,N_22671,N_21827);
nor U25323 (N_25323,N_21601,N_22702);
xnor U25324 (N_25324,N_23924,N_24523);
xnor U25325 (N_25325,N_22748,N_22025);
or U25326 (N_25326,N_24868,N_24094);
and U25327 (N_25327,N_22253,N_22548);
xnor U25328 (N_25328,N_21156,N_24825);
or U25329 (N_25329,N_23404,N_21119);
nor U25330 (N_25330,N_20649,N_23999);
nor U25331 (N_25331,N_20026,N_24355);
or U25332 (N_25332,N_22739,N_24318);
and U25333 (N_25333,N_20112,N_20948);
nor U25334 (N_25334,N_21187,N_22648);
and U25335 (N_25335,N_20670,N_21892);
xor U25336 (N_25336,N_24769,N_21264);
nor U25337 (N_25337,N_21596,N_20532);
and U25338 (N_25338,N_22241,N_22244);
xnor U25339 (N_25339,N_22138,N_21405);
nand U25340 (N_25340,N_21920,N_24760);
xnor U25341 (N_25341,N_22354,N_23284);
xnor U25342 (N_25342,N_23101,N_22612);
nor U25343 (N_25343,N_24031,N_24484);
nor U25344 (N_25344,N_21211,N_20246);
nor U25345 (N_25345,N_22440,N_21066);
or U25346 (N_25346,N_21889,N_22376);
and U25347 (N_25347,N_22578,N_20993);
xnor U25348 (N_25348,N_20415,N_23008);
xnor U25349 (N_25349,N_20947,N_24129);
and U25350 (N_25350,N_20778,N_23222);
nor U25351 (N_25351,N_22413,N_24776);
or U25352 (N_25352,N_23678,N_23592);
xor U25353 (N_25353,N_23666,N_24338);
or U25354 (N_25354,N_21337,N_23751);
and U25355 (N_25355,N_22286,N_24268);
or U25356 (N_25356,N_24891,N_23656);
nand U25357 (N_25357,N_24295,N_20924);
nor U25358 (N_25358,N_22154,N_22570);
nand U25359 (N_25359,N_21323,N_24912);
and U25360 (N_25360,N_21715,N_22027);
and U25361 (N_25361,N_23593,N_23352);
nor U25362 (N_25362,N_24966,N_22177);
or U25363 (N_25363,N_22964,N_24186);
and U25364 (N_25364,N_22122,N_22664);
and U25365 (N_25365,N_20632,N_23099);
or U25366 (N_25366,N_23643,N_22239);
nor U25367 (N_25367,N_22795,N_24904);
nand U25368 (N_25368,N_23598,N_21365);
and U25369 (N_25369,N_24573,N_23671);
or U25370 (N_25370,N_21604,N_23243);
xnor U25371 (N_25371,N_20972,N_24738);
and U25372 (N_25372,N_22372,N_23477);
nor U25373 (N_25373,N_24138,N_22086);
and U25374 (N_25374,N_24194,N_21618);
nand U25375 (N_25375,N_22893,N_20410);
xnor U25376 (N_25376,N_22087,N_22195);
nor U25377 (N_25377,N_21711,N_23201);
xnor U25378 (N_25378,N_21050,N_24319);
or U25379 (N_25379,N_24164,N_21022);
or U25380 (N_25380,N_21762,N_20465);
nor U25381 (N_25381,N_22151,N_20757);
nand U25382 (N_25382,N_21911,N_21124);
nor U25383 (N_25383,N_20341,N_24737);
nor U25384 (N_25384,N_24392,N_21732);
nor U25385 (N_25385,N_21079,N_21114);
or U25386 (N_25386,N_23683,N_22104);
and U25387 (N_25387,N_23513,N_22054);
and U25388 (N_25388,N_21367,N_20057);
nand U25389 (N_25389,N_24477,N_20090);
and U25390 (N_25390,N_24661,N_20366);
nor U25391 (N_25391,N_23398,N_20135);
xor U25392 (N_25392,N_24278,N_21808);
xor U25393 (N_25393,N_22701,N_20884);
or U25394 (N_25394,N_20648,N_20408);
or U25395 (N_25395,N_20595,N_20841);
and U25396 (N_25396,N_20323,N_20722);
and U25397 (N_25397,N_21717,N_24239);
nand U25398 (N_25398,N_21791,N_24922);
or U25399 (N_25399,N_20903,N_20480);
and U25400 (N_25400,N_21997,N_21838);
and U25401 (N_25401,N_20636,N_22791);
xor U25402 (N_25402,N_22642,N_23013);
nand U25403 (N_25403,N_21129,N_22149);
nor U25404 (N_25404,N_23677,N_23966);
or U25405 (N_25405,N_20739,N_20572);
nor U25406 (N_25406,N_22567,N_20367);
xor U25407 (N_25407,N_23328,N_22524);
nand U25408 (N_25408,N_22479,N_20417);
nand U25409 (N_25409,N_24685,N_20440);
or U25410 (N_25410,N_20626,N_20356);
nand U25411 (N_25411,N_24994,N_20463);
xnor U25412 (N_25412,N_20996,N_22564);
nand U25413 (N_25413,N_24054,N_21229);
nor U25414 (N_25414,N_21845,N_24831);
nand U25415 (N_25415,N_23968,N_21626);
nand U25416 (N_25416,N_23824,N_20423);
xor U25417 (N_25417,N_22770,N_24261);
xor U25418 (N_25418,N_23244,N_20889);
or U25419 (N_25419,N_23590,N_23631);
or U25420 (N_25420,N_22159,N_21089);
or U25421 (N_25421,N_23213,N_24024);
and U25422 (N_25422,N_24351,N_22662);
nor U25423 (N_25423,N_23571,N_22487);
or U25424 (N_25424,N_24720,N_20668);
nand U25425 (N_25425,N_20194,N_21496);
or U25426 (N_25426,N_24759,N_23164);
or U25427 (N_25427,N_24280,N_21571);
xnor U25428 (N_25428,N_21897,N_23275);
nor U25429 (N_25429,N_21967,N_20087);
or U25430 (N_25430,N_20442,N_24103);
nand U25431 (N_25431,N_24649,N_20943);
nor U25432 (N_25432,N_22968,N_20765);
xor U25433 (N_25433,N_21544,N_21883);
and U25434 (N_25434,N_20033,N_24528);
nor U25435 (N_25435,N_23637,N_22021);
nand U25436 (N_25436,N_22453,N_21103);
nand U25437 (N_25437,N_21510,N_20506);
xor U25438 (N_25438,N_24975,N_21526);
xor U25439 (N_25439,N_21439,N_20305);
nor U25440 (N_25440,N_21131,N_20692);
or U25441 (N_25441,N_20671,N_21919);
nand U25442 (N_25442,N_22072,N_22449);
xnor U25443 (N_25443,N_24091,N_24644);
or U25444 (N_25444,N_24863,N_20034);
nand U25445 (N_25445,N_23508,N_23699);
xor U25446 (N_25446,N_22992,N_24906);
or U25447 (N_25447,N_22658,N_24507);
or U25448 (N_25448,N_20427,N_21479);
or U25449 (N_25449,N_20176,N_20940);
nand U25450 (N_25450,N_20801,N_20382);
nor U25451 (N_25451,N_23723,N_22922);
nand U25452 (N_25452,N_21631,N_24320);
nor U25453 (N_25453,N_22576,N_24276);
or U25454 (N_25454,N_20961,N_20459);
or U25455 (N_25455,N_22436,N_24726);
and U25456 (N_25456,N_21290,N_21055);
xnor U25457 (N_25457,N_23794,N_22272);
or U25458 (N_25458,N_20273,N_22634);
nor U25459 (N_25459,N_24625,N_24145);
nand U25460 (N_25460,N_22118,N_22304);
and U25461 (N_25461,N_24556,N_21484);
or U25462 (N_25462,N_22473,N_20422);
nor U25463 (N_25463,N_20104,N_23853);
and U25464 (N_25464,N_20172,N_24826);
or U25465 (N_25465,N_21606,N_22687);
or U25466 (N_25466,N_24395,N_20134);
nor U25467 (N_25467,N_21790,N_21186);
nand U25468 (N_25468,N_20822,N_24941);
and U25469 (N_25469,N_21648,N_24225);
nor U25470 (N_25470,N_23464,N_21584);
nor U25471 (N_25471,N_20842,N_22596);
nor U25472 (N_25472,N_23886,N_22415);
nor U25473 (N_25473,N_20405,N_24712);
nor U25474 (N_25474,N_20467,N_21192);
or U25475 (N_25475,N_23361,N_20977);
xnor U25476 (N_25476,N_21470,N_24928);
or U25477 (N_25477,N_20326,N_24036);
and U25478 (N_25478,N_22904,N_21443);
or U25479 (N_25479,N_22534,N_20301);
and U25480 (N_25480,N_23491,N_22952);
and U25481 (N_25481,N_21321,N_23077);
or U25482 (N_25482,N_23448,N_21619);
or U25483 (N_25483,N_20954,N_21835);
or U25484 (N_25484,N_22489,N_20343);
nand U25485 (N_25485,N_23541,N_20897);
nand U25486 (N_25486,N_22360,N_20566);
xor U25487 (N_25487,N_22417,N_23254);
or U25488 (N_25488,N_20991,N_20918);
and U25489 (N_25489,N_23301,N_23321);
xor U25490 (N_25490,N_24761,N_23157);
nor U25491 (N_25491,N_24582,N_22056);
and U25492 (N_25492,N_24803,N_24705);
nor U25493 (N_25493,N_20028,N_24561);
and U25494 (N_25494,N_24232,N_21266);
and U25495 (N_25495,N_24744,N_21621);
nand U25496 (N_25496,N_22990,N_23365);
and U25497 (N_25497,N_23808,N_21227);
or U25498 (N_25498,N_22877,N_21969);
and U25499 (N_25499,N_21569,N_20274);
nor U25500 (N_25500,N_21549,N_20660);
and U25501 (N_25501,N_23027,N_24821);
nor U25502 (N_25502,N_24518,N_22788);
and U25503 (N_25503,N_24403,N_23460);
nand U25504 (N_25504,N_21137,N_23906);
xnor U25505 (N_25505,N_21878,N_22568);
nand U25506 (N_25506,N_20288,N_21909);
or U25507 (N_25507,N_22937,N_23597);
nand U25508 (N_25508,N_20169,N_21538);
and U25509 (N_25509,N_20736,N_20447);
nand U25510 (N_25510,N_23295,N_21358);
nor U25511 (N_25511,N_24315,N_20310);
xor U25512 (N_25512,N_20073,N_24438);
and U25513 (N_25513,N_23257,N_21442);
and U25514 (N_25514,N_20558,N_23556);
or U25515 (N_25515,N_22825,N_24961);
nor U25516 (N_25516,N_23069,N_20594);
xnor U25517 (N_25517,N_22359,N_24133);
nor U25518 (N_25518,N_24324,N_22076);
or U25519 (N_25519,N_20704,N_24581);
xnor U25520 (N_25520,N_24757,N_20936);
nand U25521 (N_25521,N_21966,N_22721);
and U25522 (N_25522,N_22744,N_24163);
and U25523 (N_25523,N_23675,N_23997);
nor U25524 (N_25524,N_21952,N_24572);
or U25525 (N_25525,N_23713,N_21190);
nor U25526 (N_25526,N_20345,N_21359);
xor U25527 (N_25527,N_24897,N_21212);
or U25528 (N_25528,N_23126,N_24995);
or U25529 (N_25529,N_23625,N_24082);
nor U25530 (N_25530,N_21929,N_23431);
nor U25531 (N_25531,N_20563,N_20153);
nor U25532 (N_25532,N_21152,N_22490);
or U25533 (N_25533,N_23955,N_23833);
xor U25534 (N_25534,N_24235,N_24428);
nor U25535 (N_25535,N_24134,N_24447);
nor U25536 (N_25536,N_24963,N_24955);
and U25537 (N_25537,N_20512,N_20952);
nand U25538 (N_25538,N_21304,N_20866);
or U25539 (N_25539,N_21087,N_24181);
or U25540 (N_25540,N_21928,N_22517);
or U25541 (N_25541,N_23642,N_21215);
and U25542 (N_25542,N_21315,N_23959);
nand U25543 (N_25543,N_24992,N_21347);
or U25544 (N_25544,N_23397,N_21608);
or U25545 (N_25545,N_20285,N_23658);
nor U25546 (N_25546,N_22395,N_21729);
or U25547 (N_25547,N_21265,N_23623);
xor U25548 (N_25548,N_24676,N_21387);
nand U25549 (N_25549,N_22181,N_24273);
and U25550 (N_25550,N_21609,N_23132);
nand U25551 (N_25551,N_24279,N_21168);
or U25552 (N_25552,N_23847,N_24310);
nor U25553 (N_25553,N_20125,N_24820);
xnor U25554 (N_25554,N_20351,N_24943);
nor U25555 (N_25555,N_22431,N_21644);
xor U25556 (N_25556,N_22150,N_21408);
or U25557 (N_25557,N_24371,N_21639);
xnor U25558 (N_25558,N_20839,N_21692);
nand U25559 (N_25559,N_22839,N_22256);
nor U25560 (N_25560,N_24335,N_23706);
nor U25561 (N_25561,N_24646,N_22466);
and U25562 (N_25562,N_22592,N_21853);
nand U25563 (N_25563,N_20596,N_22861);
and U25564 (N_25564,N_24118,N_24951);
xnor U25565 (N_25565,N_24952,N_22705);
nor U25566 (N_25566,N_24450,N_21918);
nor U25567 (N_25567,N_24296,N_24935);
nand U25568 (N_25568,N_24389,N_21122);
nand U25569 (N_25569,N_21313,N_22514);
nand U25570 (N_25570,N_22204,N_22680);
nor U25571 (N_25571,N_21814,N_23520);
and U25572 (N_25572,N_22652,N_22198);
xnor U25573 (N_25573,N_24286,N_23363);
nor U25574 (N_25574,N_23539,N_24023);
and U25575 (N_25575,N_22965,N_23807);
nor U25576 (N_25576,N_20813,N_24424);
and U25577 (N_25577,N_21553,N_21851);
nor U25578 (N_25578,N_20272,N_24226);
or U25579 (N_25579,N_24209,N_24215);
xor U25580 (N_25580,N_20796,N_20437);
nand U25581 (N_25581,N_22532,N_21436);
xnor U25582 (N_25582,N_20721,N_23879);
or U25583 (N_25583,N_23729,N_22722);
or U25584 (N_25584,N_21689,N_20612);
nand U25585 (N_25585,N_23866,N_22165);
xor U25586 (N_25586,N_24949,N_24298);
nor U25587 (N_25587,N_21655,N_24139);
xor U25588 (N_25588,N_22433,N_20521);
and U25589 (N_25589,N_24216,N_20755);
or U25590 (N_25590,N_20280,N_21084);
xnor U25591 (N_25591,N_21882,N_21237);
xor U25592 (N_25592,N_23920,N_23504);
nand U25593 (N_25593,N_20114,N_23992);
or U25594 (N_25594,N_24168,N_24367);
xnor U25595 (N_25595,N_21540,N_21048);
and U25596 (N_25596,N_23022,N_21423);
nor U25597 (N_25597,N_23078,N_21412);
and U25598 (N_25598,N_20456,N_20344);
and U25599 (N_25599,N_24080,N_21521);
nor U25600 (N_25600,N_23233,N_23024);
nand U25601 (N_25601,N_24327,N_23472);
and U25602 (N_25602,N_22771,N_20881);
xor U25603 (N_25603,N_24030,N_24714);
nor U25604 (N_25604,N_21749,N_23143);
nor U25605 (N_25605,N_22723,N_20123);
or U25606 (N_25606,N_21763,N_24948);
and U25607 (N_25607,N_23602,N_20475);
nor U25608 (N_25608,N_21638,N_24733);
nor U25609 (N_25609,N_20605,N_20095);
or U25610 (N_25610,N_20781,N_20313);
nor U25611 (N_25611,N_22190,N_20872);
nor U25612 (N_25612,N_21891,N_24397);
nand U25613 (N_25613,N_22942,N_24207);
nand U25614 (N_25614,N_23926,N_21707);
nand U25615 (N_25615,N_23033,N_21098);
nand U25616 (N_25616,N_23704,N_23741);
xnor U25617 (N_25617,N_23559,N_21058);
and U25618 (N_25618,N_20147,N_20635);
or U25619 (N_25619,N_23672,N_23122);
and U25620 (N_25620,N_22617,N_24406);
xnor U25621 (N_25621,N_22520,N_20204);
and U25622 (N_25622,N_22069,N_23311);
or U25623 (N_25623,N_20390,N_20577);
xnor U25624 (N_25624,N_24946,N_21861);
xnor U25625 (N_25625,N_22618,N_20603);
nand U25626 (N_25626,N_20187,N_20453);
or U25627 (N_25627,N_24307,N_21377);
nor U25628 (N_25628,N_21547,N_20609);
and U25629 (N_25629,N_20283,N_22827);
xnor U25630 (N_25630,N_22966,N_21870);
or U25631 (N_25631,N_22023,N_21730);
and U25632 (N_25632,N_24102,N_24214);
nor U25633 (N_25633,N_24543,N_23910);
or U25634 (N_25634,N_21823,N_24910);
nand U25635 (N_25635,N_21978,N_21983);
xor U25636 (N_25636,N_24690,N_23500);
and U25637 (N_25637,N_20476,N_23188);
and U25638 (N_25638,N_23525,N_24981);
nand U25639 (N_25639,N_24258,N_21522);
or U25640 (N_25640,N_24854,N_22280);
xor U25641 (N_25641,N_24743,N_24627);
or U25642 (N_25642,N_23829,N_24056);
or U25643 (N_25643,N_20847,N_24441);
xnor U25644 (N_25644,N_23473,N_24741);
and U25645 (N_25645,N_23962,N_21222);
nand U25646 (N_25646,N_23362,N_20569);
nand U25647 (N_25647,N_23944,N_22044);
or U25648 (N_25648,N_21368,N_24998);
or U25649 (N_25649,N_21165,N_23260);
nor U25650 (N_25650,N_23917,N_20416);
nand U25651 (N_25651,N_20484,N_20987);
nand U25652 (N_25652,N_20047,N_23049);
nand U25653 (N_25653,N_21704,N_20213);
nor U25654 (N_25654,N_22537,N_24346);
xnor U25655 (N_25655,N_20883,N_24606);
nor U25656 (N_25656,N_23890,N_24378);
nand U25657 (N_25657,N_22805,N_20231);
xor U25658 (N_25658,N_21480,N_24242);
xnor U25659 (N_25659,N_24850,N_20769);
or U25660 (N_25660,N_22420,N_21998);
nand U25661 (N_25661,N_24049,N_24617);
nor U25662 (N_25662,N_21663,N_21224);
nand U25663 (N_25663,N_22862,N_21041);
nand U25664 (N_25664,N_24281,N_23685);
nor U25665 (N_25665,N_24973,N_21896);
or U25666 (N_25666,N_22914,N_22814);
or U25667 (N_25667,N_22613,N_23652);
and U25668 (N_25668,N_23901,N_20579);
and U25669 (N_25669,N_20817,N_23185);
or U25670 (N_25670,N_22784,N_23900);
nor U25671 (N_25671,N_24212,N_23040);
nor U25672 (N_25672,N_22986,N_21932);
nor U25673 (N_25673,N_20229,N_23392);
nor U25674 (N_25674,N_21503,N_20782);
and U25675 (N_25675,N_21016,N_24639);
and U25676 (N_25676,N_21632,N_20767);
and U25677 (N_25677,N_21996,N_23865);
nor U25678 (N_25678,N_24585,N_20048);
nor U25679 (N_25679,N_23567,N_21507);
nor U25680 (N_25680,N_21024,N_24234);
xnor U25681 (N_25681,N_20319,N_24121);
and U25682 (N_25682,N_22005,N_23483);
and U25683 (N_25683,N_23358,N_24348);
and U25684 (N_25684,N_21714,N_23795);
and U25685 (N_25685,N_20336,N_24512);
or U25686 (N_25686,N_20585,N_23839);
nor U25687 (N_25687,N_24464,N_22624);
and U25688 (N_25688,N_21976,N_23297);
nor U25689 (N_25689,N_20260,N_20528);
xor U25690 (N_25690,N_23071,N_23595);
nand U25691 (N_25691,N_23084,N_22733);
xor U25692 (N_25692,N_22111,N_21760);
or U25693 (N_25693,N_23147,N_20877);
nor U25694 (N_25694,N_20543,N_21537);
xnor U25695 (N_25695,N_24001,N_23911);
nand U25696 (N_25696,N_24506,N_22080);
or U25697 (N_25697,N_20262,N_22823);
or U25698 (N_25698,N_20400,N_20909);
nand U25699 (N_25699,N_22673,N_24233);
and U25700 (N_25700,N_22444,N_21355);
nor U25701 (N_25701,N_21134,N_23972);
nor U25702 (N_25702,N_23679,N_22632);
or U25703 (N_25703,N_20462,N_21251);
and U25704 (N_25704,N_21719,N_20036);
xor U25705 (N_25705,N_24965,N_24983);
or U25706 (N_25706,N_24010,N_21640);
or U25707 (N_25707,N_21000,N_20523);
or U25708 (N_25708,N_23619,N_23011);
xor U25709 (N_25709,N_23494,N_24037);
nor U25710 (N_25710,N_21598,N_21872);
or U25711 (N_25711,N_21868,N_24900);
nand U25712 (N_25712,N_20161,N_23273);
or U25713 (N_25713,N_20023,N_22629);
or U25714 (N_25714,N_23463,N_21984);
nand U25715 (N_25715,N_22527,N_21570);
xnor U25716 (N_25716,N_20143,N_24866);
nor U25717 (N_25717,N_21444,N_23577);
nor U25718 (N_25718,N_23239,N_21019);
or U25719 (N_25719,N_22248,N_23991);
or U25720 (N_25720,N_22984,N_20190);
nor U25721 (N_25721,N_21685,N_22684);
nor U25722 (N_25722,N_23413,N_24544);
nor U25723 (N_25723,N_24734,N_22319);
and U25724 (N_25724,N_22365,N_24336);
and U25725 (N_25725,N_24962,N_21776);
nor U25726 (N_25726,N_23517,N_21670);
and U25727 (N_25727,N_23217,N_23904);
xor U25728 (N_25728,N_23582,N_22225);
nand U25729 (N_25729,N_23640,N_21253);
and U25730 (N_25730,N_23970,N_20074);
nor U25731 (N_25731,N_24122,N_24236);
nand U25732 (N_25732,N_24658,N_22526);
or U25733 (N_25733,N_23133,N_22075);
nand U25734 (N_25734,N_24501,N_20941);
xor U25735 (N_25735,N_24025,N_22657);
nor U25736 (N_25736,N_22626,N_24839);
nand U25737 (N_25737,N_20086,N_20383);
nand U25738 (N_25738,N_23444,N_20752);
nor U25739 (N_25739,N_22793,N_20332);
and U25740 (N_25740,N_21179,N_23424);
nand U25741 (N_25741,N_22516,N_20157);
xnor U25742 (N_25742,N_23641,N_21712);
nor U25743 (N_25743,N_22979,N_22268);
nand U25744 (N_25744,N_20072,N_24774);
nand U25745 (N_25745,N_23140,N_23106);
nand U25746 (N_25746,N_24947,N_24255);
nand U25747 (N_25747,N_20145,N_20598);
nand U25748 (N_25748,N_23315,N_20777);
nand U25749 (N_25749,N_21478,N_22009);
nor U25750 (N_25750,N_22379,N_22908);
xor U25751 (N_25751,N_20679,N_20448);
and U25752 (N_25752,N_23976,N_22367);
and U25753 (N_25753,N_21071,N_23942);
xnor U25754 (N_25754,N_21562,N_20725);
xor U25755 (N_25755,N_24481,N_21258);
and U25756 (N_25756,N_22654,N_21455);
and U25757 (N_25757,N_22529,N_23323);
nor U25758 (N_25758,N_21486,N_23802);
xor U25759 (N_25759,N_23466,N_21783);
nand U25760 (N_25760,N_21832,N_22299);
nor U25761 (N_25761,N_24722,N_22539);
or U25762 (N_25762,N_21037,N_20256);
or U25763 (N_25763,N_20450,N_21680);
and U25764 (N_25764,N_24496,N_23343);
nor U25765 (N_25765,N_20815,N_23462);
nand U25766 (N_25766,N_21171,N_24393);
nand U25767 (N_25767,N_20487,N_22872);
nor U25768 (N_25768,N_20975,N_24460);
or U25769 (N_25769,N_21822,N_22242);
xor U25770 (N_25770,N_22685,N_21199);
and U25771 (N_25771,N_24476,N_23418);
xnor U25772 (N_25772,N_20944,N_23044);
nor U25773 (N_25773,N_23804,N_24195);
or U25774 (N_25774,N_21789,N_24696);
xor U25775 (N_25775,N_20240,N_21599);
xnor U25776 (N_25776,N_20014,N_20444);
nand U25777 (N_25777,N_21748,N_21208);
or U25778 (N_25778,N_21907,N_21843);
nor U25779 (N_25779,N_21453,N_24905);
or U25780 (N_25780,N_24925,N_22951);
and U25781 (N_25781,N_24550,N_21993);
and U25782 (N_25782,N_24835,N_23584);
nor U25783 (N_25783,N_21534,N_21021);
nor U25784 (N_25784,N_21106,N_23821);
or U25785 (N_25785,N_22330,N_21279);
or U25786 (N_25786,N_23407,N_23799);
nor U25787 (N_25787,N_24125,N_21550);
and U25788 (N_25788,N_20178,N_21421);
nor U25789 (N_25789,N_22187,N_23394);
nor U25790 (N_25790,N_21456,N_24399);
xnor U25791 (N_25791,N_22553,N_21572);
or U25792 (N_25792,N_20261,N_22841);
nand U25793 (N_25793,N_21849,N_23158);
or U25794 (N_25794,N_23774,N_21325);
and U25795 (N_25795,N_20582,N_21816);
xnor U25796 (N_25796,N_24028,N_22590);
and U25797 (N_25797,N_24112,N_22983);
xnor U25798 (N_25798,N_23415,N_24456);
xor U25799 (N_25799,N_23410,N_22710);
nor U25800 (N_25800,N_20858,N_22938);
xor U25801 (N_25801,N_22847,N_23048);
nor U25802 (N_25802,N_21310,N_20296);
xor U25803 (N_25803,N_20251,N_20624);
nor U25804 (N_25804,N_23455,N_20921);
and U25805 (N_25805,N_24684,N_24557);
nand U25806 (N_25806,N_23896,N_21532);
or U25807 (N_25807,N_22586,N_22559);
and U25808 (N_25808,N_20525,N_20901);
or U25809 (N_25809,N_23420,N_22092);
or U25810 (N_25810,N_21858,N_22425);
nand U25811 (N_25811,N_20942,N_20719);
xnor U25812 (N_25812,N_23874,N_21681);
nand U25813 (N_25813,N_23851,N_23752);
and U25814 (N_25814,N_21163,N_24979);
and U25815 (N_25815,N_23744,N_24751);
nor U25816 (N_25816,N_20929,N_24435);
xnor U25817 (N_25817,N_22727,N_24075);
xnor U25818 (N_25818,N_22905,N_20698);
or U25819 (N_25819,N_23863,N_22643);
nand U25820 (N_25820,N_22736,N_22630);
nor U25821 (N_25821,N_23555,N_24791);
nand U25822 (N_25822,N_23279,N_23025);
and U25823 (N_25823,N_20193,N_20578);
or U25824 (N_25824,N_20144,N_24560);
or U25825 (N_25825,N_23083,N_24569);
or U25826 (N_25826,N_22587,N_21293);
or U25827 (N_25827,N_24576,N_24203);
or U25828 (N_25828,N_23519,N_24587);
nor U25829 (N_25829,N_22329,N_24309);
xnor U25830 (N_25830,N_23878,N_22237);
and U25831 (N_25831,N_21117,N_24603);
and U25832 (N_25832,N_24547,N_22866);
xor U25833 (N_25833,N_21731,N_20129);
or U25834 (N_25834,N_23803,N_22456);
and U25835 (N_25835,N_21857,N_23880);
xor U25836 (N_25836,N_20154,N_24069);
nand U25837 (N_25837,N_22842,N_20760);
nand U25838 (N_25838,N_21351,N_22963);
or U25839 (N_25839,N_20820,N_23936);
xnor U25840 (N_25840,N_20547,N_24816);
nor U25841 (N_25841,N_20130,N_22804);
xnor U25842 (N_25842,N_21629,N_24954);
and U25843 (N_25843,N_22310,N_21424);
or U25844 (N_25844,N_24546,N_21457);
nand U25845 (N_25845,N_22469,N_22001);
nor U25846 (N_25846,N_23489,N_24457);
xor U25847 (N_25847,N_24248,N_20481);
nand U25848 (N_25848,N_24551,N_24380);
and U25849 (N_25849,N_23241,N_20191);
xnor U25850 (N_25850,N_24051,N_23638);
xnor U25851 (N_25851,N_23700,N_22531);
and U25852 (N_25852,N_23894,N_21713);
nand U25853 (N_25853,N_23979,N_20992);
and U25854 (N_25854,N_20804,N_21985);
nand U25855 (N_25855,N_24356,N_21500);
and U25856 (N_25856,N_20223,N_20056);
xnor U25857 (N_25857,N_24000,N_22133);
and U25858 (N_25858,N_23544,N_20318);
and U25859 (N_25859,N_20016,N_21311);
or U25860 (N_25860,N_21374,N_21203);
nor U25861 (N_25861,N_21980,N_20843);
xnor U25862 (N_25862,N_24648,N_23947);
nor U25863 (N_25863,N_20333,N_20140);
xnor U25864 (N_25864,N_21587,N_20714);
or U25865 (N_25865,N_23051,N_24784);
and U25866 (N_25866,N_23216,N_23238);
nand U25867 (N_25867,N_23446,N_20166);
and U25868 (N_25868,N_22335,N_22145);
or U25869 (N_25869,N_22096,N_21318);
nand U25870 (N_25870,N_22399,N_24837);
or U25871 (N_25871,N_21968,N_20254);
nand U25872 (N_25872,N_21174,N_21452);
nor U25873 (N_25873,N_22315,N_22119);
nand U25874 (N_25874,N_20818,N_22382);
and U25875 (N_25875,N_20374,N_22621);
and U25876 (N_25876,N_24440,N_23585);
nand U25877 (N_25877,N_22696,N_23667);
nor U25878 (N_25878,N_24852,N_22502);
xor U25879 (N_25879,N_22424,N_20741);
or U25880 (N_25880,N_21874,N_22203);
nand U25881 (N_25881,N_22752,N_24610);
xnor U25882 (N_25882,N_21652,N_21092);
or U25883 (N_25883,N_22607,N_23940);
and U25884 (N_25884,N_21958,N_20926);
xnor U25885 (N_25885,N_23629,N_20619);
xor U25886 (N_25886,N_22731,N_22598);
nand U25887 (N_25887,N_22348,N_21172);
xnor U25888 (N_25888,N_21778,N_24077);
and U25889 (N_25889,N_21141,N_24875);
nor U25890 (N_25890,N_23387,N_23097);
nor U25891 (N_25891,N_22697,N_20496);
xor U25892 (N_25892,N_20559,N_24341);
xnor U25893 (N_25893,N_24656,N_21846);
xnor U25894 (N_25894,N_24176,N_20962);
xnor U25895 (N_25895,N_21516,N_24865);
nor U25896 (N_25896,N_22467,N_22480);
nor U25897 (N_25897,N_24762,N_22068);
xnor U25898 (N_25898,N_22157,N_23684);
or U25899 (N_25899,N_22577,N_21177);
or U25900 (N_25900,N_24531,N_23950);
or U25901 (N_25901,N_23026,N_21379);
and U25902 (N_25902,N_23134,N_23702);
nor U25903 (N_25903,N_24908,N_24675);
nand U25904 (N_25904,N_23633,N_21396);
nand U25905 (N_25905,N_24664,N_23128);
xor U25906 (N_25906,N_24048,N_20970);
or U25907 (N_25907,N_21828,N_20862);
or U25908 (N_25908,N_20650,N_23050);
and U25909 (N_25909,N_22512,N_22840);
nand U25910 (N_25910,N_23432,N_21196);
and U25911 (N_25911,N_24143,N_23037);
nor U25912 (N_25912,N_21939,N_21605);
or U25913 (N_25913,N_23053,N_23355);
nand U25914 (N_25914,N_24797,N_21394);
and U25915 (N_25915,N_24246,N_24206);
nor U25916 (N_25916,N_23199,N_23998);
xnor U25917 (N_25917,N_21994,N_21061);
nand U25918 (N_25918,N_23395,N_24291);
or U25919 (N_25919,N_21990,N_20402);
nor U25920 (N_25920,N_21406,N_22616);
nand U25921 (N_25921,N_23747,N_22714);
and U25922 (N_25922,N_24124,N_24593);
xnor U25923 (N_25923,N_20561,N_22000);
nand U25924 (N_25924,N_23219,N_24860);
nand U25925 (N_25925,N_20075,N_20032);
or U25926 (N_25926,N_23042,N_22611);
and U25927 (N_25927,N_21038,N_23289);
nand U25928 (N_25928,N_21362,N_21922);
nor U25929 (N_25929,N_22868,N_23790);
nand U25930 (N_25930,N_21342,N_20181);
nand U25931 (N_25931,N_22972,N_23594);
xor U25932 (N_25932,N_23971,N_24260);
or U25933 (N_25933,N_23722,N_21151);
nand U25934 (N_25934,N_24978,N_23952);
and U25935 (N_25935,N_20923,N_21697);
xor U25936 (N_25936,N_20779,N_20118);
or U25937 (N_25937,N_20728,N_22135);
xor U25938 (N_25938,N_20531,N_23163);
and U25939 (N_25939,N_24007,N_21767);
or U25940 (N_25940,N_22167,N_22130);
or U25941 (N_25941,N_22546,N_23903);
nand U25942 (N_25942,N_20357,N_20322);
nor U25943 (N_25943,N_21126,N_23495);
or U25944 (N_25944,N_20003,N_20854);
nor U25945 (N_25945,N_24401,N_22929);
or U25946 (N_25946,N_24704,N_20389);
nor U25947 (N_25947,N_23875,N_20425);
nand U25948 (N_25948,N_24063,N_22890);
or U25949 (N_25949,N_22059,N_22174);
nand U25950 (N_25950,N_21660,N_23727);
and U25951 (N_25951,N_24109,N_24843);
xor U25952 (N_25952,N_21418,N_23015);
or U25953 (N_25953,N_24615,N_20826);
and U25954 (N_25954,N_24208,N_20794);
nand U25955 (N_25955,N_22740,N_24631);
and U25956 (N_25956,N_20676,N_24220);
or U25957 (N_25957,N_22811,N_24502);
nand U25958 (N_25958,N_22428,N_21664);
and U25959 (N_25959,N_20932,N_21001);
and U25960 (N_25960,N_20838,N_23482);
nand U25961 (N_25961,N_22062,N_21003);
nor U25962 (N_25962,N_22820,N_23502);
and U25963 (N_25963,N_20379,N_24408);
nand U25964 (N_25964,N_24828,N_21947);
or U25965 (N_25965,N_22269,N_24482);
and U25966 (N_25966,N_20709,N_24192);
and U25967 (N_25967,N_20404,N_22391);
nand U25968 (N_25968,N_21683,N_21032);
nand U25969 (N_25969,N_22750,N_23695);
and U25970 (N_25970,N_20951,N_24014);
or U25971 (N_25971,N_24834,N_21241);
and U25972 (N_25972,N_20233,N_24537);
nor U25973 (N_25973,N_23166,N_21261);
xor U25974 (N_25974,N_21701,N_23719);
nor U25975 (N_25975,N_20656,N_20368);
xor U25976 (N_25976,N_22211,N_23573);
xor U25977 (N_25977,N_23212,N_24719);
nor U25978 (N_25978,N_22462,N_24283);
or U25979 (N_25979,N_20754,N_23204);
or U25980 (N_25980,N_23545,N_23644);
nor U25981 (N_25981,N_23324,N_20433);
and U25982 (N_25982,N_21975,N_22845);
xor U25983 (N_25983,N_23079,N_23030);
and U25984 (N_25984,N_21794,N_22316);
xnor U25985 (N_25985,N_21916,N_23167);
nand U25986 (N_25986,N_22064,N_24135);
and U25987 (N_25987,N_21955,N_21676);
and U25988 (N_25988,N_21779,N_23646);
nand U25989 (N_25989,N_23510,N_20832);
and U25990 (N_25990,N_22194,N_21232);
nor U25991 (N_25991,N_21879,N_24329);
xor U25992 (N_25992,N_24731,N_20985);
and U25993 (N_25993,N_24755,N_21964);
or U25994 (N_25994,N_24715,N_22519);
or U25995 (N_25995,N_21623,N_20238);
nand U25996 (N_25996,N_24364,N_23989);
nor U25997 (N_25997,N_22726,N_20946);
nor U25998 (N_25998,N_24858,N_22505);
xnor U25999 (N_25999,N_22229,N_23341);
or U26000 (N_26000,N_23198,N_24641);
or U26001 (N_26001,N_23660,N_23738);
nand U26002 (N_26002,N_20673,N_23819);
and U26003 (N_26003,N_21111,N_23960);
nor U26004 (N_26004,N_24786,N_23227);
and U26005 (N_26005,N_20589,N_23296);
xor U26006 (N_26006,N_22255,N_24416);
or U26007 (N_26007,N_24699,N_24359);
nand U26008 (N_26008,N_21875,N_21414);
nand U26009 (N_26009,N_24499,N_24771);
xnor U26010 (N_26010,N_21799,N_23414);
nand U26011 (N_26011,N_23428,N_20639);
nand U26012 (N_26012,N_24832,N_21161);
xor U26013 (N_26013,N_23845,N_24926);
and U26014 (N_26014,N_20196,N_22606);
and U26015 (N_26015,N_20949,N_20266);
and U26016 (N_26016,N_20180,N_22902);
nor U26017 (N_26017,N_20327,N_22794);
or U26018 (N_26018,N_20756,N_23850);
nand U26019 (N_26019,N_23694,N_20316);
or U26020 (N_26020,N_24936,N_21110);
nand U26021 (N_26021,N_22459,N_22495);
nor U26022 (N_26022,N_22342,N_22364);
and U26023 (N_26023,N_22222,N_20038);
nand U26024 (N_26024,N_24349,N_23797);
nand U26025 (N_26025,N_22208,N_22834);
and U26026 (N_26026,N_23052,N_24680);
xor U26027 (N_26027,N_22344,N_23181);
nor U26028 (N_26028,N_22781,N_23653);
or U26029 (N_26029,N_20451,N_24184);
and U26030 (N_26030,N_21228,N_20111);
and U26031 (N_26031,N_22446,N_22689);
and U26032 (N_26032,N_21612,N_20517);
xor U26033 (N_26033,N_20738,N_24989);
or U26034 (N_26034,N_20165,N_23786);
and U26035 (N_26035,N_21543,N_23654);
xnor U26036 (N_26036,N_21128,N_21205);
and U26037 (N_26037,N_22460,N_22883);
xnor U26038 (N_26038,N_23788,N_20493);
nand U26039 (N_26039,N_23223,N_22454);
nand U26040 (N_26040,N_20179,N_20564);
or U26041 (N_26041,N_24308,N_20269);
nor U26042 (N_26042,N_22351,N_22055);
xor U26043 (N_26043,N_22058,N_22110);
or U26044 (N_26044,N_24126,N_20329);
xnor U26045 (N_26045,N_24756,N_22173);
nor U26046 (N_26046,N_21235,N_23169);
and U26047 (N_26047,N_20835,N_21751);
xnor U26048 (N_26048,N_21216,N_23669);
nor U26049 (N_26049,N_24097,N_24702);
nor U26050 (N_26050,N_21999,N_20497);
or U26051 (N_26051,N_21720,N_22541);
xnor U26052 (N_26052,N_21149,N_20460);
nand U26053 (N_26053,N_22168,N_22756);
nand U26054 (N_26054,N_20807,N_21404);
nor U26055 (N_26055,N_22363,N_22392);
and U26056 (N_26056,N_22482,N_20378);
nor U26057 (N_26057,N_22716,N_21393);
nor U26058 (N_26058,N_22228,N_20823);
nor U26059 (N_26059,N_23172,N_20337);
xnor U26060 (N_26060,N_24174,N_23983);
or U26061 (N_26061,N_22653,N_23728);
xor U26062 (N_26062,N_20363,N_24177);
xor U26063 (N_26063,N_23630,N_23884);
nor U26064 (N_26064,N_22260,N_23116);
nand U26065 (N_26065,N_21565,N_20905);
or U26066 (N_26066,N_22747,N_23749);
and U26067 (N_26067,N_20167,N_23412);
and U26068 (N_26068,N_22676,N_23287);
or U26069 (N_26069,N_20593,N_20824);
nand U26070 (N_26070,N_23215,N_23342);
nand U26071 (N_26071,N_22535,N_22909);
nor U26072 (N_26072,N_21147,N_22728);
nand U26073 (N_26073,N_22544,N_23557);
nor U26074 (N_26074,N_23381,N_22147);
nand U26075 (N_26075,N_22878,N_21275);
nor U26076 (N_26076,N_21567,N_23221);
or U26077 (N_26077,N_22293,N_23721);
xnor U26078 (N_26078,N_20070,N_24802);
and U26079 (N_26079,N_20546,N_22143);
xor U26080 (N_26080,N_24350,N_23689);
or U26081 (N_26081,N_20995,N_22022);
xnor U26082 (N_26082,N_21946,N_23138);
xor U26083 (N_26083,N_23812,N_20339);
and U26084 (N_26084,N_23197,N_22427);
or U26085 (N_26085,N_22717,N_20792);
xnor U26086 (N_26086,N_24509,N_24415);
xnor U26087 (N_26087,N_20277,N_20912);
and U26088 (N_26088,N_24347,N_23347);
nand U26089 (N_26089,N_20768,N_23409);
xor U26090 (N_26090,N_23515,N_21081);
nor U26091 (N_26091,N_20170,N_24713);
and U26092 (N_26092,N_23070,N_21082);
or U26093 (N_26093,N_22619,N_22711);
nand U26094 (N_26094,N_22830,N_21206);
and U26095 (N_26095,N_23888,N_21908);
or U26096 (N_26096,N_21684,N_22083);
nor U26097 (N_26097,N_20930,N_23600);
and U26098 (N_26098,N_23081,N_21085);
and U26099 (N_26099,N_23913,N_23531);
nor U26100 (N_26100,N_22832,N_23461);
nand U26101 (N_26101,N_22886,N_20142);
xor U26102 (N_26102,N_20662,N_24374);
nand U26103 (N_26103,N_24534,N_21184);
nor U26104 (N_26104,N_24190,N_23760);
nor U26105 (N_26105,N_21035,N_21804);
or U26106 (N_26106,N_20518,N_23607);
xnor U26107 (N_26107,N_22871,N_23813);
xor U26108 (N_26108,N_22057,N_21746);
nor U26109 (N_26109,N_23237,N_21514);
and U26110 (N_26110,N_23977,N_22227);
nor U26111 (N_26111,N_21146,N_23360);
or U26112 (N_26112,N_24923,N_20735);
xnor U26113 (N_26113,N_20252,N_20700);
xnor U26114 (N_26114,N_24003,N_20141);
and U26115 (N_26115,N_23834,N_21489);
xnor U26116 (N_26116,N_22924,N_24806);
and U26117 (N_26117,N_24407,N_24874);
or U26118 (N_26118,N_23601,N_21933);
or U26119 (N_26119,N_22352,N_24727);
nor U26120 (N_26120,N_21625,N_24013);
and U26121 (N_26121,N_22806,N_20395);
and U26122 (N_26122,N_20094,N_21088);
nand U26123 (N_26123,N_21356,N_23986);
or U26124 (N_26124,N_24357,N_22798);
xnor U26125 (N_26125,N_22860,N_20207);
xnor U26126 (N_26126,N_20984,N_22870);
nand U26127 (N_26127,N_21166,N_24605);
and U26128 (N_26128,N_20317,N_20783);
or U26129 (N_26129,N_21504,N_20584);
and U26130 (N_26130,N_23209,N_22790);
xor U26131 (N_26131,N_21903,N_20221);
or U26132 (N_26132,N_20004,N_23160);
xor U26133 (N_26133,N_20774,N_20910);
or U26134 (N_26134,N_22192,N_20064);
xnor U26135 (N_26135,N_24391,N_22421);
and U26136 (N_26136,N_21523,N_20297);
and U26137 (N_26137,N_20136,N_24467);
xnor U26138 (N_26138,N_24698,N_23836);
xor U26139 (N_26139,N_22561,N_20498);
nor U26140 (N_26140,N_20232,N_24065);
and U26141 (N_26141,N_22692,N_20122);
nand U26142 (N_26142,N_20119,N_21806);
or U26143 (N_26143,N_20681,N_24886);
nor U26144 (N_26144,N_20483,N_23162);
and U26145 (N_26145,N_23634,N_23467);
and U26146 (N_26146,N_24497,N_22900);
or U26147 (N_26147,N_20377,N_24294);
or U26148 (N_26148,N_24478,N_20988);
nand U26149 (N_26149,N_20084,N_20644);
nand U26150 (N_26150,N_21182,N_24189);
nor U26151 (N_26151,N_24538,N_21905);
or U26152 (N_26152,N_24140,N_21691);
xor U26153 (N_26153,N_22084,N_23798);
or U26154 (N_26154,N_20499,N_24553);
or U26155 (N_26155,N_23697,N_22766);
or U26156 (N_26156,N_22501,N_21545);
or U26157 (N_26157,N_23405,N_20570);
nand U26158 (N_26158,N_20307,N_23589);
and U26159 (N_26159,N_20097,N_24446);
nor U26160 (N_26160,N_24986,N_20894);
xnor U26161 (N_26161,N_22270,N_24564);
or U26162 (N_26162,N_24152,N_22488);
xor U26163 (N_26163,N_24607,N_22859);
xor U26164 (N_26164,N_23645,N_21506);
and U26165 (N_26165,N_22809,N_23569);
xor U26166 (N_26166,N_22061,N_23974);
xnor U26167 (N_26167,N_23905,N_22036);
or U26168 (N_26168,N_23218,N_24262);
and U26169 (N_26169,N_24492,N_21233);
or U26170 (N_26170,N_23561,N_23453);
or U26171 (N_26171,N_20939,N_24873);
nor U26172 (N_26172,N_21390,N_22854);
xor U26173 (N_26173,N_22394,N_24443);
or U26174 (N_26174,N_23288,N_21590);
or U26175 (N_26175,N_24950,N_21741);
and U26176 (N_26176,N_22115,N_24890);
or U26177 (N_26177,N_22065,N_24716);
nor U26178 (N_26178,N_21236,N_20263);
and U26179 (N_26179,N_21005,N_21693);
nand U26180 (N_26180,N_22628,N_23497);
xor U26181 (N_26181,N_22090,N_24322);
nand U26182 (N_26182,N_24622,N_20829);
nor U26183 (N_26183,N_24539,N_21860);
or U26184 (N_26184,N_23359,N_20010);
nor U26185 (N_26185,N_20979,N_24466);
nor U26186 (N_26186,N_21524,N_20759);
and U26187 (N_26187,N_22646,N_20354);
xnor U26188 (N_26188,N_21678,N_22450);
nand U26189 (N_26189,N_24750,N_24045);
or U26190 (N_26190,N_20018,N_21594);
xor U26191 (N_26191,N_20574,N_23846);
and U26192 (N_26192,N_24373,N_24624);
nand U26193 (N_26193,N_23389,N_20201);
nand U26194 (N_26194,N_22779,N_23114);
or U26195 (N_26195,N_20793,N_22493);
and U26196 (N_26196,N_22441,N_20874);
or U26197 (N_26197,N_22562,N_22107);
nor U26198 (N_26198,N_24202,N_20040);
xor U26199 (N_26199,N_23208,N_24822);
xnor U26200 (N_26200,N_22807,N_21284);
nand U26201 (N_26201,N_23776,N_23736);
or U26202 (N_26202,N_22896,N_22004);
nor U26203 (N_26203,N_20661,N_22465);
or U26204 (N_26204,N_24793,N_24221);
nand U26205 (N_26205,N_21388,N_23440);
xnor U26206 (N_26206,N_22749,N_22166);
and U26207 (N_26207,N_22035,N_20568);
nor U26208 (N_26208,N_22266,N_24667);
nor U26209 (N_26209,N_21708,N_22506);
xor U26210 (N_26210,N_22231,N_23142);
or U26211 (N_26211,N_24256,N_22326);
and U26212 (N_26212,N_20606,N_20687);
nand U26213 (N_26213,N_23572,N_22214);
xnor U26214 (N_26214,N_24304,N_21139);
nand U26215 (N_26215,N_21095,N_21014);
nand U26216 (N_26216,N_20938,N_21595);
and U26217 (N_26217,N_24527,N_24314);
xnor U26218 (N_26218,N_23346,N_20281);
nor U26219 (N_26219,N_22416,N_22158);
xnor U26220 (N_26220,N_22812,N_21198);
nand U26221 (N_26221,N_22625,N_22741);
nor U26222 (N_26222,N_20409,N_23371);
nand U26223 (N_26223,N_23349,N_22970);
or U26224 (N_26224,N_24470,N_23386);
nor U26225 (N_26225,N_20411,N_23299);
nor U26226 (N_26226,N_21579,N_20421);
xor U26227 (N_26227,N_23552,N_21563);
xnor U26228 (N_26228,N_22769,N_20542);
and U26229 (N_26229,N_23400,N_24429);
or U26230 (N_26230,N_24104,N_22199);
nor U26231 (N_26231,N_22912,N_21830);
nor U26232 (N_26232,N_20293,N_23354);
and U26233 (N_26233,N_20346,N_22451);
and U26234 (N_26234,N_22835,N_20515);
and U26235 (N_26235,N_24436,N_20763);
nor U26236 (N_26236,N_21508,N_22373);
or U26237 (N_26237,N_24517,N_22934);
or U26238 (N_26238,N_21162,N_20856);
nand U26239 (N_26239,N_22822,N_21383);
nor U26240 (N_26240,N_20387,N_23272);
or U26241 (N_26241,N_23094,N_22303);
or U26242 (N_26242,N_24988,N_24017);
xor U26243 (N_26243,N_21307,N_23350);
and U26244 (N_26244,N_23258,N_24829);
nor U26245 (N_26245,N_21202,N_21160);
nor U26246 (N_26246,N_23843,N_21987);
and U26247 (N_26247,N_24901,N_20089);
and U26248 (N_26248,N_23484,N_24812);
xor U26249 (N_26249,N_21700,N_21885);
xnor U26250 (N_26250,N_22876,N_20265);
and U26251 (N_26251,N_24284,N_21561);
and U26252 (N_26252,N_22837,N_23963);
xnor U26253 (N_26253,N_20519,N_21512);
and U26254 (N_26254,N_23061,N_22333);
nor U26255 (N_26255,N_21743,N_21102);
or U26256 (N_26256,N_23016,N_22117);
nor U26257 (N_26257,N_20746,N_20956);
xnor U26258 (N_26258,N_23596,N_21578);
and U26259 (N_26259,N_22931,N_23148);
and U26260 (N_26260,N_21063,N_23711);
nand U26261 (N_26261,N_20751,N_24729);
nor U26262 (N_26262,N_23231,N_22899);
nand U26263 (N_26263,N_24495,N_23178);
nand U26264 (N_26264,N_21734,N_22063);
nand U26265 (N_26265,N_23626,N_20381);
nand U26266 (N_26266,N_24067,N_20873);
nor U26267 (N_26267,N_23075,N_22584);
xnor U26268 (N_26268,N_21913,N_20615);
and U26269 (N_26269,N_22925,N_21188);
or U26270 (N_26270,N_23731,N_22881);
and U26271 (N_26271,N_24251,N_24057);
xor U26272 (N_26272,N_23252,N_21552);
xor U26273 (N_26273,N_21906,N_20573);
nand U26274 (N_26274,N_22762,N_21115);
nor U26275 (N_26275,N_22945,N_21726);
nand U26276 (N_26276,N_20920,N_24337);
and U26277 (N_26277,N_21592,N_21633);
xnor U26278 (N_26278,N_22134,N_24612);
nor U26279 (N_26279,N_23055,N_24113);
nor U26280 (N_26280,N_21622,N_20965);
and U26281 (N_26281,N_23175,N_21334);
xnor U26282 (N_26282,N_21792,N_20534);
nor U26283 (N_26283,N_23757,N_22961);
and U26284 (N_26284,N_24778,N_21028);
nand U26285 (N_26285,N_23329,N_22355);
nor U26286 (N_26286,N_24032,N_24768);
and U26287 (N_26287,N_20658,N_23632);
nand U26288 (N_26288,N_21431,N_21842);
nor U26289 (N_26289,N_20061,N_20776);
nor U26290 (N_26290,N_23098,N_21020);
and U26291 (N_26291,N_23714,N_20737);
nor U26292 (N_26292,N_23372,N_20055);
nand U26293 (N_26293,N_23990,N_23978);
nand U26294 (N_26294,N_20065,N_24647);
nand U26295 (N_26295,N_22919,N_24765);
and U26296 (N_26296,N_23861,N_24830);
xor U26297 (N_26297,N_21943,N_21826);
or U26298 (N_26298,N_20727,N_22455);
xor U26299 (N_26299,N_21473,N_20891);
or U26300 (N_26300,N_22140,N_22941);
nor U26301 (N_26301,N_24224,N_20707);
nor U26302 (N_26302,N_20397,N_23353);
nor U26303 (N_26303,N_23730,N_21108);
and U26304 (N_26304,N_23777,N_20925);
and U26305 (N_26305,N_22353,N_22707);
xnor U26306 (N_26306,N_21286,N_20388);
and U26307 (N_26307,N_21257,N_22116);
nor U26308 (N_26308,N_20091,N_22918);
and U26309 (N_26309,N_22368,N_23426);
nor U26310 (N_26310,N_24753,N_23516);
and U26311 (N_26311,N_21065,N_22020);
nor U26312 (N_26312,N_20424,N_22953);
xor U26313 (N_26313,N_23425,N_20503);
nand U26314 (N_26314,N_24709,N_22679);
nand U26315 (N_26315,N_21170,N_21656);
nand U26316 (N_26316,N_24827,N_22659);
nor U26317 (N_26317,N_20610,N_22631);
xor U26318 (N_26318,N_21252,N_22665);
and U26319 (N_26319,N_22414,N_20653);
nor U26320 (N_26320,N_21925,N_23709);
xor U26321 (N_26321,N_20115,N_20439);
or U26322 (N_26322,N_21403,N_21703);
nand U26323 (N_26323,N_21581,N_21167);
nand U26324 (N_26324,N_21575,N_23325);
nor U26325 (N_26325,N_22602,N_22573);
xor U26326 (N_26326,N_24034,N_21189);
and U26327 (N_26327,N_21093,N_24724);
and U26328 (N_26328,N_22589,N_20732);
and U26329 (N_26329,N_23831,N_24074);
nor U26330 (N_26330,N_22545,N_21775);
nor U26331 (N_26331,N_22218,N_21158);
xnor U26332 (N_26332,N_23280,N_24205);
and U26333 (N_26333,N_23733,N_22500);
and U26334 (N_26334,N_21888,N_23304);
or U26335 (N_26335,N_23526,N_24493);
xor U26336 (N_26336,N_21727,N_20385);
and U26337 (N_26337,N_24717,N_22290);
nor U26338 (N_26338,N_21245,N_24487);
nand U26339 (N_26339,N_22867,N_24015);
nor U26340 (N_26340,N_21554,N_21505);
xnor U26341 (N_26341,N_23954,N_20174);
or U26342 (N_26342,N_20435,N_21469);
xor U26343 (N_26343,N_22977,N_24653);
and U26344 (N_26344,N_23240,N_24980);
nand U26345 (N_26345,N_24549,N_21718);
or U26346 (N_26346,N_20182,N_21254);
xnor U26347 (N_26347,N_23580,N_20674);
or U26348 (N_26348,N_20043,N_21144);
and U26349 (N_26349,N_20689,N_23316);
nand U26350 (N_26350,N_21268,N_23139);
xnor U26351 (N_26351,N_20529,N_20406);
nor U26352 (N_26352,N_23105,N_24488);
nor U26353 (N_26353,N_22936,N_22761);
or U26354 (N_26354,N_20869,N_22981);
and U26355 (N_26355,N_23265,N_22973);
or U26356 (N_26356,N_21123,N_23478);
and U26357 (N_26357,N_20937,N_20863);
xnor U26358 (N_26358,N_24902,N_21231);
and U26359 (N_26359,N_24790,N_22884);
and U26360 (N_26360,N_21200,N_21515);
or U26361 (N_26361,N_23503,N_23370);
xnor U26362 (N_26362,N_20469,N_20694);
nand U26363 (N_26363,N_22855,N_21049);
nand U26364 (N_26364,N_21306,N_21209);
xnor U26365 (N_26365,N_24984,N_21817);
nor U26366 (N_26366,N_23980,N_21871);
and U26367 (N_26367,N_24381,N_24267);
nor U26368 (N_26368,N_23112,N_23010);
and U26369 (N_26369,N_21191,N_21287);
xnor U26370 (N_26370,N_24430,N_22271);
nor U26371 (N_26371,N_21097,N_24752);
nor U26372 (N_26372,N_20833,N_22873);
nand U26373 (N_26373,N_23224,N_20850);
and U26374 (N_26374,N_20298,N_23382);
and U26375 (N_26375,N_23505,N_22975);
xnor U26376 (N_26376,N_23740,N_24372);
nor U26377 (N_26377,N_24153,N_21556);
nor U26378 (N_26378,N_23468,N_24991);
nor U26379 (N_26379,N_21051,N_20875);
xnor U26380 (N_26380,N_24005,N_20541);
or U26381 (N_26381,N_20482,N_21308);
or U26382 (N_26382,N_22374,N_22475);
and U26383 (N_26383,N_21360,N_23251);
nand U26384 (N_26384,N_20571,N_20834);
nand U26385 (N_26385,N_21802,N_22497);
and U26386 (N_26386,N_21380,N_20399);
and U26387 (N_26387,N_23266,N_22183);
xor U26388 (N_26388,N_23306,N_20360);
or U26389 (N_26389,N_21576,N_23452);
nor U26390 (N_26390,N_22600,N_21974);
nand U26391 (N_26391,N_20788,N_22894);
and U26392 (N_26392,N_22698,N_23470);
and U26393 (N_26393,N_23945,N_23703);
and U26394 (N_26394,N_24578,N_22155);
xor U26395 (N_26395,N_21671,N_24777);
nor U26396 (N_26396,N_22635,N_21818);
or U26397 (N_26397,N_20846,N_23135);
xor U26398 (N_26398,N_24050,N_21125);
nor U26399 (N_26399,N_20880,N_23627);
xnor U26400 (N_26400,N_21015,N_24953);
and U26401 (N_26401,N_24856,N_23271);
xor U26402 (N_26402,N_24018,N_20654);
and U26403 (N_26403,N_20916,N_20715);
xnor U26404 (N_26404,N_21099,N_21052);
or U26405 (N_26405,N_20186,N_23574);
nand U26406 (N_26406,N_24974,N_24361);
nor U26407 (N_26407,N_21738,N_21477);
or U26408 (N_26408,N_24660,N_24170);
or U26409 (N_26409,N_24385,N_24535);
xnor U26410 (N_26410,N_21600,N_24187);
xnor U26411 (N_26411,N_20810,N_24427);
nand U26412 (N_26412,N_21371,N_20622);
or U26413 (N_26413,N_22649,N_22396);
and U26414 (N_26414,N_21914,N_20392);
nor U26415 (N_26415,N_24305,N_22880);
and U26416 (N_26416,N_23655,N_22030);
nand U26417 (N_26417,N_24417,N_20359);
nand U26418 (N_26418,N_20968,N_23490);
and U26419 (N_26419,N_22916,N_20690);
or U26420 (N_26420,N_21810,N_23770);
xnor U26421 (N_26421,N_20117,N_20588);
xnor U26422 (N_26422,N_21890,N_22305);
or U26423 (N_26423,N_24058,N_22949);
nor U26424 (N_26424,N_20560,N_22597);
nand U26425 (N_26425,N_21573,N_22833);
or U26426 (N_26426,N_22224,N_22615);
and U26427 (N_26427,N_23889,N_21178);
nand U26428 (N_26428,N_21463,N_24934);
nand U26429 (N_26429,N_21046,N_22422);
and U26430 (N_26430,N_21539,N_23524);
xnor U26431 (N_26431,N_22343,N_22470);
nand U26432 (N_26432,N_24687,N_21750);
nand U26433 (N_26433,N_22503,N_23841);
xnor U26434 (N_26434,N_23501,N_24697);
nand U26435 (N_26435,N_22875,N_22478);
and U26436 (N_26436,N_21528,N_22015);
xnor U26437 (N_26437,N_23085,N_20011);
or U26438 (N_26438,N_23267,N_22758);
nor U26439 (N_26439,N_22060,N_21513);
or U26440 (N_26440,N_24809,N_21962);
or U26441 (N_26441,N_20078,N_20882);
or U26442 (N_26442,N_22660,N_22669);
nand U26443 (N_26443,N_23712,N_21899);
nor U26444 (N_26444,N_23479,N_24396);
nand U26445 (N_26445,N_22423,N_24855);
and U26446 (N_26446,N_21699,N_23937);
or U26447 (N_26447,N_22418,N_21574);
and U26448 (N_26448,N_24985,N_23883);
or U26449 (N_26449,N_24937,N_22831);
xor U26450 (N_26450,N_23262,N_20369);
and U26451 (N_26451,N_23661,N_23530);
or U26452 (N_26452,N_23716,N_23662);
xor U26453 (N_26453,N_23587,N_21527);
or U26454 (N_26454,N_23086,N_23210);
nor U26455 (N_26455,N_23131,N_20049);
or U26456 (N_26456,N_24244,N_20548);
or U26457 (N_26457,N_20309,N_22777);
and U26458 (N_26458,N_22754,N_21688);
or U26459 (N_26459,N_24626,N_23996);
and U26460 (N_26460,N_20928,N_24876);
or U26461 (N_26461,N_23681,N_23373);
nand U26462 (N_26462,N_23439,N_23480);
nand U26463 (N_26463,N_20959,N_22347);
or U26464 (N_26464,N_24211,N_22474);
nand U26465 (N_26465,N_23932,N_20279);
xor U26466 (N_26466,N_23207,N_20526);
nor U26467 (N_26467,N_21501,N_23109);
and U26468 (N_26468,N_21218,N_22928);
or U26469 (N_26469,N_20495,N_23334);
nand U26470 (N_26470,N_20693,N_20088);
nand U26471 (N_26471,N_24404,N_20978);
or U26472 (N_26472,N_20156,N_24026);
and U26473 (N_26473,N_21025,N_24896);
and U26474 (N_26474,N_21299,N_22397);
and U26475 (N_26475,N_21611,N_20971);
and U26476 (N_26476,N_24945,N_20931);
xnor U26477 (N_26477,N_24555,N_20042);
and U26478 (N_26478,N_24002,N_22765);
nand U26479 (N_26479,N_22507,N_20162);
and U26480 (N_26480,N_23882,N_24301);
and U26481 (N_26481,N_24651,N_20899);
xor U26482 (N_26482,N_24996,N_21702);
xor U26483 (N_26483,N_22695,N_22206);
or U26484 (N_26484,N_21107,N_20434);
nor U26485 (N_26485,N_20999,N_22002);
or U26486 (N_26486,N_24473,N_23691);
or U26487 (N_26487,N_23317,N_20749);
and U26488 (N_26488,N_21309,N_24035);
xnor U26489 (N_26489,N_23390,N_20915);
or U26490 (N_26490,N_20320,N_22105);
nor U26491 (N_26491,N_23421,N_20831);
xnor U26492 (N_26492,N_24749,N_22864);
or U26493 (N_26493,N_21054,N_21300);
nand U26494 (N_26494,N_20121,N_24084);
and U26495 (N_26495,N_20879,N_20890);
nor U26496 (N_26496,N_22543,N_22200);
nand U26497 (N_26497,N_21034,N_22389);
xor U26498 (N_26498,N_24794,N_24652);
nand U26499 (N_26499,N_22476,N_24881);
and U26500 (N_26500,N_21487,N_20302);
nand U26501 (N_26501,N_24608,N_22935);
and U26502 (N_26502,N_23117,N_22265);
nor U26503 (N_26503,N_24344,N_21239);
nor U26504 (N_26504,N_23766,N_20821);
and U26505 (N_26505,N_23570,N_20340);
or U26506 (N_26506,N_21398,N_23800);
xnor U26507 (N_26507,N_22647,N_20045);
and U26508 (N_26508,N_21086,N_23125);
xor U26509 (N_26509,N_22051,N_20647);
or U26510 (N_26510,N_21771,N_22538);
and U26511 (N_26511,N_22186,N_24775);
and U26512 (N_26512,N_22813,N_22221);
and U26513 (N_26513,N_24172,N_21795);
xnor U26514 (N_26514,N_23693,N_21116);
or U26515 (N_26515,N_23435,N_20428);
or U26516 (N_26516,N_20742,N_22637);
xnor U26517 (N_26517,N_21520,N_24159);
xnor U26518 (N_26518,N_20146,N_23344);
or U26519 (N_26519,N_24042,N_23393);
and U26520 (N_26520,N_21935,N_21752);
nand U26521 (N_26521,N_23772,N_23333);
nor U26522 (N_26522,N_22362,N_23830);
xnor U26523 (N_26523,N_23314,N_23639);
nor U26524 (N_26524,N_22078,N_20657);
xor U26525 (N_26525,N_22675,N_23537);
nand U26526 (N_26526,N_22108,N_20860);
xor U26527 (N_26527,N_24471,N_23445);
and U26528 (N_26528,N_21893,N_23023);
xor U26529 (N_26529,N_20592,N_20271);
and U26530 (N_26530,N_20945,N_21467);
nor U26531 (N_26531,N_24302,N_24842);
nand U26532 (N_26532,N_22767,N_21710);
and U26533 (N_26533,N_20811,N_21354);
nor U26534 (N_26534,N_22321,N_21223);
nor U26535 (N_26535,N_23184,N_24921);
or U26536 (N_26536,N_21636,N_20775);
nand U26537 (N_26537,N_20466,N_22552);
nand U26538 (N_26538,N_21548,N_20342);
or U26539 (N_26539,N_23419,N_22385);
nor U26540 (N_26540,N_21630,N_20334);
and U26541 (N_26541,N_20621,N_24510);
or U26542 (N_26542,N_23745,N_21934);
nand U26543 (N_26543,N_22605,N_24944);
xnor U26544 (N_26544,N_24369,N_23925);
and U26545 (N_26545,N_20530,N_24654);
nor U26546 (N_26546,N_20868,N_23509);
nand U26547 (N_26547,N_23773,N_20126);
nand U26548 (N_26548,N_23805,N_21260);
xor U26549 (N_26549,N_24833,N_20446);
xor U26550 (N_26550,N_22708,N_24453);
nand U26551 (N_26551,N_21448,N_23690);
or U26552 (N_26552,N_23064,N_23934);
or U26553 (N_26553,N_23665,N_24387);
or U26554 (N_26554,N_22819,N_24669);
and U26555 (N_26555,N_21675,N_23869);
or U26556 (N_26556,N_24942,N_24020);
and U26557 (N_26557,N_23578,N_23810);
or U26558 (N_26558,N_23002,N_23384);
nor U26559 (N_26559,N_21491,N_22663);
or U26560 (N_26560,N_22308,N_21472);
nor U26561 (N_26561,N_21642,N_24263);
xnor U26562 (N_26562,N_22800,N_20155);
or U26563 (N_26563,N_20599,N_23527);
or U26564 (N_26564,N_24522,N_24849);
nand U26565 (N_26565,N_20160,N_20787);
or U26566 (N_26566,N_21735,N_23200);
nand U26567 (N_26567,N_24218,N_21588);
and U26568 (N_26568,N_21474,N_23868);
nand U26569 (N_26569,N_23245,N_21511);
or U26570 (N_26570,N_20802,N_24526);
nand U26571 (N_26571,N_21834,N_20002);
nand U26572 (N_26572,N_21614,N_24162);
nor U26573 (N_26573,N_20412,N_21659);
nor U26574 (N_26574,N_22776,N_23001);
xnor U26575 (N_26575,N_21159,N_23485);
and U26576 (N_26576,N_24101,N_20418);
nand U26577 (N_26577,N_22720,N_24483);
xnor U26578 (N_26578,N_22797,N_23154);
xor U26579 (N_26579,N_24695,N_20200);
nand U26580 (N_26580,N_20917,N_22121);
or U26581 (N_26581,N_22550,N_22885);
nor U26582 (N_26582,N_24773,N_21042);
xor U26583 (N_26583,N_20349,N_21250);
or U26584 (N_26584,N_22357,N_20614);
xor U26585 (N_26585,N_20960,N_22682);
nand U26586 (N_26586,N_20669,N_24800);
nand U26587 (N_26587,N_21798,N_21064);
or U26588 (N_26588,N_23186,N_20876);
and U26589 (N_26589,N_24913,N_20969);
and U26590 (N_26590,N_20655,N_20362);
or U26591 (N_26591,N_23692,N_20025);
nor U26592 (N_26592,N_22073,N_24055);
or U26593 (N_26593,N_22724,N_20250);
nor U26594 (N_26594,N_23826,N_22043);
nand U26595 (N_26595,N_21357,N_23612);
nand U26596 (N_26596,N_21330,N_24508);
xor U26597 (N_26597,N_20066,N_22581);
and U26598 (N_26598,N_20457,N_21303);
nor U26599 (N_26599,N_23778,N_20688);
nor U26600 (N_26600,N_23725,N_24823);
or U26601 (N_26601,N_23356,N_24161);
xnor U26602 (N_26602,N_21971,N_22787);
nand U26603 (N_26603,N_21435,N_23782);
and U26604 (N_26604,N_22252,N_20037);
or U26605 (N_26605,N_24078,N_21437);
or U26606 (N_26606,N_22295,N_22950);
or U26607 (N_26607,N_21809,N_21801);
nand U26608 (N_26608,N_20059,N_24175);
and U26609 (N_26609,N_21977,N_21542);
nor U26610 (N_26610,N_22400,N_22863);
xnor U26611 (N_26611,N_22856,N_21012);
xor U26612 (N_26612,N_24461,N_24120);
and U26613 (N_26613,N_23481,N_23332);
and U26614 (N_26614,N_22988,N_20348);
and U26615 (N_26615,N_22955,N_23202);
and U26616 (N_26616,N_21044,N_24064);
xnor U26617 (N_26617,N_21615,N_21651);
and U26618 (N_26618,N_20120,N_20600);
and U26619 (N_26619,N_24154,N_24452);
nor U26620 (N_26620,N_21725,N_20538);
and U26621 (N_26621,N_24706,N_21389);
and U26622 (N_26622,N_20267,N_23726);
nor U26623 (N_26623,N_24516,N_24596);
xnor U26624 (N_26624,N_21482,N_23074);
nor U26625 (N_26625,N_21753,N_23173);
nand U26626 (N_26626,N_24282,N_24796);
nand U26627 (N_26627,N_24638,N_24862);
and U26628 (N_26628,N_24614,N_20234);
nand U26629 (N_26629,N_22681,N_20452);
or U26630 (N_26630,N_21960,N_21973);
nor U26631 (N_26631,N_20479,N_24678);
nand U26632 (N_26632,N_24047,N_23228);
nand U26633 (N_26633,N_22028,N_20380);
nor U26634 (N_26634,N_23168,N_22816);
or U26635 (N_26635,N_23144,N_21331);
or U26636 (N_26636,N_24758,N_20611);
nor U26637 (N_26637,N_23194,N_24325);
or U26638 (N_26638,N_21616,N_22249);
and U26639 (N_26639,N_22898,N_23471);
nand U26640 (N_26640,N_21887,N_20950);
or U26641 (N_26641,N_22789,N_20195);
nand U26642 (N_26642,N_24844,N_24853);
or U26643 (N_26643,N_22448,N_20079);
nor U26644 (N_26644,N_22202,N_22824);
and U26645 (N_26645,N_20892,N_24081);
xor U26646 (N_26646,N_24132,N_22175);
nor U26647 (N_26647,N_24060,N_20666);
or U26648 (N_26648,N_20215,N_24964);
nand U26649 (N_26649,N_22588,N_21669);
nor U26650 (N_26650,N_23717,N_24851);
xnor U26651 (N_26651,N_21754,N_21402);
and U26652 (N_26652,N_23121,N_24376);
nor U26653 (N_26653,N_22542,N_23832);
xnor U26654 (N_26654,N_20093,N_20219);
nand U26655 (N_26655,N_20100,N_21634);
and U26656 (N_26656,N_21937,N_21465);
nor U26657 (N_26657,N_20300,N_20590);
xnor U26658 (N_26658,N_21793,N_20819);
and U26659 (N_26659,N_21413,N_22136);
nor U26660 (N_26660,N_24040,N_20695);
and U26661 (N_26661,N_22381,N_20773);
xor U26662 (N_26662,N_20107,N_24384);
nand U26663 (N_26663,N_22799,N_21348);
and U26664 (N_26664,N_22306,N_23442);
and U26665 (N_26665,N_23312,N_21787);
or U26666 (N_26666,N_21855,N_21385);
or U26667 (N_26667,N_23849,N_24474);
or U26668 (N_26668,N_23891,N_24804);
or U26669 (N_26669,N_21557,N_21535);
and U26670 (N_26670,N_21765,N_23540);
and U26671 (N_26671,N_20198,N_22188);
or U26672 (N_26672,N_22037,N_24577);
or U26673 (N_26673,N_24402,N_22435);
nor U26674 (N_26674,N_22328,N_22888);
nand U26675 (N_26675,N_21797,N_23650);
xnor U26676 (N_26676,N_22591,N_20239);
xor U26677 (N_26677,N_21773,N_23753);
nor U26678 (N_26678,N_21850,N_22384);
xor U26679 (N_26679,N_21316,N_23844);
and U26680 (N_26680,N_24353,N_20292);
nand U26681 (N_26681,N_23337,N_24237);
nand U26682 (N_26682,N_22987,N_20163);
nor U26683 (N_26683,N_22377,N_24642);
or U26684 (N_26684,N_20473,N_22042);
nor U26685 (N_26685,N_23041,N_23581);
xor U26686 (N_26686,N_20210,N_24616);
and U26687 (N_26687,N_22668,N_21327);
or U26688 (N_26688,N_22910,N_21214);
nand U26689 (N_26689,N_23137,N_22623);
or U26690 (N_26690,N_24880,N_21195);
nand U26691 (N_26691,N_23965,N_22375);
xor U26692 (N_26692,N_23327,N_20109);
and U26693 (N_26693,N_24479,N_21282);
nand U26694 (N_26694,N_21070,N_23029);
or U26695 (N_26695,N_24933,N_20887);
or U26696 (N_26696,N_22106,N_24231);
or U26697 (N_26697,N_21979,N_24711);
nor U26698 (N_26698,N_21255,N_22201);
nand U26699 (N_26699,N_24311,N_21566);
xor U26700 (N_26700,N_24932,N_23302);
and U26701 (N_26701,N_24781,N_23611);
xnor U26702 (N_26702,N_20576,N_23624);
or U26703 (N_26703,N_22743,N_20311);
nand U26704 (N_26704,N_22018,N_22920);
and U26705 (N_26705,N_24182,N_21213);
nor U26706 (N_26706,N_21989,N_20150);
xnor U26707 (N_26707,N_24445,N_21643);
xor U26708 (N_26708,N_22817,N_23735);
xnor U26709 (N_26709,N_22160,N_24199);
xor U26710 (N_26710,N_20825,N_22774);
and U26711 (N_26711,N_21848,N_20800);
nand U26712 (N_26712,N_24968,N_21204);
nand U26713 (N_26713,N_21953,N_23211);
and U26714 (N_26714,N_24157,N_20253);
xnor U26715 (N_26715,N_21076,N_21519);
xor U26716 (N_26716,N_20248,N_21492);
nand U26717 (N_26717,N_22504,N_20830);
xnor U26718 (N_26718,N_23628,N_22477);
or U26719 (N_26719,N_24277,N_23651);
and U26720 (N_26720,N_24166,N_21018);
and U26721 (N_26721,N_24383,N_24451);
nor U26722 (N_26722,N_22412,N_21288);
nand U26723 (N_26723,N_23964,N_22594);
and U26724 (N_26724,N_21813,N_20245);
xor U26725 (N_26725,N_24259,N_23549);
and U26726 (N_26726,N_24039,N_24165);
or U26727 (N_26727,N_23095,N_23809);
nor U26728 (N_26728,N_21531,N_24967);
and U26729 (N_26729,N_20103,N_22691);
and U26730 (N_26730,N_24343,N_24334);
nand U26731 (N_26731,N_23034,N_22033);
nor U26732 (N_26732,N_21248,N_21460);
nand U26733 (N_26733,N_21466,N_23701);
nor U26734 (N_26734,N_20152,N_21364);
nand U26735 (N_26735,N_20845,N_21225);
and U26736 (N_26736,N_22939,N_22494);
and U26737 (N_26737,N_22818,N_20303);
or U26738 (N_26738,N_21053,N_23613);
nor U26739 (N_26739,N_22638,N_22439);
or U26740 (N_26740,N_23107,N_22164);
xnor U26741 (N_26741,N_22282,N_21138);
and U26742 (N_26742,N_23189,N_23988);
or U26743 (N_26743,N_21247,N_24919);
nor U26744 (N_26744,N_22636,N_21349);
xor U26745 (N_26745,N_21485,N_24808);
xor U26746 (N_26746,N_22672,N_24340);
xnor U26747 (N_26747,N_24358,N_22603);
nand U26748 (N_26748,N_21074,N_23088);
nor U26749 (N_26749,N_21401,N_23320);
xor U26750 (N_26750,N_20861,N_24204);
nor U26751 (N_26751,N_20008,N_21796);
and U26752 (N_26752,N_20308,N_22026);
and U26753 (N_26753,N_22772,N_22298);
xor U26754 (N_26754,N_23785,N_20994);
nor U26755 (N_26755,N_24433,N_20164);
or U26756 (N_26756,N_21132,N_20859);
xor U26757 (N_26757,N_23123,N_20419);
and U26758 (N_26758,N_22232,N_24568);
nor U26759 (N_26759,N_24098,N_21982);
or U26760 (N_26760,N_24066,N_22525);
nor U26761 (N_26761,N_24041,N_21391);
nand U26762 (N_26762,N_23806,N_22486);
xnor U26763 (N_26763,N_23068,N_21039);
nand U26764 (N_26764,N_20699,N_20128);
nand U26765 (N_26765,N_22254,N_21782);
xnor U26766 (N_26766,N_23916,N_23229);
or U26767 (N_26767,N_21628,N_22103);
nand U26768 (N_26768,N_21399,N_24782);
and U26769 (N_26769,N_23987,N_22324);
and U26770 (N_26770,N_24326,N_23686);
nand U26771 (N_26771,N_20436,N_21272);
nor U26772 (N_26772,N_23860,N_23649);
nor U26773 (N_26773,N_23036,N_23009);
nor U26774 (N_26774,N_24836,N_23475);
nand U26775 (N_26775,N_22088,N_24883);
nand U26776 (N_26776,N_21438,N_24197);
or U26777 (N_26777,N_23300,N_20429);
nand U26778 (N_26778,N_21280,N_24630);
xor U26779 (N_26779,N_24805,N_24287);
or U26780 (N_26780,N_23104,N_21772);
or U26781 (N_26781,N_21075,N_21840);
xor U26782 (N_26782,N_23090,N_20750);
nand U26783 (N_26783,N_24597,N_20536);
xnor U26784 (N_26784,N_22411,N_23553);
or U26785 (N_26785,N_22666,N_21894);
nor U26786 (N_26786,N_20132,N_23422);
nand U26787 (N_26787,N_22683,N_20489);
nand U26788 (N_26788,N_21954,N_24185);
nand U26789 (N_26789,N_20116,N_22276);
xnor U26790 (N_26790,N_21026,N_20597);
nor U26791 (N_26791,N_23401,N_22650);
nand U26792 (N_26792,N_20137,N_22370);
nor U26793 (N_26793,N_20315,N_24665);
xor U26794 (N_26794,N_23604,N_20080);
and U26795 (N_26795,N_21361,N_21461);
nand U26796 (N_26796,N_23566,N_20685);
and U26797 (N_26797,N_23000,N_23708);
nor U26798 (N_26798,N_22563,N_20031);
and U26799 (N_26799,N_23124,N_23893);
and U26800 (N_26800,N_21271,N_21963);
nand U26801 (N_26801,N_20020,N_24634);
nor U26802 (N_26802,N_24285,N_20278);
or U26803 (N_26803,N_23120,N_24693);
or U26804 (N_26804,N_23447,N_22734);
xnor U26805 (N_26805,N_24524,N_22732);
xnor U26806 (N_26806,N_21981,N_21931);
nand U26807 (N_26807,N_20852,N_20565);
nand U26808 (N_26808,N_24114,N_23993);
or U26809 (N_26809,N_20324,N_21941);
and U26810 (N_26810,N_20413,N_23789);
nor U26811 (N_26811,N_23616,N_22236);
xnor U26812 (N_26812,N_23909,N_22513);
nand U26813 (N_26813,N_24567,N_21580);
nand U26814 (N_26814,N_23499,N_24386);
or U26815 (N_26815,N_22808,N_22571);
nand U26816 (N_26816,N_22882,N_24754);
nand U26817 (N_26817,N_20365,N_20785);
or U26818 (N_26818,N_22205,N_21392);
nor U26819 (N_26819,N_23877,N_23995);
nand U26820 (N_26820,N_20646,N_23696);
nand U26821 (N_26821,N_21105,N_22651);
nor U26822 (N_26822,N_20758,N_20077);
and U26823 (N_26823,N_24811,N_21488);
or U26824 (N_26824,N_24046,N_24655);
nor U26825 (N_26825,N_22641,N_20500);
and U26826 (N_26826,N_21234,N_23082);
nand U26827 (N_26827,N_22262,N_24519);
or U26828 (N_26828,N_23856,N_20720);
xor U26829 (N_26829,N_23369,N_24562);
nor U26830 (N_26830,N_24770,N_24792);
xor U26831 (N_26831,N_23096,N_24073);
xnor U26832 (N_26832,N_24108,N_22639);
nor U26833 (N_26833,N_20177,N_21744);
nor U26834 (N_26834,N_20798,N_23259);
or U26835 (N_26835,N_24869,N_20555);
or U26836 (N_26836,N_23339,N_24150);
nand U26837 (N_26837,N_22560,N_20724);
nand U26838 (N_26838,N_23103,N_23091);
or U26839 (N_26839,N_24247,N_24745);
xor U26840 (N_26840,N_22406,N_20173);
nand U26841 (N_26841,N_23551,N_21027);
xnor U26842 (N_26842,N_21242,N_23375);
and U26843 (N_26843,N_22279,N_24532);
nor U26844 (N_26844,N_23110,N_22297);
nand U26845 (N_26845,N_24700,N_21854);
xnor U26846 (N_26846,N_23784,N_20352);
and U26847 (N_26847,N_22492,N_23828);
nand U26848 (N_26848,N_23021,N_23588);
nand U26849 (N_26849,N_23670,N_23368);
xnor U26850 (N_26850,N_24583,N_20287);
or U26851 (N_26851,N_21112,N_23775);
or U26852 (N_26852,N_24801,N_22958);
xnor U26853 (N_26853,N_23720,N_20051);
nor U26854 (N_26854,N_20491,N_24083);
nor U26855 (N_26855,N_23364,N_24814);
or U26856 (N_26856,N_21023,N_23179);
nor U26857 (N_26857,N_22067,N_22565);
xor U26858 (N_26858,N_24632,N_22302);
nor U26859 (N_26859,N_24110,N_21811);
xor U26860 (N_26860,N_20171,N_22903);
nor U26861 (N_26861,N_23764,N_22127);
xor U26862 (N_26862,N_24265,N_20335);
nand U26863 (N_26863,N_22780,N_20151);
nor U26864 (N_26864,N_22257,N_23063);
or U26865 (N_26865,N_21320,N_23310);
nand U26866 (N_26866,N_20069,N_23951);
nand U26867 (N_26867,N_20214,N_23512);
and U26868 (N_26868,N_24870,N_21194);
or U26869 (N_26869,N_20898,N_23108);
nand U26870 (N_26870,N_23781,N_21902);
and U26871 (N_26871,N_20185,N_23281);
or U26872 (N_26872,N_23058,N_22185);
nor U26873 (N_26873,N_21617,N_20870);
nor U26874 (N_26874,N_20642,N_21017);
nor U26875 (N_26875,N_22318,N_21904);
nand U26876 (N_26876,N_21104,N_23897);
or U26877 (N_26877,N_24598,N_20855);
or U26878 (N_26878,N_23767,N_21624);
and U26879 (N_26879,N_23946,N_20347);
xor U26880 (N_26880,N_24819,N_20677);
nand U26881 (N_26881,N_23196,N_23072);
nor U26882 (N_26882,N_23285,N_21344);
nor U26883 (N_26883,N_24672,N_21742);
or U26884 (N_26884,N_23858,N_22100);
nor U26885 (N_26885,N_22091,N_20212);
nand U26886 (N_26886,N_21876,N_23151);
or U26887 (N_26887,N_20664,N_23867);
and U26888 (N_26888,N_22438,N_20907);
nand U26889 (N_26889,N_23183,N_20220);
or U26890 (N_26890,N_21770,N_23176);
and U26891 (N_26891,N_24266,N_21667);
nand U26892 (N_26892,N_21530,N_21706);
xor U26893 (N_26893,N_21884,N_24086);
or U26894 (N_26894,N_22579,N_21923);
nor U26895 (N_26895,N_21942,N_20241);
and U26896 (N_26896,N_24171,N_21705);
or U26897 (N_26897,N_21558,N_20587);
nand U26898 (N_26898,N_23837,N_24503);
nand U26899 (N_26899,N_24888,N_21292);
and U26900 (N_26900,N_22334,N_23434);
xnor U26901 (N_26901,N_20222,N_23818);
or U26902 (N_26902,N_22897,N_24245);
xor U26903 (N_26903,N_21341,N_22518);
xnor U26904 (N_26904,N_21004,N_23981);
and U26905 (N_26905,N_22125,N_21301);
nand U26906 (N_26906,N_20583,N_21338);
or U26907 (N_26907,N_20618,N_21665);
nand U26908 (N_26908,N_22686,N_24650);
nor U26909 (N_26909,N_21805,N_22093);
xor U26910 (N_26910,N_22346,N_20488);
nor U26911 (N_26911,N_20068,N_22853);
xor U26912 (N_26912,N_21185,N_20627);
or U26913 (N_26913,N_24328,N_24799);
or U26914 (N_26914,N_23430,N_21529);
and U26915 (N_26915,N_23046,N_24377);
xor U26916 (N_26916,N_23912,N_20764);
nor U26917 (N_26917,N_20092,N_21430);
nand U26918 (N_26918,N_20934,N_23214);
and U26919 (N_26919,N_23290,N_20192);
nor U26920 (N_26920,N_21036,N_24269);
xnor U26921 (N_26921,N_21859,N_20911);
and U26922 (N_26922,N_24795,N_21777);
xnor U26923 (N_26923,N_23718,N_20641);
xor U26924 (N_26924,N_24982,N_20983);
and U26925 (N_26925,N_24571,N_20430);
and U26926 (N_26926,N_22997,N_24414);
or U26927 (N_26927,N_21127,N_24432);
nand U26928 (N_26928,N_23261,N_21369);
nand U26929 (N_26929,N_20358,N_23250);
nor U26930 (N_26930,N_24920,N_22582);
and U26931 (N_26931,N_21807,N_24879);
nor U26932 (N_26932,N_24602,N_24100);
and U26933 (N_26933,N_22906,N_22281);
nor U26934 (N_26934,N_22263,N_24160);
xnor U26935 (N_26935,N_23047,N_23039);
nor U26936 (N_26936,N_23514,N_22393);
xnor U26937 (N_26937,N_23076,N_20511);
nand U26938 (N_26938,N_21148,N_24117);
or U26939 (N_26939,N_23762,N_20878);
nor U26940 (N_26940,N_22081,N_20848);
and U26941 (N_26941,N_20007,N_20376);
nand U26942 (N_26942,N_23345,N_22803);
nand U26943 (N_26943,N_21497,N_24249);
nand U26944 (N_26944,N_22510,N_22751);
nand U26945 (N_26945,N_20896,N_20520);
nand U26946 (N_26946,N_24137,N_23253);
xor U26947 (N_26947,N_24494,N_24515);
or U26948 (N_26948,N_21820,N_24993);
or U26949 (N_26949,N_24409,N_21446);
nand U26950 (N_26950,N_23563,N_23668);
nor U26951 (N_26951,N_24179,N_23308);
nor U26952 (N_26952,N_21002,N_20507);
nor U26953 (N_26953,N_24659,N_22419);
and U26954 (N_26954,N_22655,N_20046);
nor U26955 (N_26955,N_21620,N_23236);
or U26956 (N_26956,N_22508,N_22274);
and U26957 (N_26957,N_20403,N_20124);
or U26958 (N_26958,N_23367,N_23852);
nand U26959 (N_26959,N_23532,N_22287);
or U26960 (N_26960,N_24894,N_22223);
and U26961 (N_26961,N_24956,N_20795);
nand U26962 (N_26962,N_23416,N_20006);
nand U26963 (N_26963,N_20330,N_20672);
and U26964 (N_26964,N_23348,N_23848);
nor U26965 (N_26965,N_23793,N_21873);
nor U26966 (N_26966,N_20885,N_21445);
nand U26967 (N_26967,N_24264,N_20321);
nand U26968 (N_26968,N_24924,N_24016);
xnor U26969 (N_26969,N_24029,N_21658);
or U26970 (N_26970,N_22251,N_24679);
nand U26971 (N_26971,N_22865,N_22212);
and U26972 (N_26972,N_22471,N_21593);
nand U26973 (N_26973,N_22549,N_20645);
nand U26974 (N_26974,N_21067,N_23177);
xor U26975 (N_26975,N_22700,N_20289);
nand U26976 (N_26976,N_24914,N_20131);
xnor U26977 (N_26977,N_24454,N_23443);
or U26978 (N_26978,N_20139,N_24147);
and U26979 (N_26979,N_24718,N_22485);
nor U26980 (N_26980,N_23674,N_20623);
or U26981 (N_26981,N_24601,N_21756);
or U26982 (N_26982,N_24588,N_24188);
nand U26983 (N_26983,N_24972,N_22468);
xor U26984 (N_26984,N_22850,N_23754);
or U26985 (N_26985,N_20299,N_23032);
nand U26986 (N_26986,N_22802,N_20683);
and U26987 (N_26987,N_23165,N_21864);
xnor U26988 (N_26988,N_24498,N_20580);
and U26989 (N_26989,N_22246,N_22327);
nor U26990 (N_26990,N_22645,N_24068);
nor U26991 (N_26991,N_23226,N_20458);
nor U26992 (N_26992,N_23768,N_22079);
or U26993 (N_26993,N_23450,N_20225);
nand U26994 (N_26994,N_24686,N_21635);
nor U26995 (N_26995,N_23038,N_20784);
and U26996 (N_26996,N_23264,N_21944);
and U26997 (N_26997,N_20386,N_22978);
nor U26998 (N_26998,N_23838,N_22156);
or U26999 (N_26999,N_23235,N_23825);
xor U27000 (N_27000,N_22247,N_24540);
nor U27001 (N_27001,N_24629,N_20148);
and U27002 (N_27002,N_21898,N_21518);
nand U27003 (N_27003,N_23523,N_20009);
or U27004 (N_27004,N_21007,N_22250);
xor U27005 (N_27005,N_20849,N_23338);
or U27006 (N_27006,N_24382,N_24210);
and U27007 (N_27007,N_24093,N_22484);
xnor U27008 (N_27008,N_21856,N_23985);
nand U27009 (N_27009,N_22703,N_21915);
or U27010 (N_27010,N_24915,N_20620);
nor U27011 (N_27011,N_20702,N_20552);
nand U27012 (N_27012,N_21673,N_21417);
nand U27013 (N_27013,N_23043,N_20553);
xor U27014 (N_27014,N_22693,N_22314);
nand U27015 (N_27015,N_20314,N_24342);
or U27016 (N_27016,N_22039,N_21995);
xnor U27017 (N_27017,N_24252,N_23307);
nand U27018 (N_27018,N_23269,N_24419);
or U27019 (N_27019,N_21867,N_21961);
or U27020 (N_27020,N_24362,N_20257);
or U27021 (N_27021,N_22742,N_21603);
xor U27022 (N_27022,N_20726,N_22557);
and U27023 (N_27023,N_21462,N_20197);
nand U27024 (N_27024,N_24426,N_21210);
nand U27025 (N_27025,N_24841,N_20063);
and U27026 (N_27026,N_23340,N_23680);
or U27027 (N_27027,N_20697,N_21201);
nor U27028 (N_27028,N_24390,N_24907);
nor U27029 (N_27029,N_23737,N_23102);
nor U27030 (N_27030,N_24692,N_24158);
nor U27031 (N_27031,N_20235,N_23535);
or U27032 (N_27032,N_21451,N_21262);
or U27033 (N_27033,N_22307,N_23145);
nand U27034 (N_27034,N_23153,N_23150);
and U27035 (N_27035,N_20206,N_24288);
xnor U27036 (N_27036,N_21094,N_22944);
and U27037 (N_27037,N_22180,N_21295);
xor U27038 (N_27038,N_20513,N_24444);
nor U27039 (N_27039,N_21350,N_24241);
nor U27040 (N_27040,N_22796,N_24130);
nor U27041 (N_27041,N_22007,N_21901);
xnor U27042 (N_27042,N_23427,N_23994);
nand U27043 (N_27043,N_22132,N_20682);
nor U27044 (N_27044,N_21083,N_23146);
nand U27045 (N_27045,N_22959,N_22322);
nor U27046 (N_27046,N_22994,N_22169);
nor U27047 (N_27047,N_20218,N_20747);
nand U27048 (N_27048,N_23193,N_20718);
nor U27049 (N_27049,N_22869,N_24889);
nor U27050 (N_27050,N_23062,N_24253);
or U27051 (N_27051,N_22730,N_24957);
or U27052 (N_27052,N_24257,N_24413);
and U27053 (N_27053,N_23385,N_22429);
nor U27054 (N_27054,N_24763,N_24878);
nor U27055 (N_27055,N_24609,N_23318);
or U27056 (N_27056,N_24533,N_24591);
nand U27057 (N_27057,N_22114,N_24885);
xnor U27058 (N_27058,N_24728,N_22437);
and U27059 (N_27059,N_23698,N_20105);
nand U27060 (N_27060,N_22162,N_23562);
nor U27061 (N_27061,N_23417,N_23615);
xnor U27062 (N_27062,N_20464,N_23006);
nor U27063 (N_27063,N_24400,N_24071);
or U27064 (N_27064,N_21674,N_21739);
nand U27065 (N_27065,N_23953,N_22123);
nand U27066 (N_27066,N_23411,N_24370);
nand U27067 (N_27067,N_24155,N_20797);
xor U27068 (N_27068,N_20030,N_24813);
and U27069 (N_27069,N_21157,N_21434);
or U27070 (N_27070,N_24688,N_21068);
nor U27071 (N_27071,N_21154,N_22555);
xnor U27072 (N_27072,N_20505,N_21661);
xnor U27073 (N_27073,N_23294,N_24999);
nand U27074 (N_27074,N_24780,N_21682);
and U27075 (N_27075,N_24330,N_20058);
xnor U27076 (N_27076,N_21221,N_22852);
nand U27077 (N_27077,N_22432,N_24545);
and U27078 (N_27078,N_20973,N_21314);
or U27079 (N_27079,N_22120,N_24011);
nand U27080 (N_27080,N_22523,N_24238);
nor U27081 (N_27081,N_20963,N_22226);
or U27082 (N_27082,N_24198,N_21646);
or U27083 (N_27083,N_24599,N_23956);
nand U27084 (N_27084,N_20980,N_24394);
xnor U27085 (N_27085,N_20586,N_21785);
xor U27086 (N_27086,N_20633,N_22760);
and U27087 (N_27087,N_22551,N_21376);
nand U27088 (N_27088,N_20438,N_24085);
xor U27089 (N_27089,N_24798,N_23935);
nor U27090 (N_27090,N_24575,N_23248);
xnor U27091 (N_27091,N_22264,N_24465);
nor U27092 (N_27092,N_23887,N_23796);
xor U27093 (N_27093,N_23763,N_20701);
nor U27094 (N_27094,N_21724,N_21641);
or U27095 (N_27095,N_24410,N_23073);
or U27096 (N_27096,N_22911,N_24019);
xor U27097 (N_27097,N_20743,N_23379);
nand U27098 (N_27098,N_22709,N_20041);
nor U27099 (N_27099,N_20268,N_21464);
or U27100 (N_27100,N_21296,N_21073);
nand U27101 (N_27101,N_20168,N_22688);
xnor U27102 (N_27102,N_20900,N_23278);
xor U27103 (N_27103,N_20158,N_24365);
nor U27104 (N_27104,N_22996,N_22112);
and U27105 (N_27105,N_22892,N_23155);
nand U27106 (N_27106,N_20398,N_23225);
or U27107 (N_27107,N_21737,N_22810);
xor U27108 (N_27108,N_20012,N_20516);
and U27109 (N_27109,N_20443,N_22974);
nand U27110 (N_27110,N_22540,N_22383);
or U27111 (N_27111,N_24146,N_23492);
or U27112 (N_27112,N_24099,N_22240);
xor U27113 (N_27113,N_21173,N_23748);
nor U27114 (N_27114,N_22595,N_21709);
nor U27115 (N_27115,N_22408,N_23113);
nand U27116 (N_27116,N_22378,N_21924);
nor U27117 (N_27117,N_22283,N_20651);
nand U27118 (N_27118,N_20772,N_24222);
xor U27119 (N_27119,N_21150,N_21564);
and U27120 (N_27120,N_21155,N_21395);
xnor U27121 (N_27121,N_22336,N_24976);
nand U27122 (N_27122,N_20957,N_21458);
and U27123 (N_27123,N_22358,N_22031);
and U27124 (N_27124,N_22050,N_21597);
xnor U27125 (N_27125,N_20373,N_20138);
nor U27126 (N_27126,N_23507,N_20276);
and U27127 (N_27127,N_20325,N_20902);
nand U27128 (N_27128,N_23817,N_20024);
nand U27129 (N_27129,N_20562,N_23474);
or U27130 (N_27130,N_20217,N_22719);
and U27131 (N_27131,N_21030,N_21328);
xor U27132 (N_27132,N_22101,N_22991);
xnor U27133 (N_27133,N_21281,N_23898);
xnor U27134 (N_27134,N_21774,N_20753);
or U27135 (N_27135,N_20964,N_22976);
or U27136 (N_27136,N_21677,N_21940);
or U27137 (N_27137,N_20617,N_22498);
xnor U27138 (N_27138,N_24128,N_23755);
nor U27139 (N_27139,N_24219,N_24178);
nand U27140 (N_27140,N_24223,N_22193);
or U27141 (N_27141,N_21419,N_24882);
nand U27142 (N_27142,N_22566,N_22238);
xor U27143 (N_27143,N_20208,N_24619);
nor U27144 (N_27144,N_23873,N_20255);
and U27145 (N_27145,N_23618,N_24332);
xor U27146 (N_27146,N_22146,N_24090);
and U27147 (N_27147,N_22575,N_24604);
nand U27148 (N_27148,N_23864,N_23486);
nand U27149 (N_27149,N_21246,N_23814);
xor U27150 (N_27150,N_20205,N_23621);
nand U27151 (N_27151,N_24579,N_20557);
or U27152 (N_27152,N_23031,N_24590);
xnor U27153 (N_27153,N_23005,N_20809);
and U27154 (N_27154,N_24554,N_24368);
nand U27155 (N_27155,N_24505,N_23498);
or U27156 (N_27156,N_21992,N_23129);
nand U27157 (N_27157,N_20844,N_21788);
or U27158 (N_27158,N_23437,N_23948);
nor U27159 (N_27159,N_23174,N_22574);
and U27160 (N_27160,N_20101,N_24707);
and U27161 (N_27161,N_22047,N_20871);
nand U27162 (N_27162,N_24566,N_22706);
xnor U27163 (N_27163,N_22430,N_24895);
or U27164 (N_27164,N_20270,N_21118);
nand U27165 (N_27165,N_21433,N_20242);
and U27166 (N_27166,N_24779,N_24504);
nor U27167 (N_27167,N_21722,N_20052);
or U27168 (N_27168,N_22331,N_20211);
and U27169 (N_27169,N_22259,N_24180);
nand U27170 (N_27170,N_22386,N_24977);
and U27171 (N_27171,N_22464,N_21238);
nor U27172 (N_27172,N_23441,N_22006);
nand U27173 (N_27173,N_22191,N_24552);
nor U27174 (N_27174,N_20710,N_20981);
nor U27175 (N_27175,N_23922,N_22729);
nor U27176 (N_27176,N_22340,N_20730);
nand U27177 (N_27177,N_24303,N_20675);
nor U27178 (N_27178,N_23399,N_22917);
nand U27179 (N_27179,N_23396,N_20766);
or U27180 (N_27180,N_22792,N_22082);
nand U27181 (N_27181,N_22113,N_20081);
or U27182 (N_27182,N_24810,N_21013);
and U27183 (N_27183,N_22821,N_22452);
nor U27184 (N_27184,N_20236,N_22946);
nor U27185 (N_27185,N_21164,N_21839);
and U27186 (N_27186,N_20524,N_24123);
nand U27187 (N_27187,N_22601,N_20244);
or U27188 (N_27188,N_22891,N_22763);
nand U27189 (N_27189,N_24939,N_20706);
nand U27190 (N_27190,N_22278,N_21972);
or U27191 (N_27191,N_20510,N_22580);
or U27192 (N_27192,N_21040,N_23823);
nand U27193 (N_27193,N_20643,N_21410);
nand U27194 (N_27194,N_21589,N_23705);
or U27195 (N_27195,N_23815,N_24173);
and U27196 (N_27196,N_22499,N_24213);
nand U27197 (N_27197,N_21193,N_23476);
and U27198 (N_27198,N_22522,N_20249);
nand U27199 (N_27199,N_20282,N_20514);
and U27200 (N_27200,N_22782,N_23274);
nand U27201 (N_27201,N_21865,N_21786);
nor U27202 (N_27202,N_21384,N_23313);
xnor U27203 (N_27203,N_21869,N_20734);
nand U27204 (N_27204,N_20071,N_22085);
nor U27205 (N_27205,N_21432,N_20638);
and U27206 (N_27206,N_23859,N_21716);
nand U27207 (N_27207,N_22815,N_20470);
and U27208 (N_27208,N_24111,N_22786);
xnor U27209 (N_27209,N_21240,N_23579);
xnor U27210 (N_27210,N_22041,N_24420);
xor U27211 (N_27211,N_24574,N_23918);
nor U27212 (N_27212,N_24398,N_22131);
or U27213 (N_27213,N_23192,N_20703);
nor U27214 (N_27214,N_23923,N_24525);
and U27215 (N_27215,N_21345,N_23881);
and U27216 (N_27216,N_22887,N_23045);
and U27217 (N_27217,N_23606,N_24708);
xnor U27218 (N_27218,N_21277,N_21181);
or U27219 (N_27219,N_21340,N_22052);
and U27220 (N_27220,N_23558,N_23093);
xor U27221 (N_27221,N_20275,N_23059);
xnor U27222 (N_27222,N_22768,N_24012);
and U27223 (N_27223,N_20601,N_20371);
nor U27224 (N_27224,N_21687,N_22849);
xnor U27225 (N_27225,N_23190,N_22235);
nand U27226 (N_27226,N_20544,N_20537);
nor U27227 (N_27227,N_22388,N_24469);
nor U27228 (N_27228,N_20691,N_20771);
xor U27229 (N_27229,N_21803,N_23130);
nand U27230 (N_27230,N_22753,N_23100);
nor U27231 (N_27231,N_23769,N_22325);
xnor U27232 (N_27232,N_20243,N_22309);
nand U27233 (N_27233,N_21142,N_24448);
nor U27234 (N_27234,N_20338,N_21312);
or U27235 (N_27235,N_24807,N_24542);
nand U27236 (N_27236,N_22182,N_22074);
and U27237 (N_27237,N_20780,N_22356);
nand U27238 (N_27238,N_24725,N_24191);
and U27239 (N_27239,N_21957,N_24824);
nor U27240 (N_27240,N_22773,N_22712);
xor U27241 (N_27241,N_23206,N_22715);
or U27242 (N_27242,N_24958,N_22536);
nor U27243 (N_27243,N_22604,N_20551);
nand U27244 (N_27244,N_21471,N_23854);
nand U27245 (N_27245,N_20535,N_20533);
nor U27246 (N_27246,N_20786,N_24272);
and U27247 (N_27247,N_23171,N_22879);
nor U27248 (N_27248,N_22933,N_22144);
and U27249 (N_27249,N_21343,N_21243);
or U27250 (N_27250,N_21135,N_23664);
nand U27251 (N_27251,N_24671,N_24730);
or U27252 (N_27252,N_22233,N_23614);
xor U27253 (N_27253,N_22401,N_21881);
xnor U27254 (N_27254,N_23469,N_23734);
nand U27255 (N_27255,N_21332,N_20904);
nor U27256 (N_27256,N_21583,N_23608);
xnor U27257 (N_27257,N_21950,N_21454);
nor U27258 (N_27258,N_21352,N_21945);
xor U27259 (N_27259,N_21297,N_23973);
and U27260 (N_27260,N_20857,N_21386);
nor U27261 (N_27261,N_24840,N_20659);
nand U27262 (N_27262,N_24674,N_22609);
and U27263 (N_27263,N_24331,N_22481);
nand U27264 (N_27264,N_23286,N_21610);
xor U27265 (N_27265,N_21450,N_20286);
xnor U27266 (N_27266,N_22220,N_21183);
or U27267 (N_27267,N_21008,N_22755);
nand U27268 (N_27268,N_23957,N_24747);
and U27269 (N_27269,N_21180,N_20652);
nor U27270 (N_27270,N_21666,N_22142);
and U27271 (N_27271,N_24909,N_22995);
nand U27272 (N_27272,N_22962,N_21219);
nor U27273 (N_27273,N_20096,N_24785);
or U27274 (N_27274,N_20604,N_24898);
and U27275 (N_27275,N_21060,N_21747);
nor U27276 (N_27276,N_22445,N_24339);
xnor U27277 (N_27277,N_21533,N_22585);
or U27278 (N_27278,N_23388,N_20976);
nand U27279 (N_27279,N_23305,N_20199);
and U27280 (N_27280,N_23232,N_20295);
nand U27281 (N_27281,N_21072,N_21764);
nor U27282 (N_27282,N_21988,N_20678);
nor U27283 (N_27283,N_20099,N_22312);
and U27284 (N_27284,N_20631,N_21429);
xnor U27285 (N_27285,N_20527,N_20895);
xnor U27286 (N_27286,N_20306,N_23377);
nand U27287 (N_27287,N_21249,N_21728);
nor U27288 (N_27288,N_24022,N_22070);
nor U27289 (N_27289,N_22667,N_21319);
nand U27290 (N_27290,N_22380,N_23066);
and U27291 (N_27291,N_20906,N_23456);
or U27292 (N_27292,N_22387,N_22094);
nor U27293 (N_27293,N_24682,N_22828);
xnor U27294 (N_27294,N_23283,N_22426);
nor U27295 (N_27295,N_23493,N_23908);
and U27296 (N_27296,N_24940,N_20711);
xnor U27297 (N_27297,N_22301,N_21586);
nand U27298 (N_27298,N_22829,N_22443);
nand U27299 (N_27299,N_20770,N_23380);
and U27300 (N_27300,N_23622,N_22129);
nand U27301 (N_27301,N_24354,N_24637);
xnor U27302 (N_27302,N_22718,N_24059);
nand U27303 (N_27303,N_22003,N_24931);
nand U27304 (N_27304,N_24228,N_21800);
xnor U27305 (N_27305,N_22407,N_21373);
and U27306 (N_27306,N_20740,N_22040);
xnor U27307 (N_27307,N_21153,N_23933);
or U27308 (N_27308,N_24313,N_20549);
xnor U27309 (N_27309,N_20328,N_24360);
or U27310 (N_27310,N_24052,N_23220);
and U27311 (N_27311,N_21836,N_24580);
nor U27312 (N_27312,N_20953,N_21582);
or U27313 (N_27313,N_23958,N_22515);
nand U27314 (N_27314,N_22152,N_20966);
and U27315 (N_27315,N_22273,N_22178);
and U27316 (N_27316,N_23862,N_24345);
nor U27317 (N_27317,N_20375,N_23811);
or U27318 (N_27318,N_23620,N_21375);
nand U27319 (N_27319,N_20616,N_22234);
xor U27320 (N_27320,N_20304,N_20468);
or U27321 (N_27321,N_22528,N_24021);
xnor U27322 (N_27322,N_23035,N_21077);
nor U27323 (N_27323,N_21305,N_24871);
and U27324 (N_27324,N_21585,N_21866);
nand U27325 (N_27325,N_20216,N_20076);
xor U27326 (N_27326,N_23682,N_24196);
nor U27327 (N_27327,N_21230,N_21936);
or U27328 (N_27328,N_23599,N_22311);
xor U27329 (N_27329,N_24861,N_23547);
or U27330 (N_27330,N_21427,N_21833);
or U27331 (N_27331,N_22230,N_23982);
or U27332 (N_27332,N_23518,N_23710);
nor U27333 (N_27333,N_22148,N_22521);
nand U27334 (N_27334,N_20098,N_24437);
and U27335 (N_27335,N_24418,N_23111);
and U27336 (N_27336,N_22989,N_20990);
xor U27337 (N_27337,N_23583,N_21031);
nor U27338 (N_27338,N_20812,N_21274);
nor U27339 (N_27339,N_22245,N_23277);
nor U27340 (N_27340,N_21695,N_22556);
xor U27341 (N_27341,N_24643,N_24735);
nor U27342 (N_27342,N_22217,N_20575);
and U27343 (N_27343,N_24694,N_21267);
or U27344 (N_27344,N_22998,N_21672);
and U27345 (N_27345,N_22725,N_22746);
nor U27346 (N_27346,N_23538,N_24959);
nor U27347 (N_27347,N_22071,N_24930);
and U27348 (N_27348,N_22704,N_24892);
or U27349 (N_27349,N_23322,N_20608);
and U27350 (N_27350,N_21428,N_20247);
nor U27351 (N_27351,N_24668,N_23761);
or U27352 (N_27352,N_21346,N_21033);
or U27353 (N_27353,N_20922,N_23984);
nand U27354 (N_27354,N_22339,N_20353);
nor U27355 (N_27355,N_20331,N_20799);
and U27356 (N_27356,N_22956,N_21607);
or U27357 (N_27357,N_22049,N_22640);
nand U27358 (N_27358,N_22572,N_23914);
nand U27359 (N_27359,N_20814,N_22947);
or U27360 (N_27360,N_21821,N_22593);
nor U27361 (N_27361,N_23780,N_24570);
and U27362 (N_27362,N_24439,N_21662);
xor U27363 (N_27363,N_22210,N_23822);
xnor U27364 (N_27364,N_20209,N_20050);
or U27365 (N_27365,N_24388,N_22019);
nand U27366 (N_27366,N_22291,N_21447);
nand U27367 (N_27367,N_22029,N_22926);
nand U27368 (N_27368,N_21509,N_20684);
or U27369 (N_27369,N_22614,N_23319);
xor U27370 (N_27370,N_21175,N_20540);
and U27371 (N_27371,N_21759,N_21259);
xnor U27372 (N_27372,N_24485,N_23303);
nor U27373 (N_27373,N_20628,N_21862);
or U27374 (N_27374,N_24141,N_23816);
xor U27375 (N_27375,N_22128,N_21339);
or U27376 (N_27376,N_20504,N_20035);
nand U27377 (N_27377,N_20060,N_21910);
and U27378 (N_27378,N_22179,N_22277);
or U27379 (N_27379,N_22012,N_21844);
xor U27380 (N_27380,N_21956,N_21900);
nand U27381 (N_27381,N_23391,N_23488);
and U27382 (N_27382,N_20396,N_20865);
nand U27383 (N_27383,N_23673,N_20085);
and U27384 (N_27384,N_20867,N_22095);
nand U27385 (N_27385,N_22930,N_24096);
nand U27386 (N_27386,N_24043,N_21698);
or U27387 (N_27387,N_24321,N_20492);
or U27388 (N_27388,N_21407,N_24788);
nand U27389 (N_27389,N_22171,N_22670);
nor U27390 (N_27390,N_24772,N_22954);
or U27391 (N_27391,N_24689,N_24072);
nand U27392 (N_27392,N_21970,N_21382);
or U27393 (N_27393,N_20184,N_20202);
and U27394 (N_27394,N_20401,N_23276);
nand U27395 (N_27395,N_24458,N_23521);
xnor U27396 (N_27396,N_21366,N_23423);
nand U27397 (N_27397,N_24766,N_24131);
and U27398 (N_27398,N_23792,N_22442);
nor U27399 (N_27399,N_21120,N_21824);
or U27400 (N_27400,N_23291,N_21113);
and U27401 (N_27401,N_23429,N_21226);
nand U27402 (N_27402,N_20927,N_20640);
or U27403 (N_27403,N_22943,N_24089);
xor U27404 (N_27404,N_20828,N_24990);
nor U27405 (N_27405,N_24884,N_21207);
and U27406 (N_27406,N_21324,N_23402);
or U27407 (N_27407,N_23065,N_20837);
nor U27408 (N_27408,N_22759,N_22243);
or U27409 (N_27409,N_21220,N_23779);
nor U27410 (N_27410,N_20393,N_20853);
or U27411 (N_27411,N_21481,N_21378);
nand U27412 (N_27412,N_24070,N_23246);
or U27413 (N_27413,N_24106,N_22172);
and U27414 (N_27414,N_20958,N_23087);
and U27415 (N_27415,N_22764,N_24783);
nand U27416 (N_27416,N_22836,N_23282);
or U27417 (N_27417,N_23820,N_23028);
and U27418 (N_27418,N_21745,N_20803);
xor U27419 (N_27419,N_20149,N_21381);
and U27420 (N_27420,N_24929,N_20933);
and U27421 (N_27421,N_23067,N_20478);
xor U27422 (N_27422,N_23403,N_20761);
xor U27423 (N_27423,N_24513,N_23636);
xnor U27424 (N_27424,N_20017,N_23542);
xor U27425 (N_27425,N_22843,N_23357);
nand U27426 (N_27426,N_22737,N_23336);
nor U27427 (N_27427,N_24787,N_24312);
xor U27428 (N_27428,N_22124,N_21551);
xor U27429 (N_27429,N_22300,N_23534);
xor U27430 (N_27430,N_22338,N_20967);
nand U27431 (N_27431,N_23378,N_23255);
nor U27432 (N_27432,N_20228,N_20717);
nand U27433 (N_27433,N_22690,N_21335);
xnor U27434 (N_27434,N_22126,N_20370);
or U27435 (N_27435,N_21285,N_24275);
xnor U27436 (N_27436,N_24375,N_22215);
xor U27437 (N_27437,N_22622,N_24872);
xor U27438 (N_27438,N_21912,N_23242);
xor U27439 (N_27439,N_23930,N_21555);
and U27440 (N_27440,N_21740,N_22610);
and U27441 (N_27441,N_21721,N_20745);
nand U27442 (N_27442,N_22509,N_20454);
nor U27443 (N_27443,N_22915,N_20461);
xnor U27444 (N_27444,N_23921,N_20607);
nand U27445 (N_27445,N_23855,N_23791);
and U27446 (N_27446,N_22608,N_21757);
and U27447 (N_27447,N_24092,N_23170);
nand U27448 (N_27448,N_21101,N_22554);
and U27449 (N_27449,N_24635,N_20013);
and U27450 (N_27450,N_23465,N_21863);
or U27451 (N_27451,N_24300,N_20893);
or U27452 (N_27452,N_24903,N_24960);
or U27453 (N_27453,N_21278,N_22405);
or U27454 (N_27454,N_21409,N_22350);
and U27455 (N_27455,N_23870,N_21831);
nor U27456 (N_27456,N_22034,N_23565);
or U27457 (N_27457,N_24119,N_22547);
xor U27458 (N_27458,N_21130,N_22851);
nor U27459 (N_27459,N_23374,N_20284);
and U27460 (N_27460,N_24217,N_20665);
and U27461 (N_27461,N_21654,N_21422);
xnor U27462 (N_27462,N_20556,N_22014);
xor U27463 (N_27463,N_23487,N_21411);
and U27464 (N_27464,N_23783,N_23732);
nand U27465 (N_27465,N_23408,N_21577);
and U27466 (N_27466,N_21502,N_23857);
nor U27467 (N_27467,N_23617,N_20663);
or U27468 (N_27468,N_23609,N_23771);
or U27469 (N_27469,N_23827,N_20914);
or U27470 (N_27470,N_24333,N_21917);
or U27471 (N_27471,N_20384,N_23335);
nand U27472 (N_27472,N_20189,N_22066);
and U27473 (N_27473,N_22403,N_20955);
and U27474 (N_27474,N_24620,N_21217);
nor U27475 (N_27475,N_21298,N_22011);
nor U27476 (N_27476,N_24167,N_24613);
xnor U27477 (N_27477,N_24254,N_21650);
and U27478 (N_27478,N_22620,N_20816);
nand U27479 (N_27479,N_23383,N_21780);
nor U27480 (N_27480,N_21781,N_23293);
nand U27481 (N_27481,N_24565,N_22390);
or U27482 (N_27482,N_20705,N_23127);
nand U27483 (N_27483,N_21657,N_22163);
nor U27484 (N_27484,N_23092,N_20986);
or U27485 (N_27485,N_22209,N_23943);
or U27486 (N_27486,N_21769,N_22161);
xor U27487 (N_27487,N_20022,N_22713);
and U27488 (N_27488,N_22434,N_23610);
nor U27489 (N_27489,N_22341,N_23451);
nand U27490 (N_27490,N_21468,N_20989);
nand U27491 (N_27491,N_21370,N_22294);
nand U27492 (N_27492,N_24352,N_20188);
and U27493 (N_27493,N_22184,N_20044);
xor U27494 (N_27494,N_22284,N_23663);
and U27495 (N_27495,N_23554,N_22267);
nor U27496 (N_27496,N_24592,N_24088);
xnor U27497 (N_27497,N_20502,N_21645);
and U27498 (N_27498,N_24270,N_20000);
nor U27499 (N_27499,N_24683,N_24636);
nand U27500 (N_27500,N_24963,N_22051);
xor U27501 (N_27501,N_20499,N_22666);
nor U27502 (N_27502,N_23352,N_22381);
nand U27503 (N_27503,N_23375,N_24838);
nor U27504 (N_27504,N_21753,N_23558);
nand U27505 (N_27505,N_23228,N_20481);
or U27506 (N_27506,N_21004,N_23670);
or U27507 (N_27507,N_21896,N_22694);
or U27508 (N_27508,N_21116,N_23080);
xor U27509 (N_27509,N_23663,N_24421);
and U27510 (N_27510,N_24007,N_24942);
xnor U27511 (N_27511,N_21890,N_22692);
or U27512 (N_27512,N_20823,N_22605);
nand U27513 (N_27513,N_21776,N_24459);
nor U27514 (N_27514,N_23088,N_24387);
nor U27515 (N_27515,N_21318,N_23317);
and U27516 (N_27516,N_22274,N_23886);
or U27517 (N_27517,N_24332,N_20038);
nor U27518 (N_27518,N_21455,N_24505);
or U27519 (N_27519,N_24892,N_23438);
xor U27520 (N_27520,N_22290,N_20682);
nand U27521 (N_27521,N_21666,N_21138);
xnor U27522 (N_27522,N_23171,N_22584);
or U27523 (N_27523,N_20730,N_20053);
and U27524 (N_27524,N_23661,N_21945);
xnor U27525 (N_27525,N_21170,N_24622);
and U27526 (N_27526,N_23282,N_22991);
xor U27527 (N_27527,N_20317,N_22679);
xnor U27528 (N_27528,N_23998,N_20599);
nand U27529 (N_27529,N_24704,N_20290);
xnor U27530 (N_27530,N_23698,N_22549);
or U27531 (N_27531,N_23174,N_22572);
nor U27532 (N_27532,N_21550,N_21032);
nand U27533 (N_27533,N_24723,N_23083);
and U27534 (N_27534,N_21410,N_22633);
xor U27535 (N_27535,N_21792,N_21266);
nor U27536 (N_27536,N_23793,N_24974);
and U27537 (N_27537,N_22274,N_24589);
nor U27538 (N_27538,N_23849,N_22356);
and U27539 (N_27539,N_24683,N_22059);
xnor U27540 (N_27540,N_23620,N_24967);
or U27541 (N_27541,N_24810,N_23715);
xor U27542 (N_27542,N_24505,N_24662);
nand U27543 (N_27543,N_22094,N_22838);
nor U27544 (N_27544,N_20316,N_24785);
xor U27545 (N_27545,N_20045,N_20642);
and U27546 (N_27546,N_24398,N_20441);
nor U27547 (N_27547,N_24010,N_20658);
and U27548 (N_27548,N_24485,N_21466);
nand U27549 (N_27549,N_20426,N_23613);
or U27550 (N_27550,N_22218,N_23582);
or U27551 (N_27551,N_21427,N_23405);
and U27552 (N_27552,N_22202,N_20792);
or U27553 (N_27553,N_22772,N_20899);
nand U27554 (N_27554,N_22734,N_22934);
xor U27555 (N_27555,N_22514,N_20663);
nand U27556 (N_27556,N_22791,N_24937);
and U27557 (N_27557,N_23320,N_21735);
and U27558 (N_27558,N_21332,N_24583);
xor U27559 (N_27559,N_23893,N_24743);
nor U27560 (N_27560,N_21616,N_22309);
xnor U27561 (N_27561,N_22923,N_20947);
or U27562 (N_27562,N_24107,N_21540);
nand U27563 (N_27563,N_21044,N_23205);
or U27564 (N_27564,N_24745,N_21585);
nand U27565 (N_27565,N_20963,N_23121);
and U27566 (N_27566,N_23920,N_24648);
nand U27567 (N_27567,N_20110,N_20725);
nor U27568 (N_27568,N_23317,N_24248);
nand U27569 (N_27569,N_23341,N_22925);
and U27570 (N_27570,N_20913,N_23912);
or U27571 (N_27571,N_21237,N_20567);
xnor U27572 (N_27572,N_21312,N_20367);
or U27573 (N_27573,N_21202,N_24466);
nand U27574 (N_27574,N_24617,N_20543);
and U27575 (N_27575,N_22676,N_20619);
nand U27576 (N_27576,N_21277,N_24460);
and U27577 (N_27577,N_24123,N_23840);
nand U27578 (N_27578,N_22423,N_24079);
nor U27579 (N_27579,N_21901,N_24663);
nand U27580 (N_27580,N_20444,N_23233);
nor U27581 (N_27581,N_22289,N_22715);
and U27582 (N_27582,N_22039,N_24383);
xnor U27583 (N_27583,N_23452,N_22706);
nor U27584 (N_27584,N_23870,N_24740);
or U27585 (N_27585,N_20670,N_20874);
nand U27586 (N_27586,N_24890,N_24325);
and U27587 (N_27587,N_24937,N_23939);
or U27588 (N_27588,N_22531,N_23509);
nor U27589 (N_27589,N_23904,N_20643);
nand U27590 (N_27590,N_22479,N_22507);
or U27591 (N_27591,N_23466,N_22727);
or U27592 (N_27592,N_20962,N_22464);
nor U27593 (N_27593,N_24122,N_23039);
and U27594 (N_27594,N_20346,N_22093);
xor U27595 (N_27595,N_22155,N_23690);
and U27596 (N_27596,N_20159,N_24934);
xnor U27597 (N_27597,N_20613,N_21678);
and U27598 (N_27598,N_21488,N_23695);
or U27599 (N_27599,N_24794,N_22100);
nand U27600 (N_27600,N_22319,N_23627);
nand U27601 (N_27601,N_24102,N_20625);
nand U27602 (N_27602,N_20688,N_22565);
xor U27603 (N_27603,N_20824,N_20858);
nor U27604 (N_27604,N_20767,N_21308);
nor U27605 (N_27605,N_20367,N_20098);
and U27606 (N_27606,N_23921,N_22010);
xnor U27607 (N_27607,N_24978,N_21252);
or U27608 (N_27608,N_20293,N_21000);
nand U27609 (N_27609,N_24071,N_20016);
and U27610 (N_27610,N_22141,N_21762);
nand U27611 (N_27611,N_24153,N_20910);
and U27612 (N_27612,N_22397,N_22448);
nor U27613 (N_27613,N_20568,N_22355);
or U27614 (N_27614,N_21141,N_24888);
nand U27615 (N_27615,N_24697,N_24066);
and U27616 (N_27616,N_20670,N_22955);
or U27617 (N_27617,N_22431,N_24548);
nand U27618 (N_27618,N_24148,N_22936);
or U27619 (N_27619,N_22068,N_23983);
or U27620 (N_27620,N_21670,N_22110);
nand U27621 (N_27621,N_21093,N_20983);
nor U27622 (N_27622,N_24354,N_23443);
and U27623 (N_27623,N_21224,N_21021);
xor U27624 (N_27624,N_24962,N_23527);
nor U27625 (N_27625,N_24228,N_24824);
xor U27626 (N_27626,N_24628,N_22567);
and U27627 (N_27627,N_22787,N_21447);
and U27628 (N_27628,N_24789,N_20920);
nand U27629 (N_27629,N_23661,N_20516);
and U27630 (N_27630,N_22592,N_21844);
nand U27631 (N_27631,N_22802,N_22831);
nand U27632 (N_27632,N_21674,N_22614);
xnor U27633 (N_27633,N_24721,N_24407);
nor U27634 (N_27634,N_22273,N_22897);
or U27635 (N_27635,N_24005,N_24254);
nand U27636 (N_27636,N_20082,N_20997);
nor U27637 (N_27637,N_23958,N_22126);
and U27638 (N_27638,N_22049,N_23653);
xor U27639 (N_27639,N_22505,N_23924);
or U27640 (N_27640,N_22096,N_24686);
nand U27641 (N_27641,N_21346,N_23450);
nor U27642 (N_27642,N_20234,N_21189);
xor U27643 (N_27643,N_22118,N_23421);
nor U27644 (N_27644,N_20360,N_23051);
nand U27645 (N_27645,N_21761,N_24768);
nand U27646 (N_27646,N_22396,N_21680);
and U27647 (N_27647,N_24529,N_24277);
and U27648 (N_27648,N_20542,N_21528);
nand U27649 (N_27649,N_24470,N_23860);
nand U27650 (N_27650,N_21856,N_21914);
xnor U27651 (N_27651,N_22513,N_23863);
and U27652 (N_27652,N_23611,N_21526);
xor U27653 (N_27653,N_22352,N_24810);
and U27654 (N_27654,N_20166,N_23124);
or U27655 (N_27655,N_20044,N_20112);
nand U27656 (N_27656,N_20641,N_21391);
nor U27657 (N_27657,N_20251,N_20284);
nand U27658 (N_27658,N_24738,N_21029);
nand U27659 (N_27659,N_20254,N_22431);
nand U27660 (N_27660,N_21564,N_24168);
nor U27661 (N_27661,N_23869,N_22489);
xor U27662 (N_27662,N_21320,N_22288);
nor U27663 (N_27663,N_21373,N_24951);
xor U27664 (N_27664,N_21360,N_20230);
and U27665 (N_27665,N_23487,N_24792);
or U27666 (N_27666,N_21985,N_22904);
and U27667 (N_27667,N_21388,N_21007);
or U27668 (N_27668,N_20104,N_22397);
or U27669 (N_27669,N_22719,N_20333);
and U27670 (N_27670,N_24244,N_24951);
xnor U27671 (N_27671,N_21591,N_23935);
xnor U27672 (N_27672,N_20034,N_24165);
xor U27673 (N_27673,N_20354,N_22309);
and U27674 (N_27674,N_23570,N_20946);
nor U27675 (N_27675,N_24519,N_24115);
nor U27676 (N_27676,N_21535,N_21700);
xor U27677 (N_27677,N_24878,N_22419);
nand U27678 (N_27678,N_20050,N_22158);
nor U27679 (N_27679,N_22134,N_20144);
xnor U27680 (N_27680,N_20431,N_23334);
xnor U27681 (N_27681,N_21686,N_23171);
nor U27682 (N_27682,N_23634,N_21094);
and U27683 (N_27683,N_24602,N_22845);
or U27684 (N_27684,N_20678,N_22813);
and U27685 (N_27685,N_23619,N_20652);
or U27686 (N_27686,N_20917,N_23621);
or U27687 (N_27687,N_20060,N_20025);
xnor U27688 (N_27688,N_21159,N_22113);
or U27689 (N_27689,N_20065,N_20688);
or U27690 (N_27690,N_20092,N_22392);
and U27691 (N_27691,N_21179,N_24236);
nand U27692 (N_27692,N_23574,N_22991);
nor U27693 (N_27693,N_20187,N_22225);
and U27694 (N_27694,N_20112,N_22532);
or U27695 (N_27695,N_20530,N_23657);
xor U27696 (N_27696,N_20022,N_20709);
nor U27697 (N_27697,N_23107,N_23150);
and U27698 (N_27698,N_23622,N_24997);
nor U27699 (N_27699,N_21172,N_22192);
xnor U27700 (N_27700,N_24160,N_24809);
and U27701 (N_27701,N_24235,N_22467);
or U27702 (N_27702,N_22354,N_22978);
and U27703 (N_27703,N_21320,N_23420);
xnor U27704 (N_27704,N_23636,N_21487);
nand U27705 (N_27705,N_20519,N_21590);
and U27706 (N_27706,N_24221,N_22752);
nor U27707 (N_27707,N_23359,N_22234);
xor U27708 (N_27708,N_24798,N_23400);
nand U27709 (N_27709,N_24003,N_23343);
or U27710 (N_27710,N_21904,N_22512);
nand U27711 (N_27711,N_23560,N_21790);
or U27712 (N_27712,N_22024,N_24747);
xnor U27713 (N_27713,N_22053,N_22769);
xnor U27714 (N_27714,N_23775,N_21588);
nor U27715 (N_27715,N_20191,N_21068);
nor U27716 (N_27716,N_23077,N_23017);
or U27717 (N_27717,N_24443,N_21783);
or U27718 (N_27718,N_24183,N_24408);
nand U27719 (N_27719,N_21228,N_22117);
nor U27720 (N_27720,N_21271,N_24334);
or U27721 (N_27721,N_23323,N_24496);
nor U27722 (N_27722,N_21445,N_21679);
and U27723 (N_27723,N_23225,N_23528);
and U27724 (N_27724,N_20294,N_24188);
xor U27725 (N_27725,N_21734,N_22361);
and U27726 (N_27726,N_23414,N_23197);
or U27727 (N_27727,N_23451,N_24623);
and U27728 (N_27728,N_21326,N_21640);
xnor U27729 (N_27729,N_23238,N_20095);
xnor U27730 (N_27730,N_21085,N_23007);
xnor U27731 (N_27731,N_23053,N_22699);
xor U27732 (N_27732,N_20946,N_23047);
nor U27733 (N_27733,N_22473,N_22091);
nand U27734 (N_27734,N_21282,N_24249);
nand U27735 (N_27735,N_22483,N_24865);
nor U27736 (N_27736,N_24564,N_23471);
nand U27737 (N_27737,N_23021,N_20547);
nand U27738 (N_27738,N_20690,N_20397);
xor U27739 (N_27739,N_22437,N_23743);
xnor U27740 (N_27740,N_21583,N_20326);
xor U27741 (N_27741,N_24753,N_23062);
xnor U27742 (N_27742,N_22184,N_22121);
nand U27743 (N_27743,N_20835,N_22826);
nand U27744 (N_27744,N_20393,N_23570);
nor U27745 (N_27745,N_21676,N_21240);
xor U27746 (N_27746,N_22913,N_23226);
or U27747 (N_27747,N_21001,N_20069);
and U27748 (N_27748,N_20493,N_24344);
or U27749 (N_27749,N_20547,N_21769);
xor U27750 (N_27750,N_24831,N_21329);
nor U27751 (N_27751,N_20027,N_23753);
nor U27752 (N_27752,N_22391,N_24500);
xnor U27753 (N_27753,N_21846,N_23696);
xnor U27754 (N_27754,N_20456,N_22823);
or U27755 (N_27755,N_20599,N_23929);
and U27756 (N_27756,N_22582,N_23474);
or U27757 (N_27757,N_24951,N_20683);
xnor U27758 (N_27758,N_21063,N_23558);
nor U27759 (N_27759,N_24379,N_20857);
nand U27760 (N_27760,N_20063,N_23661);
xnor U27761 (N_27761,N_23774,N_24907);
nor U27762 (N_27762,N_20904,N_21880);
xor U27763 (N_27763,N_21893,N_22952);
nor U27764 (N_27764,N_21128,N_23277);
nor U27765 (N_27765,N_20193,N_20715);
and U27766 (N_27766,N_20454,N_24153);
or U27767 (N_27767,N_20716,N_20745);
nor U27768 (N_27768,N_23233,N_20469);
nor U27769 (N_27769,N_21598,N_20532);
or U27770 (N_27770,N_21719,N_24850);
or U27771 (N_27771,N_23523,N_23313);
xor U27772 (N_27772,N_22494,N_20860);
xor U27773 (N_27773,N_20024,N_24522);
nand U27774 (N_27774,N_24104,N_23996);
and U27775 (N_27775,N_22673,N_23975);
and U27776 (N_27776,N_22592,N_21975);
nand U27777 (N_27777,N_22109,N_21003);
or U27778 (N_27778,N_24404,N_21852);
or U27779 (N_27779,N_22950,N_24503);
nand U27780 (N_27780,N_23917,N_22063);
and U27781 (N_27781,N_23947,N_23260);
xor U27782 (N_27782,N_24454,N_21125);
and U27783 (N_27783,N_22512,N_20795);
nand U27784 (N_27784,N_23110,N_20355);
and U27785 (N_27785,N_20721,N_20473);
xnor U27786 (N_27786,N_22128,N_20715);
nand U27787 (N_27787,N_23630,N_21565);
nor U27788 (N_27788,N_20990,N_24436);
or U27789 (N_27789,N_20220,N_22813);
xor U27790 (N_27790,N_24541,N_21397);
nand U27791 (N_27791,N_23562,N_23027);
or U27792 (N_27792,N_20111,N_21131);
xnor U27793 (N_27793,N_24568,N_21441);
xnor U27794 (N_27794,N_21586,N_23538);
or U27795 (N_27795,N_21793,N_20333);
nand U27796 (N_27796,N_23303,N_20225);
or U27797 (N_27797,N_21860,N_23074);
or U27798 (N_27798,N_24174,N_23774);
or U27799 (N_27799,N_20819,N_22352);
and U27800 (N_27800,N_20351,N_21254);
xnor U27801 (N_27801,N_24185,N_24721);
and U27802 (N_27802,N_22158,N_20397);
nand U27803 (N_27803,N_21972,N_23884);
nor U27804 (N_27804,N_24471,N_21671);
or U27805 (N_27805,N_24270,N_22862);
nor U27806 (N_27806,N_21230,N_24247);
or U27807 (N_27807,N_20369,N_21691);
or U27808 (N_27808,N_24091,N_23400);
nor U27809 (N_27809,N_23255,N_24739);
nor U27810 (N_27810,N_23819,N_24329);
xor U27811 (N_27811,N_20369,N_22143);
nor U27812 (N_27812,N_22433,N_20263);
or U27813 (N_27813,N_21341,N_22971);
nand U27814 (N_27814,N_20422,N_21707);
and U27815 (N_27815,N_24752,N_21941);
or U27816 (N_27816,N_21361,N_21068);
and U27817 (N_27817,N_22837,N_24957);
nor U27818 (N_27818,N_22965,N_20329);
nor U27819 (N_27819,N_24465,N_22703);
xor U27820 (N_27820,N_23859,N_21066);
or U27821 (N_27821,N_21128,N_23114);
nor U27822 (N_27822,N_22784,N_22555);
xor U27823 (N_27823,N_22025,N_23328);
nor U27824 (N_27824,N_23495,N_23277);
xor U27825 (N_27825,N_23282,N_24227);
xnor U27826 (N_27826,N_24766,N_24693);
and U27827 (N_27827,N_22639,N_21224);
xnor U27828 (N_27828,N_23677,N_22478);
nor U27829 (N_27829,N_20574,N_21740);
or U27830 (N_27830,N_22565,N_22630);
nor U27831 (N_27831,N_21128,N_22366);
nor U27832 (N_27832,N_20086,N_21392);
nand U27833 (N_27833,N_24031,N_24897);
nand U27834 (N_27834,N_21592,N_24151);
nor U27835 (N_27835,N_21655,N_21256);
nand U27836 (N_27836,N_24605,N_22238);
nor U27837 (N_27837,N_20157,N_24564);
xnor U27838 (N_27838,N_21301,N_24367);
nor U27839 (N_27839,N_21069,N_23228);
and U27840 (N_27840,N_23357,N_21159);
and U27841 (N_27841,N_20745,N_23953);
xor U27842 (N_27842,N_20671,N_22880);
or U27843 (N_27843,N_22655,N_22002);
and U27844 (N_27844,N_21227,N_23782);
and U27845 (N_27845,N_21638,N_20486);
nor U27846 (N_27846,N_21521,N_23951);
and U27847 (N_27847,N_24641,N_21066);
nor U27848 (N_27848,N_23853,N_22337);
xor U27849 (N_27849,N_22781,N_23083);
or U27850 (N_27850,N_20138,N_23395);
xnor U27851 (N_27851,N_22467,N_21060);
nor U27852 (N_27852,N_22716,N_23637);
or U27853 (N_27853,N_21616,N_23933);
nor U27854 (N_27854,N_22702,N_22425);
and U27855 (N_27855,N_23561,N_21890);
nor U27856 (N_27856,N_23784,N_23322);
and U27857 (N_27857,N_24581,N_21316);
nand U27858 (N_27858,N_23279,N_21543);
and U27859 (N_27859,N_24431,N_23472);
and U27860 (N_27860,N_22318,N_23369);
and U27861 (N_27861,N_24612,N_24866);
or U27862 (N_27862,N_22254,N_21410);
and U27863 (N_27863,N_22967,N_20082);
or U27864 (N_27864,N_22113,N_24042);
and U27865 (N_27865,N_21027,N_24323);
or U27866 (N_27866,N_21661,N_20611);
nor U27867 (N_27867,N_23398,N_23607);
nor U27868 (N_27868,N_20654,N_24032);
xor U27869 (N_27869,N_23368,N_24353);
or U27870 (N_27870,N_24816,N_20673);
or U27871 (N_27871,N_23646,N_24055);
nand U27872 (N_27872,N_22327,N_23614);
nor U27873 (N_27873,N_23665,N_24444);
and U27874 (N_27874,N_21039,N_20977);
or U27875 (N_27875,N_23453,N_21925);
nand U27876 (N_27876,N_21143,N_23162);
and U27877 (N_27877,N_24470,N_24196);
xor U27878 (N_27878,N_24984,N_20170);
nand U27879 (N_27879,N_23604,N_23972);
and U27880 (N_27880,N_24761,N_21312);
nand U27881 (N_27881,N_22662,N_20270);
and U27882 (N_27882,N_22895,N_22529);
nor U27883 (N_27883,N_23231,N_24388);
nor U27884 (N_27884,N_23660,N_22356);
or U27885 (N_27885,N_24826,N_22547);
or U27886 (N_27886,N_21412,N_24097);
and U27887 (N_27887,N_24005,N_23032);
nor U27888 (N_27888,N_22567,N_21372);
nand U27889 (N_27889,N_20317,N_20333);
nor U27890 (N_27890,N_23049,N_20283);
and U27891 (N_27891,N_23013,N_22843);
nand U27892 (N_27892,N_22453,N_23568);
xnor U27893 (N_27893,N_23047,N_20505);
nor U27894 (N_27894,N_20374,N_24668);
nor U27895 (N_27895,N_20555,N_24096);
or U27896 (N_27896,N_24892,N_23463);
nor U27897 (N_27897,N_24831,N_24519);
nand U27898 (N_27898,N_20488,N_21035);
nor U27899 (N_27899,N_23552,N_23939);
nand U27900 (N_27900,N_20605,N_20660);
nor U27901 (N_27901,N_24809,N_22751);
nor U27902 (N_27902,N_20064,N_20388);
nor U27903 (N_27903,N_21376,N_20789);
or U27904 (N_27904,N_22793,N_21567);
or U27905 (N_27905,N_21323,N_23233);
xnor U27906 (N_27906,N_23808,N_21168);
nand U27907 (N_27907,N_21459,N_24444);
nor U27908 (N_27908,N_21518,N_23702);
xor U27909 (N_27909,N_22810,N_20462);
and U27910 (N_27910,N_23094,N_20202);
nor U27911 (N_27911,N_23217,N_23270);
xor U27912 (N_27912,N_20107,N_24288);
nand U27913 (N_27913,N_22888,N_22536);
xnor U27914 (N_27914,N_21904,N_24594);
or U27915 (N_27915,N_23143,N_24586);
or U27916 (N_27916,N_21942,N_23972);
or U27917 (N_27917,N_21346,N_24944);
xor U27918 (N_27918,N_20565,N_23702);
and U27919 (N_27919,N_23603,N_24606);
or U27920 (N_27920,N_24487,N_21429);
xnor U27921 (N_27921,N_20928,N_20247);
nor U27922 (N_27922,N_22150,N_24633);
xnor U27923 (N_27923,N_21733,N_22357);
nor U27924 (N_27924,N_24313,N_20340);
xnor U27925 (N_27925,N_21683,N_22577);
nand U27926 (N_27926,N_21405,N_22200);
nand U27927 (N_27927,N_24798,N_21858);
and U27928 (N_27928,N_23007,N_23230);
or U27929 (N_27929,N_21933,N_22389);
or U27930 (N_27930,N_20697,N_21339);
xor U27931 (N_27931,N_24641,N_20501);
xnor U27932 (N_27932,N_20735,N_22684);
and U27933 (N_27933,N_23087,N_21617);
or U27934 (N_27934,N_22573,N_20139);
xor U27935 (N_27935,N_21081,N_22165);
nor U27936 (N_27936,N_21951,N_23475);
nor U27937 (N_27937,N_24464,N_20809);
nand U27938 (N_27938,N_24893,N_24033);
xor U27939 (N_27939,N_23410,N_23110);
nor U27940 (N_27940,N_21472,N_24104);
or U27941 (N_27941,N_24140,N_21118);
and U27942 (N_27942,N_22636,N_24357);
nand U27943 (N_27943,N_22906,N_22161);
and U27944 (N_27944,N_21556,N_23264);
or U27945 (N_27945,N_21358,N_20498);
xor U27946 (N_27946,N_24717,N_20973);
nor U27947 (N_27947,N_21688,N_20187);
nand U27948 (N_27948,N_20353,N_24845);
and U27949 (N_27949,N_21468,N_23283);
and U27950 (N_27950,N_20943,N_24628);
and U27951 (N_27951,N_21906,N_23529);
nor U27952 (N_27952,N_22926,N_22991);
or U27953 (N_27953,N_20463,N_24028);
nor U27954 (N_27954,N_22241,N_22378);
nor U27955 (N_27955,N_20010,N_21389);
xnor U27956 (N_27956,N_24451,N_24559);
nand U27957 (N_27957,N_20870,N_23156);
nand U27958 (N_27958,N_22029,N_20134);
nor U27959 (N_27959,N_22759,N_24124);
or U27960 (N_27960,N_24474,N_21709);
xor U27961 (N_27961,N_22168,N_21421);
xor U27962 (N_27962,N_21909,N_22922);
and U27963 (N_27963,N_21115,N_20129);
and U27964 (N_27964,N_24524,N_22862);
nor U27965 (N_27965,N_22330,N_24085);
nand U27966 (N_27966,N_21345,N_22984);
xor U27967 (N_27967,N_24083,N_24783);
nand U27968 (N_27968,N_24530,N_24575);
nor U27969 (N_27969,N_23371,N_22223);
xnor U27970 (N_27970,N_23244,N_21395);
or U27971 (N_27971,N_24622,N_24980);
nor U27972 (N_27972,N_24747,N_21644);
nand U27973 (N_27973,N_23158,N_20993);
or U27974 (N_27974,N_20749,N_21170);
xnor U27975 (N_27975,N_22549,N_20366);
xor U27976 (N_27976,N_21817,N_20461);
and U27977 (N_27977,N_21254,N_24258);
or U27978 (N_27978,N_20969,N_22311);
xnor U27979 (N_27979,N_22732,N_21622);
xor U27980 (N_27980,N_22415,N_21665);
xor U27981 (N_27981,N_21373,N_21901);
and U27982 (N_27982,N_20346,N_20286);
or U27983 (N_27983,N_20300,N_21700);
or U27984 (N_27984,N_24902,N_24227);
and U27985 (N_27985,N_23581,N_22683);
or U27986 (N_27986,N_23468,N_22922);
or U27987 (N_27987,N_20998,N_24157);
and U27988 (N_27988,N_23925,N_22975);
nand U27989 (N_27989,N_23815,N_20798);
xnor U27990 (N_27990,N_21762,N_20003);
or U27991 (N_27991,N_20249,N_20473);
nor U27992 (N_27992,N_20672,N_24353);
nor U27993 (N_27993,N_24419,N_24974);
nor U27994 (N_27994,N_23535,N_21443);
xor U27995 (N_27995,N_22114,N_23511);
or U27996 (N_27996,N_22183,N_23474);
nand U27997 (N_27997,N_20956,N_23971);
and U27998 (N_27998,N_21791,N_20096);
xnor U27999 (N_27999,N_23794,N_21173);
xor U28000 (N_28000,N_22504,N_23939);
nand U28001 (N_28001,N_24012,N_24671);
or U28002 (N_28002,N_24025,N_24737);
and U28003 (N_28003,N_20843,N_20135);
nand U28004 (N_28004,N_21448,N_24228);
nor U28005 (N_28005,N_24387,N_24918);
or U28006 (N_28006,N_24932,N_23254);
nor U28007 (N_28007,N_20119,N_21975);
or U28008 (N_28008,N_24761,N_22543);
xnor U28009 (N_28009,N_20214,N_24201);
or U28010 (N_28010,N_21825,N_20420);
nand U28011 (N_28011,N_24115,N_23502);
and U28012 (N_28012,N_24084,N_22324);
nor U28013 (N_28013,N_22958,N_24726);
nor U28014 (N_28014,N_24212,N_22274);
nand U28015 (N_28015,N_20075,N_21403);
nor U28016 (N_28016,N_23531,N_20439);
xnor U28017 (N_28017,N_21011,N_24837);
xor U28018 (N_28018,N_24545,N_21230);
xor U28019 (N_28019,N_24007,N_24486);
and U28020 (N_28020,N_21436,N_21308);
xor U28021 (N_28021,N_23160,N_21754);
xnor U28022 (N_28022,N_21309,N_23818);
and U28023 (N_28023,N_22400,N_24646);
nand U28024 (N_28024,N_24741,N_22466);
or U28025 (N_28025,N_21413,N_21226);
and U28026 (N_28026,N_23749,N_22357);
or U28027 (N_28027,N_23110,N_21632);
xnor U28028 (N_28028,N_22255,N_22749);
or U28029 (N_28029,N_22849,N_23531);
or U28030 (N_28030,N_20831,N_21023);
nor U28031 (N_28031,N_20666,N_20280);
nor U28032 (N_28032,N_20621,N_24611);
or U28033 (N_28033,N_22647,N_21453);
xor U28034 (N_28034,N_23464,N_20100);
nor U28035 (N_28035,N_22587,N_22627);
xnor U28036 (N_28036,N_21487,N_24673);
nand U28037 (N_28037,N_21740,N_23827);
nand U28038 (N_28038,N_21307,N_22222);
and U28039 (N_28039,N_24381,N_21853);
or U28040 (N_28040,N_22820,N_24852);
and U28041 (N_28041,N_23065,N_22022);
nor U28042 (N_28042,N_23329,N_23657);
nor U28043 (N_28043,N_23777,N_24254);
or U28044 (N_28044,N_20644,N_24308);
and U28045 (N_28045,N_22820,N_22590);
xnor U28046 (N_28046,N_20908,N_21317);
nand U28047 (N_28047,N_23380,N_21762);
or U28048 (N_28048,N_22183,N_22393);
or U28049 (N_28049,N_22652,N_21986);
and U28050 (N_28050,N_24499,N_21752);
xor U28051 (N_28051,N_22875,N_20256);
nor U28052 (N_28052,N_24304,N_23151);
nor U28053 (N_28053,N_24818,N_20129);
nor U28054 (N_28054,N_21153,N_20967);
or U28055 (N_28055,N_20773,N_24851);
and U28056 (N_28056,N_22553,N_22347);
nand U28057 (N_28057,N_24623,N_24472);
or U28058 (N_28058,N_20390,N_23170);
and U28059 (N_28059,N_21871,N_20395);
xnor U28060 (N_28060,N_24459,N_21129);
nand U28061 (N_28061,N_24419,N_24761);
nor U28062 (N_28062,N_21525,N_21486);
and U28063 (N_28063,N_20168,N_23468);
nand U28064 (N_28064,N_23187,N_21087);
nor U28065 (N_28065,N_24185,N_20161);
or U28066 (N_28066,N_20028,N_23144);
xnor U28067 (N_28067,N_24309,N_22933);
xor U28068 (N_28068,N_20696,N_22972);
or U28069 (N_28069,N_21539,N_20176);
and U28070 (N_28070,N_22070,N_22350);
nor U28071 (N_28071,N_21727,N_22234);
nor U28072 (N_28072,N_20017,N_20212);
or U28073 (N_28073,N_24335,N_23560);
and U28074 (N_28074,N_22577,N_20795);
and U28075 (N_28075,N_22873,N_22186);
or U28076 (N_28076,N_22217,N_23651);
and U28077 (N_28077,N_23340,N_21714);
nor U28078 (N_28078,N_22856,N_20192);
nand U28079 (N_28079,N_20618,N_21766);
or U28080 (N_28080,N_24217,N_20072);
nor U28081 (N_28081,N_22064,N_20915);
or U28082 (N_28082,N_22605,N_20358);
and U28083 (N_28083,N_20892,N_24698);
and U28084 (N_28084,N_24812,N_20860);
xnor U28085 (N_28085,N_22715,N_20367);
nand U28086 (N_28086,N_20671,N_20126);
nand U28087 (N_28087,N_20021,N_21740);
or U28088 (N_28088,N_22743,N_24381);
xnor U28089 (N_28089,N_21167,N_21729);
nand U28090 (N_28090,N_20427,N_24362);
or U28091 (N_28091,N_20996,N_20071);
nor U28092 (N_28092,N_23119,N_21320);
nor U28093 (N_28093,N_23031,N_23079);
nand U28094 (N_28094,N_21456,N_22920);
xnor U28095 (N_28095,N_24077,N_24226);
and U28096 (N_28096,N_22854,N_20595);
and U28097 (N_28097,N_23296,N_22300);
nand U28098 (N_28098,N_23573,N_20908);
xor U28099 (N_28099,N_23478,N_20999);
and U28100 (N_28100,N_23731,N_24263);
and U28101 (N_28101,N_20549,N_22242);
nand U28102 (N_28102,N_23282,N_22635);
nand U28103 (N_28103,N_23932,N_23022);
and U28104 (N_28104,N_23003,N_21988);
xor U28105 (N_28105,N_20898,N_24150);
and U28106 (N_28106,N_23053,N_23867);
xor U28107 (N_28107,N_23776,N_22219);
or U28108 (N_28108,N_23474,N_22820);
or U28109 (N_28109,N_23162,N_22033);
nor U28110 (N_28110,N_20738,N_21691);
xnor U28111 (N_28111,N_21633,N_24223);
xor U28112 (N_28112,N_20460,N_22162);
xor U28113 (N_28113,N_22613,N_24269);
xor U28114 (N_28114,N_24524,N_22734);
and U28115 (N_28115,N_23719,N_23742);
nand U28116 (N_28116,N_22605,N_22148);
and U28117 (N_28117,N_20842,N_22941);
nor U28118 (N_28118,N_24873,N_24937);
nand U28119 (N_28119,N_21556,N_22027);
or U28120 (N_28120,N_23840,N_21812);
nor U28121 (N_28121,N_21383,N_24227);
and U28122 (N_28122,N_22798,N_20004);
xor U28123 (N_28123,N_21697,N_23459);
xor U28124 (N_28124,N_21606,N_21252);
xor U28125 (N_28125,N_22268,N_23982);
and U28126 (N_28126,N_23442,N_20624);
nor U28127 (N_28127,N_22958,N_22605);
nor U28128 (N_28128,N_22949,N_24329);
xnor U28129 (N_28129,N_24000,N_21525);
xor U28130 (N_28130,N_22126,N_21099);
nand U28131 (N_28131,N_22136,N_23918);
and U28132 (N_28132,N_21905,N_22604);
nand U28133 (N_28133,N_21583,N_22298);
and U28134 (N_28134,N_22586,N_22810);
and U28135 (N_28135,N_24534,N_22915);
nor U28136 (N_28136,N_22872,N_22384);
nand U28137 (N_28137,N_24859,N_24164);
nor U28138 (N_28138,N_20792,N_24888);
nand U28139 (N_28139,N_22194,N_22083);
and U28140 (N_28140,N_20305,N_23579);
nand U28141 (N_28141,N_22819,N_21969);
xor U28142 (N_28142,N_24282,N_22105);
nor U28143 (N_28143,N_23814,N_20790);
or U28144 (N_28144,N_20994,N_24160);
nor U28145 (N_28145,N_22678,N_23980);
nor U28146 (N_28146,N_20221,N_20052);
xnor U28147 (N_28147,N_21269,N_22252);
and U28148 (N_28148,N_23906,N_20021);
xor U28149 (N_28149,N_21041,N_21017);
nand U28150 (N_28150,N_22504,N_22016);
nand U28151 (N_28151,N_22190,N_23225);
or U28152 (N_28152,N_23635,N_20277);
and U28153 (N_28153,N_20561,N_23173);
xor U28154 (N_28154,N_23235,N_21728);
or U28155 (N_28155,N_23746,N_24043);
or U28156 (N_28156,N_22247,N_24012);
xnor U28157 (N_28157,N_22900,N_23284);
and U28158 (N_28158,N_22552,N_22332);
nor U28159 (N_28159,N_23103,N_20338);
xor U28160 (N_28160,N_22970,N_20965);
nor U28161 (N_28161,N_20108,N_22336);
or U28162 (N_28162,N_22342,N_22636);
or U28163 (N_28163,N_23707,N_23085);
xor U28164 (N_28164,N_23098,N_23752);
xnor U28165 (N_28165,N_20855,N_24363);
nand U28166 (N_28166,N_22532,N_21446);
or U28167 (N_28167,N_22304,N_23522);
or U28168 (N_28168,N_24386,N_23137);
nand U28169 (N_28169,N_24258,N_21948);
and U28170 (N_28170,N_24578,N_24271);
nor U28171 (N_28171,N_22133,N_23768);
or U28172 (N_28172,N_21852,N_24492);
and U28173 (N_28173,N_20670,N_20406);
nand U28174 (N_28174,N_22653,N_24950);
or U28175 (N_28175,N_20233,N_20321);
xnor U28176 (N_28176,N_21800,N_21940);
nor U28177 (N_28177,N_21093,N_20299);
nor U28178 (N_28178,N_23302,N_23446);
nor U28179 (N_28179,N_21905,N_24687);
nand U28180 (N_28180,N_24423,N_24193);
or U28181 (N_28181,N_21278,N_23328);
nand U28182 (N_28182,N_20041,N_23330);
and U28183 (N_28183,N_22904,N_22680);
nand U28184 (N_28184,N_23131,N_21204);
nand U28185 (N_28185,N_24728,N_22112);
or U28186 (N_28186,N_21107,N_24701);
nor U28187 (N_28187,N_21855,N_21429);
nor U28188 (N_28188,N_21125,N_20454);
nand U28189 (N_28189,N_20631,N_20084);
or U28190 (N_28190,N_24610,N_24507);
and U28191 (N_28191,N_22825,N_20986);
or U28192 (N_28192,N_21547,N_21772);
nand U28193 (N_28193,N_20986,N_24792);
nand U28194 (N_28194,N_23022,N_24074);
or U28195 (N_28195,N_21938,N_23377);
nor U28196 (N_28196,N_21730,N_20205);
or U28197 (N_28197,N_21290,N_22873);
nor U28198 (N_28198,N_21867,N_23094);
or U28199 (N_28199,N_20670,N_20057);
and U28200 (N_28200,N_24452,N_23975);
nand U28201 (N_28201,N_21946,N_22910);
or U28202 (N_28202,N_24733,N_24856);
and U28203 (N_28203,N_21445,N_20938);
xor U28204 (N_28204,N_20392,N_22326);
xor U28205 (N_28205,N_23838,N_23414);
and U28206 (N_28206,N_21292,N_20337);
xnor U28207 (N_28207,N_21987,N_21544);
xor U28208 (N_28208,N_22690,N_20533);
xor U28209 (N_28209,N_20935,N_22331);
and U28210 (N_28210,N_24940,N_21510);
nand U28211 (N_28211,N_23210,N_23614);
nor U28212 (N_28212,N_22975,N_22375);
or U28213 (N_28213,N_22743,N_21295);
nand U28214 (N_28214,N_21062,N_21177);
nor U28215 (N_28215,N_20987,N_20570);
xor U28216 (N_28216,N_20982,N_20477);
xor U28217 (N_28217,N_22893,N_22027);
nor U28218 (N_28218,N_24534,N_21565);
nor U28219 (N_28219,N_21019,N_23257);
nor U28220 (N_28220,N_20392,N_22129);
or U28221 (N_28221,N_24091,N_24941);
or U28222 (N_28222,N_22546,N_24708);
nand U28223 (N_28223,N_20059,N_23749);
nor U28224 (N_28224,N_21350,N_24671);
xnor U28225 (N_28225,N_24549,N_20412);
xnor U28226 (N_28226,N_21610,N_24392);
nor U28227 (N_28227,N_23626,N_20462);
or U28228 (N_28228,N_20999,N_21746);
nor U28229 (N_28229,N_23156,N_21428);
nor U28230 (N_28230,N_22115,N_23914);
and U28231 (N_28231,N_20732,N_24077);
and U28232 (N_28232,N_21489,N_20719);
nand U28233 (N_28233,N_21499,N_21436);
or U28234 (N_28234,N_24175,N_21509);
nand U28235 (N_28235,N_20069,N_20643);
nor U28236 (N_28236,N_22484,N_21747);
xnor U28237 (N_28237,N_20606,N_21154);
nor U28238 (N_28238,N_21530,N_24083);
and U28239 (N_28239,N_20530,N_23508);
nand U28240 (N_28240,N_20517,N_22583);
nand U28241 (N_28241,N_23426,N_20319);
nor U28242 (N_28242,N_23141,N_20626);
xor U28243 (N_28243,N_20164,N_22985);
xor U28244 (N_28244,N_21728,N_22290);
xor U28245 (N_28245,N_21818,N_24818);
or U28246 (N_28246,N_24853,N_24669);
xnor U28247 (N_28247,N_20570,N_20942);
nand U28248 (N_28248,N_23154,N_21574);
nand U28249 (N_28249,N_23684,N_21089);
nand U28250 (N_28250,N_24497,N_21355);
nand U28251 (N_28251,N_23281,N_24862);
xnor U28252 (N_28252,N_21349,N_21668);
xor U28253 (N_28253,N_22975,N_24526);
or U28254 (N_28254,N_22050,N_21564);
nor U28255 (N_28255,N_24453,N_24861);
nand U28256 (N_28256,N_20514,N_22118);
xor U28257 (N_28257,N_21408,N_23640);
and U28258 (N_28258,N_23807,N_20914);
and U28259 (N_28259,N_22165,N_21825);
xnor U28260 (N_28260,N_20316,N_23265);
and U28261 (N_28261,N_22964,N_22132);
and U28262 (N_28262,N_23693,N_24743);
xor U28263 (N_28263,N_22525,N_21926);
nand U28264 (N_28264,N_22093,N_24987);
nor U28265 (N_28265,N_24898,N_22588);
xor U28266 (N_28266,N_20282,N_21886);
nor U28267 (N_28267,N_22397,N_20466);
nor U28268 (N_28268,N_22975,N_22182);
nor U28269 (N_28269,N_20223,N_22812);
or U28270 (N_28270,N_21597,N_22697);
nand U28271 (N_28271,N_22553,N_20326);
nor U28272 (N_28272,N_24905,N_22113);
xor U28273 (N_28273,N_23359,N_23156);
xor U28274 (N_28274,N_21882,N_23082);
and U28275 (N_28275,N_23369,N_24379);
or U28276 (N_28276,N_20159,N_22722);
and U28277 (N_28277,N_22997,N_20909);
and U28278 (N_28278,N_22570,N_23912);
nand U28279 (N_28279,N_21328,N_20768);
and U28280 (N_28280,N_22781,N_21929);
and U28281 (N_28281,N_24666,N_22852);
nand U28282 (N_28282,N_23017,N_20693);
nor U28283 (N_28283,N_24316,N_22212);
or U28284 (N_28284,N_24139,N_21005);
and U28285 (N_28285,N_20798,N_21276);
or U28286 (N_28286,N_20678,N_23096);
nor U28287 (N_28287,N_24445,N_20076);
and U28288 (N_28288,N_21847,N_23171);
or U28289 (N_28289,N_20331,N_22676);
xor U28290 (N_28290,N_24992,N_20390);
nand U28291 (N_28291,N_21659,N_21851);
xor U28292 (N_28292,N_23136,N_20955);
xor U28293 (N_28293,N_24156,N_22835);
nor U28294 (N_28294,N_21110,N_20925);
or U28295 (N_28295,N_23641,N_24685);
and U28296 (N_28296,N_23996,N_22321);
and U28297 (N_28297,N_24885,N_21784);
or U28298 (N_28298,N_22828,N_20981);
nand U28299 (N_28299,N_23045,N_24819);
or U28300 (N_28300,N_24292,N_24096);
nand U28301 (N_28301,N_23883,N_23273);
or U28302 (N_28302,N_21977,N_23637);
nor U28303 (N_28303,N_24866,N_24510);
nand U28304 (N_28304,N_23409,N_22004);
or U28305 (N_28305,N_21908,N_20500);
nor U28306 (N_28306,N_23828,N_23266);
nand U28307 (N_28307,N_22592,N_21653);
nand U28308 (N_28308,N_24913,N_24560);
and U28309 (N_28309,N_22001,N_24288);
and U28310 (N_28310,N_23166,N_21119);
nand U28311 (N_28311,N_21269,N_22161);
or U28312 (N_28312,N_22589,N_24997);
xor U28313 (N_28313,N_22038,N_22560);
and U28314 (N_28314,N_23695,N_21870);
or U28315 (N_28315,N_20802,N_21751);
and U28316 (N_28316,N_23059,N_20524);
xnor U28317 (N_28317,N_22913,N_21928);
nand U28318 (N_28318,N_24117,N_22701);
nand U28319 (N_28319,N_20200,N_22095);
nor U28320 (N_28320,N_24058,N_22655);
or U28321 (N_28321,N_24451,N_20157);
nor U28322 (N_28322,N_24992,N_24238);
nor U28323 (N_28323,N_21775,N_24425);
nor U28324 (N_28324,N_22538,N_21326);
nand U28325 (N_28325,N_23445,N_21183);
nand U28326 (N_28326,N_23900,N_23550);
and U28327 (N_28327,N_20694,N_22383);
and U28328 (N_28328,N_22213,N_20106);
and U28329 (N_28329,N_20178,N_24134);
nor U28330 (N_28330,N_22877,N_24938);
nor U28331 (N_28331,N_21505,N_20670);
or U28332 (N_28332,N_23577,N_24629);
and U28333 (N_28333,N_24632,N_22557);
xor U28334 (N_28334,N_22814,N_22601);
nor U28335 (N_28335,N_23213,N_20510);
nor U28336 (N_28336,N_24945,N_23930);
nand U28337 (N_28337,N_23112,N_21388);
or U28338 (N_28338,N_24063,N_22954);
nor U28339 (N_28339,N_20046,N_22790);
or U28340 (N_28340,N_24307,N_23136);
or U28341 (N_28341,N_24179,N_20818);
or U28342 (N_28342,N_24463,N_23300);
or U28343 (N_28343,N_20759,N_21878);
and U28344 (N_28344,N_20718,N_21767);
nand U28345 (N_28345,N_21127,N_21226);
and U28346 (N_28346,N_24639,N_21499);
nand U28347 (N_28347,N_20303,N_20313);
xor U28348 (N_28348,N_24724,N_22616);
and U28349 (N_28349,N_22745,N_20568);
nand U28350 (N_28350,N_23626,N_20852);
or U28351 (N_28351,N_24749,N_22330);
nor U28352 (N_28352,N_24166,N_22349);
xor U28353 (N_28353,N_24459,N_21232);
xor U28354 (N_28354,N_24592,N_23541);
xnor U28355 (N_28355,N_21828,N_23371);
or U28356 (N_28356,N_23849,N_22797);
and U28357 (N_28357,N_23892,N_22893);
nand U28358 (N_28358,N_23465,N_23684);
nor U28359 (N_28359,N_22419,N_23988);
xor U28360 (N_28360,N_24678,N_21147);
and U28361 (N_28361,N_22879,N_21293);
or U28362 (N_28362,N_20224,N_24929);
and U28363 (N_28363,N_24994,N_24202);
or U28364 (N_28364,N_22031,N_23838);
and U28365 (N_28365,N_21277,N_24061);
and U28366 (N_28366,N_24052,N_20542);
and U28367 (N_28367,N_23442,N_20007);
xnor U28368 (N_28368,N_24881,N_24587);
or U28369 (N_28369,N_24519,N_23542);
nor U28370 (N_28370,N_21986,N_24294);
nand U28371 (N_28371,N_22337,N_23407);
or U28372 (N_28372,N_23209,N_22465);
or U28373 (N_28373,N_23862,N_23742);
nor U28374 (N_28374,N_23630,N_21547);
or U28375 (N_28375,N_22313,N_22429);
nand U28376 (N_28376,N_22846,N_20356);
nor U28377 (N_28377,N_20554,N_24630);
nor U28378 (N_28378,N_20047,N_24544);
nor U28379 (N_28379,N_23806,N_21361);
nor U28380 (N_28380,N_21182,N_23733);
nor U28381 (N_28381,N_21863,N_23428);
nor U28382 (N_28382,N_23381,N_21479);
xor U28383 (N_28383,N_21573,N_21553);
or U28384 (N_28384,N_22379,N_22648);
nor U28385 (N_28385,N_20330,N_20916);
and U28386 (N_28386,N_20123,N_23413);
or U28387 (N_28387,N_23090,N_24662);
xor U28388 (N_28388,N_21113,N_24497);
nand U28389 (N_28389,N_21806,N_20293);
and U28390 (N_28390,N_22567,N_22295);
xnor U28391 (N_28391,N_23751,N_22490);
xnor U28392 (N_28392,N_20313,N_21576);
nor U28393 (N_28393,N_22060,N_20416);
nand U28394 (N_28394,N_21674,N_20850);
nand U28395 (N_28395,N_22270,N_22427);
and U28396 (N_28396,N_21044,N_24198);
or U28397 (N_28397,N_24982,N_23338);
and U28398 (N_28398,N_21022,N_22784);
and U28399 (N_28399,N_23444,N_21044);
or U28400 (N_28400,N_21706,N_23544);
and U28401 (N_28401,N_23523,N_21488);
or U28402 (N_28402,N_20037,N_20826);
nand U28403 (N_28403,N_20593,N_21897);
xor U28404 (N_28404,N_23037,N_23791);
nor U28405 (N_28405,N_23453,N_21792);
nand U28406 (N_28406,N_20014,N_24917);
nor U28407 (N_28407,N_24716,N_22190);
or U28408 (N_28408,N_21949,N_23005);
xor U28409 (N_28409,N_24274,N_20381);
and U28410 (N_28410,N_20970,N_21517);
and U28411 (N_28411,N_21690,N_24576);
and U28412 (N_28412,N_20035,N_20942);
or U28413 (N_28413,N_23141,N_24383);
nand U28414 (N_28414,N_23554,N_21529);
or U28415 (N_28415,N_22259,N_20738);
nand U28416 (N_28416,N_23811,N_20088);
and U28417 (N_28417,N_23023,N_22823);
xor U28418 (N_28418,N_24617,N_24324);
nand U28419 (N_28419,N_24075,N_22794);
xor U28420 (N_28420,N_24550,N_21244);
xnor U28421 (N_28421,N_22604,N_24752);
and U28422 (N_28422,N_21383,N_22998);
xor U28423 (N_28423,N_22578,N_21431);
xor U28424 (N_28424,N_24966,N_20298);
or U28425 (N_28425,N_24929,N_23397);
or U28426 (N_28426,N_21998,N_20811);
or U28427 (N_28427,N_21676,N_23828);
nand U28428 (N_28428,N_22938,N_20963);
xor U28429 (N_28429,N_22998,N_23634);
and U28430 (N_28430,N_24081,N_24603);
nand U28431 (N_28431,N_21848,N_23454);
or U28432 (N_28432,N_23061,N_20867);
nand U28433 (N_28433,N_24339,N_23516);
and U28434 (N_28434,N_24432,N_21786);
nor U28435 (N_28435,N_22765,N_24927);
and U28436 (N_28436,N_22037,N_22034);
or U28437 (N_28437,N_23519,N_21832);
and U28438 (N_28438,N_24033,N_23234);
nand U28439 (N_28439,N_21173,N_22616);
nand U28440 (N_28440,N_23615,N_20363);
or U28441 (N_28441,N_24091,N_21282);
nand U28442 (N_28442,N_23169,N_23531);
or U28443 (N_28443,N_21626,N_24109);
nand U28444 (N_28444,N_20802,N_22508);
nand U28445 (N_28445,N_23787,N_24025);
or U28446 (N_28446,N_23938,N_24886);
nand U28447 (N_28447,N_22789,N_23057);
or U28448 (N_28448,N_20778,N_23023);
xnor U28449 (N_28449,N_23376,N_22689);
xor U28450 (N_28450,N_23463,N_23128);
or U28451 (N_28451,N_23589,N_23812);
nand U28452 (N_28452,N_20488,N_23779);
or U28453 (N_28453,N_24721,N_23649);
or U28454 (N_28454,N_22367,N_23227);
xor U28455 (N_28455,N_20764,N_21263);
and U28456 (N_28456,N_24225,N_21732);
nor U28457 (N_28457,N_23645,N_21144);
nand U28458 (N_28458,N_21576,N_21324);
and U28459 (N_28459,N_21297,N_20116);
nor U28460 (N_28460,N_23861,N_24977);
nand U28461 (N_28461,N_20314,N_24855);
nor U28462 (N_28462,N_20893,N_20362);
or U28463 (N_28463,N_23706,N_24808);
xor U28464 (N_28464,N_24113,N_20929);
nand U28465 (N_28465,N_24174,N_21490);
nand U28466 (N_28466,N_23399,N_23375);
nor U28467 (N_28467,N_23211,N_20802);
nor U28468 (N_28468,N_24449,N_23175);
xnor U28469 (N_28469,N_20987,N_21070);
or U28470 (N_28470,N_20748,N_23643);
or U28471 (N_28471,N_20139,N_22159);
xor U28472 (N_28472,N_20793,N_24926);
nor U28473 (N_28473,N_22043,N_20381);
or U28474 (N_28474,N_22117,N_20669);
xor U28475 (N_28475,N_22356,N_21166);
and U28476 (N_28476,N_22788,N_20863);
xnor U28477 (N_28477,N_22719,N_24213);
xnor U28478 (N_28478,N_21963,N_21635);
nand U28479 (N_28479,N_23321,N_22530);
nand U28480 (N_28480,N_20100,N_21985);
and U28481 (N_28481,N_20791,N_22935);
and U28482 (N_28482,N_20134,N_22706);
or U28483 (N_28483,N_23695,N_24208);
xor U28484 (N_28484,N_22003,N_22568);
or U28485 (N_28485,N_21215,N_20029);
or U28486 (N_28486,N_23355,N_21088);
nor U28487 (N_28487,N_23417,N_23828);
xnor U28488 (N_28488,N_24069,N_23360);
xnor U28489 (N_28489,N_22117,N_21744);
nand U28490 (N_28490,N_22422,N_24269);
and U28491 (N_28491,N_24236,N_20955);
and U28492 (N_28492,N_20800,N_20516);
nor U28493 (N_28493,N_23295,N_24711);
or U28494 (N_28494,N_22607,N_23177);
xnor U28495 (N_28495,N_22932,N_21979);
or U28496 (N_28496,N_24336,N_20502);
nor U28497 (N_28497,N_24885,N_23308);
or U28498 (N_28498,N_21097,N_23723);
and U28499 (N_28499,N_20571,N_23862);
and U28500 (N_28500,N_21335,N_23113);
nor U28501 (N_28501,N_20487,N_24269);
nand U28502 (N_28502,N_23333,N_22934);
xnor U28503 (N_28503,N_20644,N_24843);
xor U28504 (N_28504,N_20347,N_20282);
or U28505 (N_28505,N_20728,N_22539);
xnor U28506 (N_28506,N_23849,N_21967);
xor U28507 (N_28507,N_22728,N_20949);
xnor U28508 (N_28508,N_24215,N_20903);
nor U28509 (N_28509,N_20891,N_23982);
or U28510 (N_28510,N_24516,N_24427);
xor U28511 (N_28511,N_22868,N_22069);
xnor U28512 (N_28512,N_20084,N_23894);
nor U28513 (N_28513,N_24518,N_20178);
xor U28514 (N_28514,N_20557,N_21102);
or U28515 (N_28515,N_20107,N_23209);
and U28516 (N_28516,N_21016,N_23699);
nor U28517 (N_28517,N_22304,N_23280);
nand U28518 (N_28518,N_22986,N_20287);
nor U28519 (N_28519,N_22831,N_23102);
nand U28520 (N_28520,N_21090,N_23615);
nand U28521 (N_28521,N_20421,N_24350);
and U28522 (N_28522,N_20986,N_23759);
xor U28523 (N_28523,N_21206,N_22807);
nand U28524 (N_28524,N_20423,N_23935);
xor U28525 (N_28525,N_22494,N_22178);
xor U28526 (N_28526,N_21563,N_20378);
nor U28527 (N_28527,N_21716,N_21004);
xnor U28528 (N_28528,N_21317,N_24486);
and U28529 (N_28529,N_23611,N_21637);
or U28530 (N_28530,N_22734,N_22101);
nor U28531 (N_28531,N_21560,N_21868);
or U28532 (N_28532,N_20701,N_21082);
or U28533 (N_28533,N_24745,N_20898);
or U28534 (N_28534,N_20520,N_21705);
xnor U28535 (N_28535,N_23027,N_21305);
nand U28536 (N_28536,N_24504,N_22393);
or U28537 (N_28537,N_24823,N_21472);
xnor U28538 (N_28538,N_21270,N_24032);
nor U28539 (N_28539,N_24153,N_22086);
xor U28540 (N_28540,N_20357,N_20157);
nand U28541 (N_28541,N_23937,N_23141);
or U28542 (N_28542,N_22892,N_24432);
xnor U28543 (N_28543,N_21997,N_20181);
xor U28544 (N_28544,N_23559,N_21871);
nand U28545 (N_28545,N_21627,N_23572);
nand U28546 (N_28546,N_20550,N_24941);
or U28547 (N_28547,N_20035,N_22680);
nor U28548 (N_28548,N_20659,N_21636);
nor U28549 (N_28549,N_23617,N_24458);
xor U28550 (N_28550,N_23330,N_21981);
xor U28551 (N_28551,N_23470,N_22718);
or U28552 (N_28552,N_21692,N_21930);
xnor U28553 (N_28553,N_24598,N_21735);
xor U28554 (N_28554,N_21038,N_21376);
nor U28555 (N_28555,N_23897,N_22576);
nand U28556 (N_28556,N_22427,N_21274);
nand U28557 (N_28557,N_20423,N_22161);
nand U28558 (N_28558,N_22855,N_23998);
nor U28559 (N_28559,N_24681,N_21771);
xnor U28560 (N_28560,N_24624,N_22256);
and U28561 (N_28561,N_22821,N_23271);
nand U28562 (N_28562,N_22069,N_21264);
xnor U28563 (N_28563,N_21769,N_24107);
nand U28564 (N_28564,N_23724,N_21848);
nand U28565 (N_28565,N_23241,N_24046);
xor U28566 (N_28566,N_21673,N_24388);
or U28567 (N_28567,N_21558,N_22460);
and U28568 (N_28568,N_20496,N_22662);
or U28569 (N_28569,N_21917,N_24931);
and U28570 (N_28570,N_22530,N_23445);
or U28571 (N_28571,N_20044,N_24191);
nor U28572 (N_28572,N_20835,N_23496);
and U28573 (N_28573,N_23830,N_21551);
nand U28574 (N_28574,N_23537,N_20709);
or U28575 (N_28575,N_21177,N_21411);
nand U28576 (N_28576,N_22175,N_23564);
or U28577 (N_28577,N_23595,N_21498);
xor U28578 (N_28578,N_21325,N_24190);
xnor U28579 (N_28579,N_23386,N_22863);
nor U28580 (N_28580,N_20198,N_24643);
and U28581 (N_28581,N_20031,N_23726);
nor U28582 (N_28582,N_22304,N_23294);
nand U28583 (N_28583,N_23054,N_22531);
xor U28584 (N_28584,N_22591,N_20460);
and U28585 (N_28585,N_24645,N_20784);
nor U28586 (N_28586,N_24335,N_20708);
nand U28587 (N_28587,N_20133,N_21277);
and U28588 (N_28588,N_24030,N_23497);
xnor U28589 (N_28589,N_24149,N_24787);
xnor U28590 (N_28590,N_22795,N_23521);
xnor U28591 (N_28591,N_23421,N_20800);
nand U28592 (N_28592,N_23582,N_24705);
xnor U28593 (N_28593,N_21582,N_22096);
or U28594 (N_28594,N_22260,N_23871);
and U28595 (N_28595,N_21729,N_23381);
nand U28596 (N_28596,N_22489,N_23411);
and U28597 (N_28597,N_21113,N_23627);
xnor U28598 (N_28598,N_22381,N_23955);
and U28599 (N_28599,N_20667,N_22663);
or U28600 (N_28600,N_24547,N_21525);
and U28601 (N_28601,N_20767,N_24943);
or U28602 (N_28602,N_21142,N_20604);
nor U28603 (N_28603,N_22202,N_23277);
nor U28604 (N_28604,N_21174,N_23216);
nand U28605 (N_28605,N_22949,N_24612);
xor U28606 (N_28606,N_20643,N_23568);
nand U28607 (N_28607,N_21319,N_23617);
nand U28608 (N_28608,N_22479,N_22692);
or U28609 (N_28609,N_23118,N_20980);
and U28610 (N_28610,N_24715,N_22434);
or U28611 (N_28611,N_20676,N_20235);
or U28612 (N_28612,N_20005,N_23974);
xnor U28613 (N_28613,N_21083,N_21135);
xnor U28614 (N_28614,N_23702,N_24231);
and U28615 (N_28615,N_22005,N_24577);
or U28616 (N_28616,N_20718,N_23726);
and U28617 (N_28617,N_22371,N_20172);
nor U28618 (N_28618,N_20140,N_22434);
or U28619 (N_28619,N_23402,N_22654);
or U28620 (N_28620,N_24545,N_20542);
nor U28621 (N_28621,N_20241,N_23191);
xnor U28622 (N_28622,N_24505,N_24343);
or U28623 (N_28623,N_21631,N_24818);
or U28624 (N_28624,N_22760,N_22306);
or U28625 (N_28625,N_23137,N_22868);
or U28626 (N_28626,N_21164,N_23658);
xnor U28627 (N_28627,N_24423,N_23860);
nor U28628 (N_28628,N_24538,N_23190);
xnor U28629 (N_28629,N_23687,N_24720);
nand U28630 (N_28630,N_23694,N_23679);
or U28631 (N_28631,N_20478,N_23273);
nor U28632 (N_28632,N_23550,N_24025);
nor U28633 (N_28633,N_21914,N_23027);
xor U28634 (N_28634,N_21085,N_20975);
xnor U28635 (N_28635,N_22705,N_22878);
and U28636 (N_28636,N_24091,N_20945);
nor U28637 (N_28637,N_20029,N_21657);
nor U28638 (N_28638,N_21126,N_22645);
nand U28639 (N_28639,N_24537,N_20586);
and U28640 (N_28640,N_24194,N_24189);
nand U28641 (N_28641,N_21042,N_21490);
and U28642 (N_28642,N_23755,N_20195);
nor U28643 (N_28643,N_22251,N_22410);
nand U28644 (N_28644,N_20833,N_20277);
or U28645 (N_28645,N_20831,N_20594);
nor U28646 (N_28646,N_24308,N_24940);
nand U28647 (N_28647,N_20959,N_23353);
nand U28648 (N_28648,N_22041,N_20241);
or U28649 (N_28649,N_23611,N_24067);
nand U28650 (N_28650,N_23751,N_22521);
nor U28651 (N_28651,N_23766,N_22915);
xnor U28652 (N_28652,N_22250,N_20688);
xor U28653 (N_28653,N_22819,N_20587);
or U28654 (N_28654,N_21132,N_23994);
xnor U28655 (N_28655,N_20482,N_22070);
nor U28656 (N_28656,N_21904,N_22221);
nand U28657 (N_28657,N_21624,N_22125);
nor U28658 (N_28658,N_21843,N_22227);
and U28659 (N_28659,N_22692,N_23714);
nor U28660 (N_28660,N_21971,N_20040);
nand U28661 (N_28661,N_22987,N_22796);
xnor U28662 (N_28662,N_23378,N_21519);
and U28663 (N_28663,N_24309,N_20533);
nand U28664 (N_28664,N_23661,N_22674);
or U28665 (N_28665,N_21474,N_24691);
and U28666 (N_28666,N_20624,N_23549);
and U28667 (N_28667,N_22812,N_24593);
nor U28668 (N_28668,N_22189,N_22601);
and U28669 (N_28669,N_21404,N_20732);
xor U28670 (N_28670,N_22737,N_21562);
nand U28671 (N_28671,N_23195,N_24380);
nor U28672 (N_28672,N_24866,N_22221);
and U28673 (N_28673,N_20054,N_22808);
xnor U28674 (N_28674,N_23088,N_21555);
and U28675 (N_28675,N_22315,N_22238);
nand U28676 (N_28676,N_24323,N_22372);
and U28677 (N_28677,N_22034,N_20010);
or U28678 (N_28678,N_21309,N_20630);
and U28679 (N_28679,N_23545,N_24892);
nor U28680 (N_28680,N_23361,N_22973);
nor U28681 (N_28681,N_21140,N_24209);
or U28682 (N_28682,N_22791,N_24970);
or U28683 (N_28683,N_24844,N_24547);
or U28684 (N_28684,N_22296,N_22678);
nor U28685 (N_28685,N_24246,N_24460);
and U28686 (N_28686,N_24347,N_23231);
or U28687 (N_28687,N_24024,N_24616);
xnor U28688 (N_28688,N_21276,N_21932);
nor U28689 (N_28689,N_22416,N_20118);
xnor U28690 (N_28690,N_21174,N_23664);
or U28691 (N_28691,N_23014,N_21008);
and U28692 (N_28692,N_24883,N_21378);
nand U28693 (N_28693,N_24817,N_21212);
and U28694 (N_28694,N_20428,N_23009);
or U28695 (N_28695,N_24211,N_23780);
nand U28696 (N_28696,N_21208,N_22272);
xor U28697 (N_28697,N_24319,N_21487);
nand U28698 (N_28698,N_23607,N_24242);
and U28699 (N_28699,N_21604,N_21591);
nand U28700 (N_28700,N_23603,N_23723);
nand U28701 (N_28701,N_24902,N_20985);
xor U28702 (N_28702,N_20255,N_20268);
nand U28703 (N_28703,N_21933,N_23096);
xor U28704 (N_28704,N_22224,N_23813);
xor U28705 (N_28705,N_20563,N_20497);
and U28706 (N_28706,N_23583,N_23736);
or U28707 (N_28707,N_22243,N_23469);
and U28708 (N_28708,N_21507,N_21145);
and U28709 (N_28709,N_24561,N_22974);
nand U28710 (N_28710,N_20159,N_24453);
or U28711 (N_28711,N_21797,N_21382);
xor U28712 (N_28712,N_23476,N_21192);
or U28713 (N_28713,N_21010,N_20844);
and U28714 (N_28714,N_23599,N_24558);
nand U28715 (N_28715,N_21271,N_22329);
nand U28716 (N_28716,N_24910,N_20457);
nand U28717 (N_28717,N_20373,N_20871);
nor U28718 (N_28718,N_22494,N_24661);
nand U28719 (N_28719,N_24390,N_23671);
xor U28720 (N_28720,N_22010,N_24286);
or U28721 (N_28721,N_22249,N_20035);
nand U28722 (N_28722,N_23865,N_23155);
and U28723 (N_28723,N_22026,N_21652);
xor U28724 (N_28724,N_21538,N_21265);
xor U28725 (N_28725,N_24842,N_22691);
nor U28726 (N_28726,N_21610,N_23842);
nand U28727 (N_28727,N_24728,N_23835);
nor U28728 (N_28728,N_20540,N_20358);
nor U28729 (N_28729,N_20031,N_20872);
or U28730 (N_28730,N_24440,N_21600);
nor U28731 (N_28731,N_21544,N_20546);
or U28732 (N_28732,N_23579,N_22370);
and U28733 (N_28733,N_23150,N_24415);
xnor U28734 (N_28734,N_22618,N_22384);
xor U28735 (N_28735,N_20502,N_22706);
nand U28736 (N_28736,N_23361,N_22023);
or U28737 (N_28737,N_22731,N_22031);
xor U28738 (N_28738,N_24858,N_22038);
and U28739 (N_28739,N_21933,N_24653);
or U28740 (N_28740,N_20742,N_20024);
and U28741 (N_28741,N_21032,N_20017);
nand U28742 (N_28742,N_23763,N_21918);
and U28743 (N_28743,N_23852,N_24389);
nor U28744 (N_28744,N_21434,N_23007);
and U28745 (N_28745,N_22711,N_24861);
nand U28746 (N_28746,N_24587,N_21224);
or U28747 (N_28747,N_20797,N_22368);
or U28748 (N_28748,N_22801,N_23833);
or U28749 (N_28749,N_23646,N_22616);
nand U28750 (N_28750,N_23870,N_21191);
nand U28751 (N_28751,N_21611,N_20251);
xor U28752 (N_28752,N_24464,N_20812);
or U28753 (N_28753,N_20852,N_21831);
xor U28754 (N_28754,N_24447,N_23673);
or U28755 (N_28755,N_24877,N_20188);
xor U28756 (N_28756,N_24627,N_24977);
nor U28757 (N_28757,N_20038,N_24859);
or U28758 (N_28758,N_22026,N_23486);
xnor U28759 (N_28759,N_22026,N_23779);
and U28760 (N_28760,N_24507,N_21950);
nand U28761 (N_28761,N_22050,N_23002);
and U28762 (N_28762,N_23192,N_21582);
or U28763 (N_28763,N_21331,N_22155);
nor U28764 (N_28764,N_23890,N_22619);
nor U28765 (N_28765,N_22205,N_20292);
and U28766 (N_28766,N_21625,N_22590);
or U28767 (N_28767,N_21556,N_21756);
and U28768 (N_28768,N_22405,N_23711);
nand U28769 (N_28769,N_23005,N_23336);
nor U28770 (N_28770,N_23311,N_22329);
nor U28771 (N_28771,N_22901,N_23458);
or U28772 (N_28772,N_24583,N_22714);
or U28773 (N_28773,N_22737,N_23019);
and U28774 (N_28774,N_24080,N_23022);
or U28775 (N_28775,N_24235,N_20412);
and U28776 (N_28776,N_21291,N_23967);
and U28777 (N_28777,N_24960,N_22852);
or U28778 (N_28778,N_24738,N_22096);
nor U28779 (N_28779,N_22975,N_23008);
nand U28780 (N_28780,N_20785,N_23471);
or U28781 (N_28781,N_24416,N_20037);
or U28782 (N_28782,N_20557,N_22807);
or U28783 (N_28783,N_24983,N_23484);
nand U28784 (N_28784,N_21221,N_24077);
or U28785 (N_28785,N_22392,N_20137);
nand U28786 (N_28786,N_22535,N_20276);
nor U28787 (N_28787,N_23858,N_23788);
and U28788 (N_28788,N_24321,N_21953);
xor U28789 (N_28789,N_22064,N_20375);
and U28790 (N_28790,N_20777,N_23177);
nor U28791 (N_28791,N_23657,N_23058);
nand U28792 (N_28792,N_20661,N_20474);
xor U28793 (N_28793,N_23960,N_24472);
nor U28794 (N_28794,N_24820,N_22110);
nor U28795 (N_28795,N_22540,N_22572);
and U28796 (N_28796,N_22914,N_24550);
nand U28797 (N_28797,N_24437,N_22256);
or U28798 (N_28798,N_22513,N_20468);
nand U28799 (N_28799,N_22268,N_20614);
and U28800 (N_28800,N_22037,N_20168);
nor U28801 (N_28801,N_20244,N_20785);
and U28802 (N_28802,N_20193,N_21456);
xor U28803 (N_28803,N_23879,N_24475);
xnor U28804 (N_28804,N_23385,N_22979);
and U28805 (N_28805,N_20007,N_22521);
nor U28806 (N_28806,N_23060,N_21023);
or U28807 (N_28807,N_22434,N_21612);
nor U28808 (N_28808,N_23116,N_22726);
nor U28809 (N_28809,N_21812,N_24635);
and U28810 (N_28810,N_23821,N_22797);
and U28811 (N_28811,N_22341,N_20538);
or U28812 (N_28812,N_23402,N_22004);
xnor U28813 (N_28813,N_23941,N_20090);
xnor U28814 (N_28814,N_24013,N_20726);
and U28815 (N_28815,N_24725,N_24528);
nand U28816 (N_28816,N_24828,N_21273);
nand U28817 (N_28817,N_24091,N_22820);
nor U28818 (N_28818,N_22702,N_23294);
xnor U28819 (N_28819,N_23709,N_21576);
nand U28820 (N_28820,N_21352,N_23696);
nand U28821 (N_28821,N_23349,N_21887);
nand U28822 (N_28822,N_23398,N_24690);
or U28823 (N_28823,N_20287,N_21809);
or U28824 (N_28824,N_23874,N_24676);
xnor U28825 (N_28825,N_21272,N_21159);
nand U28826 (N_28826,N_21486,N_22521);
or U28827 (N_28827,N_24358,N_21181);
nor U28828 (N_28828,N_21412,N_21946);
xor U28829 (N_28829,N_23747,N_21025);
or U28830 (N_28830,N_21998,N_24387);
nor U28831 (N_28831,N_20894,N_23672);
and U28832 (N_28832,N_22895,N_23380);
and U28833 (N_28833,N_22869,N_23695);
nor U28834 (N_28834,N_23580,N_24137);
or U28835 (N_28835,N_22456,N_20061);
and U28836 (N_28836,N_24843,N_20510);
nor U28837 (N_28837,N_23884,N_24070);
nand U28838 (N_28838,N_24447,N_24119);
xor U28839 (N_28839,N_22447,N_21729);
or U28840 (N_28840,N_24651,N_23331);
nand U28841 (N_28841,N_20330,N_21945);
and U28842 (N_28842,N_23220,N_21725);
xnor U28843 (N_28843,N_23098,N_22404);
nor U28844 (N_28844,N_20289,N_22185);
xor U28845 (N_28845,N_21296,N_24528);
or U28846 (N_28846,N_22820,N_20036);
and U28847 (N_28847,N_23358,N_23515);
nor U28848 (N_28848,N_24178,N_24981);
and U28849 (N_28849,N_21642,N_22141);
or U28850 (N_28850,N_24565,N_20657);
and U28851 (N_28851,N_23380,N_20558);
and U28852 (N_28852,N_20364,N_24138);
or U28853 (N_28853,N_22754,N_23227);
and U28854 (N_28854,N_22840,N_20516);
and U28855 (N_28855,N_22179,N_21622);
nor U28856 (N_28856,N_21545,N_22334);
or U28857 (N_28857,N_23722,N_22669);
and U28858 (N_28858,N_20976,N_21108);
and U28859 (N_28859,N_22159,N_21141);
nand U28860 (N_28860,N_23060,N_22797);
xnor U28861 (N_28861,N_22409,N_24602);
nor U28862 (N_28862,N_20605,N_22357);
nand U28863 (N_28863,N_20228,N_22943);
nor U28864 (N_28864,N_20630,N_20480);
and U28865 (N_28865,N_24476,N_21370);
or U28866 (N_28866,N_24461,N_22481);
xnor U28867 (N_28867,N_22056,N_20014);
or U28868 (N_28868,N_21762,N_24673);
or U28869 (N_28869,N_24507,N_21969);
or U28870 (N_28870,N_23051,N_21586);
nor U28871 (N_28871,N_24410,N_24044);
nor U28872 (N_28872,N_21077,N_21740);
and U28873 (N_28873,N_23231,N_20680);
or U28874 (N_28874,N_24561,N_20502);
nor U28875 (N_28875,N_23094,N_24527);
xnor U28876 (N_28876,N_24350,N_24551);
and U28877 (N_28877,N_20317,N_22230);
or U28878 (N_28878,N_20339,N_22607);
or U28879 (N_28879,N_21416,N_20995);
and U28880 (N_28880,N_24869,N_21402);
or U28881 (N_28881,N_20034,N_24774);
xnor U28882 (N_28882,N_20154,N_22669);
and U28883 (N_28883,N_23639,N_24322);
nand U28884 (N_28884,N_23677,N_20289);
nand U28885 (N_28885,N_23236,N_23694);
nor U28886 (N_28886,N_22567,N_23966);
or U28887 (N_28887,N_23712,N_23913);
and U28888 (N_28888,N_21314,N_22931);
or U28889 (N_28889,N_20850,N_22494);
xor U28890 (N_28890,N_20733,N_23526);
xnor U28891 (N_28891,N_20766,N_24302);
or U28892 (N_28892,N_24823,N_21157);
and U28893 (N_28893,N_21711,N_23301);
nand U28894 (N_28894,N_21222,N_23229);
or U28895 (N_28895,N_22116,N_23873);
or U28896 (N_28896,N_20876,N_20105);
and U28897 (N_28897,N_24926,N_23042);
and U28898 (N_28898,N_22648,N_22670);
xnor U28899 (N_28899,N_20599,N_21552);
nand U28900 (N_28900,N_22040,N_24443);
and U28901 (N_28901,N_21818,N_20423);
and U28902 (N_28902,N_22533,N_23761);
xor U28903 (N_28903,N_22174,N_24644);
nor U28904 (N_28904,N_22206,N_23277);
xnor U28905 (N_28905,N_24379,N_20300);
and U28906 (N_28906,N_22759,N_21128);
and U28907 (N_28907,N_21399,N_23948);
nor U28908 (N_28908,N_21707,N_23906);
or U28909 (N_28909,N_20515,N_20432);
nand U28910 (N_28910,N_22171,N_20250);
or U28911 (N_28911,N_23351,N_24380);
and U28912 (N_28912,N_22124,N_20024);
or U28913 (N_28913,N_24804,N_22771);
nor U28914 (N_28914,N_20093,N_22467);
nor U28915 (N_28915,N_23111,N_21072);
xnor U28916 (N_28916,N_23377,N_21480);
nand U28917 (N_28917,N_21349,N_21220);
nand U28918 (N_28918,N_20909,N_24181);
xor U28919 (N_28919,N_23605,N_22093);
or U28920 (N_28920,N_24504,N_24229);
or U28921 (N_28921,N_24231,N_21848);
nand U28922 (N_28922,N_21232,N_20880);
and U28923 (N_28923,N_23196,N_22921);
or U28924 (N_28924,N_24686,N_23240);
and U28925 (N_28925,N_22630,N_20117);
nand U28926 (N_28926,N_20287,N_20989);
xnor U28927 (N_28927,N_21243,N_21532);
xor U28928 (N_28928,N_21855,N_22479);
and U28929 (N_28929,N_20071,N_22296);
and U28930 (N_28930,N_21716,N_23181);
and U28931 (N_28931,N_20376,N_24840);
and U28932 (N_28932,N_24865,N_22031);
nand U28933 (N_28933,N_21597,N_21194);
and U28934 (N_28934,N_20681,N_23513);
xor U28935 (N_28935,N_22223,N_21108);
nand U28936 (N_28936,N_22647,N_22872);
or U28937 (N_28937,N_20102,N_20465);
or U28938 (N_28938,N_20244,N_20653);
xor U28939 (N_28939,N_22372,N_20339);
nor U28940 (N_28940,N_21511,N_20214);
xor U28941 (N_28941,N_21029,N_23977);
or U28942 (N_28942,N_23702,N_23885);
xor U28943 (N_28943,N_22581,N_23666);
and U28944 (N_28944,N_20226,N_24298);
and U28945 (N_28945,N_22356,N_22851);
or U28946 (N_28946,N_22776,N_21910);
xor U28947 (N_28947,N_20190,N_20005);
and U28948 (N_28948,N_23191,N_23997);
nand U28949 (N_28949,N_24919,N_24896);
nand U28950 (N_28950,N_22951,N_20985);
xnor U28951 (N_28951,N_23140,N_21489);
nand U28952 (N_28952,N_21465,N_23375);
nand U28953 (N_28953,N_21320,N_23016);
nor U28954 (N_28954,N_21985,N_21460);
and U28955 (N_28955,N_24620,N_24701);
nor U28956 (N_28956,N_23102,N_24992);
or U28957 (N_28957,N_23548,N_20834);
xnor U28958 (N_28958,N_20950,N_20452);
nand U28959 (N_28959,N_21432,N_23409);
nand U28960 (N_28960,N_24219,N_24401);
nor U28961 (N_28961,N_22313,N_20906);
or U28962 (N_28962,N_23286,N_20651);
xor U28963 (N_28963,N_22429,N_23361);
xnor U28964 (N_28964,N_20981,N_21958);
nand U28965 (N_28965,N_21707,N_23411);
nor U28966 (N_28966,N_23366,N_22006);
nor U28967 (N_28967,N_21168,N_22066);
and U28968 (N_28968,N_20021,N_21004);
xor U28969 (N_28969,N_24089,N_24071);
nor U28970 (N_28970,N_22284,N_22470);
xor U28971 (N_28971,N_22848,N_24287);
and U28972 (N_28972,N_22697,N_22894);
xnor U28973 (N_28973,N_21411,N_24437);
xnor U28974 (N_28974,N_23157,N_24872);
nand U28975 (N_28975,N_23246,N_20937);
nand U28976 (N_28976,N_23664,N_23502);
and U28977 (N_28977,N_22285,N_24377);
and U28978 (N_28978,N_22203,N_20743);
and U28979 (N_28979,N_22808,N_20562);
xnor U28980 (N_28980,N_21553,N_22624);
nand U28981 (N_28981,N_21634,N_20208);
nor U28982 (N_28982,N_20698,N_23357);
nor U28983 (N_28983,N_23912,N_24484);
xnor U28984 (N_28984,N_23877,N_22660);
xor U28985 (N_28985,N_21030,N_22349);
nor U28986 (N_28986,N_21210,N_24597);
and U28987 (N_28987,N_22102,N_23514);
xnor U28988 (N_28988,N_20543,N_21178);
or U28989 (N_28989,N_24884,N_20330);
xor U28990 (N_28990,N_20275,N_24349);
nand U28991 (N_28991,N_20040,N_22360);
nand U28992 (N_28992,N_21090,N_22104);
xnor U28993 (N_28993,N_21890,N_20563);
nor U28994 (N_28994,N_24780,N_23190);
nand U28995 (N_28995,N_23495,N_23516);
or U28996 (N_28996,N_24093,N_24838);
nor U28997 (N_28997,N_20832,N_24897);
or U28998 (N_28998,N_23024,N_22655);
and U28999 (N_28999,N_23991,N_24694);
nor U29000 (N_29000,N_22079,N_23030);
xor U29001 (N_29001,N_23533,N_23886);
xor U29002 (N_29002,N_21325,N_23011);
xor U29003 (N_29003,N_23151,N_23646);
xnor U29004 (N_29004,N_22327,N_22008);
nand U29005 (N_29005,N_22169,N_22758);
nand U29006 (N_29006,N_23576,N_20191);
and U29007 (N_29007,N_21468,N_23932);
nor U29008 (N_29008,N_20648,N_22047);
nand U29009 (N_29009,N_22493,N_21705);
nand U29010 (N_29010,N_21686,N_24715);
nand U29011 (N_29011,N_24474,N_24452);
or U29012 (N_29012,N_22393,N_21222);
nand U29013 (N_29013,N_24257,N_23392);
nor U29014 (N_29014,N_23036,N_23124);
nand U29015 (N_29015,N_20051,N_21122);
nand U29016 (N_29016,N_24873,N_24727);
or U29017 (N_29017,N_20436,N_23945);
nand U29018 (N_29018,N_23111,N_22031);
xor U29019 (N_29019,N_24906,N_23848);
nand U29020 (N_29020,N_23306,N_24474);
xnor U29021 (N_29021,N_20512,N_20824);
or U29022 (N_29022,N_22901,N_22219);
nor U29023 (N_29023,N_20969,N_21674);
nor U29024 (N_29024,N_21518,N_20949);
nor U29025 (N_29025,N_20897,N_20692);
and U29026 (N_29026,N_22564,N_22651);
nor U29027 (N_29027,N_22741,N_24575);
nor U29028 (N_29028,N_22163,N_22970);
nand U29029 (N_29029,N_23194,N_22871);
nor U29030 (N_29030,N_21921,N_22606);
xor U29031 (N_29031,N_21022,N_21351);
and U29032 (N_29032,N_21414,N_21191);
and U29033 (N_29033,N_20553,N_22962);
xor U29034 (N_29034,N_24076,N_21012);
nand U29035 (N_29035,N_22067,N_24334);
or U29036 (N_29036,N_20034,N_24409);
nand U29037 (N_29037,N_20449,N_22266);
nor U29038 (N_29038,N_23591,N_24400);
and U29039 (N_29039,N_23107,N_20620);
and U29040 (N_29040,N_22905,N_24570);
nor U29041 (N_29041,N_22644,N_22261);
nand U29042 (N_29042,N_20026,N_20915);
xnor U29043 (N_29043,N_20554,N_22253);
xor U29044 (N_29044,N_23043,N_23105);
or U29045 (N_29045,N_24516,N_24894);
nand U29046 (N_29046,N_22984,N_22572);
or U29047 (N_29047,N_22740,N_20911);
nor U29048 (N_29048,N_22754,N_23215);
nand U29049 (N_29049,N_20180,N_21250);
nand U29050 (N_29050,N_24185,N_24255);
or U29051 (N_29051,N_20544,N_20666);
xor U29052 (N_29052,N_24081,N_24659);
or U29053 (N_29053,N_24694,N_22766);
and U29054 (N_29054,N_23755,N_24213);
nor U29055 (N_29055,N_24516,N_22314);
xor U29056 (N_29056,N_21819,N_20217);
or U29057 (N_29057,N_23918,N_24284);
nor U29058 (N_29058,N_24631,N_22923);
and U29059 (N_29059,N_21773,N_20356);
and U29060 (N_29060,N_23130,N_23947);
or U29061 (N_29061,N_24267,N_23484);
nor U29062 (N_29062,N_21082,N_21209);
and U29063 (N_29063,N_24778,N_21015);
or U29064 (N_29064,N_23636,N_20472);
and U29065 (N_29065,N_20418,N_24429);
nor U29066 (N_29066,N_24396,N_21445);
xnor U29067 (N_29067,N_22040,N_22521);
or U29068 (N_29068,N_23678,N_23340);
nand U29069 (N_29069,N_23177,N_20793);
xor U29070 (N_29070,N_20452,N_24445);
xor U29071 (N_29071,N_24486,N_24517);
and U29072 (N_29072,N_20884,N_21232);
xor U29073 (N_29073,N_22550,N_24310);
and U29074 (N_29074,N_22012,N_24787);
nor U29075 (N_29075,N_21405,N_22254);
or U29076 (N_29076,N_21212,N_21715);
xor U29077 (N_29077,N_24510,N_21372);
and U29078 (N_29078,N_22929,N_23748);
or U29079 (N_29079,N_23370,N_24744);
and U29080 (N_29080,N_21241,N_22259);
nand U29081 (N_29081,N_23884,N_21396);
and U29082 (N_29082,N_22729,N_24487);
nand U29083 (N_29083,N_24342,N_20324);
xor U29084 (N_29084,N_22322,N_24994);
xnor U29085 (N_29085,N_20513,N_24564);
and U29086 (N_29086,N_21710,N_24697);
or U29087 (N_29087,N_21471,N_24903);
or U29088 (N_29088,N_22767,N_21195);
or U29089 (N_29089,N_22438,N_20020);
or U29090 (N_29090,N_24722,N_22060);
or U29091 (N_29091,N_20134,N_21117);
xor U29092 (N_29092,N_22321,N_20297);
nor U29093 (N_29093,N_22817,N_22881);
nor U29094 (N_29094,N_23861,N_20531);
and U29095 (N_29095,N_21779,N_22552);
and U29096 (N_29096,N_24846,N_20784);
xor U29097 (N_29097,N_21947,N_24387);
xnor U29098 (N_29098,N_22075,N_23442);
or U29099 (N_29099,N_22320,N_23979);
or U29100 (N_29100,N_22404,N_22237);
xnor U29101 (N_29101,N_21399,N_21007);
nand U29102 (N_29102,N_24904,N_20227);
and U29103 (N_29103,N_22842,N_23595);
and U29104 (N_29104,N_20982,N_23646);
nand U29105 (N_29105,N_22255,N_21295);
xor U29106 (N_29106,N_24807,N_23997);
nand U29107 (N_29107,N_23524,N_21281);
or U29108 (N_29108,N_24490,N_21590);
nand U29109 (N_29109,N_20875,N_23449);
nor U29110 (N_29110,N_21685,N_22169);
and U29111 (N_29111,N_21329,N_23494);
and U29112 (N_29112,N_20236,N_22971);
nand U29113 (N_29113,N_23975,N_21864);
and U29114 (N_29114,N_23388,N_20525);
or U29115 (N_29115,N_21317,N_23590);
nand U29116 (N_29116,N_22268,N_22228);
and U29117 (N_29117,N_21066,N_22091);
or U29118 (N_29118,N_24826,N_22312);
or U29119 (N_29119,N_22615,N_22004);
xnor U29120 (N_29120,N_23371,N_20541);
and U29121 (N_29121,N_20447,N_24075);
nand U29122 (N_29122,N_21748,N_21606);
or U29123 (N_29123,N_21899,N_20163);
nand U29124 (N_29124,N_20623,N_22676);
or U29125 (N_29125,N_20774,N_20940);
nor U29126 (N_29126,N_21075,N_20963);
nand U29127 (N_29127,N_24021,N_21622);
or U29128 (N_29128,N_20440,N_22021);
or U29129 (N_29129,N_21925,N_21815);
nand U29130 (N_29130,N_22009,N_21804);
nor U29131 (N_29131,N_24260,N_22911);
xnor U29132 (N_29132,N_23125,N_20796);
or U29133 (N_29133,N_22288,N_21999);
or U29134 (N_29134,N_21836,N_20459);
or U29135 (N_29135,N_20023,N_20024);
or U29136 (N_29136,N_24841,N_24347);
nand U29137 (N_29137,N_23104,N_24922);
nor U29138 (N_29138,N_23060,N_21570);
or U29139 (N_29139,N_22938,N_21622);
and U29140 (N_29140,N_24953,N_20727);
and U29141 (N_29141,N_24637,N_21212);
nand U29142 (N_29142,N_20677,N_22661);
xnor U29143 (N_29143,N_23653,N_23436);
and U29144 (N_29144,N_20735,N_23845);
or U29145 (N_29145,N_21071,N_20477);
nand U29146 (N_29146,N_23705,N_23282);
and U29147 (N_29147,N_23045,N_20530);
nor U29148 (N_29148,N_24238,N_23331);
nor U29149 (N_29149,N_22776,N_23106);
or U29150 (N_29150,N_24013,N_20006);
and U29151 (N_29151,N_24705,N_20366);
nor U29152 (N_29152,N_23601,N_21494);
and U29153 (N_29153,N_23628,N_22254);
and U29154 (N_29154,N_24342,N_21148);
nand U29155 (N_29155,N_22363,N_22471);
nor U29156 (N_29156,N_22362,N_20345);
and U29157 (N_29157,N_22860,N_20889);
xor U29158 (N_29158,N_20775,N_20788);
nor U29159 (N_29159,N_21313,N_23115);
xor U29160 (N_29160,N_21973,N_20854);
nor U29161 (N_29161,N_22101,N_20102);
and U29162 (N_29162,N_21845,N_23695);
or U29163 (N_29163,N_23559,N_21392);
nor U29164 (N_29164,N_21509,N_24759);
nand U29165 (N_29165,N_23923,N_23635);
or U29166 (N_29166,N_20962,N_24408);
xor U29167 (N_29167,N_23254,N_23529);
nand U29168 (N_29168,N_20343,N_22226);
xor U29169 (N_29169,N_20028,N_24550);
xnor U29170 (N_29170,N_24170,N_22865);
xor U29171 (N_29171,N_22179,N_23069);
nor U29172 (N_29172,N_22241,N_23053);
and U29173 (N_29173,N_22121,N_23623);
and U29174 (N_29174,N_23443,N_23687);
or U29175 (N_29175,N_21122,N_20102);
xnor U29176 (N_29176,N_22424,N_22683);
xor U29177 (N_29177,N_20454,N_21375);
or U29178 (N_29178,N_24069,N_23063);
xnor U29179 (N_29179,N_24280,N_21191);
nand U29180 (N_29180,N_21432,N_23708);
and U29181 (N_29181,N_23920,N_24316);
nor U29182 (N_29182,N_20871,N_23750);
and U29183 (N_29183,N_20402,N_23426);
and U29184 (N_29184,N_22868,N_21530);
nor U29185 (N_29185,N_24173,N_23406);
xnor U29186 (N_29186,N_20313,N_24164);
nand U29187 (N_29187,N_22667,N_21895);
xor U29188 (N_29188,N_20151,N_20043);
xor U29189 (N_29189,N_24894,N_23271);
or U29190 (N_29190,N_23058,N_22826);
nor U29191 (N_29191,N_24838,N_20068);
nand U29192 (N_29192,N_24017,N_24269);
and U29193 (N_29193,N_20097,N_20350);
xor U29194 (N_29194,N_23899,N_21067);
nor U29195 (N_29195,N_20652,N_22950);
or U29196 (N_29196,N_24718,N_21100);
nand U29197 (N_29197,N_20818,N_22870);
or U29198 (N_29198,N_21181,N_21782);
nand U29199 (N_29199,N_23928,N_21067);
nand U29200 (N_29200,N_23783,N_20031);
and U29201 (N_29201,N_21598,N_20148);
or U29202 (N_29202,N_23159,N_24484);
or U29203 (N_29203,N_21984,N_23472);
and U29204 (N_29204,N_24886,N_24149);
nor U29205 (N_29205,N_22252,N_23119);
nor U29206 (N_29206,N_23435,N_23277);
nand U29207 (N_29207,N_21975,N_21769);
and U29208 (N_29208,N_22657,N_23454);
and U29209 (N_29209,N_21795,N_24341);
xor U29210 (N_29210,N_21191,N_20618);
or U29211 (N_29211,N_24898,N_24884);
nor U29212 (N_29212,N_24712,N_21151);
xor U29213 (N_29213,N_24252,N_20294);
nand U29214 (N_29214,N_22834,N_20456);
or U29215 (N_29215,N_23662,N_20865);
and U29216 (N_29216,N_24737,N_22903);
and U29217 (N_29217,N_20508,N_22136);
nor U29218 (N_29218,N_24910,N_22552);
nor U29219 (N_29219,N_24488,N_21725);
nand U29220 (N_29220,N_23426,N_20524);
or U29221 (N_29221,N_21468,N_21051);
or U29222 (N_29222,N_23634,N_23623);
nand U29223 (N_29223,N_21551,N_23523);
nand U29224 (N_29224,N_22202,N_24691);
or U29225 (N_29225,N_22030,N_24320);
or U29226 (N_29226,N_22871,N_21860);
nor U29227 (N_29227,N_21089,N_24896);
and U29228 (N_29228,N_23754,N_22475);
nand U29229 (N_29229,N_23270,N_22161);
nor U29230 (N_29230,N_24654,N_24440);
nand U29231 (N_29231,N_23819,N_21911);
xnor U29232 (N_29232,N_20196,N_21034);
or U29233 (N_29233,N_22747,N_23268);
nand U29234 (N_29234,N_21796,N_23658);
or U29235 (N_29235,N_23890,N_23256);
xor U29236 (N_29236,N_21863,N_24670);
or U29237 (N_29237,N_20304,N_24288);
nor U29238 (N_29238,N_21726,N_20428);
nand U29239 (N_29239,N_20673,N_22349);
nor U29240 (N_29240,N_21084,N_21283);
or U29241 (N_29241,N_23840,N_20455);
nand U29242 (N_29242,N_22637,N_22512);
nor U29243 (N_29243,N_22241,N_24177);
and U29244 (N_29244,N_24259,N_23889);
or U29245 (N_29245,N_23430,N_20734);
nor U29246 (N_29246,N_20535,N_24627);
or U29247 (N_29247,N_22730,N_23829);
xnor U29248 (N_29248,N_23676,N_21012);
nand U29249 (N_29249,N_20125,N_23383);
nor U29250 (N_29250,N_23167,N_22486);
nand U29251 (N_29251,N_23000,N_23445);
nor U29252 (N_29252,N_20742,N_21546);
or U29253 (N_29253,N_24491,N_21495);
xnor U29254 (N_29254,N_22337,N_21086);
or U29255 (N_29255,N_20599,N_23811);
and U29256 (N_29256,N_22945,N_24568);
xor U29257 (N_29257,N_21583,N_24106);
or U29258 (N_29258,N_24409,N_21241);
xor U29259 (N_29259,N_20735,N_21989);
or U29260 (N_29260,N_24456,N_22342);
nand U29261 (N_29261,N_22552,N_23765);
nor U29262 (N_29262,N_23601,N_20106);
and U29263 (N_29263,N_22162,N_20526);
nand U29264 (N_29264,N_24384,N_23466);
nand U29265 (N_29265,N_24157,N_20744);
nor U29266 (N_29266,N_23760,N_22813);
nor U29267 (N_29267,N_24812,N_21898);
or U29268 (N_29268,N_21758,N_21670);
xnor U29269 (N_29269,N_20432,N_24262);
nand U29270 (N_29270,N_24027,N_22415);
and U29271 (N_29271,N_23307,N_20800);
nor U29272 (N_29272,N_23148,N_24296);
nor U29273 (N_29273,N_21739,N_24551);
xnor U29274 (N_29274,N_21063,N_21591);
nand U29275 (N_29275,N_20591,N_22575);
nor U29276 (N_29276,N_20958,N_23180);
nand U29277 (N_29277,N_23911,N_22088);
or U29278 (N_29278,N_22944,N_21998);
xnor U29279 (N_29279,N_22065,N_20950);
xnor U29280 (N_29280,N_24919,N_24922);
and U29281 (N_29281,N_22944,N_21785);
and U29282 (N_29282,N_20846,N_24250);
nand U29283 (N_29283,N_23971,N_21089);
or U29284 (N_29284,N_23794,N_21071);
or U29285 (N_29285,N_24560,N_22788);
xnor U29286 (N_29286,N_20889,N_23391);
nand U29287 (N_29287,N_23151,N_20208);
nand U29288 (N_29288,N_23240,N_23633);
nor U29289 (N_29289,N_24930,N_21437);
nand U29290 (N_29290,N_20277,N_24515);
and U29291 (N_29291,N_21089,N_21014);
nor U29292 (N_29292,N_20118,N_21525);
or U29293 (N_29293,N_22938,N_22696);
or U29294 (N_29294,N_24191,N_24812);
or U29295 (N_29295,N_23863,N_23084);
nand U29296 (N_29296,N_24269,N_21844);
nand U29297 (N_29297,N_23831,N_20579);
and U29298 (N_29298,N_23788,N_21301);
nor U29299 (N_29299,N_23407,N_24026);
nor U29300 (N_29300,N_20046,N_20769);
or U29301 (N_29301,N_22413,N_21323);
nand U29302 (N_29302,N_20114,N_24902);
nand U29303 (N_29303,N_23676,N_23851);
xor U29304 (N_29304,N_22774,N_23497);
nand U29305 (N_29305,N_24887,N_22899);
or U29306 (N_29306,N_24626,N_24691);
and U29307 (N_29307,N_22750,N_22027);
xnor U29308 (N_29308,N_23323,N_23310);
nand U29309 (N_29309,N_21452,N_21538);
or U29310 (N_29310,N_23285,N_22023);
and U29311 (N_29311,N_22431,N_23141);
and U29312 (N_29312,N_22636,N_23577);
xnor U29313 (N_29313,N_23041,N_21991);
nand U29314 (N_29314,N_21330,N_24582);
or U29315 (N_29315,N_23774,N_23488);
or U29316 (N_29316,N_23958,N_20002);
and U29317 (N_29317,N_22421,N_24625);
nor U29318 (N_29318,N_24023,N_22044);
nor U29319 (N_29319,N_20004,N_20504);
or U29320 (N_29320,N_24105,N_22817);
or U29321 (N_29321,N_22128,N_23321);
nor U29322 (N_29322,N_21365,N_23130);
nand U29323 (N_29323,N_24428,N_20669);
or U29324 (N_29324,N_24388,N_21871);
or U29325 (N_29325,N_20245,N_24444);
and U29326 (N_29326,N_23612,N_22791);
or U29327 (N_29327,N_24878,N_20202);
nand U29328 (N_29328,N_23349,N_24328);
nand U29329 (N_29329,N_21745,N_21571);
xor U29330 (N_29330,N_21039,N_24232);
or U29331 (N_29331,N_23586,N_22761);
xor U29332 (N_29332,N_22174,N_20585);
and U29333 (N_29333,N_21901,N_21232);
nand U29334 (N_29334,N_20615,N_20304);
and U29335 (N_29335,N_20958,N_21045);
nor U29336 (N_29336,N_20455,N_21701);
and U29337 (N_29337,N_24915,N_22219);
nand U29338 (N_29338,N_21584,N_22637);
and U29339 (N_29339,N_23010,N_20571);
and U29340 (N_29340,N_23307,N_21620);
and U29341 (N_29341,N_22416,N_22858);
xnor U29342 (N_29342,N_21895,N_22602);
or U29343 (N_29343,N_24908,N_23662);
xor U29344 (N_29344,N_24393,N_21763);
nor U29345 (N_29345,N_22468,N_22484);
nand U29346 (N_29346,N_20604,N_24312);
nor U29347 (N_29347,N_21863,N_23949);
nand U29348 (N_29348,N_22064,N_23646);
nor U29349 (N_29349,N_20105,N_21126);
and U29350 (N_29350,N_22545,N_21606);
xnor U29351 (N_29351,N_22313,N_24851);
nand U29352 (N_29352,N_23708,N_21466);
nor U29353 (N_29353,N_23238,N_23617);
nand U29354 (N_29354,N_20907,N_22240);
xor U29355 (N_29355,N_21918,N_20905);
xor U29356 (N_29356,N_20039,N_20779);
nor U29357 (N_29357,N_21850,N_22448);
nor U29358 (N_29358,N_24068,N_20366);
and U29359 (N_29359,N_21007,N_22083);
and U29360 (N_29360,N_21606,N_24190);
or U29361 (N_29361,N_23268,N_20078);
nor U29362 (N_29362,N_24344,N_22575);
and U29363 (N_29363,N_23975,N_20062);
nand U29364 (N_29364,N_24562,N_22588);
and U29365 (N_29365,N_22276,N_20771);
nor U29366 (N_29366,N_21121,N_24003);
xor U29367 (N_29367,N_22491,N_20822);
and U29368 (N_29368,N_23575,N_21459);
or U29369 (N_29369,N_24171,N_24841);
nand U29370 (N_29370,N_23921,N_23282);
nand U29371 (N_29371,N_22327,N_22870);
nand U29372 (N_29372,N_22108,N_24252);
and U29373 (N_29373,N_20943,N_24715);
nor U29374 (N_29374,N_22209,N_22403);
xnor U29375 (N_29375,N_21044,N_23279);
and U29376 (N_29376,N_23645,N_20325);
xnor U29377 (N_29377,N_24094,N_20146);
nor U29378 (N_29378,N_22780,N_24507);
nand U29379 (N_29379,N_24313,N_21947);
nor U29380 (N_29380,N_23579,N_21558);
nand U29381 (N_29381,N_22308,N_21158);
nor U29382 (N_29382,N_20598,N_21827);
nand U29383 (N_29383,N_23527,N_23626);
or U29384 (N_29384,N_23208,N_22503);
nand U29385 (N_29385,N_23450,N_21279);
nand U29386 (N_29386,N_23728,N_23976);
nor U29387 (N_29387,N_23085,N_24724);
xnor U29388 (N_29388,N_24324,N_23228);
nand U29389 (N_29389,N_23742,N_20804);
nor U29390 (N_29390,N_21491,N_21781);
nor U29391 (N_29391,N_21722,N_23864);
or U29392 (N_29392,N_21897,N_21610);
nor U29393 (N_29393,N_23172,N_21761);
or U29394 (N_29394,N_21318,N_24648);
nand U29395 (N_29395,N_20864,N_23414);
nand U29396 (N_29396,N_23659,N_22529);
nand U29397 (N_29397,N_24224,N_21098);
or U29398 (N_29398,N_23077,N_22649);
nand U29399 (N_29399,N_24778,N_20261);
xnor U29400 (N_29400,N_23700,N_21939);
nand U29401 (N_29401,N_22790,N_20474);
or U29402 (N_29402,N_21503,N_22047);
xnor U29403 (N_29403,N_24670,N_23683);
nor U29404 (N_29404,N_20196,N_21813);
nor U29405 (N_29405,N_24424,N_20597);
nor U29406 (N_29406,N_23503,N_23643);
nor U29407 (N_29407,N_20460,N_21100);
nand U29408 (N_29408,N_22839,N_22259);
xor U29409 (N_29409,N_21592,N_21182);
or U29410 (N_29410,N_20247,N_21376);
nand U29411 (N_29411,N_22034,N_21636);
nand U29412 (N_29412,N_24910,N_24420);
xor U29413 (N_29413,N_22625,N_20520);
and U29414 (N_29414,N_21565,N_23792);
and U29415 (N_29415,N_23081,N_21306);
xor U29416 (N_29416,N_24244,N_23843);
or U29417 (N_29417,N_21157,N_24208);
and U29418 (N_29418,N_20220,N_21497);
nor U29419 (N_29419,N_20956,N_22455);
or U29420 (N_29420,N_20399,N_22407);
nand U29421 (N_29421,N_23900,N_24859);
nand U29422 (N_29422,N_21082,N_20228);
nand U29423 (N_29423,N_24869,N_24229);
and U29424 (N_29424,N_22263,N_20710);
or U29425 (N_29425,N_22710,N_21270);
or U29426 (N_29426,N_23545,N_22827);
or U29427 (N_29427,N_23501,N_22472);
or U29428 (N_29428,N_23277,N_24343);
xnor U29429 (N_29429,N_23959,N_24045);
nor U29430 (N_29430,N_21116,N_23007);
nor U29431 (N_29431,N_23176,N_20842);
nand U29432 (N_29432,N_24253,N_21274);
nor U29433 (N_29433,N_24289,N_24058);
and U29434 (N_29434,N_21211,N_23229);
xor U29435 (N_29435,N_21090,N_24698);
or U29436 (N_29436,N_23767,N_21128);
nor U29437 (N_29437,N_21981,N_20085);
or U29438 (N_29438,N_21926,N_23554);
xnor U29439 (N_29439,N_21200,N_20954);
xnor U29440 (N_29440,N_20185,N_20369);
xor U29441 (N_29441,N_20052,N_20345);
and U29442 (N_29442,N_21112,N_24128);
and U29443 (N_29443,N_20268,N_23789);
xor U29444 (N_29444,N_23616,N_20170);
nand U29445 (N_29445,N_21103,N_23670);
or U29446 (N_29446,N_23674,N_20155);
nor U29447 (N_29447,N_23991,N_22234);
and U29448 (N_29448,N_23963,N_23198);
or U29449 (N_29449,N_20159,N_22835);
and U29450 (N_29450,N_20424,N_20281);
nor U29451 (N_29451,N_24027,N_24327);
xnor U29452 (N_29452,N_24842,N_21577);
nor U29453 (N_29453,N_21549,N_22795);
xnor U29454 (N_29454,N_22332,N_24504);
or U29455 (N_29455,N_21316,N_21413);
and U29456 (N_29456,N_22399,N_23262);
and U29457 (N_29457,N_24820,N_20478);
xor U29458 (N_29458,N_23119,N_23982);
or U29459 (N_29459,N_24763,N_23436);
xor U29460 (N_29460,N_24566,N_22432);
or U29461 (N_29461,N_21297,N_21570);
nand U29462 (N_29462,N_20936,N_24925);
and U29463 (N_29463,N_23292,N_22617);
nor U29464 (N_29464,N_21318,N_22164);
nand U29465 (N_29465,N_24719,N_23751);
xnor U29466 (N_29466,N_24672,N_24162);
and U29467 (N_29467,N_21693,N_20392);
xor U29468 (N_29468,N_20314,N_20838);
nor U29469 (N_29469,N_23085,N_22720);
or U29470 (N_29470,N_23989,N_24055);
nor U29471 (N_29471,N_21821,N_21409);
nand U29472 (N_29472,N_23348,N_21031);
nor U29473 (N_29473,N_24812,N_22354);
xnor U29474 (N_29474,N_23683,N_21341);
or U29475 (N_29475,N_23437,N_24198);
xor U29476 (N_29476,N_23167,N_24063);
or U29477 (N_29477,N_20546,N_22053);
xnor U29478 (N_29478,N_24423,N_23771);
xnor U29479 (N_29479,N_22427,N_21768);
and U29480 (N_29480,N_21123,N_23116);
or U29481 (N_29481,N_24243,N_21720);
and U29482 (N_29482,N_24323,N_21792);
nand U29483 (N_29483,N_24374,N_22327);
nand U29484 (N_29484,N_22764,N_20798);
or U29485 (N_29485,N_24374,N_21824);
and U29486 (N_29486,N_21093,N_24389);
or U29487 (N_29487,N_24034,N_22908);
nand U29488 (N_29488,N_22376,N_22196);
xor U29489 (N_29489,N_24089,N_20968);
and U29490 (N_29490,N_23055,N_24357);
xor U29491 (N_29491,N_22364,N_22007);
xnor U29492 (N_29492,N_24668,N_22035);
or U29493 (N_29493,N_21908,N_20379);
or U29494 (N_29494,N_23890,N_21345);
nor U29495 (N_29495,N_22647,N_22875);
xnor U29496 (N_29496,N_23494,N_20666);
nand U29497 (N_29497,N_22674,N_23678);
nor U29498 (N_29498,N_21764,N_21410);
and U29499 (N_29499,N_20135,N_20147);
and U29500 (N_29500,N_24577,N_21886);
or U29501 (N_29501,N_23521,N_23999);
nor U29502 (N_29502,N_22324,N_20594);
nor U29503 (N_29503,N_23866,N_24564);
nor U29504 (N_29504,N_24550,N_22686);
xnor U29505 (N_29505,N_20500,N_21931);
nor U29506 (N_29506,N_24230,N_22506);
xnor U29507 (N_29507,N_24326,N_20281);
xor U29508 (N_29508,N_21860,N_21411);
xor U29509 (N_29509,N_24151,N_20850);
and U29510 (N_29510,N_20617,N_21129);
and U29511 (N_29511,N_22763,N_21612);
nor U29512 (N_29512,N_22973,N_21103);
nand U29513 (N_29513,N_20205,N_24771);
and U29514 (N_29514,N_24300,N_23356);
nand U29515 (N_29515,N_20483,N_20198);
nor U29516 (N_29516,N_21479,N_24060);
nand U29517 (N_29517,N_24385,N_22567);
xnor U29518 (N_29518,N_24895,N_20923);
xor U29519 (N_29519,N_20817,N_24177);
and U29520 (N_29520,N_22539,N_20120);
and U29521 (N_29521,N_23961,N_22529);
nand U29522 (N_29522,N_24926,N_22427);
xnor U29523 (N_29523,N_20284,N_22484);
nand U29524 (N_29524,N_22155,N_24236);
xor U29525 (N_29525,N_23582,N_22909);
xnor U29526 (N_29526,N_20886,N_20186);
and U29527 (N_29527,N_23537,N_21155);
nand U29528 (N_29528,N_20134,N_21784);
xor U29529 (N_29529,N_21123,N_21697);
xnor U29530 (N_29530,N_22401,N_22002);
and U29531 (N_29531,N_23613,N_24782);
xnor U29532 (N_29532,N_21247,N_23674);
nand U29533 (N_29533,N_22742,N_20149);
nor U29534 (N_29534,N_20742,N_24449);
nand U29535 (N_29535,N_22307,N_21765);
nor U29536 (N_29536,N_20390,N_22161);
nand U29537 (N_29537,N_20302,N_22231);
or U29538 (N_29538,N_24393,N_23614);
nor U29539 (N_29539,N_22793,N_22765);
xnor U29540 (N_29540,N_23402,N_24071);
nor U29541 (N_29541,N_20551,N_22912);
nand U29542 (N_29542,N_23339,N_23947);
xor U29543 (N_29543,N_24662,N_24159);
or U29544 (N_29544,N_21511,N_24615);
or U29545 (N_29545,N_22683,N_23876);
and U29546 (N_29546,N_23939,N_22137);
xnor U29547 (N_29547,N_20071,N_23818);
nand U29548 (N_29548,N_23195,N_20580);
and U29549 (N_29549,N_24192,N_21491);
nand U29550 (N_29550,N_20094,N_24928);
or U29551 (N_29551,N_23647,N_22568);
nand U29552 (N_29552,N_23127,N_22337);
nor U29553 (N_29553,N_23515,N_20666);
nand U29554 (N_29554,N_24202,N_20266);
nand U29555 (N_29555,N_22668,N_22933);
xor U29556 (N_29556,N_24066,N_21510);
nor U29557 (N_29557,N_20913,N_22960);
nand U29558 (N_29558,N_24997,N_24950);
xnor U29559 (N_29559,N_22101,N_20361);
nand U29560 (N_29560,N_23547,N_21861);
or U29561 (N_29561,N_21202,N_23876);
nand U29562 (N_29562,N_24261,N_23563);
or U29563 (N_29563,N_22293,N_20359);
nand U29564 (N_29564,N_20065,N_23800);
nor U29565 (N_29565,N_20142,N_24892);
and U29566 (N_29566,N_24447,N_23223);
nor U29567 (N_29567,N_23323,N_23062);
nor U29568 (N_29568,N_23083,N_20147);
or U29569 (N_29569,N_20176,N_20579);
or U29570 (N_29570,N_23768,N_22380);
and U29571 (N_29571,N_22509,N_24205);
or U29572 (N_29572,N_21214,N_20670);
nand U29573 (N_29573,N_21675,N_23973);
xnor U29574 (N_29574,N_23410,N_22683);
or U29575 (N_29575,N_22254,N_21001);
xor U29576 (N_29576,N_20509,N_23997);
nor U29577 (N_29577,N_22161,N_24704);
and U29578 (N_29578,N_24675,N_22095);
xor U29579 (N_29579,N_24291,N_21168);
xnor U29580 (N_29580,N_22705,N_23098);
nor U29581 (N_29581,N_21283,N_20276);
or U29582 (N_29582,N_21933,N_20715);
nor U29583 (N_29583,N_21973,N_22315);
nand U29584 (N_29584,N_21109,N_24112);
xor U29585 (N_29585,N_23833,N_23815);
xor U29586 (N_29586,N_23134,N_22830);
nor U29587 (N_29587,N_20050,N_20335);
nand U29588 (N_29588,N_22826,N_20152);
and U29589 (N_29589,N_24369,N_20422);
nor U29590 (N_29590,N_23126,N_21685);
or U29591 (N_29591,N_24369,N_20221);
and U29592 (N_29592,N_22310,N_22688);
nor U29593 (N_29593,N_20099,N_23797);
and U29594 (N_29594,N_21736,N_22161);
or U29595 (N_29595,N_22102,N_21505);
and U29596 (N_29596,N_21120,N_20582);
and U29597 (N_29597,N_21299,N_21921);
nor U29598 (N_29598,N_23012,N_21608);
and U29599 (N_29599,N_21671,N_20180);
nor U29600 (N_29600,N_23250,N_22751);
nand U29601 (N_29601,N_20681,N_20001);
and U29602 (N_29602,N_20373,N_21849);
and U29603 (N_29603,N_23506,N_20248);
xor U29604 (N_29604,N_20922,N_20726);
or U29605 (N_29605,N_22308,N_24699);
nor U29606 (N_29606,N_21728,N_20290);
xor U29607 (N_29607,N_24476,N_23466);
nor U29608 (N_29608,N_24933,N_20287);
or U29609 (N_29609,N_22766,N_24510);
nor U29610 (N_29610,N_23793,N_20651);
xnor U29611 (N_29611,N_23299,N_21660);
or U29612 (N_29612,N_21605,N_24975);
nand U29613 (N_29613,N_22911,N_21087);
nand U29614 (N_29614,N_23107,N_24473);
or U29615 (N_29615,N_23010,N_20566);
nor U29616 (N_29616,N_21827,N_22760);
and U29617 (N_29617,N_21370,N_23335);
xnor U29618 (N_29618,N_22652,N_21414);
or U29619 (N_29619,N_23653,N_22429);
and U29620 (N_29620,N_20037,N_23630);
nor U29621 (N_29621,N_22848,N_21244);
nand U29622 (N_29622,N_21115,N_21314);
nand U29623 (N_29623,N_21847,N_21617);
xnor U29624 (N_29624,N_21204,N_23718);
xnor U29625 (N_29625,N_24743,N_23062);
nor U29626 (N_29626,N_21281,N_20108);
or U29627 (N_29627,N_23577,N_22093);
or U29628 (N_29628,N_24126,N_21256);
nand U29629 (N_29629,N_20250,N_22989);
and U29630 (N_29630,N_20899,N_23260);
nor U29631 (N_29631,N_21448,N_20455);
and U29632 (N_29632,N_21848,N_22894);
nor U29633 (N_29633,N_22095,N_24586);
or U29634 (N_29634,N_23949,N_20872);
nor U29635 (N_29635,N_21521,N_24987);
xor U29636 (N_29636,N_20925,N_21744);
nor U29637 (N_29637,N_22231,N_23059);
nor U29638 (N_29638,N_21710,N_21916);
xnor U29639 (N_29639,N_23625,N_21155);
nor U29640 (N_29640,N_22425,N_23237);
and U29641 (N_29641,N_20042,N_20808);
or U29642 (N_29642,N_20266,N_24628);
and U29643 (N_29643,N_24492,N_20808);
nor U29644 (N_29644,N_21742,N_24005);
nor U29645 (N_29645,N_21928,N_22315);
and U29646 (N_29646,N_20378,N_20165);
nand U29647 (N_29647,N_24759,N_22733);
nor U29648 (N_29648,N_23916,N_23561);
nand U29649 (N_29649,N_22869,N_20805);
or U29650 (N_29650,N_21589,N_20873);
nor U29651 (N_29651,N_24228,N_22044);
xnor U29652 (N_29652,N_23392,N_20084);
and U29653 (N_29653,N_24907,N_23099);
or U29654 (N_29654,N_21513,N_20824);
nor U29655 (N_29655,N_23837,N_20024);
or U29656 (N_29656,N_24717,N_24496);
or U29657 (N_29657,N_23634,N_24634);
nor U29658 (N_29658,N_20746,N_22930);
xnor U29659 (N_29659,N_21012,N_24470);
nor U29660 (N_29660,N_20164,N_22546);
and U29661 (N_29661,N_23320,N_20167);
and U29662 (N_29662,N_20376,N_21718);
or U29663 (N_29663,N_21841,N_22573);
xor U29664 (N_29664,N_22765,N_23833);
or U29665 (N_29665,N_21806,N_21673);
xor U29666 (N_29666,N_20298,N_20242);
xnor U29667 (N_29667,N_21652,N_20168);
or U29668 (N_29668,N_22842,N_24188);
xnor U29669 (N_29669,N_22773,N_23276);
or U29670 (N_29670,N_20912,N_20954);
nand U29671 (N_29671,N_20774,N_24755);
nand U29672 (N_29672,N_21869,N_24464);
or U29673 (N_29673,N_24237,N_22844);
and U29674 (N_29674,N_20897,N_23260);
or U29675 (N_29675,N_22380,N_23134);
and U29676 (N_29676,N_21891,N_24852);
xnor U29677 (N_29677,N_24937,N_23048);
and U29678 (N_29678,N_20426,N_24368);
and U29679 (N_29679,N_24096,N_22690);
xnor U29680 (N_29680,N_21716,N_24864);
and U29681 (N_29681,N_20447,N_22886);
nand U29682 (N_29682,N_24835,N_22649);
or U29683 (N_29683,N_22037,N_23212);
nand U29684 (N_29684,N_24287,N_20868);
or U29685 (N_29685,N_20654,N_24782);
nand U29686 (N_29686,N_24201,N_21630);
nor U29687 (N_29687,N_22433,N_23945);
and U29688 (N_29688,N_21419,N_22416);
nor U29689 (N_29689,N_20241,N_24626);
xor U29690 (N_29690,N_23449,N_21826);
nand U29691 (N_29691,N_23786,N_20031);
and U29692 (N_29692,N_21191,N_20387);
or U29693 (N_29693,N_24481,N_23322);
and U29694 (N_29694,N_22344,N_23445);
xnor U29695 (N_29695,N_20912,N_20608);
or U29696 (N_29696,N_23193,N_22248);
or U29697 (N_29697,N_21452,N_22198);
xnor U29698 (N_29698,N_23344,N_21835);
xnor U29699 (N_29699,N_23360,N_23682);
xnor U29700 (N_29700,N_24474,N_22623);
nand U29701 (N_29701,N_21272,N_21081);
and U29702 (N_29702,N_21470,N_22040);
nor U29703 (N_29703,N_23772,N_23697);
nor U29704 (N_29704,N_24158,N_24203);
nand U29705 (N_29705,N_20262,N_23337);
or U29706 (N_29706,N_22105,N_23491);
nand U29707 (N_29707,N_22511,N_21980);
xor U29708 (N_29708,N_20874,N_21393);
and U29709 (N_29709,N_21680,N_20041);
xor U29710 (N_29710,N_24971,N_23027);
and U29711 (N_29711,N_21856,N_24711);
and U29712 (N_29712,N_22303,N_24006);
nor U29713 (N_29713,N_20008,N_20151);
or U29714 (N_29714,N_20695,N_23356);
nand U29715 (N_29715,N_23533,N_20757);
or U29716 (N_29716,N_20317,N_21586);
and U29717 (N_29717,N_21052,N_20598);
and U29718 (N_29718,N_20330,N_22026);
nand U29719 (N_29719,N_20167,N_21989);
xnor U29720 (N_29720,N_23954,N_22250);
or U29721 (N_29721,N_24180,N_20735);
xor U29722 (N_29722,N_21457,N_21122);
xor U29723 (N_29723,N_23233,N_20880);
nand U29724 (N_29724,N_23050,N_23121);
nand U29725 (N_29725,N_20349,N_20222);
or U29726 (N_29726,N_22269,N_23903);
nand U29727 (N_29727,N_21692,N_22566);
nand U29728 (N_29728,N_23984,N_24519);
nand U29729 (N_29729,N_22283,N_20891);
nand U29730 (N_29730,N_21117,N_23869);
xnor U29731 (N_29731,N_20337,N_22301);
nor U29732 (N_29732,N_24557,N_20736);
or U29733 (N_29733,N_22037,N_24609);
nand U29734 (N_29734,N_20460,N_24829);
nor U29735 (N_29735,N_24395,N_21926);
or U29736 (N_29736,N_24903,N_23848);
xnor U29737 (N_29737,N_24042,N_24551);
xor U29738 (N_29738,N_22225,N_24901);
and U29739 (N_29739,N_23797,N_22764);
nand U29740 (N_29740,N_21886,N_23174);
or U29741 (N_29741,N_20508,N_21032);
xor U29742 (N_29742,N_21138,N_22793);
nand U29743 (N_29743,N_24625,N_21615);
nor U29744 (N_29744,N_23127,N_22018);
xor U29745 (N_29745,N_24694,N_22404);
and U29746 (N_29746,N_23524,N_24313);
and U29747 (N_29747,N_23505,N_22055);
or U29748 (N_29748,N_21556,N_24505);
xor U29749 (N_29749,N_21325,N_23391);
nor U29750 (N_29750,N_21081,N_21877);
nand U29751 (N_29751,N_24834,N_24781);
or U29752 (N_29752,N_24784,N_24343);
and U29753 (N_29753,N_22844,N_20024);
or U29754 (N_29754,N_21817,N_22424);
xor U29755 (N_29755,N_20443,N_24104);
nand U29756 (N_29756,N_23508,N_21647);
and U29757 (N_29757,N_20180,N_24457);
xnor U29758 (N_29758,N_21132,N_24678);
and U29759 (N_29759,N_21813,N_22032);
nand U29760 (N_29760,N_21196,N_22318);
nand U29761 (N_29761,N_22811,N_22843);
and U29762 (N_29762,N_22233,N_22273);
nor U29763 (N_29763,N_21014,N_21077);
or U29764 (N_29764,N_20686,N_23881);
or U29765 (N_29765,N_20169,N_24546);
xor U29766 (N_29766,N_20014,N_21163);
or U29767 (N_29767,N_21578,N_21105);
xnor U29768 (N_29768,N_24058,N_21382);
or U29769 (N_29769,N_22470,N_22544);
or U29770 (N_29770,N_22048,N_24181);
xnor U29771 (N_29771,N_22869,N_24134);
and U29772 (N_29772,N_20403,N_23022);
and U29773 (N_29773,N_20405,N_21783);
nor U29774 (N_29774,N_20613,N_24280);
and U29775 (N_29775,N_22165,N_21999);
nor U29776 (N_29776,N_23651,N_20834);
and U29777 (N_29777,N_20243,N_23532);
xor U29778 (N_29778,N_22166,N_21958);
nor U29779 (N_29779,N_21272,N_21827);
and U29780 (N_29780,N_24254,N_21318);
nor U29781 (N_29781,N_22322,N_20771);
xnor U29782 (N_29782,N_23818,N_24794);
nand U29783 (N_29783,N_20938,N_21755);
xor U29784 (N_29784,N_23347,N_22320);
and U29785 (N_29785,N_21679,N_24006);
and U29786 (N_29786,N_20544,N_22681);
and U29787 (N_29787,N_20499,N_20481);
and U29788 (N_29788,N_21356,N_20431);
or U29789 (N_29789,N_24591,N_21805);
xor U29790 (N_29790,N_21055,N_20743);
nor U29791 (N_29791,N_22846,N_20509);
nor U29792 (N_29792,N_20116,N_22964);
xnor U29793 (N_29793,N_22690,N_23178);
or U29794 (N_29794,N_24551,N_24916);
or U29795 (N_29795,N_22013,N_20377);
xor U29796 (N_29796,N_20400,N_21756);
xor U29797 (N_29797,N_24092,N_23848);
xor U29798 (N_29798,N_24835,N_22510);
nor U29799 (N_29799,N_24496,N_23879);
or U29800 (N_29800,N_23479,N_23922);
xnor U29801 (N_29801,N_24663,N_21519);
or U29802 (N_29802,N_20952,N_23832);
or U29803 (N_29803,N_23111,N_23196);
xnor U29804 (N_29804,N_22124,N_21752);
xor U29805 (N_29805,N_24196,N_20353);
and U29806 (N_29806,N_23945,N_23507);
nand U29807 (N_29807,N_24715,N_20979);
nand U29808 (N_29808,N_23289,N_23770);
nor U29809 (N_29809,N_20292,N_21539);
nand U29810 (N_29810,N_23980,N_21599);
nor U29811 (N_29811,N_20241,N_21950);
xnor U29812 (N_29812,N_23916,N_22146);
nand U29813 (N_29813,N_23714,N_24086);
nand U29814 (N_29814,N_22177,N_22212);
or U29815 (N_29815,N_20727,N_22816);
or U29816 (N_29816,N_20672,N_24371);
nor U29817 (N_29817,N_22338,N_24574);
or U29818 (N_29818,N_22718,N_21183);
and U29819 (N_29819,N_22787,N_23519);
or U29820 (N_29820,N_21539,N_23636);
xor U29821 (N_29821,N_21344,N_21295);
nor U29822 (N_29822,N_20917,N_21397);
and U29823 (N_29823,N_21115,N_22663);
xor U29824 (N_29824,N_21420,N_24022);
or U29825 (N_29825,N_22558,N_23031);
nand U29826 (N_29826,N_21222,N_21766);
nand U29827 (N_29827,N_22004,N_20077);
xor U29828 (N_29828,N_23413,N_24660);
nor U29829 (N_29829,N_21362,N_22499);
xor U29830 (N_29830,N_22823,N_24576);
or U29831 (N_29831,N_23991,N_20083);
or U29832 (N_29832,N_23651,N_24257);
or U29833 (N_29833,N_21042,N_22221);
nand U29834 (N_29834,N_21178,N_20871);
or U29835 (N_29835,N_20539,N_21573);
and U29836 (N_29836,N_24052,N_20796);
and U29837 (N_29837,N_20315,N_21145);
nor U29838 (N_29838,N_20482,N_20571);
or U29839 (N_29839,N_22457,N_23646);
or U29840 (N_29840,N_22342,N_24941);
and U29841 (N_29841,N_22620,N_22880);
nor U29842 (N_29842,N_21538,N_24672);
xor U29843 (N_29843,N_21773,N_24161);
nand U29844 (N_29844,N_22186,N_22300);
nand U29845 (N_29845,N_23116,N_24443);
or U29846 (N_29846,N_20962,N_23166);
xor U29847 (N_29847,N_20469,N_21096);
xor U29848 (N_29848,N_23128,N_24681);
xnor U29849 (N_29849,N_22044,N_22340);
and U29850 (N_29850,N_22342,N_20239);
and U29851 (N_29851,N_24770,N_21679);
xnor U29852 (N_29852,N_22160,N_22883);
xor U29853 (N_29853,N_20415,N_24347);
or U29854 (N_29854,N_23499,N_21323);
and U29855 (N_29855,N_24838,N_24493);
and U29856 (N_29856,N_24619,N_24496);
xor U29857 (N_29857,N_23682,N_22408);
and U29858 (N_29858,N_20332,N_20816);
or U29859 (N_29859,N_24946,N_24843);
or U29860 (N_29860,N_20727,N_23394);
nor U29861 (N_29861,N_23559,N_22765);
or U29862 (N_29862,N_21061,N_22444);
and U29863 (N_29863,N_21011,N_20846);
and U29864 (N_29864,N_20731,N_22431);
nor U29865 (N_29865,N_22222,N_21723);
nand U29866 (N_29866,N_23180,N_21519);
nand U29867 (N_29867,N_23066,N_24610);
xnor U29868 (N_29868,N_22919,N_22799);
or U29869 (N_29869,N_22510,N_21890);
or U29870 (N_29870,N_22787,N_20104);
and U29871 (N_29871,N_23330,N_24987);
and U29872 (N_29872,N_22476,N_20772);
nor U29873 (N_29873,N_22328,N_24251);
nor U29874 (N_29874,N_23744,N_23779);
and U29875 (N_29875,N_22789,N_24537);
and U29876 (N_29876,N_24279,N_22178);
xor U29877 (N_29877,N_23273,N_24828);
and U29878 (N_29878,N_23172,N_23051);
xnor U29879 (N_29879,N_20813,N_24450);
nor U29880 (N_29880,N_23201,N_20701);
or U29881 (N_29881,N_23610,N_24864);
xor U29882 (N_29882,N_22144,N_21841);
or U29883 (N_29883,N_22423,N_22004);
or U29884 (N_29884,N_22883,N_24030);
xor U29885 (N_29885,N_22699,N_22963);
xor U29886 (N_29886,N_22485,N_23675);
and U29887 (N_29887,N_24858,N_22488);
or U29888 (N_29888,N_20908,N_24425);
and U29889 (N_29889,N_24632,N_23916);
nand U29890 (N_29890,N_24592,N_21857);
nor U29891 (N_29891,N_23176,N_20197);
and U29892 (N_29892,N_20546,N_22135);
xnor U29893 (N_29893,N_22363,N_21317);
xnor U29894 (N_29894,N_22126,N_24336);
or U29895 (N_29895,N_23156,N_22319);
nand U29896 (N_29896,N_22125,N_23830);
nand U29897 (N_29897,N_21066,N_20764);
nor U29898 (N_29898,N_24564,N_21697);
xor U29899 (N_29899,N_20891,N_23785);
and U29900 (N_29900,N_22873,N_22316);
nand U29901 (N_29901,N_24447,N_20957);
nor U29902 (N_29902,N_24663,N_21072);
nor U29903 (N_29903,N_24446,N_21092);
and U29904 (N_29904,N_20561,N_22945);
xor U29905 (N_29905,N_24052,N_22119);
xnor U29906 (N_29906,N_22230,N_21477);
xnor U29907 (N_29907,N_22949,N_24807);
xnor U29908 (N_29908,N_20460,N_22308);
nand U29909 (N_29909,N_24257,N_22049);
nand U29910 (N_29910,N_23399,N_23838);
nand U29911 (N_29911,N_23208,N_23049);
nor U29912 (N_29912,N_22271,N_20216);
and U29913 (N_29913,N_22603,N_24172);
xnor U29914 (N_29914,N_22575,N_24599);
xnor U29915 (N_29915,N_20205,N_22275);
nor U29916 (N_29916,N_23220,N_22962);
nand U29917 (N_29917,N_23214,N_24867);
nand U29918 (N_29918,N_23622,N_20718);
nor U29919 (N_29919,N_23339,N_22074);
or U29920 (N_29920,N_22577,N_21099);
nand U29921 (N_29921,N_20101,N_22257);
xor U29922 (N_29922,N_20760,N_22122);
nor U29923 (N_29923,N_23145,N_22156);
nor U29924 (N_29924,N_22912,N_20848);
nand U29925 (N_29925,N_22352,N_21312);
nor U29926 (N_29926,N_20526,N_21507);
or U29927 (N_29927,N_23819,N_24640);
nor U29928 (N_29928,N_21450,N_21512);
xnor U29929 (N_29929,N_22699,N_22424);
or U29930 (N_29930,N_20380,N_24549);
xnor U29931 (N_29931,N_21981,N_20193);
or U29932 (N_29932,N_23485,N_24028);
and U29933 (N_29933,N_24405,N_23278);
or U29934 (N_29934,N_23948,N_21386);
nor U29935 (N_29935,N_21378,N_24924);
and U29936 (N_29936,N_20681,N_21386);
nor U29937 (N_29937,N_21593,N_20766);
nand U29938 (N_29938,N_21862,N_21034);
and U29939 (N_29939,N_24304,N_24795);
xor U29940 (N_29940,N_20868,N_23066);
xor U29941 (N_29941,N_24302,N_24776);
xor U29942 (N_29942,N_24015,N_22697);
nor U29943 (N_29943,N_22947,N_23169);
or U29944 (N_29944,N_23657,N_22133);
and U29945 (N_29945,N_24971,N_23338);
or U29946 (N_29946,N_23560,N_20731);
xnor U29947 (N_29947,N_21709,N_23485);
and U29948 (N_29948,N_21639,N_23642);
xor U29949 (N_29949,N_22918,N_21459);
or U29950 (N_29950,N_24511,N_20791);
nand U29951 (N_29951,N_21031,N_21300);
nor U29952 (N_29952,N_24807,N_23531);
nand U29953 (N_29953,N_21504,N_20537);
xor U29954 (N_29954,N_24490,N_24868);
nand U29955 (N_29955,N_20558,N_20042);
xnor U29956 (N_29956,N_21002,N_20617);
nor U29957 (N_29957,N_23542,N_20589);
and U29958 (N_29958,N_23889,N_23510);
nor U29959 (N_29959,N_22766,N_20340);
nor U29960 (N_29960,N_20184,N_24457);
nor U29961 (N_29961,N_22195,N_23306);
and U29962 (N_29962,N_20965,N_23797);
or U29963 (N_29963,N_24835,N_23850);
nand U29964 (N_29964,N_22642,N_23567);
nand U29965 (N_29965,N_20961,N_20745);
nand U29966 (N_29966,N_24212,N_24337);
or U29967 (N_29967,N_21834,N_20936);
xor U29968 (N_29968,N_21693,N_22261);
nand U29969 (N_29969,N_23290,N_24483);
xnor U29970 (N_29970,N_20618,N_24362);
nand U29971 (N_29971,N_20377,N_22856);
or U29972 (N_29972,N_24559,N_21596);
and U29973 (N_29973,N_23802,N_24657);
and U29974 (N_29974,N_20535,N_20748);
and U29975 (N_29975,N_22109,N_23306);
and U29976 (N_29976,N_21443,N_22231);
and U29977 (N_29977,N_21554,N_23215);
xnor U29978 (N_29978,N_21843,N_24937);
or U29979 (N_29979,N_20865,N_23459);
xor U29980 (N_29980,N_21548,N_24529);
nor U29981 (N_29981,N_20503,N_22334);
nand U29982 (N_29982,N_24115,N_22335);
or U29983 (N_29983,N_20367,N_21152);
nor U29984 (N_29984,N_21129,N_22691);
nand U29985 (N_29985,N_22937,N_22620);
nor U29986 (N_29986,N_24900,N_20411);
nand U29987 (N_29987,N_24121,N_20075);
and U29988 (N_29988,N_22721,N_22531);
xor U29989 (N_29989,N_22548,N_23319);
nor U29990 (N_29990,N_24168,N_23952);
nor U29991 (N_29991,N_23132,N_20996);
nor U29992 (N_29992,N_21916,N_21802);
or U29993 (N_29993,N_24735,N_20131);
or U29994 (N_29994,N_23821,N_20321);
nand U29995 (N_29995,N_20031,N_23393);
nor U29996 (N_29996,N_23137,N_21293);
nand U29997 (N_29997,N_21606,N_24090);
and U29998 (N_29998,N_21060,N_23953);
and U29999 (N_29999,N_23381,N_24627);
nand UO_0 (O_0,N_27453,N_29942);
nand UO_1 (O_1,N_29642,N_27636);
or UO_2 (O_2,N_26139,N_27186);
or UO_3 (O_3,N_25676,N_26451);
nand UO_4 (O_4,N_26244,N_25426);
and UO_5 (O_5,N_29393,N_29361);
xnor UO_6 (O_6,N_28968,N_29202);
xnor UO_7 (O_7,N_29417,N_25588);
nor UO_8 (O_8,N_28660,N_28658);
nand UO_9 (O_9,N_27708,N_29205);
or UO_10 (O_10,N_27570,N_26958);
nor UO_11 (O_11,N_26201,N_29043);
nand UO_12 (O_12,N_25995,N_29036);
xor UO_13 (O_13,N_26229,N_26785);
or UO_14 (O_14,N_27883,N_26365);
and UO_15 (O_15,N_26484,N_28380);
nand UO_16 (O_16,N_26513,N_28400);
xor UO_17 (O_17,N_28457,N_25419);
nand UO_18 (O_18,N_29892,N_27845);
or UO_19 (O_19,N_28464,N_27656);
and UO_20 (O_20,N_25497,N_29444);
xnor UO_21 (O_21,N_26611,N_29551);
nor UO_22 (O_22,N_29875,N_29402);
xnor UO_23 (O_23,N_28750,N_25884);
and UO_24 (O_24,N_27319,N_28482);
or UO_25 (O_25,N_25727,N_27584);
and UO_26 (O_26,N_26447,N_29323);
nor UO_27 (O_27,N_27162,N_26178);
nor UO_28 (O_28,N_25091,N_29163);
nand UO_29 (O_29,N_25992,N_27258);
and UO_30 (O_30,N_25404,N_29459);
nor UO_31 (O_31,N_25334,N_26974);
xnor UO_32 (O_32,N_27265,N_29285);
and UO_33 (O_33,N_26502,N_27642);
or UO_34 (O_34,N_25962,N_25406);
xnor UO_35 (O_35,N_27448,N_27715);
xor UO_36 (O_36,N_25658,N_26890);
and UO_37 (O_37,N_27658,N_28070);
nor UO_38 (O_38,N_28440,N_28358);
nor UO_39 (O_39,N_29179,N_27219);
or UO_40 (O_40,N_25433,N_26246);
nor UO_41 (O_41,N_25200,N_27490);
or UO_42 (O_42,N_28107,N_27901);
and UO_43 (O_43,N_25759,N_25247);
or UO_44 (O_44,N_25609,N_26211);
nor UO_45 (O_45,N_27796,N_26427);
xnor UO_46 (O_46,N_25869,N_27864);
and UO_47 (O_47,N_26358,N_29501);
nor UO_48 (O_48,N_27235,N_29208);
nand UO_49 (O_49,N_26571,N_28251);
xnor UO_50 (O_50,N_26522,N_28198);
xor UO_51 (O_51,N_27723,N_29616);
xnor UO_52 (O_52,N_25624,N_27014);
and UO_53 (O_53,N_28415,N_27176);
or UO_54 (O_54,N_28870,N_25225);
or UO_55 (O_55,N_28035,N_28797);
nand UO_56 (O_56,N_28887,N_28231);
xor UO_57 (O_57,N_27260,N_27602);
and UO_58 (O_58,N_26405,N_27418);
or UO_59 (O_59,N_29269,N_27193);
nor UO_60 (O_60,N_29692,N_27984);
nand UO_61 (O_61,N_27142,N_28915);
nand UO_62 (O_62,N_27679,N_28616);
and UO_63 (O_63,N_28071,N_28328);
nor UO_64 (O_64,N_28523,N_29870);
and UO_65 (O_65,N_29856,N_27902);
xor UO_66 (O_66,N_25029,N_29093);
nand UO_67 (O_67,N_29087,N_25523);
xnor UO_68 (O_68,N_27197,N_25399);
or UO_69 (O_69,N_25720,N_28486);
nand UO_70 (O_70,N_26384,N_28346);
nand UO_71 (O_71,N_29528,N_27112);
xor UO_72 (O_72,N_27590,N_26177);
and UO_73 (O_73,N_29084,N_27023);
nor UO_74 (O_74,N_25876,N_27420);
nand UO_75 (O_75,N_27261,N_27056);
nor UO_76 (O_76,N_26896,N_26337);
nand UO_77 (O_77,N_29288,N_25753);
or UO_78 (O_78,N_26830,N_25361);
nand UO_79 (O_79,N_27930,N_28253);
and UO_80 (O_80,N_25871,N_29407);
and UO_81 (O_81,N_26776,N_25826);
and UO_82 (O_82,N_26908,N_27093);
or UO_83 (O_83,N_25474,N_29320);
nor UO_84 (O_84,N_29681,N_25765);
xor UO_85 (O_85,N_25343,N_26921);
or UO_86 (O_86,N_25654,N_27588);
nand UO_87 (O_87,N_25709,N_25887);
xnor UO_88 (O_88,N_29236,N_26321);
nand UO_89 (O_89,N_27704,N_25446);
and UO_90 (O_90,N_29369,N_28869);
nor UO_91 (O_91,N_25304,N_26375);
or UO_92 (O_92,N_26560,N_26909);
xnor UO_93 (O_93,N_26023,N_26910);
xor UO_94 (O_94,N_27717,N_26757);
and UO_95 (O_95,N_29447,N_28683);
nor UO_96 (O_96,N_27810,N_27196);
nand UO_97 (O_97,N_28962,N_27172);
nand UO_98 (O_98,N_28708,N_28285);
xnor UO_99 (O_99,N_26968,N_25283);
xor UO_100 (O_100,N_28418,N_28094);
and UO_101 (O_101,N_27218,N_27863);
or UO_102 (O_102,N_26866,N_28734);
and UO_103 (O_103,N_28883,N_25987);
or UO_104 (O_104,N_28377,N_28850);
nand UO_105 (O_105,N_27557,N_26149);
nor UO_106 (O_106,N_25662,N_27151);
and UO_107 (O_107,N_27101,N_27394);
nand UO_108 (O_108,N_26193,N_26243);
nand UO_109 (O_109,N_25472,N_26312);
and UO_110 (O_110,N_26225,N_29900);
xor UO_111 (O_111,N_25859,N_27545);
or UO_112 (O_112,N_27586,N_26683);
or UO_113 (O_113,N_29063,N_27647);
nor UO_114 (O_114,N_26599,N_27856);
nand UO_115 (O_115,N_28884,N_27956);
nand UO_116 (O_116,N_27664,N_27379);
nand UO_117 (O_117,N_25599,N_28643);
nor UO_118 (O_118,N_29325,N_27039);
or UO_119 (O_119,N_28038,N_29289);
and UO_120 (O_120,N_26079,N_27285);
or UO_121 (O_121,N_26763,N_25597);
nor UO_122 (O_122,N_26441,N_29070);
or UO_123 (O_123,N_25882,N_29086);
nor UO_124 (O_124,N_29675,N_29316);
xnor UO_125 (O_125,N_27412,N_28714);
nand UO_126 (O_126,N_25217,N_27225);
xor UO_127 (O_127,N_28012,N_27215);
xnor UO_128 (O_128,N_26999,N_27478);
and UO_129 (O_129,N_26873,N_26794);
xnor UO_130 (O_130,N_25619,N_28450);
xor UO_131 (O_131,N_28446,N_27009);
and UO_132 (O_132,N_26829,N_26736);
nor UO_133 (O_133,N_27955,N_26542);
or UO_134 (O_134,N_26681,N_26073);
xnor UO_135 (O_135,N_27690,N_29431);
xnor UO_136 (O_136,N_29116,N_25355);
or UO_137 (O_137,N_27061,N_26378);
or UO_138 (O_138,N_27734,N_26996);
or UO_139 (O_139,N_25006,N_27538);
nand UO_140 (O_140,N_26477,N_28858);
nor UO_141 (O_141,N_26479,N_29074);
and UO_142 (O_142,N_25603,N_27696);
nor UO_143 (O_143,N_25848,N_25927);
or UO_144 (O_144,N_29371,N_28013);
nor UO_145 (O_145,N_27026,N_26418);
or UO_146 (O_146,N_26342,N_25023);
nand UO_147 (O_147,N_28972,N_26732);
and UO_148 (O_148,N_29143,N_26005);
and UO_149 (O_149,N_28008,N_28654);
and UO_150 (O_150,N_26644,N_29618);
or UO_151 (O_151,N_25818,N_28156);
xnor UO_152 (O_152,N_26902,N_25965);
and UO_153 (O_153,N_26582,N_25596);
nor UO_154 (O_154,N_27019,N_27029);
nor UO_155 (O_155,N_27236,N_27695);
nor UO_156 (O_156,N_26602,N_25566);
xor UO_157 (O_157,N_26624,N_28599);
and UO_158 (O_158,N_27800,N_25844);
or UO_159 (O_159,N_29854,N_27848);
or UO_160 (O_160,N_25671,N_27416);
nand UO_161 (O_161,N_25099,N_28257);
xnor UO_162 (O_162,N_28526,N_25739);
or UO_163 (O_163,N_28103,N_26435);
nor UO_164 (O_164,N_26099,N_26898);
nor UO_165 (O_165,N_27686,N_25112);
nor UO_166 (O_166,N_25109,N_26221);
or UO_167 (O_167,N_27229,N_25241);
or UO_168 (O_168,N_27034,N_28731);
and UO_169 (O_169,N_28437,N_27119);
and UO_170 (O_170,N_29984,N_29621);
nor UO_171 (O_171,N_28501,N_26165);
and UO_172 (O_172,N_25194,N_28067);
nor UO_173 (O_173,N_25274,N_26617);
nand UO_174 (O_174,N_29295,N_28987);
and UO_175 (O_175,N_26381,N_28260);
and UO_176 (O_176,N_29889,N_27812);
nor UO_177 (O_177,N_26042,N_26145);
nor UO_178 (O_178,N_25368,N_29919);
or UO_179 (O_179,N_29249,N_28164);
and UO_180 (O_180,N_27605,N_27498);
or UO_181 (O_181,N_28002,N_25617);
nor UO_182 (O_182,N_25953,N_26704);
and UO_183 (O_183,N_25829,N_28955);
xnor UO_184 (O_184,N_29643,N_26360);
and UO_185 (O_185,N_26938,N_28097);
and UO_186 (O_186,N_25397,N_26702);
and UO_187 (O_187,N_25989,N_27890);
or UO_188 (O_188,N_27910,N_29281);
and UO_189 (O_189,N_27731,N_28529);
nand UO_190 (O_190,N_29510,N_27541);
nor UO_191 (O_191,N_26595,N_28354);
and UO_192 (O_192,N_28846,N_29917);
nor UO_193 (O_193,N_29630,N_29071);
nand UO_194 (O_194,N_29965,N_29506);
and UO_195 (O_195,N_29581,N_26865);
xnor UO_196 (O_196,N_29301,N_28502);
nand UO_197 (O_197,N_27514,N_28997);
nor UO_198 (O_198,N_28027,N_25010);
xor UO_199 (O_199,N_26392,N_26603);
nand UO_200 (O_200,N_28689,N_26678);
or UO_201 (O_201,N_27702,N_25684);
and UO_202 (O_202,N_26296,N_27778);
nand UO_203 (O_203,N_27371,N_25439);
xor UO_204 (O_204,N_25268,N_25713);
or UO_205 (O_205,N_27608,N_27736);
and UO_206 (O_206,N_27899,N_28514);
and UO_207 (O_207,N_25550,N_29363);
xor UO_208 (O_208,N_29136,N_29791);
xnor UO_209 (O_209,N_28867,N_27638);
or UO_210 (O_210,N_26848,N_26469);
and UO_211 (O_211,N_28622,N_29026);
and UO_212 (O_212,N_26182,N_29005);
nor UO_213 (O_213,N_27949,N_28715);
nor UO_214 (O_214,N_29536,N_28556);
nor UO_215 (O_215,N_29037,N_27456);
nor UO_216 (O_216,N_25388,N_26333);
or UO_217 (O_217,N_27222,N_29662);
and UO_218 (O_218,N_29048,N_28385);
nor UO_219 (O_219,N_29461,N_29445);
and UO_220 (O_220,N_29016,N_26416);
and UO_221 (O_221,N_25245,N_27592);
and UO_222 (O_222,N_29319,N_27402);
xnor UO_223 (O_223,N_25712,N_25934);
or UO_224 (O_224,N_29066,N_26199);
xnor UO_225 (O_225,N_27583,N_29736);
xor UO_226 (O_226,N_28911,N_28311);
nor UO_227 (O_227,N_27935,N_26457);
or UO_228 (O_228,N_29674,N_27515);
nor UO_229 (O_229,N_26555,N_25578);
xor UO_230 (O_230,N_29644,N_29851);
nand UO_231 (O_231,N_29709,N_29129);
nand UO_232 (O_232,N_25246,N_26738);
or UO_233 (O_233,N_27031,N_27944);
nor UO_234 (O_234,N_26942,N_29180);
or UO_235 (O_235,N_25847,N_29822);
nor UO_236 (O_236,N_29985,N_26798);
or UO_237 (O_237,N_28995,N_26911);
nand UO_238 (O_238,N_29812,N_27269);
nor UO_239 (O_239,N_27669,N_25401);
and UO_240 (O_240,N_27512,N_26289);
xor UO_241 (O_241,N_26626,N_26121);
nand UO_242 (O_242,N_25754,N_26656);
and UO_243 (O_243,N_27079,N_26129);
nor UO_244 (O_244,N_26092,N_27170);
xnor UO_245 (O_245,N_29771,N_28859);
nand UO_246 (O_246,N_25453,N_25986);
xnor UO_247 (O_247,N_29195,N_25798);
nor UO_248 (O_248,N_27655,N_28906);
or UO_249 (O_249,N_26450,N_28563);
and UO_250 (O_250,N_29126,N_27182);
xnor UO_251 (O_251,N_27415,N_25340);
and UO_252 (O_252,N_25849,N_29031);
nand UO_253 (O_253,N_29811,N_27594);
or UO_254 (O_254,N_27133,N_28037);
nor UO_255 (O_255,N_26818,N_29803);
nor UO_256 (O_256,N_28936,N_28001);
and UO_257 (O_257,N_29602,N_28109);
nand UO_258 (O_258,N_27979,N_26060);
and UO_259 (O_259,N_26114,N_26979);
and UO_260 (O_260,N_28227,N_28417);
or UO_261 (O_261,N_29305,N_25137);
nor UO_262 (O_262,N_29814,N_28119);
xnor UO_263 (O_263,N_29555,N_28165);
and UO_264 (O_264,N_26294,N_25152);
and UO_265 (O_265,N_27872,N_25900);
xor UO_266 (O_266,N_27759,N_28876);
nand UO_267 (O_267,N_25428,N_26284);
xnor UO_268 (O_268,N_28706,N_28294);
nor UO_269 (O_269,N_29543,N_29708);
xor UO_270 (O_270,N_25297,N_27967);
or UO_271 (O_271,N_28748,N_25998);
xor UO_272 (O_272,N_26947,N_25155);
xor UO_273 (O_273,N_26847,N_26329);
nor UO_274 (O_274,N_25776,N_29523);
nand UO_275 (O_275,N_28180,N_27429);
and UO_276 (O_276,N_28712,N_27818);
nor UO_277 (O_277,N_29092,N_26003);
xor UO_278 (O_278,N_28639,N_26147);
nor UO_279 (O_279,N_27572,N_29580);
nand UO_280 (O_280,N_28934,N_28412);
nor UO_281 (O_281,N_25298,N_27621);
nand UO_282 (O_282,N_27414,N_26837);
or UO_283 (O_283,N_27068,N_29106);
or UO_284 (O_284,N_25630,N_25956);
nand UO_285 (O_285,N_28776,N_29122);
xor UO_286 (O_286,N_28626,N_28146);
nor UO_287 (O_287,N_28894,N_25567);
nor UO_288 (O_288,N_29415,N_26609);
and UO_289 (O_289,N_26103,N_27343);
xor UO_290 (O_290,N_28844,N_29167);
and UO_291 (O_291,N_29650,N_28447);
or UO_292 (O_292,N_29482,N_29585);
xor UO_293 (O_293,N_29570,N_29411);
nor UO_294 (O_294,N_28878,N_29717);
xnor UO_295 (O_295,N_25158,N_25809);
nor UO_296 (O_296,N_26639,N_25950);
nor UO_297 (O_297,N_26916,N_25094);
nand UO_298 (O_298,N_25434,N_29833);
and UO_299 (O_299,N_26547,N_27296);
xor UO_300 (O_300,N_26623,N_27318);
or UO_301 (O_301,N_25352,N_28549);
or UO_302 (O_302,N_26945,N_29437);
nor UO_303 (O_303,N_25376,N_29428);
nand UO_304 (O_304,N_25269,N_26089);
and UO_305 (O_305,N_26980,N_27393);
or UO_306 (O_306,N_29255,N_29409);
and UO_307 (O_307,N_25276,N_28709);
xor UO_308 (O_308,N_27975,N_28247);
nand UO_309 (O_309,N_25092,N_28981);
xor UO_310 (O_310,N_29552,N_28537);
nor UO_311 (O_311,N_29209,N_25301);
xnor UO_312 (O_312,N_27190,N_29133);
and UO_313 (O_313,N_27641,N_26382);
or UO_314 (O_314,N_25050,N_27086);
and UO_315 (O_315,N_26748,N_26081);
xnor UO_316 (O_316,N_27110,N_28342);
nand UO_317 (O_317,N_29112,N_28738);
xnor UO_318 (O_318,N_28416,N_29292);
xor UO_319 (O_319,N_25885,N_29328);
nand UO_320 (O_320,N_26929,N_28895);
xor UO_321 (O_321,N_25808,N_27614);
xor UO_322 (O_322,N_27918,N_28596);
nor UO_323 (O_323,N_29750,N_25792);
nor UO_324 (O_324,N_25448,N_25024);
nor UO_325 (O_325,N_26948,N_28275);
or UO_326 (O_326,N_26057,N_29800);
and UO_327 (O_327,N_29671,N_27965);
nand UO_328 (O_328,N_28186,N_26606);
xor UO_329 (O_329,N_28226,N_26552);
nand UO_330 (O_330,N_26912,N_25057);
and UO_331 (O_331,N_29924,N_25466);
or UO_332 (O_332,N_26297,N_28816);
and UO_333 (O_333,N_28133,N_28885);
or UO_334 (O_334,N_27003,N_29384);
or UO_335 (O_335,N_25761,N_28589);
or UO_336 (O_336,N_29680,N_25003);
nand UO_337 (O_337,N_28000,N_29219);
and UO_338 (O_338,N_26927,N_28522);
nor UO_339 (O_339,N_27740,N_27064);
xnor UO_340 (O_340,N_26207,N_25275);
nor UO_341 (O_341,N_26585,N_25103);
xnor UO_342 (O_342,N_26868,N_29574);
and UO_343 (O_343,N_26307,N_26357);
xnor UO_344 (O_344,N_29313,N_27062);
and UO_345 (O_345,N_27551,N_27861);
xor UO_346 (O_346,N_28413,N_29769);
nor UO_347 (O_347,N_28703,N_27568);
or UO_348 (O_348,N_27832,N_26701);
nand UO_349 (O_349,N_25892,N_29367);
and UO_350 (O_350,N_29819,N_27113);
and UO_351 (O_351,N_28839,N_27687);
nand UO_352 (O_352,N_27733,N_25613);
nand UO_353 (O_353,N_26616,N_27326);
xor UO_354 (O_354,N_28312,N_27482);
xnor UO_355 (O_355,N_27785,N_25004);
or UO_356 (O_356,N_27510,N_26462);
nand UO_357 (O_357,N_29089,N_26588);
and UO_358 (O_358,N_25178,N_26975);
xor UO_359 (O_359,N_27879,N_28806);
xnor UO_360 (O_360,N_28980,N_29562);
nor UO_361 (O_361,N_26150,N_27105);
nor UO_362 (O_362,N_27829,N_29840);
xor UO_363 (O_363,N_26541,N_26671);
xor UO_364 (O_364,N_26467,N_26721);
nor UO_365 (O_365,N_26412,N_26925);
nand UO_366 (O_366,N_25312,N_26593);
nor UO_367 (O_367,N_26914,N_26490);
xor UO_368 (O_368,N_27537,N_29563);
and UO_369 (O_369,N_26710,N_27248);
nor UO_370 (O_370,N_27012,N_29608);
or UO_371 (O_371,N_25438,N_25110);
xnor UO_372 (O_372,N_28280,N_26863);
or UO_373 (O_373,N_27206,N_28462);
nor UO_374 (O_374,N_28079,N_25536);
nor UO_375 (O_375,N_28106,N_29573);
nand UO_376 (O_376,N_26119,N_29332);
xnor UO_377 (O_377,N_25483,N_29583);
nor UO_378 (O_378,N_27253,N_26728);
nor UO_379 (O_379,N_29741,N_27834);
xor UO_380 (O_380,N_25173,N_29049);
or UO_381 (O_381,N_29120,N_28893);
xor UO_382 (O_382,N_26459,N_26401);
nor UO_383 (O_383,N_26670,N_28136);
and UO_384 (O_384,N_29279,N_25125);
and UO_385 (O_385,N_27065,N_25602);
and UO_386 (O_386,N_25034,N_29438);
and UO_387 (O_387,N_29137,N_29619);
and UO_388 (O_388,N_26161,N_29025);
xor UO_389 (O_389,N_25175,N_25515);
xnor UO_390 (O_390,N_29162,N_29507);
nand UO_391 (O_391,N_26148,N_25394);
nor UO_392 (O_392,N_28252,N_28834);
or UO_393 (O_393,N_29879,N_29718);
nor UO_394 (O_394,N_26063,N_27574);
or UO_395 (O_395,N_27938,N_27223);
and UO_396 (O_396,N_29184,N_25445);
nor UO_397 (O_397,N_27180,N_28054);
and UO_398 (O_398,N_29704,N_28498);
nor UO_399 (O_399,N_29233,N_29535);
xnor UO_400 (O_400,N_28579,N_25834);
nor UO_401 (O_401,N_25387,N_29511);
and UO_402 (O_402,N_27509,N_28115);
xor UO_403 (O_403,N_25559,N_26471);
xor UO_404 (O_404,N_28336,N_26138);
nor UO_405 (O_405,N_29469,N_29189);
nand UO_406 (O_406,N_25943,N_27615);
or UO_407 (O_407,N_28686,N_25345);
xnor UO_408 (O_408,N_28384,N_25842);
or UO_409 (O_409,N_26966,N_29142);
xnor UO_410 (O_410,N_25918,N_28242);
xnor UO_411 (O_411,N_27092,N_26510);
xnor UO_412 (O_412,N_27722,N_27880);
or UO_413 (O_413,N_26128,N_25947);
and UO_414 (O_414,N_25941,N_29916);
xnor UO_415 (O_415,N_25585,N_25317);
nor UO_416 (O_416,N_27808,N_29374);
nor UO_417 (O_417,N_27838,N_26044);
and UO_418 (O_418,N_29982,N_25413);
and UO_419 (O_419,N_28456,N_25393);
nor UO_420 (O_420,N_27960,N_25048);
xor UO_421 (O_421,N_29419,N_25743);
and UO_422 (O_422,N_25942,N_28477);
nor UO_423 (O_423,N_28154,N_26027);
nand UO_424 (O_424,N_25086,N_29028);
and UO_425 (O_425,N_25915,N_25456);
or UO_426 (O_426,N_28082,N_25000);
nand UO_427 (O_427,N_26242,N_27929);
xnor UO_428 (O_428,N_27606,N_28988);
xnor UO_429 (O_429,N_27657,N_28974);
and UO_430 (O_430,N_25652,N_27617);
xnor UO_431 (O_431,N_29270,N_26176);
nor UO_432 (O_432,N_29828,N_26105);
or UO_433 (O_433,N_26587,N_26117);
nor UO_434 (O_434,N_28408,N_29429);
xnor UO_435 (O_435,N_26400,N_27238);
xnor UO_436 (O_436,N_25074,N_29705);
or UO_437 (O_437,N_26833,N_27966);
and UO_438 (O_438,N_25382,N_27611);
and UO_439 (O_439,N_29390,N_27814);
nor UO_440 (O_440,N_27015,N_26781);
nor UO_441 (O_441,N_28078,N_25349);
xor UO_442 (O_442,N_26247,N_25243);
xor UO_443 (O_443,N_28753,N_29972);
nor UO_444 (O_444,N_26526,N_25416);
nor UO_445 (O_445,N_26796,N_29935);
and UO_446 (O_446,N_25698,N_29891);
or UO_447 (O_447,N_25669,N_28249);
nand UO_448 (O_448,N_26920,N_26677);
nor UO_449 (O_449,N_27072,N_29841);
nand UO_450 (O_450,N_26222,N_28817);
or UO_451 (O_451,N_27220,N_27524);
nor UO_452 (O_452,N_29809,N_29829);
xor UO_453 (O_453,N_26167,N_27873);
xor UO_454 (O_454,N_28979,N_28258);
nor UO_455 (O_455,N_28190,N_29051);
nand UO_456 (O_456,N_26851,N_27575);
nor UO_457 (O_457,N_26108,N_28073);
nor UO_458 (O_458,N_28566,N_28527);
or UO_459 (O_459,N_28825,N_26152);
nor UO_460 (O_460,N_28835,N_28487);
or UO_461 (O_461,N_29915,N_28454);
or UO_462 (O_462,N_27751,N_25375);
and UO_463 (O_463,N_27550,N_25678);
and UO_464 (O_464,N_25210,N_26420);
nor UO_465 (O_465,N_29000,N_28497);
and UO_466 (O_466,N_29353,N_27203);
or UO_467 (O_467,N_29383,N_28395);
nor UO_468 (O_468,N_26126,N_29350);
or UO_469 (O_469,N_27457,N_27970);
or UO_470 (O_470,N_26933,N_29201);
nor UO_471 (O_471,N_28810,N_27480);
and UO_472 (O_472,N_25486,N_26046);
nand UO_473 (O_473,N_25628,N_27505);
and UO_474 (O_474,N_28960,N_29186);
xor UO_475 (O_475,N_28657,N_28396);
nor UO_476 (O_476,N_26335,N_29962);
nand UO_477 (O_477,N_26112,N_28234);
or UO_478 (O_478,N_25066,N_25161);
nor UO_479 (O_479,N_29584,N_29685);
nor UO_480 (O_480,N_29654,N_25664);
or UO_481 (O_481,N_28239,N_26989);
xor UO_482 (O_482,N_25513,N_25539);
and UO_483 (O_483,N_26577,N_29192);
or UO_484 (O_484,N_28552,N_26354);
xor UO_485 (O_485,N_27000,N_27836);
and UO_486 (O_486,N_27153,N_26518);
or UO_487 (O_487,N_27802,N_29321);
or UO_488 (O_488,N_25093,N_29941);
nand UO_489 (O_489,N_26004,N_28646);
and UO_490 (O_490,N_28667,N_27302);
nand UO_491 (O_491,N_28304,N_27817);
nand UO_492 (O_492,N_26430,N_29657);
xor UO_493 (O_493,N_28325,N_28187);
nor UO_494 (O_494,N_27920,N_29597);
nor UO_495 (O_495,N_29273,N_29577);
nand UO_496 (O_496,N_28003,N_27948);
or UO_497 (O_497,N_29146,N_27988);
xnor UO_498 (O_498,N_27694,N_25823);
nand UO_499 (O_499,N_27764,N_29725);
nand UO_500 (O_500,N_29238,N_26218);
xnor UO_501 (O_501,N_25746,N_27522);
and UO_502 (O_502,N_29781,N_25281);
nand UO_503 (O_503,N_26276,N_25725);
or UO_504 (O_504,N_27782,N_26698);
and UO_505 (O_505,N_25756,N_26647);
or UO_506 (O_506,N_27174,N_29022);
nor UO_507 (O_507,N_25586,N_25360);
xnor UO_508 (O_508,N_26517,N_25148);
nor UO_509 (O_509,N_29241,N_25287);
xor UO_510 (O_510,N_28754,N_29156);
nor UO_511 (O_511,N_27511,N_29914);
nor UO_512 (O_512,N_25396,N_26694);
xnor UO_513 (O_513,N_28744,N_25493);
nand UO_514 (O_514,N_25136,N_25102);
nand UO_515 (O_515,N_25377,N_25997);
and UO_516 (O_516,N_25499,N_25171);
or UO_517 (O_517,N_27531,N_29612);
xor UO_518 (O_518,N_29520,N_28168);
or UO_519 (O_519,N_25059,N_25068);
and UO_520 (O_520,N_26960,N_29886);
xor UO_521 (O_521,N_28814,N_26836);
and UO_522 (O_522,N_27911,N_28388);
or UO_523 (O_523,N_29212,N_25799);
or UO_524 (O_524,N_28625,N_27396);
nor UO_525 (O_525,N_27451,N_25675);
or UO_526 (O_526,N_29798,N_28954);
xnor UO_527 (O_527,N_29450,N_27578);
nand UO_528 (O_528,N_28381,N_28856);
xor UO_529 (O_529,N_26185,N_25556);
nor UO_530 (O_530,N_27725,N_29387);
nor UO_531 (O_531,N_27573,N_28977);
nor UO_532 (O_532,N_29046,N_29243);
nor UO_533 (O_533,N_25790,N_26531);
nor UO_534 (O_534,N_29850,N_26731);
or UO_535 (O_535,N_25740,N_27630);
xor UO_536 (O_536,N_25702,N_27987);
or UO_537 (O_537,N_26041,N_29107);
and UO_538 (O_538,N_26424,N_29091);
and UO_539 (O_539,N_28085,N_27906);
xor UO_540 (O_540,N_26561,N_28882);
nor UO_541 (O_541,N_26767,N_29754);
nor UO_542 (O_542,N_26220,N_29380);
or UO_543 (O_543,N_28047,N_26433);
nor UO_544 (O_544,N_27436,N_28888);
xor UO_545 (O_545,N_26488,N_29442);
nand UO_546 (O_546,N_29069,N_26969);
and UO_547 (O_547,N_26095,N_26771);
or UO_548 (O_548,N_26376,N_28910);
nand UO_549 (O_549,N_28036,N_25521);
xnor UO_550 (O_550,N_26772,N_26621);
or UO_551 (O_551,N_29446,N_29748);
xnor UO_552 (O_552,N_27866,N_27772);
nand UO_553 (O_553,N_26308,N_25895);
or UO_554 (O_554,N_27652,N_25151);
xnor UO_555 (O_555,N_29954,N_29902);
xnor UO_556 (O_556,N_28364,N_28015);
nor UO_557 (O_557,N_28794,N_26846);
nor UO_558 (O_558,N_25160,N_26071);
or UO_559 (O_559,N_29923,N_29226);
nor UO_560 (O_560,N_28718,N_28393);
nor UO_561 (O_561,N_29277,N_28819);
nand UO_562 (O_562,N_25025,N_28404);
nor UO_563 (O_563,N_29435,N_28765);
or UO_564 (O_564,N_29403,N_27523);
and UO_565 (O_565,N_26391,N_27329);
or UO_566 (O_566,N_29111,N_29177);
nor UO_567 (O_567,N_28533,N_25321);
and UO_568 (O_568,N_27465,N_25665);
and UO_569 (O_569,N_27250,N_29790);
or UO_570 (O_570,N_25633,N_27213);
xor UO_571 (O_571,N_27312,N_25323);
and UO_572 (O_572,N_26859,N_25810);
nor UO_573 (O_573,N_26876,N_26120);
or UO_574 (O_574,N_29877,N_26087);
and UO_575 (O_575,N_27707,N_29634);
xnor UO_576 (O_576,N_25543,N_28143);
and UO_577 (O_577,N_29149,N_28763);
or UO_578 (O_578,N_29525,N_25666);
nor UO_579 (O_579,N_26931,N_28268);
nand UO_580 (O_580,N_27757,N_29569);
xnor UO_581 (O_581,N_28751,N_29307);
nand UO_582 (O_582,N_25039,N_25314);
and UO_583 (O_583,N_28046,N_28110);
nand UO_584 (O_584,N_29679,N_28099);
and UO_585 (O_585,N_26637,N_26202);
xnor UO_586 (O_586,N_26699,N_26840);
and UO_587 (O_587,N_26810,N_25335);
nand UO_588 (O_588,N_28219,N_29933);
and UO_589 (O_589,N_29477,N_26649);
nor UO_590 (O_590,N_26153,N_26714);
nand UO_591 (O_591,N_26867,N_29050);
nor UO_592 (O_592,N_25459,N_27828);
nor UO_593 (O_593,N_28310,N_28976);
nand UO_594 (O_594,N_29542,N_28340);
and UO_595 (O_595,N_29689,N_27789);
xnor UO_596 (O_596,N_26667,N_25289);
and UO_597 (O_597,N_29694,N_26913);
nor UO_598 (O_598,N_25409,N_26000);
nand UO_599 (O_599,N_27900,N_28939);
and UO_600 (O_600,N_28719,N_25511);
xor UO_601 (O_601,N_29259,N_26156);
xor UO_602 (O_602,N_26862,N_28746);
or UO_603 (O_603,N_29047,N_25014);
nor UO_604 (O_604,N_27990,N_29855);
and UO_605 (O_605,N_25477,N_28889);
xnor UO_606 (O_606,N_25667,N_26596);
xor UO_607 (O_607,N_27981,N_28049);
xnor UO_608 (O_608,N_27937,N_29100);
nor UO_609 (O_609,N_25398,N_29247);
or UO_610 (O_610,N_28640,N_25249);
xor UO_611 (O_611,N_25570,N_27292);
and UO_612 (O_612,N_26919,N_28308);
nor UO_613 (O_613,N_27275,N_28397);
and UO_614 (O_614,N_25612,N_29715);
nand UO_615 (O_615,N_25108,N_27390);
xor UO_616 (O_616,N_29695,N_29947);
nand UO_617 (O_617,N_29733,N_26788);
or UO_618 (O_618,N_29365,N_25035);
and UO_619 (O_619,N_28237,N_29866);
nand UO_620 (O_620,N_26259,N_26695);
nor UO_621 (O_621,N_27827,N_28363);
or UO_622 (O_622,N_28273,N_28595);
or UO_623 (O_623,N_28407,N_28240);
and UO_624 (O_624,N_26409,N_28445);
nand UO_625 (O_625,N_26566,N_25498);
or UO_626 (O_626,N_29789,N_26532);
nand UO_627 (O_627,N_28448,N_28574);
and UO_628 (O_628,N_28578,N_29197);
and UO_629 (O_629,N_29003,N_27534);
or UO_630 (O_630,N_29948,N_28830);
nor UO_631 (O_631,N_29424,N_28682);
xnor UO_632 (O_632,N_25085,N_27137);
and UO_633 (O_633,N_29742,N_26643);
nor UO_634 (O_634,N_25372,N_25165);
nor UO_635 (O_635,N_27972,N_26675);
and UO_636 (O_636,N_27886,N_26495);
or UO_637 (O_637,N_25768,N_26397);
or UO_638 (O_638,N_28431,N_29989);
nand UO_639 (O_639,N_29073,N_26527);
xnor UO_640 (O_640,N_26696,N_27527);
nor UO_641 (O_641,N_25028,N_26986);
nor UO_642 (O_642,N_29375,N_26250);
and UO_643 (O_643,N_26632,N_26184);
nor UO_644 (O_644,N_28785,N_29728);
or UO_645 (O_645,N_27618,N_29139);
xnor UO_646 (O_646,N_26483,N_29466);
and UO_647 (O_647,N_26066,N_28499);
and UO_648 (O_648,N_27805,N_26514);
nand UO_649 (O_649,N_28194,N_27486);
or UO_650 (O_650,N_27425,N_25016);
xnor UO_651 (O_651,N_28619,N_28843);
nor UO_652 (O_652,N_29519,N_28973);
and UO_653 (O_653,N_25512,N_29860);
xnor UO_654 (O_654,N_28601,N_29055);
and UO_655 (O_655,N_27471,N_25075);
nand UO_656 (O_656,N_25378,N_26516);
nand UO_657 (O_657,N_28438,N_29844);
xnor UO_658 (O_658,N_28842,N_26144);
nor UO_659 (O_659,N_29966,N_28700);
or UO_660 (O_660,N_25021,N_25971);
nand UO_661 (O_661,N_27701,N_26586);
nand UO_662 (O_662,N_26729,N_26515);
or UO_663 (O_663,N_25206,N_25901);
nand UO_664 (O_664,N_25679,N_25751);
or UO_665 (O_665,N_27591,N_27066);
xnor UO_666 (O_666,N_29082,N_25858);
xor UO_667 (O_667,N_27738,N_29169);
nand UO_668 (O_668,N_26098,N_25182);
and UO_669 (O_669,N_29611,N_25555);
nand UO_670 (O_670,N_26834,N_26937);
nor UO_671 (O_671,N_28287,N_25629);
nor UO_672 (O_672,N_25076,N_26351);
and UO_673 (O_673,N_25518,N_28929);
xnor UO_674 (O_674,N_26805,N_29468);
xor UO_675 (O_675,N_29213,N_27971);
nor UO_676 (O_676,N_28214,N_28017);
and UO_677 (O_677,N_28161,N_29687);
xnor UO_678 (O_678,N_28163,N_28841);
nor UO_679 (O_679,N_28236,N_28353);
or UO_680 (O_680,N_25470,N_29835);
nor UO_681 (O_681,N_25747,N_25157);
nand UO_682 (O_682,N_26991,N_29955);
xor UO_683 (O_683,N_26319,N_26750);
nor UO_684 (O_684,N_29347,N_27347);
or UO_685 (O_685,N_25222,N_25408);
and UO_686 (O_686,N_27692,N_27912);
or UO_687 (O_687,N_25199,N_29714);
xnor UO_688 (O_688,N_27132,N_27720);
or UO_689 (O_689,N_27484,N_26480);
and UO_690 (O_690,N_25861,N_26191);
xnor UO_691 (O_691,N_26449,N_29496);
or UO_692 (O_692,N_27579,N_27317);
nand UO_693 (O_693,N_28383,N_29970);
nor UO_694 (O_694,N_27876,N_26348);
xnor UO_695 (O_695,N_26760,N_26583);
nor UO_696 (O_696,N_28760,N_25935);
or UO_697 (O_697,N_25229,N_29959);
and UO_698 (O_698,N_26343,N_27766);
and UO_699 (O_699,N_28826,N_29837);
or UO_700 (O_700,N_28374,N_25526);
and UO_701 (O_701,N_26151,N_27387);
or UO_702 (O_702,N_28056,N_29757);
or UO_703 (O_703,N_27299,N_29494);
nor UO_704 (O_704,N_26832,N_29842);
nor UO_705 (O_705,N_26858,N_28673);
nor UO_706 (O_706,N_25909,N_29888);
and UO_707 (O_707,N_29792,N_26174);
or UO_708 (O_708,N_25139,N_26752);
nor UO_709 (O_709,N_28182,N_28624);
or UO_710 (O_710,N_27087,N_28875);
nor UO_711 (O_711,N_25945,N_27869);
xnor UO_712 (O_712,N_25204,N_27926);
nand UO_713 (O_713,N_29294,N_25379);
xor UO_714 (O_714,N_25828,N_25285);
xor UO_715 (O_715,N_27085,N_26627);
xnor UO_716 (O_716,N_29593,N_29436);
and UO_717 (O_717,N_29926,N_26745);
nand UO_718 (O_718,N_27107,N_29802);
xnor UO_719 (O_719,N_25681,N_25936);
nand UO_720 (O_720,N_28941,N_29623);
nor UO_721 (O_721,N_28178,N_25073);
nor UO_722 (O_722,N_28392,N_26700);
and UO_723 (O_723,N_29227,N_26625);
or UO_724 (O_724,N_26429,N_29336);
xnor UO_725 (O_725,N_28773,N_28986);
nor UO_726 (O_726,N_25052,N_25063);
nor UO_727 (O_727,N_29503,N_27205);
xnor UO_728 (O_728,N_29318,N_26336);
and UO_729 (O_729,N_27525,N_25412);
nor UO_730 (O_730,N_26075,N_27765);
nor UO_731 (O_731,N_25991,N_28953);
nor UO_732 (O_732,N_28005,N_26198);
or UO_733 (O_733,N_25659,N_28348);
or UO_734 (O_734,N_26496,N_28569);
or UO_735 (O_735,N_26111,N_27489);
or UO_736 (O_736,N_27377,N_26264);
xor UO_737 (O_737,N_25687,N_28796);
nand UO_738 (O_738,N_27826,N_25886);
and UO_739 (O_739,N_27499,N_26088);
xor UO_740 (O_740,N_27809,N_25994);
or UO_741 (O_741,N_26132,N_29040);
xnor UO_742 (O_742,N_27272,N_26634);
xor UO_743 (O_743,N_29274,N_26508);
or UO_744 (O_744,N_28195,N_28697);
or UO_745 (O_745,N_28727,N_27850);
nand UO_746 (O_746,N_28197,N_25134);
xnor UO_747 (O_747,N_29863,N_29665);
xnor UO_748 (O_748,N_27350,N_28548);
nand UO_749 (O_749,N_29413,N_28945);
xnor UO_750 (O_750,N_27342,N_29498);
xor UO_751 (O_751,N_25514,N_28274);
or UO_752 (O_752,N_25963,N_29672);
nand UO_753 (O_753,N_25369,N_26661);
xnor UO_754 (O_754,N_27114,N_25984);
nor UO_755 (O_755,N_29558,N_27013);
nor UO_756 (O_756,N_26754,N_29684);
nand UO_757 (O_757,N_28641,N_27455);
xnor UO_758 (O_758,N_25913,N_28590);
xor UO_759 (O_759,N_26819,N_26460);
and UO_760 (O_760,N_27308,N_29944);
and UO_761 (O_761,N_27544,N_29346);
xor UO_762 (O_762,N_29160,N_25100);
xor UO_763 (O_763,N_28301,N_26298);
xnor UO_764 (O_764,N_28824,N_28908);
and UO_765 (O_765,N_27947,N_27428);
or UO_766 (O_766,N_25288,N_26536);
xor UO_767 (O_767,N_27171,N_26238);
or UO_768 (O_768,N_27487,N_27624);
nor UO_769 (O_769,N_27337,N_25336);
xor UO_770 (O_770,N_29395,N_29992);
nor UO_771 (O_771,N_26870,N_25820);
nand UO_772 (O_772,N_25706,N_25038);
and UO_773 (O_773,N_27131,N_29398);
and UO_774 (O_774,N_26169,N_25185);
nand UO_775 (O_775,N_26197,N_28766);
nand UO_776 (O_776,N_28091,N_28542);
nor UO_777 (O_777,N_28064,N_26172);
and UO_778 (O_778,N_28044,N_28653);
or UO_779 (O_779,N_28927,N_25390);
nand UO_780 (O_780,N_29078,N_26256);
nand UO_781 (O_781,N_29816,N_26491);
xnor UO_782 (O_782,N_28365,N_25789);
nor UO_783 (O_783,N_26882,N_29788);
nor UO_784 (O_784,N_28801,N_25026);
nand UO_785 (O_785,N_27674,N_28932);
xnor UO_786 (O_786,N_25485,N_27152);
or UO_787 (O_787,N_29978,N_29322);
xnor UO_788 (O_788,N_25686,N_25546);
or UO_789 (O_789,N_26628,N_27585);
nand UO_790 (O_790,N_29836,N_28792);
nor UO_791 (O_791,N_29628,N_27356);
nand UO_792 (O_792,N_27622,N_25772);
nand UO_793 (O_793,N_28157,N_27120);
or UO_794 (O_794,N_27683,N_26347);
or UO_795 (O_795,N_25771,N_26021);
nand UO_796 (O_796,N_28904,N_28019);
and UO_797 (O_797,N_28545,N_29286);
or UO_798 (O_798,N_28679,N_25816);
xor UO_799 (O_799,N_26850,N_29980);
nor UO_800 (O_800,N_29234,N_27936);
or UO_801 (O_801,N_25049,N_27871);
or UO_802 (O_802,N_29682,N_29015);
or UO_803 (O_803,N_25560,N_25650);
or UO_804 (O_804,N_27813,N_29620);
and UO_805 (O_805,N_27676,N_27992);
nor UO_806 (O_806,N_28125,N_28931);
or UO_807 (O_807,N_25267,N_29181);
or UO_808 (O_808,N_27858,N_28769);
nor UO_809 (O_809,N_28089,N_28716);
and UO_810 (O_810,N_25855,N_25797);
nand UO_811 (O_811,N_26278,N_25270);
or UO_812 (O_812,N_29934,N_27548);
xnor UO_813 (O_813,N_29691,N_27841);
xor UO_814 (O_814,N_28919,N_29230);
and UO_815 (O_815,N_27355,N_29033);
xnor UO_816 (O_816,N_27406,N_28225);
nor UO_817 (O_817,N_26403,N_27191);
and UO_818 (O_818,N_26672,N_27851);
nor UO_819 (O_819,N_29486,N_28483);
nand UO_820 (O_820,N_29072,N_26971);
nor UO_821 (O_821,N_26891,N_25192);
or UO_822 (O_822,N_27673,N_29404);
or UO_823 (O_823,N_27045,N_29925);
nor UO_824 (O_824,N_25614,N_29565);
nor UO_825 (O_825,N_25359,N_25670);
nor UO_826 (O_826,N_26175,N_26054);
nor UO_827 (O_827,N_28485,N_25547);
nand UO_828 (O_828,N_28892,N_27922);
xor UO_829 (O_829,N_26183,N_25201);
nand UO_830 (O_830,N_28799,N_29755);
nand UO_831 (O_831,N_27999,N_27710);
nand UO_832 (O_832,N_28496,N_29737);
nor UO_833 (O_833,N_28695,N_25775);
or UO_834 (O_834,N_27122,N_26963);
and UO_835 (O_835,N_26755,N_28224);
xnor UO_836 (O_836,N_29421,N_28117);
nand UO_837 (O_837,N_28255,N_28860);
or UO_838 (O_838,N_29102,N_26765);
xnor UO_839 (O_839,N_26083,N_27755);
nor UO_840 (O_840,N_28933,N_26888);
or UO_841 (O_841,N_27159,N_25089);
xor UO_842 (O_842,N_27280,N_29918);
xnor UO_843 (O_843,N_28460,N_29853);
nor UO_844 (O_844,N_27040,N_27976);
or UO_845 (O_845,N_29443,N_26546);
nor UO_846 (O_846,N_25691,N_29882);
nor UO_847 (O_847,N_29232,N_27049);
nor UO_848 (O_848,N_27057,N_28322);
or UO_849 (O_849,N_25719,N_26486);
nand UO_850 (O_850,N_26537,N_29721);
and UO_851 (O_851,N_28600,N_26410);
nand UO_852 (O_852,N_27256,N_26260);
nand UO_853 (O_853,N_25535,N_27898);
xor UO_854 (O_854,N_29199,N_27047);
or UO_855 (O_855,N_25627,N_29818);
and UO_856 (O_856,N_29971,N_27773);
and UO_857 (O_857,N_27689,N_25031);
or UO_858 (O_858,N_26650,N_26597);
xnor UO_859 (O_859,N_26318,N_28508);
nand UO_860 (O_860,N_28733,N_25538);
nor UO_861 (O_861,N_28409,N_29538);
and UO_862 (O_862,N_26653,N_29878);
nor UO_863 (O_863,N_25423,N_29872);
and UO_864 (O_864,N_28629,N_28331);
nand UO_865 (O_865,N_26507,N_27070);
or UO_866 (O_866,N_26421,N_29004);
or UO_867 (O_867,N_25604,N_26164);
nor UO_868 (O_868,N_29767,N_26812);
nand UO_869 (O_869,N_29210,N_28004);
and UO_870 (O_870,N_29271,N_25047);
xnor UO_871 (O_871,N_27417,N_25878);
xnor UO_872 (O_872,N_27865,N_29314);
nand UO_873 (O_873,N_29716,N_25896);
nor UO_874 (O_874,N_25697,N_25065);
and UO_875 (O_875,N_25582,N_25311);
xor UO_876 (O_876,N_28222,N_29054);
or UO_877 (O_877,N_26086,N_27637);
nand UO_878 (O_878,N_26716,N_29309);
or UO_879 (O_879,N_26135,N_28638);
xnor UO_880 (O_880,N_26511,N_25933);
or UO_881 (O_881,N_26949,N_29391);
xor UO_882 (O_882,N_26470,N_27380);
xnor UO_883 (O_883,N_29348,N_29379);
and UO_884 (O_884,N_26655,N_29700);
or UO_885 (O_885,N_27892,N_28861);
xor UO_886 (O_886,N_25118,N_27150);
nand UO_887 (O_887,N_26823,N_26320);
xnor UO_888 (O_888,N_29995,N_26317);
and UO_889 (O_889,N_26463,N_26815);
nand UO_890 (O_890,N_25342,N_27894);
and UO_891 (O_891,N_26524,N_29766);
or UO_892 (O_892,N_25167,N_25371);
nand UO_893 (O_893,N_25785,N_26759);
xor UO_894 (O_894,N_26346,N_28737);
and UO_895 (O_895,N_29090,N_29561);
nor UO_896 (O_896,N_26268,N_25517);
nand UO_897 (O_897,N_26031,N_28655);
xnor UO_898 (O_898,N_25280,N_28048);
xor UO_899 (O_899,N_28293,N_26828);
or UO_900 (O_900,N_29683,N_28630);
xor UO_901 (O_901,N_26852,N_26324);
nand UO_902 (O_902,N_26953,N_25051);
and UO_903 (O_903,N_28100,N_27662);
nor UO_904 (O_904,N_29487,N_27395);
nand UO_905 (O_905,N_29368,N_25032);
xor UO_906 (O_906,N_28261,N_25782);
nor UO_907 (O_907,N_25264,N_25879);
xor UO_908 (O_908,N_25447,N_28315);
nor UO_909 (O_909,N_26924,N_25320);
or UO_910 (O_910,N_29377,N_25930);
nor UO_911 (O_911,N_27753,N_27316);
nand UO_912 (O_912,N_29480,N_25575);
nor UO_913 (O_913,N_29931,N_26730);
nor UO_914 (O_914,N_29785,N_25273);
nor UO_915 (O_915,N_26367,N_25142);
xnor UO_916 (O_916,N_26528,N_25163);
nor UO_917 (O_917,N_25189,N_25519);
or UO_918 (O_918,N_25080,N_25951);
nor UO_919 (O_919,N_26040,N_26173);
or UO_920 (O_920,N_26774,N_26905);
nor UO_921 (O_921,N_28120,N_29588);
xor UO_922 (O_922,N_29027,N_26777);
or UO_923 (O_923,N_29996,N_29744);
nor UO_924 (O_924,N_28518,N_28434);
and UO_925 (O_925,N_26252,N_29176);
or UO_926 (O_926,N_25959,N_26982);
and UO_927 (O_927,N_26045,N_27684);
xor UO_928 (O_928,N_25707,N_27323);
nor UO_929 (O_929,N_25757,N_25054);
and UO_930 (O_930,N_29796,N_26640);
or UO_931 (O_931,N_25350,N_25354);
nor UO_932 (O_932,N_26258,N_25833);
nor UO_933 (O_933,N_27539,N_28343);
xnor UO_934 (O_934,N_26442,N_28840);
nand UO_935 (O_935,N_28970,N_27210);
and UO_936 (O_936,N_29532,N_29617);
and UO_937 (O_937,N_26226,N_26778);
or UO_938 (O_938,N_26026,N_26016);
xor UO_939 (O_939,N_28808,N_25463);
and UO_940 (O_940,N_28228,N_28648);
or UO_941 (O_941,N_27135,N_29625);
nand UO_942 (O_942,N_26478,N_27516);
nor UO_943 (O_943,N_28467,N_29052);
nor UO_944 (O_944,N_25316,N_27776);
or UO_945 (O_945,N_29337,N_29957);
and UO_946 (O_946,N_26241,N_27361);
xnor UO_947 (O_947,N_28998,N_28615);
and UO_948 (O_948,N_27860,N_29010);
nor UO_949 (O_949,N_26301,N_25082);
and UO_950 (O_950,N_28351,N_25079);
xor UO_951 (O_951,N_27164,N_28800);
nand UO_952 (O_952,N_29342,N_28032);
xor UO_953 (O_953,N_29539,N_28196);
or UO_954 (O_954,N_26768,N_26456);
nor UO_955 (O_955,N_26692,N_27496);
nand UO_956 (O_956,N_25502,N_28367);
nor UO_957 (O_957,N_25718,N_27044);
or UO_958 (O_958,N_26262,N_29666);
or UO_959 (O_959,N_26802,N_29776);
or UO_960 (O_960,N_29756,N_28665);
nand UO_961 (O_961,N_25870,N_25769);
nand UO_962 (O_962,N_28965,N_28691);
nor UO_963 (O_963,N_28191,N_26610);
nor UO_964 (O_964,N_29724,N_29250);
xor UO_965 (O_965,N_29655,N_27022);
xnor UO_966 (O_966,N_27954,N_25916);
or UO_967 (O_967,N_28756,N_26439);
nand UO_968 (O_968,N_26339,N_26554);
or UO_969 (O_969,N_27833,N_27520);
nand UO_970 (O_970,N_26465,N_26895);
nor UO_971 (O_971,N_26885,N_26082);
and UO_972 (O_972,N_26287,N_28928);
nand UO_973 (O_973,N_29589,N_28685);
xor UO_974 (O_974,N_26557,N_27160);
xnor UO_975 (O_975,N_27914,N_25850);
or UO_976 (O_976,N_27650,N_27462);
nor UO_977 (O_977,N_27629,N_25703);
xnor UO_978 (O_978,N_27058,N_27224);
xor UO_979 (O_979,N_26017,N_28775);
nor UO_980 (O_980,N_26530,N_25418);
nor UO_981 (O_981,N_28551,N_26856);
nand UO_982 (O_982,N_25045,N_28558);
and UO_983 (O_983,N_26162,N_27632);
or UO_984 (O_984,N_26540,N_29110);
xnor UO_985 (O_985,N_25460,N_29432);
xnor UO_986 (O_986,N_29825,N_26615);
or UO_987 (O_987,N_27046,N_27139);
xor UO_988 (O_988,N_26251,N_25207);
or UO_989 (O_989,N_25471,N_29020);
nor UO_990 (O_990,N_25813,N_25450);
and UO_991 (O_991,N_26380,N_25980);
xnor UO_992 (O_992,N_25966,N_29330);
and UO_993 (O_993,N_28903,N_26281);
and UO_994 (O_994,N_29595,N_27739);
or UO_995 (O_995,N_25598,N_25770);
nor UO_996 (O_996,N_27577,N_25146);
nand UO_997 (O_997,N_28041,N_26826);
and UO_998 (O_998,N_29153,N_27090);
xor UO_999 (O_999,N_25122,N_28725);
nor UO_1000 (O_1000,N_27384,N_29278);
or UO_1001 (O_1001,N_29981,N_28349);
xor UO_1002 (O_1002,N_26654,N_26419);
nor UO_1003 (O_1003,N_28220,N_29373);
nand UO_1004 (O_1004,N_25405,N_26733);
or UO_1005 (O_1005,N_26453,N_27106);
xor UO_1006 (O_1006,N_29458,N_29221);
xnor UO_1007 (O_1007,N_25634,N_27270);
and UO_1008 (O_1008,N_27678,N_26770);
or UO_1009 (O_1009,N_27616,N_27821);
or UO_1010 (O_1010,N_28018,N_26266);
or UO_1011 (O_1011,N_25783,N_26806);
nand UO_1012 (O_1012,N_26458,N_29341);
and UO_1013 (O_1013,N_28181,N_25279);
nor UO_1014 (O_1014,N_26097,N_26506);
xnor UO_1015 (O_1015,N_27996,N_28914);
xnor UO_1016 (O_1016,N_25774,N_27351);
or UO_1017 (O_1017,N_29763,N_29920);
xnor UO_1018 (O_1018,N_28930,N_26930);
and UO_1019 (O_1019,N_25688,N_29104);
and UO_1020 (O_1020,N_28539,N_26309);
xnor UO_1021 (O_1021,N_28992,N_27424);
nor UO_1022 (O_1022,N_29497,N_29312);
xor UO_1023 (O_1023,N_28742,N_26691);
or UO_1024 (O_1024,N_26096,N_29566);
nor UO_1025 (O_1025,N_26200,N_29364);
nor UO_1026 (O_1026,N_25700,N_26512);
nand UO_1027 (O_1027,N_25784,N_26345);
and UO_1028 (O_1028,N_25819,N_27028);
or UO_1029 (O_1029,N_25730,N_28525);
and UO_1030 (O_1030,N_25805,N_29607);
or UO_1031 (O_1031,N_26423,N_27032);
and UO_1032 (O_1032,N_25607,N_25530);
nand UO_1033 (O_1033,N_29370,N_28455);
or UO_1034 (O_1034,N_25801,N_28250);
or UO_1035 (O_1035,N_27533,N_27835);
and UO_1036 (O_1036,N_27108,N_25138);
xnor UO_1037 (O_1037,N_26166,N_25906);
nand UO_1038 (O_1038,N_29610,N_25190);
nand UO_1039 (O_1039,N_29646,N_29940);
or UO_1040 (O_1040,N_27074,N_28461);
nor UO_1041 (O_1041,N_27430,N_26104);
and UO_1042 (O_1042,N_28339,N_28868);
nand UO_1043 (O_1043,N_28123,N_27401);
xor UO_1044 (O_1044,N_26428,N_25979);
xnor UO_1045 (O_1045,N_25968,N_28583);
nor UO_1046 (O_1046,N_25778,N_28169);
nand UO_1047 (O_1047,N_26398,N_29490);
or UO_1048 (O_1048,N_29298,N_25714);
and UO_1049 (O_1049,N_27228,N_25531);
and UO_1050 (O_1050,N_28598,N_27977);
or UO_1051 (O_1051,N_25128,N_26881);
or UO_1052 (O_1052,N_26928,N_27408);
and UO_1053 (O_1053,N_25507,N_26438);
and UO_1054 (O_1054,N_27569,N_27994);
nor UO_1055 (O_1055,N_27754,N_25012);
nand UO_1056 (O_1056,N_25851,N_28740);
nand UO_1057 (O_1057,N_26797,N_26291);
xnor UO_1058 (O_1058,N_29752,N_28218);
nand UO_1059 (O_1059,N_29382,N_29009);
nand UO_1060 (O_1060,N_27277,N_26501);
nand UO_1061 (O_1061,N_27452,N_25019);
nor UO_1062 (O_1062,N_26113,N_27762);
nor UO_1063 (O_1063,N_26385,N_27595);
xnor UO_1064 (O_1064,N_27158,N_28764);
nand UO_1065 (O_1065,N_29622,N_28803);
nor UO_1066 (O_1066,N_26070,N_29222);
or UO_1067 (O_1067,N_29795,N_27240);
and UO_1068 (O_1068,N_28848,N_29706);
nor UO_1069 (O_1069,N_28547,N_28474);
and UO_1070 (O_1070,N_27237,N_26038);
nor UO_1071 (O_1071,N_29132,N_26970);
xor UO_1072 (O_1072,N_27354,N_28721);
nor UO_1073 (O_1073,N_26849,N_27633);
nor UO_1074 (O_1074,N_25357,N_27706);
xor UO_1075 (O_1075,N_27002,N_29673);
nor UO_1076 (O_1076,N_28978,N_29324);
nand UO_1077 (O_1077,N_27742,N_26579);
or UO_1078 (O_1078,N_25491,N_28122);
nand UO_1079 (O_1079,N_28898,N_28264);
and UO_1080 (O_1080,N_27908,N_25240);
xnor UO_1081 (O_1081,N_27345,N_27691);
nand UO_1082 (O_1082,N_28444,N_26959);
xor UO_1083 (O_1083,N_26997,N_26564);
nand UO_1084 (O_1084,N_27519,N_27052);
nand UO_1085 (O_1085,N_25364,N_27083);
nor UO_1086 (O_1086,N_28329,N_27867);
and UO_1087 (O_1087,N_29598,N_28333);
xnor UO_1088 (O_1088,N_28254,N_29578);
and UO_1089 (O_1089,N_25339,N_27078);
nand UO_1090 (O_1090,N_25081,N_28292);
and UO_1091 (O_1091,N_28130,N_27998);
nand UO_1092 (O_1092,N_28033,N_26313);
nand UO_1093 (O_1093,N_29760,N_28661);
and UO_1094 (O_1094,N_26065,N_25745);
or UO_1095 (O_1095,N_27115,N_27521);
xor UO_1096 (O_1096,N_25571,N_27094);
and UO_1097 (O_1097,N_25465,N_29786);
or UO_1098 (O_1098,N_26723,N_26485);
and UO_1099 (O_1099,N_26838,N_27798);
nor UO_1100 (O_1100,N_25324,N_26255);
nand UO_1101 (O_1101,N_28305,N_28469);
xnor UO_1102 (O_1102,N_25410,N_25011);
or UO_1103 (O_1103,N_25055,N_26824);
nor UO_1104 (O_1104,N_29514,N_27144);
nor UO_1105 (O_1105,N_26601,N_27071);
nor UO_1106 (O_1106,N_27716,N_26283);
xor UO_1107 (O_1107,N_29758,N_25508);
nand UO_1108 (O_1108,N_29381,N_29426);
nor UO_1109 (O_1109,N_26835,N_26208);
or UO_1110 (O_1110,N_26981,N_28058);
and UO_1111 (O_1111,N_29284,N_26789);
and UO_1112 (O_1112,N_28215,N_27837);
nand UO_1113 (O_1113,N_28957,N_25147);
or UO_1114 (O_1114,N_25856,N_29774);
xnor UO_1115 (O_1115,N_27903,N_25233);
nand UO_1116 (O_1116,N_27145,N_27467);
and UO_1117 (O_1117,N_27232,N_28429);
or UO_1118 (O_1118,N_26192,N_28337);
and UO_1119 (O_1119,N_26267,N_25891);
nand UO_1120 (O_1120,N_25758,N_28778);
nand UO_1121 (O_1121,N_25854,N_29560);
or UO_1122 (O_1122,N_25990,N_29567);
and UO_1123 (O_1123,N_25133,N_25370);
and UO_1124 (O_1124,N_25524,N_26521);
or UO_1125 (O_1125,N_27069,N_29734);
nor UO_1126 (O_1126,N_27969,N_29698);
nor UO_1127 (O_1127,N_25857,N_26664);
xor UO_1128 (O_1128,N_29095,N_29546);
nand UO_1129 (O_1129,N_27426,N_27806);
xnor UO_1130 (O_1130,N_25890,N_25964);
nor UO_1131 (O_1131,N_26932,N_28577);
nor UO_1132 (O_1132,N_29953,N_28006);
and UO_1133 (O_1133,N_28372,N_25346);
nand UO_1134 (O_1134,N_28947,N_28345);
xnor UO_1135 (O_1135,N_28059,N_28172);
nor UO_1136 (O_1136,N_26303,N_28057);
nor UO_1137 (O_1137,N_27877,N_26223);
nand UO_1138 (O_1138,N_26753,N_25668);
or UO_1139 (O_1139,N_26594,N_26340);
nor UO_1140 (O_1140,N_26941,N_29500);
xnor UO_1141 (O_1141,N_25473,N_25407);
nor UO_1142 (O_1142,N_27705,N_28183);
xnor UO_1143 (O_1143,N_29491,N_25672);
nor UO_1144 (O_1144,N_28774,N_25931);
or UO_1145 (O_1145,N_27247,N_27752);
nand UO_1146 (O_1146,N_28503,N_27340);
or UO_1147 (O_1147,N_27663,N_28592);
or UO_1148 (O_1148,N_28573,N_28880);
nand UO_1149 (O_1149,N_25981,N_27041);
nor UO_1150 (O_1150,N_25631,N_27825);
nor UO_1151 (O_1151,N_29641,N_27788);
and UO_1152 (O_1152,N_25564,N_28871);
or UO_1153 (O_1153,N_28124,N_27905);
nand UO_1154 (O_1154,N_27076,N_26141);
and UO_1155 (O_1155,N_25462,N_28366);
and UO_1156 (O_1156,N_25198,N_27230);
and UO_1157 (O_1157,N_26907,N_27005);
nor UO_1158 (O_1158,N_29575,N_28489);
nand UO_1159 (O_1159,N_25860,N_26374);
nand UO_1160 (O_1160,N_29327,N_25777);
and UO_1161 (O_1161,N_26235,N_28847);
or UO_1162 (O_1162,N_26068,N_29912);
nand UO_1163 (O_1163,N_27889,N_27291);
and UO_1164 (O_1164,N_28813,N_29867);
nor UO_1165 (O_1165,N_26872,N_27051);
or UO_1166 (O_1166,N_29360,N_27719);
nand UO_1167 (O_1167,N_26055,N_29975);
nand UO_1168 (O_1168,N_25944,N_28083);
nand UO_1169 (O_1169,N_28296,N_25351);
nor UO_1170 (O_1170,N_26314,N_29591);
nand UO_1171 (O_1171,N_29150,N_25183);
or UO_1172 (O_1172,N_26237,N_25581);
xor UO_1173 (O_1173,N_27276,N_27744);
or UO_1174 (O_1174,N_27381,N_26473);
xor UO_1175 (O_1175,N_28428,N_25326);
nor UO_1176 (O_1176,N_29824,N_26037);
or UO_1177 (O_1177,N_27983,N_26645);
nand UO_1178 (O_1178,N_25208,N_28650);
xor UO_1179 (O_1179,N_29639,N_25802);
xor UO_1180 (O_1180,N_27301,N_25363);
xor UO_1181 (O_1181,N_25952,N_29457);
xor UO_1182 (O_1182,N_27290,N_29508);
or UO_1183 (O_1183,N_26827,N_28676);
and UO_1184 (O_1184,N_26302,N_25143);
or UO_1185 (O_1185,N_27801,N_25286);
nand UO_1186 (O_1186,N_29937,N_26693);
nor UO_1187 (O_1187,N_26269,N_28877);
nor UO_1188 (O_1188,N_28401,N_29385);
nor UO_1189 (O_1189,N_29159,N_26187);
xor UO_1190 (O_1190,N_25414,N_28045);
nand UO_1191 (O_1191,N_25338,N_26843);
nand UO_1192 (O_1192,N_29640,N_25641);
nand UO_1193 (O_1193,N_26431,N_26076);
nand UO_1194 (O_1194,N_28594,N_29451);
and UO_1195 (O_1195,N_28690,N_25516);
or UO_1196 (O_1196,N_27644,N_28770);
and UO_1197 (O_1197,N_28283,N_27376);
or UO_1198 (O_1198,N_28062,N_29729);
or UO_1199 (O_1199,N_27370,N_27362);
and UO_1200 (O_1200,N_25825,N_29175);
xnor UO_1201 (O_1201,N_25041,N_28532);
or UO_1202 (O_1202,N_29720,N_28963);
nand UO_1203 (O_1203,N_28096,N_27974);
nand UO_1204 (O_1204,N_26426,N_26605);
xor UO_1205 (O_1205,N_29315,N_29799);
or UO_1206 (O_1206,N_27846,N_29997);
and UO_1207 (O_1207,N_29187,N_28223);
xnor UO_1208 (O_1208,N_27993,N_27274);
and UO_1209 (O_1209,N_27483,N_29121);
xor UO_1210 (O_1210,N_27743,N_29986);
or UO_1211 (O_1211,N_29765,N_27146);
and UO_1212 (O_1212,N_28724,N_25046);
nor UO_1213 (O_1213,N_28131,N_25253);
or UO_1214 (O_1214,N_25786,N_29151);
nor UO_1215 (O_1215,N_25744,N_28554);
nand UO_1216 (O_1216,N_29077,N_29549);
nor UO_1217 (O_1217,N_27643,N_27140);
nand UO_1218 (O_1218,N_29235,N_25156);
or UO_1219 (O_1219,N_28424,N_29518);
and UO_1220 (O_1220,N_26787,N_28212);
xnor UO_1221 (O_1221,N_28167,N_27259);
xnor UO_1222 (O_1222,N_27945,N_28588);
xnor UO_1223 (O_1223,N_26454,N_27931);
or UO_1224 (O_1224,N_29062,N_25087);
nand UO_1225 (O_1225,N_29108,N_26967);
nand UO_1226 (O_1226,N_28323,N_26735);
and UO_1227 (O_1227,N_25572,N_28711);
or UO_1228 (O_1228,N_29207,N_25001);
xor UO_1229 (O_1229,N_29280,N_25226);
xnor UO_1230 (O_1230,N_27518,N_29310);
nand UO_1231 (O_1231,N_28787,N_25568);
or UO_1232 (O_1232,N_27365,N_29138);
xor UO_1233 (O_1233,N_28680,N_26804);
and UO_1234 (O_1234,N_27540,N_25549);
or UO_1235 (O_1235,N_28442,N_28705);
or UO_1236 (O_1236,N_26822,N_26662);
xor UO_1237 (O_1237,N_25008,N_27989);
nor UO_1238 (O_1238,N_28314,N_26978);
nor UO_1239 (O_1239,N_26493,N_28838);
or UO_1240 (O_1240,N_25611,N_26519);
nor UO_1241 (O_1241,N_28603,N_28783);
xor UO_1242 (O_1242,N_26725,N_25736);
xor UO_1243 (O_1243,N_26234,N_29475);
and UO_1244 (O_1244,N_26466,N_29257);
and UO_1245 (O_1245,N_28593,N_28277);
or UO_1246 (O_1246,N_25898,N_25729);
or UO_1247 (O_1247,N_28610,N_26575);
nand UO_1248 (O_1248,N_25425,N_25088);
nor UO_1249 (O_1249,N_29416,N_29983);
xor UO_1250 (O_1250,N_29801,N_25788);
xnor UO_1251 (O_1251,N_29547,N_29039);
nor UO_1252 (O_1252,N_26411,N_27433);
xnor UO_1253 (O_1253,N_28571,N_26352);
xor UO_1254 (O_1254,N_25977,N_27383);
and UO_1255 (O_1255,N_27882,N_26893);
and UO_1256 (O_1256,N_25618,N_27951);
and UO_1257 (O_1257,N_26520,N_25954);
or UO_1258 (O_1258,N_28102,N_29372);
or UO_1259 (O_1259,N_27010,N_25975);
xnor UO_1260 (O_1260,N_29410,N_29119);
nand UO_1261 (O_1261,N_26180,N_27598);
or UO_1262 (O_1262,N_25583,N_29001);
and UO_1263 (O_1263,N_28617,N_26353);
xnor UO_1264 (O_1264,N_27060,N_28298);
nor UO_1265 (O_1265,N_26977,N_28530);
xor UO_1266 (O_1266,N_25302,N_29349);
nand UO_1267 (O_1267,N_28757,N_26190);
xor UO_1268 (O_1268,N_26652,N_28105);
nand UO_1269 (O_1269,N_26373,N_26985);
nor UO_1270 (O_1270,N_25221,N_29456);
and UO_1271 (O_1271,N_28155,N_26101);
nand UO_1272 (O_1272,N_26814,N_27952);
nor UO_1273 (O_1273,N_27328,N_25174);
nand UO_1274 (O_1274,N_28235,N_27526);
xnor UO_1275 (O_1275,N_25912,N_28907);
nand UO_1276 (O_1276,N_25561,N_29173);
and UO_1277 (O_1277,N_27242,N_29231);
xor UO_1278 (O_1278,N_25812,N_25803);
nand UO_1279 (O_1279,N_25940,N_26906);
or UO_1280 (O_1280,N_28678,N_26020);
and UO_1281 (O_1281,N_27311,N_25643);
xnor UO_1282 (O_1282,N_28207,N_27604);
and UO_1283 (O_1283,N_25764,N_26476);
xor UO_1284 (O_1284,N_29225,N_25441);
xnor UO_1285 (O_1285,N_29730,N_25993);
xor UO_1286 (O_1286,N_28126,N_26286);
nor UO_1287 (O_1287,N_27968,N_29502);
nand UO_1288 (O_1288,N_28728,N_25800);
nand UO_1289 (O_1289,N_25717,N_28635);
or UO_1290 (O_1290,N_28982,N_29060);
nand UO_1291 (O_1291,N_25488,N_27567);
nand UO_1292 (O_1292,N_28996,N_28022);
or UO_1293 (O_1293,N_29462,N_29440);
xnor UO_1294 (O_1294,N_26123,N_28162);
xor UO_1295 (O_1295,N_29751,N_25793);
and UO_1296 (O_1296,N_25696,N_29969);
xor UO_1297 (O_1297,N_29648,N_26687);
and UO_1298 (O_1298,N_28565,N_29861);
and UO_1299 (O_1299,N_27784,N_26271);
xnor UO_1300 (O_1300,N_25454,N_28741);
and UO_1301 (O_1301,N_26713,N_27303);
xor UO_1302 (O_1302,N_29433,N_27018);
nor UO_1303 (O_1303,N_26012,N_28890);
nand UO_1304 (O_1304,N_28811,N_25303);
xor UO_1305 (O_1305,N_26159,N_28702);
xor UO_1306 (O_1306,N_28956,N_25852);
nor UO_1307 (O_1307,N_27404,N_25132);
nor UO_1308 (O_1308,N_27640,N_28007);
and UO_1309 (O_1309,N_28710,N_29079);
nand UO_1310 (O_1310,N_25866,N_25695);
or UO_1311 (O_1311,N_25307,N_25605);
or UO_1312 (O_1312,N_26740,N_26751);
or UO_1313 (O_1313,N_29263,N_28637);
and UO_1314 (O_1314,N_26668,N_25121);
nor UO_1315 (O_1315,N_29254,N_25166);
nand UO_1316 (O_1316,N_27891,N_29664);
and UO_1317 (O_1317,N_29710,N_25648);
nand UO_1318 (O_1318,N_27596,N_28694);
nand UO_1319 (O_1319,N_25432,N_27050);
xor UO_1320 (O_1320,N_27004,N_28784);
xor UO_1321 (O_1321,N_25271,N_28436);
and UO_1322 (O_1322,N_26666,N_27528);
xor UO_1323 (O_1323,N_27399,N_29174);
nand UO_1324 (O_1324,N_25365,N_29834);
nor UO_1325 (O_1325,N_26227,N_26370);
and UO_1326 (O_1326,N_28677,N_29504);
or UO_1327 (O_1327,N_25894,N_25715);
nand UO_1328 (O_1328,N_25748,N_27366);
or UO_1329 (O_1329,N_26253,N_26795);
nand UO_1330 (O_1330,N_25529,N_29329);
or UO_1331 (O_1331,N_25899,N_28318);
nand UO_1332 (O_1332,N_26808,N_29857);
nand UO_1333 (O_1333,N_27542,N_26922);
and UO_1334 (O_1334,N_26782,N_28465);
and UO_1335 (O_1335,N_25978,N_27273);
or UO_1336 (O_1336,N_29215,N_28659);
nor UO_1337 (O_1337,N_29830,N_29554);
or UO_1338 (O_1338,N_26002,N_25211);
nand UO_1339 (O_1339,N_26325,N_25442);
xnor UO_1340 (O_1340,N_26983,N_25193);
nand UO_1341 (O_1341,N_27756,N_26899);
and UO_1342 (O_1342,N_28043,N_28946);
nor UO_1343 (O_1343,N_29101,N_26591);
or UO_1344 (O_1344,N_25313,N_29224);
nand UO_1345 (O_1345,N_25608,N_29843);
nor UO_1346 (O_1346,N_27635,N_26053);
xor UO_1347 (O_1347,N_27403,N_28823);
nand UO_1348 (O_1348,N_28762,N_26689);
xor UO_1349 (O_1349,N_29873,N_29903);
and UO_1350 (O_1350,N_28484,N_29299);
and UO_1351 (O_1351,N_27353,N_25711);
and UO_1352 (O_1352,N_29478,N_26934);
nand UO_1353 (O_1353,N_28730,N_26219);
and UO_1354 (O_1354,N_26943,N_28422);
nor UO_1355 (O_1355,N_25616,N_29688);
nor UO_1356 (O_1356,N_25176,N_29967);
or UO_1357 (O_1357,N_25392,N_28994);
or UO_1358 (O_1358,N_29103,N_26444);
nand UO_1359 (O_1359,N_28505,N_29326);
xor UO_1360 (O_1360,N_27870,N_26305);
or UO_1361 (O_1361,N_26669,N_26697);
nand UO_1362 (O_1362,N_26050,N_25479);
nand UO_1363 (O_1363,N_27446,N_27991);
or UO_1364 (O_1364,N_28942,N_28669);
nand UO_1365 (O_1365,N_28543,N_28300);
xnor UO_1366 (O_1366,N_27868,N_27924);
or UO_1367 (O_1367,N_25083,N_25005);
or UO_1368 (O_1368,N_28791,N_25252);
nor UO_1369 (O_1369,N_29056,N_27116);
xor UO_1370 (O_1370,N_26362,N_29059);
nand UO_1371 (O_1371,N_25637,N_26903);
and UO_1372 (O_1372,N_25385,N_26734);
and UO_1373 (O_1373,N_26181,N_29331);
or UO_1374 (O_1374,N_28605,N_26525);
nand UO_1375 (O_1375,N_26951,N_25374);
and UO_1376 (O_1376,N_25056,N_28815);
or UO_1377 (O_1377,N_25437,N_27300);
or UO_1378 (O_1378,N_28185,N_25996);
or UO_1379 (O_1379,N_28864,N_25234);
xnor UO_1380 (O_1380,N_25655,N_29495);
xor UO_1381 (O_1381,N_28350,N_27407);
or UO_1382 (O_1382,N_26727,N_25875);
xor UO_1383 (O_1383,N_27593,N_26756);
nand UO_1384 (O_1384,N_25164,N_28390);
or UO_1385 (O_1385,N_28623,N_26674);
xnor UO_1386 (O_1386,N_27822,N_26686);
and UO_1387 (O_1387,N_26014,N_29035);
xnor UO_1388 (O_1388,N_28606,N_28520);
xnor UO_1389 (O_1389,N_27397,N_28698);
or UO_1390 (O_1390,N_28391,N_29529);
nor UO_1391 (O_1391,N_28580,N_27748);
and UO_1392 (O_1392,N_27008,N_25318);
nor UO_1393 (O_1393,N_29245,N_28361);
and UO_1394 (O_1394,N_29723,N_29782);
and UO_1395 (O_1395,N_25402,N_26280);
xnor UO_1396 (O_1396,N_26535,N_26706);
nor UO_1397 (O_1397,N_25728,N_26549);
nor UO_1398 (O_1398,N_27582,N_29592);
xor UO_1399 (O_1399,N_25742,N_29152);
and UO_1400 (O_1400,N_26894,N_28544);
xor UO_1401 (O_1401,N_27129,N_28829);
or UO_1402 (O_1402,N_25386,N_28399);
or UO_1403 (O_1403,N_25970,N_25098);
and UO_1404 (O_1404,N_27126,N_28009);
and UO_1405 (O_1405,N_28913,N_26679);
xor UO_1406 (O_1406,N_27439,N_29609);
nand UO_1407 (O_1407,N_27431,N_26769);
xnor UO_1408 (O_1408,N_26273,N_28201);
or UO_1409 (O_1409,N_28341,N_28865);
and UO_1410 (O_1410,N_29454,N_27712);
and UO_1411 (O_1411,N_25347,N_25639);
xnor UO_1412 (O_1412,N_29290,N_29296);
nand UO_1413 (O_1413,N_27915,N_29656);
nand UO_1414 (O_1414,N_29778,N_27163);
xnor UO_1415 (O_1415,N_29472,N_29540);
xor UO_1416 (O_1416,N_25685,N_28095);
xor UO_1417 (O_1417,N_26875,N_27405);
nand UO_1418 (O_1418,N_26984,N_26383);
nand UO_1419 (O_1419,N_28736,N_25553);
and UO_1420 (O_1420,N_28674,N_27597);
nor UO_1421 (O_1421,N_29653,N_29645);
or UO_1422 (O_1422,N_28290,N_27358);
or UO_1423 (O_1423,N_27461,N_26142);
xor UO_1424 (O_1424,N_27941,N_26957);
nor UO_1425 (O_1425,N_27339,N_25573);
or UO_1426 (O_1426,N_27711,N_26010);
nand UO_1427 (O_1427,N_28137,N_28211);
and UO_1428 (O_1428,N_25620,N_27730);
and UO_1429 (O_1429,N_28662,N_29388);
and UO_1430 (O_1430,N_29845,N_29537);
or UO_1431 (O_1431,N_26039,N_29633);
nand UO_1432 (O_1432,N_28387,N_26935);
xnor UO_1433 (O_1433,N_27950,N_28232);
or UO_1434 (O_1434,N_29686,N_28609);
and UO_1435 (O_1435,N_25710,N_27157);
nor UO_1436 (O_1436,N_26726,N_27100);
or UO_1437 (O_1437,N_25982,N_27934);
or UO_1438 (O_1438,N_29453,N_25923);
nand UO_1439 (O_1439,N_29929,N_25839);
xor UO_1440 (O_1440,N_25558,N_28262);
and UO_1441 (O_1441,N_25590,N_27075);
and UO_1442 (O_1442,N_29663,N_28014);
or UO_1443 (O_1443,N_27245,N_28969);
or UO_1444 (O_1444,N_29012,N_25595);
nor UO_1445 (O_1445,N_26534,N_27469);
nor UO_1446 (O_1446,N_27294,N_29045);
nor UO_1447 (O_1447,N_27627,N_28999);
nor UO_1448 (O_1448,N_29182,N_27458);
nor UO_1449 (O_1449,N_27216,N_29198);
xnor UO_1450 (O_1450,N_26569,N_28233);
and UO_1451 (O_1451,N_26883,N_28330);
nand UO_1452 (O_1452,N_25254,N_25640);
and UO_1453 (O_1453,N_26196,N_29311);
nor UO_1454 (O_1454,N_25958,N_28747);
xnor UO_1455 (O_1455,N_25762,N_26955);
xor UO_1456 (O_1456,N_28561,N_28327);
nor UO_1457 (O_1457,N_26489,N_29761);
xnor UO_1458 (O_1458,N_29722,N_26436);
xnor UO_1459 (O_1459,N_26630,N_26612);
nor UO_1460 (O_1460,N_25863,N_27333);
or UO_1461 (O_1461,N_25272,N_29533);
nand UO_1462 (O_1462,N_28990,N_25310);
nand UO_1463 (O_1463,N_28087,N_28481);
or UO_1464 (O_1464,N_25251,N_26622);
xnor UO_1465 (O_1465,N_28821,N_27234);
and UO_1466 (O_1466,N_28352,N_29303);
and UO_1467 (O_1467,N_28309,N_28127);
nor UO_1468 (O_1468,N_25946,N_27059);
nor UO_1469 (O_1469,N_26295,N_26213);
nor UO_1470 (O_1470,N_27410,N_25421);
nand UO_1471 (O_1471,N_26163,N_26072);
and UO_1472 (O_1472,N_25305,N_27194);
xnor UO_1473 (O_1473,N_26332,N_25907);
or UO_1474 (O_1474,N_26590,N_25908);
and UO_1475 (O_1475,N_28536,N_25677);
or UO_1476 (O_1476,N_25027,N_28681);
nand UO_1477 (O_1477,N_26249,N_29041);
xnor UO_1478 (O_1478,N_27422,N_29239);
xnor UO_1479 (O_1479,N_26861,N_25476);
nand UO_1480 (O_1480,N_26758,N_29378);
nand UO_1481 (O_1481,N_27479,N_26598);
xnor UO_1482 (O_1482,N_27607,N_28410);
xnor UO_1483 (O_1483,N_29526,N_29065);
nor UO_1484 (O_1484,N_29961,N_26494);
or UO_1485 (O_1485,N_26533,N_29272);
or UO_1486 (O_1486,N_29124,N_26825);
or UO_1487 (O_1487,N_29135,N_28302);
or UO_1488 (O_1488,N_27811,N_27307);
nand UO_1489 (O_1489,N_25150,N_29743);
nand UO_1490 (O_1490,N_25817,N_29246);
or UO_1491 (O_1491,N_27670,N_27475);
nor UO_1492 (O_1492,N_29613,N_27267);
or UO_1493 (O_1493,N_28202,N_28585);
nand UO_1494 (O_1494,N_29044,N_27713);
xor UO_1495 (O_1495,N_28206,N_27504);
and UO_1496 (O_1496,N_28531,N_27495);
and UO_1497 (O_1497,N_27389,N_25495);
xnor UO_1498 (O_1498,N_25911,N_26030);
nor UO_1499 (O_1499,N_26224,N_26341);
nand UO_1500 (O_1500,N_26310,N_27799);
or UO_1501 (O_1501,N_25224,N_26592);
and UO_1502 (O_1502,N_27155,N_27697);
xnor UO_1503 (O_1503,N_26749,N_26722);
xor UO_1504 (O_1504,N_25111,N_26168);
or UO_1505 (O_1505,N_28369,N_27239);
and UO_1506 (O_1506,N_27862,N_28901);
nand UO_1507 (O_1507,N_29911,N_28937);
xnor UO_1508 (O_1508,N_29678,N_25868);
nand UO_1509 (O_1509,N_26377,N_29434);
nand UO_1510 (O_1510,N_28836,N_25440);
and UO_1511 (O_1511,N_29118,N_27775);
or UO_1512 (O_1512,N_26887,N_25062);
xnor UO_1513 (O_1513,N_27306,N_27136);
or UO_1514 (O_1514,N_25843,N_25084);
xor UO_1515 (O_1515,N_27183,N_29218);
nor UO_1516 (O_1516,N_28922,N_26811);
or UO_1517 (O_1517,N_28818,N_28394);
nand UO_1518 (O_1518,N_27501,N_28088);
nor UO_1519 (O_1519,N_25760,N_26388);
and UO_1520 (O_1520,N_27961,N_27917);
xor UO_1521 (O_1521,N_28265,N_29690);
or UO_1522 (O_1522,N_28752,N_26171);
and UO_1523 (O_1523,N_26372,N_28335);
and UO_1524 (O_1524,N_28317,N_25645);
xnor UO_1525 (O_1525,N_25389,N_29999);
xnor UO_1526 (O_1526,N_25299,N_27786);
nand UO_1527 (O_1527,N_25635,N_28075);
or UO_1528 (O_1528,N_26279,N_25461);
nand UO_1529 (O_1529,N_28612,N_26551);
xnor UO_1530 (O_1530,N_29354,N_25227);
nor UO_1531 (O_1531,N_25926,N_29007);
nand UO_1532 (O_1532,N_28478,N_29747);
or UO_1533 (O_1533,N_26817,N_25580);
and UO_1534 (O_1534,N_27211,N_25403);
or UO_1535 (O_1535,N_28031,N_26322);
nor UO_1536 (O_1536,N_26049,N_28055);
xnor UO_1537 (O_1537,N_25140,N_28398);
or UO_1538 (O_1538,N_25306,N_25216);
nand UO_1539 (O_1539,N_28028,N_25649);
nand UO_1540 (O_1540,N_27895,N_27252);
xor UO_1541 (O_1541,N_28984,N_29148);
xnor UO_1542 (O_1542,N_27143,N_28591);
or UO_1543 (O_1543,N_29064,N_28238);
or UO_1544 (O_1544,N_26793,N_28118);
and UO_1545 (O_1545,N_29631,N_26263);
nand UO_1546 (O_1546,N_27625,N_26904);
nand UO_1547 (O_1547,N_27599,N_26366);
and UO_1548 (O_1548,N_25116,N_26636);
or UO_1549 (O_1549,N_29256,N_29596);
and UO_1550 (O_1550,N_28204,N_28092);
nor UO_1551 (O_1551,N_25457,N_28948);
xor UO_1552 (O_1552,N_28782,N_29624);
xnor UO_1553 (O_1553,N_25348,N_25213);
or UO_1554 (O_1554,N_26742,N_27378);
nor UO_1555 (O_1555,N_28739,N_26635);
and UO_1556 (O_1556,N_29762,N_26739);
or UO_1557 (O_1557,N_28278,N_28320);
nor UO_1558 (O_1558,N_25159,N_28199);
and UO_1559 (O_1559,N_28179,N_26350);
or UO_1560 (O_1560,N_28150,N_25367);
nor UO_1561 (O_1561,N_27226,N_29002);
and UO_1562 (O_1562,N_25236,N_29287);
and UO_1563 (O_1563,N_26803,N_25888);
nor UO_1564 (O_1564,N_27780,N_27913);
nor UO_1565 (O_1565,N_26992,N_29821);
nand UO_1566 (O_1566,N_26673,N_25263);
xor UO_1567 (O_1567,N_26015,N_26059);
nand UO_1568 (O_1568,N_28546,N_25862);
nand UO_1569 (O_1569,N_28267,N_29988);
nor UO_1570 (O_1570,N_26492,N_25853);
and UO_1571 (O_1571,N_27185,N_25105);
and UO_1572 (O_1572,N_27063,N_27027);
and UO_1573 (O_1573,N_28205,N_28512);
xnor UO_1574 (O_1574,N_25417,N_27792);
and UO_1575 (O_1575,N_27820,N_25037);
or UO_1576 (O_1576,N_25337,N_28670);
nor UO_1577 (O_1577,N_29283,N_27400);
and UO_1578 (O_1578,N_28671,N_26052);
nand UO_1579 (O_1579,N_28313,N_25228);
nor UO_1580 (O_1580,N_26642,N_26326);
and UO_1581 (O_1581,N_26878,N_26069);
or UO_1582 (O_1582,N_25258,N_26504);
nor UO_1583 (O_1583,N_26124,N_28145);
and UO_1584 (O_1584,N_27671,N_27195);
nor UO_1585 (O_1585,N_25841,N_27613);
nor UO_1586 (O_1586,N_27314,N_27958);
xor UO_1587 (O_1587,N_26684,N_25154);
nand UO_1588 (O_1588,N_26663,N_25284);
and UO_1589 (O_1589,N_25949,N_26011);
xor UO_1590 (O_1590,N_28971,N_25929);
xor UO_1591 (O_1591,N_25131,N_27349);
nor UO_1592 (O_1592,N_28949,N_28081);
nor UO_1593 (O_1593,N_28111,N_27770);
and UO_1594 (O_1594,N_27289,N_28475);
or UO_1595 (O_1595,N_25864,N_28488);
or UO_1596 (O_1596,N_29171,N_28509);
and UO_1597 (O_1597,N_29275,N_26122);
xor UO_1598 (O_1598,N_26078,N_27609);
nand UO_1599 (O_1599,N_25807,N_28221);
xor UO_1600 (O_1600,N_28524,N_28065);
or UO_1601 (O_1601,N_25292,N_27391);
xnor UO_1602 (O_1602,N_27878,N_29516);
or UO_1603 (O_1603,N_29904,N_28135);
nor UO_1604 (O_1604,N_25145,N_28433);
xor UO_1605 (O_1605,N_29787,N_28852);
xor UO_1606 (O_1606,N_28332,N_25120);
xnor UO_1607 (O_1607,N_28559,N_25328);
and UO_1608 (O_1608,N_26567,N_28786);
nor UO_1609 (O_1609,N_25646,N_25496);
and UO_1610 (O_1610,N_26443,N_27565);
or UO_1611 (O_1611,N_26415,N_28647);
xnor UO_1612 (O_1612,N_28983,N_28357);
nand UO_1613 (O_1613,N_27470,N_25780);
nand UO_1614 (O_1614,N_28068,N_25464);
xor UO_1615 (O_1615,N_26886,N_26008);
nand UO_1616 (O_1616,N_28735,N_29099);
or UO_1617 (O_1617,N_27718,N_29898);
or UO_1618 (O_1618,N_28177,N_26277);
nand UO_1619 (O_1619,N_26248,N_29262);
or UO_1620 (O_1620,N_27677,N_28151);
nand UO_1621 (O_1621,N_29125,N_28053);
xor UO_1622 (O_1622,N_28371,N_26160);
nand UO_1623 (O_1623,N_29939,N_28833);
nand UO_1624 (O_1624,N_28299,N_26880);
or UO_1625 (O_1625,N_28076,N_27443);
nand UO_1626 (O_1626,N_28854,N_25914);
and UO_1627 (O_1627,N_29871,N_27442);
and UO_1628 (O_1628,N_28039,N_27468);
nand UO_1629 (O_1629,N_27073,N_25557);
or UO_1630 (O_1630,N_25362,N_25353);
nand UO_1631 (O_1631,N_25202,N_29773);
nor UO_1632 (O_1632,N_25293,N_26316);
xnor UO_1633 (O_1633,N_27603,N_26744);
xor UO_1634 (O_1634,N_28926,N_28289);
or UO_1635 (O_1635,N_28355,N_26446);
nor UO_1636 (O_1636,N_28080,N_29807);
and UO_1637 (O_1637,N_28403,N_25973);
nor UO_1638 (O_1638,N_29264,N_27558);
nand UO_1639 (O_1639,N_29206,N_28160);
or UO_1640 (O_1640,N_25548,N_26497);
xor UO_1641 (O_1641,N_25569,N_25309);
nand UO_1642 (O_1642,N_26864,N_27959);
nor UO_1643 (O_1643,N_28713,N_25903);
nand UO_1644 (O_1644,N_28896,N_28511);
nor UO_1645 (O_1645,N_28476,N_25877);
nand UO_1646 (O_1646,N_28905,N_27973);
xor UO_1647 (O_1647,N_27454,N_29968);
nor UO_1648 (O_1648,N_29134,N_25541);
nand UO_1649 (O_1649,N_26813,N_28192);
and UO_1650 (O_1650,N_27888,N_29594);
xor UO_1651 (O_1651,N_25723,N_29293);
nand UO_1652 (O_1652,N_27330,N_25527);
xor UO_1653 (O_1653,N_28535,N_27513);
nor UO_1654 (O_1654,N_29806,N_25731);
or UO_1655 (O_1655,N_27793,N_25278);
nor UO_1656 (O_1656,N_26364,N_25721);
or UO_1657 (O_1657,N_25897,N_26665);
nand UO_1658 (O_1658,N_26871,N_27815);
nand UO_1659 (O_1659,N_27554,N_29351);
xor UO_1660 (O_1660,N_25022,N_26874);
nand UO_1661 (O_1661,N_28967,N_28809);
xnor UO_1662 (O_1662,N_29228,N_29097);
nor UO_1663 (O_1663,N_26954,N_27485);
nor UO_1664 (O_1664,N_29302,N_27413);
nand UO_1665 (O_1665,N_25544,N_27134);
nand UO_1666 (O_1666,N_27320,N_27262);
and UO_1667 (O_1667,N_25215,N_28142);
xor UO_1668 (O_1668,N_29963,N_28128);
nor UO_1669 (O_1669,N_27552,N_28555);
nor UO_1670 (O_1670,N_29921,N_29746);
and UO_1671 (O_1671,N_27217,N_26855);
or UO_1672 (O_1672,N_25149,N_26118);
nor UO_1673 (O_1673,N_25295,N_27038);
or UO_1674 (O_1674,N_28628,N_25716);
nand UO_1675 (O_1675,N_28188,N_26007);
xnor UO_1676 (O_1676,N_25315,N_26195);
or UO_1677 (O_1677,N_25699,N_25705);
nor UO_1678 (O_1678,N_26965,N_25967);
and UO_1679 (O_1679,N_26783,N_29267);
nand UO_1680 (O_1680,N_25795,N_26578);
xor UO_1681 (O_1681,N_27566,N_25905);
nand UO_1682 (O_1682,N_25796,N_27580);
nand UO_1683 (O_1683,N_27214,N_28010);
xor UO_1684 (O_1684,N_26445,N_28420);
nor UO_1685 (O_1685,N_27897,N_25061);
and UO_1686 (O_1686,N_25327,N_27175);
nand UO_1687 (O_1687,N_25846,N_28777);
or UO_1688 (O_1688,N_29196,N_29727);
or UO_1689 (O_1689,N_25219,N_25325);
or UO_1690 (O_1690,N_26236,N_25036);
and UO_1691 (O_1691,N_26022,N_28029);
xor UO_1692 (O_1692,N_27923,N_25889);
xnor UO_1693 (O_1693,N_28586,N_29677);
nor UO_1694 (O_1694,N_25880,N_26437);
nand UO_1695 (O_1695,N_28176,N_28767);
xor UO_1696 (O_1696,N_26035,N_28024);
or UO_1697 (O_1697,N_28720,N_26831);
and UO_1698 (O_1698,N_25469,N_26311);
nor UO_1699 (O_1699,N_25071,N_25053);
nand UO_1700 (O_1700,N_28761,N_26056);
or UO_1701 (O_1701,N_27309,N_27386);
and UO_1702 (O_1702,N_29203,N_29908);
nor UO_1703 (O_1703,N_29408,N_25400);
or UO_1704 (O_1704,N_29144,N_29603);
or UO_1705 (O_1705,N_28668,N_25579);
nand UO_1706 (O_1706,N_28129,N_27325);
or UO_1707 (O_1707,N_26461,N_29161);
and UO_1708 (O_1708,N_28688,N_28772);
or UO_1709 (O_1709,N_25587,N_26344);
and UO_1710 (O_1710,N_27843,N_29229);
nand UO_1711 (O_1711,N_29749,N_28964);
nand UO_1712 (O_1712,N_26976,N_27506);
nor UO_1713 (O_1713,N_29083,N_29732);
and UO_1714 (O_1714,N_28649,N_28651);
or UO_1715 (O_1715,N_29869,N_26559);
nor UO_1716 (O_1716,N_26051,N_29076);
and UO_1717 (O_1717,N_26841,N_28832);
nor UO_1718 (O_1718,N_28449,N_25811);
nand UO_1719 (O_1719,N_29880,N_26879);
nor UO_1720 (O_1720,N_26402,N_25381);
nor UO_1721 (O_1721,N_29386,N_29604);
xor UO_1722 (O_1722,N_27497,N_29340);
nor UO_1723 (O_1723,N_26157,N_27324);
or UO_1724 (O_1724,N_29471,N_26961);
or UO_1725 (O_1725,N_28244,N_29579);
and UO_1726 (O_1726,N_26509,N_28303);
nor UO_1727 (O_1727,N_27021,N_25384);
nor UO_1728 (O_1728,N_26013,N_25653);
xnor UO_1729 (O_1729,N_27264,N_25467);
nand UO_1730 (O_1730,N_27492,N_29460);
and UO_1731 (O_1731,N_27546,N_26936);
nand UO_1732 (O_1732,N_25694,N_25130);
nor UO_1733 (O_1733,N_27043,N_27117);
and UO_1734 (O_1734,N_26800,N_25625);
nor UO_1735 (O_1735,N_28570,N_28307);
or UO_1736 (O_1736,N_27760,N_29185);
and UO_1737 (O_1737,N_25622,N_28656);
and UO_1738 (O_1738,N_26293,N_29614);
or UO_1739 (O_1739,N_27177,N_27221);
and UO_1740 (O_1740,N_26390,N_29178);
nand UO_1741 (O_1741,N_27178,N_25924);
nor UO_1742 (O_1742,N_29557,N_28066);
or UO_1743 (O_1743,N_27103,N_28405);
nand UO_1744 (O_1744,N_26472,N_26019);
nand UO_1745 (O_1745,N_26395,N_28359);
nand UO_1746 (O_1746,N_25451,N_27042);
or UO_1747 (O_1747,N_29034,N_25692);
nor UO_1748 (O_1748,N_27666,N_29636);
or UO_1749 (O_1749,N_28411,N_25755);
xor UO_1750 (O_1750,N_26257,N_29014);
and UO_1751 (O_1751,N_29887,N_29397);
nor UO_1752 (O_1752,N_25127,N_26393);
xnor UO_1753 (O_1753,N_25179,N_27367);
xor UO_1754 (O_1754,N_28025,N_29345);
and UO_1755 (O_1755,N_28991,N_26869);
or UO_1756 (O_1756,N_26270,N_29544);
nor UO_1757 (O_1757,N_25574,N_26408);
nor UO_1758 (O_1758,N_26205,N_26274);
nand UO_1759 (O_1759,N_27435,N_27555);
nand UO_1760 (O_1760,N_25872,N_28074);
xnor UO_1761 (O_1761,N_28463,N_25822);
xnor UO_1762 (O_1762,N_28804,N_26025);
xor UO_1763 (O_1763,N_29994,N_29670);
nand UO_1764 (O_1764,N_25452,N_28541);
and UO_1765 (O_1765,N_29425,N_25277);
nor UO_1766 (O_1766,N_28780,N_28286);
or UO_1767 (O_1767,N_29548,N_27517);
or UO_1768 (O_1768,N_29147,N_26233);
nor UO_1769 (O_1769,N_28614,N_27564);
nor UO_1770 (O_1770,N_29661,N_26363);
nand UO_1771 (O_1771,N_27444,N_25333);
and UO_1772 (O_1772,N_27791,N_29731);
nor UO_1773 (O_1773,N_27560,N_25651);
and UO_1774 (O_1774,N_25458,N_27104);
nor UO_1775 (O_1775,N_27288,N_27997);
nand UO_1776 (O_1776,N_26058,N_25787);
and UO_1777 (O_1777,N_28636,N_28582);
and UO_1778 (O_1778,N_27279,N_27855);
and UO_1779 (O_1779,N_27771,N_29699);
or UO_1780 (O_1780,N_28441,N_25593);
or UO_1781 (O_1781,N_25955,N_27099);
and UO_1782 (O_1782,N_25919,N_26029);
nor UO_1783 (O_1783,N_27769,N_29884);
xor UO_1784 (O_1784,N_27761,N_29783);
nand UO_1785 (O_1785,N_28144,N_28828);
nor UO_1786 (O_1786,N_28414,N_28722);
nor UO_1787 (O_1787,N_25601,N_29651);
nand UO_1788 (O_1788,N_25682,N_29017);
and UO_1789 (O_1789,N_26077,N_27359);
nor UO_1790 (O_1790,N_29098,N_25069);
or UO_1791 (O_1791,N_29804,N_25920);
nor UO_1792 (O_1792,N_29140,N_29463);
xor UO_1793 (O_1793,N_27904,N_27364);
nand UO_1794 (O_1794,N_27084,N_29011);
nor UO_1795 (O_1795,N_25545,N_27543);
xnor UO_1796 (O_1796,N_28704,N_25043);
nor UO_1797 (O_1797,N_25917,N_28935);
nand UO_1798 (O_1798,N_25708,N_26474);
or UO_1799 (O_1799,N_28663,N_27493);
nand UO_1800 (O_1800,N_28282,N_29647);
nor UO_1801 (O_1801,N_25429,N_29979);
and UO_1802 (O_1802,N_26584,N_27797);
xor UO_1803 (O_1803,N_29127,N_25009);
and UO_1804 (O_1804,N_25734,N_27830);
nor UO_1805 (O_1805,N_28788,N_25528);
xor UO_1806 (O_1806,N_27803,N_27907);
xor UO_1807 (O_1807,N_27536,N_25733);
nor UO_1808 (O_1808,N_29876,N_28881);
and UO_1809 (O_1809,N_28141,N_27964);
nor UO_1810 (O_1810,N_29067,N_25621);
or UO_1811 (O_1811,N_28379,N_26995);
or UO_1812 (O_1812,N_27007,N_28568);
and UO_1813 (O_1813,N_27198,N_26799);
xor UO_1814 (O_1814,N_29427,N_25256);
or UO_1815 (O_1815,N_29488,N_29190);
nor UO_1816 (O_1816,N_29430,N_25565);
or UO_1817 (O_1817,N_26860,N_29805);
nor UO_1818 (O_1818,N_25732,N_26717);
nand UO_1819 (O_1819,N_27816,N_27227);
xnor UO_1820 (O_1820,N_25481,N_26231);
nor UO_1821 (O_1821,N_28538,N_26988);
xor UO_1822 (O_1822,N_27388,N_28086);
xor UO_1823 (O_1823,N_26232,N_25576);
nor UO_1824 (O_1824,N_27654,N_27946);
or UO_1825 (O_1825,N_28897,N_29467);
or UO_1826 (O_1826,N_27795,N_29606);
nor UO_1827 (O_1827,N_25921,N_29473);
nor UO_1828 (O_1828,N_28050,N_27161);
nor UO_1829 (O_1829,N_27466,N_25197);
nor UO_1830 (O_1830,N_27699,N_27750);
or UO_1831 (O_1831,N_26034,N_25169);
nor UO_1832 (O_1832,N_27995,N_27659);
and UO_1833 (O_1833,N_25235,N_29141);
nor UO_1834 (O_1834,N_29515,N_29357);
or UO_1835 (O_1835,N_27450,N_27036);
and UO_1836 (O_1836,N_27488,N_29753);
xor UO_1837 (O_1837,N_25013,N_27620);
xnor UO_1838 (O_1838,N_26791,N_28729);
and UO_1839 (O_1839,N_29220,N_27202);
and UO_1840 (O_1840,N_25095,N_25449);
nor UO_1841 (O_1841,N_26239,N_29401);
or UO_1842 (O_1842,N_25503,N_29032);
nand UO_1843 (O_1843,N_29901,N_26127);
nor UO_1844 (O_1844,N_28173,N_28862);
or UO_1845 (O_1845,N_25606,N_25218);
nand UO_1846 (O_1846,N_29096,N_27507);
xor UO_1847 (O_1847,N_27887,N_28272);
and UO_1848 (O_1848,N_27653,N_25308);
or UO_1849 (O_1849,N_25255,N_26544);
and UO_1850 (O_1850,N_25492,N_26300);
nand UO_1851 (O_1851,N_26618,N_28802);
or UO_1852 (O_1852,N_28918,N_28023);
or UO_1853 (O_1853,N_27332,N_28279);
or UO_1854 (O_1854,N_25455,N_28269);
nor UO_1855 (O_1855,N_26048,N_28266);
xor UO_1856 (O_1856,N_29105,N_29894);
nor UO_1857 (O_1857,N_29927,N_26761);
xor UO_1858 (O_1858,N_28213,N_26529);
and UO_1859 (O_1859,N_28121,N_25490);
xnor UO_1860 (O_1860,N_27088,N_25126);
nor UO_1861 (O_1861,N_28021,N_28961);
and UO_1862 (O_1862,N_27561,N_25443);
nand UO_1863 (O_1863,N_27794,N_27661);
and UO_1864 (O_1864,N_27449,N_29772);
nor UO_1865 (O_1865,N_29626,N_26641);
nand UO_1866 (O_1866,N_26956,N_29605);
xor UO_1867 (O_1867,N_28855,N_28938);
nand UO_1868 (O_1868,N_27628,N_26228);
or UO_1869 (O_1869,N_25266,N_29601);
nand UO_1870 (O_1870,N_26962,N_25509);
and UO_1871 (O_1871,N_25636,N_27556);
nor UO_1872 (O_1872,N_28666,N_25520);
or UO_1873 (O_1873,N_29412,N_28284);
and UO_1874 (O_1874,N_25657,N_29465);
and UO_1875 (O_1875,N_27287,N_25663);
nor UO_1876 (O_1876,N_28607,N_27668);
and UO_1877 (O_1877,N_27121,N_25726);
and UO_1878 (O_1878,N_27156,N_26952);
nor UO_1879 (O_1879,N_26792,N_27819);
or UO_1880 (O_1880,N_25925,N_27208);
xor UO_1881 (O_1881,N_28134,N_29827);
or UO_1882 (O_1882,N_25983,N_27885);
and UO_1883 (O_1883,N_28376,N_26724);
nor UO_1884 (O_1884,N_29400,N_27728);
and UO_1885 (O_1885,N_26265,N_27698);
and UO_1886 (O_1886,N_25988,N_25835);
xnor UO_1887 (O_1887,N_27249,N_25749);
or UO_1888 (O_1888,N_26064,N_29719);
nor UO_1889 (O_1889,N_27688,N_27576);
xor UO_1890 (O_1890,N_27831,N_26839);
nor UO_1891 (O_1891,N_25489,N_26475);
nand UO_1892 (O_1892,N_29193,N_25104);
or UO_1893 (O_1893,N_29599,N_25482);
nor UO_1894 (O_1894,N_27385,N_29131);
nand UO_1895 (O_1895,N_27763,N_27859);
xor UO_1896 (O_1896,N_26146,N_29990);
and UO_1897 (O_1897,N_28159,N_26993);
and UO_1898 (O_1898,N_28494,N_25724);
or UO_1899 (O_1899,N_27254,N_27665);
or UO_1900 (O_1900,N_25763,N_27165);
nor UO_1901 (O_1901,N_27257,N_27925);
nor UO_1902 (O_1902,N_29945,N_29505);
nand UO_1903 (O_1903,N_25752,N_29905);
and UO_1904 (O_1904,N_26186,N_26394);
xnor UO_1905 (O_1905,N_26690,N_27173);
and UO_1906 (O_1906,N_28375,N_27774);
nor UO_1907 (O_1907,N_27854,N_27932);
xnor UO_1908 (O_1908,N_26646,N_29492);
nor UO_1909 (O_1909,N_25259,N_26950);
and UO_1910 (O_1910,N_25331,N_25420);
xnor UO_1911 (O_1911,N_28923,N_29906);
nor UO_1912 (O_1912,N_26737,N_29343);
xnor UO_1913 (O_1913,N_26568,N_28248);
or UO_1914 (O_1914,N_26189,N_25504);
xnor UO_1915 (O_1915,N_28781,N_27703);
nor UO_1916 (O_1916,N_26660,N_29587);
nand UO_1917 (O_1917,N_28985,N_27685);
nor UO_1918 (O_1918,N_27823,N_27374);
or UO_1919 (O_1919,N_26282,N_29883);
or UO_1920 (O_1920,N_25096,N_28620);
nand UO_1921 (O_1921,N_25188,N_26604);
xnor UO_1922 (O_1922,N_27721,N_25203);
or UO_1923 (O_1923,N_29019,N_25431);
or UO_1924 (O_1924,N_27154,N_27727);
xor UO_1925 (O_1925,N_28951,N_29846);
or UO_1926 (O_1926,N_25058,N_25220);
xor UO_1927 (O_1927,N_26359,N_29291);
and UO_1928 (O_1928,N_26809,N_29735);
or UO_1929 (O_1929,N_29513,N_26994);
nand UO_1930 (O_1930,N_25436,N_27271);
nand UO_1931 (O_1931,N_29170,N_29276);
and UO_1932 (O_1932,N_28208,N_28425);
nor UO_1933 (O_1933,N_25341,N_26389);
nand UO_1934 (O_1934,N_29058,N_25106);
nor UO_1935 (O_1935,N_27187,N_29258);
xnor UO_1936 (O_1936,N_27639,N_28430);
or UO_1937 (O_1937,N_28831,N_26715);
nor UO_1938 (O_1938,N_26801,N_29669);
or UO_1939 (O_1939,N_28575,N_29376);
and UO_1940 (O_1940,N_28793,N_26648);
nand UO_1941 (O_1941,N_28389,N_28288);
xnor UO_1942 (O_1942,N_25184,N_26203);
nor UO_1943 (O_1943,N_27781,N_26434);
or UO_1944 (O_1944,N_29864,N_27006);
nor UO_1945 (O_1945,N_27375,N_27147);
and UO_1946 (O_1946,N_26254,N_25533);
nor UO_1947 (O_1947,N_29240,N_27874);
and UO_1948 (O_1948,N_27804,N_28171);
and UO_1949 (O_1949,N_27168,N_28200);
nand UO_1950 (O_1950,N_27138,N_26703);
xor UO_1951 (O_1951,N_29977,N_26892);
xnor UO_1952 (O_1952,N_25262,N_25115);
nand UO_1953 (O_1953,N_25124,N_29943);
nand UO_1954 (O_1954,N_27982,N_28241);
and UO_1955 (O_1955,N_26006,N_26558);
or UO_1956 (O_1956,N_28132,N_27438);
or UO_1957 (O_1957,N_28243,N_25468);
nor UO_1958 (O_1958,N_29418,N_27201);
nor UO_1959 (O_1959,N_26154,N_26464);
nor UO_1960 (O_1960,N_29414,N_26422);
nand UO_1961 (O_1961,N_28471,N_27091);
or UO_1962 (O_1962,N_26334,N_26917);
or UO_1963 (O_1963,N_27581,N_29166);
and UO_1964 (O_1964,N_26500,N_29362);
and UO_1965 (O_1965,N_26130,N_28768);
nand UO_1966 (O_1966,N_27130,N_26946);
nand UO_1967 (O_1967,N_25537,N_27729);
nand UO_1968 (O_1968,N_25638,N_28263);
xnor UO_1969 (O_1969,N_26261,N_27460);
xor UO_1970 (O_1970,N_27200,N_27102);
nand UO_1971 (O_1971,N_26680,N_28378);
or UO_1972 (O_1972,N_29211,N_25589);
nand UO_1973 (O_1973,N_29251,N_25600);
xnor UO_1974 (O_1974,N_25478,N_29713);
xor UO_1975 (O_1975,N_28567,N_28152);
xor UO_1976 (O_1976,N_25129,N_28743);
and UO_1977 (O_1977,N_27209,N_28506);
or UO_1978 (O_1978,N_28755,N_26807);
or UO_1979 (O_1979,N_28540,N_27953);
xor UO_1980 (O_1980,N_26288,N_29115);
and UO_1981 (O_1981,N_28334,N_29545);
xor UO_1982 (O_1982,N_27233,N_28693);
and UO_1983 (O_1983,N_25985,N_28723);
xor UO_1984 (O_1984,N_27246,N_27985);
nand UO_1985 (O_1985,N_27741,N_26102);
or UO_1986 (O_1986,N_27336,N_25186);
nor UO_1987 (O_1987,N_29145,N_29930);
and UO_1988 (O_1988,N_27857,N_29223);
nand UO_1989 (O_1989,N_27282,N_28453);
xnor UO_1990 (O_1990,N_25172,N_26570);
nor UO_1991 (O_1991,N_28597,N_26918);
and UO_1992 (O_1992,N_27011,N_27709);
and UO_1993 (O_1993,N_29485,N_25250);
xor UO_1994 (O_1994,N_27502,N_28104);
or UO_1995 (O_1995,N_26973,N_25522);
and UO_1996 (O_1996,N_29768,N_25791);
xor UO_1997 (O_1997,N_27409,N_28699);
and UO_1998 (O_1998,N_29448,N_26275);
nor UO_1999 (O_1999,N_29701,N_25874);
xnor UO_2000 (O_2000,N_29057,N_27341);
or UO_2001 (O_2001,N_27921,N_26651);
nand UO_2002 (O_2002,N_27927,N_27660);
and UO_2003 (O_2003,N_27631,N_28368);
nand UO_2004 (O_2004,N_28975,N_29113);
or UO_2005 (O_2005,N_25815,N_27787);
xor UO_2006 (O_2006,N_29023,N_25827);
or UO_2007 (O_2007,N_29261,N_27204);
and UO_2008 (O_2008,N_28912,N_26877);
nand UO_2009 (O_2009,N_26543,N_25260);
nor UO_2010 (O_2010,N_26844,N_29564);
and UO_2011 (O_2011,N_28386,N_25660);
nor UO_2012 (O_2012,N_29615,N_29586);
or UO_2013 (O_2013,N_27111,N_25135);
nor UO_2014 (O_2014,N_26565,N_27571);
nor UO_2015 (O_2015,N_26330,N_25294);
xor UO_2016 (O_2016,N_25196,N_27758);
and UO_2017 (O_2017,N_26915,N_27626);
nor UO_2018 (O_2018,N_26369,N_28822);
or UO_2019 (O_2019,N_28472,N_25647);
nor UO_2020 (O_2020,N_27128,N_27199);
and UO_2021 (O_2021,N_26115,N_25831);
and UO_2022 (O_2022,N_28113,N_28479);
nand UO_2023 (O_2023,N_28432,N_27207);
nor UO_2024 (O_2024,N_29993,N_26707);
xnor UO_2025 (O_2025,N_25237,N_29868);
xnor UO_2026 (O_2026,N_27037,N_29659);
or UO_2027 (O_2027,N_25212,N_29922);
xnor UO_2028 (O_2028,N_28360,N_29572);
or UO_2029 (O_2029,N_29797,N_29658);
and UO_2030 (O_2030,N_25153,N_28632);
nand UO_2031 (O_2031,N_26292,N_26328);
nand UO_2032 (O_2032,N_28749,N_29897);
nand UO_2033 (O_2033,N_27587,N_27030);
and UO_2034 (O_2034,N_28517,N_29946);
nand UO_2035 (O_2035,N_26972,N_25542);
or UO_2036 (O_2036,N_28459,N_28519);
nand UO_2037 (O_2037,N_28886,N_25532);
nand UO_2038 (O_2038,N_25837,N_25814);
nand UO_2039 (O_2039,N_26091,N_27231);
and UO_2040 (O_2040,N_27749,N_28316);
nand UO_2041 (O_2041,N_25195,N_27474);
and UO_2042 (O_2042,N_28040,N_29483);
and UO_2043 (O_2043,N_27747,N_25626);
nand UO_2044 (O_2044,N_28940,N_27601);
nand UO_2045 (O_2045,N_27963,N_27281);
nor UO_2046 (O_2046,N_28170,N_26417);
nand UO_2047 (O_2047,N_25415,N_29165);
nand UO_2048 (O_2048,N_28158,N_29392);
nand UO_2049 (O_2049,N_29693,N_29667);
or UO_2050 (O_2050,N_27589,N_26720);
and UO_2051 (O_2051,N_27807,N_25487);
or UO_2052 (O_2052,N_25356,N_26215);
nor UO_2053 (O_2053,N_27313,N_28798);
and UO_2054 (O_2054,N_28642,N_28989);
and UO_2055 (O_2055,N_26109,N_28872);
nand UO_2056 (O_2056,N_27672,N_26633);
and UO_2057 (O_2057,N_26889,N_25540);
nor UO_2058 (O_2058,N_29910,N_29865);
or UO_2059 (O_2059,N_28426,N_28827);
nand UO_2060 (O_2060,N_29893,N_26816);
and UO_2061 (O_2061,N_28795,N_27940);
nor UO_2062 (O_2062,N_25007,N_27978);
or UO_2063 (O_2063,N_29627,N_25554);
or UO_2064 (O_2064,N_26404,N_28423);
or UO_2065 (O_2065,N_26573,N_29128);
nand UO_2066 (O_2066,N_29474,N_28495);
xnor UO_2067 (O_2067,N_29358,N_27980);
nor UO_2068 (O_2068,N_27648,N_27986);
nor UO_2069 (O_2069,N_29531,N_25291);
or UO_2070 (O_2070,N_26553,N_25064);
or UO_2071 (O_2071,N_27777,N_28576);
nand UO_2072 (O_2072,N_27473,N_25976);
nor UO_2073 (O_2073,N_29952,N_28042);
nand UO_2074 (O_2074,N_29550,N_27352);
xor UO_2075 (O_2075,N_26448,N_29075);
nor UO_2076 (O_2076,N_25141,N_28899);
and UO_2077 (O_2077,N_26572,N_27459);
or UO_2078 (O_2078,N_27189,N_27463);
and UO_2079 (O_2079,N_28480,N_25957);
nand UO_2080 (O_2080,N_26926,N_28584);
nor UO_2081 (O_2081,N_29499,N_29030);
nand UO_2082 (O_2082,N_28016,N_26209);
or UO_2083 (O_2083,N_25577,N_29172);
or UO_2084 (O_2084,N_29333,N_28101);
or UO_2085 (O_2085,N_29422,N_29652);
xnor UO_2086 (O_2086,N_27127,N_26657);
or UO_2087 (O_2087,N_28458,N_29439);
nand UO_2088 (O_2088,N_25017,N_28270);
xor UO_2089 (O_2089,N_26134,N_29817);
xnor UO_2090 (O_2090,N_29668,N_25330);
or UO_2091 (O_2091,N_26036,N_28439);
nor UO_2092 (O_2092,N_29839,N_27853);
and UO_2093 (O_2093,N_28030,N_29712);
nand UO_2094 (O_2094,N_28696,N_29808);
nand UO_2095 (O_2095,N_25214,N_28675);
nor UO_2096 (O_2096,N_25300,N_29389);
nand UO_2097 (O_2097,N_25097,N_28608);
xor UO_2098 (O_2098,N_29085,N_26629);
nand UO_2099 (O_2099,N_27441,N_28627);
nand UO_2100 (O_2100,N_29949,N_26581);
or UO_2101 (O_2101,N_28406,N_26747);
or UO_2102 (O_2102,N_28271,N_29527);
xnor UO_2103 (O_2103,N_27680,N_29632);
or UO_2104 (O_2104,N_28256,N_28644);
or UO_2105 (O_2105,N_26990,N_29214);
nand UO_2106 (O_2106,N_28849,N_29268);
xor UO_2107 (O_2107,N_25974,N_25845);
or UO_2108 (O_2108,N_26432,N_27746);
nor UO_2109 (O_2109,N_28147,N_26676);
xnor UO_2110 (O_2110,N_25534,N_25722);
and UO_2111 (O_2111,N_28291,N_25506);
xnor UO_2112 (O_2112,N_26106,N_28726);
xnor UO_2113 (O_2113,N_25114,N_26214);
and UO_2114 (O_2114,N_27167,N_29956);
nor UO_2115 (O_2115,N_28306,N_27179);
or UO_2116 (O_2116,N_27098,N_27477);
or UO_2117 (O_2117,N_25767,N_29576);
nor UO_2118 (O_2118,N_26688,N_28645);
nor UO_2119 (O_2119,N_27053,N_26614);
nand UO_2120 (O_2120,N_28452,N_26638);
nor UO_2121 (O_2121,N_25701,N_26762);
or UO_2122 (O_2122,N_28295,N_25191);
xnor UO_2123 (O_2123,N_26711,N_29300);
nand UO_2124 (O_2124,N_28245,N_28326);
nor UO_2125 (O_2125,N_25893,N_25883);
or UO_2126 (O_2126,N_26386,N_29909);
and UO_2127 (O_2127,N_29394,N_29018);
and UO_2128 (O_2128,N_27472,N_28060);
xor UO_2129 (O_2129,N_25435,N_29874);
xor UO_2130 (O_2130,N_28382,N_28944);
and UO_2131 (O_2131,N_26067,N_27714);
and UO_2132 (O_2132,N_28209,N_26094);
xnor UO_2133 (O_2133,N_29265,N_27933);
xnor UO_2134 (O_2134,N_25480,N_26158);
nor UO_2135 (O_2135,N_26563,N_27634);
and UO_2136 (O_2136,N_29061,N_27909);
nor UO_2137 (O_2137,N_29464,N_27651);
or UO_2138 (O_2138,N_25838,N_28090);
xnor UO_2139 (O_2139,N_27682,N_29859);
and UO_2140 (O_2140,N_26425,N_27315);
xor UO_2141 (O_2141,N_27020,N_26080);
or UO_2142 (O_2142,N_25230,N_28759);
nor UO_2143 (O_2143,N_25510,N_28874);
or UO_2144 (O_2144,N_28562,N_26613);
xor UO_2145 (O_2145,N_29517,N_25015);
nor UO_2146 (O_2146,N_28468,N_25960);
nand UO_2147 (O_2147,N_27344,N_29726);
and UO_2148 (O_2148,N_25366,N_28902);
nand UO_2149 (O_2149,N_28510,N_28958);
and UO_2150 (O_2150,N_27844,N_26964);
or UO_2151 (O_2151,N_26356,N_25865);
nor UO_2152 (O_2152,N_26299,N_29521);
nand UO_2153 (O_2153,N_27255,N_27166);
nand UO_2154 (O_2154,N_27942,N_28373);
and UO_2155 (O_2155,N_26043,N_27732);
or UO_2156 (O_2156,N_25750,N_27681);
nor UO_2157 (O_2157,N_26136,N_25344);
xor UO_2158 (O_2158,N_25840,N_27346);
or UO_2159 (O_2159,N_25972,N_29697);
nand UO_2160 (O_2160,N_28909,N_29266);
or UO_2161 (O_2161,N_28857,N_28564);
or UO_2162 (O_2162,N_25322,N_29481);
and UO_2163 (O_2163,N_25296,N_26368);
nand UO_2164 (O_2164,N_27916,N_26944);
xor UO_2165 (O_2165,N_25444,N_29123);
xor UO_2166 (O_2166,N_27503,N_25424);
and UO_2167 (O_2167,N_28421,N_27437);
nor UO_2168 (O_2168,N_29405,N_27243);
nand UO_2169 (O_2169,N_25632,N_25290);
and UO_2170 (O_2170,N_26608,N_27089);
or UO_2171 (O_2171,N_25836,N_28139);
or UO_2172 (O_2172,N_29928,N_28553);
and UO_2173 (O_2173,N_25592,N_27368);
or UO_2174 (O_2174,N_29974,N_26361);
and UO_2175 (O_2175,N_29524,N_29764);
and UO_2176 (O_2176,N_25794,N_26786);
nand UO_2177 (O_2177,N_29899,N_29973);
nor UO_2178 (O_2178,N_27095,N_29556);
xnor UO_2179 (O_2179,N_28993,N_28419);
or UO_2180 (O_2180,N_25741,N_25939);
nor UO_2181 (O_2181,N_27109,N_28812);
and UO_2182 (O_2182,N_29896,N_29509);
nand UO_2183 (O_2183,N_28707,N_27033);
xnor UO_2184 (O_2184,N_26396,N_29950);
or UO_2185 (O_2185,N_27419,N_25922);
or UO_2186 (O_2186,N_25430,N_29297);
xnor UO_2187 (O_2187,N_29932,N_25180);
and UO_2188 (O_2188,N_26743,N_26718);
xor UO_2189 (O_2189,N_28717,N_26845);
xor UO_2190 (O_2190,N_28347,N_26884);
nor UO_2191 (O_2191,N_27251,N_26619);
nor UO_2192 (O_2192,N_28621,N_29794);
and UO_2193 (O_2193,N_27148,N_28217);
xor UO_2194 (O_2194,N_28093,N_25551);
xor UO_2195 (O_2195,N_27024,N_29779);
nor UO_2196 (O_2196,N_27372,N_29635);
xnor UO_2197 (O_2197,N_29308,N_27646);
nor UO_2198 (O_2198,N_29204,N_28193);
nor UO_2199 (O_2199,N_28077,N_28230);
nor UO_2200 (O_2200,N_28837,N_29338);
or UO_2201 (O_2201,N_29366,N_29130);
xnor UO_2202 (O_2202,N_26137,N_25242);
or UO_2203 (O_2203,N_29541,N_27875);
and UO_2204 (O_2204,N_29553,N_26290);
or UO_2205 (O_2205,N_29306,N_25395);
and UO_2206 (O_2206,N_26414,N_29489);
xor UO_2207 (O_2207,N_25248,N_28758);
and UO_2208 (O_2208,N_25232,N_29660);
and UO_2209 (O_2209,N_25881,N_25642);
nand UO_2210 (O_2210,N_25427,N_27283);
nor UO_2211 (O_2211,N_28851,N_29335);
nor UO_2212 (O_2212,N_26545,N_25591);
and UO_2213 (O_2213,N_26131,N_27896);
or UO_2214 (O_2214,N_26285,N_25319);
nor UO_2215 (O_2215,N_27080,N_25773);
nand UO_2216 (O_2216,N_27440,N_29987);
and UO_2217 (O_2217,N_27962,N_29399);
xnor UO_2218 (O_2218,N_29852,N_26821);
and UO_2219 (O_2219,N_28513,N_26897);
nand UO_2220 (O_2220,N_28140,N_27619);
or UO_2221 (O_2221,N_26468,N_29707);
or UO_2222 (O_2222,N_26304,N_28516);
nand UO_2223 (O_2223,N_28745,N_28891);
and UO_2224 (O_2224,N_27675,N_26523);
or UO_2225 (O_2225,N_27067,N_29080);
xnor UO_2226 (O_2226,N_26784,N_29810);
nor UO_2227 (O_2227,N_27286,N_29282);
xor UO_2228 (O_2228,N_27881,N_29356);
nor UO_2229 (O_2229,N_26407,N_26452);
xnor UO_2230 (O_2230,N_29629,N_29008);
nand UO_2231 (O_2231,N_29168,N_27884);
nor UO_2232 (O_2232,N_27535,N_25584);
or UO_2233 (O_2233,N_26589,N_27266);
or UO_2234 (O_2234,N_28153,N_29770);
nor UO_2235 (O_2235,N_29194,N_29493);
nor UO_2236 (O_2236,N_27667,N_29998);
nand UO_2237 (O_2237,N_28203,N_29793);
nand UO_2238 (O_2238,N_28490,N_26773);
nand UO_2239 (O_2239,N_25282,N_26210);
or UO_2240 (O_2240,N_26355,N_26538);
xnor UO_2241 (O_2241,N_28344,N_27768);
nor UO_2242 (O_2242,N_29885,N_27421);
xnor UO_2243 (O_2243,N_27327,N_28166);
or UO_2244 (O_2244,N_26658,N_26001);
xor UO_2245 (O_2245,N_29155,N_26110);
or UO_2246 (O_2246,N_28435,N_29157);
or UO_2247 (O_2247,N_25563,N_27321);
nor UO_2248 (O_2248,N_28026,N_29253);
xnor UO_2249 (O_2249,N_29455,N_26607);
or UO_2250 (O_2250,N_29739,N_28061);
nor UO_2251 (O_2251,N_27553,N_28618);
and UO_2252 (O_2252,N_25937,N_25806);
and UO_2253 (O_2253,N_26155,N_26009);
or UO_2254 (O_2254,N_26620,N_27529);
and UO_2255 (O_2255,N_29339,N_28427);
and UO_2256 (O_2256,N_27612,N_25737);
xnor UO_2257 (O_2257,N_25044,N_29396);
or UO_2258 (O_2258,N_27559,N_26047);
xor UO_2259 (O_2259,N_27188,N_26708);
or UO_2260 (O_2260,N_25689,N_25779);
nand UO_2261 (O_2261,N_28634,N_26033);
or UO_2262 (O_2262,N_26709,N_25060);
and UO_2263 (O_2263,N_25358,N_29826);
and UO_2264 (O_2264,N_29029,N_26216);
xor UO_2265 (O_2265,N_29780,N_27331);
and UO_2266 (O_2266,N_27369,N_27149);
nand UO_2267 (O_2267,N_28692,N_29738);
xnor UO_2268 (O_2268,N_25170,N_25144);
nand UO_2269 (O_2269,N_28879,N_25904);
and UO_2270 (O_2270,N_27600,N_29237);
or UO_2271 (O_2271,N_26212,N_26481);
and UO_2272 (O_2272,N_27957,N_28732);
nor UO_2273 (O_2273,N_26406,N_28210);
and UO_2274 (O_2274,N_25505,N_29759);
and UO_2275 (O_2275,N_26741,N_25209);
nor UO_2276 (O_2276,N_27476,N_27645);
nor UO_2277 (O_2277,N_27563,N_27824);
or UO_2278 (O_2278,N_27532,N_28916);
nand UO_2279 (O_2279,N_26779,N_26719);
xnor UO_2280 (O_2280,N_29862,N_28602);
or UO_2281 (O_2281,N_27842,N_29406);
or UO_2282 (O_2282,N_28451,N_29649);
nand UO_2283 (O_2283,N_29470,N_28402);
nand UO_2284 (O_2284,N_29183,N_28338);
or UO_2285 (O_2285,N_25766,N_29815);
xnor UO_2286 (O_2286,N_28807,N_27610);
xnor UO_2287 (O_2287,N_29094,N_28108);
xor UO_2288 (O_2288,N_29964,N_29512);
xor UO_2289 (O_2289,N_28507,N_28550);
nor UO_2290 (O_2290,N_25683,N_29559);
nand UO_2291 (O_2291,N_27001,N_29960);
xnor UO_2292 (O_2292,N_28664,N_29702);
nor UO_2293 (O_2293,N_29164,N_29936);
or UO_2294 (O_2294,N_27693,N_27305);
xnor UO_2295 (O_2295,N_25168,N_27373);
xor UO_2296 (O_2296,N_28297,N_27411);
nand UO_2297 (O_2297,N_29895,N_27530);
or UO_2298 (O_2298,N_27125,N_25644);
nand UO_2299 (O_2299,N_28116,N_25999);
or UO_2300 (O_2300,N_26548,N_26084);
nor UO_2301 (O_2301,N_25615,N_26487);
or UO_2302 (O_2302,N_28771,N_26780);
nand UO_2303 (O_2303,N_29021,N_26194);
nand UO_2304 (O_2304,N_29991,N_28863);
nor UO_2305 (O_2305,N_28443,N_26562);
xnor UO_2306 (O_2306,N_27745,N_29188);
or UO_2307 (O_2307,N_25329,N_26093);
nor UO_2308 (O_2308,N_28370,N_27244);
or UO_2309 (O_2309,N_26556,N_25910);
nor UO_2310 (O_2310,N_26331,N_25162);
nor UO_2311 (O_2311,N_25373,N_25205);
nor UO_2312 (O_2312,N_29191,N_28063);
and UO_2313 (O_2313,N_27562,N_29352);
nor UO_2314 (O_2314,N_27382,N_25494);
nand UO_2315 (O_2315,N_27726,N_25610);
xor UO_2316 (O_2316,N_27097,N_25680);
nand UO_2317 (O_2317,N_29703,N_29568);
nand UO_2318 (O_2318,N_25422,N_29006);
xnor UO_2319 (O_2319,N_26188,N_28324);
or UO_2320 (O_2320,N_25832,N_26133);
xor UO_2321 (O_2321,N_25674,N_28845);
and UO_2322 (O_2322,N_26371,N_26240);
nor UO_2323 (O_2323,N_25690,N_27447);
or UO_2324 (O_2324,N_28189,N_27357);
and UO_2325 (O_2325,N_28148,N_25562);
or UO_2326 (O_2326,N_27464,N_26820);
xnor UO_2327 (O_2327,N_25177,N_25113);
xnor UO_2328 (O_2328,N_28920,N_27035);
nand UO_2329 (O_2329,N_28229,N_26204);
nand UO_2330 (O_2330,N_26018,N_26399);
nand UO_2331 (O_2331,N_25077,N_25107);
and UO_2332 (O_2332,N_25040,N_27118);
or UO_2333 (O_2333,N_27928,N_25623);
and UO_2334 (O_2334,N_25552,N_29847);
and UO_2335 (O_2335,N_29958,N_29832);
and UO_2336 (O_2336,N_25500,N_25018);
nand UO_2337 (O_2337,N_28175,N_27298);
nand UO_2338 (O_2338,N_28528,N_27054);
or UO_2339 (O_2339,N_27212,N_27491);
or UO_2340 (O_2340,N_27016,N_27096);
nand UO_2341 (O_2341,N_28114,N_25265);
nor UO_2342 (O_2342,N_29745,N_28011);
and UO_2343 (O_2343,N_26685,N_29590);
nor UO_2344 (O_2344,N_28789,N_28866);
nand UO_2345 (O_2345,N_26503,N_27623);
xor UO_2346 (O_2346,N_26580,N_27184);
nor UO_2347 (O_2347,N_25238,N_27839);
nor UO_2348 (O_2348,N_26116,N_29334);
or UO_2349 (O_2349,N_28917,N_25475);
xnor UO_2350 (O_2350,N_28321,N_29252);
nor UO_2351 (O_2351,N_27445,N_26539);
nand UO_2352 (O_2352,N_26998,N_29530);
and UO_2353 (O_2353,N_26387,N_26705);
xor UO_2354 (O_2354,N_29907,N_28572);
or UO_2355 (O_2355,N_27943,N_26125);
nand UO_2356 (O_2356,N_26939,N_29976);
nor UO_2357 (O_2357,N_28112,N_28820);
xor UO_2358 (O_2358,N_28500,N_28466);
xnor UO_2359 (O_2359,N_29890,N_27055);
and UO_2360 (O_2360,N_26413,N_28020);
and UO_2361 (O_2361,N_27481,N_26170);
or UO_2362 (O_2362,N_25123,N_25223);
and UO_2363 (O_2363,N_27123,N_27398);
nand UO_2364 (O_2364,N_25824,N_25411);
or UO_2365 (O_2365,N_28633,N_26085);
nor UO_2366 (O_2366,N_25661,N_29260);
or UO_2367 (O_2367,N_26323,N_25383);
nand UO_2368 (O_2368,N_28921,N_28873);
nand UO_2369 (O_2369,N_25030,N_29637);
and UO_2370 (O_2370,N_26550,N_28925);
xnor UO_2371 (O_2371,N_28504,N_27304);
xnor UO_2372 (O_2372,N_25187,N_29534);
or UO_2373 (O_2373,N_27735,N_29244);
nand UO_2374 (O_2374,N_25938,N_28805);
nor UO_2375 (O_2375,N_26631,N_29081);
xor UO_2376 (O_2376,N_26217,N_27077);
nor UO_2377 (O_2377,N_28587,N_25501);
xor UO_2378 (O_2378,N_28072,N_26574);
nand UO_2379 (O_2379,N_28611,N_29582);
nand UO_2380 (O_2380,N_26857,N_28138);
and UO_2381 (O_2381,N_29711,N_28900);
nand UO_2382 (O_2382,N_26379,N_25020);
or UO_2383 (O_2383,N_26746,N_25002);
xor UO_2384 (O_2384,N_27500,N_26107);
nand UO_2385 (O_2385,N_27048,N_28515);
and UO_2386 (O_2386,N_28652,N_29088);
or UO_2387 (O_2387,N_28281,N_28581);
or UO_2388 (O_2388,N_28631,N_26140);
xnor UO_2389 (O_2389,N_28084,N_29775);
or UO_2390 (O_2390,N_25948,N_26659);
or UO_2391 (O_2391,N_29813,N_29951);
xor UO_2392 (O_2392,N_26499,N_27840);
and UO_2393 (O_2393,N_29013,N_29676);
or UO_2394 (O_2394,N_27549,N_27434);
nor UO_2395 (O_2395,N_25072,N_25257);
or UO_2396 (O_2396,N_29638,N_29042);
or UO_2397 (O_2397,N_29359,N_29848);
nor UO_2398 (O_2398,N_29441,N_26100);
nand UO_2399 (O_2399,N_26600,N_25042);
xnor UO_2400 (O_2400,N_25484,N_27893);
nand UO_2401 (O_2401,N_26682,N_29831);
and UO_2402 (O_2402,N_28853,N_29217);
and UO_2403 (O_2403,N_27081,N_29317);
nor UO_2404 (O_2404,N_29476,N_25261);
xnor UO_2405 (O_2405,N_28493,N_29823);
nor UO_2406 (O_2406,N_25928,N_25391);
or UO_2407 (O_2407,N_25781,N_29420);
nor UO_2408 (O_2408,N_28098,N_29355);
or UO_2409 (O_2409,N_27017,N_28959);
nor UO_2410 (O_2410,N_25969,N_27508);
xor UO_2411 (O_2411,N_26349,N_26775);
nand UO_2412 (O_2412,N_29158,N_25738);
nand UO_2413 (O_2413,N_29068,N_28966);
or UO_2414 (O_2414,N_29740,N_29479);
and UO_2415 (O_2415,N_25735,N_29820);
nor UO_2416 (O_2416,N_28069,N_26766);
and UO_2417 (O_2417,N_27847,N_27849);
xor UO_2418 (O_2418,N_28560,N_29881);
nand UO_2419 (O_2419,N_27141,N_26245);
nor UO_2420 (O_2420,N_29344,N_28534);
nand UO_2421 (O_2421,N_27335,N_27297);
or UO_2422 (O_2422,N_26790,N_28149);
and UO_2423 (O_2423,N_29452,N_28034);
nor UO_2424 (O_2424,N_26306,N_25932);
or UO_2425 (O_2425,N_26505,N_27293);
xor UO_2426 (O_2426,N_25821,N_25181);
nor UO_2427 (O_2427,N_26143,N_25332);
nor UO_2428 (O_2428,N_25525,N_27310);
or UO_2429 (O_2429,N_25873,N_27427);
or UO_2430 (O_2430,N_27423,N_29109);
nor UO_2431 (O_2431,N_27284,N_25078);
xor UO_2432 (O_2432,N_27192,N_29154);
nand UO_2433 (O_2433,N_26940,N_28356);
xnor UO_2434 (O_2434,N_27649,N_26327);
or UO_2435 (O_2435,N_29248,N_28687);
and UO_2436 (O_2436,N_28924,N_25830);
and UO_2437 (O_2437,N_29053,N_25380);
or UO_2438 (O_2438,N_25101,N_27724);
or UO_2439 (O_2439,N_28672,N_28362);
or UO_2440 (O_2440,N_28174,N_26206);
nand UO_2441 (O_2441,N_29200,N_29938);
nand UO_2442 (O_2442,N_29114,N_29784);
xor UO_2443 (O_2443,N_29522,N_29449);
nand UO_2444 (O_2444,N_25902,N_27181);
xnor UO_2445 (O_2445,N_28491,N_26482);
nor UO_2446 (O_2446,N_27338,N_29024);
and UO_2447 (O_2447,N_28259,N_27169);
nand UO_2448 (O_2448,N_28319,N_28613);
and UO_2449 (O_2449,N_28557,N_29849);
and UO_2450 (O_2450,N_28701,N_26230);
nor UO_2451 (O_2451,N_28184,N_25090);
or UO_2452 (O_2452,N_28943,N_29696);
or UO_2453 (O_2453,N_28276,N_28950);
xor UO_2454 (O_2454,N_26576,N_28473);
nand UO_2455 (O_2455,N_29304,N_25961);
and UO_2456 (O_2456,N_28684,N_26987);
and UO_2457 (O_2457,N_25117,N_26853);
and UO_2458 (O_2458,N_27322,N_28790);
or UO_2459 (O_2459,N_27334,N_28604);
and UO_2460 (O_2460,N_29216,N_28470);
or UO_2461 (O_2461,N_26074,N_25867);
or UO_2462 (O_2462,N_26455,N_27767);
and UO_2463 (O_2463,N_28052,N_28246);
xnor UO_2464 (O_2464,N_29038,N_26179);
nor UO_2465 (O_2465,N_26024,N_27700);
xor UO_2466 (O_2466,N_25656,N_25594);
nor UO_2467 (O_2467,N_27919,N_26712);
xnor UO_2468 (O_2468,N_26338,N_28952);
nor UO_2469 (O_2469,N_25804,N_27547);
nand UO_2470 (O_2470,N_27268,N_28521);
xnor UO_2471 (O_2471,N_29777,N_29838);
and UO_2472 (O_2472,N_27432,N_29484);
and UO_2473 (O_2473,N_27790,N_26923);
or UO_2474 (O_2474,N_27783,N_26901);
and UO_2475 (O_2475,N_27295,N_26440);
xor UO_2476 (O_2476,N_25704,N_27852);
nor UO_2477 (O_2477,N_26062,N_26028);
nand UO_2478 (O_2478,N_26498,N_29600);
nor UO_2479 (O_2479,N_27263,N_27348);
xor UO_2480 (O_2480,N_27939,N_27025);
and UO_2481 (O_2481,N_29242,N_27363);
and UO_2482 (O_2482,N_25231,N_25033);
nand UO_2483 (O_2483,N_27392,N_25239);
and UO_2484 (O_2484,N_26061,N_27278);
and UO_2485 (O_2485,N_29117,N_27082);
and UO_2486 (O_2486,N_26315,N_28492);
or UO_2487 (O_2487,N_26272,N_28779);
and UO_2488 (O_2488,N_28216,N_25244);
xnor UO_2489 (O_2489,N_25693,N_26090);
or UO_2490 (O_2490,N_26032,N_27779);
or UO_2491 (O_2491,N_27737,N_27360);
xor UO_2492 (O_2492,N_26854,N_25070);
xnor UO_2493 (O_2493,N_28051,N_25673);
and UO_2494 (O_2494,N_25119,N_29423);
nand UO_2495 (O_2495,N_26842,N_25067);
nand UO_2496 (O_2496,N_27124,N_29858);
nor UO_2497 (O_2497,N_26764,N_26900);
and UO_2498 (O_2498,N_29571,N_27494);
and UO_2499 (O_2499,N_27241,N_29913);
nand UO_2500 (O_2500,N_26039,N_27890);
nor UO_2501 (O_2501,N_25412,N_28313);
nand UO_2502 (O_2502,N_29538,N_26801);
xor UO_2503 (O_2503,N_25658,N_29044);
nand UO_2504 (O_2504,N_25109,N_29575);
nand UO_2505 (O_2505,N_25317,N_29137);
xnor UO_2506 (O_2506,N_28191,N_26997);
and UO_2507 (O_2507,N_27522,N_25343);
or UO_2508 (O_2508,N_29467,N_26733);
and UO_2509 (O_2509,N_28645,N_28936);
nor UO_2510 (O_2510,N_28152,N_29080);
nand UO_2511 (O_2511,N_26054,N_28111);
and UO_2512 (O_2512,N_28742,N_25973);
nand UO_2513 (O_2513,N_26700,N_26327);
xor UO_2514 (O_2514,N_25246,N_28358);
xnor UO_2515 (O_2515,N_27884,N_25095);
nor UO_2516 (O_2516,N_27979,N_27935);
and UO_2517 (O_2517,N_26008,N_27676);
xnor UO_2518 (O_2518,N_29227,N_25432);
or UO_2519 (O_2519,N_29855,N_29311);
nor UO_2520 (O_2520,N_28237,N_26383);
and UO_2521 (O_2521,N_26059,N_28431);
and UO_2522 (O_2522,N_28403,N_28102);
nand UO_2523 (O_2523,N_27700,N_26800);
xnor UO_2524 (O_2524,N_27000,N_26830);
nand UO_2525 (O_2525,N_29099,N_29983);
or UO_2526 (O_2526,N_27205,N_25284);
nand UO_2527 (O_2527,N_29069,N_28532);
or UO_2528 (O_2528,N_25304,N_28511);
nor UO_2529 (O_2529,N_26474,N_25846);
nor UO_2530 (O_2530,N_29216,N_25382);
nand UO_2531 (O_2531,N_27505,N_25056);
nand UO_2532 (O_2532,N_29347,N_28824);
nor UO_2533 (O_2533,N_29764,N_29732);
nand UO_2534 (O_2534,N_29611,N_28938);
or UO_2535 (O_2535,N_26640,N_25467);
nor UO_2536 (O_2536,N_29873,N_25995);
or UO_2537 (O_2537,N_29229,N_27611);
xnor UO_2538 (O_2538,N_27545,N_26764);
nand UO_2539 (O_2539,N_25789,N_26249);
xnor UO_2540 (O_2540,N_29375,N_25364);
xor UO_2541 (O_2541,N_29439,N_26827);
xor UO_2542 (O_2542,N_26950,N_26127);
nor UO_2543 (O_2543,N_28284,N_26452);
and UO_2544 (O_2544,N_25542,N_27338);
nand UO_2545 (O_2545,N_25920,N_29853);
nand UO_2546 (O_2546,N_29186,N_29534);
or UO_2547 (O_2547,N_27528,N_25872);
nor UO_2548 (O_2548,N_25138,N_25211);
and UO_2549 (O_2549,N_29233,N_27093);
nand UO_2550 (O_2550,N_28418,N_29513);
and UO_2551 (O_2551,N_27095,N_27170);
and UO_2552 (O_2552,N_28253,N_29741);
nor UO_2553 (O_2553,N_29324,N_29835);
xnor UO_2554 (O_2554,N_25122,N_28368);
or UO_2555 (O_2555,N_25945,N_27248);
nor UO_2556 (O_2556,N_25945,N_27352);
nand UO_2557 (O_2557,N_26791,N_25591);
xor UO_2558 (O_2558,N_25312,N_27619);
or UO_2559 (O_2559,N_28602,N_27399);
and UO_2560 (O_2560,N_29150,N_25073);
and UO_2561 (O_2561,N_26095,N_25277);
and UO_2562 (O_2562,N_27332,N_25647);
and UO_2563 (O_2563,N_29388,N_27459);
nand UO_2564 (O_2564,N_28406,N_25958);
xor UO_2565 (O_2565,N_25288,N_27003);
nand UO_2566 (O_2566,N_29615,N_28774);
nor UO_2567 (O_2567,N_29122,N_28888);
or UO_2568 (O_2568,N_26872,N_29708);
or UO_2569 (O_2569,N_27866,N_26464);
or UO_2570 (O_2570,N_29775,N_25759);
or UO_2571 (O_2571,N_25998,N_29220);
xnor UO_2572 (O_2572,N_28755,N_27903);
and UO_2573 (O_2573,N_26907,N_29699);
xnor UO_2574 (O_2574,N_26168,N_25138);
and UO_2575 (O_2575,N_25388,N_28723);
and UO_2576 (O_2576,N_26414,N_26029);
nor UO_2577 (O_2577,N_28355,N_27807);
xnor UO_2578 (O_2578,N_25237,N_26355);
nor UO_2579 (O_2579,N_27589,N_25014);
xnor UO_2580 (O_2580,N_28894,N_29219);
nand UO_2581 (O_2581,N_28120,N_29860);
nand UO_2582 (O_2582,N_25613,N_27387);
nor UO_2583 (O_2583,N_28677,N_29161);
nor UO_2584 (O_2584,N_27325,N_28535);
nor UO_2585 (O_2585,N_29875,N_26912);
nor UO_2586 (O_2586,N_28131,N_29451);
nor UO_2587 (O_2587,N_25211,N_27823);
xnor UO_2588 (O_2588,N_26062,N_28915);
or UO_2589 (O_2589,N_26956,N_25579);
xor UO_2590 (O_2590,N_29512,N_28932);
nand UO_2591 (O_2591,N_28903,N_28056);
xnor UO_2592 (O_2592,N_29898,N_27789);
nor UO_2593 (O_2593,N_27068,N_26978);
and UO_2594 (O_2594,N_25561,N_29130);
nand UO_2595 (O_2595,N_27512,N_28648);
or UO_2596 (O_2596,N_25753,N_27761);
xor UO_2597 (O_2597,N_26901,N_28560);
and UO_2598 (O_2598,N_26524,N_27376);
nand UO_2599 (O_2599,N_27289,N_29131);
nor UO_2600 (O_2600,N_29372,N_25820);
or UO_2601 (O_2601,N_25718,N_26328);
xor UO_2602 (O_2602,N_29630,N_26889);
nand UO_2603 (O_2603,N_28276,N_29832);
or UO_2604 (O_2604,N_29940,N_28654);
nor UO_2605 (O_2605,N_29079,N_27560);
nand UO_2606 (O_2606,N_25460,N_25163);
and UO_2607 (O_2607,N_27203,N_25738);
nand UO_2608 (O_2608,N_27763,N_26425);
nor UO_2609 (O_2609,N_28803,N_29747);
nand UO_2610 (O_2610,N_27852,N_26961);
and UO_2611 (O_2611,N_26525,N_25559);
and UO_2612 (O_2612,N_27417,N_26855);
nand UO_2613 (O_2613,N_26344,N_25192);
or UO_2614 (O_2614,N_27046,N_27991);
nand UO_2615 (O_2615,N_26588,N_27853);
or UO_2616 (O_2616,N_29027,N_29810);
or UO_2617 (O_2617,N_26783,N_28093);
xor UO_2618 (O_2618,N_25427,N_28825);
or UO_2619 (O_2619,N_28610,N_25884);
xor UO_2620 (O_2620,N_28062,N_25976);
or UO_2621 (O_2621,N_25923,N_25575);
xnor UO_2622 (O_2622,N_27236,N_27539);
xnor UO_2623 (O_2623,N_26721,N_26762);
or UO_2624 (O_2624,N_29253,N_27245);
xnor UO_2625 (O_2625,N_27795,N_25682);
nand UO_2626 (O_2626,N_26114,N_25135);
nand UO_2627 (O_2627,N_26542,N_26021);
or UO_2628 (O_2628,N_28417,N_28746);
and UO_2629 (O_2629,N_27411,N_29540);
nand UO_2630 (O_2630,N_25439,N_26054);
nand UO_2631 (O_2631,N_28018,N_28950);
and UO_2632 (O_2632,N_29793,N_27102);
nor UO_2633 (O_2633,N_27060,N_25071);
nor UO_2634 (O_2634,N_29173,N_26570);
nor UO_2635 (O_2635,N_26871,N_28245);
nor UO_2636 (O_2636,N_25302,N_27547);
nand UO_2637 (O_2637,N_29794,N_29849);
xnor UO_2638 (O_2638,N_29599,N_26435);
xnor UO_2639 (O_2639,N_28916,N_27425);
and UO_2640 (O_2640,N_29595,N_29354);
nand UO_2641 (O_2641,N_28841,N_27016);
nor UO_2642 (O_2642,N_25792,N_27303);
and UO_2643 (O_2643,N_26106,N_29355);
nor UO_2644 (O_2644,N_28458,N_28413);
and UO_2645 (O_2645,N_27431,N_28294);
nand UO_2646 (O_2646,N_25634,N_27848);
xnor UO_2647 (O_2647,N_28348,N_26705);
and UO_2648 (O_2648,N_25492,N_26297);
or UO_2649 (O_2649,N_29656,N_25854);
and UO_2650 (O_2650,N_29230,N_28601);
and UO_2651 (O_2651,N_25656,N_25481);
or UO_2652 (O_2652,N_27265,N_25424);
and UO_2653 (O_2653,N_25512,N_29776);
or UO_2654 (O_2654,N_27017,N_29967);
nand UO_2655 (O_2655,N_29018,N_29296);
xnor UO_2656 (O_2656,N_27806,N_25323);
nand UO_2657 (O_2657,N_26355,N_25125);
nand UO_2658 (O_2658,N_28245,N_28926);
and UO_2659 (O_2659,N_27907,N_29449);
nand UO_2660 (O_2660,N_28655,N_27504);
nand UO_2661 (O_2661,N_28725,N_25733);
and UO_2662 (O_2662,N_26131,N_26377);
xor UO_2663 (O_2663,N_27551,N_28389);
and UO_2664 (O_2664,N_29267,N_29364);
or UO_2665 (O_2665,N_25152,N_25193);
xnor UO_2666 (O_2666,N_27924,N_26539);
xor UO_2667 (O_2667,N_28707,N_29387);
xnor UO_2668 (O_2668,N_27314,N_26745);
nand UO_2669 (O_2669,N_27908,N_27605);
xor UO_2670 (O_2670,N_29972,N_28448);
and UO_2671 (O_2671,N_28429,N_29384);
and UO_2672 (O_2672,N_28175,N_26840);
or UO_2673 (O_2673,N_25800,N_26676);
xnor UO_2674 (O_2674,N_26917,N_25165);
and UO_2675 (O_2675,N_26805,N_27129);
xnor UO_2676 (O_2676,N_26322,N_25715);
nand UO_2677 (O_2677,N_28940,N_28243);
or UO_2678 (O_2678,N_29918,N_29062);
and UO_2679 (O_2679,N_27668,N_28147);
and UO_2680 (O_2680,N_27235,N_25953);
and UO_2681 (O_2681,N_27593,N_25024);
nor UO_2682 (O_2682,N_26469,N_29067);
or UO_2683 (O_2683,N_25055,N_26067);
nor UO_2684 (O_2684,N_29694,N_28349);
xnor UO_2685 (O_2685,N_27691,N_28630);
or UO_2686 (O_2686,N_29787,N_29109);
or UO_2687 (O_2687,N_28454,N_28193);
nor UO_2688 (O_2688,N_29392,N_28784);
xor UO_2689 (O_2689,N_26193,N_27903);
and UO_2690 (O_2690,N_26629,N_26080);
nor UO_2691 (O_2691,N_27230,N_28059);
xor UO_2692 (O_2692,N_28272,N_27893);
or UO_2693 (O_2693,N_28897,N_29945);
nor UO_2694 (O_2694,N_26802,N_26176);
nand UO_2695 (O_2695,N_25259,N_26807);
xor UO_2696 (O_2696,N_28338,N_29066);
xor UO_2697 (O_2697,N_29663,N_28361);
and UO_2698 (O_2698,N_28718,N_28741);
nor UO_2699 (O_2699,N_25866,N_29189);
or UO_2700 (O_2700,N_27986,N_29636);
nor UO_2701 (O_2701,N_29077,N_26920);
and UO_2702 (O_2702,N_28488,N_28080);
nand UO_2703 (O_2703,N_29704,N_29959);
nand UO_2704 (O_2704,N_28489,N_25720);
or UO_2705 (O_2705,N_26054,N_27939);
nor UO_2706 (O_2706,N_27553,N_26743);
or UO_2707 (O_2707,N_27955,N_25603);
nor UO_2708 (O_2708,N_25620,N_29453);
or UO_2709 (O_2709,N_26596,N_27174);
xor UO_2710 (O_2710,N_25239,N_26384);
xor UO_2711 (O_2711,N_26119,N_26296);
nor UO_2712 (O_2712,N_28675,N_29865);
nor UO_2713 (O_2713,N_26795,N_29112);
nor UO_2714 (O_2714,N_29956,N_29860);
nor UO_2715 (O_2715,N_28445,N_27868);
xnor UO_2716 (O_2716,N_27326,N_25729);
nand UO_2717 (O_2717,N_27082,N_25062);
or UO_2718 (O_2718,N_25128,N_28261);
and UO_2719 (O_2719,N_28387,N_25098);
nor UO_2720 (O_2720,N_29085,N_27356);
or UO_2721 (O_2721,N_27754,N_28854);
and UO_2722 (O_2722,N_26815,N_26046);
nand UO_2723 (O_2723,N_26700,N_27638);
xor UO_2724 (O_2724,N_27365,N_27809);
nand UO_2725 (O_2725,N_27706,N_29954);
nand UO_2726 (O_2726,N_25226,N_29643);
and UO_2727 (O_2727,N_27469,N_26893);
or UO_2728 (O_2728,N_28751,N_27059);
or UO_2729 (O_2729,N_28561,N_28312);
nand UO_2730 (O_2730,N_26552,N_27575);
xnor UO_2731 (O_2731,N_29220,N_25287);
nor UO_2732 (O_2732,N_26822,N_27875);
xor UO_2733 (O_2733,N_28780,N_29429);
nand UO_2734 (O_2734,N_26013,N_27343);
or UO_2735 (O_2735,N_25718,N_25628);
nand UO_2736 (O_2736,N_25104,N_25061);
nand UO_2737 (O_2737,N_27667,N_28422);
or UO_2738 (O_2738,N_28996,N_28418);
or UO_2739 (O_2739,N_26169,N_29522);
or UO_2740 (O_2740,N_29238,N_29569);
xor UO_2741 (O_2741,N_28763,N_27420);
nand UO_2742 (O_2742,N_29487,N_25590);
or UO_2743 (O_2743,N_29151,N_27398);
xor UO_2744 (O_2744,N_26399,N_26336);
nor UO_2745 (O_2745,N_28953,N_27204);
nor UO_2746 (O_2746,N_25906,N_29623);
and UO_2747 (O_2747,N_29931,N_26431);
nand UO_2748 (O_2748,N_26891,N_27455);
or UO_2749 (O_2749,N_26366,N_27750);
nor UO_2750 (O_2750,N_25787,N_28219);
xor UO_2751 (O_2751,N_26139,N_28456);
nor UO_2752 (O_2752,N_26530,N_25778);
or UO_2753 (O_2753,N_29765,N_25367);
nand UO_2754 (O_2754,N_25419,N_29168);
xnor UO_2755 (O_2755,N_25696,N_26502);
xor UO_2756 (O_2756,N_26682,N_26847);
and UO_2757 (O_2757,N_28025,N_25727);
or UO_2758 (O_2758,N_25027,N_27834);
nand UO_2759 (O_2759,N_25088,N_25721);
and UO_2760 (O_2760,N_25109,N_26393);
or UO_2761 (O_2761,N_25554,N_25496);
nand UO_2762 (O_2762,N_29292,N_28178);
nand UO_2763 (O_2763,N_26679,N_25315);
or UO_2764 (O_2764,N_29453,N_25655);
nor UO_2765 (O_2765,N_26324,N_29494);
and UO_2766 (O_2766,N_27142,N_29323);
and UO_2767 (O_2767,N_29259,N_28720);
nand UO_2768 (O_2768,N_25976,N_27758);
nor UO_2769 (O_2769,N_27183,N_28592);
and UO_2770 (O_2770,N_28795,N_29837);
nand UO_2771 (O_2771,N_28634,N_27217);
xor UO_2772 (O_2772,N_25558,N_29436);
nor UO_2773 (O_2773,N_25094,N_26826);
xor UO_2774 (O_2774,N_27650,N_28897);
xnor UO_2775 (O_2775,N_29096,N_25418);
nor UO_2776 (O_2776,N_26560,N_27439);
nor UO_2777 (O_2777,N_29342,N_29722);
nand UO_2778 (O_2778,N_29935,N_28450);
nor UO_2779 (O_2779,N_27237,N_28274);
xor UO_2780 (O_2780,N_27951,N_25381);
nand UO_2781 (O_2781,N_25939,N_26298);
nor UO_2782 (O_2782,N_25814,N_25084);
nor UO_2783 (O_2783,N_29260,N_27131);
xor UO_2784 (O_2784,N_26580,N_27687);
xor UO_2785 (O_2785,N_29802,N_27337);
or UO_2786 (O_2786,N_29292,N_27095);
and UO_2787 (O_2787,N_26106,N_29987);
or UO_2788 (O_2788,N_27378,N_25997);
nor UO_2789 (O_2789,N_27723,N_25324);
xor UO_2790 (O_2790,N_26637,N_29378);
nand UO_2791 (O_2791,N_25306,N_25789);
nor UO_2792 (O_2792,N_26737,N_26433);
and UO_2793 (O_2793,N_25274,N_25020);
xor UO_2794 (O_2794,N_26310,N_25679);
xnor UO_2795 (O_2795,N_25547,N_26457);
nand UO_2796 (O_2796,N_28145,N_28647);
nand UO_2797 (O_2797,N_27000,N_26142);
and UO_2798 (O_2798,N_25911,N_26263);
xnor UO_2799 (O_2799,N_29657,N_29060);
and UO_2800 (O_2800,N_26875,N_26085);
nor UO_2801 (O_2801,N_25629,N_25693);
or UO_2802 (O_2802,N_26043,N_26357);
or UO_2803 (O_2803,N_29981,N_27322);
or UO_2804 (O_2804,N_25656,N_28185);
or UO_2805 (O_2805,N_28970,N_27176);
nor UO_2806 (O_2806,N_28816,N_26400);
nand UO_2807 (O_2807,N_27111,N_26516);
xnor UO_2808 (O_2808,N_29210,N_28353);
nand UO_2809 (O_2809,N_26878,N_28465);
nor UO_2810 (O_2810,N_28519,N_26207);
nand UO_2811 (O_2811,N_25115,N_26687);
nand UO_2812 (O_2812,N_29814,N_28463);
xor UO_2813 (O_2813,N_26635,N_29374);
and UO_2814 (O_2814,N_28048,N_27282);
or UO_2815 (O_2815,N_28071,N_29779);
xor UO_2816 (O_2816,N_29568,N_25293);
nand UO_2817 (O_2817,N_28439,N_26961);
nand UO_2818 (O_2818,N_25308,N_25306);
nand UO_2819 (O_2819,N_26004,N_27222);
nor UO_2820 (O_2820,N_27638,N_28198);
and UO_2821 (O_2821,N_26642,N_28322);
nand UO_2822 (O_2822,N_29349,N_27682);
nor UO_2823 (O_2823,N_29729,N_26798);
nand UO_2824 (O_2824,N_26811,N_26653);
and UO_2825 (O_2825,N_28418,N_28469);
and UO_2826 (O_2826,N_26340,N_28005);
nand UO_2827 (O_2827,N_27606,N_29479);
nor UO_2828 (O_2828,N_26131,N_28195);
nor UO_2829 (O_2829,N_29505,N_26577);
or UO_2830 (O_2830,N_27315,N_29223);
nand UO_2831 (O_2831,N_25644,N_28469);
or UO_2832 (O_2832,N_28355,N_26253);
and UO_2833 (O_2833,N_26346,N_26080);
or UO_2834 (O_2834,N_28638,N_27867);
nor UO_2835 (O_2835,N_29095,N_29418);
nor UO_2836 (O_2836,N_25397,N_28046);
nor UO_2837 (O_2837,N_26104,N_26417);
nand UO_2838 (O_2838,N_27994,N_26149);
and UO_2839 (O_2839,N_25841,N_25301);
and UO_2840 (O_2840,N_29678,N_25540);
nand UO_2841 (O_2841,N_28340,N_28026);
nor UO_2842 (O_2842,N_28140,N_26002);
and UO_2843 (O_2843,N_27487,N_28956);
nand UO_2844 (O_2844,N_28394,N_25130);
nand UO_2845 (O_2845,N_29418,N_25982);
or UO_2846 (O_2846,N_25732,N_28797);
nand UO_2847 (O_2847,N_27675,N_25033);
nor UO_2848 (O_2848,N_26202,N_26375);
or UO_2849 (O_2849,N_28443,N_29007);
nand UO_2850 (O_2850,N_27625,N_26224);
xor UO_2851 (O_2851,N_26117,N_29921);
nor UO_2852 (O_2852,N_28611,N_26830);
nor UO_2853 (O_2853,N_26525,N_27337);
or UO_2854 (O_2854,N_25554,N_27283);
xor UO_2855 (O_2855,N_26388,N_26695);
xnor UO_2856 (O_2856,N_28618,N_25973);
nand UO_2857 (O_2857,N_29203,N_25592);
xor UO_2858 (O_2858,N_26974,N_28519);
nand UO_2859 (O_2859,N_27227,N_26741);
or UO_2860 (O_2860,N_28145,N_28402);
xor UO_2861 (O_2861,N_25771,N_25648);
and UO_2862 (O_2862,N_27953,N_26627);
nand UO_2863 (O_2863,N_29216,N_27590);
xor UO_2864 (O_2864,N_25914,N_26062);
nand UO_2865 (O_2865,N_26895,N_27242);
xor UO_2866 (O_2866,N_27284,N_25324);
nand UO_2867 (O_2867,N_25642,N_26146);
nor UO_2868 (O_2868,N_26611,N_27249);
nor UO_2869 (O_2869,N_28428,N_27632);
or UO_2870 (O_2870,N_28892,N_29281);
nor UO_2871 (O_2871,N_29202,N_25616);
nand UO_2872 (O_2872,N_25407,N_26991);
xnor UO_2873 (O_2873,N_29025,N_27920);
xnor UO_2874 (O_2874,N_29461,N_26382);
nand UO_2875 (O_2875,N_25918,N_25851);
and UO_2876 (O_2876,N_29636,N_26057);
or UO_2877 (O_2877,N_29922,N_26662);
and UO_2878 (O_2878,N_29794,N_25908);
nor UO_2879 (O_2879,N_26211,N_29593);
or UO_2880 (O_2880,N_25930,N_27044);
xnor UO_2881 (O_2881,N_29062,N_25267);
nor UO_2882 (O_2882,N_29376,N_29657);
xor UO_2883 (O_2883,N_29057,N_29740);
nand UO_2884 (O_2884,N_27000,N_28606);
nand UO_2885 (O_2885,N_28013,N_29030);
xor UO_2886 (O_2886,N_26362,N_29558);
or UO_2887 (O_2887,N_29111,N_29493);
xor UO_2888 (O_2888,N_26218,N_25641);
nor UO_2889 (O_2889,N_25497,N_29280);
nor UO_2890 (O_2890,N_28045,N_28322);
nor UO_2891 (O_2891,N_29028,N_29598);
or UO_2892 (O_2892,N_26154,N_25623);
or UO_2893 (O_2893,N_26573,N_28604);
nand UO_2894 (O_2894,N_29474,N_29485);
and UO_2895 (O_2895,N_29093,N_28603);
nand UO_2896 (O_2896,N_29504,N_27889);
and UO_2897 (O_2897,N_27485,N_25638);
nor UO_2898 (O_2898,N_25966,N_25784);
or UO_2899 (O_2899,N_29248,N_25031);
xor UO_2900 (O_2900,N_25768,N_27989);
or UO_2901 (O_2901,N_26550,N_28176);
nand UO_2902 (O_2902,N_26615,N_25997);
xor UO_2903 (O_2903,N_28901,N_29903);
nor UO_2904 (O_2904,N_28179,N_25676);
xnor UO_2905 (O_2905,N_27475,N_28913);
or UO_2906 (O_2906,N_28975,N_25951);
xnor UO_2907 (O_2907,N_29606,N_26251);
or UO_2908 (O_2908,N_29209,N_26417);
nand UO_2909 (O_2909,N_29379,N_26404);
nor UO_2910 (O_2910,N_25703,N_28946);
nor UO_2911 (O_2911,N_25748,N_26989);
nor UO_2912 (O_2912,N_27179,N_25496);
nand UO_2913 (O_2913,N_26401,N_28871);
and UO_2914 (O_2914,N_25064,N_28651);
nor UO_2915 (O_2915,N_26216,N_29326);
nor UO_2916 (O_2916,N_28673,N_27142);
xnor UO_2917 (O_2917,N_25013,N_25346);
nor UO_2918 (O_2918,N_28980,N_25817);
or UO_2919 (O_2919,N_25557,N_25352);
xnor UO_2920 (O_2920,N_28478,N_27607);
and UO_2921 (O_2921,N_28895,N_26969);
nand UO_2922 (O_2922,N_25322,N_25481);
and UO_2923 (O_2923,N_27966,N_26117);
or UO_2924 (O_2924,N_28253,N_28934);
nand UO_2925 (O_2925,N_27212,N_29923);
or UO_2926 (O_2926,N_28928,N_28413);
xor UO_2927 (O_2927,N_27679,N_26611);
xnor UO_2928 (O_2928,N_25027,N_26411);
nand UO_2929 (O_2929,N_25421,N_26281);
xnor UO_2930 (O_2930,N_26504,N_26602);
nand UO_2931 (O_2931,N_28060,N_29078);
and UO_2932 (O_2932,N_25948,N_25608);
nor UO_2933 (O_2933,N_25846,N_25357);
or UO_2934 (O_2934,N_27861,N_25478);
and UO_2935 (O_2935,N_27259,N_28242);
nor UO_2936 (O_2936,N_28348,N_26414);
xor UO_2937 (O_2937,N_29866,N_25918);
xnor UO_2938 (O_2938,N_27716,N_26944);
nor UO_2939 (O_2939,N_29598,N_29074);
xor UO_2940 (O_2940,N_25873,N_25320);
nand UO_2941 (O_2941,N_25029,N_26076);
xor UO_2942 (O_2942,N_29170,N_27671);
xor UO_2943 (O_2943,N_29717,N_27342);
nor UO_2944 (O_2944,N_27016,N_28587);
nor UO_2945 (O_2945,N_25668,N_27211);
xor UO_2946 (O_2946,N_28951,N_25914);
xor UO_2947 (O_2947,N_28295,N_29135);
or UO_2948 (O_2948,N_26150,N_25565);
xor UO_2949 (O_2949,N_29387,N_28123);
nor UO_2950 (O_2950,N_25881,N_28612);
xor UO_2951 (O_2951,N_26797,N_26853);
nand UO_2952 (O_2952,N_26291,N_26965);
nor UO_2953 (O_2953,N_28236,N_27625);
and UO_2954 (O_2954,N_26416,N_25344);
nor UO_2955 (O_2955,N_25683,N_27435);
nand UO_2956 (O_2956,N_25103,N_26661);
or UO_2957 (O_2957,N_25699,N_29369);
and UO_2958 (O_2958,N_27846,N_26707);
and UO_2959 (O_2959,N_26736,N_25537);
nand UO_2960 (O_2960,N_28752,N_26574);
xor UO_2961 (O_2961,N_27590,N_25144);
xor UO_2962 (O_2962,N_29808,N_27036);
xnor UO_2963 (O_2963,N_28093,N_28894);
or UO_2964 (O_2964,N_26947,N_25795);
xnor UO_2965 (O_2965,N_25101,N_29407);
nor UO_2966 (O_2966,N_26266,N_28818);
or UO_2967 (O_2967,N_29707,N_25605);
xnor UO_2968 (O_2968,N_29561,N_28863);
and UO_2969 (O_2969,N_28663,N_27564);
or UO_2970 (O_2970,N_25685,N_27228);
nor UO_2971 (O_2971,N_28340,N_26956);
and UO_2972 (O_2972,N_27189,N_26096);
or UO_2973 (O_2973,N_29239,N_27168);
and UO_2974 (O_2974,N_27474,N_26129);
and UO_2975 (O_2975,N_25949,N_29674);
nand UO_2976 (O_2976,N_27660,N_29694);
and UO_2977 (O_2977,N_26445,N_27750);
nand UO_2978 (O_2978,N_27187,N_26438);
xor UO_2979 (O_2979,N_26069,N_26011);
and UO_2980 (O_2980,N_25952,N_26605);
xnor UO_2981 (O_2981,N_27845,N_25713);
xnor UO_2982 (O_2982,N_29304,N_25196);
xor UO_2983 (O_2983,N_26802,N_25147);
or UO_2984 (O_2984,N_26547,N_25087);
nand UO_2985 (O_2985,N_26902,N_25214);
or UO_2986 (O_2986,N_26615,N_26767);
or UO_2987 (O_2987,N_26138,N_27639);
nor UO_2988 (O_2988,N_25043,N_25796);
nor UO_2989 (O_2989,N_27309,N_28448);
nor UO_2990 (O_2990,N_29970,N_29602);
and UO_2991 (O_2991,N_26895,N_29357);
or UO_2992 (O_2992,N_25115,N_26828);
and UO_2993 (O_2993,N_25196,N_25264);
and UO_2994 (O_2994,N_28072,N_28112);
nor UO_2995 (O_2995,N_25923,N_28918);
xnor UO_2996 (O_2996,N_29951,N_27140);
nor UO_2997 (O_2997,N_26843,N_28850);
or UO_2998 (O_2998,N_25799,N_25120);
nand UO_2999 (O_2999,N_27556,N_25250);
or UO_3000 (O_3000,N_29787,N_28446);
and UO_3001 (O_3001,N_28217,N_27877);
nor UO_3002 (O_3002,N_29173,N_26274);
nand UO_3003 (O_3003,N_25305,N_29030);
nor UO_3004 (O_3004,N_28492,N_25322);
xnor UO_3005 (O_3005,N_27316,N_27102);
xnor UO_3006 (O_3006,N_25674,N_29624);
nand UO_3007 (O_3007,N_28375,N_27964);
or UO_3008 (O_3008,N_25871,N_29051);
or UO_3009 (O_3009,N_28080,N_29686);
xor UO_3010 (O_3010,N_29356,N_28356);
xor UO_3011 (O_3011,N_25114,N_25136);
nand UO_3012 (O_3012,N_25563,N_25344);
nand UO_3013 (O_3013,N_27371,N_28614);
nor UO_3014 (O_3014,N_25694,N_28391);
xnor UO_3015 (O_3015,N_27993,N_29377);
and UO_3016 (O_3016,N_25581,N_27409);
and UO_3017 (O_3017,N_28804,N_26284);
or UO_3018 (O_3018,N_29849,N_29158);
nor UO_3019 (O_3019,N_28274,N_26654);
xnor UO_3020 (O_3020,N_28530,N_29535);
or UO_3021 (O_3021,N_27648,N_25037);
nand UO_3022 (O_3022,N_28717,N_27284);
and UO_3023 (O_3023,N_29020,N_28354);
nand UO_3024 (O_3024,N_28767,N_27185);
nor UO_3025 (O_3025,N_27846,N_27923);
xor UO_3026 (O_3026,N_25553,N_26095);
nor UO_3027 (O_3027,N_26772,N_27378);
xnor UO_3028 (O_3028,N_28974,N_29643);
nor UO_3029 (O_3029,N_26873,N_26357);
and UO_3030 (O_3030,N_28024,N_26136);
and UO_3031 (O_3031,N_25185,N_28248);
or UO_3032 (O_3032,N_29531,N_25530);
nand UO_3033 (O_3033,N_25273,N_27021);
nor UO_3034 (O_3034,N_26204,N_28720);
or UO_3035 (O_3035,N_26518,N_28450);
and UO_3036 (O_3036,N_27154,N_25160);
nand UO_3037 (O_3037,N_25254,N_29206);
nor UO_3038 (O_3038,N_28690,N_29403);
nor UO_3039 (O_3039,N_29831,N_27779);
or UO_3040 (O_3040,N_27728,N_27405);
xnor UO_3041 (O_3041,N_26934,N_29155);
or UO_3042 (O_3042,N_25016,N_27762);
xor UO_3043 (O_3043,N_25203,N_27015);
nand UO_3044 (O_3044,N_25590,N_27325);
nor UO_3045 (O_3045,N_29109,N_29494);
and UO_3046 (O_3046,N_27622,N_29071);
xor UO_3047 (O_3047,N_29076,N_27818);
and UO_3048 (O_3048,N_25431,N_27561);
and UO_3049 (O_3049,N_26344,N_28148);
xor UO_3050 (O_3050,N_25909,N_27522);
or UO_3051 (O_3051,N_27525,N_28550);
nand UO_3052 (O_3052,N_29177,N_26227);
xnor UO_3053 (O_3053,N_28471,N_27417);
nand UO_3054 (O_3054,N_26045,N_28211);
nor UO_3055 (O_3055,N_27705,N_26931);
nor UO_3056 (O_3056,N_28042,N_27467);
and UO_3057 (O_3057,N_27258,N_29502);
nand UO_3058 (O_3058,N_26484,N_26541);
nand UO_3059 (O_3059,N_26284,N_26846);
xor UO_3060 (O_3060,N_25546,N_25322);
nor UO_3061 (O_3061,N_28081,N_28890);
xor UO_3062 (O_3062,N_27121,N_28991);
nand UO_3063 (O_3063,N_27324,N_25482);
or UO_3064 (O_3064,N_25181,N_27239);
or UO_3065 (O_3065,N_27936,N_29610);
and UO_3066 (O_3066,N_27932,N_28899);
nand UO_3067 (O_3067,N_29842,N_27112);
or UO_3068 (O_3068,N_26677,N_25540);
xor UO_3069 (O_3069,N_28828,N_26665);
nand UO_3070 (O_3070,N_28150,N_25706);
nor UO_3071 (O_3071,N_26390,N_26746);
nor UO_3072 (O_3072,N_25492,N_27417);
xnor UO_3073 (O_3073,N_28999,N_28836);
xor UO_3074 (O_3074,N_27342,N_27384);
nor UO_3075 (O_3075,N_27086,N_29446);
and UO_3076 (O_3076,N_27050,N_26795);
nand UO_3077 (O_3077,N_27408,N_29247);
or UO_3078 (O_3078,N_26544,N_26838);
nor UO_3079 (O_3079,N_28616,N_26685);
xor UO_3080 (O_3080,N_26492,N_26967);
xnor UO_3081 (O_3081,N_27923,N_27060);
xor UO_3082 (O_3082,N_28431,N_27592);
and UO_3083 (O_3083,N_29014,N_28702);
and UO_3084 (O_3084,N_28312,N_27047);
nor UO_3085 (O_3085,N_27908,N_27713);
or UO_3086 (O_3086,N_29745,N_28525);
or UO_3087 (O_3087,N_29566,N_28923);
nand UO_3088 (O_3088,N_29781,N_26208);
nand UO_3089 (O_3089,N_25568,N_28668);
nor UO_3090 (O_3090,N_29029,N_25853);
nor UO_3091 (O_3091,N_27968,N_25885);
or UO_3092 (O_3092,N_26628,N_28925);
nor UO_3093 (O_3093,N_25868,N_25192);
and UO_3094 (O_3094,N_27678,N_28105);
nand UO_3095 (O_3095,N_26721,N_26647);
or UO_3096 (O_3096,N_27865,N_25940);
nand UO_3097 (O_3097,N_27987,N_28164);
or UO_3098 (O_3098,N_25117,N_27912);
nand UO_3099 (O_3099,N_25500,N_28285);
xnor UO_3100 (O_3100,N_25232,N_25171);
nor UO_3101 (O_3101,N_25335,N_25281);
nand UO_3102 (O_3102,N_26651,N_25118);
xnor UO_3103 (O_3103,N_28997,N_26778);
or UO_3104 (O_3104,N_28745,N_28007);
or UO_3105 (O_3105,N_25661,N_28190);
nand UO_3106 (O_3106,N_28770,N_25230);
xor UO_3107 (O_3107,N_27884,N_27933);
xor UO_3108 (O_3108,N_25688,N_27885);
or UO_3109 (O_3109,N_27121,N_29887);
nor UO_3110 (O_3110,N_29492,N_26229);
xor UO_3111 (O_3111,N_29972,N_28489);
and UO_3112 (O_3112,N_28018,N_29612);
nor UO_3113 (O_3113,N_26887,N_27062);
nor UO_3114 (O_3114,N_27476,N_27382);
xnor UO_3115 (O_3115,N_25747,N_29097);
nand UO_3116 (O_3116,N_26512,N_27943);
xnor UO_3117 (O_3117,N_26748,N_26227);
and UO_3118 (O_3118,N_27588,N_25647);
and UO_3119 (O_3119,N_27248,N_25497);
or UO_3120 (O_3120,N_26479,N_26895);
nor UO_3121 (O_3121,N_25351,N_25714);
nand UO_3122 (O_3122,N_29542,N_29512);
xor UO_3123 (O_3123,N_27352,N_28822);
or UO_3124 (O_3124,N_25174,N_26470);
nor UO_3125 (O_3125,N_29619,N_28629);
and UO_3126 (O_3126,N_28398,N_27931);
or UO_3127 (O_3127,N_27028,N_25116);
nor UO_3128 (O_3128,N_29675,N_29079);
xnor UO_3129 (O_3129,N_25999,N_25520);
or UO_3130 (O_3130,N_26864,N_25168);
nand UO_3131 (O_3131,N_27459,N_29373);
nand UO_3132 (O_3132,N_26138,N_28188);
and UO_3133 (O_3133,N_28789,N_26787);
nor UO_3134 (O_3134,N_29499,N_29072);
and UO_3135 (O_3135,N_27081,N_25645);
and UO_3136 (O_3136,N_28621,N_27575);
nand UO_3137 (O_3137,N_27997,N_28750);
or UO_3138 (O_3138,N_28188,N_27794);
and UO_3139 (O_3139,N_28572,N_29840);
nor UO_3140 (O_3140,N_28498,N_25519);
or UO_3141 (O_3141,N_25611,N_27317);
or UO_3142 (O_3142,N_29874,N_28494);
and UO_3143 (O_3143,N_29612,N_27213);
nor UO_3144 (O_3144,N_28291,N_29045);
xor UO_3145 (O_3145,N_26297,N_26725);
nand UO_3146 (O_3146,N_29135,N_27530);
and UO_3147 (O_3147,N_25090,N_27415);
and UO_3148 (O_3148,N_29383,N_26198);
or UO_3149 (O_3149,N_28743,N_27171);
nand UO_3150 (O_3150,N_25538,N_26323);
nor UO_3151 (O_3151,N_29387,N_28171);
or UO_3152 (O_3152,N_27745,N_28946);
nor UO_3153 (O_3153,N_29470,N_28480);
nor UO_3154 (O_3154,N_26119,N_29651);
nand UO_3155 (O_3155,N_25112,N_29913);
or UO_3156 (O_3156,N_28343,N_25676);
or UO_3157 (O_3157,N_28744,N_25593);
xnor UO_3158 (O_3158,N_28419,N_26392);
xor UO_3159 (O_3159,N_26271,N_26679);
xor UO_3160 (O_3160,N_29184,N_26569);
and UO_3161 (O_3161,N_28082,N_28575);
xnor UO_3162 (O_3162,N_29869,N_25229);
or UO_3163 (O_3163,N_27345,N_27871);
and UO_3164 (O_3164,N_28792,N_26711);
nor UO_3165 (O_3165,N_25140,N_25078);
nand UO_3166 (O_3166,N_27633,N_29989);
nand UO_3167 (O_3167,N_28034,N_25156);
nor UO_3168 (O_3168,N_29039,N_28973);
nand UO_3169 (O_3169,N_27108,N_25855);
or UO_3170 (O_3170,N_25324,N_27140);
nand UO_3171 (O_3171,N_25991,N_27508);
nor UO_3172 (O_3172,N_25917,N_27034);
and UO_3173 (O_3173,N_29769,N_26041);
nor UO_3174 (O_3174,N_27490,N_29701);
nand UO_3175 (O_3175,N_25010,N_25108);
and UO_3176 (O_3176,N_28302,N_27052);
nor UO_3177 (O_3177,N_27082,N_28847);
nor UO_3178 (O_3178,N_26500,N_25982);
or UO_3179 (O_3179,N_29140,N_29128);
nand UO_3180 (O_3180,N_25293,N_26556);
nand UO_3181 (O_3181,N_27176,N_26476);
xor UO_3182 (O_3182,N_27754,N_27830);
or UO_3183 (O_3183,N_27751,N_26785);
xnor UO_3184 (O_3184,N_29841,N_27604);
and UO_3185 (O_3185,N_28953,N_29089);
nand UO_3186 (O_3186,N_29376,N_29923);
xor UO_3187 (O_3187,N_28340,N_27264);
and UO_3188 (O_3188,N_27491,N_25494);
nand UO_3189 (O_3189,N_26385,N_26903);
xnor UO_3190 (O_3190,N_26146,N_28226);
nor UO_3191 (O_3191,N_29691,N_29823);
nand UO_3192 (O_3192,N_26099,N_29697);
xnor UO_3193 (O_3193,N_28157,N_26492);
or UO_3194 (O_3194,N_27750,N_25394);
xnor UO_3195 (O_3195,N_27823,N_29176);
nor UO_3196 (O_3196,N_25354,N_29004);
xor UO_3197 (O_3197,N_29179,N_26324);
xnor UO_3198 (O_3198,N_29527,N_27381);
nor UO_3199 (O_3199,N_25307,N_28625);
xnor UO_3200 (O_3200,N_29689,N_29843);
nor UO_3201 (O_3201,N_26010,N_25387);
or UO_3202 (O_3202,N_26626,N_29618);
and UO_3203 (O_3203,N_28693,N_25931);
nor UO_3204 (O_3204,N_27630,N_25476);
nor UO_3205 (O_3205,N_28265,N_29631);
or UO_3206 (O_3206,N_29632,N_26971);
nand UO_3207 (O_3207,N_27631,N_29629);
nor UO_3208 (O_3208,N_27450,N_28409);
and UO_3209 (O_3209,N_27130,N_25885);
xnor UO_3210 (O_3210,N_25178,N_28959);
and UO_3211 (O_3211,N_27103,N_27798);
nor UO_3212 (O_3212,N_26463,N_25037);
xnor UO_3213 (O_3213,N_29396,N_25126);
and UO_3214 (O_3214,N_27954,N_27192);
and UO_3215 (O_3215,N_26525,N_26002);
nand UO_3216 (O_3216,N_25160,N_29342);
xnor UO_3217 (O_3217,N_26377,N_27850);
and UO_3218 (O_3218,N_28551,N_25441);
and UO_3219 (O_3219,N_28531,N_27096);
and UO_3220 (O_3220,N_26770,N_28279);
xor UO_3221 (O_3221,N_26851,N_27714);
or UO_3222 (O_3222,N_26112,N_27542);
nand UO_3223 (O_3223,N_27674,N_29179);
xor UO_3224 (O_3224,N_27722,N_28520);
and UO_3225 (O_3225,N_29490,N_26673);
or UO_3226 (O_3226,N_26892,N_26987);
xor UO_3227 (O_3227,N_25275,N_25885);
or UO_3228 (O_3228,N_25451,N_29237);
nand UO_3229 (O_3229,N_29370,N_26297);
and UO_3230 (O_3230,N_27849,N_25993);
xor UO_3231 (O_3231,N_28425,N_28082);
xnor UO_3232 (O_3232,N_26087,N_26691);
nand UO_3233 (O_3233,N_28108,N_28695);
and UO_3234 (O_3234,N_27162,N_25329);
and UO_3235 (O_3235,N_27307,N_29133);
nor UO_3236 (O_3236,N_28639,N_25529);
nand UO_3237 (O_3237,N_27480,N_25009);
nor UO_3238 (O_3238,N_29812,N_27446);
or UO_3239 (O_3239,N_27331,N_29235);
nand UO_3240 (O_3240,N_26863,N_27900);
or UO_3241 (O_3241,N_25705,N_28733);
or UO_3242 (O_3242,N_26527,N_27364);
xnor UO_3243 (O_3243,N_28172,N_27697);
xor UO_3244 (O_3244,N_29750,N_28537);
and UO_3245 (O_3245,N_26128,N_27030);
and UO_3246 (O_3246,N_27879,N_25705);
and UO_3247 (O_3247,N_27533,N_28640);
and UO_3248 (O_3248,N_29068,N_25050);
and UO_3249 (O_3249,N_28449,N_29064);
or UO_3250 (O_3250,N_27792,N_28903);
nand UO_3251 (O_3251,N_27775,N_28533);
xor UO_3252 (O_3252,N_29252,N_28405);
and UO_3253 (O_3253,N_27222,N_29248);
xor UO_3254 (O_3254,N_25617,N_25470);
and UO_3255 (O_3255,N_27926,N_28473);
and UO_3256 (O_3256,N_29381,N_25771);
or UO_3257 (O_3257,N_26514,N_25675);
nand UO_3258 (O_3258,N_29532,N_29714);
nor UO_3259 (O_3259,N_27106,N_28562);
or UO_3260 (O_3260,N_26727,N_28181);
nand UO_3261 (O_3261,N_25358,N_27281);
or UO_3262 (O_3262,N_25671,N_29697);
or UO_3263 (O_3263,N_26818,N_26925);
and UO_3264 (O_3264,N_29253,N_29011);
xnor UO_3265 (O_3265,N_27024,N_28556);
nand UO_3266 (O_3266,N_29015,N_25517);
nand UO_3267 (O_3267,N_27617,N_28750);
or UO_3268 (O_3268,N_28283,N_27432);
nor UO_3269 (O_3269,N_28131,N_26041);
or UO_3270 (O_3270,N_27128,N_28765);
and UO_3271 (O_3271,N_26344,N_26602);
nor UO_3272 (O_3272,N_29751,N_29927);
nand UO_3273 (O_3273,N_27066,N_26115);
nor UO_3274 (O_3274,N_26639,N_25483);
or UO_3275 (O_3275,N_27432,N_29960);
and UO_3276 (O_3276,N_26204,N_29390);
xnor UO_3277 (O_3277,N_29100,N_25012);
xnor UO_3278 (O_3278,N_27520,N_26250);
nand UO_3279 (O_3279,N_28097,N_26754);
nor UO_3280 (O_3280,N_27714,N_29350);
nor UO_3281 (O_3281,N_25295,N_28751);
xnor UO_3282 (O_3282,N_25081,N_28996);
nand UO_3283 (O_3283,N_26843,N_27893);
nand UO_3284 (O_3284,N_28284,N_27249);
nand UO_3285 (O_3285,N_29321,N_26444);
nor UO_3286 (O_3286,N_29500,N_29101);
and UO_3287 (O_3287,N_27655,N_26900);
nor UO_3288 (O_3288,N_28737,N_29090);
nor UO_3289 (O_3289,N_27763,N_27508);
nor UO_3290 (O_3290,N_25245,N_26227);
or UO_3291 (O_3291,N_29670,N_29373);
or UO_3292 (O_3292,N_26897,N_25367);
nor UO_3293 (O_3293,N_26595,N_25845);
or UO_3294 (O_3294,N_27572,N_29983);
nor UO_3295 (O_3295,N_26224,N_28684);
nand UO_3296 (O_3296,N_25534,N_26398);
and UO_3297 (O_3297,N_27081,N_26190);
or UO_3298 (O_3298,N_29794,N_28882);
nand UO_3299 (O_3299,N_26591,N_25618);
nor UO_3300 (O_3300,N_28229,N_25876);
xnor UO_3301 (O_3301,N_28220,N_26704);
nor UO_3302 (O_3302,N_29350,N_28045);
or UO_3303 (O_3303,N_25544,N_25727);
xnor UO_3304 (O_3304,N_25072,N_29632);
xnor UO_3305 (O_3305,N_29760,N_29475);
or UO_3306 (O_3306,N_28072,N_28526);
and UO_3307 (O_3307,N_25759,N_27173);
or UO_3308 (O_3308,N_25729,N_26072);
and UO_3309 (O_3309,N_25118,N_26839);
xor UO_3310 (O_3310,N_28734,N_29058);
or UO_3311 (O_3311,N_27524,N_28458);
nor UO_3312 (O_3312,N_26647,N_26596);
nor UO_3313 (O_3313,N_28700,N_27375);
nor UO_3314 (O_3314,N_25033,N_26919);
and UO_3315 (O_3315,N_29422,N_29147);
xnor UO_3316 (O_3316,N_28626,N_26873);
and UO_3317 (O_3317,N_26566,N_25982);
nor UO_3318 (O_3318,N_28533,N_28757);
or UO_3319 (O_3319,N_28213,N_25869);
xnor UO_3320 (O_3320,N_28980,N_27530);
xor UO_3321 (O_3321,N_25936,N_26415);
nand UO_3322 (O_3322,N_25859,N_28781);
xnor UO_3323 (O_3323,N_28334,N_25011);
nand UO_3324 (O_3324,N_29237,N_27993);
nand UO_3325 (O_3325,N_29594,N_29293);
nor UO_3326 (O_3326,N_26141,N_26150);
nor UO_3327 (O_3327,N_29695,N_28937);
xor UO_3328 (O_3328,N_28003,N_29300);
and UO_3329 (O_3329,N_25217,N_29665);
nor UO_3330 (O_3330,N_25699,N_26930);
nand UO_3331 (O_3331,N_28507,N_27524);
nor UO_3332 (O_3332,N_28878,N_26777);
nor UO_3333 (O_3333,N_26430,N_28353);
and UO_3334 (O_3334,N_28350,N_26395);
nor UO_3335 (O_3335,N_25237,N_28523);
nor UO_3336 (O_3336,N_28027,N_25969);
nor UO_3337 (O_3337,N_29570,N_26955);
or UO_3338 (O_3338,N_25004,N_27520);
nor UO_3339 (O_3339,N_28872,N_25877);
xor UO_3340 (O_3340,N_27959,N_27246);
nand UO_3341 (O_3341,N_29252,N_28276);
nor UO_3342 (O_3342,N_25094,N_28127);
nand UO_3343 (O_3343,N_26307,N_27061);
xor UO_3344 (O_3344,N_28008,N_25954);
nand UO_3345 (O_3345,N_29722,N_29101);
xnor UO_3346 (O_3346,N_27149,N_29134);
or UO_3347 (O_3347,N_26209,N_29506);
or UO_3348 (O_3348,N_27008,N_27721);
nor UO_3349 (O_3349,N_29087,N_26943);
and UO_3350 (O_3350,N_26434,N_27041);
nor UO_3351 (O_3351,N_25717,N_28469);
nor UO_3352 (O_3352,N_26018,N_28076);
xor UO_3353 (O_3353,N_29079,N_28167);
nor UO_3354 (O_3354,N_26223,N_29711);
xor UO_3355 (O_3355,N_27111,N_27829);
or UO_3356 (O_3356,N_25839,N_27010);
and UO_3357 (O_3357,N_29254,N_28763);
nand UO_3358 (O_3358,N_26126,N_28842);
nand UO_3359 (O_3359,N_25026,N_28235);
and UO_3360 (O_3360,N_25395,N_28841);
nand UO_3361 (O_3361,N_28770,N_26155);
or UO_3362 (O_3362,N_25203,N_29231);
nand UO_3363 (O_3363,N_25002,N_29317);
or UO_3364 (O_3364,N_27632,N_26388);
and UO_3365 (O_3365,N_28677,N_28842);
nand UO_3366 (O_3366,N_26678,N_27611);
or UO_3367 (O_3367,N_28545,N_28424);
nand UO_3368 (O_3368,N_27695,N_26180);
and UO_3369 (O_3369,N_26120,N_26816);
and UO_3370 (O_3370,N_28484,N_28345);
and UO_3371 (O_3371,N_25644,N_25013);
or UO_3372 (O_3372,N_28708,N_29605);
or UO_3373 (O_3373,N_26629,N_28504);
or UO_3374 (O_3374,N_28202,N_25349);
xor UO_3375 (O_3375,N_26173,N_29309);
and UO_3376 (O_3376,N_29893,N_27247);
nand UO_3377 (O_3377,N_25039,N_26907);
and UO_3378 (O_3378,N_29728,N_25719);
xor UO_3379 (O_3379,N_29111,N_27106);
or UO_3380 (O_3380,N_29921,N_25092);
or UO_3381 (O_3381,N_25706,N_25802);
nor UO_3382 (O_3382,N_26842,N_25333);
nor UO_3383 (O_3383,N_25766,N_29837);
nor UO_3384 (O_3384,N_25059,N_27080);
nand UO_3385 (O_3385,N_26369,N_29686);
nand UO_3386 (O_3386,N_25323,N_28183);
nor UO_3387 (O_3387,N_27081,N_25854);
xnor UO_3388 (O_3388,N_28760,N_27622);
and UO_3389 (O_3389,N_29442,N_29701);
xnor UO_3390 (O_3390,N_25304,N_29686);
and UO_3391 (O_3391,N_26866,N_27864);
nand UO_3392 (O_3392,N_29813,N_28581);
and UO_3393 (O_3393,N_26431,N_25002);
nand UO_3394 (O_3394,N_27852,N_25687);
and UO_3395 (O_3395,N_29279,N_27132);
xor UO_3396 (O_3396,N_26369,N_25695);
nand UO_3397 (O_3397,N_25691,N_28634);
or UO_3398 (O_3398,N_28996,N_27999);
and UO_3399 (O_3399,N_27302,N_28630);
nand UO_3400 (O_3400,N_27039,N_26276);
xnor UO_3401 (O_3401,N_27950,N_29449);
nand UO_3402 (O_3402,N_26266,N_28240);
nand UO_3403 (O_3403,N_29540,N_29079);
nor UO_3404 (O_3404,N_27537,N_29666);
xnor UO_3405 (O_3405,N_25355,N_25754);
or UO_3406 (O_3406,N_25197,N_29971);
xnor UO_3407 (O_3407,N_25818,N_27759);
and UO_3408 (O_3408,N_27980,N_28952);
and UO_3409 (O_3409,N_27716,N_25536);
or UO_3410 (O_3410,N_27463,N_25097);
xnor UO_3411 (O_3411,N_27013,N_27236);
xor UO_3412 (O_3412,N_27613,N_29615);
or UO_3413 (O_3413,N_25732,N_29520);
or UO_3414 (O_3414,N_29669,N_28174);
nand UO_3415 (O_3415,N_28492,N_27431);
nand UO_3416 (O_3416,N_27952,N_25197);
nor UO_3417 (O_3417,N_27821,N_26405);
nand UO_3418 (O_3418,N_25474,N_25417);
nor UO_3419 (O_3419,N_27707,N_28358);
or UO_3420 (O_3420,N_27621,N_29306);
nand UO_3421 (O_3421,N_26812,N_25987);
nor UO_3422 (O_3422,N_26509,N_27910);
xor UO_3423 (O_3423,N_28087,N_29376);
and UO_3424 (O_3424,N_26097,N_25041);
or UO_3425 (O_3425,N_29431,N_27665);
nor UO_3426 (O_3426,N_26144,N_26555);
nor UO_3427 (O_3427,N_28898,N_29130);
nand UO_3428 (O_3428,N_28337,N_29752);
or UO_3429 (O_3429,N_29940,N_29599);
nand UO_3430 (O_3430,N_28581,N_29382);
nor UO_3431 (O_3431,N_28997,N_29150);
or UO_3432 (O_3432,N_28480,N_27760);
nor UO_3433 (O_3433,N_25820,N_26191);
nand UO_3434 (O_3434,N_28897,N_28713);
nor UO_3435 (O_3435,N_25991,N_29386);
and UO_3436 (O_3436,N_28431,N_27754);
or UO_3437 (O_3437,N_27817,N_29563);
or UO_3438 (O_3438,N_27790,N_25370);
nor UO_3439 (O_3439,N_25444,N_25681);
nand UO_3440 (O_3440,N_28350,N_26457);
and UO_3441 (O_3441,N_25083,N_26128);
and UO_3442 (O_3442,N_26980,N_28607);
nand UO_3443 (O_3443,N_25961,N_26224);
nor UO_3444 (O_3444,N_26545,N_27276);
xnor UO_3445 (O_3445,N_28653,N_25488);
nand UO_3446 (O_3446,N_29959,N_27235);
xnor UO_3447 (O_3447,N_28108,N_25175);
nor UO_3448 (O_3448,N_28686,N_28765);
nand UO_3449 (O_3449,N_25772,N_27165);
xor UO_3450 (O_3450,N_26275,N_28574);
nor UO_3451 (O_3451,N_25705,N_27635);
nor UO_3452 (O_3452,N_25735,N_26927);
and UO_3453 (O_3453,N_28148,N_29861);
and UO_3454 (O_3454,N_27550,N_25113);
nand UO_3455 (O_3455,N_29947,N_28656);
or UO_3456 (O_3456,N_28480,N_25939);
or UO_3457 (O_3457,N_28200,N_27791);
xnor UO_3458 (O_3458,N_26951,N_27113);
nor UO_3459 (O_3459,N_29850,N_29984);
xor UO_3460 (O_3460,N_25637,N_29157);
and UO_3461 (O_3461,N_27964,N_29580);
nand UO_3462 (O_3462,N_27515,N_26930);
xor UO_3463 (O_3463,N_27966,N_27765);
and UO_3464 (O_3464,N_27143,N_26919);
xnor UO_3465 (O_3465,N_28268,N_25918);
nand UO_3466 (O_3466,N_29087,N_27376);
nor UO_3467 (O_3467,N_29240,N_26396);
and UO_3468 (O_3468,N_29095,N_28044);
and UO_3469 (O_3469,N_29572,N_27668);
xor UO_3470 (O_3470,N_27277,N_26540);
xor UO_3471 (O_3471,N_29926,N_27219);
xnor UO_3472 (O_3472,N_29956,N_27320);
nand UO_3473 (O_3473,N_28761,N_27310);
and UO_3474 (O_3474,N_28416,N_25330);
nand UO_3475 (O_3475,N_26853,N_27102);
nor UO_3476 (O_3476,N_29885,N_26231);
xor UO_3477 (O_3477,N_29092,N_27323);
or UO_3478 (O_3478,N_25898,N_25407);
nor UO_3479 (O_3479,N_27807,N_28428);
nor UO_3480 (O_3480,N_25782,N_26478);
and UO_3481 (O_3481,N_26259,N_25921);
or UO_3482 (O_3482,N_28774,N_27463);
nand UO_3483 (O_3483,N_28844,N_28792);
xnor UO_3484 (O_3484,N_26620,N_28712);
or UO_3485 (O_3485,N_29203,N_25462);
xnor UO_3486 (O_3486,N_26524,N_26126);
xnor UO_3487 (O_3487,N_26125,N_27619);
or UO_3488 (O_3488,N_29263,N_28606);
xnor UO_3489 (O_3489,N_27118,N_28770);
nand UO_3490 (O_3490,N_26484,N_25259);
nand UO_3491 (O_3491,N_29064,N_29275);
nor UO_3492 (O_3492,N_28366,N_29611);
nand UO_3493 (O_3493,N_27898,N_25170);
xnor UO_3494 (O_3494,N_25027,N_29388);
xnor UO_3495 (O_3495,N_27857,N_27315);
nand UO_3496 (O_3496,N_28215,N_27409);
and UO_3497 (O_3497,N_27918,N_27498);
xor UO_3498 (O_3498,N_26399,N_26276);
nor UO_3499 (O_3499,N_25496,N_25894);
endmodule