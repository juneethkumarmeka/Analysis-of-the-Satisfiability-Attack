module basic_2500_25000_3000_40_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_202,In_782);
nor U1 (N_1,In_1840,In_2040);
nor U2 (N_2,In_653,In_1302);
nand U3 (N_3,In_961,In_628);
or U4 (N_4,In_276,In_150);
or U5 (N_5,In_742,In_1642);
nand U6 (N_6,In_1745,In_1783);
nor U7 (N_7,In_1925,In_2062);
nor U8 (N_8,In_915,In_959);
xnor U9 (N_9,In_1993,In_113);
and U10 (N_10,In_359,In_2270);
nand U11 (N_11,In_2000,In_478);
nor U12 (N_12,In_428,In_691);
nand U13 (N_13,In_123,In_1702);
or U14 (N_14,In_2106,In_442);
nand U15 (N_15,In_1777,In_284);
or U16 (N_16,In_208,In_258);
or U17 (N_17,In_1493,In_787);
nand U18 (N_18,In_1873,In_1359);
nor U19 (N_19,In_764,In_1661);
nand U20 (N_20,In_2412,In_1435);
xnor U21 (N_21,In_1985,In_605);
nand U22 (N_22,In_2170,In_2260);
xor U23 (N_23,In_2288,In_1259);
and U24 (N_24,In_55,In_2207);
xor U25 (N_25,In_1608,In_1081);
and U26 (N_26,In_1185,In_1257);
xor U27 (N_27,In_900,In_2131);
nand U28 (N_28,In_281,In_802);
or U29 (N_29,In_1950,In_1013);
and U30 (N_30,In_2026,In_1271);
nor U31 (N_31,In_1789,In_1674);
nor U32 (N_32,In_2182,In_907);
or U33 (N_33,In_1947,In_749);
and U34 (N_34,In_1656,In_806);
and U35 (N_35,In_2033,In_1072);
nand U36 (N_36,In_917,In_77);
nand U37 (N_37,In_332,In_2343);
nand U38 (N_38,In_2462,In_1550);
and U39 (N_39,In_2328,In_1500);
or U40 (N_40,In_680,In_761);
nand U41 (N_41,In_325,In_257);
or U42 (N_42,In_1148,In_1347);
and U43 (N_43,In_186,In_2410);
nand U44 (N_44,In_4,In_972);
nand U45 (N_45,In_304,In_1971);
or U46 (N_46,In_1209,In_1831);
nor U47 (N_47,In_2169,In_738);
or U48 (N_48,In_2161,In_1235);
and U49 (N_49,In_760,In_786);
or U50 (N_50,In_33,In_1590);
xnor U51 (N_51,In_2437,In_1996);
and U52 (N_52,In_1844,In_1002);
or U53 (N_53,In_647,In_448);
or U54 (N_54,In_25,In_389);
nor U55 (N_55,In_937,In_1427);
and U56 (N_56,In_1677,In_1887);
nor U57 (N_57,In_1513,In_1516);
xor U58 (N_58,In_1059,In_37);
nand U59 (N_59,In_328,In_918);
nand U60 (N_60,In_2333,In_1834);
and U61 (N_61,In_930,In_2396);
nand U62 (N_62,In_388,In_600);
nand U63 (N_63,In_1801,In_661);
or U64 (N_64,In_1439,In_450);
and U65 (N_65,In_356,In_1680);
or U66 (N_66,In_1956,In_336);
and U67 (N_67,In_2360,In_461);
or U68 (N_68,In_1217,In_2453);
xnor U69 (N_69,In_558,In_1450);
nor U70 (N_70,In_125,In_97);
or U71 (N_71,In_1662,In_41);
nor U72 (N_72,In_2355,In_866);
nor U73 (N_73,In_1463,In_1653);
nor U74 (N_74,In_1068,In_1093);
or U75 (N_75,In_1491,In_2481);
and U76 (N_76,In_1157,In_1260);
nor U77 (N_77,In_527,In_1420);
and U78 (N_78,In_1647,In_1248);
nor U79 (N_79,In_1095,In_1096);
nand U80 (N_80,In_1116,In_1042);
nand U81 (N_81,In_2084,In_2168);
and U82 (N_82,In_855,In_1696);
or U83 (N_83,In_403,In_429);
and U84 (N_84,In_1903,In_2198);
and U85 (N_85,In_1876,In_1180);
nand U86 (N_86,In_1786,In_1268);
and U87 (N_87,In_1543,In_2374);
nor U88 (N_88,In_1141,In_2175);
or U89 (N_89,In_968,In_546);
or U90 (N_90,In_2022,In_1365);
xor U91 (N_91,In_2031,In_1153);
and U92 (N_92,In_2467,In_1699);
or U93 (N_93,In_220,In_744);
or U94 (N_94,In_503,In_91);
nor U95 (N_95,In_1430,In_1142);
nand U96 (N_96,In_620,In_921);
or U97 (N_97,In_1713,In_22);
nor U98 (N_98,In_1084,In_550);
or U99 (N_99,In_2457,In_920);
nand U100 (N_100,In_0,In_626);
or U101 (N_101,In_2298,In_1555);
nor U102 (N_102,In_165,In_121);
nand U103 (N_103,In_1426,In_603);
nand U104 (N_104,In_1117,In_166);
nand U105 (N_105,In_616,In_801);
xnor U106 (N_106,In_705,In_510);
or U107 (N_107,In_2116,In_939);
or U108 (N_108,In_583,In_47);
and U109 (N_109,In_140,In_1459);
nor U110 (N_110,In_272,In_1310);
nand U111 (N_111,In_94,In_2471);
nor U112 (N_112,In_979,In_1571);
and U113 (N_113,In_2302,In_110);
or U114 (N_114,In_2266,In_1232);
and U115 (N_115,In_1867,In_1058);
nor U116 (N_116,In_805,In_1584);
nor U117 (N_117,In_2127,In_557);
nand U118 (N_118,In_247,In_631);
nand U119 (N_119,In_1949,In_1175);
or U120 (N_120,In_441,In_864);
nor U121 (N_121,In_981,In_739);
and U122 (N_122,In_1221,In_2265);
or U123 (N_123,In_1685,In_658);
and U124 (N_124,In_142,In_2217);
or U125 (N_125,In_2054,In_544);
and U126 (N_126,In_1418,In_1075);
nand U127 (N_127,In_1955,In_1007);
nand U128 (N_128,In_1936,In_1613);
xnor U129 (N_129,In_1684,In_2006);
or U130 (N_130,In_2386,In_2129);
or U131 (N_131,In_76,In_783);
nand U132 (N_132,In_30,In_886);
nor U133 (N_133,In_2398,In_2101);
xor U134 (N_134,In_1901,In_214);
nand U135 (N_135,In_678,In_2494);
and U136 (N_136,In_2289,In_858);
or U137 (N_137,In_809,In_2269);
nor U138 (N_138,In_1795,In_624);
or U139 (N_139,In_2388,In_2189);
nor U140 (N_140,In_596,In_1462);
xnor U141 (N_141,In_241,In_1546);
nand U142 (N_142,In_1962,In_1055);
nand U143 (N_143,In_2153,In_1186);
or U144 (N_144,In_351,In_913);
or U145 (N_145,In_1863,In_435);
and U146 (N_146,In_1630,In_66);
nand U147 (N_147,In_1758,In_521);
nand U148 (N_148,In_2475,In_529);
or U149 (N_149,In_2145,In_1110);
or U150 (N_150,In_242,In_992);
or U151 (N_151,In_2090,In_1527);
nand U152 (N_152,In_704,In_1510);
nand U153 (N_153,In_1234,In_1780);
nor U154 (N_154,In_1978,In_2316);
and U155 (N_155,In_372,In_2183);
and U156 (N_156,In_1280,In_201);
nand U157 (N_157,In_1165,In_692);
nand U158 (N_158,In_2213,In_1849);
nand U159 (N_159,In_1161,In_2144);
and U160 (N_160,In_794,In_563);
or U161 (N_161,In_2309,In_836);
nand U162 (N_162,In_1779,In_2258);
nor U163 (N_163,In_2439,In_2402);
and U164 (N_164,In_2195,In_1698);
and U165 (N_165,In_1963,In_2185);
nand U166 (N_166,In_1670,In_236);
xor U167 (N_167,In_1385,In_1600);
nor U168 (N_168,In_79,In_1253);
nand U169 (N_169,In_2294,In_158);
nor U170 (N_170,In_1835,In_1124);
nand U171 (N_171,In_2291,In_1891);
nor U172 (N_172,In_2435,In_634);
and U173 (N_173,In_151,In_2202);
and U174 (N_174,In_177,In_1397);
or U175 (N_175,In_1968,In_2034);
or U176 (N_176,In_2177,In_1335);
xnor U177 (N_177,In_433,In_1281);
nor U178 (N_178,In_1554,In_1298);
nor U179 (N_179,In_537,In_1511);
and U180 (N_180,In_873,In_686);
nand U181 (N_181,In_100,In_1746);
xor U182 (N_182,In_1039,In_2201);
or U183 (N_183,In_536,In_2488);
xnor U184 (N_184,In_1718,In_784);
or U185 (N_185,In_1370,In_2262);
nand U186 (N_186,In_1118,In_2391);
and U187 (N_187,In_101,In_538);
or U188 (N_188,In_2303,In_339);
xnor U189 (N_189,In_2357,In_384);
nor U190 (N_190,In_714,In_460);
or U191 (N_191,In_1899,In_133);
and U192 (N_192,In_2070,In_1415);
nand U193 (N_193,In_1393,In_1318);
nand U194 (N_194,In_1731,In_103);
or U195 (N_195,In_1877,In_2468);
or U196 (N_196,In_1297,In_846);
nor U197 (N_197,In_1448,In_2419);
and U198 (N_198,In_2075,In_951);
nand U199 (N_199,In_1791,In_1805);
nor U200 (N_200,In_530,In_769);
or U201 (N_201,In_1040,In_2397);
or U202 (N_202,In_1063,In_361);
xnor U203 (N_203,In_927,In_1275);
nor U204 (N_204,In_93,In_1885);
nand U205 (N_205,In_1562,In_2060);
and U206 (N_206,In_607,In_2134);
and U207 (N_207,In_643,In_1255);
nand U208 (N_208,In_1005,In_1595);
nor U209 (N_209,In_1011,In_561);
and U210 (N_210,In_908,In_497);
nand U211 (N_211,In_1472,In_1770);
nand U212 (N_212,In_1808,In_1614);
or U213 (N_213,In_1473,In_698);
nand U214 (N_214,In_2267,In_509);
nor U215 (N_215,In_1464,In_2059);
nor U216 (N_216,In_2130,In_932);
nand U217 (N_217,In_1803,In_10);
nand U218 (N_218,In_1693,In_1576);
nor U219 (N_219,In_49,In_40);
or U220 (N_220,In_1788,In_1105);
nor U221 (N_221,In_1998,In_2152);
nor U222 (N_222,In_2451,In_1727);
nand U223 (N_223,In_1277,In_61);
and U224 (N_224,In_2231,In_1665);
and U225 (N_225,In_820,In_1889);
nand U226 (N_226,In_516,In_2404);
nand U227 (N_227,In_1062,In_1200);
and U228 (N_228,In_1482,In_1193);
or U229 (N_229,In_1089,In_482);
or U230 (N_230,In_2256,In_819);
nor U231 (N_231,In_925,In_421);
or U232 (N_232,In_762,In_1012);
and U233 (N_233,In_947,In_2124);
nor U234 (N_234,In_1874,In_31);
or U235 (N_235,In_2214,In_1181);
xor U236 (N_236,In_48,In_1765);
nor U237 (N_237,In_2301,In_953);
nor U238 (N_238,In_615,In_1577);
nor U239 (N_239,In_2018,In_941);
and U240 (N_240,In_1194,In_1961);
nand U241 (N_241,In_1037,In_1994);
nand U242 (N_242,In_1402,In_1797);
nor U243 (N_243,In_1564,In_1091);
and U244 (N_244,In_1502,In_1158);
nor U245 (N_245,In_171,In_206);
or U246 (N_246,In_173,In_976);
nor U247 (N_247,In_1732,In_2465);
nor U248 (N_248,In_2380,In_713);
xnor U249 (N_249,In_386,In_1659);
xor U250 (N_250,In_1669,In_969);
nand U251 (N_251,In_1563,In_1658);
nand U252 (N_252,In_513,In_1348);
nor U253 (N_253,In_552,In_574);
and U254 (N_254,In_2208,In_883);
or U255 (N_255,In_2341,In_1568);
and U256 (N_256,In_526,In_598);
or U257 (N_257,In_1536,In_68);
nand U258 (N_258,In_730,In_2227);
nand U259 (N_259,In_38,In_973);
and U260 (N_260,In_1150,In_2035);
nor U261 (N_261,In_1673,In_2354);
nor U262 (N_262,In_1289,In_19);
nand U263 (N_263,In_70,In_2276);
nand U264 (N_264,In_1060,In_777);
and U265 (N_265,In_2192,In_85);
or U266 (N_266,In_1616,In_2320);
or U267 (N_267,In_994,In_190);
nor U268 (N_268,In_639,In_444);
and U269 (N_269,In_1167,In_2491);
and U270 (N_270,In_619,In_1541);
nor U271 (N_271,In_2204,In_793);
or U272 (N_272,In_1958,In_1846);
and U273 (N_273,In_2017,In_1220);
nand U274 (N_274,In_1640,In_392);
or U275 (N_275,In_1131,In_840);
xor U276 (N_276,In_344,In_1822);
or U277 (N_277,In_96,In_1090);
nand U278 (N_278,In_492,In_1977);
nand U279 (N_279,In_697,In_104);
nand U280 (N_280,In_321,In_995);
or U281 (N_281,In_2155,In_455);
nor U282 (N_282,In_660,In_899);
and U283 (N_283,In_2331,In_248);
nand U284 (N_284,In_2203,In_1242);
nand U285 (N_285,In_807,In_709);
or U286 (N_286,In_205,In_1441);
or U287 (N_287,In_1990,In_423);
and U288 (N_288,In_2064,In_1497);
or U289 (N_289,In_1315,In_823);
nand U290 (N_290,In_545,In_571);
nand U291 (N_291,In_1306,In_445);
or U292 (N_292,In_716,In_1114);
nand U293 (N_293,In_1303,In_295);
and U294 (N_294,In_1355,In_1307);
nand U295 (N_295,In_1195,In_1300);
or U296 (N_296,In_2012,In_611);
or U297 (N_297,In_581,In_1847);
or U298 (N_298,In_145,In_1811);
xnor U299 (N_299,In_185,In_632);
nor U300 (N_300,In_1083,In_1778);
nand U301 (N_301,In_1319,In_1556);
nand U302 (N_302,In_724,In_81);
and U303 (N_303,In_7,In_2326);
nor U304 (N_304,In_139,In_1351);
or U305 (N_305,In_2339,In_115);
nor U306 (N_306,In_2048,In_2080);
nand U307 (N_307,In_2077,In_1744);
xnor U308 (N_308,In_1076,In_2240);
or U309 (N_309,In_1773,In_1061);
nand U310 (N_310,In_1969,In_1440);
nor U311 (N_311,In_2337,In_1810);
or U312 (N_312,In_244,In_2181);
nand U313 (N_313,In_193,In_153);
nand U314 (N_314,In_2098,In_1241);
nand U315 (N_315,In_904,In_531);
nand U316 (N_316,In_1833,In_207);
nand U317 (N_317,In_876,In_826);
or U318 (N_318,In_1905,In_888);
nand U319 (N_319,In_610,In_1612);
nor U320 (N_320,In_1292,In_1982);
nand U321 (N_321,In_309,In_1941);
nor U322 (N_322,In_837,In_1445);
and U323 (N_323,In_743,In_1276);
nor U324 (N_324,In_1154,In_67);
nand U325 (N_325,In_2236,In_1757);
and U326 (N_326,In_1787,In_288);
or U327 (N_327,In_1841,In_1585);
or U328 (N_328,In_1092,In_1251);
or U329 (N_329,In_748,In_320);
and U330 (N_330,In_1373,In_180);
nor U331 (N_331,In_2009,In_2366);
or U332 (N_332,In_1760,In_1624);
and U333 (N_333,In_2450,In_609);
nor U334 (N_334,In_128,In_737);
xor U335 (N_335,In_2078,In_938);
xor U336 (N_336,In_656,In_533);
nor U337 (N_337,In_1311,In_374);
xor U338 (N_338,In_1528,In_948);
and U339 (N_339,In_2358,In_2187);
and U340 (N_340,In_825,In_1660);
or U341 (N_341,In_2283,In_1937);
nor U342 (N_342,In_798,In_418);
nor U343 (N_343,In_725,In_1073);
or U344 (N_344,In_1654,In_65);
and U345 (N_345,In_52,In_1631);
and U346 (N_346,In_494,In_2164);
xor U347 (N_347,In_168,In_1363);
nor U348 (N_348,In_1304,In_446);
or U349 (N_349,In_1372,In_745);
nor U350 (N_350,In_2307,In_2497);
nand U351 (N_351,In_2495,In_1987);
xor U352 (N_352,In_2212,In_1605);
and U353 (N_353,In_221,In_1160);
nor U354 (N_354,In_114,In_1162);
nor U355 (N_355,In_1552,In_2125);
nand U356 (N_356,In_1646,In_931);
or U357 (N_357,In_780,In_11);
or U358 (N_358,In_1471,In_1479);
xnor U359 (N_359,In_1223,In_326);
and U360 (N_360,In_282,In_1572);
and U361 (N_361,In_1676,In_1171);
nor U362 (N_362,In_2209,In_1717);
or U363 (N_363,In_2329,In_519);
nand U364 (N_364,In_1320,In_850);
or U365 (N_365,In_532,In_1458);
and U366 (N_366,In_1768,In_256);
nand U367 (N_367,In_2010,In_2032);
nor U368 (N_368,In_375,In_1883);
nand U369 (N_369,In_2378,In_2186);
and U370 (N_370,In_2338,In_1628);
nor U371 (N_371,In_2206,In_1829);
xor U372 (N_372,In_129,In_914);
and U373 (N_373,In_1030,In_302);
nor U374 (N_374,In_2193,In_2150);
and U375 (N_375,In_1299,In_1679);
or U376 (N_376,In_1112,In_756);
nor U377 (N_377,In_1703,In_1398);
nor U378 (N_378,In_778,In_928);
xnor U379 (N_379,In_2139,In_1858);
nand U380 (N_380,In_813,In_2381);
or U381 (N_381,In_1414,In_2489);
nor U382 (N_382,In_75,In_2091);
nand U383 (N_383,In_1137,In_414);
xnor U384 (N_384,In_694,In_1125);
nor U385 (N_385,In_1918,In_1378);
or U386 (N_386,In_175,In_1444);
nand U387 (N_387,In_222,In_1409);
nor U388 (N_388,In_1864,In_1535);
or U389 (N_389,In_617,In_240);
and U390 (N_390,In_174,In_2041);
and U391 (N_391,In_1317,In_1524);
and U392 (N_392,In_1191,In_2093);
or U393 (N_393,In_1443,In_881);
nor U394 (N_394,In_63,In_2238);
nand U395 (N_395,In_2245,In_132);
or U396 (N_396,In_520,In_1845);
and U397 (N_397,In_1050,In_614);
and U398 (N_398,In_1617,In_1515);
nand U399 (N_399,In_2321,In_2418);
nor U400 (N_400,In_822,In_1328);
nor U401 (N_401,In_1029,In_874);
and U402 (N_402,In_269,In_548);
nand U403 (N_403,In_1283,In_1484);
nand U404 (N_404,In_323,In_483);
nor U405 (N_405,In_898,In_997);
nand U406 (N_406,In_1145,In_861);
xor U407 (N_407,In_1880,In_1591);
xor U408 (N_408,In_499,In_728);
nor U409 (N_409,In_112,In_1270);
and U410 (N_410,In_2484,In_568);
and U411 (N_411,In_1044,In_1923);
and U412 (N_412,In_810,In_667);
nor U413 (N_413,In_2036,In_1751);
nand U414 (N_414,In_465,In_508);
or U415 (N_415,In_1868,In_2389);
nand U416 (N_416,In_1329,In_2230);
xnor U417 (N_417,In_355,In_1313);
and U418 (N_418,In_573,In_1336);
nor U419 (N_419,In_365,In_766);
or U420 (N_420,In_51,In_2021);
nand U421 (N_421,In_2233,In_1570);
and U422 (N_422,In_679,In_1399);
and U423 (N_423,In_715,In_1231);
nand U424 (N_424,In_1566,In_905);
nand U425 (N_425,In_602,In_135);
or U426 (N_426,In_923,In_2426);
nand U427 (N_427,In_1417,In_747);
and U428 (N_428,In_1166,In_1279);
nor U429 (N_429,In_229,In_331);
and U430 (N_430,In_566,In_1331);
nor U431 (N_431,In_1853,In_1294);
nor U432 (N_432,In_2016,In_1774);
or U433 (N_433,In_343,In_1875);
nor U434 (N_434,In_595,In_14);
and U435 (N_435,In_795,In_2007);
and U436 (N_436,In_46,In_2443);
nor U437 (N_437,In_1939,In_181);
nor U438 (N_438,In_1466,In_1859);
or U439 (N_439,In_2382,In_2414);
nand U440 (N_440,In_172,In_791);
or U441 (N_441,In_916,In_2440);
and U442 (N_442,In_26,In_2349);
or U443 (N_443,In_456,In_2157);
nor U444 (N_444,In_498,In_2332);
nand U445 (N_445,In_991,In_1775);
or U446 (N_446,In_690,In_1043);
xnor U447 (N_447,In_1496,In_253);
and U448 (N_448,In_1610,In_5);
or U449 (N_449,In_1986,In_470);
and U450 (N_450,In_99,In_1999);
nand U451 (N_451,In_107,In_922);
nor U452 (N_452,In_223,In_2030);
nor U453 (N_453,In_1130,In_1664);
nand U454 (N_454,In_2194,In_1052);
nor U455 (N_455,In_1721,In_1032);
nor U456 (N_456,In_2472,In_753);
nand U457 (N_457,In_597,In_2478);
nor U458 (N_458,In_329,In_1477);
and U459 (N_459,In_1225,In_2120);
nand U460 (N_460,In_32,In_1263);
xor U461 (N_461,In_1755,In_1433);
nor U462 (N_462,In_260,In_27);
nand U463 (N_463,In_940,In_1377);
or U464 (N_464,In_891,In_261);
and U465 (N_465,In_949,In_1269);
and U466 (N_466,In_831,In_1369);
or U467 (N_467,In_872,In_1817);
nand U468 (N_468,In_682,In_234);
nor U469 (N_469,In_466,In_2137);
nor U470 (N_470,In_757,In_522);
or U471 (N_471,In_1588,In_182);
and U472 (N_472,In_431,In_2191);
nand U473 (N_473,In_496,In_2352);
and U474 (N_474,In_2135,In_1057);
xor U475 (N_475,In_1431,In_1386);
nand U476 (N_476,In_224,In_1470);
or U477 (N_477,In_1520,In_2148);
and U478 (N_478,In_2087,In_2411);
and U479 (N_479,In_1632,In_2460);
xor U480 (N_480,In_1682,In_2480);
and U481 (N_481,In_1467,In_1623);
nand U482 (N_482,In_1284,In_2133);
nor U483 (N_483,In_1113,In_146);
nor U484 (N_484,In_670,In_397);
nand U485 (N_485,In_2222,In_334);
and U486 (N_486,In_2049,In_946);
and U487 (N_487,In_1785,In_426);
nor U488 (N_488,In_842,In_1813);
and U489 (N_489,In_870,In_1547);
or U490 (N_490,In_1565,In_2401);
nor U491 (N_491,In_1362,In_227);
nand U492 (N_492,In_1933,In_2141);
nor U493 (N_493,In_477,In_1667);
and U494 (N_494,In_975,In_382);
or U495 (N_495,In_1338,In_1379);
xor U496 (N_496,In_369,In_985);
nor U497 (N_497,In_2094,In_771);
nand U498 (N_498,In_2052,In_188);
nor U499 (N_499,In_983,In_342);
xnor U500 (N_500,In_1014,In_1210);
or U501 (N_501,In_277,In_1697);
and U502 (N_502,In_1047,In_1724);
or U503 (N_503,In_1020,In_911);
and U504 (N_504,In_835,In_1951);
or U505 (N_505,In_9,In_1080);
nor U506 (N_506,In_1395,In_1038);
and U507 (N_507,In_1079,In_1004);
nor U508 (N_508,In_542,In_2002);
nor U509 (N_509,In_138,In_1465);
and U510 (N_510,In_999,In_966);
and U511 (N_511,In_452,In_960);
and U512 (N_512,In_1750,In_353);
or U513 (N_513,In_1715,In_1487);
or U514 (N_514,In_84,In_1266);
and U515 (N_515,In_2243,In_912);
nand U516 (N_516,In_1689,In_347);
xnor U517 (N_517,In_1690,In_1273);
or U518 (N_518,In_2250,In_849);
or U519 (N_519,In_1326,In_1442);
nor U520 (N_520,In_539,In_1558);
or U521 (N_521,In_268,In_729);
nand U522 (N_522,In_512,In_1321);
or U523 (N_523,In_187,In_1957);
and U524 (N_524,In_310,In_606);
xor U525 (N_525,In_1368,In_1754);
and U526 (N_526,In_2039,In_45);
nand U527 (N_527,In_1519,In_1506);
or U528 (N_528,In_1827,In_1018);
and U529 (N_529,In_1578,In_1262);
nor U530 (N_530,In_1135,In_1367);
or U531 (N_531,In_540,In_889);
or U532 (N_532,In_120,In_638);
nor U533 (N_533,In_480,In_2028);
nand U534 (N_534,In_218,In_1837);
and U535 (N_535,In_1389,In_651);
nand U536 (N_536,In_1371,In_1719);
nand U537 (N_537,In_534,In_42);
nor U538 (N_538,In_853,In_1078);
nor U539 (N_539,In_1026,In_773);
or U540 (N_540,In_1192,In_1776);
nor U541 (N_541,In_2272,In_2455);
nand U542 (N_542,In_2074,In_1278);
nand U543 (N_543,In_2261,In_567);
xor U544 (N_544,In_238,In_2459);
and U545 (N_545,In_1622,In_1478);
nor U546 (N_546,In_2104,In_1400);
or U547 (N_547,In_28,In_1169);
xor U548 (N_548,In_572,In_722);
or U549 (N_549,In_2477,In_2197);
and U550 (N_550,In_2050,In_2372);
nand U551 (N_551,In_1122,In_1187);
or U552 (N_552,In_1295,In_2284);
nor U553 (N_553,In_1384,In_488);
or U554 (N_554,In_60,In_83);
nor U555 (N_555,In_1759,In_2038);
nor U556 (N_556,In_1587,In_1504);
and U557 (N_557,In_1207,In_865);
and U558 (N_558,In_1753,In_1976);
nand U559 (N_559,In_841,In_350);
nor U560 (N_560,In_126,In_1107);
and U561 (N_561,In_1529,In_349);
nor U562 (N_562,In_902,In_1657);
and U563 (N_563,In_950,In_394);
xnor U564 (N_564,In_2271,In_1598);
or U565 (N_565,In_1388,In_2115);
or U566 (N_566,In_645,In_2051);
and U567 (N_567,In_1354,In_514);
nand U568 (N_568,In_385,In_1729);
and U569 (N_569,In_1940,In_462);
nand U570 (N_570,In_1922,In_589);
or U571 (N_571,In_2263,In_934);
and U572 (N_572,In_1521,In_988);
and U573 (N_573,In_1641,In_2433);
or U574 (N_574,In_2199,In_593);
and U575 (N_575,In_1820,In_1008);
nand U576 (N_576,In_1553,In_1282);
and U577 (N_577,In_2399,In_2369);
nor U578 (N_578,In_1914,In_1839);
nand U579 (N_579,In_1010,In_824);
nor U580 (N_580,In_525,In_897);
xnor U581 (N_581,In_648,In_1592);
nor U582 (N_582,In_1767,In_1992);
and U583 (N_583,In_2011,In_1024);
nand U584 (N_584,In_1074,In_1035);
nor U585 (N_585,In_2422,In_35);
and U586 (N_586,In_1375,In_2300);
xnor U587 (N_587,In_957,In_2470);
and U588 (N_588,In_54,In_1077);
and U589 (N_589,In_803,In_2493);
nand U590 (N_590,In_2046,In_2082);
nand U591 (N_591,In_2149,In_1015);
nor U592 (N_592,In_2483,In_476);
or U593 (N_593,In_90,In_1419);
and U594 (N_594,In_367,In_1944);
nand U595 (N_595,In_1539,In_821);
xor U596 (N_596,In_2416,In_1714);
and U597 (N_597,In_348,In_1293);
and U598 (N_598,In_671,In_578);
nor U599 (N_599,In_1085,In_1842);
and U600 (N_600,In_438,In_731);
or U601 (N_601,In_621,In_629);
nor U602 (N_602,In_2306,In_584);
or U603 (N_603,In_313,In_491);
or U604 (N_604,In_700,In_1522);
or U605 (N_605,In_2442,In_2448);
or U606 (N_606,In_559,In_2045);
nand U607 (N_607,In_1589,In_677);
nand U608 (N_608,In_306,In_1021);
nor U609 (N_609,In_3,In_2);
xnor U610 (N_610,In_755,In_1064);
and U611 (N_611,In_1988,In_279);
nor U612 (N_612,In_687,In_2085);
nand U613 (N_613,In_1240,In_1542);
xor U614 (N_614,In_1048,In_1651);
or U615 (N_615,In_1843,In_1639);
nand U616 (N_616,In_1671,In_2285);
nand U617 (N_617,In_2424,In_1239);
and U618 (N_618,In_654,In_732);
and U619 (N_619,In_1256,In_1561);
xnor U620 (N_620,In_693,In_759);
xor U621 (N_621,In_2109,In_316);
nand U622 (N_622,In_147,In_2296);
and U623 (N_623,In_160,In_1560);
nand U624 (N_624,In_1537,In_1686);
and U625 (N_625,N_274,N_200);
xnor U626 (N_626,N_173,N_345);
or U627 (N_627,In_2097,In_685);
or U628 (N_628,In_582,N_278);
and U629 (N_629,In_2224,N_380);
and U630 (N_630,N_178,N_238);
nor U631 (N_631,N_343,N_584);
or U632 (N_632,In_893,N_622);
nand U633 (N_633,N_6,In_1428);
or U634 (N_634,N_495,N_379);
nand U635 (N_635,In_1025,In_585);
nor U636 (N_636,In_649,N_369);
nor U637 (N_637,In_1214,N_138);
nor U638 (N_638,In_2143,N_318);
and U639 (N_639,In_1618,In_1151);
nor U640 (N_640,N_519,N_20);
nand U641 (N_641,In_586,In_2117);
xnor U642 (N_642,In_1663,N_98);
nand U643 (N_643,N_172,In_2123);
and U644 (N_644,In_676,In_856);
or U645 (N_645,In_929,N_558);
or U646 (N_646,N_270,In_857);
nor U647 (N_647,In_106,In_1747);
nor U648 (N_648,In_1573,In_776);
or U649 (N_649,N_605,N_578);
and U650 (N_650,In_2171,In_2279);
nor U651 (N_651,In_170,In_473);
nand U652 (N_652,In_1216,N_514);
nand U653 (N_653,N_280,N_180);
or U654 (N_654,N_552,In_2056);
or U655 (N_655,In_1183,N_498);
nand U656 (N_656,In_2223,In_362);
nand U657 (N_657,In_555,In_1738);
xnor U658 (N_658,In_910,In_1108);
nor U659 (N_659,In_1850,N_491);
nor U660 (N_660,In_854,In_2274);
or U661 (N_661,In_901,In_324);
nand U662 (N_662,N_300,In_327);
nor U663 (N_663,In_298,N_441);
nand U664 (N_664,N_230,In_1668);
and U665 (N_665,In_2063,N_31);
and U666 (N_666,In_1247,N_428);
and U667 (N_667,In_1915,In_2293);
xor U668 (N_668,In_1648,In_664);
and U669 (N_669,In_1423,N_327);
nor U670 (N_670,In_1935,In_1394);
and U671 (N_671,In_2069,N_118);
nor U672 (N_672,In_303,In_1182);
nand U673 (N_673,In_1953,In_1490);
nor U674 (N_674,In_1119,In_1254);
nand U675 (N_675,In_955,In_102);
or U676 (N_676,In_2241,N_84);
nand U677 (N_677,In_2147,In_869);
or U678 (N_678,In_2394,In_1163);
nor U679 (N_679,In_1330,N_160);
or U680 (N_680,In_58,In_1908);
or U681 (N_681,In_1594,In_926);
or U682 (N_682,N_165,In_2255);
nor U683 (N_683,In_1649,In_1229);
nor U684 (N_684,In_1265,In_2165);
or U685 (N_685,In_1989,In_495);
xnor U686 (N_686,N_225,In_210);
and U687 (N_687,In_319,N_335);
and U688 (N_688,In_655,In_1053);
nand U689 (N_689,In_1902,N_467);
or U690 (N_690,N_459,In_1712);
or U691 (N_691,In_1404,N_94);
xor U692 (N_692,In_2027,N_338);
and U693 (N_693,In_862,In_2370);
xor U694 (N_694,N_271,In_2373);
nor U695 (N_695,N_110,N_356);
nand U696 (N_696,N_279,In_1737);
or U697 (N_697,N_290,N_472);
and U698 (N_698,N_227,N_568);
or U699 (N_699,In_2392,In_1410);
nor U700 (N_700,In_1218,In_2447);
or U701 (N_701,In_1782,In_2430);
or U702 (N_702,N_105,In_1425);
and U703 (N_703,In_2496,In_1579);
and U704 (N_704,N_496,N_26);
nand U705 (N_705,N_607,N_388);
nor U706 (N_706,N_146,N_102);
nand U707 (N_707,In_1067,In_2146);
nand U708 (N_708,N_59,In_896);
or U709 (N_709,In_2220,In_1695);
or U710 (N_710,N_396,In_2438);
nor U711 (N_711,N_358,In_2473);
and U712 (N_712,In_1818,In_162);
xnor U713 (N_713,In_919,In_829);
xor U714 (N_714,N_326,N_331);
nand U715 (N_715,In_167,N_422);
nand U716 (N_716,N_246,N_560);
nor U717 (N_717,N_420,N_393);
or U718 (N_718,N_608,N_257);
nand U719 (N_719,N_372,In_318);
nor U720 (N_720,In_239,N_128);
nor U721 (N_721,In_993,In_734);
nand U722 (N_722,N_44,In_2359);
nor U723 (N_723,N_10,N_32);
and U724 (N_724,In_2113,In_417);
nor U725 (N_725,N_166,In_2066);
or U726 (N_726,In_2431,N_196);
xnor U727 (N_727,N_337,In_1895);
or U728 (N_728,In_2482,N_233);
nand U729 (N_729,N_573,In_1603);
xnor U730 (N_730,N_235,N_297);
or U731 (N_731,N_402,In_1143);
or U732 (N_732,In_2228,N_304);
nand U733 (N_733,In_987,In_451);
nand U734 (N_734,N_370,In_2346);
or U735 (N_735,In_2121,N_56);
or U736 (N_736,In_1476,In_80);
or U737 (N_737,In_560,In_36);
or U738 (N_738,In_228,N_399);
xor U739 (N_739,N_286,In_420);
nand U740 (N_740,In_1049,In_301);
or U741 (N_741,N_72,In_189);
nor U742 (N_742,N_470,In_2384);
nor U743 (N_743,In_109,In_24);
and U744 (N_744,N_332,In_1332);
and U745 (N_745,N_186,In_2368);
or U746 (N_746,N_556,In_964);
xnor U747 (N_747,In_1870,N_464);
and U748 (N_748,In_1518,In_263);
or U749 (N_749,N_489,In_1099);
and U750 (N_750,In_29,N_535);
and U751 (N_751,In_1109,In_2180);
and U752 (N_752,In_1645,In_2452);
and U753 (N_753,N_61,In_1358);
nor U754 (N_754,In_368,In_57);
and U755 (N_755,In_1756,In_381);
xor U756 (N_756,N_592,In_903);
nand U757 (N_757,N_534,In_1892);
or U758 (N_758,In_1802,In_1337);
or U759 (N_759,In_710,In_1323);
and U760 (N_760,In_1678,In_1041);
nor U761 (N_761,In_1736,In_1346);
nor U762 (N_762,In_2485,N_259);
nand U763 (N_763,In_1794,In_1655);
and U764 (N_764,In_2314,In_1189);
and U765 (N_765,In_1480,N_328);
xnor U766 (N_766,In_1828,In_1920);
nand U767 (N_767,In_127,In_2043);
nor U768 (N_768,In_1483,In_2342);
or U769 (N_769,N_551,In_399);
or U770 (N_770,In_852,N_502);
or U771 (N_771,In_1942,N_435);
and U772 (N_772,In_1694,In_50);
xnor U773 (N_773,N_507,In_314);
or U774 (N_774,N_154,N_453);
or U775 (N_775,In_471,In_393);
xor U776 (N_776,In_1446,In_74);
nand U777 (N_777,In_1879,N_96);
and U778 (N_778,N_155,In_2348);
nor U779 (N_779,N_312,In_2273);
nor U780 (N_780,N_1,N_376);
and U781 (N_781,In_1621,N_291);
nand U782 (N_782,In_1826,In_1492);
nand U783 (N_783,In_1197,In_1526);
and U784 (N_784,In_1551,In_1000);
nand U785 (N_785,In_1405,In_2029);
and U786 (N_786,N_42,In_2415);
nor U787 (N_787,In_1396,In_1006);
nor U788 (N_788,N_281,In_1392);
nor U789 (N_789,In_2079,In_1374);
or U790 (N_790,N_481,In_1911);
nor U791 (N_791,In_53,In_333);
or U792 (N_792,In_44,In_1406);
or U793 (N_793,In_2281,N_430);
or U794 (N_794,In_974,In_400);
and U795 (N_795,In_467,In_412);
nor U796 (N_796,In_1602,In_315);
nor U797 (N_797,N_212,N_25);
nor U798 (N_798,N_197,In_287);
nand U799 (N_799,N_273,N_148);
xnor U800 (N_800,In_2068,In_1711);
and U801 (N_801,N_103,In_204);
or U802 (N_802,In_2219,N_226);
and U803 (N_803,In_541,In_1196);
nand U804 (N_804,In_774,In_1238);
and U805 (N_805,N_360,N_251);
xnor U806 (N_806,N_95,N_559);
xnor U807 (N_807,N_161,In_1314);
nand U808 (N_808,N_624,In_750);
and U809 (N_809,N_357,In_156);
and U810 (N_810,N_213,In_1730);
nor U811 (N_811,In_562,N_383);
or U812 (N_812,N_127,In_1882);
nor U813 (N_813,N_473,In_2166);
or U814 (N_814,In_1129,In_2282);
and U815 (N_815,N_619,In_1505);
nand U816 (N_816,N_142,In_2119);
nor U817 (N_817,In_2347,N_236);
nand U818 (N_818,In_579,In_458);
nand U819 (N_819,In_1422,In_650);
nor U820 (N_820,N_124,N_438);
or U821 (N_821,In_291,In_735);
nor U822 (N_822,In_689,In_484);
xnor U823 (N_823,In_2425,In_1340);
nor U824 (N_824,N_210,In_2413);
or U825 (N_825,N_598,In_701);
nor U826 (N_826,In_1559,In_164);
and U827 (N_827,N_508,In_2407);
xnor U828 (N_828,In_675,N_67);
nor U829 (N_829,In_346,N_113);
nand U830 (N_830,In_12,N_342);
nand U831 (N_831,N_503,N_545);
nor U832 (N_832,N_179,In_1627);
and U833 (N_833,In_322,In_1946);
nor U834 (N_834,N_29,In_1742);
nor U835 (N_835,N_194,In_366);
nand U836 (N_836,In_989,N_384);
and U837 (N_837,In_378,In_2138);
xor U838 (N_838,N_28,In_2449);
and U839 (N_839,In_652,In_13);
nor U840 (N_840,In_2176,In_1190);
and U841 (N_841,N_205,In_1691);
or U842 (N_842,In_1927,In_231);
nor U843 (N_843,In_785,N_46);
xor U844 (N_844,In_254,In_1357);
or U845 (N_845,N_253,N_595);
or U846 (N_846,In_1688,In_1896);
nor U847 (N_847,In_1871,In_410);
or U848 (N_848,N_80,In_64);
nand U849 (N_849,In_2463,In_2428);
or U850 (N_850,In_1945,In_270);
nor U851 (N_851,N_207,N_319);
or U852 (N_852,N_572,N_70);
nand U853 (N_853,In_255,In_250);
or U854 (N_854,In_271,In_2427);
or U855 (N_855,N_89,N_135);
nand U856 (N_856,In_16,In_1033);
nor U857 (N_857,N_133,In_213);
and U858 (N_858,In_1421,In_1474);
or U859 (N_859,N_38,In_2136);
and U860 (N_860,N_269,In_2096);
and U861 (N_861,In_88,In_243);
or U862 (N_862,In_119,In_800);
xor U863 (N_863,N_482,In_1028);
nand U864 (N_864,N_576,In_56);
nor U865 (N_865,N_314,N_292);
or U866 (N_866,In_2008,In_130);
xnor U867 (N_867,In_149,In_2334);
nand U868 (N_868,N_49,In_1607);
and U869 (N_869,In_1291,In_1666);
xor U870 (N_870,In_594,N_287);
nand U871 (N_871,In_2083,In_275);
nand U872 (N_872,N_66,In_1115);
nand U873 (N_873,In_612,In_1056);
nand U874 (N_874,In_134,In_73);
and U875 (N_875,In_1188,In_1334);
nor U876 (N_876,In_117,In_1792);
nand U877 (N_877,In_1633,In_2365);
nand U878 (N_878,In_1960,N_3);
and U879 (N_879,In_2350,N_22);
and U880 (N_880,In_1475,In_549);
nand U881 (N_881,N_488,In_1485);
xor U882 (N_882,N_333,In_209);
or U883 (N_883,In_1009,In_727);
or U884 (N_884,In_851,N_408);
or U885 (N_885,In_1954,In_768);
nand U886 (N_886,N_367,In_2037);
or U887 (N_887,In_2053,N_513);
xnor U888 (N_888,In_2408,In_1147);
and U889 (N_889,In_1339,N_204);
nand U890 (N_890,In_1934,N_512);
xor U891 (N_891,In_868,In_936);
and U892 (N_892,In_879,In_746);
nand U893 (N_893,In_1230,N_323);
nand U894 (N_894,In_274,In_1333);
and U895 (N_895,N_168,In_845);
or U896 (N_896,N_35,In_1548);
nor U897 (N_897,In_486,In_1261);
nor U898 (N_898,In_604,N_583);
nand U899 (N_899,In_2174,In_1912);
nor U900 (N_900,In_754,In_1507);
or U901 (N_901,In_1692,N_248);
nand U902 (N_902,In_885,N_449);
or U903 (N_903,In_2058,In_2311);
and U904 (N_904,N_17,N_264);
nor U905 (N_905,In_59,In_1869);
nand U906 (N_906,N_177,In_1725);
nor U907 (N_907,In_1296,In_2379);
or U908 (N_908,N_403,In_1910);
and U909 (N_909,In_2268,N_533);
nand U910 (N_910,In_1233,N_541);
nor U911 (N_911,In_2188,In_1704);
nor U912 (N_912,In_1288,N_322);
and U913 (N_913,N_442,In_1133);
xor U914 (N_914,N_283,In_625);
nor U915 (N_915,N_366,In_1264);
nor U916 (N_916,In_1931,In_1503);
nor U917 (N_917,In_98,N_579);
nor U918 (N_918,N_65,N_462);
or U919 (N_919,In_1540,In_124);
nand U920 (N_920,In_2088,N_336);
nor U921 (N_921,N_613,In_543);
nand U922 (N_922,N_445,In_1416);
nand U923 (N_923,In_843,N_523);
and U924 (N_924,In_1252,N_108);
xor U925 (N_925,In_419,In_1486);
and U926 (N_926,In_1997,N_52);
or U927 (N_927,In_554,N_381);
nor U928 (N_928,In_859,In_17);
nand U929 (N_929,N_599,In_396);
or U930 (N_930,N_219,In_1898);
and U931 (N_931,In_967,In_300);
nor U932 (N_932,In_622,In_1761);
nor U933 (N_933,In_2237,In_1489);
and U934 (N_934,In_767,In_148);
nand U935 (N_935,N_418,In_449);
xnor U936 (N_936,N_601,In_2178);
and U937 (N_937,In_1733,N_590);
xnor U938 (N_938,In_818,N_85);
or U939 (N_939,In_1488,N_382);
and U940 (N_940,In_413,N_394);
nor U941 (N_941,N_54,In_457);
nor U942 (N_942,In_2118,N_474);
nand U943 (N_943,In_2235,In_2226);
nor U944 (N_944,N_121,In_335);
and U945 (N_945,N_609,In_984);
nand U946 (N_946,In_2286,N_272);
and U947 (N_947,In_1128,In_1532);
nand U948 (N_948,N_215,In_2200);
nor U949 (N_949,In_1635,In_2205);
nor U950 (N_950,N_518,In_475);
nand U951 (N_951,In_630,In_1781);
or U952 (N_952,N_530,In_511);
xor U953 (N_953,In_437,In_1722);
nand U954 (N_954,N_71,In_2456);
nand U955 (N_955,In_500,In_1620);
or U956 (N_956,N_305,In_2253);
nor U957 (N_957,N_436,In_1352);
and U958 (N_958,In_1894,In_217);
and U959 (N_959,In_882,In_2356);
nor U960 (N_960,N_256,In_1709);
or U961 (N_961,N_190,In_1309);
and U962 (N_962,N_51,In_1436);
or U963 (N_963,In_952,N_43);
xor U964 (N_964,In_200,In_2385);
and U965 (N_965,N_567,N_234);
nand U966 (N_966,In_62,In_517);
and U967 (N_967,In_2406,In_781);
and U968 (N_968,N_340,In_1088);
nand U969 (N_969,N_506,In_1226);
xnor U970 (N_970,N_143,In_1814);
nand U971 (N_971,N_139,In_118);
nand U972 (N_972,N_424,N_117);
or U973 (N_973,In_1222,In_360);
and U974 (N_974,In_195,In_673);
or U975 (N_975,In_942,In_1383);
xor U976 (N_976,In_1973,N_199);
or U977 (N_977,N_245,N_86);
nor U978 (N_978,In_895,In_1643);
nor U979 (N_979,In_1675,In_474);
nand U980 (N_980,In_1878,In_1966);
nor U981 (N_981,In_405,N_603);
or U982 (N_982,In_2383,In_1198);
nand U983 (N_983,In_646,N_400);
or U984 (N_984,N_16,In_788);
nor U985 (N_985,In_1403,In_892);
or U986 (N_986,In_2367,In_1173);
or U987 (N_987,In_668,In_2122);
nand U988 (N_988,N_63,In_1701);
nand U989 (N_989,In_2336,In_909);
or U990 (N_990,N_525,In_2251);
and U991 (N_991,In_1027,In_2249);
and U992 (N_992,In_2225,N_159);
or U993 (N_993,N_604,In_1205);
nand U994 (N_994,In_1019,In_830);
or U995 (N_995,In_772,In_1199);
xnor U996 (N_996,N_50,N_294);
nor U997 (N_997,In_1316,N_183);
xnor U998 (N_998,In_2015,In_1382);
and U999 (N_999,In_341,In_1728);
nand U1000 (N_1000,N_131,N_504);
xor U1001 (N_1001,N_122,In_2278);
nor U1002 (N_1002,N_554,In_1272);
or U1003 (N_1003,In_371,In_515);
or U1004 (N_1004,In_143,In_796);
and U1005 (N_1005,In_2196,In_2001);
or U1006 (N_1006,N_184,N_516);
nor U1007 (N_1007,In_196,N_359);
and U1008 (N_1008,In_20,In_1710);
and U1009 (N_1009,N_377,In_39);
and U1010 (N_1010,In_2005,N_526);
nand U1011 (N_1011,In_2229,N_451);
nor U1012 (N_1012,In_259,N_371);
or U1013 (N_1013,In_1380,In_1412);
nor U1014 (N_1014,In_233,In_2042);
or U1015 (N_1015,N_497,In_763);
and U1016 (N_1016,In_672,In_1159);
nand U1017 (N_1017,N_412,In_440);
nor U1018 (N_1018,N_374,N_589);
and U1019 (N_1019,In_1111,In_2179);
nor U1020 (N_1020,In_2325,N_47);
or U1021 (N_1021,In_1816,N_162);
xnor U1022 (N_1022,In_790,In_1126);
nor U1023 (N_1023,In_1127,N_0);
or U1024 (N_1024,In_1387,In_479);
and U1025 (N_1025,In_1762,In_1634);
nand U1026 (N_1026,In_2065,N_591);
and U1027 (N_1027,N_282,N_203);
or U1028 (N_1028,In_2436,In_1825);
and U1029 (N_1029,In_2003,In_1948);
nor U1030 (N_1030,In_1907,In_1203);
and U1031 (N_1031,In_587,In_1391);
or U1032 (N_1032,In_996,In_2499);
and U1033 (N_1033,In_506,In_1807);
or U1034 (N_1034,In_1350,In_799);
or U1035 (N_1035,In_2099,N_434);
nor U1036 (N_1036,In_1929,N_373);
and U1037 (N_1037,In_1848,In_1821);
nor U1038 (N_1038,In_1700,N_306);
and U1039 (N_1039,N_254,In_1723);
or U1040 (N_1040,In_1305,In_232);
xor U1041 (N_1041,In_720,N_618);
and U1042 (N_1042,In_1772,In_867);
or U1043 (N_1043,N_487,N_192);
or U1044 (N_1044,N_243,N_265);
and U1045 (N_1045,N_405,In_1752);
nand U1046 (N_1046,In_1799,In_2444);
or U1047 (N_1047,N_107,In_2476);
and U1048 (N_1048,In_2434,N_252);
nor U1049 (N_1049,In_2025,In_1308);
or U1050 (N_1050,In_718,In_1741);
nand U1051 (N_1051,N_387,In_945);
or U1052 (N_1052,N_170,In_1545);
and U1053 (N_1053,In_1740,In_2421);
nand U1054 (N_1054,In_285,N_365);
nand U1055 (N_1055,In_1065,In_847);
nor U1056 (N_1056,In_245,N_21);
nand U1057 (N_1057,N_73,In_286);
nor U1058 (N_1058,N_150,In_1512);
nor U1059 (N_1059,In_1149,In_659);
and U1060 (N_1060,N_458,In_2172);
and U1061 (N_1061,N_228,In_1132);
and U1062 (N_1062,N_60,In_2377);
nor U1063 (N_1063,In_1208,In_1913);
and U1064 (N_1064,In_1832,N_562);
or U1065 (N_1065,In_34,In_377);
or U1066 (N_1066,In_252,N_454);
or U1067 (N_1067,N_361,N_262);
and U1068 (N_1068,In_2461,N_268);
and U1069 (N_1069,N_389,In_1349);
or U1070 (N_1070,N_267,N_484);
and U1071 (N_1071,N_39,In_2254);
nor U1072 (N_1072,In_1051,N_145);
nand U1073 (N_1073,In_108,N_69);
nor U1074 (N_1074,In_507,In_1094);
nor U1075 (N_1075,N_296,In_2299);
nand U1076 (N_1076,In_2160,In_1861);
nand U1077 (N_1077,N_433,In_1164);
nor U1078 (N_1078,In_2047,N_501);
and U1079 (N_1079,In_528,In_2151);
or U1080 (N_1080,N_100,N_2);
nor U1081 (N_1081,In_1860,In_278);
nor U1082 (N_1082,In_137,N_55);
nor U1083 (N_1083,In_1637,In_523);
and U1084 (N_1084,In_267,N_34);
nand U1085 (N_1085,In_1581,N_275);
and U1086 (N_1086,In_1286,In_1045);
nor U1087 (N_1087,N_623,In_439);
xor U1088 (N_1088,N_364,In_1134);
nand U1089 (N_1089,N_320,In_1569);
and U1090 (N_1090,In_1031,N_615);
nor U1091 (N_1091,In_283,In_289);
xor U1092 (N_1092,N_14,In_1916);
and U1093 (N_1093,In_1574,N_415);
nor U1094 (N_1094,N_532,In_1784);
xnor U1095 (N_1095,In_1376,In_978);
and U1096 (N_1096,In_1830,In_1054);
and U1097 (N_1097,N_531,N_62);
nor U1098 (N_1098,In_1582,N_597);
nand U1099 (N_1099,N_316,In_8);
nand U1100 (N_1100,N_537,In_427);
or U1101 (N_1101,In_1176,In_2014);
or U1102 (N_1102,In_15,N_237);
nand U1103 (N_1103,In_469,In_1);
nor U1104 (N_1104,In_2071,N_446);
and U1105 (N_1105,In_2221,In_808);
and U1106 (N_1106,In_1508,In_1549);
and U1107 (N_1107,N_307,In_963);
or U1108 (N_1108,N_325,N_477);
and U1109 (N_1109,N_409,In_2044);
nor U1110 (N_1110,In_623,N_460);
nor U1111 (N_1111,In_1604,In_1557);
or U1112 (N_1112,In_2335,In_95);
nand U1113 (N_1113,N_499,In_230);
nand U1114 (N_1114,In_2102,In_591);
or U1115 (N_1115,In_1213,In_890);
or U1116 (N_1116,N_429,In_1201);
or U1117 (N_1117,N_427,N_153);
or U1118 (N_1118,N_9,In_169);
or U1119 (N_1119,In_1991,N_351);
and U1120 (N_1120,In_711,N_119);
and U1121 (N_1121,N_33,In_1228);
nor U1122 (N_1122,In_2232,N_486);
and U1123 (N_1123,In_877,In_2154);
nor U1124 (N_1124,In_1036,In_415);
nand U1125 (N_1125,N_109,In_82);
xor U1126 (N_1126,In_575,N_398);
and U1127 (N_1127,In_2423,In_1606);
nor U1128 (N_1128,In_2252,N_104);
xor U1129 (N_1129,N_217,In_1638);
nor U1130 (N_1130,In_1437,In_447);
nor U1131 (N_1131,In_2114,In_590);
or U1132 (N_1132,In_924,In_1838);
or U1133 (N_1133,In_2081,N_247);
nor U1134 (N_1134,N_255,In_2264);
nor U1135 (N_1135,In_176,N_557);
or U1136 (N_1136,N_392,In_736);
and U1137 (N_1137,In_69,In_2454);
nor U1138 (N_1138,In_501,N_24);
or U1139 (N_1139,In_266,In_657);
or U1140 (N_1140,In_1170,In_556);
nor U1141 (N_1141,In_159,N_524);
nand U1142 (N_1142,N_239,In_407);
and U1143 (N_1143,In_1249,In_212);
nor U1144 (N_1144,In_1156,In_2319);
nand U1145 (N_1145,In_409,In_1206);
xor U1146 (N_1146,In_398,N_417);
nor U1147 (N_1147,In_1178,N_261);
nor U1148 (N_1148,In_1743,In_194);
or U1149 (N_1149,N_432,In_297);
and U1150 (N_1150,In_464,N_355);
and U1151 (N_1151,N_45,N_208);
and U1152 (N_1152,In_906,In_1102);
nor U1153 (N_1153,N_244,N_444);
nand U1154 (N_1154,N_140,N_517);
nand U1155 (N_1155,In_1514,In_2353);
nand U1156 (N_1156,In_797,In_1457);
and U1157 (N_1157,In_665,In_577);
nand U1158 (N_1158,In_1926,In_311);
or U1159 (N_1159,In_391,N_544);
nand U1160 (N_1160,In_2322,N_299);
or U1161 (N_1161,In_641,In_875);
or U1162 (N_1162,In_459,In_2247);
and U1163 (N_1163,In_2364,N_522);
nand U1164 (N_1164,N_99,In_1451);
and U1165 (N_1165,In_1735,N_187);
xor U1166 (N_1166,In_1865,In_684);
xor U1167 (N_1167,N_401,In_219);
nor U1168 (N_1168,N_90,In_1287);
and U1169 (N_1169,In_1886,In_2405);
and U1170 (N_1170,In_1001,In_1979);
or U1171 (N_1171,In_1434,In_1179);
xnor U1172 (N_1172,In_1172,N_149);
nor U1173 (N_1173,N_548,In_1790);
nor U1174 (N_1174,N_346,In_141);
or U1175 (N_1175,In_535,In_43);
xnor U1176 (N_1176,N_75,N_123);
and U1177 (N_1177,In_1938,In_1851);
and U1178 (N_1178,In_1101,In_380);
nor U1179 (N_1179,In_733,In_2446);
nand U1180 (N_1180,N_577,In_827);
xnor U1181 (N_1181,In_23,In_1959);
xnor U1182 (N_1182,N_222,In_1586);
or U1183 (N_1183,In_2375,N_341);
xor U1184 (N_1184,N_258,N_315);
and U1185 (N_1185,In_1066,In_2403);
and U1186 (N_1186,N_448,In_395);
and U1187 (N_1187,In_2211,N_600);
nor U1188 (N_1188,In_273,N_529);
or U1189 (N_1189,In_666,In_406);
nand U1190 (N_1190,In_553,In_2295);
nor U1191 (N_1191,N_593,In_1258);
or U1192 (N_1192,In_956,In_2158);
nor U1193 (N_1193,In_432,N_350);
nand U1194 (N_1194,N_476,In_1023);
and U1195 (N_1195,In_1413,N_362);
nor U1196 (N_1196,In_1763,N_53);
and U1197 (N_1197,In_633,In_1069);
nand U1198 (N_1198,N_27,N_457);
nor U1199 (N_1199,N_201,N_211);
nor U1200 (N_1200,In_163,In_1683);
nor U1201 (N_1201,In_1981,In_1970);
or U1202 (N_1202,In_1530,In_2324);
or U1203 (N_1203,In_1136,In_2297);
nand U1204 (N_1204,N_621,In_1237);
and U1205 (N_1205,N_301,In_2376);
or U1206 (N_1206,In_2393,In_370);
and U1207 (N_1207,In_1104,In_111);
nor U1208 (N_1208,In_547,In_1924);
and U1209 (N_1209,In_770,In_203);
or U1210 (N_1210,In_1071,In_2156);
and U1211 (N_1211,In_1046,In_1764);
xor U1212 (N_1212,In_237,N_485);
nor U1213 (N_1213,In_434,In_719);
nor U1214 (N_1214,In_2363,In_1364);
nor U1215 (N_1215,N_413,In_1342);
nand U1216 (N_1216,N_542,N_284);
or U1217 (N_1217,N_91,In_2163);
nor U1218 (N_1218,N_181,In_1819);
nand U1219 (N_1219,In_1893,N_106);
nand U1220 (N_1220,In_1952,In_1855);
and U1221 (N_1221,N_347,N_30);
nor U1222 (N_1222,In_2498,N_147);
xor U1223 (N_1223,N_15,In_1856);
and U1224 (N_1224,In_1884,N_443);
and U1225 (N_1225,In_358,In_958);
or U1226 (N_1226,In_296,In_1619);
and U1227 (N_1227,In_1411,N_469);
nand U1228 (N_1228,N_182,N_152);
nand U1229 (N_1229,In_430,In_1366);
nor U1230 (N_1230,In_1429,In_2290);
nand U1231 (N_1231,In_2162,N_617);
nand U1232 (N_1232,In_588,N_285);
or U1233 (N_1233,N_550,N_144);
nand U1234 (N_1234,In_1452,In_871);
nor U1235 (N_1235,N_276,In_944);
xor U1236 (N_1236,In_312,In_982);
and U1237 (N_1237,In_226,N_575);
nand U1238 (N_1238,In_613,In_839);
and U1239 (N_1239,In_468,In_943);
nor U1240 (N_1240,N_240,In_1267);
or U1241 (N_1241,In_216,N_266);
nor U1242 (N_1242,In_1824,N_391);
nand U1243 (N_1243,In_618,In_2362);
nor U1244 (N_1244,N_232,In_1123);
nor U1245 (N_1245,In_1070,N_520);
nor U1246 (N_1246,In_337,In_518);
nor U1247 (N_1247,In_1301,In_1888);
nor U1248 (N_1248,In_2072,N_425);
or U1249 (N_1249,In_1236,In_1629);
nor U1250 (N_1250,N_1071,N_511);
and U1251 (N_1251,N_779,N_125);
nand U1252 (N_1252,N_718,N_1112);
nand U1253 (N_1253,N_1244,In_2108);
nand U1254 (N_1254,N_1245,N_970);
xnor U1255 (N_1255,N_1018,N_811);
nor U1256 (N_1256,In_2487,In_1322);
or U1257 (N_1257,N_375,N_349);
nand U1258 (N_1258,N_1161,N_1204);
nand U1259 (N_1259,N_414,N_1111);
xor U1260 (N_1260,In_1932,N_450);
or U1261 (N_1261,In_1900,In_2310);
xor U1262 (N_1262,N_1095,N_945);
nand U1263 (N_1263,In_453,In_1184);
and U1264 (N_1264,N_727,N_733);
or U1265 (N_1265,In_504,N_807);
xor U1266 (N_1266,In_1812,N_13);
xor U1267 (N_1267,In_1082,In_1447);
or U1268 (N_1268,In_416,In_1890);
nand U1269 (N_1269,N_695,In_860);
xnor U1270 (N_1270,N_1034,N_221);
and U1271 (N_1271,In_1146,In_338);
nor U1272 (N_1272,N_1058,In_815);
nand U1273 (N_1273,N_397,N_972);
nand U1274 (N_1274,N_1076,N_757);
nand U1275 (N_1275,In_2073,N_1192);
nand U1276 (N_1276,N_1249,In_642);
nand U1277 (N_1277,N_977,N_1114);
or U1278 (N_1278,N_925,In_1525);
and U1279 (N_1279,N_78,N_1134);
or U1280 (N_1280,N_766,In_1155);
nand U1281 (N_1281,N_761,N_1087);
nor U1282 (N_1282,N_804,N_461);
xor U1283 (N_1283,N_1053,In_1599);
and U1284 (N_1284,N_627,In_472);
nor U1285 (N_1285,In_1567,N_933);
or U1286 (N_1286,N_1131,In_1531);
nor U1287 (N_1287,In_1836,N_724);
nand U1288 (N_1288,In_1438,In_702);
and U1289 (N_1289,N_1031,N_1202);
xnor U1290 (N_1290,N_680,N_157);
or U1291 (N_1291,In_838,In_155);
and U1292 (N_1292,N_581,In_635);
and U1293 (N_1293,In_814,N_1165);
xnor U1294 (N_1294,N_633,N_1122);
nor U1295 (N_1295,N_395,N_836);
and U1296 (N_1296,N_1092,N_1070);
xor U1297 (N_1297,N_93,N_1189);
nor U1298 (N_1298,In_2340,N_1032);
nand U1299 (N_1299,In_980,N_801);
or U1300 (N_1300,In_2023,N_797);
nor U1301 (N_1301,N_841,N_1046);
nor U1302 (N_1302,N_709,N_827);
nor U1303 (N_1303,N_985,In_1872);
nand U1304 (N_1304,N_795,N_185);
nor U1305 (N_1305,In_280,N_419);
nor U1306 (N_1306,N_840,N_1080);
or U1307 (N_1307,In_1285,N_1166);
and U1308 (N_1308,N_574,In_741);
nor U1309 (N_1309,In_292,N_772);
nand U1310 (N_1310,N_1041,In_2308);
and U1311 (N_1311,N_981,N_792);
nand U1312 (N_1312,N_720,N_892);
nand U1313 (N_1313,N_1026,In_569);
nor U1314 (N_1314,In_443,In_2242);
or U1315 (N_1315,N_913,N_437);
nor U1316 (N_1316,In_971,N_819);
nand U1317 (N_1317,In_1204,In_1509);
nand U1318 (N_1318,N_938,N_1239);
and U1319 (N_1319,N_1175,N_1225);
nor U1320 (N_1320,N_991,In_2287);
and U1321 (N_1321,In_1734,In_1361);
nor U1322 (N_1322,In_197,N_1052);
nor U1323 (N_1323,N_1027,N_824);
xnor U1324 (N_1324,N_302,N_404);
and U1325 (N_1325,N_313,In_1343);
and U1326 (N_1326,N_348,In_493);
and U1327 (N_1327,In_1857,N_390);
nand U1328 (N_1328,N_493,In_1984);
and U1329 (N_1329,N_1160,N_954);
xnor U1330 (N_1330,In_1494,N_1221);
and U1331 (N_1331,N_1180,In_1983);
nor U1332 (N_1332,N_134,N_587);
nor U1333 (N_1333,In_215,In_1965);
nor U1334 (N_1334,In_706,N_363);
and U1335 (N_1335,N_191,In_2067);
and U1336 (N_1336,In_408,N_740);
or U1337 (N_1337,N_758,In_580);
nand U1338 (N_1338,N_675,N_632);
nor U1339 (N_1339,In_1219,In_1815);
nand U1340 (N_1340,In_1245,N_1194);
and U1341 (N_1341,In_990,In_2218);
nor U1342 (N_1342,N_767,N_962);
or U1343 (N_1343,In_935,N_321);
nand U1344 (N_1344,N_721,In_2132);
and U1345 (N_1345,N_921,N_288);
nand U1346 (N_1346,In_1424,In_2239);
nor U1347 (N_1347,In_751,N_521);
or U1348 (N_1348,N_478,In_637);
nor U1349 (N_1349,N_903,N_964);
xor U1350 (N_1350,N_866,N_1182);
nor U1351 (N_1351,N_353,N_1002);
and U1352 (N_1352,N_1164,N_714);
nor U1353 (N_1353,N_465,In_1771);
or U1354 (N_1354,N_1098,N_1113);
and U1355 (N_1355,N_672,N_510);
and U1356 (N_1356,N_421,N_871);
or U1357 (N_1357,In_986,N_585);
xnor U1358 (N_1358,In_1495,N_169);
nor U1359 (N_1359,N_1209,N_1060);
xnor U1360 (N_1360,N_8,In_265);
nor U1361 (N_1361,N_198,N_1106);
nand U1362 (N_1362,In_2013,In_1243);
nand U1363 (N_1363,N_1136,In_2095);
nand U1364 (N_1364,N_800,In_1804);
or U1365 (N_1365,N_802,In_1341);
or U1366 (N_1366,N_339,N_1061);
or U1367 (N_1367,N_762,N_746);
nand U1368 (N_1368,N_637,In_1469);
nand U1369 (N_1369,N_940,N_76);
and U1370 (N_1370,In_644,N_723);
and U1371 (N_1371,In_2445,In_707);
or U1372 (N_1372,N_958,In_2019);
nor U1373 (N_1373,N_1174,In_1906);
nand U1374 (N_1374,In_2313,N_961);
nand U1375 (N_1375,In_357,N_976);
nand U1376 (N_1376,In_2100,In_1290);
xor U1377 (N_1377,N_1188,N_1101);
nor U1378 (N_1378,In_758,In_2076);
nand U1379 (N_1379,N_1228,N_1000);
nor U1380 (N_1380,In_2216,N_781);
nand U1381 (N_1381,In_1769,In_712);
nor U1382 (N_1382,N_406,N_1075);
nand U1383 (N_1383,In_608,N_943);
nand U1384 (N_1384,N_658,N_468);
and U1385 (N_1385,N_897,N_858);
and U1386 (N_1386,N_411,In_1461);
and U1387 (N_1387,N_645,N_754);
or U1388 (N_1388,N_423,N_527);
nor U1389 (N_1389,In_2210,N_639);
nor U1390 (N_1390,In_717,In_152);
or U1391 (N_1391,N_873,In_1456);
nor U1392 (N_1392,In_2110,N_1105);
nor U1393 (N_1393,N_1213,N_1073);
nand U1394 (N_1394,N_844,N_697);
and U1395 (N_1395,In_390,In_2275);
or U1396 (N_1396,N_630,N_895);
nor U1397 (N_1397,In_2395,In_1726);
nand U1398 (N_1398,N_1104,In_2323);
and U1399 (N_1399,N_670,N_955);
nand U1400 (N_1400,In_1897,In_1681);
and U1401 (N_1401,In_1930,N_483);
nand U1402 (N_1402,N_1062,N_755);
and U1403 (N_1403,N_1133,N_826);
xnor U1404 (N_1404,N_683,N_158);
and U1405 (N_1405,N_1121,N_1196);
xnor U1406 (N_1406,In_246,N_855);
and U1407 (N_1407,N_691,N_1096);
nor U1408 (N_1408,In_1212,N_997);
nand U1409 (N_1409,N_854,N_1181);
and U1410 (N_1410,N_864,N_1033);
xor U1411 (N_1411,N_982,N_701);
and U1412 (N_1412,In_1796,N_959);
nor U1413 (N_1413,N_768,In_2107);
and U1414 (N_1414,N_136,N_1235);
nand U1415 (N_1415,N_999,N_674);
and U1416 (N_1416,In_1626,N_606);
nand U1417 (N_1417,In_2140,In_1106);
and U1418 (N_1418,N_640,In_1356);
nor U1419 (N_1419,N_1001,N_664);
nand U1420 (N_1420,N_1097,In_2466);
or U1421 (N_1421,N_1064,In_2317);
xor U1422 (N_1422,In_1468,N_1132);
nand U1423 (N_1423,N_1012,N_856);
nor U1424 (N_1424,N_463,N_1015);
nor U1425 (N_1425,N_950,In_1174);
and U1426 (N_1426,N_687,In_789);
or U1427 (N_1427,N_651,In_1625);
and U1428 (N_1428,N_773,N_769);
nand U1429 (N_1429,N_116,N_678);
or U1430 (N_1430,N_1203,N_823);
nor U1431 (N_1431,In_1601,In_965);
or U1432 (N_1432,N_996,N_1066);
or U1433 (N_1433,In_662,N_547);
nor U1434 (N_1434,N_825,In_1866);
nor U1435 (N_1435,N_1057,N_920);
or U1436 (N_1436,N_635,In_1139);
nand U1437 (N_1437,N_588,In_1224);
nor U1438 (N_1438,N_1247,In_2105);
nor U1439 (N_1439,In_1928,N_132);
and U1440 (N_1440,In_884,N_1059);
and U1441 (N_1441,N_561,In_962);
or U1442 (N_1442,N_765,N_713);
and U1443 (N_1443,N_475,N_842);
and U1444 (N_1444,In_71,In_1980);
and U1445 (N_1445,N_876,N_1067);
nor U1446 (N_1446,In_696,In_2244);
nor U1447 (N_1447,N_900,In_1793);
nand U1448 (N_1448,N_1009,In_199);
nand U1449 (N_1449,In_192,N_129);
or U1450 (N_1450,In_2055,N_1216);
and U1451 (N_1451,In_490,In_1544);
and U1452 (N_1452,N_923,N_1215);
and U1453 (N_1453,In_487,N_12);
and U1454 (N_1454,N_1238,N_466);
or U1455 (N_1455,N_368,In_1022);
or U1456 (N_1456,N_692,N_1191);
and U1457 (N_1457,N_918,N_1047);
or U1458 (N_1458,In_1327,N_87);
nand U1459 (N_1459,In_2259,N_126);
or U1460 (N_1460,In_1324,N_993);
nor U1461 (N_1461,In_401,N_859);
nand U1462 (N_1462,N_298,In_1538);
or U1463 (N_1463,N_77,N_995);
and U1464 (N_1464,N_820,N_835);
nand U1465 (N_1465,In_1103,N_805);
xor U1466 (N_1466,N_666,N_1155);
nand U1467 (N_1467,In_1003,In_2215);
nand U1468 (N_1468,In_387,N_742);
or U1469 (N_1469,N_553,N_839);
and U1470 (N_1470,N_747,N_1127);
and U1471 (N_1471,In_364,N_277);
nand U1472 (N_1472,N_922,In_2126);
nand U1473 (N_1473,In_1611,N_555);
and U1474 (N_1474,N_969,N_308);
nor U1475 (N_1475,In_1144,In_592);
xor U1476 (N_1476,In_330,N_1030);
nand U1477 (N_1477,In_489,N_764);
and U1478 (N_1478,N_917,N_960);
and U1479 (N_1479,N_974,In_1453);
nor U1480 (N_1480,N_775,N_546);
and U1481 (N_1481,N_163,In_179);
xor U1482 (N_1482,N_1120,N_705);
nor U1483 (N_1483,N_654,In_78);
and U1484 (N_1484,N_906,N_696);
nand U1485 (N_1485,N_5,N_846);
and U1486 (N_1486,N_1025,N_655);
nor U1487 (N_1487,N_1223,N_965);
nand U1488 (N_1488,N_1170,N_1162);
nor U1489 (N_1489,N_657,In_352);
xnor U1490 (N_1490,N_1214,In_379);
and U1491 (N_1491,N_447,N_1019);
nand U1492 (N_1492,In_505,N_879);
and U1493 (N_1493,In_225,In_2479);
nor U1494 (N_1494,N_649,N_1197);
and U1495 (N_1495,N_886,N_1117);
or U1496 (N_1496,N_164,N_716);
and U1497 (N_1497,N_893,N_979);
nor U1498 (N_1498,N_798,N_957);
or U1499 (N_1499,In_411,In_1636);
nor U1500 (N_1500,N_156,N_1081);
nand U1501 (N_1501,N_852,N_828);
nand U1502 (N_1502,N_887,N_681);
nand U1503 (N_1503,In_1687,In_105);
or U1504 (N_1504,In_674,N_209);
or U1505 (N_1505,N_810,N_295);
xnor U1506 (N_1506,N_908,N_249);
nor U1507 (N_1507,N_809,In_1121);
nor U1508 (N_1508,N_751,In_89);
nand U1509 (N_1509,N_845,N_1011);
or U1510 (N_1510,In_1975,In_2420);
and U1511 (N_1511,N_1008,In_1227);
nand U1512 (N_1512,N_410,N_1100);
xor U1513 (N_1513,N_37,N_898);
nor U1514 (N_1514,In_834,N_966);
nand U1515 (N_1515,In_2004,N_582);
nand U1516 (N_1516,In_1455,N_188);
and U1517 (N_1517,N_354,N_1163);
and U1518 (N_1518,In_2248,In_1097);
nor U1519 (N_1519,N_1039,N_571);
and U1520 (N_1520,N_662,In_463);
and U1521 (N_1521,N_1050,N_141);
and U1522 (N_1522,In_2492,N_1118);
nor U1523 (N_1523,In_1597,N_83);
xor U1524 (N_1524,N_647,N_785);
or U1525 (N_1525,N_223,N_515);
and U1526 (N_1526,In_1034,In_454);
and U1527 (N_1527,N_480,N_1024);
nand U1528 (N_1528,N_137,N_719);
nand U1529 (N_1529,N_471,N_869);
nand U1530 (N_1530,In_1449,N_872);
nand U1531 (N_1531,N_565,N_229);
nand U1532 (N_1532,N_878,In_6);
xnor U1533 (N_1533,N_880,N_814);
nor U1534 (N_1534,N_1130,In_1100);
nand U1535 (N_1535,In_2345,In_2304);
nor U1536 (N_1536,In_1533,N_586);
nor U1537 (N_1537,In_1498,N_1079);
nor U1538 (N_1538,N_1148,N_648);
nor U1539 (N_1539,N_88,N_120);
nor U1540 (N_1540,N_973,In_863);
nand U1541 (N_1541,In_436,In_1862);
or U1542 (N_1542,N_1158,N_1190);
and U1543 (N_1543,In_2173,In_122);
nand U1544 (N_1544,N_875,N_951);
or U1545 (N_1545,In_2318,N_1231);
and U1546 (N_1546,N_1094,In_601);
nand U1547 (N_1547,N_1010,In_424);
nand U1548 (N_1548,N_684,N_570);
and U1549 (N_1549,N_569,In_345);
nand U1550 (N_1550,In_262,N_912);
nand U1551 (N_1551,N_833,N_1038);
or U1552 (N_1552,N_813,N_896);
nor U1553 (N_1553,N_770,In_1523);
nor U1554 (N_1554,In_2167,N_849);
nand U1555 (N_1555,N_812,In_1716);
nor U1556 (N_1556,N_1108,N_919);
and U1557 (N_1557,N_750,N_703);
nand U1558 (N_1558,N_536,N_92);
and U1559 (N_1559,N_888,N_1206);
nor U1560 (N_1560,N_1049,N_987);
and U1561 (N_1561,N_1102,N_860);
nor U1562 (N_1562,N_628,N_528);
or U1563 (N_1563,N_1085,In_2092);
or U1564 (N_1564,N_791,In_1098);
nor U1565 (N_1565,N_815,N_1054);
and U1566 (N_1566,N_745,In_404);
or U1567 (N_1567,N_494,N_848);
or U1568 (N_1568,N_1226,N_1141);
xor U1569 (N_1569,N_796,N_717);
nor U1570 (N_1570,In_1246,N_890);
and U1571 (N_1571,N_794,N_1007);
and U1572 (N_1572,In_1152,In_184);
and U1573 (N_1573,N_735,In_183);
nor U1574 (N_1574,N_58,N_756);
nand U1575 (N_1575,N_1234,In_191);
nand U1576 (N_1576,N_97,N_602);
nor U1577 (N_1577,N_806,N_744);
or U1578 (N_1578,In_2246,In_1766);
nand U1579 (N_1579,N_656,N_853);
or U1580 (N_1580,N_1167,N_668);
or U1581 (N_1581,N_949,N_57);
nor U1582 (N_1582,In_354,N_760);
or U1583 (N_1583,N_1065,In_2441);
xnor U1584 (N_1584,In_1534,N_594);
nor U1585 (N_1585,N_1156,In_2387);
nand U1586 (N_1586,In_18,In_1244);
or U1587 (N_1587,N_847,N_174);
and U1588 (N_1588,N_216,N_832);
or U1589 (N_1589,In_317,N_611);
or U1590 (N_1590,N_946,N_650);
nor U1591 (N_1591,In_765,N_710);
and U1592 (N_1592,In_1353,In_1708);
nor U1593 (N_1593,In_695,N_883);
and U1594 (N_1594,In_894,In_2390);
nor U1595 (N_1595,N_625,N_712);
xnor U1596 (N_1596,N_786,In_1250);
nor U1597 (N_1597,N_505,In_502);
nand U1598 (N_1598,N_490,N_748);
nor U1599 (N_1599,N_1037,N_612);
or U1600 (N_1600,In_290,In_2417);
and U1601 (N_1601,In_1432,N_818);
and U1602 (N_1602,N_41,In_2061);
nand U1603 (N_1603,In_1575,N_706);
and U1604 (N_1604,N_431,In_1401);
nand U1605 (N_1605,In_2020,N_324);
nand U1606 (N_1606,N_731,N_1004);
or U1607 (N_1607,N_975,N_596);
nor U1608 (N_1608,In_792,N_1022);
or U1609 (N_1609,In_752,N_111);
or U1610 (N_1610,N_659,N_1176);
or U1611 (N_1611,In_1596,In_1800);
nor U1612 (N_1612,In_1644,N_646);
or U1613 (N_1613,N_189,N_690);
nor U1614 (N_1614,N_941,N_426);
or U1615 (N_1615,N_782,N_1138);
nand U1616 (N_1616,In_249,N_1153);
nor U1617 (N_1617,In_264,In_2330);
or U1618 (N_1618,N_1044,In_2315);
or U1619 (N_1619,N_1199,N_998);
and U1620 (N_1620,In_1972,In_1739);
or U1621 (N_1621,N_439,In_157);
nand U1622 (N_1622,N_11,N_1144);
nand U1623 (N_1623,N_1126,N_679);
nand U1624 (N_1624,N_693,In_422);
nand U1625 (N_1625,N_1183,N_310);
or U1626 (N_1626,N_739,N_289);
and U1627 (N_1627,In_178,N_787);
nand U1628 (N_1628,In_211,N_40);
or U1629 (N_1629,In_627,N_1029);
nor U1630 (N_1630,N_708,N_260);
nor U1631 (N_1631,N_1035,N_1179);
xor U1632 (N_1632,In_2361,In_2327);
or U1633 (N_1633,N_330,In_551);
or U1634 (N_1634,N_171,In_1593);
nand U1635 (N_1635,N_1227,N_971);
xnor U1636 (N_1636,N_1091,N_309);
and U1637 (N_1637,N_722,In_1274);
and U1638 (N_1638,N_882,N_677);
nand U1639 (N_1639,N_905,In_1823);
or U1640 (N_1640,In_2112,In_1016);
or U1641 (N_1641,N_68,In_1211);
or U1642 (N_1642,N_1171,In_1215);
or U1643 (N_1643,N_620,N_994);
and U1644 (N_1644,In_1705,N_334);
or U1645 (N_1645,In_481,N_538);
nand U1646 (N_1646,In_1345,N_990);
or U1647 (N_1647,N_130,N_749);
or U1648 (N_1648,N_688,N_1077);
xnor U1649 (N_1649,In_880,In_599);
or U1650 (N_1650,In_2474,In_564);
or U1651 (N_1651,In_131,N_1129);
or U1652 (N_1652,N_682,In_72);
nor U1653 (N_1653,N_704,N_885);
nor U1654 (N_1654,N_817,In_1120);
nand U1655 (N_1655,In_299,N_19);
or U1656 (N_1656,N_1123,N_863);
and U1657 (N_1657,N_830,N_948);
nand U1658 (N_1658,N_1143,N_753);
nand U1659 (N_1659,N_986,N_563);
or U1660 (N_1660,In_844,N_774);
xor U1661 (N_1661,N_455,In_144);
nand U1662 (N_1662,N_1028,In_1749);
nor U1663 (N_1663,In_87,N_1074);
nand U1664 (N_1664,N_944,N_638);
nand U1665 (N_1665,N_653,N_1211);
nand U1666 (N_1666,N_661,In_308);
nor U1667 (N_1667,N_924,N_7);
and U1668 (N_1668,N_1219,N_1014);
nand U1669 (N_1669,In_1909,In_1381);
or U1670 (N_1670,N_1237,N_195);
and U1671 (N_1671,N_1142,N_771);
and U1672 (N_1672,N_175,N_777);
nand U1673 (N_1673,In_2292,N_48);
xnor U1674 (N_1674,N_1055,N_851);
and U1675 (N_1675,N_1205,In_402);
or U1676 (N_1676,N_610,In_376);
and U1677 (N_1677,N_1208,N_81);
xor U1678 (N_1678,In_2234,N_1193);
and U1679 (N_1679,N_202,In_1517);
or U1680 (N_1680,N_218,N_293);
nand U1681 (N_1681,N_702,N_694);
xor U1682 (N_1682,N_386,In_1650);
nand U1683 (N_1683,N_634,N_932);
nor U1684 (N_1684,N_115,N_1236);
nand U1685 (N_1685,In_2429,In_1177);
and U1686 (N_1686,In_954,N_1154);
or U1687 (N_1687,N_911,N_311);
nor U1688 (N_1688,N_867,N_1241);
and U1689 (N_1689,In_2184,In_2458);
or U1690 (N_1690,In_640,N_352);
and U1691 (N_1691,N_937,In_1202);
nand U1692 (N_1692,In_86,N_789);
nor U1693 (N_1693,N_936,In_2089);
and U1694 (N_1694,N_899,N_1232);
nor U1695 (N_1695,N_780,N_884);
and U1696 (N_1696,N_1178,N_669);
or U1697 (N_1697,In_1919,N_543);
nor U1698 (N_1698,N_652,In_570);
or U1699 (N_1699,N_1217,N_909);
nand U1700 (N_1700,In_294,In_1798);
nand U1701 (N_1701,N_834,In_116);
and U1702 (N_1702,N_831,N_928);
nor U1703 (N_1703,In_1407,N_479);
or U1704 (N_1704,In_2486,N_644);
nor U1705 (N_1705,N_4,N_1157);
or U1706 (N_1706,N_1005,N_1210);
nand U1707 (N_1707,In_1499,In_2409);
nand U1708 (N_1708,N_1135,N_980);
nor U1709 (N_1709,N_1220,N_686);
nand U1710 (N_1710,In_779,N_1173);
or U1711 (N_1711,N_1086,In_636);
and U1712 (N_1712,In_1943,N_636);
or U1713 (N_1713,N_978,N_1124);
nor U1714 (N_1714,In_293,In_2024);
nand U1715 (N_1715,In_1967,N_1084);
and U1716 (N_1716,In_154,N_1099);
and U1717 (N_1717,N_1116,N_1119);
nand U1718 (N_1718,N_1017,N_616);
or U1719 (N_1719,In_161,In_21);
or U1720 (N_1720,N_736,N_82);
and U1721 (N_1721,N_151,In_565);
nor U1722 (N_1722,N_1242,N_1224);
or U1723 (N_1723,In_524,N_626);
or U1724 (N_1724,N_816,N_79);
nand U1725 (N_1725,In_848,N_1185);
or U1726 (N_1726,N_1090,In_1609);
nor U1727 (N_1727,N_101,N_1093);
and U1728 (N_1728,In_1325,N_707);
xnor U1729 (N_1729,N_566,N_1201);
and U1730 (N_1730,In_977,N_1243);
or U1731 (N_1731,In_1921,N_220);
or U1732 (N_1732,N_788,In_812);
or U1733 (N_1733,N_752,N_915);
nand U1734 (N_1734,In_878,N_1212);
nand U1735 (N_1735,N_715,In_2371);
nor U1736 (N_1736,In_307,In_136);
and U1737 (N_1737,N_934,In_2280);
or U1738 (N_1738,In_1501,N_1207);
or U1739 (N_1739,N_1068,N_685);
and U1740 (N_1740,N_1198,N_1233);
and U1741 (N_1741,In_726,N_1043);
nand U1742 (N_1742,N_988,N_1109);
nand U1743 (N_1743,N_952,In_1454);
nand U1744 (N_1744,In_1806,N_904);
and U1745 (N_1745,In_688,N_698);
or U1746 (N_1746,N_829,N_790);
and U1747 (N_1747,N_74,N_1168);
nor U1748 (N_1748,N_663,N_861);
or U1749 (N_1749,In_703,In_92);
or U1750 (N_1750,N_784,N_1083);
or U1751 (N_1751,N_967,In_775);
nand U1752 (N_1752,N_907,In_2277);
and U1753 (N_1753,In_2190,N_641);
or U1754 (N_1754,In_699,N_1036);
nor U1755 (N_1755,N_416,In_2111);
nor U1756 (N_1756,N_935,In_816);
and U1757 (N_1757,N_734,N_631);
nor U1758 (N_1758,N_1003,In_198);
and U1759 (N_1759,In_663,N_378);
nor U1760 (N_1760,N_838,N_241);
nor U1761 (N_1761,N_509,N_931);
nor U1762 (N_1762,N_953,In_2312);
xor U1763 (N_1763,N_699,N_407);
or U1764 (N_1764,N_1177,N_737);
nand U1765 (N_1765,In_1360,N_992);
nor U1766 (N_1766,N_456,In_832);
xor U1767 (N_1767,In_340,N_732);
nor U1768 (N_1768,N_580,N_874);
or U1769 (N_1769,N_759,N_1200);
nor U1770 (N_1770,N_889,In_2490);
and U1771 (N_1771,N_1150,N_929);
and U1772 (N_1772,N_1072,N_112);
nor U1773 (N_1773,In_2257,N_329);
nor U1774 (N_1774,N_901,N_725);
nor U1775 (N_1775,N_1006,N_916);
nor U1776 (N_1776,In_1964,N_793);
and U1777 (N_1777,N_1082,In_1460);
xnor U1778 (N_1778,N_857,N_726);
nand U1779 (N_1779,In_1881,N_865);
nor U1780 (N_1780,N_1147,N_539);
or U1781 (N_1781,N_843,N_1186);
nand U1782 (N_1782,In_485,N_1103);
nor U1783 (N_1783,In_1720,N_540);
nand U1784 (N_1784,In_373,N_23);
nor U1785 (N_1785,N_1222,N_689);
and U1786 (N_1786,In_576,N_1246);
and U1787 (N_1787,In_383,N_939);
and U1788 (N_1788,N_862,N_729);
or U1789 (N_1789,In_1652,N_18);
or U1790 (N_1790,N_891,In_1086);
nand U1791 (N_1791,In_1904,N_242);
nor U1792 (N_1792,N_870,In_1854);
or U1793 (N_1793,N_799,N_114);
or U1794 (N_1794,N_984,N_1023);
or U1795 (N_1795,N_868,In_1917);
or U1796 (N_1796,N_877,N_942);
and U1797 (N_1797,N_1125,N_947);
nand U1798 (N_1798,N_1063,N_549);
nand U1799 (N_1799,N_1021,N_1230);
nor U1800 (N_1800,In_251,N_711);
and U1801 (N_1801,N_214,N_1020);
and U1802 (N_1802,N_983,N_963);
and U1803 (N_1803,In_681,N_629);
nand U1804 (N_1804,N_673,N_894);
and U1805 (N_1805,In_2103,In_970);
and U1806 (N_1806,In_1087,In_669);
nand U1807 (N_1807,N_614,N_741);
nor U1808 (N_1808,N_193,In_1408);
nor U1809 (N_1809,N_822,N_1045);
nand U1810 (N_1810,In_363,N_206);
xnor U1811 (N_1811,N_968,N_927);
nand U1812 (N_1812,N_808,In_1995);
nor U1813 (N_1813,In_1707,In_425);
nor U1814 (N_1814,N_1128,N_642);
and U1815 (N_1815,N_1137,In_804);
nand U1816 (N_1816,In_887,N_926);
nand U1817 (N_1817,N_902,N_317);
nor U1818 (N_1818,In_1748,N_385);
nor U1819 (N_1819,N_1184,In_1672);
and U1820 (N_1820,N_344,In_2159);
nor U1821 (N_1821,In_1390,N_989);
and U1822 (N_1822,In_1706,N_837);
xnor U1823 (N_1823,In_1312,N_1013);
or U1824 (N_1824,N_263,N_1056);
nand U1825 (N_1825,In_740,N_1048);
xnor U1826 (N_1826,N_1218,In_817);
and U1827 (N_1827,N_730,In_305);
xnor U1828 (N_1828,N_1110,N_667);
nor U1829 (N_1829,N_1088,N_1146);
nand U1830 (N_1830,In_721,N_1139);
nand U1831 (N_1831,N_850,N_1240);
and U1832 (N_1832,N_660,N_303);
nand U1833 (N_1833,In_1809,N_440);
nand U1834 (N_1834,In_811,In_1583);
and U1835 (N_1835,In_2351,N_881);
nor U1836 (N_1836,In_1974,N_231);
or U1837 (N_1837,N_1187,N_821);
nor U1838 (N_1838,In_2305,In_708);
nor U1839 (N_1839,In_1615,N_564);
nor U1840 (N_1840,In_2432,In_2464);
nand U1841 (N_1841,N_1151,In_2344);
or U1842 (N_1842,N_1140,N_700);
xor U1843 (N_1843,N_1149,In_1852);
and U1844 (N_1844,N_1089,N_1145);
or U1845 (N_1845,In_235,In_1344);
and U1846 (N_1846,In_2086,N_1115);
or U1847 (N_1847,N_665,N_36);
or U1848 (N_1848,In_2142,N_1051);
nor U1849 (N_1849,N_1229,N_763);
xnor U1850 (N_1850,N_1248,N_1040);
nand U1851 (N_1851,N_803,N_64);
or U1852 (N_1852,In_2128,In_2057);
nand U1853 (N_1853,N_176,N_167);
and U1854 (N_1854,N_910,N_914);
and U1855 (N_1855,N_224,N_500);
or U1856 (N_1856,N_778,N_643);
or U1857 (N_1857,In_998,In_833);
nor U1858 (N_1858,N_1152,In_1138);
or U1859 (N_1859,In_2400,N_1195);
and U1860 (N_1860,N_492,N_728);
xor U1861 (N_1861,N_250,N_1172);
nor U1862 (N_1862,N_676,In_1481);
and U1863 (N_1863,N_783,In_933);
or U1864 (N_1864,In_1168,N_743);
and U1865 (N_1865,N_1042,N_1078);
and U1866 (N_1866,N_738,N_956);
nor U1867 (N_1867,In_828,N_671);
nand U1868 (N_1868,In_723,N_776);
nand U1869 (N_1869,In_1140,N_1169);
xor U1870 (N_1870,N_452,N_1159);
and U1871 (N_1871,N_930,In_2469);
or U1872 (N_1872,N_1016,In_1580);
xor U1873 (N_1873,In_683,N_1069);
and U1874 (N_1874,N_1107,In_1017);
xnor U1875 (N_1875,N_1647,N_1434);
nor U1876 (N_1876,N_1449,N_1452);
or U1877 (N_1877,N_1429,N_1373);
nand U1878 (N_1878,N_1354,N_1704);
or U1879 (N_1879,N_1769,N_1637);
and U1880 (N_1880,N_1321,N_1722);
and U1881 (N_1881,N_1353,N_1765);
and U1882 (N_1882,N_1306,N_1817);
nor U1883 (N_1883,N_1280,N_1690);
and U1884 (N_1884,N_1663,N_1500);
and U1885 (N_1885,N_1796,N_1778);
or U1886 (N_1886,N_1518,N_1784);
and U1887 (N_1887,N_1813,N_1764);
or U1888 (N_1888,N_1274,N_1686);
nor U1889 (N_1889,N_1399,N_1498);
nand U1890 (N_1890,N_1506,N_1617);
nor U1891 (N_1891,N_1619,N_1517);
nand U1892 (N_1892,N_1466,N_1867);
nor U1893 (N_1893,N_1364,N_1341);
nor U1894 (N_1894,N_1393,N_1467);
or U1895 (N_1895,N_1851,N_1379);
nor U1896 (N_1896,N_1657,N_1456);
nor U1897 (N_1897,N_1572,N_1610);
nor U1898 (N_1898,N_1747,N_1795);
nand U1899 (N_1899,N_1872,N_1603);
nor U1900 (N_1900,N_1630,N_1433);
nor U1901 (N_1901,N_1329,N_1347);
and U1902 (N_1902,N_1675,N_1719);
and U1903 (N_1903,N_1601,N_1305);
nor U1904 (N_1904,N_1471,N_1385);
or U1905 (N_1905,N_1730,N_1563);
and U1906 (N_1906,N_1438,N_1258);
and U1907 (N_1907,N_1840,N_1622);
or U1908 (N_1908,N_1855,N_1411);
and U1909 (N_1909,N_1758,N_1299);
xor U1910 (N_1910,N_1343,N_1776);
nor U1911 (N_1911,N_1394,N_1502);
nand U1912 (N_1912,N_1609,N_1763);
xnor U1913 (N_1913,N_1391,N_1461);
nor U1914 (N_1914,N_1741,N_1279);
nand U1915 (N_1915,N_1549,N_1574);
and U1916 (N_1916,N_1799,N_1579);
and U1917 (N_1917,N_1465,N_1412);
and U1918 (N_1918,N_1281,N_1398);
nand U1919 (N_1919,N_1738,N_1616);
or U1920 (N_1920,N_1697,N_1486);
nand U1921 (N_1921,N_1863,N_1360);
or U1922 (N_1922,N_1265,N_1313);
or U1923 (N_1923,N_1535,N_1315);
or U1924 (N_1924,N_1590,N_1821);
nand U1925 (N_1925,N_1389,N_1636);
or U1926 (N_1926,N_1816,N_1402);
nor U1927 (N_1927,N_1284,N_1684);
or U1928 (N_1928,N_1372,N_1370);
nand U1929 (N_1929,N_1767,N_1832);
nand U1930 (N_1930,N_1665,N_1542);
nand U1931 (N_1931,N_1800,N_1621);
nor U1932 (N_1932,N_1294,N_1302);
nor U1933 (N_1933,N_1653,N_1287);
nand U1934 (N_1934,N_1290,N_1331);
or U1935 (N_1935,N_1860,N_1357);
and U1936 (N_1936,N_1253,N_1442);
nor U1937 (N_1937,N_1825,N_1654);
and U1938 (N_1938,N_1476,N_1462);
nand U1939 (N_1939,N_1252,N_1560);
xor U1940 (N_1940,N_1345,N_1333);
nor U1941 (N_1941,N_1569,N_1323);
and U1942 (N_1942,N_1628,N_1717);
nand U1943 (N_1943,N_1596,N_1599);
xnor U1944 (N_1944,N_1514,N_1858);
or U1945 (N_1945,N_1678,N_1640);
nor U1946 (N_1946,N_1849,N_1516);
and U1947 (N_1947,N_1519,N_1311);
xnor U1948 (N_1948,N_1735,N_1807);
nor U1949 (N_1949,N_1699,N_1631);
or U1950 (N_1950,N_1645,N_1511);
xnor U1951 (N_1951,N_1251,N_1723);
nor U1952 (N_1952,N_1854,N_1557);
nor U1953 (N_1953,N_1325,N_1777);
and U1954 (N_1954,N_1819,N_1862);
nor U1955 (N_1955,N_1541,N_1614);
xnor U1956 (N_1956,N_1576,N_1836);
nand U1957 (N_1957,N_1499,N_1413);
nand U1958 (N_1958,N_1760,N_1839);
nand U1959 (N_1959,N_1787,N_1696);
nand U1960 (N_1960,N_1419,N_1822);
nor U1961 (N_1961,N_1425,N_1676);
or U1962 (N_1962,N_1859,N_1446);
or U1963 (N_1963,N_1505,N_1629);
nor U1964 (N_1964,N_1841,N_1779);
nand U1965 (N_1965,N_1602,N_1304);
nor U1966 (N_1966,N_1856,N_1538);
nor U1967 (N_1967,N_1320,N_1406);
nor U1968 (N_1968,N_1369,N_1520);
nand U1969 (N_1969,N_1423,N_1529);
nor U1970 (N_1970,N_1527,N_1383);
nor U1971 (N_1971,N_1612,N_1532);
nand U1972 (N_1972,N_1454,N_1484);
nor U1973 (N_1973,N_1358,N_1706);
nor U1974 (N_1974,N_1559,N_1340);
nor U1975 (N_1975,N_1568,N_1754);
or U1976 (N_1976,N_1300,N_1613);
nand U1977 (N_1977,N_1432,N_1403);
nor U1978 (N_1978,N_1582,N_1427);
nand U1979 (N_1979,N_1288,N_1533);
nor U1980 (N_1980,N_1267,N_1750);
nand U1981 (N_1981,N_1753,N_1826);
and U1982 (N_1982,N_1550,N_1314);
or U1983 (N_1983,N_1838,N_1464);
or U1984 (N_1984,N_1384,N_1578);
nor U1985 (N_1985,N_1297,N_1873);
and U1986 (N_1986,N_1457,N_1459);
or U1987 (N_1987,N_1745,N_1426);
and U1988 (N_1988,N_1509,N_1565);
or U1989 (N_1989,N_1521,N_1319);
xor U1990 (N_1990,N_1495,N_1477);
nor U1991 (N_1991,N_1436,N_1618);
and U1992 (N_1992,N_1667,N_1556);
nor U1993 (N_1993,N_1482,N_1303);
or U1994 (N_1994,N_1539,N_1554);
or U1995 (N_1995,N_1573,N_1536);
nand U1996 (N_1996,N_1714,N_1277);
or U1997 (N_1997,N_1749,N_1605);
nand U1998 (N_1998,N_1386,N_1455);
and U1999 (N_1999,N_1285,N_1392);
nor U2000 (N_2000,N_1381,N_1338);
nand U2001 (N_2001,N_1720,N_1635);
or U2002 (N_2002,N_1448,N_1526);
nor U2003 (N_2003,N_1700,N_1830);
nor U2004 (N_2004,N_1847,N_1592);
and U2005 (N_2005,N_1673,N_1591);
or U2006 (N_2006,N_1707,N_1790);
nor U2007 (N_2007,N_1264,N_1395);
or U2008 (N_2008,N_1632,N_1296);
nor U2009 (N_2009,N_1301,N_1600);
nand U2010 (N_2010,N_1512,N_1701);
nand U2011 (N_2011,N_1365,N_1473);
nand U2012 (N_2012,N_1780,N_1694);
nand U2013 (N_2013,N_1334,N_1510);
and U2014 (N_2014,N_1724,N_1416);
nand U2015 (N_2015,N_1570,N_1848);
and U2016 (N_2016,N_1803,N_1857);
nand U2017 (N_2017,N_1740,N_1755);
nor U2018 (N_2018,N_1558,N_1275);
nor U2019 (N_2019,N_1668,N_1528);
nor U2020 (N_2020,N_1814,N_1674);
xor U2021 (N_2021,N_1792,N_1677);
or U2022 (N_2022,N_1481,N_1833);
nor U2023 (N_2023,N_1827,N_1713);
or U2024 (N_2024,N_1659,N_1418);
nor U2025 (N_2025,N_1414,N_1782);
or U2026 (N_2026,N_1260,N_1404);
nor U2027 (N_2027,N_1439,N_1344);
or U2028 (N_2028,N_1312,N_1501);
or U2029 (N_2029,N_1405,N_1781);
or U2030 (N_2030,N_1443,N_1843);
and U2031 (N_2031,N_1655,N_1831);
and U2032 (N_2032,N_1447,N_1829);
nor U2033 (N_2033,N_1837,N_1430);
nor U2034 (N_2034,N_1846,N_1768);
or U2035 (N_2035,N_1698,N_1742);
nor U2036 (N_2036,N_1437,N_1731);
nor U2037 (N_2037,N_1815,N_1259);
and U2038 (N_2038,N_1366,N_1567);
and U2039 (N_2039,N_1522,N_1598);
or U2040 (N_2040,N_1339,N_1480);
nor U2041 (N_2041,N_1546,N_1408);
nor U2042 (N_2042,N_1809,N_1588);
nand U2043 (N_2043,N_1734,N_1739);
xnor U2044 (N_2044,N_1773,N_1656);
nor U2045 (N_2045,N_1774,N_1692);
and U2046 (N_2046,N_1861,N_1607);
nor U2047 (N_2047,N_1363,N_1269);
nand U2048 (N_2048,N_1497,N_1871);
xnor U2049 (N_2049,N_1472,N_1322);
nand U2050 (N_2050,N_1270,N_1444);
and U2051 (N_2051,N_1548,N_1869);
and U2052 (N_2052,N_1615,N_1670);
or U2053 (N_2053,N_1593,N_1695);
and U2054 (N_2054,N_1804,N_1496);
nand U2055 (N_2055,N_1708,N_1828);
and U2056 (N_2056,N_1711,N_1718);
or U2057 (N_2057,N_1737,N_1382);
nand U2058 (N_2058,N_1691,N_1547);
nor U2059 (N_2059,N_1494,N_1337);
nor U2060 (N_2060,N_1682,N_1748);
and U2061 (N_2061,N_1865,N_1587);
or U2062 (N_2062,N_1431,N_1606);
and U2063 (N_2063,N_1652,N_1709);
nand U2064 (N_2064,N_1770,N_1633);
and U2065 (N_2065,N_1783,N_1661);
and U2066 (N_2066,N_1309,N_1488);
nand U2067 (N_2067,N_1440,N_1853);
nand U2068 (N_2068,N_1746,N_1672);
or U2069 (N_2069,N_1376,N_1664);
xor U2070 (N_2070,N_1255,N_1483);
nand U2071 (N_2071,N_1620,N_1283);
xor U2072 (N_2072,N_1660,N_1864);
or U2073 (N_2073,N_1318,N_1651);
or U2074 (N_2074,N_1292,N_1254);
xnor U2075 (N_2075,N_1543,N_1451);
nor U2076 (N_2076,N_1324,N_1789);
nand U2077 (N_2077,N_1608,N_1555);
xor U2078 (N_2078,N_1375,N_1504);
or U2079 (N_2079,N_1327,N_1643);
or U2080 (N_2080,N_1348,N_1401);
nand U2081 (N_2081,N_1400,N_1797);
or U2082 (N_2082,N_1727,N_1415);
and U2083 (N_2083,N_1646,N_1638);
and U2084 (N_2084,N_1421,N_1371);
nand U2085 (N_2085,N_1293,N_1842);
nor U2086 (N_2086,N_1396,N_1705);
xor U2087 (N_2087,N_1263,N_1295);
or U2088 (N_2088,N_1458,N_1352);
nor U2089 (N_2089,N_1564,N_1537);
nand U2090 (N_2090,N_1575,N_1553);
or U2091 (N_2091,N_1328,N_1531);
or U2092 (N_2092,N_1649,N_1766);
nand U2093 (N_2093,N_1688,N_1387);
nor U2094 (N_2094,N_1487,N_1361);
nor U2095 (N_2095,N_1489,N_1650);
or U2096 (N_2096,N_1810,N_1725);
and U2097 (N_2097,N_1390,N_1793);
nand U2098 (N_2098,N_1420,N_1798);
xnor U2099 (N_2099,N_1586,N_1335);
and U2100 (N_2100,N_1491,N_1669);
and U2101 (N_2101,N_1681,N_1756);
and U2102 (N_2102,N_1307,N_1627);
nand U2103 (N_2103,N_1479,N_1485);
or U2104 (N_2104,N_1445,N_1762);
nand U2105 (N_2105,N_1515,N_1641);
nand U2106 (N_2106,N_1351,N_1424);
and U2107 (N_2107,N_1785,N_1332);
nor U2108 (N_2108,N_1256,N_1662);
nor U2109 (N_2109,N_1571,N_1470);
or U2110 (N_2110,N_1410,N_1823);
nand U2111 (N_2111,N_1752,N_1595);
nor U2112 (N_2112,N_1759,N_1751);
and U2113 (N_2113,N_1820,N_1671);
or U2114 (N_2114,N_1503,N_1453);
nand U2115 (N_2115,N_1729,N_1693);
or U2116 (N_2116,N_1468,N_1566);
nand U2117 (N_2117,N_1786,N_1604);
nor U2118 (N_2118,N_1811,N_1577);
xor U2119 (N_2119,N_1583,N_1870);
and U2120 (N_2120,N_1703,N_1644);
or U2121 (N_2121,N_1530,N_1584);
nand U2122 (N_2122,N_1624,N_1262);
and U2123 (N_2123,N_1475,N_1791);
or U2124 (N_2124,N_1844,N_1733);
and U2125 (N_2125,N_1544,N_1374);
xnor U2126 (N_2126,N_1278,N_1625);
nor U2127 (N_2127,N_1450,N_1525);
nand U2128 (N_2128,N_1562,N_1580);
or U2129 (N_2129,N_1585,N_1702);
or U2130 (N_2130,N_1802,N_1469);
nor U2131 (N_2131,N_1824,N_1812);
or U2132 (N_2132,N_1732,N_1639);
nand U2133 (N_2133,N_1289,N_1409);
nor U2134 (N_2134,N_1623,N_1428);
and U2135 (N_2135,N_1524,N_1845);
or U2136 (N_2136,N_1378,N_1310);
nand U2137 (N_2137,N_1552,N_1397);
and U2138 (N_2138,N_1710,N_1545);
nor U2139 (N_2139,N_1866,N_1597);
and U2140 (N_2140,N_1634,N_1407);
and U2141 (N_2141,N_1250,N_1523);
or U2142 (N_2142,N_1689,N_1794);
nand U2143 (N_2143,N_1330,N_1282);
nand U2144 (N_2144,N_1772,N_1658);
or U2145 (N_2145,N_1771,N_1367);
or U2146 (N_2146,N_1493,N_1463);
nand U2147 (N_2147,N_1272,N_1744);
nand U2148 (N_2148,N_1336,N_1490);
and U2149 (N_2149,N_1492,N_1271);
and U2150 (N_2150,N_1346,N_1757);
or U2151 (N_2151,N_1362,N_1551);
nand U2152 (N_2152,N_1680,N_1326);
or U2153 (N_2153,N_1868,N_1743);
nand U2154 (N_2154,N_1350,N_1441);
nand U2155 (N_2155,N_1355,N_1850);
and U2156 (N_2156,N_1728,N_1721);
or U2157 (N_2157,N_1835,N_1268);
xor U2158 (N_2158,N_1417,N_1377);
nor U2159 (N_2159,N_1257,N_1261);
nor U2160 (N_2160,N_1666,N_1648);
nor U2161 (N_2161,N_1460,N_1715);
xnor U2162 (N_2162,N_1380,N_1594);
nand U2163 (N_2163,N_1298,N_1736);
xnor U2164 (N_2164,N_1507,N_1712);
nor U2165 (N_2165,N_1508,N_1801);
or U2166 (N_2166,N_1775,N_1818);
nor U2167 (N_2167,N_1356,N_1852);
xnor U2168 (N_2168,N_1581,N_1534);
and U2169 (N_2169,N_1683,N_1716);
nand U2170 (N_2170,N_1834,N_1679);
xnor U2171 (N_2171,N_1286,N_1874);
and U2172 (N_2172,N_1726,N_1266);
and U2173 (N_2173,N_1642,N_1273);
or U2174 (N_2174,N_1422,N_1308);
nor U2175 (N_2175,N_1388,N_1806);
and U2176 (N_2176,N_1291,N_1589);
or U2177 (N_2177,N_1435,N_1540);
nor U2178 (N_2178,N_1808,N_1788);
nand U2179 (N_2179,N_1349,N_1359);
or U2180 (N_2180,N_1342,N_1316);
or U2181 (N_2181,N_1687,N_1368);
or U2182 (N_2182,N_1478,N_1317);
nor U2183 (N_2183,N_1611,N_1805);
nand U2184 (N_2184,N_1513,N_1561);
nor U2185 (N_2185,N_1685,N_1276);
and U2186 (N_2186,N_1626,N_1761);
and U2187 (N_2187,N_1474,N_1325);
nand U2188 (N_2188,N_1420,N_1414);
or U2189 (N_2189,N_1872,N_1340);
nor U2190 (N_2190,N_1663,N_1354);
nor U2191 (N_2191,N_1507,N_1721);
nand U2192 (N_2192,N_1344,N_1409);
nand U2193 (N_2193,N_1425,N_1496);
nand U2194 (N_2194,N_1477,N_1398);
and U2195 (N_2195,N_1780,N_1727);
nor U2196 (N_2196,N_1822,N_1766);
and U2197 (N_2197,N_1534,N_1800);
xor U2198 (N_2198,N_1594,N_1663);
nor U2199 (N_2199,N_1428,N_1447);
nor U2200 (N_2200,N_1701,N_1303);
nand U2201 (N_2201,N_1768,N_1785);
nor U2202 (N_2202,N_1770,N_1307);
nand U2203 (N_2203,N_1622,N_1554);
xnor U2204 (N_2204,N_1788,N_1810);
or U2205 (N_2205,N_1666,N_1785);
nand U2206 (N_2206,N_1571,N_1393);
or U2207 (N_2207,N_1548,N_1525);
and U2208 (N_2208,N_1604,N_1846);
nand U2209 (N_2209,N_1671,N_1768);
and U2210 (N_2210,N_1640,N_1772);
or U2211 (N_2211,N_1822,N_1541);
nand U2212 (N_2212,N_1299,N_1794);
nand U2213 (N_2213,N_1394,N_1855);
xnor U2214 (N_2214,N_1456,N_1505);
nand U2215 (N_2215,N_1318,N_1789);
and U2216 (N_2216,N_1402,N_1251);
nor U2217 (N_2217,N_1578,N_1422);
and U2218 (N_2218,N_1485,N_1756);
or U2219 (N_2219,N_1642,N_1303);
xnor U2220 (N_2220,N_1511,N_1477);
or U2221 (N_2221,N_1432,N_1397);
nand U2222 (N_2222,N_1451,N_1840);
or U2223 (N_2223,N_1743,N_1698);
or U2224 (N_2224,N_1510,N_1627);
nor U2225 (N_2225,N_1376,N_1762);
and U2226 (N_2226,N_1628,N_1678);
nand U2227 (N_2227,N_1715,N_1846);
nor U2228 (N_2228,N_1445,N_1505);
xor U2229 (N_2229,N_1304,N_1824);
xnor U2230 (N_2230,N_1371,N_1847);
or U2231 (N_2231,N_1320,N_1643);
xor U2232 (N_2232,N_1317,N_1551);
nand U2233 (N_2233,N_1609,N_1702);
nand U2234 (N_2234,N_1612,N_1707);
xnor U2235 (N_2235,N_1817,N_1292);
xor U2236 (N_2236,N_1363,N_1848);
nor U2237 (N_2237,N_1289,N_1450);
and U2238 (N_2238,N_1431,N_1449);
or U2239 (N_2239,N_1669,N_1375);
xnor U2240 (N_2240,N_1814,N_1438);
nand U2241 (N_2241,N_1760,N_1271);
or U2242 (N_2242,N_1516,N_1831);
xor U2243 (N_2243,N_1533,N_1297);
nor U2244 (N_2244,N_1627,N_1509);
or U2245 (N_2245,N_1816,N_1448);
and U2246 (N_2246,N_1519,N_1671);
nand U2247 (N_2247,N_1388,N_1835);
or U2248 (N_2248,N_1703,N_1285);
nand U2249 (N_2249,N_1518,N_1296);
xor U2250 (N_2250,N_1564,N_1595);
xor U2251 (N_2251,N_1689,N_1588);
xnor U2252 (N_2252,N_1503,N_1756);
nand U2253 (N_2253,N_1647,N_1251);
nand U2254 (N_2254,N_1713,N_1603);
and U2255 (N_2255,N_1604,N_1663);
xnor U2256 (N_2256,N_1873,N_1652);
xnor U2257 (N_2257,N_1531,N_1475);
or U2258 (N_2258,N_1409,N_1438);
nand U2259 (N_2259,N_1802,N_1288);
and U2260 (N_2260,N_1536,N_1438);
nor U2261 (N_2261,N_1700,N_1363);
or U2262 (N_2262,N_1857,N_1779);
nor U2263 (N_2263,N_1630,N_1704);
nand U2264 (N_2264,N_1731,N_1529);
xor U2265 (N_2265,N_1584,N_1324);
nand U2266 (N_2266,N_1735,N_1378);
nor U2267 (N_2267,N_1783,N_1871);
nand U2268 (N_2268,N_1451,N_1767);
and U2269 (N_2269,N_1786,N_1278);
or U2270 (N_2270,N_1702,N_1763);
and U2271 (N_2271,N_1365,N_1335);
and U2272 (N_2272,N_1555,N_1282);
nand U2273 (N_2273,N_1541,N_1701);
nor U2274 (N_2274,N_1419,N_1815);
xnor U2275 (N_2275,N_1757,N_1811);
nor U2276 (N_2276,N_1585,N_1569);
xor U2277 (N_2277,N_1280,N_1742);
nor U2278 (N_2278,N_1774,N_1281);
or U2279 (N_2279,N_1567,N_1647);
or U2280 (N_2280,N_1521,N_1330);
nor U2281 (N_2281,N_1674,N_1330);
nand U2282 (N_2282,N_1741,N_1362);
nand U2283 (N_2283,N_1720,N_1398);
nor U2284 (N_2284,N_1457,N_1403);
nor U2285 (N_2285,N_1304,N_1325);
nor U2286 (N_2286,N_1747,N_1282);
nor U2287 (N_2287,N_1430,N_1757);
nor U2288 (N_2288,N_1580,N_1832);
or U2289 (N_2289,N_1841,N_1469);
or U2290 (N_2290,N_1719,N_1417);
xnor U2291 (N_2291,N_1302,N_1507);
nand U2292 (N_2292,N_1783,N_1653);
or U2293 (N_2293,N_1824,N_1600);
or U2294 (N_2294,N_1853,N_1561);
nand U2295 (N_2295,N_1421,N_1395);
or U2296 (N_2296,N_1336,N_1657);
or U2297 (N_2297,N_1786,N_1533);
nand U2298 (N_2298,N_1521,N_1614);
and U2299 (N_2299,N_1689,N_1614);
nor U2300 (N_2300,N_1426,N_1640);
and U2301 (N_2301,N_1470,N_1671);
and U2302 (N_2302,N_1383,N_1580);
xor U2303 (N_2303,N_1827,N_1637);
and U2304 (N_2304,N_1792,N_1580);
nor U2305 (N_2305,N_1567,N_1664);
and U2306 (N_2306,N_1711,N_1576);
nand U2307 (N_2307,N_1743,N_1641);
nor U2308 (N_2308,N_1368,N_1804);
or U2309 (N_2309,N_1744,N_1335);
nor U2310 (N_2310,N_1388,N_1620);
and U2311 (N_2311,N_1749,N_1412);
nor U2312 (N_2312,N_1591,N_1548);
nor U2313 (N_2313,N_1481,N_1327);
or U2314 (N_2314,N_1563,N_1348);
xnor U2315 (N_2315,N_1453,N_1282);
or U2316 (N_2316,N_1471,N_1420);
nor U2317 (N_2317,N_1578,N_1457);
or U2318 (N_2318,N_1738,N_1338);
nor U2319 (N_2319,N_1443,N_1300);
nand U2320 (N_2320,N_1652,N_1312);
or U2321 (N_2321,N_1679,N_1315);
or U2322 (N_2322,N_1729,N_1759);
nand U2323 (N_2323,N_1728,N_1873);
nor U2324 (N_2324,N_1537,N_1663);
nand U2325 (N_2325,N_1646,N_1773);
xor U2326 (N_2326,N_1505,N_1346);
and U2327 (N_2327,N_1423,N_1874);
and U2328 (N_2328,N_1718,N_1734);
nor U2329 (N_2329,N_1777,N_1369);
or U2330 (N_2330,N_1358,N_1695);
or U2331 (N_2331,N_1600,N_1353);
or U2332 (N_2332,N_1360,N_1796);
or U2333 (N_2333,N_1476,N_1449);
xnor U2334 (N_2334,N_1775,N_1667);
and U2335 (N_2335,N_1833,N_1487);
nor U2336 (N_2336,N_1845,N_1364);
or U2337 (N_2337,N_1567,N_1848);
or U2338 (N_2338,N_1334,N_1633);
xnor U2339 (N_2339,N_1846,N_1640);
nand U2340 (N_2340,N_1773,N_1336);
and U2341 (N_2341,N_1784,N_1715);
xor U2342 (N_2342,N_1873,N_1732);
nand U2343 (N_2343,N_1718,N_1539);
or U2344 (N_2344,N_1612,N_1295);
nor U2345 (N_2345,N_1340,N_1653);
nand U2346 (N_2346,N_1664,N_1489);
or U2347 (N_2347,N_1691,N_1634);
and U2348 (N_2348,N_1363,N_1756);
nand U2349 (N_2349,N_1716,N_1413);
nand U2350 (N_2350,N_1748,N_1678);
xor U2351 (N_2351,N_1715,N_1324);
or U2352 (N_2352,N_1786,N_1705);
nand U2353 (N_2353,N_1400,N_1714);
or U2354 (N_2354,N_1389,N_1628);
or U2355 (N_2355,N_1411,N_1665);
and U2356 (N_2356,N_1733,N_1465);
and U2357 (N_2357,N_1433,N_1621);
or U2358 (N_2358,N_1866,N_1484);
or U2359 (N_2359,N_1649,N_1555);
xor U2360 (N_2360,N_1616,N_1587);
nand U2361 (N_2361,N_1858,N_1469);
or U2362 (N_2362,N_1702,N_1446);
or U2363 (N_2363,N_1633,N_1544);
nand U2364 (N_2364,N_1465,N_1267);
nand U2365 (N_2365,N_1773,N_1866);
xor U2366 (N_2366,N_1800,N_1374);
nand U2367 (N_2367,N_1509,N_1576);
nor U2368 (N_2368,N_1387,N_1765);
xnor U2369 (N_2369,N_1382,N_1436);
xor U2370 (N_2370,N_1536,N_1687);
nor U2371 (N_2371,N_1616,N_1678);
and U2372 (N_2372,N_1305,N_1309);
xor U2373 (N_2373,N_1562,N_1685);
and U2374 (N_2374,N_1581,N_1306);
nand U2375 (N_2375,N_1865,N_1548);
nand U2376 (N_2376,N_1363,N_1598);
nor U2377 (N_2377,N_1869,N_1543);
and U2378 (N_2378,N_1649,N_1552);
xor U2379 (N_2379,N_1324,N_1370);
nand U2380 (N_2380,N_1773,N_1643);
or U2381 (N_2381,N_1300,N_1432);
and U2382 (N_2382,N_1366,N_1289);
nand U2383 (N_2383,N_1322,N_1744);
nand U2384 (N_2384,N_1294,N_1792);
or U2385 (N_2385,N_1781,N_1666);
nor U2386 (N_2386,N_1760,N_1862);
xnor U2387 (N_2387,N_1539,N_1828);
nor U2388 (N_2388,N_1824,N_1563);
and U2389 (N_2389,N_1856,N_1584);
xor U2390 (N_2390,N_1617,N_1599);
nor U2391 (N_2391,N_1547,N_1718);
nor U2392 (N_2392,N_1612,N_1806);
nor U2393 (N_2393,N_1617,N_1521);
xor U2394 (N_2394,N_1872,N_1765);
and U2395 (N_2395,N_1639,N_1641);
nand U2396 (N_2396,N_1822,N_1643);
nand U2397 (N_2397,N_1791,N_1349);
nand U2398 (N_2398,N_1689,N_1849);
or U2399 (N_2399,N_1690,N_1761);
nand U2400 (N_2400,N_1669,N_1444);
and U2401 (N_2401,N_1582,N_1332);
nor U2402 (N_2402,N_1770,N_1641);
nand U2403 (N_2403,N_1289,N_1621);
nor U2404 (N_2404,N_1385,N_1722);
nor U2405 (N_2405,N_1749,N_1423);
nor U2406 (N_2406,N_1295,N_1783);
and U2407 (N_2407,N_1453,N_1308);
and U2408 (N_2408,N_1766,N_1485);
or U2409 (N_2409,N_1627,N_1622);
and U2410 (N_2410,N_1648,N_1816);
or U2411 (N_2411,N_1301,N_1511);
nand U2412 (N_2412,N_1787,N_1610);
and U2413 (N_2413,N_1826,N_1502);
nor U2414 (N_2414,N_1454,N_1677);
and U2415 (N_2415,N_1274,N_1637);
nor U2416 (N_2416,N_1263,N_1602);
nand U2417 (N_2417,N_1272,N_1307);
or U2418 (N_2418,N_1579,N_1350);
or U2419 (N_2419,N_1772,N_1869);
or U2420 (N_2420,N_1640,N_1767);
nand U2421 (N_2421,N_1338,N_1635);
or U2422 (N_2422,N_1641,N_1702);
xnor U2423 (N_2423,N_1633,N_1335);
or U2424 (N_2424,N_1863,N_1735);
and U2425 (N_2425,N_1467,N_1511);
and U2426 (N_2426,N_1674,N_1307);
or U2427 (N_2427,N_1500,N_1820);
nor U2428 (N_2428,N_1490,N_1398);
and U2429 (N_2429,N_1703,N_1749);
and U2430 (N_2430,N_1592,N_1763);
xor U2431 (N_2431,N_1456,N_1850);
nand U2432 (N_2432,N_1315,N_1469);
nor U2433 (N_2433,N_1845,N_1293);
xnor U2434 (N_2434,N_1645,N_1380);
nand U2435 (N_2435,N_1581,N_1566);
nor U2436 (N_2436,N_1634,N_1859);
or U2437 (N_2437,N_1407,N_1815);
xor U2438 (N_2438,N_1334,N_1752);
nand U2439 (N_2439,N_1573,N_1563);
nor U2440 (N_2440,N_1788,N_1787);
and U2441 (N_2441,N_1434,N_1371);
xor U2442 (N_2442,N_1842,N_1410);
and U2443 (N_2443,N_1270,N_1321);
and U2444 (N_2444,N_1503,N_1764);
nor U2445 (N_2445,N_1660,N_1604);
nand U2446 (N_2446,N_1804,N_1325);
or U2447 (N_2447,N_1854,N_1341);
or U2448 (N_2448,N_1298,N_1622);
or U2449 (N_2449,N_1861,N_1293);
nor U2450 (N_2450,N_1453,N_1644);
or U2451 (N_2451,N_1426,N_1769);
or U2452 (N_2452,N_1749,N_1574);
nand U2453 (N_2453,N_1520,N_1375);
or U2454 (N_2454,N_1539,N_1630);
nand U2455 (N_2455,N_1704,N_1688);
nor U2456 (N_2456,N_1493,N_1278);
nor U2457 (N_2457,N_1808,N_1728);
or U2458 (N_2458,N_1821,N_1772);
nor U2459 (N_2459,N_1576,N_1464);
or U2460 (N_2460,N_1614,N_1574);
and U2461 (N_2461,N_1713,N_1291);
and U2462 (N_2462,N_1423,N_1426);
and U2463 (N_2463,N_1834,N_1394);
nor U2464 (N_2464,N_1861,N_1554);
nand U2465 (N_2465,N_1573,N_1600);
or U2466 (N_2466,N_1811,N_1716);
and U2467 (N_2467,N_1494,N_1327);
nand U2468 (N_2468,N_1632,N_1404);
nand U2469 (N_2469,N_1789,N_1555);
nand U2470 (N_2470,N_1340,N_1284);
and U2471 (N_2471,N_1441,N_1707);
nand U2472 (N_2472,N_1626,N_1335);
and U2473 (N_2473,N_1565,N_1815);
or U2474 (N_2474,N_1474,N_1744);
nand U2475 (N_2475,N_1425,N_1455);
xnor U2476 (N_2476,N_1295,N_1619);
nand U2477 (N_2477,N_1548,N_1620);
nand U2478 (N_2478,N_1607,N_1390);
and U2479 (N_2479,N_1753,N_1635);
xnor U2480 (N_2480,N_1522,N_1709);
nor U2481 (N_2481,N_1701,N_1827);
nor U2482 (N_2482,N_1650,N_1690);
nor U2483 (N_2483,N_1563,N_1798);
nand U2484 (N_2484,N_1264,N_1363);
or U2485 (N_2485,N_1609,N_1804);
or U2486 (N_2486,N_1676,N_1464);
nand U2487 (N_2487,N_1689,N_1637);
and U2488 (N_2488,N_1353,N_1735);
and U2489 (N_2489,N_1288,N_1607);
nand U2490 (N_2490,N_1386,N_1730);
and U2491 (N_2491,N_1453,N_1694);
or U2492 (N_2492,N_1355,N_1845);
nand U2493 (N_2493,N_1692,N_1464);
nor U2494 (N_2494,N_1407,N_1816);
or U2495 (N_2495,N_1765,N_1519);
or U2496 (N_2496,N_1335,N_1409);
nor U2497 (N_2497,N_1695,N_1264);
or U2498 (N_2498,N_1331,N_1340);
and U2499 (N_2499,N_1773,N_1521);
nand U2500 (N_2500,N_1910,N_2397);
nand U2501 (N_2501,N_1976,N_2423);
and U2502 (N_2502,N_1915,N_2055);
or U2503 (N_2503,N_2030,N_2283);
and U2504 (N_2504,N_2332,N_2226);
or U2505 (N_2505,N_2150,N_2118);
nand U2506 (N_2506,N_2077,N_2378);
and U2507 (N_2507,N_2348,N_2167);
and U2508 (N_2508,N_1986,N_2040);
and U2509 (N_2509,N_2379,N_2024);
nor U2510 (N_2510,N_2087,N_2488);
and U2511 (N_2511,N_2170,N_2486);
and U2512 (N_2512,N_2002,N_2009);
nor U2513 (N_2513,N_2103,N_1877);
xor U2514 (N_2514,N_2176,N_1970);
xnor U2515 (N_2515,N_2490,N_1999);
or U2516 (N_2516,N_2480,N_2147);
or U2517 (N_2517,N_2338,N_2257);
xor U2518 (N_2518,N_2126,N_2107);
nor U2519 (N_2519,N_2327,N_2006);
and U2520 (N_2520,N_2148,N_2431);
nor U2521 (N_2521,N_2000,N_1901);
or U2522 (N_2522,N_2154,N_2161);
nand U2523 (N_2523,N_2197,N_2031);
and U2524 (N_2524,N_2068,N_2230);
or U2525 (N_2525,N_2325,N_2191);
nor U2526 (N_2526,N_2497,N_2174);
or U2527 (N_2527,N_2053,N_2375);
or U2528 (N_2528,N_2393,N_2437);
and U2529 (N_2529,N_1994,N_1929);
and U2530 (N_2530,N_1920,N_2198);
nand U2531 (N_2531,N_2452,N_2285);
nor U2532 (N_2532,N_2487,N_2043);
nand U2533 (N_2533,N_1971,N_2451);
nand U2534 (N_2534,N_2259,N_2020);
xor U2535 (N_2535,N_1905,N_2182);
or U2536 (N_2536,N_1947,N_1963);
or U2537 (N_2537,N_2036,N_2240);
nand U2538 (N_2538,N_2410,N_1941);
or U2539 (N_2539,N_2404,N_2304);
nor U2540 (N_2540,N_2474,N_2142);
nand U2541 (N_2541,N_1933,N_2398);
nand U2542 (N_2542,N_2218,N_1890);
xnor U2543 (N_2543,N_2234,N_2162);
nand U2544 (N_2544,N_2268,N_2491);
xor U2545 (N_2545,N_2199,N_2008);
or U2546 (N_2546,N_2242,N_2172);
xor U2547 (N_2547,N_2387,N_2323);
nor U2548 (N_2548,N_2157,N_1892);
nand U2549 (N_2549,N_2428,N_2231);
and U2550 (N_2550,N_1965,N_1880);
or U2551 (N_2551,N_2391,N_2111);
and U2552 (N_2552,N_2448,N_1896);
nand U2553 (N_2553,N_2116,N_2371);
or U2554 (N_2554,N_2493,N_2467);
and U2555 (N_2555,N_2311,N_2244);
and U2556 (N_2556,N_2331,N_2214);
and U2557 (N_2557,N_2012,N_1876);
nand U2558 (N_2558,N_2134,N_2196);
nor U2559 (N_2559,N_1930,N_2415);
nand U2560 (N_2560,N_2440,N_2295);
nand U2561 (N_2561,N_2365,N_1995);
and U2562 (N_2562,N_2388,N_2027);
or U2563 (N_2563,N_2035,N_1949);
and U2564 (N_2564,N_1902,N_2194);
nand U2565 (N_2565,N_2237,N_2446);
nor U2566 (N_2566,N_2402,N_1875);
nand U2567 (N_2567,N_2101,N_2334);
or U2568 (N_2568,N_2203,N_2289);
nand U2569 (N_2569,N_2168,N_2224);
xor U2570 (N_2570,N_2372,N_1962);
nand U2571 (N_2571,N_2245,N_1980);
and U2572 (N_2572,N_2290,N_2427);
nor U2573 (N_2573,N_1990,N_2460);
or U2574 (N_2574,N_1975,N_2100);
nand U2575 (N_2575,N_1900,N_2344);
nor U2576 (N_2576,N_2314,N_2337);
nor U2577 (N_2577,N_2125,N_2355);
nor U2578 (N_2578,N_2269,N_1934);
nor U2579 (N_2579,N_2246,N_2110);
and U2580 (N_2580,N_2457,N_1881);
nor U2581 (N_2581,N_2347,N_2065);
nand U2582 (N_2582,N_2275,N_2319);
and U2583 (N_2583,N_2112,N_2128);
or U2584 (N_2584,N_2156,N_2106);
nand U2585 (N_2585,N_2321,N_2376);
nand U2586 (N_2586,N_2326,N_1908);
nand U2587 (N_2587,N_2345,N_2294);
xnor U2588 (N_2588,N_1909,N_1993);
and U2589 (N_2589,N_1959,N_1984);
nor U2590 (N_2590,N_2408,N_1950);
and U2591 (N_2591,N_2207,N_2265);
nand U2592 (N_2592,N_2281,N_2466);
nor U2593 (N_2593,N_2438,N_2233);
nor U2594 (N_2594,N_2351,N_1985);
nand U2595 (N_2595,N_2318,N_2016);
nand U2596 (N_2596,N_2113,N_2146);
nand U2597 (N_2597,N_1907,N_2076);
xnor U2598 (N_2598,N_2322,N_2114);
and U2599 (N_2599,N_2071,N_2310);
nor U2600 (N_2600,N_2444,N_2179);
or U2601 (N_2601,N_2346,N_2132);
nand U2602 (N_2602,N_2336,N_2091);
nor U2603 (N_2603,N_2343,N_2014);
and U2604 (N_2604,N_2436,N_2165);
nand U2605 (N_2605,N_2274,N_2001);
nand U2606 (N_2606,N_1893,N_2028);
nor U2607 (N_2607,N_1987,N_2047);
nor U2608 (N_2608,N_2416,N_2382);
xor U2609 (N_2609,N_1997,N_2117);
nand U2610 (N_2610,N_1996,N_1919);
nand U2611 (N_2611,N_2256,N_1939);
nand U2612 (N_2612,N_2241,N_2190);
or U2613 (N_2613,N_2164,N_1887);
or U2614 (N_2614,N_1917,N_2258);
xor U2615 (N_2615,N_2038,N_1938);
or U2616 (N_2616,N_2477,N_2026);
xnor U2617 (N_2617,N_2039,N_2158);
and U2618 (N_2618,N_2227,N_1982);
or U2619 (N_2619,N_2048,N_2229);
or U2620 (N_2620,N_2478,N_2263);
nor U2621 (N_2621,N_2064,N_2249);
nand U2622 (N_2622,N_2042,N_2209);
or U2623 (N_2623,N_1911,N_1957);
xor U2624 (N_2624,N_2472,N_1989);
xnor U2625 (N_2625,N_2187,N_2456);
nor U2626 (N_2626,N_2296,N_1977);
nor U2627 (N_2627,N_1958,N_2449);
xor U2628 (N_2628,N_2186,N_2359);
or U2629 (N_2629,N_1953,N_2354);
and U2630 (N_2630,N_1967,N_2088);
nand U2631 (N_2631,N_2280,N_2080);
nand U2632 (N_2632,N_2284,N_2075);
and U2633 (N_2633,N_2481,N_1912);
nor U2634 (N_2634,N_2181,N_2183);
nor U2635 (N_2635,N_2369,N_2219);
nor U2636 (N_2636,N_2211,N_2023);
and U2637 (N_2637,N_2094,N_2430);
nor U2638 (N_2638,N_2056,N_2352);
xnor U2639 (N_2639,N_2368,N_1918);
nand U2640 (N_2640,N_2173,N_2115);
and U2641 (N_2641,N_2377,N_2180);
xnor U2642 (N_2642,N_2407,N_2098);
xnor U2643 (N_2643,N_2145,N_2300);
nor U2644 (N_2644,N_1886,N_2037);
or U2645 (N_2645,N_1926,N_2350);
and U2646 (N_2646,N_1937,N_2122);
nor U2647 (N_2647,N_1974,N_2262);
nor U2648 (N_2648,N_1894,N_2223);
or U2649 (N_2649,N_2342,N_2089);
nor U2650 (N_2650,N_2271,N_2130);
nor U2651 (N_2651,N_2386,N_2413);
nor U2652 (N_2652,N_1966,N_1906);
or U2653 (N_2653,N_2086,N_2069);
nor U2654 (N_2654,N_2137,N_2252);
xor U2655 (N_2655,N_1914,N_2072);
xnor U2656 (N_2656,N_2066,N_2489);
and U2657 (N_2657,N_1882,N_2235);
nand U2658 (N_2658,N_2339,N_2215);
and U2659 (N_2659,N_2090,N_2054);
and U2660 (N_2660,N_2236,N_2034);
and U2661 (N_2661,N_2140,N_2019);
nand U2662 (N_2662,N_1992,N_2239);
or U2663 (N_2663,N_2044,N_2160);
nand U2664 (N_2664,N_2193,N_2045);
and U2665 (N_2665,N_2374,N_2184);
nor U2666 (N_2666,N_2455,N_2250);
nor U2667 (N_2667,N_1935,N_2277);
xnor U2668 (N_2668,N_2210,N_2135);
xnor U2669 (N_2669,N_2383,N_2461);
or U2670 (N_2670,N_1879,N_2426);
nand U2671 (N_2671,N_2389,N_2313);
or U2672 (N_2672,N_2073,N_2029);
nor U2673 (N_2673,N_2356,N_2070);
nor U2674 (N_2674,N_2264,N_2303);
nand U2675 (N_2675,N_2495,N_2051);
or U2676 (N_2676,N_2022,N_2366);
and U2677 (N_2677,N_1946,N_2419);
nor U2678 (N_2678,N_2308,N_2171);
nor U2679 (N_2679,N_2059,N_2412);
or U2680 (N_2680,N_2057,N_2120);
nor U2681 (N_2681,N_1942,N_2276);
nand U2682 (N_2682,N_2373,N_1981);
nand U2683 (N_2683,N_2129,N_2033);
and U2684 (N_2684,N_1940,N_2367);
or U2685 (N_2685,N_2124,N_2248);
nand U2686 (N_2686,N_2138,N_2409);
nor U2687 (N_2687,N_1898,N_2251);
nand U2688 (N_2688,N_2400,N_2330);
nand U2689 (N_2689,N_2084,N_2153);
nand U2690 (N_2690,N_2061,N_2266);
nor U2691 (N_2691,N_2464,N_2309);
or U2692 (N_2692,N_2443,N_2121);
nand U2693 (N_2693,N_2381,N_2195);
nor U2694 (N_2694,N_2447,N_2499);
nor U2695 (N_2695,N_2434,N_2058);
nand U2696 (N_2696,N_2429,N_2151);
xor U2697 (N_2697,N_2445,N_1904);
nand U2698 (N_2698,N_2025,N_2149);
xor U2699 (N_2699,N_2204,N_2166);
nor U2700 (N_2700,N_1960,N_2010);
nand U2701 (N_2701,N_2425,N_1954);
and U2702 (N_2702,N_2050,N_2093);
or U2703 (N_2703,N_2032,N_1888);
nor U2704 (N_2704,N_2370,N_2096);
nand U2705 (N_2705,N_2328,N_2483);
or U2706 (N_2706,N_2353,N_2278);
xor U2707 (N_2707,N_2238,N_2305);
or U2708 (N_2708,N_1927,N_2155);
nand U2709 (N_2709,N_2450,N_2060);
and U2710 (N_2710,N_2232,N_2291);
and U2711 (N_2711,N_2013,N_1979);
and U2712 (N_2712,N_2017,N_2473);
and U2713 (N_2713,N_2441,N_1913);
or U2714 (N_2714,N_2399,N_2163);
nor U2715 (N_2715,N_1951,N_2357);
or U2716 (N_2716,N_2270,N_1955);
nor U2717 (N_2717,N_1924,N_1903);
or U2718 (N_2718,N_2418,N_1936);
nor U2719 (N_2719,N_2018,N_2463);
nor U2720 (N_2720,N_2469,N_1964);
or U2721 (N_2721,N_1948,N_1978);
or U2722 (N_2722,N_2217,N_2401);
nand U2723 (N_2723,N_2052,N_2143);
nand U2724 (N_2724,N_2333,N_2062);
and U2725 (N_2725,N_2216,N_2261);
xor U2726 (N_2726,N_1956,N_1895);
nor U2727 (N_2727,N_2363,N_2095);
nand U2728 (N_2728,N_2222,N_1878);
and U2729 (N_2729,N_2127,N_2206);
nor U2730 (N_2730,N_2225,N_2405);
nor U2731 (N_2731,N_2159,N_2081);
or U2732 (N_2732,N_2189,N_1969);
or U2733 (N_2733,N_1889,N_2260);
and U2734 (N_2734,N_1952,N_2175);
nor U2735 (N_2735,N_2079,N_2435);
and U2736 (N_2736,N_2074,N_2208);
and U2737 (N_2737,N_2299,N_2394);
nor U2738 (N_2738,N_1922,N_2341);
nor U2739 (N_2739,N_1916,N_2364);
nor U2740 (N_2740,N_1931,N_2141);
and U2741 (N_2741,N_2004,N_2384);
xor U2742 (N_2742,N_2152,N_1899);
xor U2743 (N_2743,N_2139,N_2097);
nor U2744 (N_2744,N_2411,N_2272);
or U2745 (N_2745,N_2432,N_2335);
nand U2746 (N_2746,N_2200,N_2470);
xnor U2747 (N_2747,N_1973,N_1944);
xnor U2748 (N_2748,N_2462,N_2293);
nand U2749 (N_2749,N_2201,N_1943);
nand U2750 (N_2750,N_2482,N_2267);
or U2751 (N_2751,N_2453,N_2092);
or U2752 (N_2752,N_2144,N_2243);
or U2753 (N_2753,N_2485,N_2273);
or U2754 (N_2754,N_2083,N_2015);
or U2755 (N_2755,N_2498,N_2104);
and U2756 (N_2756,N_2254,N_2302);
or U2757 (N_2757,N_2247,N_2005);
and U2758 (N_2758,N_2105,N_2324);
nand U2759 (N_2759,N_2292,N_2424);
and U2760 (N_2760,N_2421,N_2177);
or U2761 (N_2761,N_2360,N_2420);
or U2762 (N_2762,N_2192,N_2003);
nor U2763 (N_2763,N_2253,N_2492);
or U2764 (N_2764,N_2479,N_2316);
nor U2765 (N_2765,N_2317,N_2109);
or U2766 (N_2766,N_2306,N_2286);
nand U2767 (N_2767,N_2255,N_2403);
nand U2768 (N_2768,N_2282,N_2380);
and U2769 (N_2769,N_2131,N_2119);
or U2770 (N_2770,N_2361,N_2312);
and U2771 (N_2771,N_2422,N_2301);
and U2772 (N_2772,N_1945,N_1925);
nand U2773 (N_2773,N_1961,N_2475);
nand U2774 (N_2774,N_2169,N_2067);
or U2775 (N_2775,N_2414,N_2349);
and U2776 (N_2776,N_2496,N_2329);
or U2777 (N_2777,N_2205,N_2102);
or U2778 (N_2778,N_2315,N_2279);
nor U2779 (N_2779,N_2046,N_2288);
or U2780 (N_2780,N_2484,N_1921);
nand U2781 (N_2781,N_2396,N_2078);
or U2782 (N_2782,N_2041,N_1891);
or U2783 (N_2783,N_2454,N_2320);
nor U2784 (N_2784,N_1972,N_2385);
nor U2785 (N_2785,N_2221,N_2063);
and U2786 (N_2786,N_2136,N_2202);
and U2787 (N_2787,N_2433,N_2108);
nand U2788 (N_2788,N_2228,N_2340);
nor U2789 (N_2789,N_1883,N_2395);
xnor U2790 (N_2790,N_1884,N_2442);
xor U2791 (N_2791,N_1991,N_2471);
or U2792 (N_2792,N_2494,N_2458);
or U2793 (N_2793,N_2358,N_1968);
and U2794 (N_2794,N_2439,N_1932);
nand U2795 (N_2795,N_1897,N_2298);
or U2796 (N_2796,N_2082,N_1885);
or U2797 (N_2797,N_2459,N_2133);
xor U2798 (N_2798,N_2185,N_2476);
or U2799 (N_2799,N_2213,N_2220);
or U2800 (N_2800,N_2465,N_2287);
nor U2801 (N_2801,N_2021,N_2307);
nand U2802 (N_2802,N_2099,N_2390);
and U2803 (N_2803,N_1983,N_1988);
and U2804 (N_2804,N_1928,N_2178);
nor U2805 (N_2805,N_2085,N_2297);
nor U2806 (N_2806,N_2188,N_2011);
nor U2807 (N_2807,N_2362,N_2123);
and U2808 (N_2808,N_2212,N_2417);
nor U2809 (N_2809,N_2392,N_2007);
nand U2810 (N_2810,N_2049,N_2406);
or U2811 (N_2811,N_1923,N_1998);
or U2812 (N_2812,N_2468,N_1941);
nor U2813 (N_2813,N_2123,N_2032);
or U2814 (N_2814,N_2108,N_2449);
and U2815 (N_2815,N_2076,N_2072);
or U2816 (N_2816,N_2491,N_1907);
or U2817 (N_2817,N_2005,N_2182);
nor U2818 (N_2818,N_2313,N_2278);
and U2819 (N_2819,N_2178,N_2289);
nor U2820 (N_2820,N_2218,N_2119);
nor U2821 (N_2821,N_2223,N_2202);
nand U2822 (N_2822,N_1915,N_2396);
or U2823 (N_2823,N_2312,N_2281);
or U2824 (N_2824,N_2334,N_2028);
nand U2825 (N_2825,N_2124,N_2064);
and U2826 (N_2826,N_2104,N_2066);
nor U2827 (N_2827,N_2240,N_2486);
nor U2828 (N_2828,N_2255,N_2307);
or U2829 (N_2829,N_2394,N_2122);
nor U2830 (N_2830,N_2295,N_2267);
nand U2831 (N_2831,N_2361,N_2015);
nor U2832 (N_2832,N_2422,N_2054);
xnor U2833 (N_2833,N_2090,N_2111);
nor U2834 (N_2834,N_2311,N_2150);
nor U2835 (N_2835,N_2197,N_2438);
xor U2836 (N_2836,N_1951,N_2463);
or U2837 (N_2837,N_2401,N_2019);
and U2838 (N_2838,N_2171,N_1929);
or U2839 (N_2839,N_2039,N_1946);
nor U2840 (N_2840,N_2092,N_2302);
nor U2841 (N_2841,N_2288,N_2152);
or U2842 (N_2842,N_2103,N_1885);
nand U2843 (N_2843,N_2376,N_2487);
xor U2844 (N_2844,N_1923,N_1884);
or U2845 (N_2845,N_1967,N_2040);
nand U2846 (N_2846,N_2182,N_2494);
nor U2847 (N_2847,N_2191,N_2193);
and U2848 (N_2848,N_2139,N_2069);
and U2849 (N_2849,N_1940,N_2421);
xnor U2850 (N_2850,N_1987,N_2301);
nand U2851 (N_2851,N_2432,N_2298);
or U2852 (N_2852,N_1885,N_2036);
nor U2853 (N_2853,N_2073,N_2248);
nand U2854 (N_2854,N_1912,N_2289);
or U2855 (N_2855,N_2421,N_2474);
or U2856 (N_2856,N_2064,N_1901);
nand U2857 (N_2857,N_2316,N_2014);
nand U2858 (N_2858,N_1906,N_2339);
xnor U2859 (N_2859,N_2044,N_2307);
nand U2860 (N_2860,N_2422,N_2292);
nor U2861 (N_2861,N_2189,N_1940);
or U2862 (N_2862,N_2027,N_2011);
nand U2863 (N_2863,N_2313,N_2307);
and U2864 (N_2864,N_1902,N_2020);
nand U2865 (N_2865,N_2484,N_2256);
or U2866 (N_2866,N_1899,N_2046);
and U2867 (N_2867,N_2269,N_2403);
xnor U2868 (N_2868,N_2234,N_2194);
and U2869 (N_2869,N_2437,N_2016);
nor U2870 (N_2870,N_2430,N_2177);
xnor U2871 (N_2871,N_2470,N_2373);
nand U2872 (N_2872,N_2063,N_2177);
nor U2873 (N_2873,N_2497,N_1902);
nor U2874 (N_2874,N_2315,N_2218);
xor U2875 (N_2875,N_2183,N_2075);
or U2876 (N_2876,N_1988,N_2138);
and U2877 (N_2877,N_1889,N_2291);
and U2878 (N_2878,N_2483,N_2301);
xnor U2879 (N_2879,N_1940,N_2403);
nand U2880 (N_2880,N_2289,N_2198);
xnor U2881 (N_2881,N_2051,N_1942);
or U2882 (N_2882,N_2000,N_2328);
nor U2883 (N_2883,N_1897,N_1960);
nor U2884 (N_2884,N_2383,N_2082);
nor U2885 (N_2885,N_2079,N_2385);
nand U2886 (N_2886,N_2478,N_2115);
and U2887 (N_2887,N_2105,N_1936);
and U2888 (N_2888,N_1984,N_2265);
xor U2889 (N_2889,N_2289,N_2243);
or U2890 (N_2890,N_2482,N_2263);
nor U2891 (N_2891,N_2194,N_2497);
nand U2892 (N_2892,N_2434,N_2170);
nand U2893 (N_2893,N_2417,N_2427);
nand U2894 (N_2894,N_2293,N_1912);
and U2895 (N_2895,N_2290,N_2165);
and U2896 (N_2896,N_2313,N_2046);
xor U2897 (N_2897,N_2238,N_2278);
and U2898 (N_2898,N_2101,N_2496);
xor U2899 (N_2899,N_2448,N_2380);
nand U2900 (N_2900,N_2087,N_2213);
nor U2901 (N_2901,N_2478,N_2266);
nand U2902 (N_2902,N_2401,N_1916);
xor U2903 (N_2903,N_2063,N_2051);
or U2904 (N_2904,N_2496,N_2362);
nor U2905 (N_2905,N_1897,N_1999);
nor U2906 (N_2906,N_1961,N_2199);
nor U2907 (N_2907,N_2459,N_2099);
nor U2908 (N_2908,N_2086,N_1913);
xnor U2909 (N_2909,N_2482,N_2138);
and U2910 (N_2910,N_2253,N_2474);
nor U2911 (N_2911,N_2408,N_2467);
nor U2912 (N_2912,N_2442,N_2361);
nor U2913 (N_2913,N_2166,N_1985);
nor U2914 (N_2914,N_2025,N_2488);
and U2915 (N_2915,N_2140,N_2317);
nand U2916 (N_2916,N_2377,N_2482);
nor U2917 (N_2917,N_1999,N_2157);
nor U2918 (N_2918,N_1974,N_2068);
nand U2919 (N_2919,N_1932,N_2233);
or U2920 (N_2920,N_2305,N_2495);
nor U2921 (N_2921,N_2371,N_2125);
nand U2922 (N_2922,N_2102,N_1944);
nor U2923 (N_2923,N_2122,N_1984);
or U2924 (N_2924,N_2124,N_1902);
nand U2925 (N_2925,N_2121,N_2007);
nor U2926 (N_2926,N_1945,N_2275);
nand U2927 (N_2927,N_2153,N_1880);
nand U2928 (N_2928,N_2257,N_2354);
or U2929 (N_2929,N_2391,N_2332);
and U2930 (N_2930,N_2142,N_2169);
nor U2931 (N_2931,N_2142,N_2070);
xnor U2932 (N_2932,N_2282,N_2271);
nand U2933 (N_2933,N_1950,N_2029);
nand U2934 (N_2934,N_1903,N_2203);
nand U2935 (N_2935,N_1882,N_2154);
and U2936 (N_2936,N_1917,N_2497);
and U2937 (N_2937,N_2047,N_2101);
nor U2938 (N_2938,N_1954,N_2252);
xor U2939 (N_2939,N_1946,N_1875);
nor U2940 (N_2940,N_1899,N_1969);
and U2941 (N_2941,N_2408,N_2481);
xor U2942 (N_2942,N_2115,N_2365);
and U2943 (N_2943,N_2295,N_1982);
and U2944 (N_2944,N_2321,N_2452);
and U2945 (N_2945,N_2249,N_2160);
nand U2946 (N_2946,N_2218,N_2489);
or U2947 (N_2947,N_2158,N_2155);
xnor U2948 (N_2948,N_2202,N_2469);
or U2949 (N_2949,N_1907,N_1883);
or U2950 (N_2950,N_2090,N_2344);
nand U2951 (N_2951,N_2289,N_2109);
nor U2952 (N_2952,N_1909,N_2429);
nand U2953 (N_2953,N_2068,N_2484);
xor U2954 (N_2954,N_2066,N_1941);
and U2955 (N_2955,N_2378,N_2468);
or U2956 (N_2956,N_2205,N_2203);
nor U2957 (N_2957,N_2235,N_2139);
or U2958 (N_2958,N_2006,N_2340);
nor U2959 (N_2959,N_2033,N_2352);
or U2960 (N_2960,N_1890,N_2006);
or U2961 (N_2961,N_2035,N_2428);
nor U2962 (N_2962,N_2265,N_2489);
nand U2963 (N_2963,N_2336,N_2398);
or U2964 (N_2964,N_1909,N_1917);
and U2965 (N_2965,N_2381,N_2318);
or U2966 (N_2966,N_1909,N_2059);
or U2967 (N_2967,N_1976,N_2143);
and U2968 (N_2968,N_2440,N_2345);
nand U2969 (N_2969,N_2440,N_1885);
nand U2970 (N_2970,N_1926,N_2010);
or U2971 (N_2971,N_1880,N_2056);
nand U2972 (N_2972,N_2110,N_1906);
nor U2973 (N_2973,N_1879,N_2308);
and U2974 (N_2974,N_2343,N_2241);
or U2975 (N_2975,N_2105,N_2221);
nor U2976 (N_2976,N_2058,N_1965);
nand U2977 (N_2977,N_2151,N_2103);
nand U2978 (N_2978,N_1965,N_2363);
nor U2979 (N_2979,N_2066,N_2241);
nor U2980 (N_2980,N_2348,N_2385);
nor U2981 (N_2981,N_1907,N_2441);
nor U2982 (N_2982,N_2015,N_2110);
xnor U2983 (N_2983,N_2183,N_2355);
and U2984 (N_2984,N_2301,N_2458);
nand U2985 (N_2985,N_2407,N_2154);
nand U2986 (N_2986,N_2262,N_1985);
or U2987 (N_2987,N_1918,N_2079);
and U2988 (N_2988,N_1987,N_2339);
nor U2989 (N_2989,N_2099,N_1968);
and U2990 (N_2990,N_1983,N_2150);
xor U2991 (N_2991,N_2117,N_2244);
xnor U2992 (N_2992,N_2302,N_2113);
and U2993 (N_2993,N_2313,N_2321);
and U2994 (N_2994,N_2107,N_1987);
nor U2995 (N_2995,N_2486,N_2467);
or U2996 (N_2996,N_2148,N_2280);
and U2997 (N_2997,N_2335,N_2173);
or U2998 (N_2998,N_2387,N_2410);
and U2999 (N_2999,N_2325,N_2059);
or U3000 (N_3000,N_2142,N_2315);
nand U3001 (N_3001,N_2091,N_2397);
or U3002 (N_3002,N_1930,N_2038);
and U3003 (N_3003,N_1904,N_1905);
nor U3004 (N_3004,N_2023,N_2136);
nor U3005 (N_3005,N_2470,N_2327);
nor U3006 (N_3006,N_2332,N_2175);
nor U3007 (N_3007,N_2385,N_2452);
nand U3008 (N_3008,N_2453,N_2413);
or U3009 (N_3009,N_1904,N_2099);
nand U3010 (N_3010,N_1960,N_2468);
nand U3011 (N_3011,N_1972,N_1915);
and U3012 (N_3012,N_2314,N_2429);
nand U3013 (N_3013,N_2496,N_2098);
or U3014 (N_3014,N_2385,N_2296);
or U3015 (N_3015,N_2098,N_2287);
and U3016 (N_3016,N_2053,N_2482);
or U3017 (N_3017,N_1893,N_2113);
nor U3018 (N_3018,N_1976,N_2214);
nand U3019 (N_3019,N_1879,N_2156);
xnor U3020 (N_3020,N_2441,N_2094);
nor U3021 (N_3021,N_2350,N_2087);
nor U3022 (N_3022,N_2488,N_2189);
and U3023 (N_3023,N_2227,N_2424);
nand U3024 (N_3024,N_2101,N_2248);
nand U3025 (N_3025,N_2365,N_2419);
nand U3026 (N_3026,N_1996,N_2150);
and U3027 (N_3027,N_2461,N_2444);
and U3028 (N_3028,N_2311,N_1957);
and U3029 (N_3029,N_2006,N_2208);
nor U3030 (N_3030,N_2297,N_2207);
nor U3031 (N_3031,N_1928,N_2120);
nand U3032 (N_3032,N_2004,N_2059);
and U3033 (N_3033,N_2201,N_2165);
nand U3034 (N_3034,N_1932,N_2033);
or U3035 (N_3035,N_2311,N_2354);
or U3036 (N_3036,N_2101,N_2201);
and U3037 (N_3037,N_2342,N_1961);
and U3038 (N_3038,N_2200,N_2060);
and U3039 (N_3039,N_2400,N_1994);
and U3040 (N_3040,N_2358,N_2323);
nand U3041 (N_3041,N_2336,N_2391);
nor U3042 (N_3042,N_2237,N_2061);
and U3043 (N_3043,N_2439,N_2356);
or U3044 (N_3044,N_1952,N_2353);
nand U3045 (N_3045,N_2259,N_2157);
and U3046 (N_3046,N_2428,N_2054);
nand U3047 (N_3047,N_2403,N_1925);
nand U3048 (N_3048,N_2272,N_1974);
nand U3049 (N_3049,N_1907,N_2194);
or U3050 (N_3050,N_2346,N_2323);
and U3051 (N_3051,N_2208,N_2188);
or U3052 (N_3052,N_2130,N_2282);
or U3053 (N_3053,N_2297,N_2145);
nor U3054 (N_3054,N_2159,N_2012);
nor U3055 (N_3055,N_2211,N_2040);
xor U3056 (N_3056,N_2245,N_1927);
nor U3057 (N_3057,N_2214,N_2384);
nand U3058 (N_3058,N_1916,N_2393);
or U3059 (N_3059,N_1887,N_2262);
or U3060 (N_3060,N_2317,N_2024);
and U3061 (N_3061,N_2491,N_2275);
nor U3062 (N_3062,N_1940,N_2006);
and U3063 (N_3063,N_1941,N_1900);
nor U3064 (N_3064,N_2409,N_2126);
nand U3065 (N_3065,N_2380,N_2022);
or U3066 (N_3066,N_2493,N_2107);
and U3067 (N_3067,N_1901,N_2008);
or U3068 (N_3068,N_2432,N_2019);
or U3069 (N_3069,N_2375,N_2310);
nor U3070 (N_3070,N_2478,N_2254);
xnor U3071 (N_3071,N_2198,N_2086);
nor U3072 (N_3072,N_2498,N_2492);
or U3073 (N_3073,N_2126,N_2277);
nor U3074 (N_3074,N_2069,N_2047);
xor U3075 (N_3075,N_2235,N_2293);
and U3076 (N_3076,N_2201,N_2495);
xor U3077 (N_3077,N_2107,N_2390);
xor U3078 (N_3078,N_2158,N_2352);
nand U3079 (N_3079,N_2345,N_2306);
xnor U3080 (N_3080,N_2459,N_2355);
or U3081 (N_3081,N_2096,N_2332);
and U3082 (N_3082,N_2400,N_2479);
nor U3083 (N_3083,N_2420,N_2335);
or U3084 (N_3084,N_2296,N_2320);
nor U3085 (N_3085,N_2278,N_1920);
or U3086 (N_3086,N_2490,N_1894);
nor U3087 (N_3087,N_2019,N_2273);
and U3088 (N_3088,N_2117,N_2253);
or U3089 (N_3089,N_2376,N_2351);
or U3090 (N_3090,N_2094,N_2250);
or U3091 (N_3091,N_2016,N_2397);
or U3092 (N_3092,N_1898,N_2062);
nor U3093 (N_3093,N_1954,N_2110);
and U3094 (N_3094,N_2422,N_2375);
nand U3095 (N_3095,N_2036,N_2221);
nor U3096 (N_3096,N_1881,N_2396);
nand U3097 (N_3097,N_2021,N_2263);
nand U3098 (N_3098,N_2360,N_2477);
nor U3099 (N_3099,N_2353,N_2301);
xor U3100 (N_3100,N_2146,N_2396);
or U3101 (N_3101,N_2246,N_2410);
nand U3102 (N_3102,N_1908,N_2016);
nor U3103 (N_3103,N_2156,N_2452);
nor U3104 (N_3104,N_2446,N_2216);
nand U3105 (N_3105,N_1932,N_1935);
xor U3106 (N_3106,N_1893,N_2096);
or U3107 (N_3107,N_2074,N_2086);
xnor U3108 (N_3108,N_2048,N_2224);
nand U3109 (N_3109,N_2493,N_2149);
or U3110 (N_3110,N_2298,N_1957);
and U3111 (N_3111,N_2169,N_2406);
and U3112 (N_3112,N_2443,N_1944);
nand U3113 (N_3113,N_2436,N_2129);
nor U3114 (N_3114,N_1912,N_2303);
nor U3115 (N_3115,N_2484,N_2441);
and U3116 (N_3116,N_2312,N_2430);
nand U3117 (N_3117,N_2153,N_1985);
xnor U3118 (N_3118,N_2260,N_2153);
and U3119 (N_3119,N_2480,N_2331);
nand U3120 (N_3120,N_2374,N_2204);
nor U3121 (N_3121,N_1979,N_2056);
or U3122 (N_3122,N_2085,N_2445);
and U3123 (N_3123,N_2032,N_1894);
nand U3124 (N_3124,N_2485,N_2009);
nand U3125 (N_3125,N_2892,N_2821);
nor U3126 (N_3126,N_2734,N_2745);
xnor U3127 (N_3127,N_2597,N_2930);
xor U3128 (N_3128,N_2800,N_2767);
nand U3129 (N_3129,N_2656,N_3106);
nand U3130 (N_3130,N_3074,N_2657);
nand U3131 (N_3131,N_2620,N_2851);
xnor U3132 (N_3132,N_2525,N_2839);
nor U3133 (N_3133,N_2996,N_2625);
xnor U3134 (N_3134,N_2601,N_2995);
or U3135 (N_3135,N_2901,N_2738);
nand U3136 (N_3136,N_2565,N_2651);
xnor U3137 (N_3137,N_2621,N_2772);
or U3138 (N_3138,N_2542,N_2722);
nand U3139 (N_3139,N_3043,N_2872);
xor U3140 (N_3140,N_2580,N_2764);
nor U3141 (N_3141,N_2773,N_2677);
xnor U3142 (N_3142,N_2889,N_2724);
nor U3143 (N_3143,N_3105,N_2627);
nor U3144 (N_3144,N_2810,N_2850);
or U3145 (N_3145,N_2719,N_2750);
nand U3146 (N_3146,N_3119,N_3047);
nor U3147 (N_3147,N_2557,N_2575);
and U3148 (N_3148,N_3013,N_2523);
nor U3149 (N_3149,N_3021,N_2529);
nand U3150 (N_3150,N_2970,N_2546);
nand U3151 (N_3151,N_2923,N_2989);
or U3152 (N_3152,N_2687,N_2743);
and U3153 (N_3153,N_2667,N_2538);
and U3154 (N_3154,N_3020,N_2862);
xnor U3155 (N_3155,N_2781,N_2793);
nor U3156 (N_3156,N_3098,N_2711);
nor U3157 (N_3157,N_2512,N_2938);
xnor U3158 (N_3158,N_3014,N_2683);
or U3159 (N_3159,N_2501,N_2791);
nor U3160 (N_3160,N_3005,N_2804);
nor U3161 (N_3161,N_2552,N_2547);
or U3162 (N_3162,N_3115,N_2927);
or U3163 (N_3163,N_2785,N_2689);
or U3164 (N_3164,N_2912,N_2991);
or U3165 (N_3165,N_2961,N_2818);
and U3166 (N_3166,N_2720,N_2606);
nand U3167 (N_3167,N_2618,N_3110);
and U3168 (N_3168,N_3058,N_2631);
or U3169 (N_3169,N_2690,N_2803);
nor U3170 (N_3170,N_2582,N_3104);
nand U3171 (N_3171,N_2762,N_3083);
or U3172 (N_3172,N_2572,N_2929);
or U3173 (N_3173,N_3015,N_3076);
or U3174 (N_3174,N_2515,N_2902);
nand U3175 (N_3175,N_3009,N_2957);
nand U3176 (N_3176,N_2685,N_3017);
and U3177 (N_3177,N_3007,N_2884);
xnor U3178 (N_3178,N_2693,N_2858);
nor U3179 (N_3179,N_2635,N_2681);
and U3180 (N_3180,N_3045,N_2533);
nor U3181 (N_3181,N_2654,N_2945);
nand U3182 (N_3182,N_2954,N_2502);
xor U3183 (N_3183,N_3026,N_2900);
nor U3184 (N_3184,N_2798,N_3027);
nand U3185 (N_3185,N_2934,N_3031);
and U3186 (N_3186,N_2587,N_2647);
or U3187 (N_3187,N_2511,N_2973);
nand U3188 (N_3188,N_2865,N_3070);
nand U3189 (N_3189,N_2895,N_2917);
or U3190 (N_3190,N_2562,N_3002);
nand U3191 (N_3191,N_2983,N_2866);
xnor U3192 (N_3192,N_2553,N_2691);
nand U3193 (N_3193,N_2758,N_2664);
or U3194 (N_3194,N_3064,N_3008);
nand U3195 (N_3195,N_2932,N_2586);
nor U3196 (N_3196,N_2644,N_3010);
nor U3197 (N_3197,N_2613,N_3036);
xnor U3198 (N_3198,N_3032,N_3089);
nor U3199 (N_3199,N_2779,N_3082);
or U3200 (N_3200,N_3030,N_3060);
nor U3201 (N_3201,N_2857,N_2518);
nand U3202 (N_3202,N_2801,N_2759);
nor U3203 (N_3203,N_2964,N_2633);
or U3204 (N_3204,N_3117,N_2795);
or U3205 (N_3205,N_2675,N_2561);
nand U3206 (N_3206,N_2976,N_2638);
or U3207 (N_3207,N_3011,N_2579);
or U3208 (N_3208,N_2765,N_2829);
nand U3209 (N_3209,N_2662,N_2636);
nand U3210 (N_3210,N_2668,N_2897);
or U3211 (N_3211,N_3109,N_2814);
nor U3212 (N_3212,N_2949,N_2963);
and U3213 (N_3213,N_2527,N_2898);
or U3214 (N_3214,N_2864,N_2770);
nand U3215 (N_3215,N_2840,N_2893);
or U3216 (N_3216,N_3001,N_2761);
or U3217 (N_3217,N_2676,N_2922);
nor U3218 (N_3218,N_2706,N_2595);
nor U3219 (N_3219,N_2640,N_3016);
and U3220 (N_3220,N_2521,N_2506);
nor U3221 (N_3221,N_2737,N_2548);
nor U3222 (N_3222,N_2926,N_2933);
nand U3223 (N_3223,N_2918,N_2704);
and U3224 (N_3224,N_2740,N_2522);
or U3225 (N_3225,N_2555,N_2659);
nand U3226 (N_3226,N_2571,N_2948);
nand U3227 (N_3227,N_2725,N_2746);
nor U3228 (N_3228,N_3059,N_2500);
nor U3229 (N_3229,N_3056,N_3022);
nor U3230 (N_3230,N_2890,N_2747);
nor U3231 (N_3231,N_2695,N_2678);
or U3232 (N_3232,N_2710,N_2824);
xnor U3233 (N_3233,N_2653,N_2739);
and U3234 (N_3234,N_2870,N_2838);
nor U3235 (N_3235,N_2888,N_2652);
nor U3236 (N_3236,N_2972,N_2891);
nand U3237 (N_3237,N_3123,N_2760);
or U3238 (N_3238,N_3108,N_2741);
nand U3239 (N_3239,N_2728,N_2835);
or U3240 (N_3240,N_3071,N_2554);
nand U3241 (N_3241,N_2585,N_2703);
or U3242 (N_3242,N_3034,N_3039);
nand U3243 (N_3243,N_2777,N_2602);
and U3244 (N_3244,N_3116,N_3075);
nand U3245 (N_3245,N_2592,N_2830);
or U3246 (N_3246,N_3093,N_2962);
and U3247 (N_3247,N_2569,N_2783);
nand U3248 (N_3248,N_2763,N_2910);
and U3249 (N_3249,N_2573,N_2655);
or U3250 (N_3250,N_3087,N_3084);
nand U3251 (N_3251,N_2503,N_3073);
nor U3252 (N_3252,N_2697,N_2673);
and U3253 (N_3253,N_2827,N_2622);
xnor U3254 (N_3254,N_2806,N_2637);
or U3255 (N_3255,N_3038,N_2992);
and U3256 (N_3256,N_3063,N_2873);
nand U3257 (N_3257,N_2576,N_3061);
and U3258 (N_3258,N_2849,N_2952);
and U3259 (N_3259,N_2990,N_2817);
nor U3260 (N_3260,N_2813,N_2843);
nand U3261 (N_3261,N_2903,N_2812);
nor U3262 (N_3262,N_2874,N_3086);
nand U3263 (N_3263,N_2596,N_2713);
or U3264 (N_3264,N_3049,N_2846);
nor U3265 (N_3265,N_2610,N_2836);
or U3266 (N_3266,N_2563,N_2568);
nand U3267 (N_3267,N_2574,N_2679);
nor U3268 (N_3268,N_3078,N_2699);
or U3269 (N_3269,N_2646,N_2977);
and U3270 (N_3270,N_2768,N_2540);
and U3271 (N_3271,N_3054,N_2986);
nand U3272 (N_3272,N_2560,N_2550);
and U3273 (N_3273,N_2978,N_3023);
and U3274 (N_3274,N_2841,N_2670);
and U3275 (N_3275,N_2634,N_2507);
nand U3276 (N_3276,N_2784,N_2950);
nor U3277 (N_3277,N_2985,N_2535);
nor U3278 (N_3278,N_2714,N_2794);
or U3279 (N_3279,N_2680,N_3051);
and U3280 (N_3280,N_2811,N_3044);
nor U3281 (N_3281,N_2614,N_3114);
or U3282 (N_3282,N_2854,N_2701);
and U3283 (N_3283,N_2578,N_2965);
nor U3284 (N_3284,N_2643,N_3006);
nor U3285 (N_3285,N_3112,N_2796);
nand U3286 (N_3286,N_3018,N_2751);
nor U3287 (N_3287,N_2756,N_2942);
and U3288 (N_3288,N_2534,N_3003);
or U3289 (N_3289,N_2820,N_3065);
and U3290 (N_3290,N_2921,N_2649);
and U3291 (N_3291,N_2974,N_2551);
and U3292 (N_3292,N_2726,N_2604);
nor U3293 (N_3293,N_2959,N_2896);
nand U3294 (N_3294,N_3042,N_2982);
nand U3295 (N_3295,N_2639,N_3069);
nand U3296 (N_3296,N_2882,N_2732);
nand U3297 (N_3297,N_3028,N_2729);
or U3298 (N_3298,N_2789,N_3088);
nand U3299 (N_3299,N_2567,N_2530);
or U3300 (N_3300,N_2826,N_2847);
nor U3301 (N_3301,N_2536,N_2940);
xor U3302 (N_3302,N_3055,N_2886);
nand U3303 (N_3303,N_3085,N_2907);
and U3304 (N_3304,N_3029,N_2988);
nor U3305 (N_3305,N_2859,N_2861);
nor U3306 (N_3306,N_2909,N_2581);
nand U3307 (N_3307,N_2539,N_2871);
or U3308 (N_3308,N_2947,N_2845);
nand U3309 (N_3309,N_2730,N_2626);
nand U3310 (N_3310,N_3019,N_2570);
nand U3311 (N_3311,N_2612,N_3101);
nor U3312 (N_3312,N_2808,N_3124);
nor U3313 (N_3313,N_3040,N_2709);
and U3314 (N_3314,N_2509,N_2915);
nand U3315 (N_3315,N_3050,N_2943);
nor U3316 (N_3316,N_2899,N_2832);
nor U3317 (N_3317,N_3095,N_2516);
nor U3318 (N_3318,N_2831,N_2559);
and U3319 (N_3319,N_2733,N_2834);
nand U3320 (N_3320,N_2956,N_2969);
and U3321 (N_3321,N_2630,N_2744);
or U3322 (N_3322,N_3090,N_2925);
nor U3323 (N_3323,N_3068,N_3062);
and U3324 (N_3324,N_2876,N_3092);
nand U3325 (N_3325,N_2543,N_3052);
nor U3326 (N_3326,N_3057,N_2520);
and U3327 (N_3327,N_2788,N_2526);
nand U3328 (N_3328,N_2894,N_3000);
and U3329 (N_3329,N_2881,N_2920);
and U3330 (N_3330,N_3107,N_2844);
nand U3331 (N_3331,N_3079,N_2686);
nand U3332 (N_3332,N_2999,N_2615);
nor U3333 (N_3333,N_2782,N_2603);
xnor U3334 (N_3334,N_2828,N_2708);
and U3335 (N_3335,N_2774,N_2674);
nand U3336 (N_3336,N_2936,N_2805);
xor U3337 (N_3337,N_2877,N_2584);
and U3338 (N_3338,N_3103,N_2624);
and U3339 (N_3339,N_2944,N_2532);
and U3340 (N_3340,N_2855,N_2698);
or U3341 (N_3341,N_2755,N_3094);
or U3342 (N_3342,N_2757,N_2931);
or U3343 (N_3343,N_2809,N_3025);
nand U3344 (N_3344,N_2519,N_2807);
xnor U3345 (N_3345,N_2694,N_3080);
nand U3346 (N_3346,N_3053,N_3041);
xor U3347 (N_3347,N_2611,N_2863);
or U3348 (N_3348,N_2752,N_2853);
nor U3349 (N_3349,N_2955,N_2684);
nor U3350 (N_3350,N_2692,N_2537);
or U3351 (N_3351,N_2508,N_3048);
and U3352 (N_3352,N_2905,N_2669);
or U3353 (N_3353,N_2967,N_2632);
or U3354 (N_3354,N_2993,N_2875);
and U3355 (N_3355,N_2769,N_2629);
nand U3356 (N_3356,N_2517,N_2868);
or U3357 (N_3357,N_2504,N_2717);
nor U3358 (N_3358,N_3121,N_2556);
xor U3359 (N_3359,N_2776,N_2797);
and U3360 (N_3360,N_3120,N_2524);
nor U3361 (N_3361,N_2642,N_3122);
nor U3362 (N_3362,N_2528,N_2658);
nor U3363 (N_3363,N_2593,N_3081);
nor U3364 (N_3364,N_2975,N_2682);
or U3365 (N_3365,N_3077,N_2867);
nand U3366 (N_3366,N_2754,N_2702);
nand U3367 (N_3367,N_2981,N_2911);
xnor U3368 (N_3368,N_2608,N_2577);
and U3369 (N_3369,N_2531,N_2705);
nor U3370 (N_3370,N_2939,N_2825);
or U3371 (N_3371,N_2815,N_3100);
or U3372 (N_3372,N_2786,N_2913);
nand U3373 (N_3373,N_2696,N_2766);
or U3374 (N_3374,N_2998,N_2816);
and U3375 (N_3375,N_2727,N_2661);
or U3376 (N_3376,N_2609,N_2598);
nand U3377 (N_3377,N_3033,N_2914);
nand U3378 (N_3378,N_2802,N_2980);
or U3379 (N_3379,N_2749,N_2748);
or U3380 (N_3380,N_3067,N_2619);
nor U3381 (N_3381,N_2979,N_3004);
xnor U3382 (N_3382,N_3096,N_2663);
nor U3383 (N_3383,N_2617,N_3091);
nor U3384 (N_3384,N_2833,N_3118);
nand U3385 (N_3385,N_2648,N_3046);
or U3386 (N_3386,N_2822,N_2721);
or U3387 (N_3387,N_2966,N_2984);
nand U3388 (N_3388,N_2819,N_2672);
and U3389 (N_3389,N_2885,N_3111);
or U3390 (N_3390,N_2505,N_2666);
or U3391 (N_3391,N_2545,N_2968);
or U3392 (N_3392,N_2887,N_2645);
and U3393 (N_3393,N_2715,N_2600);
xnor U3394 (N_3394,N_3024,N_2823);
nand U3395 (N_3395,N_3113,N_2607);
nand U3396 (N_3396,N_2916,N_2544);
or U3397 (N_3397,N_2792,N_3035);
or U3398 (N_3398,N_2878,N_2660);
nand U3399 (N_3399,N_2771,N_2946);
xor U3400 (N_3400,N_3097,N_2971);
xor U3401 (N_3401,N_3037,N_2780);
and U3402 (N_3402,N_2549,N_2735);
nand U3403 (N_3403,N_2514,N_2790);
nor U3404 (N_3404,N_2775,N_2953);
nand U3405 (N_3405,N_2558,N_2712);
and U3406 (N_3406,N_2958,N_2987);
xnor U3407 (N_3407,N_2513,N_2951);
nor U3408 (N_3408,N_2641,N_2700);
and U3409 (N_3409,N_2628,N_2842);
or U3410 (N_3410,N_3072,N_2924);
or U3411 (N_3411,N_2848,N_2860);
nand U3412 (N_3412,N_2837,N_2906);
nand U3413 (N_3413,N_2605,N_2583);
and U3414 (N_3414,N_2994,N_2869);
nor U3415 (N_3415,N_3012,N_2566);
and U3416 (N_3416,N_3099,N_2919);
nor U3417 (N_3417,N_2731,N_2778);
nand U3418 (N_3418,N_2852,N_2564);
or U3419 (N_3419,N_2879,N_2941);
and U3420 (N_3420,N_2937,N_2650);
nand U3421 (N_3421,N_2594,N_2591);
nor U3422 (N_3422,N_2856,N_2599);
xor U3423 (N_3423,N_2960,N_2883);
or U3424 (N_3424,N_2665,N_2616);
and U3425 (N_3425,N_2541,N_2787);
nand U3426 (N_3426,N_2716,N_2510);
and U3427 (N_3427,N_2588,N_2589);
or U3428 (N_3428,N_3102,N_2997);
or U3429 (N_3429,N_2688,N_2935);
nand U3430 (N_3430,N_2736,N_2904);
or U3431 (N_3431,N_2671,N_2799);
nand U3432 (N_3432,N_3066,N_2880);
nand U3433 (N_3433,N_2590,N_2928);
nand U3434 (N_3434,N_2742,N_2908);
nor U3435 (N_3435,N_2753,N_2707);
nor U3436 (N_3436,N_2623,N_2723);
and U3437 (N_3437,N_2718,N_2788);
nand U3438 (N_3438,N_3046,N_2707);
and U3439 (N_3439,N_2609,N_2770);
nand U3440 (N_3440,N_2694,N_3110);
nand U3441 (N_3441,N_2837,N_2975);
nand U3442 (N_3442,N_2638,N_3047);
xnor U3443 (N_3443,N_3108,N_3077);
nand U3444 (N_3444,N_2505,N_2786);
nand U3445 (N_3445,N_2505,N_2682);
nor U3446 (N_3446,N_3054,N_2945);
or U3447 (N_3447,N_2579,N_2549);
and U3448 (N_3448,N_2816,N_3032);
nor U3449 (N_3449,N_2626,N_2864);
nand U3450 (N_3450,N_2748,N_2695);
and U3451 (N_3451,N_2890,N_3076);
or U3452 (N_3452,N_2568,N_2680);
nor U3453 (N_3453,N_2574,N_2974);
or U3454 (N_3454,N_2603,N_2794);
nand U3455 (N_3455,N_2643,N_2854);
and U3456 (N_3456,N_2907,N_2792);
nand U3457 (N_3457,N_2941,N_2571);
and U3458 (N_3458,N_2566,N_2930);
nor U3459 (N_3459,N_2577,N_2972);
and U3460 (N_3460,N_2724,N_2923);
nand U3461 (N_3461,N_2558,N_2563);
and U3462 (N_3462,N_3013,N_3094);
nor U3463 (N_3463,N_2638,N_2614);
or U3464 (N_3464,N_2729,N_2631);
nand U3465 (N_3465,N_2696,N_2856);
nand U3466 (N_3466,N_2707,N_2738);
xor U3467 (N_3467,N_2590,N_2864);
and U3468 (N_3468,N_3093,N_2528);
xor U3469 (N_3469,N_3068,N_2941);
nor U3470 (N_3470,N_3097,N_2985);
nand U3471 (N_3471,N_2972,N_2942);
and U3472 (N_3472,N_2628,N_2512);
or U3473 (N_3473,N_3119,N_2800);
or U3474 (N_3474,N_2836,N_2599);
nor U3475 (N_3475,N_2754,N_2843);
or U3476 (N_3476,N_2850,N_3025);
or U3477 (N_3477,N_2945,N_3057);
nand U3478 (N_3478,N_2715,N_2652);
or U3479 (N_3479,N_2502,N_3036);
or U3480 (N_3480,N_2894,N_2837);
nor U3481 (N_3481,N_2847,N_2623);
nor U3482 (N_3482,N_2740,N_2911);
nand U3483 (N_3483,N_2911,N_2512);
or U3484 (N_3484,N_2645,N_2823);
and U3485 (N_3485,N_2643,N_3106);
nor U3486 (N_3486,N_2687,N_2803);
nand U3487 (N_3487,N_2630,N_2515);
and U3488 (N_3488,N_2564,N_3111);
nor U3489 (N_3489,N_3090,N_2980);
and U3490 (N_3490,N_2697,N_2724);
and U3491 (N_3491,N_2791,N_2729);
and U3492 (N_3492,N_3035,N_3002);
and U3493 (N_3493,N_2870,N_2728);
or U3494 (N_3494,N_2669,N_2562);
nor U3495 (N_3495,N_2694,N_2906);
nand U3496 (N_3496,N_3064,N_2574);
or U3497 (N_3497,N_3070,N_3033);
or U3498 (N_3498,N_2823,N_2744);
nor U3499 (N_3499,N_2665,N_2611);
and U3500 (N_3500,N_2852,N_2630);
nand U3501 (N_3501,N_2785,N_3000);
or U3502 (N_3502,N_3076,N_2983);
and U3503 (N_3503,N_2744,N_2589);
or U3504 (N_3504,N_2538,N_2966);
xnor U3505 (N_3505,N_2786,N_3037);
or U3506 (N_3506,N_3036,N_2676);
and U3507 (N_3507,N_2960,N_2916);
and U3508 (N_3508,N_3003,N_3008);
or U3509 (N_3509,N_2964,N_2938);
xnor U3510 (N_3510,N_2968,N_2615);
nand U3511 (N_3511,N_2555,N_2986);
and U3512 (N_3512,N_2900,N_2834);
and U3513 (N_3513,N_2714,N_2551);
nand U3514 (N_3514,N_2974,N_2979);
nand U3515 (N_3515,N_2810,N_2837);
xor U3516 (N_3516,N_2532,N_2791);
nand U3517 (N_3517,N_2671,N_3100);
nor U3518 (N_3518,N_2900,N_2940);
and U3519 (N_3519,N_2683,N_2726);
xnor U3520 (N_3520,N_2907,N_2624);
and U3521 (N_3521,N_2503,N_2971);
nand U3522 (N_3522,N_2765,N_2669);
and U3523 (N_3523,N_2545,N_3107);
nor U3524 (N_3524,N_2744,N_2590);
xnor U3525 (N_3525,N_2755,N_2905);
nor U3526 (N_3526,N_2612,N_3022);
or U3527 (N_3527,N_2881,N_3055);
and U3528 (N_3528,N_2687,N_2720);
and U3529 (N_3529,N_3091,N_2967);
or U3530 (N_3530,N_3109,N_3056);
nor U3531 (N_3531,N_2748,N_2977);
nand U3532 (N_3532,N_2946,N_2547);
or U3533 (N_3533,N_3019,N_2684);
and U3534 (N_3534,N_3060,N_3054);
nor U3535 (N_3535,N_2999,N_3098);
nand U3536 (N_3536,N_2614,N_2815);
nor U3537 (N_3537,N_3114,N_2638);
xor U3538 (N_3538,N_2583,N_3037);
xor U3539 (N_3539,N_2860,N_3046);
or U3540 (N_3540,N_2904,N_2938);
nand U3541 (N_3541,N_2610,N_2852);
xnor U3542 (N_3542,N_2597,N_3013);
or U3543 (N_3543,N_2743,N_2910);
nand U3544 (N_3544,N_2846,N_2967);
or U3545 (N_3545,N_2931,N_2727);
and U3546 (N_3546,N_2999,N_2812);
or U3547 (N_3547,N_2962,N_2571);
and U3548 (N_3548,N_3096,N_2899);
or U3549 (N_3549,N_2980,N_3047);
or U3550 (N_3550,N_2662,N_2766);
nand U3551 (N_3551,N_2666,N_2664);
and U3552 (N_3552,N_2845,N_2708);
nand U3553 (N_3553,N_2586,N_3054);
or U3554 (N_3554,N_2992,N_3041);
and U3555 (N_3555,N_2776,N_2871);
or U3556 (N_3556,N_2786,N_2790);
or U3557 (N_3557,N_2670,N_2890);
nor U3558 (N_3558,N_2989,N_2837);
or U3559 (N_3559,N_2653,N_2808);
xnor U3560 (N_3560,N_2654,N_2594);
and U3561 (N_3561,N_3120,N_2704);
xnor U3562 (N_3562,N_2927,N_2584);
and U3563 (N_3563,N_2624,N_2506);
nand U3564 (N_3564,N_2905,N_3103);
nand U3565 (N_3565,N_2548,N_2614);
and U3566 (N_3566,N_2638,N_2721);
nand U3567 (N_3567,N_2805,N_2592);
xnor U3568 (N_3568,N_2764,N_2637);
nand U3569 (N_3569,N_2584,N_2907);
and U3570 (N_3570,N_2818,N_2809);
xnor U3571 (N_3571,N_2806,N_2748);
nand U3572 (N_3572,N_2768,N_2917);
nor U3573 (N_3573,N_2748,N_3001);
or U3574 (N_3574,N_3020,N_2662);
and U3575 (N_3575,N_3026,N_2803);
nand U3576 (N_3576,N_2875,N_2792);
or U3577 (N_3577,N_2777,N_3096);
or U3578 (N_3578,N_2576,N_3071);
nor U3579 (N_3579,N_3005,N_2891);
xor U3580 (N_3580,N_3078,N_2778);
or U3581 (N_3581,N_2853,N_3099);
nand U3582 (N_3582,N_2964,N_2612);
and U3583 (N_3583,N_3085,N_2810);
or U3584 (N_3584,N_3085,N_3047);
nand U3585 (N_3585,N_3089,N_2844);
or U3586 (N_3586,N_2639,N_2520);
nand U3587 (N_3587,N_2980,N_2855);
nand U3588 (N_3588,N_2509,N_2806);
or U3589 (N_3589,N_3119,N_2765);
nand U3590 (N_3590,N_2705,N_2706);
nor U3591 (N_3591,N_3017,N_2654);
xnor U3592 (N_3592,N_2895,N_3043);
nor U3593 (N_3593,N_2713,N_2549);
or U3594 (N_3594,N_2847,N_3014);
or U3595 (N_3595,N_2731,N_2947);
nand U3596 (N_3596,N_3048,N_2883);
nand U3597 (N_3597,N_2647,N_2812);
nand U3598 (N_3598,N_2541,N_2781);
or U3599 (N_3599,N_2746,N_2535);
nor U3600 (N_3600,N_3028,N_3062);
nor U3601 (N_3601,N_2634,N_2983);
nor U3602 (N_3602,N_2765,N_2748);
and U3603 (N_3603,N_2981,N_2650);
nand U3604 (N_3604,N_2503,N_2811);
nand U3605 (N_3605,N_2643,N_2763);
and U3606 (N_3606,N_2608,N_2806);
nor U3607 (N_3607,N_2568,N_2808);
nand U3608 (N_3608,N_2637,N_2886);
or U3609 (N_3609,N_2675,N_2993);
or U3610 (N_3610,N_2941,N_2593);
or U3611 (N_3611,N_2737,N_2736);
nand U3612 (N_3612,N_2992,N_3073);
xnor U3613 (N_3613,N_2927,N_2944);
and U3614 (N_3614,N_3047,N_2792);
or U3615 (N_3615,N_2942,N_2552);
nand U3616 (N_3616,N_3092,N_2795);
nand U3617 (N_3617,N_2888,N_3041);
nand U3618 (N_3618,N_2783,N_2922);
nand U3619 (N_3619,N_3025,N_3116);
and U3620 (N_3620,N_2784,N_2979);
nand U3621 (N_3621,N_2701,N_3062);
or U3622 (N_3622,N_2758,N_2757);
and U3623 (N_3623,N_2917,N_2857);
or U3624 (N_3624,N_3090,N_2649);
nor U3625 (N_3625,N_3023,N_2822);
or U3626 (N_3626,N_2575,N_2754);
nor U3627 (N_3627,N_2937,N_2954);
and U3628 (N_3628,N_2718,N_2572);
nand U3629 (N_3629,N_2876,N_2733);
and U3630 (N_3630,N_2976,N_2859);
or U3631 (N_3631,N_2777,N_2972);
nand U3632 (N_3632,N_2881,N_2645);
nor U3633 (N_3633,N_3025,N_2720);
nand U3634 (N_3634,N_3014,N_2517);
or U3635 (N_3635,N_2920,N_2873);
or U3636 (N_3636,N_3105,N_2984);
nor U3637 (N_3637,N_2993,N_2688);
and U3638 (N_3638,N_2553,N_3026);
or U3639 (N_3639,N_2914,N_2553);
xor U3640 (N_3640,N_2597,N_2849);
nand U3641 (N_3641,N_3028,N_2836);
nand U3642 (N_3642,N_2735,N_2813);
nand U3643 (N_3643,N_3037,N_3034);
nand U3644 (N_3644,N_3015,N_3094);
and U3645 (N_3645,N_2626,N_2647);
xor U3646 (N_3646,N_2704,N_3002);
and U3647 (N_3647,N_2547,N_3099);
nor U3648 (N_3648,N_2613,N_2725);
nand U3649 (N_3649,N_2828,N_2648);
nand U3650 (N_3650,N_2599,N_2990);
nor U3651 (N_3651,N_3093,N_2779);
nor U3652 (N_3652,N_2864,N_2936);
and U3653 (N_3653,N_2659,N_2996);
and U3654 (N_3654,N_2630,N_2571);
or U3655 (N_3655,N_2717,N_2593);
nand U3656 (N_3656,N_2821,N_2918);
nor U3657 (N_3657,N_2734,N_2900);
or U3658 (N_3658,N_2872,N_2590);
nor U3659 (N_3659,N_2821,N_2973);
or U3660 (N_3660,N_2697,N_2733);
xor U3661 (N_3661,N_2574,N_2938);
and U3662 (N_3662,N_2736,N_3047);
nor U3663 (N_3663,N_2638,N_2818);
or U3664 (N_3664,N_3055,N_3034);
xor U3665 (N_3665,N_2760,N_2956);
or U3666 (N_3666,N_2504,N_2774);
or U3667 (N_3667,N_2907,N_3032);
nor U3668 (N_3668,N_2512,N_2815);
nor U3669 (N_3669,N_2803,N_3035);
and U3670 (N_3670,N_3094,N_2718);
nor U3671 (N_3671,N_2650,N_2951);
or U3672 (N_3672,N_2576,N_2958);
and U3673 (N_3673,N_2903,N_2983);
or U3674 (N_3674,N_2629,N_2787);
and U3675 (N_3675,N_2616,N_2628);
or U3676 (N_3676,N_2601,N_2837);
nor U3677 (N_3677,N_2706,N_2767);
nor U3678 (N_3678,N_2895,N_2822);
and U3679 (N_3679,N_3089,N_2627);
and U3680 (N_3680,N_2780,N_2792);
and U3681 (N_3681,N_2619,N_2954);
xnor U3682 (N_3682,N_2560,N_2814);
nand U3683 (N_3683,N_2656,N_2574);
or U3684 (N_3684,N_3111,N_3065);
nand U3685 (N_3685,N_3010,N_2662);
and U3686 (N_3686,N_2596,N_2561);
or U3687 (N_3687,N_2646,N_2578);
and U3688 (N_3688,N_2964,N_3006);
and U3689 (N_3689,N_2592,N_2777);
nor U3690 (N_3690,N_2826,N_2959);
nand U3691 (N_3691,N_2531,N_2553);
and U3692 (N_3692,N_2748,N_3015);
and U3693 (N_3693,N_2859,N_2974);
xnor U3694 (N_3694,N_2873,N_2840);
and U3695 (N_3695,N_2794,N_2743);
nand U3696 (N_3696,N_2969,N_2947);
nor U3697 (N_3697,N_3044,N_3107);
nor U3698 (N_3698,N_2537,N_2627);
or U3699 (N_3699,N_2735,N_3086);
nor U3700 (N_3700,N_2719,N_2864);
and U3701 (N_3701,N_2993,N_2621);
nand U3702 (N_3702,N_3048,N_2754);
and U3703 (N_3703,N_2564,N_2700);
nor U3704 (N_3704,N_3010,N_2927);
nand U3705 (N_3705,N_2738,N_2678);
xor U3706 (N_3706,N_3032,N_3035);
or U3707 (N_3707,N_2799,N_2911);
nand U3708 (N_3708,N_3117,N_2797);
and U3709 (N_3709,N_2869,N_2647);
nand U3710 (N_3710,N_2770,N_2759);
nor U3711 (N_3711,N_2917,N_2848);
nor U3712 (N_3712,N_2926,N_2835);
nor U3713 (N_3713,N_2507,N_2648);
nand U3714 (N_3714,N_3048,N_2876);
or U3715 (N_3715,N_2801,N_2545);
nor U3716 (N_3716,N_3048,N_2852);
or U3717 (N_3717,N_2528,N_2641);
or U3718 (N_3718,N_3110,N_2866);
and U3719 (N_3719,N_2501,N_2983);
nand U3720 (N_3720,N_3068,N_2517);
xnor U3721 (N_3721,N_2784,N_3042);
nand U3722 (N_3722,N_2899,N_3027);
or U3723 (N_3723,N_2747,N_2764);
nand U3724 (N_3724,N_2956,N_3035);
or U3725 (N_3725,N_3043,N_2628);
and U3726 (N_3726,N_2997,N_3023);
and U3727 (N_3727,N_2720,N_2821);
nor U3728 (N_3728,N_3104,N_3058);
xnor U3729 (N_3729,N_2595,N_2503);
and U3730 (N_3730,N_2909,N_2528);
and U3731 (N_3731,N_2845,N_2790);
or U3732 (N_3732,N_3058,N_2803);
nor U3733 (N_3733,N_2630,N_2813);
and U3734 (N_3734,N_2755,N_2976);
nand U3735 (N_3735,N_2599,N_2841);
and U3736 (N_3736,N_2573,N_2880);
nor U3737 (N_3737,N_2704,N_2869);
or U3738 (N_3738,N_2781,N_2735);
xor U3739 (N_3739,N_2728,N_2646);
nand U3740 (N_3740,N_2579,N_2703);
xor U3741 (N_3741,N_3015,N_3010);
nor U3742 (N_3742,N_2919,N_2970);
and U3743 (N_3743,N_2793,N_3004);
and U3744 (N_3744,N_2584,N_2598);
nor U3745 (N_3745,N_2880,N_2872);
nand U3746 (N_3746,N_2529,N_2965);
nor U3747 (N_3747,N_2737,N_3056);
nand U3748 (N_3748,N_2609,N_2810);
or U3749 (N_3749,N_2769,N_2990);
nor U3750 (N_3750,N_3639,N_3187);
nor U3751 (N_3751,N_3598,N_3228);
or U3752 (N_3752,N_3267,N_3447);
nor U3753 (N_3753,N_3180,N_3182);
and U3754 (N_3754,N_3226,N_3610);
or U3755 (N_3755,N_3464,N_3177);
xnor U3756 (N_3756,N_3149,N_3133);
and U3757 (N_3757,N_3452,N_3379);
nor U3758 (N_3758,N_3463,N_3643);
nand U3759 (N_3759,N_3481,N_3150);
nor U3760 (N_3760,N_3352,N_3293);
nor U3761 (N_3761,N_3420,N_3305);
nand U3762 (N_3762,N_3685,N_3460);
or U3763 (N_3763,N_3176,N_3551);
or U3764 (N_3764,N_3314,N_3188);
nand U3765 (N_3765,N_3148,N_3430);
nor U3766 (N_3766,N_3222,N_3327);
or U3767 (N_3767,N_3278,N_3317);
or U3768 (N_3768,N_3656,N_3241);
or U3769 (N_3769,N_3213,N_3642);
xor U3770 (N_3770,N_3545,N_3436);
or U3771 (N_3771,N_3147,N_3408);
xnor U3772 (N_3772,N_3698,N_3720);
or U3773 (N_3773,N_3345,N_3723);
nand U3774 (N_3774,N_3313,N_3662);
and U3775 (N_3775,N_3393,N_3599);
nor U3776 (N_3776,N_3494,N_3385);
nor U3777 (N_3777,N_3183,N_3312);
xor U3778 (N_3778,N_3139,N_3467);
nor U3779 (N_3779,N_3397,N_3633);
nor U3780 (N_3780,N_3570,N_3432);
or U3781 (N_3781,N_3740,N_3357);
nor U3782 (N_3782,N_3692,N_3675);
and U3783 (N_3783,N_3462,N_3636);
and U3784 (N_3784,N_3302,N_3279);
or U3785 (N_3785,N_3664,N_3324);
or U3786 (N_3786,N_3128,N_3528);
xnor U3787 (N_3787,N_3207,N_3624);
nand U3788 (N_3788,N_3678,N_3703);
nand U3789 (N_3789,N_3414,N_3632);
or U3790 (N_3790,N_3550,N_3718);
and U3791 (N_3791,N_3697,N_3287);
and U3792 (N_3792,N_3547,N_3405);
nand U3793 (N_3793,N_3355,N_3282);
and U3794 (N_3794,N_3523,N_3693);
nor U3795 (N_3795,N_3349,N_3386);
and U3796 (N_3796,N_3371,N_3295);
and U3797 (N_3797,N_3360,N_3392);
nor U3798 (N_3798,N_3660,N_3384);
nor U3799 (N_3799,N_3574,N_3377);
nand U3800 (N_3800,N_3328,N_3344);
and U3801 (N_3801,N_3529,N_3546);
nor U3802 (N_3802,N_3588,N_3509);
or U3803 (N_3803,N_3206,N_3250);
nand U3804 (N_3804,N_3567,N_3707);
or U3805 (N_3805,N_3215,N_3517);
and U3806 (N_3806,N_3332,N_3361);
nand U3807 (N_3807,N_3638,N_3419);
nor U3808 (N_3808,N_3726,N_3519);
and U3809 (N_3809,N_3434,N_3343);
nand U3810 (N_3810,N_3339,N_3614);
nor U3811 (N_3811,N_3522,N_3189);
xor U3812 (N_3812,N_3644,N_3484);
or U3813 (N_3813,N_3554,N_3508);
and U3814 (N_3814,N_3389,N_3172);
and U3815 (N_3815,N_3672,N_3158);
and U3816 (N_3816,N_3291,N_3422);
and U3817 (N_3817,N_3445,N_3260);
or U3818 (N_3818,N_3184,N_3704);
and U3819 (N_3819,N_3425,N_3671);
and U3820 (N_3820,N_3457,N_3233);
or U3821 (N_3821,N_3560,N_3333);
or U3822 (N_3822,N_3716,N_3435);
nor U3823 (N_3823,N_3504,N_3265);
and U3824 (N_3824,N_3244,N_3252);
and U3825 (N_3825,N_3364,N_3272);
nand U3826 (N_3826,N_3301,N_3347);
xor U3827 (N_3827,N_3266,N_3410);
nor U3828 (N_3828,N_3673,N_3475);
xnor U3829 (N_3829,N_3627,N_3648);
nor U3830 (N_3830,N_3261,N_3510);
or U3831 (N_3831,N_3503,N_3590);
nor U3832 (N_3832,N_3359,N_3729);
and U3833 (N_3833,N_3309,N_3251);
or U3834 (N_3834,N_3273,N_3211);
and U3835 (N_3835,N_3142,N_3380);
xor U3836 (N_3836,N_3398,N_3477);
and U3837 (N_3837,N_3695,N_3471);
and U3838 (N_3838,N_3227,N_3338);
nor U3839 (N_3839,N_3443,N_3229);
or U3840 (N_3840,N_3540,N_3466);
and U3841 (N_3841,N_3428,N_3701);
xor U3842 (N_3842,N_3369,N_3394);
nor U3843 (N_3843,N_3498,N_3195);
and U3844 (N_3844,N_3275,N_3606);
and U3845 (N_3845,N_3334,N_3442);
or U3846 (N_3846,N_3353,N_3492);
nand U3847 (N_3847,N_3595,N_3711);
or U3848 (N_3848,N_3513,N_3541);
nand U3849 (N_3849,N_3518,N_3637);
nor U3850 (N_3850,N_3308,N_3271);
nand U3851 (N_3851,N_3238,N_3247);
and U3852 (N_3852,N_3391,N_3476);
and U3853 (N_3853,N_3378,N_3179);
or U3854 (N_3854,N_3520,N_3253);
and U3855 (N_3855,N_3634,N_3444);
and U3856 (N_3856,N_3131,N_3365);
and U3857 (N_3857,N_3134,N_3322);
and U3858 (N_3858,N_3431,N_3576);
nor U3859 (N_3859,N_3363,N_3631);
nor U3860 (N_3860,N_3449,N_3555);
or U3861 (N_3861,N_3186,N_3525);
or U3862 (N_3862,N_3423,N_3502);
and U3863 (N_3863,N_3256,N_3283);
or U3864 (N_3864,N_3573,N_3416);
nand U3865 (N_3865,N_3381,N_3346);
and U3866 (N_3866,N_3412,N_3137);
nand U3867 (N_3867,N_3713,N_3127);
or U3868 (N_3868,N_3200,N_3496);
and U3869 (N_3869,N_3641,N_3246);
nor U3870 (N_3870,N_3372,N_3561);
nand U3871 (N_3871,N_3629,N_3342);
or U3872 (N_3872,N_3714,N_3126);
nor U3873 (N_3873,N_3198,N_3292);
or U3874 (N_3874,N_3375,N_3203);
nor U3875 (N_3875,N_3231,N_3712);
nor U3876 (N_3876,N_3297,N_3285);
and U3877 (N_3877,N_3699,N_3173);
nand U3878 (N_3878,N_3427,N_3132);
and U3879 (N_3879,N_3366,N_3684);
nand U3880 (N_3880,N_3592,N_3168);
and U3881 (N_3881,N_3732,N_3663);
xnor U3882 (N_3882,N_3565,N_3535);
nand U3883 (N_3883,N_3748,N_3737);
or U3884 (N_3884,N_3583,N_3415);
nor U3885 (N_3885,N_3611,N_3608);
nand U3886 (N_3886,N_3243,N_3580);
and U3887 (N_3887,N_3264,N_3609);
nor U3888 (N_3888,N_3268,N_3249);
nand U3889 (N_3889,N_3744,N_3153);
and U3890 (N_3890,N_3376,N_3601);
nand U3891 (N_3891,N_3426,N_3646);
or U3892 (N_3892,N_3532,N_3319);
and U3893 (N_3893,N_3569,N_3501);
and U3894 (N_3894,N_3387,N_3237);
nand U3895 (N_3895,N_3269,N_3482);
nand U3896 (N_3896,N_3263,N_3157);
nor U3897 (N_3897,N_3331,N_3225);
or U3898 (N_3898,N_3708,N_3474);
or U3899 (N_3899,N_3563,N_3485);
or U3900 (N_3900,N_3329,N_3669);
nand U3901 (N_3901,N_3141,N_3654);
or U3902 (N_3902,N_3557,N_3676);
nor U3903 (N_3903,N_3691,N_3323);
and U3904 (N_3904,N_3450,N_3600);
nor U3905 (N_3905,N_3196,N_3303);
nand U3906 (N_3906,N_3626,N_3356);
xor U3907 (N_3907,N_3497,N_3650);
nand U3908 (N_3908,N_3728,N_3454);
and U3909 (N_3909,N_3326,N_3719);
xor U3910 (N_3910,N_3280,N_3690);
and U3911 (N_3911,N_3505,N_3739);
xor U3912 (N_3912,N_3284,N_3539);
and U3913 (N_3913,N_3399,N_3512);
or U3914 (N_3914,N_3533,N_3245);
nor U3915 (N_3915,N_3579,N_3688);
xnor U3916 (N_3916,N_3402,N_3165);
and U3917 (N_3917,N_3706,N_3694);
nand U3918 (N_3918,N_3167,N_3162);
nor U3919 (N_3919,N_3459,N_3612);
nand U3920 (N_3920,N_3407,N_3299);
or U3921 (N_3921,N_3527,N_3479);
or U3922 (N_3922,N_3288,N_3151);
and U3923 (N_3923,N_3568,N_3204);
and U3924 (N_3924,N_3129,N_3163);
xnor U3925 (N_3925,N_3161,N_3388);
or U3926 (N_3926,N_3191,N_3613);
and U3927 (N_3927,N_3727,N_3201);
nor U3928 (N_3928,N_3155,N_3461);
or U3929 (N_3929,N_3446,N_3473);
xnor U3930 (N_3930,N_3651,N_3679);
and U3931 (N_3931,N_3236,N_3607);
nand U3932 (N_3932,N_3469,N_3337);
nor U3933 (N_3933,N_3653,N_3548);
or U3934 (N_3934,N_3506,N_3749);
nor U3935 (N_3935,N_3373,N_3438);
nor U3936 (N_3936,N_3248,N_3483);
and U3937 (N_3937,N_3559,N_3166);
nand U3938 (N_3938,N_3683,N_3530);
nor U3939 (N_3939,N_3526,N_3170);
or U3940 (N_3940,N_3586,N_3478);
and U3941 (N_3941,N_3400,N_3722);
xor U3942 (N_3942,N_3205,N_3647);
nand U3943 (N_3943,N_3370,N_3325);
xnor U3944 (N_3944,N_3175,N_3318);
and U3945 (N_3945,N_3521,N_3440);
or U3946 (N_3946,N_3138,N_3725);
nor U3947 (N_3947,N_3491,N_3310);
nor U3948 (N_3948,N_3307,N_3593);
or U3949 (N_3949,N_3731,N_3700);
nand U3950 (N_3950,N_3193,N_3255);
nand U3951 (N_3951,N_3351,N_3390);
nand U3952 (N_3952,N_3382,N_3194);
xnor U3953 (N_3953,N_3316,N_3589);
and U3954 (N_3954,N_3667,N_3232);
nand U3955 (N_3955,N_3152,N_3741);
or U3956 (N_3956,N_3709,N_3144);
nor U3957 (N_3957,N_3511,N_3680);
or U3958 (N_3958,N_3335,N_3514);
nand U3959 (N_3959,N_3321,N_3619);
xnor U3960 (N_3960,N_3686,N_3235);
nand U3961 (N_3961,N_3665,N_3689);
nor U3962 (N_3962,N_3617,N_3458);
nor U3963 (N_3963,N_3499,N_3544);
nor U3964 (N_3964,N_3635,N_3210);
nor U3965 (N_3965,N_3724,N_3217);
nand U3966 (N_3966,N_3705,N_3571);
nor U3967 (N_3967,N_3216,N_3621);
nand U3968 (N_3968,N_3262,N_3674);
or U3969 (N_3969,N_3401,N_3451);
and U3970 (N_3970,N_3738,N_3710);
and U3971 (N_3971,N_3411,N_3572);
nand U3972 (N_3972,N_3336,N_3413);
nor U3973 (N_3973,N_3625,N_3224);
nor U3974 (N_3974,N_3300,N_3218);
xnor U3975 (N_3975,N_3585,N_3298);
nor U3976 (N_3976,N_3696,N_3668);
nand U3977 (N_3977,N_3330,N_3556);
or U3978 (N_3978,N_3618,N_3296);
and U3979 (N_3979,N_3362,N_3136);
nor U3980 (N_3980,N_3418,N_3562);
and U3981 (N_3981,N_3615,N_3178);
or U3982 (N_3982,N_3742,N_3597);
nand U3983 (N_3983,N_3240,N_3156);
and U3984 (N_3984,N_3659,N_3320);
or U3985 (N_3985,N_3367,N_3197);
nor U3986 (N_3986,N_3487,N_3290);
xnor U3987 (N_3987,N_3396,N_3682);
xor U3988 (N_3988,N_3181,N_3630);
and U3989 (N_3989,N_3140,N_3395);
or U3990 (N_3990,N_3456,N_3677);
nand U3991 (N_3991,N_3577,N_3439);
or U3992 (N_3992,N_3645,N_3605);
or U3993 (N_3993,N_3259,N_3640);
xnor U3994 (N_3994,N_3208,N_3745);
and U3995 (N_3995,N_3406,N_3721);
or U3996 (N_3996,N_3516,N_3274);
nor U3997 (N_3997,N_3135,N_3587);
nor U3998 (N_3998,N_3164,N_3537);
and U3999 (N_3999,N_3169,N_3202);
or U4000 (N_4000,N_3566,N_3223);
nor U4001 (N_4001,N_3733,N_3214);
and U4002 (N_4002,N_3616,N_3421);
nand U4003 (N_4003,N_3289,N_3277);
xnor U4004 (N_4004,N_3130,N_3582);
or U4005 (N_4005,N_3424,N_3455);
xor U4006 (N_4006,N_3154,N_3437);
and U4007 (N_4007,N_3661,N_3486);
and U4008 (N_4008,N_3687,N_3276);
nor U4009 (N_4009,N_3220,N_3575);
or U4010 (N_4010,N_3604,N_3649);
xnor U4011 (N_4011,N_3374,N_3143);
and U4012 (N_4012,N_3340,N_3159);
and U4013 (N_4013,N_3531,N_3468);
nor U4014 (N_4014,N_3652,N_3603);
or U4015 (N_4015,N_3500,N_3311);
and U4016 (N_4016,N_3534,N_3242);
nor U4017 (N_4017,N_3552,N_3596);
nand U4018 (N_4018,N_3542,N_3146);
or U4019 (N_4019,N_3348,N_3623);
or U4020 (N_4020,N_3453,N_3591);
or U4021 (N_4021,N_3524,N_3234);
and U4022 (N_4022,N_3304,N_3239);
nor U4023 (N_4023,N_3145,N_3581);
nor U4024 (N_4024,N_3441,N_3209);
or U4025 (N_4025,N_3409,N_3306);
or U4026 (N_4026,N_3199,N_3746);
or U4027 (N_4027,N_3558,N_3417);
and U4028 (N_4028,N_3472,N_3602);
nor U4029 (N_4029,N_3350,N_3507);
nand U4030 (N_4030,N_3354,N_3553);
nor U4031 (N_4031,N_3254,N_3125);
xor U4032 (N_4032,N_3717,N_3358);
or U4033 (N_4033,N_3192,N_3270);
and U4034 (N_4034,N_3230,N_3564);
and U4035 (N_4035,N_3536,N_3429);
nand U4036 (N_4036,N_3489,N_3383);
nand U4037 (N_4037,N_3730,N_3190);
nand U4038 (N_4038,N_3171,N_3403);
nor U4039 (N_4039,N_3221,N_3655);
nor U4040 (N_4040,N_3465,N_3620);
or U4041 (N_4041,N_3433,N_3736);
nor U4042 (N_4042,N_3578,N_3702);
nand U4043 (N_4043,N_3480,N_3743);
and U4044 (N_4044,N_3258,N_3515);
or U4045 (N_4045,N_3670,N_3549);
nor U4046 (N_4046,N_3493,N_3490);
and U4047 (N_4047,N_3448,N_3257);
or U4048 (N_4048,N_3495,N_3734);
nor U4049 (N_4049,N_3543,N_3735);
and U4050 (N_4050,N_3404,N_3212);
and U4051 (N_4051,N_3628,N_3315);
nor U4052 (N_4052,N_3666,N_3281);
nand U4053 (N_4053,N_3584,N_3368);
nand U4054 (N_4054,N_3747,N_3160);
nor U4055 (N_4055,N_3594,N_3488);
or U4056 (N_4056,N_3185,N_3538);
nor U4057 (N_4057,N_3715,N_3341);
nand U4058 (N_4058,N_3174,N_3219);
and U4059 (N_4059,N_3658,N_3622);
nor U4060 (N_4060,N_3294,N_3681);
and U4061 (N_4061,N_3657,N_3470);
nand U4062 (N_4062,N_3286,N_3246);
xor U4063 (N_4063,N_3446,N_3582);
and U4064 (N_4064,N_3229,N_3633);
xor U4065 (N_4065,N_3144,N_3681);
nand U4066 (N_4066,N_3521,N_3520);
or U4067 (N_4067,N_3273,N_3193);
nor U4068 (N_4068,N_3228,N_3654);
nand U4069 (N_4069,N_3573,N_3127);
or U4070 (N_4070,N_3233,N_3172);
nand U4071 (N_4071,N_3211,N_3590);
xor U4072 (N_4072,N_3496,N_3439);
nand U4073 (N_4073,N_3634,N_3638);
or U4074 (N_4074,N_3583,N_3543);
nor U4075 (N_4075,N_3742,N_3586);
xnor U4076 (N_4076,N_3291,N_3429);
or U4077 (N_4077,N_3372,N_3454);
and U4078 (N_4078,N_3476,N_3253);
or U4079 (N_4079,N_3165,N_3537);
nand U4080 (N_4080,N_3239,N_3392);
xor U4081 (N_4081,N_3671,N_3744);
nor U4082 (N_4082,N_3187,N_3286);
or U4083 (N_4083,N_3335,N_3620);
and U4084 (N_4084,N_3137,N_3178);
and U4085 (N_4085,N_3392,N_3526);
xnor U4086 (N_4086,N_3332,N_3549);
or U4087 (N_4087,N_3375,N_3732);
xor U4088 (N_4088,N_3322,N_3367);
and U4089 (N_4089,N_3717,N_3397);
and U4090 (N_4090,N_3586,N_3585);
or U4091 (N_4091,N_3726,N_3598);
nor U4092 (N_4092,N_3351,N_3501);
or U4093 (N_4093,N_3592,N_3305);
and U4094 (N_4094,N_3228,N_3460);
and U4095 (N_4095,N_3431,N_3390);
nand U4096 (N_4096,N_3461,N_3147);
or U4097 (N_4097,N_3519,N_3170);
nor U4098 (N_4098,N_3362,N_3695);
and U4099 (N_4099,N_3645,N_3290);
and U4100 (N_4100,N_3398,N_3125);
and U4101 (N_4101,N_3288,N_3444);
and U4102 (N_4102,N_3394,N_3711);
nand U4103 (N_4103,N_3414,N_3614);
xor U4104 (N_4104,N_3210,N_3214);
and U4105 (N_4105,N_3402,N_3715);
nand U4106 (N_4106,N_3562,N_3657);
nor U4107 (N_4107,N_3492,N_3673);
nor U4108 (N_4108,N_3517,N_3746);
and U4109 (N_4109,N_3560,N_3129);
and U4110 (N_4110,N_3186,N_3346);
nand U4111 (N_4111,N_3164,N_3154);
nor U4112 (N_4112,N_3222,N_3599);
or U4113 (N_4113,N_3338,N_3615);
and U4114 (N_4114,N_3231,N_3748);
xor U4115 (N_4115,N_3147,N_3433);
nand U4116 (N_4116,N_3389,N_3413);
nor U4117 (N_4117,N_3746,N_3299);
and U4118 (N_4118,N_3701,N_3293);
and U4119 (N_4119,N_3319,N_3210);
xnor U4120 (N_4120,N_3317,N_3507);
and U4121 (N_4121,N_3742,N_3554);
and U4122 (N_4122,N_3600,N_3271);
or U4123 (N_4123,N_3327,N_3584);
and U4124 (N_4124,N_3477,N_3715);
nand U4125 (N_4125,N_3129,N_3278);
nand U4126 (N_4126,N_3348,N_3126);
or U4127 (N_4127,N_3394,N_3247);
nor U4128 (N_4128,N_3333,N_3746);
or U4129 (N_4129,N_3150,N_3353);
nor U4130 (N_4130,N_3466,N_3290);
or U4131 (N_4131,N_3416,N_3718);
nor U4132 (N_4132,N_3482,N_3564);
or U4133 (N_4133,N_3237,N_3653);
nand U4134 (N_4134,N_3254,N_3426);
or U4135 (N_4135,N_3209,N_3321);
nor U4136 (N_4136,N_3400,N_3704);
and U4137 (N_4137,N_3589,N_3256);
or U4138 (N_4138,N_3213,N_3159);
and U4139 (N_4139,N_3236,N_3348);
xor U4140 (N_4140,N_3646,N_3526);
xor U4141 (N_4141,N_3305,N_3539);
or U4142 (N_4142,N_3472,N_3366);
and U4143 (N_4143,N_3698,N_3585);
or U4144 (N_4144,N_3641,N_3205);
and U4145 (N_4145,N_3423,N_3433);
nand U4146 (N_4146,N_3174,N_3668);
nand U4147 (N_4147,N_3229,N_3496);
nand U4148 (N_4148,N_3240,N_3404);
or U4149 (N_4149,N_3671,N_3329);
nor U4150 (N_4150,N_3523,N_3421);
and U4151 (N_4151,N_3610,N_3578);
and U4152 (N_4152,N_3696,N_3607);
nand U4153 (N_4153,N_3503,N_3738);
xnor U4154 (N_4154,N_3132,N_3393);
or U4155 (N_4155,N_3680,N_3623);
and U4156 (N_4156,N_3317,N_3243);
and U4157 (N_4157,N_3293,N_3315);
nand U4158 (N_4158,N_3391,N_3607);
and U4159 (N_4159,N_3661,N_3158);
nor U4160 (N_4160,N_3192,N_3290);
nand U4161 (N_4161,N_3193,N_3660);
nand U4162 (N_4162,N_3497,N_3314);
nand U4163 (N_4163,N_3544,N_3670);
or U4164 (N_4164,N_3688,N_3192);
and U4165 (N_4165,N_3714,N_3728);
nor U4166 (N_4166,N_3634,N_3210);
and U4167 (N_4167,N_3696,N_3664);
xor U4168 (N_4168,N_3267,N_3681);
and U4169 (N_4169,N_3193,N_3395);
nor U4170 (N_4170,N_3454,N_3613);
and U4171 (N_4171,N_3625,N_3536);
and U4172 (N_4172,N_3191,N_3233);
and U4173 (N_4173,N_3561,N_3413);
and U4174 (N_4174,N_3734,N_3239);
and U4175 (N_4175,N_3615,N_3217);
and U4176 (N_4176,N_3586,N_3253);
nor U4177 (N_4177,N_3336,N_3743);
nand U4178 (N_4178,N_3286,N_3545);
nand U4179 (N_4179,N_3419,N_3437);
nor U4180 (N_4180,N_3543,N_3636);
nand U4181 (N_4181,N_3367,N_3351);
or U4182 (N_4182,N_3571,N_3209);
and U4183 (N_4183,N_3546,N_3656);
or U4184 (N_4184,N_3527,N_3254);
and U4185 (N_4185,N_3273,N_3155);
nand U4186 (N_4186,N_3598,N_3256);
nor U4187 (N_4187,N_3219,N_3273);
nor U4188 (N_4188,N_3495,N_3307);
xor U4189 (N_4189,N_3658,N_3500);
xor U4190 (N_4190,N_3265,N_3603);
nand U4191 (N_4191,N_3378,N_3583);
nor U4192 (N_4192,N_3381,N_3317);
nand U4193 (N_4193,N_3481,N_3698);
or U4194 (N_4194,N_3410,N_3231);
or U4195 (N_4195,N_3202,N_3561);
xnor U4196 (N_4196,N_3196,N_3455);
nor U4197 (N_4197,N_3558,N_3574);
nand U4198 (N_4198,N_3471,N_3137);
nor U4199 (N_4199,N_3189,N_3549);
nand U4200 (N_4200,N_3741,N_3600);
or U4201 (N_4201,N_3190,N_3745);
nor U4202 (N_4202,N_3717,N_3569);
and U4203 (N_4203,N_3480,N_3349);
and U4204 (N_4204,N_3382,N_3593);
or U4205 (N_4205,N_3410,N_3741);
or U4206 (N_4206,N_3348,N_3231);
xnor U4207 (N_4207,N_3676,N_3645);
or U4208 (N_4208,N_3463,N_3511);
nor U4209 (N_4209,N_3727,N_3178);
nand U4210 (N_4210,N_3480,N_3211);
xnor U4211 (N_4211,N_3595,N_3220);
or U4212 (N_4212,N_3562,N_3316);
and U4213 (N_4213,N_3514,N_3373);
nor U4214 (N_4214,N_3523,N_3703);
or U4215 (N_4215,N_3692,N_3154);
and U4216 (N_4216,N_3728,N_3607);
and U4217 (N_4217,N_3251,N_3682);
nor U4218 (N_4218,N_3726,N_3516);
and U4219 (N_4219,N_3179,N_3445);
and U4220 (N_4220,N_3643,N_3357);
or U4221 (N_4221,N_3558,N_3622);
xor U4222 (N_4222,N_3656,N_3376);
and U4223 (N_4223,N_3744,N_3147);
nand U4224 (N_4224,N_3615,N_3314);
xor U4225 (N_4225,N_3556,N_3225);
or U4226 (N_4226,N_3491,N_3187);
nand U4227 (N_4227,N_3530,N_3235);
or U4228 (N_4228,N_3606,N_3358);
and U4229 (N_4229,N_3391,N_3367);
nand U4230 (N_4230,N_3641,N_3701);
or U4231 (N_4231,N_3498,N_3209);
nor U4232 (N_4232,N_3443,N_3149);
xnor U4233 (N_4233,N_3495,N_3201);
nand U4234 (N_4234,N_3661,N_3299);
nand U4235 (N_4235,N_3543,N_3492);
and U4236 (N_4236,N_3666,N_3672);
xnor U4237 (N_4237,N_3356,N_3504);
xnor U4238 (N_4238,N_3388,N_3287);
or U4239 (N_4239,N_3652,N_3372);
nor U4240 (N_4240,N_3156,N_3727);
or U4241 (N_4241,N_3547,N_3586);
xnor U4242 (N_4242,N_3391,N_3232);
nor U4243 (N_4243,N_3677,N_3253);
or U4244 (N_4244,N_3295,N_3345);
nand U4245 (N_4245,N_3340,N_3562);
or U4246 (N_4246,N_3281,N_3705);
nand U4247 (N_4247,N_3268,N_3749);
nand U4248 (N_4248,N_3248,N_3206);
nor U4249 (N_4249,N_3393,N_3310);
and U4250 (N_4250,N_3403,N_3633);
nand U4251 (N_4251,N_3363,N_3343);
or U4252 (N_4252,N_3526,N_3722);
and U4253 (N_4253,N_3236,N_3468);
nand U4254 (N_4254,N_3306,N_3569);
or U4255 (N_4255,N_3440,N_3603);
and U4256 (N_4256,N_3562,N_3180);
nand U4257 (N_4257,N_3211,N_3346);
and U4258 (N_4258,N_3313,N_3501);
or U4259 (N_4259,N_3546,N_3691);
xor U4260 (N_4260,N_3669,N_3249);
nor U4261 (N_4261,N_3221,N_3204);
or U4262 (N_4262,N_3679,N_3278);
nor U4263 (N_4263,N_3323,N_3544);
and U4264 (N_4264,N_3393,N_3286);
and U4265 (N_4265,N_3337,N_3535);
and U4266 (N_4266,N_3199,N_3251);
or U4267 (N_4267,N_3310,N_3600);
nor U4268 (N_4268,N_3420,N_3184);
nand U4269 (N_4269,N_3386,N_3429);
or U4270 (N_4270,N_3684,N_3632);
nand U4271 (N_4271,N_3334,N_3615);
or U4272 (N_4272,N_3691,N_3376);
and U4273 (N_4273,N_3524,N_3492);
or U4274 (N_4274,N_3597,N_3569);
nor U4275 (N_4275,N_3138,N_3444);
or U4276 (N_4276,N_3464,N_3721);
and U4277 (N_4277,N_3603,N_3500);
or U4278 (N_4278,N_3187,N_3142);
nor U4279 (N_4279,N_3462,N_3220);
nand U4280 (N_4280,N_3405,N_3749);
nand U4281 (N_4281,N_3629,N_3375);
nand U4282 (N_4282,N_3268,N_3170);
and U4283 (N_4283,N_3646,N_3336);
or U4284 (N_4284,N_3590,N_3746);
or U4285 (N_4285,N_3241,N_3449);
nand U4286 (N_4286,N_3559,N_3591);
nor U4287 (N_4287,N_3186,N_3273);
and U4288 (N_4288,N_3373,N_3443);
nand U4289 (N_4289,N_3697,N_3403);
nand U4290 (N_4290,N_3454,N_3167);
nor U4291 (N_4291,N_3482,N_3336);
or U4292 (N_4292,N_3407,N_3516);
nor U4293 (N_4293,N_3206,N_3488);
or U4294 (N_4294,N_3747,N_3672);
or U4295 (N_4295,N_3473,N_3139);
or U4296 (N_4296,N_3564,N_3426);
nor U4297 (N_4297,N_3467,N_3181);
and U4298 (N_4298,N_3551,N_3284);
nor U4299 (N_4299,N_3212,N_3354);
nor U4300 (N_4300,N_3377,N_3271);
nor U4301 (N_4301,N_3413,N_3195);
xor U4302 (N_4302,N_3549,N_3160);
xor U4303 (N_4303,N_3288,N_3372);
and U4304 (N_4304,N_3430,N_3528);
nand U4305 (N_4305,N_3606,N_3404);
nor U4306 (N_4306,N_3733,N_3136);
nand U4307 (N_4307,N_3319,N_3143);
nand U4308 (N_4308,N_3129,N_3745);
nand U4309 (N_4309,N_3720,N_3268);
nor U4310 (N_4310,N_3287,N_3258);
and U4311 (N_4311,N_3229,N_3181);
or U4312 (N_4312,N_3284,N_3152);
and U4313 (N_4313,N_3707,N_3163);
or U4314 (N_4314,N_3146,N_3582);
or U4315 (N_4315,N_3671,N_3674);
and U4316 (N_4316,N_3161,N_3470);
or U4317 (N_4317,N_3639,N_3512);
nand U4318 (N_4318,N_3590,N_3191);
nor U4319 (N_4319,N_3468,N_3430);
and U4320 (N_4320,N_3380,N_3660);
or U4321 (N_4321,N_3610,N_3630);
and U4322 (N_4322,N_3221,N_3573);
nand U4323 (N_4323,N_3738,N_3305);
and U4324 (N_4324,N_3624,N_3534);
or U4325 (N_4325,N_3733,N_3684);
nor U4326 (N_4326,N_3683,N_3153);
nor U4327 (N_4327,N_3596,N_3572);
xnor U4328 (N_4328,N_3643,N_3303);
and U4329 (N_4329,N_3697,N_3435);
and U4330 (N_4330,N_3648,N_3420);
nor U4331 (N_4331,N_3620,N_3479);
or U4332 (N_4332,N_3134,N_3414);
nand U4333 (N_4333,N_3320,N_3744);
or U4334 (N_4334,N_3429,N_3685);
nand U4335 (N_4335,N_3668,N_3218);
or U4336 (N_4336,N_3678,N_3650);
nor U4337 (N_4337,N_3617,N_3269);
nor U4338 (N_4338,N_3332,N_3219);
xnor U4339 (N_4339,N_3366,N_3652);
nand U4340 (N_4340,N_3219,N_3650);
or U4341 (N_4341,N_3182,N_3279);
and U4342 (N_4342,N_3251,N_3688);
and U4343 (N_4343,N_3163,N_3307);
xor U4344 (N_4344,N_3466,N_3503);
and U4345 (N_4345,N_3334,N_3337);
xnor U4346 (N_4346,N_3215,N_3154);
nor U4347 (N_4347,N_3518,N_3669);
xor U4348 (N_4348,N_3749,N_3228);
nor U4349 (N_4349,N_3461,N_3125);
or U4350 (N_4350,N_3710,N_3281);
nor U4351 (N_4351,N_3488,N_3269);
nor U4352 (N_4352,N_3142,N_3697);
or U4353 (N_4353,N_3292,N_3171);
nor U4354 (N_4354,N_3257,N_3241);
nand U4355 (N_4355,N_3606,N_3362);
nor U4356 (N_4356,N_3692,N_3204);
and U4357 (N_4357,N_3257,N_3683);
xor U4358 (N_4358,N_3284,N_3279);
and U4359 (N_4359,N_3265,N_3744);
xor U4360 (N_4360,N_3161,N_3372);
nor U4361 (N_4361,N_3271,N_3436);
nand U4362 (N_4362,N_3720,N_3140);
nand U4363 (N_4363,N_3515,N_3335);
nor U4364 (N_4364,N_3294,N_3432);
nor U4365 (N_4365,N_3599,N_3469);
or U4366 (N_4366,N_3355,N_3407);
or U4367 (N_4367,N_3589,N_3698);
and U4368 (N_4368,N_3468,N_3552);
nor U4369 (N_4369,N_3719,N_3426);
nor U4370 (N_4370,N_3173,N_3641);
nor U4371 (N_4371,N_3378,N_3424);
xnor U4372 (N_4372,N_3530,N_3429);
nor U4373 (N_4373,N_3608,N_3294);
nor U4374 (N_4374,N_3384,N_3546);
or U4375 (N_4375,N_4123,N_3867);
xnor U4376 (N_4376,N_4179,N_3959);
nand U4377 (N_4377,N_4020,N_4274);
or U4378 (N_4378,N_3995,N_4358);
or U4379 (N_4379,N_4226,N_4026);
nor U4380 (N_4380,N_4202,N_3869);
nand U4381 (N_4381,N_4366,N_4253);
and U4382 (N_4382,N_3899,N_4332);
nand U4383 (N_4383,N_3921,N_3793);
and U4384 (N_4384,N_3883,N_4003);
or U4385 (N_4385,N_4095,N_4014);
and U4386 (N_4386,N_4067,N_4133);
and U4387 (N_4387,N_4333,N_3879);
xor U4388 (N_4388,N_3754,N_3837);
nand U4389 (N_4389,N_4197,N_4359);
xnor U4390 (N_4390,N_3827,N_4374);
nand U4391 (N_4391,N_4069,N_3884);
nor U4392 (N_4392,N_3839,N_4278);
or U4393 (N_4393,N_3777,N_3902);
nand U4394 (N_4394,N_4127,N_4313);
and U4395 (N_4395,N_4032,N_4171);
nand U4396 (N_4396,N_4331,N_3911);
or U4397 (N_4397,N_4025,N_3949);
and U4398 (N_4398,N_4311,N_4183);
nand U4399 (N_4399,N_4009,N_4206);
or U4400 (N_4400,N_4010,N_4364);
or U4401 (N_4401,N_3938,N_3752);
nand U4402 (N_4402,N_3922,N_3954);
or U4403 (N_4403,N_4157,N_4156);
nand U4404 (N_4404,N_3891,N_4022);
and U4405 (N_4405,N_3905,N_4262);
nand U4406 (N_4406,N_4139,N_3831);
or U4407 (N_4407,N_4212,N_4237);
nor U4408 (N_4408,N_4135,N_3858);
nand U4409 (N_4409,N_3943,N_3807);
and U4410 (N_4410,N_3835,N_3920);
and U4411 (N_4411,N_3800,N_4343);
nor U4412 (N_4412,N_4265,N_3773);
and U4413 (N_4413,N_3889,N_4070);
nor U4414 (N_4414,N_4349,N_3951);
nand U4415 (N_4415,N_3814,N_3989);
nor U4416 (N_4416,N_4338,N_4074);
xor U4417 (N_4417,N_3763,N_3919);
nor U4418 (N_4418,N_4007,N_4341);
nand U4419 (N_4419,N_4131,N_3770);
or U4420 (N_4420,N_4002,N_3799);
or U4421 (N_4421,N_3974,N_4292);
or U4422 (N_4422,N_3817,N_3767);
or U4423 (N_4423,N_3782,N_4172);
or U4424 (N_4424,N_4016,N_3964);
xor U4425 (N_4425,N_4094,N_4117);
nand U4426 (N_4426,N_3930,N_4239);
nor U4427 (N_4427,N_4231,N_4120);
and U4428 (N_4428,N_4291,N_3977);
nand U4429 (N_4429,N_4255,N_4245);
xor U4430 (N_4430,N_4177,N_4254);
and U4431 (N_4431,N_4325,N_3789);
and U4432 (N_4432,N_4097,N_4057);
or U4433 (N_4433,N_4270,N_4115);
or U4434 (N_4434,N_4147,N_4145);
nand U4435 (N_4435,N_4090,N_4207);
and U4436 (N_4436,N_3790,N_4164);
nand U4437 (N_4437,N_4196,N_4345);
nor U4438 (N_4438,N_4160,N_4142);
nand U4439 (N_4439,N_4089,N_4114);
or U4440 (N_4440,N_3804,N_4034);
or U4441 (N_4441,N_4299,N_4310);
nor U4442 (N_4442,N_4042,N_4283);
nor U4443 (N_4443,N_3998,N_4256);
nor U4444 (N_4444,N_3841,N_4109);
or U4445 (N_4445,N_3874,N_4031);
nand U4446 (N_4446,N_3971,N_3776);
or U4447 (N_4447,N_4213,N_3960);
nor U4448 (N_4448,N_4252,N_3872);
or U4449 (N_4449,N_3957,N_4087);
or U4450 (N_4450,N_3941,N_4223);
nor U4451 (N_4451,N_3882,N_4225);
or U4452 (N_4452,N_4055,N_3991);
nor U4453 (N_4453,N_4339,N_3842);
or U4454 (N_4454,N_4039,N_3870);
and U4455 (N_4455,N_4280,N_4054);
nor U4456 (N_4456,N_4173,N_3927);
nand U4457 (N_4457,N_3986,N_4049);
and U4458 (N_4458,N_4232,N_3942);
xor U4459 (N_4459,N_3893,N_3918);
nand U4460 (N_4460,N_3791,N_4065);
nor U4461 (N_4461,N_3945,N_4053);
or U4462 (N_4462,N_3979,N_3786);
xnor U4463 (N_4463,N_4084,N_4050);
and U4464 (N_4464,N_3952,N_3908);
and U4465 (N_4465,N_4104,N_4106);
or U4466 (N_4466,N_4161,N_4222);
nor U4467 (N_4467,N_3821,N_3778);
or U4468 (N_4468,N_3751,N_4337);
or U4469 (N_4469,N_4352,N_3912);
and U4470 (N_4470,N_4201,N_4144);
nor U4471 (N_4471,N_4368,N_4129);
nor U4472 (N_4472,N_4308,N_3826);
and U4473 (N_4473,N_4085,N_3833);
or U4474 (N_4474,N_4344,N_3864);
or U4475 (N_4475,N_4361,N_3997);
and U4476 (N_4476,N_4059,N_3978);
or U4477 (N_4477,N_4019,N_4121);
or U4478 (N_4478,N_3990,N_4346);
or U4479 (N_4479,N_4169,N_4249);
nand U4480 (N_4480,N_3823,N_4351);
nand U4481 (N_4481,N_4219,N_3885);
or U4482 (N_4482,N_4367,N_4282);
or U4483 (N_4483,N_3876,N_3802);
xnor U4484 (N_4484,N_4218,N_3788);
nor U4485 (N_4485,N_3753,N_4152);
or U4486 (N_4486,N_4108,N_3853);
or U4487 (N_4487,N_4111,N_4369);
nand U4488 (N_4488,N_4304,N_3984);
or U4489 (N_4489,N_3828,N_4174);
nor U4490 (N_4490,N_4190,N_4229);
nor U4491 (N_4491,N_3796,N_3987);
or U4492 (N_4492,N_3822,N_4098);
and U4493 (N_4493,N_4058,N_3975);
or U4494 (N_4494,N_4072,N_4321);
and U4495 (N_4495,N_4008,N_4113);
and U4496 (N_4496,N_3969,N_3848);
nand U4497 (N_4497,N_4241,N_4167);
xnor U4498 (N_4498,N_3966,N_4228);
nand U4499 (N_4499,N_3967,N_3985);
and U4500 (N_4500,N_4363,N_4146);
nor U4501 (N_4501,N_3774,N_3963);
or U4502 (N_4502,N_4078,N_4182);
nor U4503 (N_4503,N_4051,N_3801);
and U4504 (N_4504,N_3897,N_3926);
nor U4505 (N_4505,N_4315,N_3878);
nor U4506 (N_4506,N_4040,N_4186);
nand U4507 (N_4507,N_4302,N_4119);
nand U4508 (N_4508,N_4150,N_4336);
xor U4509 (N_4509,N_4200,N_3898);
and U4510 (N_4510,N_4091,N_4236);
nor U4511 (N_4511,N_3760,N_3944);
and U4512 (N_4512,N_4356,N_3787);
nand U4513 (N_4513,N_3937,N_4261);
or U4514 (N_4514,N_3907,N_4300);
or U4515 (N_4515,N_3766,N_4163);
or U4516 (N_4516,N_4077,N_4083);
or U4517 (N_4517,N_4134,N_4162);
nor U4518 (N_4518,N_3913,N_4248);
or U4519 (N_4519,N_4357,N_3772);
xnor U4520 (N_4520,N_3815,N_4092);
nor U4521 (N_4521,N_4191,N_3946);
and U4522 (N_4522,N_3909,N_3780);
or U4523 (N_4523,N_3843,N_3775);
nand U4524 (N_4524,N_3803,N_4317);
nand U4525 (N_4525,N_4000,N_4056);
nor U4526 (N_4526,N_4189,N_3820);
nor U4527 (N_4527,N_4244,N_4187);
nand U4528 (N_4528,N_4220,N_3762);
nand U4529 (N_4529,N_3765,N_4012);
or U4530 (N_4530,N_4260,N_4132);
nand U4531 (N_4531,N_3769,N_3994);
nand U4532 (N_4532,N_4021,N_4140);
or U4533 (N_4533,N_4073,N_4159);
nor U4534 (N_4534,N_3976,N_3759);
and U4535 (N_4535,N_4296,N_3890);
xnor U4536 (N_4536,N_3866,N_3955);
and U4537 (N_4537,N_4100,N_3813);
nand U4538 (N_4538,N_4041,N_4024);
nor U4539 (N_4539,N_4234,N_4326);
or U4540 (N_4540,N_4214,N_3923);
or U4541 (N_4541,N_3939,N_4118);
nor U4542 (N_4542,N_4284,N_4099);
and U4543 (N_4543,N_3901,N_4038);
nor U4544 (N_4544,N_4355,N_4168);
and U4545 (N_4545,N_3917,N_4347);
nand U4546 (N_4546,N_4153,N_4075);
nand U4547 (N_4547,N_4045,N_4327);
nor U4548 (N_4548,N_4175,N_3850);
or U4549 (N_4549,N_3940,N_4210);
and U4550 (N_4550,N_3904,N_4030);
and U4551 (N_4551,N_4081,N_4107);
nand U4552 (N_4552,N_4350,N_4303);
xnor U4553 (N_4553,N_4348,N_4126);
or U4554 (N_4554,N_3755,N_4060);
or U4555 (N_4555,N_4063,N_3906);
and U4556 (N_4556,N_4093,N_4110);
xnor U4557 (N_4557,N_3834,N_4312);
nor U4558 (N_4558,N_3849,N_4329);
and U4559 (N_4559,N_3925,N_4103);
nor U4560 (N_4560,N_4243,N_3900);
nor U4561 (N_4561,N_4068,N_4340);
and U4562 (N_4562,N_4166,N_4216);
or U4563 (N_4563,N_4155,N_4240);
nand U4564 (N_4564,N_4086,N_3914);
nand U4565 (N_4565,N_3862,N_3851);
or U4566 (N_4566,N_4136,N_4023);
and U4567 (N_4567,N_3783,N_4354);
or U4568 (N_4568,N_4297,N_3924);
nand U4569 (N_4569,N_4076,N_4288);
xor U4570 (N_4570,N_4365,N_3928);
nor U4571 (N_4571,N_3825,N_4047);
nand U4572 (N_4572,N_4215,N_3805);
xnor U4573 (N_4573,N_3797,N_3916);
xor U4574 (N_4574,N_4180,N_4029);
or U4575 (N_4575,N_4017,N_4044);
or U4576 (N_4576,N_4247,N_4185);
xnor U4577 (N_4577,N_4246,N_4165);
nor U4578 (N_4578,N_3947,N_4148);
nor U4579 (N_4579,N_4143,N_3996);
nor U4580 (N_4580,N_4273,N_3950);
or U4581 (N_4581,N_4353,N_4211);
nor U4582 (N_4582,N_3962,N_4004);
nor U4583 (N_4583,N_4170,N_3761);
nor U4584 (N_4584,N_4001,N_3794);
xor U4585 (N_4585,N_4046,N_3953);
xor U4586 (N_4586,N_3896,N_4124);
or U4587 (N_4587,N_4360,N_4221);
nor U4588 (N_4588,N_3811,N_4322);
xor U4589 (N_4589,N_4285,N_3968);
nor U4590 (N_4590,N_3829,N_4289);
xnor U4591 (N_4591,N_3750,N_4372);
or U4592 (N_4592,N_3856,N_4209);
or U4593 (N_4593,N_4251,N_4176);
nor U4594 (N_4594,N_3863,N_4275);
xor U4595 (N_4595,N_4192,N_4027);
and U4596 (N_4596,N_4141,N_3880);
nand U4597 (N_4597,N_3808,N_4006);
nor U4598 (N_4598,N_3792,N_4370);
and U4599 (N_4599,N_4316,N_3781);
or U4600 (N_4600,N_4307,N_4328);
nand U4601 (N_4601,N_4264,N_4323);
xor U4602 (N_4602,N_4324,N_3903);
and U4603 (N_4603,N_3973,N_3993);
nand U4604 (N_4604,N_4263,N_4224);
or U4605 (N_4605,N_4309,N_4235);
xor U4606 (N_4606,N_4102,N_4018);
nand U4607 (N_4607,N_3795,N_4005);
nor U4608 (N_4608,N_4314,N_4305);
nand U4609 (N_4609,N_4293,N_4306);
xor U4610 (N_4610,N_3809,N_3875);
nor U4611 (N_4611,N_3857,N_4335);
or U4612 (N_4612,N_4362,N_3806);
or U4613 (N_4613,N_4330,N_4154);
nor U4614 (N_4614,N_4178,N_4062);
or U4615 (N_4615,N_4258,N_3840);
and U4616 (N_4616,N_4277,N_3865);
nand U4617 (N_4617,N_4112,N_3934);
nor U4618 (N_4618,N_4061,N_3886);
or U4619 (N_4619,N_3956,N_3816);
xnor U4620 (N_4620,N_3784,N_3881);
and U4621 (N_4621,N_3892,N_4188);
or U4622 (N_4622,N_4373,N_4208);
or U4623 (N_4623,N_3948,N_4204);
and U4624 (N_4624,N_4071,N_3818);
nor U4625 (N_4625,N_4088,N_3972);
xor U4626 (N_4626,N_4272,N_3758);
and U4627 (N_4627,N_4266,N_4319);
and U4628 (N_4628,N_4194,N_4130);
nor U4629 (N_4629,N_3868,N_4257);
or U4630 (N_4630,N_3982,N_3757);
and U4631 (N_4631,N_4294,N_4199);
nor U4632 (N_4632,N_3873,N_4230);
xor U4633 (N_4633,N_4043,N_4082);
nand U4634 (N_4634,N_3965,N_3983);
nor U4635 (N_4635,N_4203,N_3970);
and U4636 (N_4636,N_3838,N_3824);
and U4637 (N_4637,N_4125,N_4064);
and U4638 (N_4638,N_3819,N_4320);
and U4639 (N_4639,N_4105,N_3861);
or U4640 (N_4640,N_3798,N_4334);
and U4641 (N_4641,N_4036,N_3771);
and U4642 (N_4642,N_3845,N_3785);
xnor U4643 (N_4643,N_4279,N_4122);
and U4644 (N_4644,N_4015,N_4301);
nand U4645 (N_4645,N_3832,N_3895);
or U4646 (N_4646,N_4268,N_4198);
or U4647 (N_4647,N_3932,N_4101);
or U4648 (N_4648,N_4151,N_3846);
xnor U4649 (N_4649,N_4227,N_4116);
or U4650 (N_4650,N_3981,N_3929);
and U4651 (N_4651,N_4138,N_3859);
or U4652 (N_4652,N_3992,N_4267);
nor U4653 (N_4653,N_4013,N_3830);
nor U4654 (N_4654,N_4096,N_3844);
and U4655 (N_4655,N_4048,N_4137);
xor U4656 (N_4656,N_4181,N_4080);
nor U4657 (N_4657,N_3958,N_4052);
nor U4658 (N_4658,N_4033,N_3768);
or U4659 (N_4659,N_4158,N_4271);
or U4660 (N_4660,N_4184,N_3961);
and U4661 (N_4661,N_4286,N_3888);
nor U4662 (N_4662,N_3980,N_4342);
and U4663 (N_4663,N_3812,N_3931);
and U4664 (N_4664,N_3810,N_3999);
nand U4665 (N_4665,N_4276,N_3860);
nor U4666 (N_4666,N_4066,N_3871);
and U4667 (N_4667,N_4035,N_3988);
and U4668 (N_4668,N_4217,N_3779);
nor U4669 (N_4669,N_4295,N_3887);
or U4670 (N_4670,N_3935,N_3877);
nand U4671 (N_4671,N_4287,N_4195);
or U4672 (N_4672,N_3936,N_4242);
xor U4673 (N_4673,N_3933,N_3910);
and U4674 (N_4674,N_4028,N_4250);
nor U4675 (N_4675,N_3756,N_3855);
or U4676 (N_4676,N_3894,N_3836);
or U4677 (N_4677,N_3915,N_3847);
or U4678 (N_4678,N_4318,N_4037);
nand U4679 (N_4679,N_4371,N_4290);
nor U4680 (N_4680,N_4233,N_3852);
or U4681 (N_4681,N_4259,N_4269);
or U4682 (N_4682,N_3764,N_3854);
nand U4683 (N_4683,N_4281,N_4298);
nand U4684 (N_4684,N_4205,N_4193);
or U4685 (N_4685,N_4011,N_4149);
nand U4686 (N_4686,N_4079,N_4238);
or U4687 (N_4687,N_4128,N_3969);
nand U4688 (N_4688,N_3786,N_3873);
or U4689 (N_4689,N_3752,N_4010);
or U4690 (N_4690,N_4300,N_3769);
and U4691 (N_4691,N_3949,N_3859);
nand U4692 (N_4692,N_3962,N_4083);
nand U4693 (N_4693,N_4046,N_4079);
or U4694 (N_4694,N_4068,N_3852);
nor U4695 (N_4695,N_4036,N_3971);
and U4696 (N_4696,N_4044,N_4045);
nand U4697 (N_4697,N_4309,N_4121);
or U4698 (N_4698,N_4065,N_3785);
nor U4699 (N_4699,N_4011,N_4031);
or U4700 (N_4700,N_4341,N_4239);
or U4701 (N_4701,N_4034,N_3985);
nor U4702 (N_4702,N_3913,N_3899);
or U4703 (N_4703,N_3822,N_3997);
and U4704 (N_4704,N_4239,N_3774);
or U4705 (N_4705,N_3973,N_4153);
nor U4706 (N_4706,N_4169,N_3816);
or U4707 (N_4707,N_3769,N_3990);
nand U4708 (N_4708,N_4050,N_4072);
or U4709 (N_4709,N_3966,N_3819);
and U4710 (N_4710,N_3911,N_3906);
nand U4711 (N_4711,N_4236,N_3798);
or U4712 (N_4712,N_3852,N_3827);
and U4713 (N_4713,N_4059,N_4224);
and U4714 (N_4714,N_3928,N_3971);
and U4715 (N_4715,N_3917,N_4127);
nand U4716 (N_4716,N_3852,N_3843);
nor U4717 (N_4717,N_3912,N_4304);
nand U4718 (N_4718,N_4291,N_4202);
nand U4719 (N_4719,N_4237,N_3889);
nand U4720 (N_4720,N_3767,N_4197);
nand U4721 (N_4721,N_4093,N_4038);
or U4722 (N_4722,N_3919,N_4303);
and U4723 (N_4723,N_3917,N_3805);
nor U4724 (N_4724,N_4121,N_3955);
and U4725 (N_4725,N_4043,N_4353);
nand U4726 (N_4726,N_4296,N_4209);
or U4727 (N_4727,N_4217,N_4201);
or U4728 (N_4728,N_3757,N_4106);
nor U4729 (N_4729,N_4269,N_3926);
and U4730 (N_4730,N_3751,N_4093);
nand U4731 (N_4731,N_3812,N_4311);
xor U4732 (N_4732,N_4286,N_4254);
nor U4733 (N_4733,N_4229,N_3955);
xor U4734 (N_4734,N_4120,N_3854);
and U4735 (N_4735,N_3863,N_4253);
and U4736 (N_4736,N_4332,N_4170);
or U4737 (N_4737,N_4260,N_4272);
nor U4738 (N_4738,N_3847,N_3828);
nand U4739 (N_4739,N_3967,N_3776);
xnor U4740 (N_4740,N_4027,N_4255);
and U4741 (N_4741,N_4201,N_3986);
nor U4742 (N_4742,N_4152,N_3920);
xnor U4743 (N_4743,N_3872,N_4293);
xor U4744 (N_4744,N_3831,N_4096);
nand U4745 (N_4745,N_4111,N_4202);
nor U4746 (N_4746,N_3762,N_3845);
and U4747 (N_4747,N_3765,N_4161);
or U4748 (N_4748,N_3821,N_3861);
nor U4749 (N_4749,N_3798,N_3873);
xnor U4750 (N_4750,N_3980,N_4333);
nand U4751 (N_4751,N_4330,N_3918);
nand U4752 (N_4752,N_3758,N_4168);
or U4753 (N_4753,N_3893,N_4341);
nor U4754 (N_4754,N_4327,N_3819);
nor U4755 (N_4755,N_4233,N_4060);
and U4756 (N_4756,N_4108,N_3832);
or U4757 (N_4757,N_4269,N_4149);
or U4758 (N_4758,N_4062,N_4241);
nor U4759 (N_4759,N_4319,N_4249);
nand U4760 (N_4760,N_3939,N_4323);
or U4761 (N_4761,N_4348,N_4196);
nor U4762 (N_4762,N_3819,N_4197);
and U4763 (N_4763,N_4267,N_3770);
nor U4764 (N_4764,N_4319,N_3850);
and U4765 (N_4765,N_4329,N_3835);
xor U4766 (N_4766,N_4291,N_4061);
or U4767 (N_4767,N_3812,N_4144);
xnor U4768 (N_4768,N_3965,N_3923);
xor U4769 (N_4769,N_3860,N_4074);
nor U4770 (N_4770,N_3870,N_4066);
or U4771 (N_4771,N_3803,N_4254);
xnor U4772 (N_4772,N_4251,N_3799);
nor U4773 (N_4773,N_4026,N_4054);
nor U4774 (N_4774,N_4284,N_3886);
or U4775 (N_4775,N_3940,N_3819);
nand U4776 (N_4776,N_4175,N_4068);
nor U4777 (N_4777,N_3911,N_3796);
nand U4778 (N_4778,N_4329,N_3865);
nor U4779 (N_4779,N_4164,N_3798);
nor U4780 (N_4780,N_3892,N_3970);
and U4781 (N_4781,N_4297,N_4072);
nand U4782 (N_4782,N_4019,N_3979);
and U4783 (N_4783,N_4225,N_4031);
or U4784 (N_4784,N_4374,N_3948);
nand U4785 (N_4785,N_3873,N_4018);
xor U4786 (N_4786,N_4044,N_4145);
and U4787 (N_4787,N_3760,N_4138);
nand U4788 (N_4788,N_4241,N_3836);
nand U4789 (N_4789,N_3827,N_3805);
and U4790 (N_4790,N_4104,N_3946);
nand U4791 (N_4791,N_3956,N_3824);
nand U4792 (N_4792,N_3881,N_4126);
and U4793 (N_4793,N_4358,N_4280);
xnor U4794 (N_4794,N_4144,N_4200);
nor U4795 (N_4795,N_4186,N_4154);
nand U4796 (N_4796,N_3842,N_4349);
and U4797 (N_4797,N_4305,N_4361);
or U4798 (N_4798,N_3897,N_4324);
nor U4799 (N_4799,N_4340,N_4177);
and U4800 (N_4800,N_4306,N_4212);
and U4801 (N_4801,N_3949,N_4125);
or U4802 (N_4802,N_3962,N_4152);
xor U4803 (N_4803,N_4151,N_4159);
or U4804 (N_4804,N_4289,N_4351);
nand U4805 (N_4805,N_3975,N_3942);
xor U4806 (N_4806,N_3824,N_3931);
nand U4807 (N_4807,N_3836,N_3815);
xnor U4808 (N_4808,N_3918,N_4071);
nor U4809 (N_4809,N_4152,N_4044);
nand U4810 (N_4810,N_3963,N_4036);
nor U4811 (N_4811,N_3960,N_4046);
nor U4812 (N_4812,N_3945,N_3988);
nor U4813 (N_4813,N_4342,N_3852);
and U4814 (N_4814,N_4366,N_3997);
nor U4815 (N_4815,N_4361,N_3824);
nand U4816 (N_4816,N_3959,N_3763);
and U4817 (N_4817,N_4200,N_3825);
xor U4818 (N_4818,N_4111,N_3775);
nor U4819 (N_4819,N_4142,N_3829);
nand U4820 (N_4820,N_4058,N_3761);
xor U4821 (N_4821,N_4200,N_4125);
nand U4822 (N_4822,N_4356,N_4166);
nor U4823 (N_4823,N_3852,N_4112);
or U4824 (N_4824,N_4069,N_4027);
or U4825 (N_4825,N_3950,N_3770);
and U4826 (N_4826,N_4110,N_3883);
nand U4827 (N_4827,N_4066,N_3826);
or U4828 (N_4828,N_3944,N_3948);
or U4829 (N_4829,N_4233,N_4251);
or U4830 (N_4830,N_4136,N_3970);
and U4831 (N_4831,N_4193,N_3801);
nor U4832 (N_4832,N_3806,N_4255);
and U4833 (N_4833,N_3782,N_3799);
or U4834 (N_4834,N_4242,N_4285);
nor U4835 (N_4835,N_4132,N_4328);
nor U4836 (N_4836,N_4104,N_3760);
nand U4837 (N_4837,N_4275,N_4365);
nand U4838 (N_4838,N_4243,N_4030);
or U4839 (N_4839,N_4274,N_4210);
or U4840 (N_4840,N_4179,N_4229);
nor U4841 (N_4841,N_4146,N_3910);
or U4842 (N_4842,N_4093,N_3958);
nand U4843 (N_4843,N_4061,N_4247);
nand U4844 (N_4844,N_4041,N_3829);
or U4845 (N_4845,N_3911,N_4031);
or U4846 (N_4846,N_4166,N_4357);
and U4847 (N_4847,N_4141,N_3968);
nor U4848 (N_4848,N_3828,N_4055);
nor U4849 (N_4849,N_4176,N_4125);
nand U4850 (N_4850,N_4237,N_3816);
nor U4851 (N_4851,N_4209,N_3991);
nand U4852 (N_4852,N_4296,N_3806);
nand U4853 (N_4853,N_3982,N_3980);
xnor U4854 (N_4854,N_4371,N_4216);
and U4855 (N_4855,N_3977,N_3756);
or U4856 (N_4856,N_3865,N_4246);
or U4857 (N_4857,N_4294,N_4084);
and U4858 (N_4858,N_4036,N_4070);
or U4859 (N_4859,N_3767,N_3978);
or U4860 (N_4860,N_4272,N_3789);
nor U4861 (N_4861,N_4158,N_4015);
nand U4862 (N_4862,N_4266,N_4023);
or U4863 (N_4863,N_4035,N_4333);
and U4864 (N_4864,N_3866,N_3821);
or U4865 (N_4865,N_4158,N_4021);
nor U4866 (N_4866,N_4121,N_4174);
or U4867 (N_4867,N_3849,N_4061);
or U4868 (N_4868,N_3944,N_4131);
and U4869 (N_4869,N_4119,N_4207);
nand U4870 (N_4870,N_4148,N_3863);
and U4871 (N_4871,N_3930,N_3920);
nor U4872 (N_4872,N_4184,N_4246);
nor U4873 (N_4873,N_3959,N_4066);
and U4874 (N_4874,N_4173,N_3905);
and U4875 (N_4875,N_4364,N_3928);
nor U4876 (N_4876,N_4374,N_4134);
nand U4877 (N_4877,N_4361,N_4331);
nand U4878 (N_4878,N_4038,N_3954);
and U4879 (N_4879,N_3799,N_4211);
nor U4880 (N_4880,N_4280,N_4166);
nor U4881 (N_4881,N_4091,N_4329);
and U4882 (N_4882,N_4242,N_4192);
or U4883 (N_4883,N_3897,N_4167);
or U4884 (N_4884,N_3773,N_4228);
and U4885 (N_4885,N_4013,N_4167);
and U4886 (N_4886,N_4166,N_3942);
or U4887 (N_4887,N_4294,N_4311);
xnor U4888 (N_4888,N_3869,N_4075);
or U4889 (N_4889,N_4001,N_4324);
and U4890 (N_4890,N_3847,N_3950);
or U4891 (N_4891,N_4334,N_3780);
and U4892 (N_4892,N_4220,N_4369);
nand U4893 (N_4893,N_4371,N_3825);
nand U4894 (N_4894,N_4143,N_4336);
and U4895 (N_4895,N_4266,N_3815);
nor U4896 (N_4896,N_3763,N_4282);
or U4897 (N_4897,N_4212,N_4170);
or U4898 (N_4898,N_4341,N_3999);
nor U4899 (N_4899,N_3949,N_4076);
nor U4900 (N_4900,N_4366,N_4115);
nor U4901 (N_4901,N_3956,N_3871);
or U4902 (N_4902,N_4271,N_4355);
nand U4903 (N_4903,N_3917,N_3811);
and U4904 (N_4904,N_4339,N_4151);
or U4905 (N_4905,N_4199,N_3977);
and U4906 (N_4906,N_3992,N_4285);
nor U4907 (N_4907,N_3871,N_4277);
and U4908 (N_4908,N_3843,N_3990);
and U4909 (N_4909,N_4079,N_4235);
and U4910 (N_4910,N_4195,N_4266);
or U4911 (N_4911,N_4160,N_4303);
or U4912 (N_4912,N_3890,N_3874);
or U4913 (N_4913,N_4353,N_4321);
nor U4914 (N_4914,N_3839,N_4041);
and U4915 (N_4915,N_4341,N_4356);
nand U4916 (N_4916,N_3767,N_4102);
nor U4917 (N_4917,N_3909,N_4196);
nor U4918 (N_4918,N_3826,N_4364);
nor U4919 (N_4919,N_4085,N_4184);
or U4920 (N_4920,N_4075,N_3886);
nand U4921 (N_4921,N_4297,N_4341);
nor U4922 (N_4922,N_4260,N_4057);
or U4923 (N_4923,N_4109,N_3949);
nand U4924 (N_4924,N_3911,N_3952);
nor U4925 (N_4925,N_4184,N_3755);
or U4926 (N_4926,N_4268,N_3751);
or U4927 (N_4927,N_3974,N_4065);
nor U4928 (N_4928,N_3947,N_4359);
and U4929 (N_4929,N_4210,N_4308);
nor U4930 (N_4930,N_3866,N_4173);
xor U4931 (N_4931,N_3854,N_4132);
or U4932 (N_4932,N_4198,N_3957);
nor U4933 (N_4933,N_4343,N_4293);
or U4934 (N_4934,N_3868,N_4351);
nor U4935 (N_4935,N_3951,N_3763);
or U4936 (N_4936,N_4014,N_4253);
xor U4937 (N_4937,N_3830,N_3786);
nand U4938 (N_4938,N_3904,N_4122);
and U4939 (N_4939,N_3940,N_3793);
nand U4940 (N_4940,N_3795,N_3916);
xnor U4941 (N_4941,N_4200,N_4070);
or U4942 (N_4942,N_4134,N_4336);
nor U4943 (N_4943,N_3912,N_3842);
or U4944 (N_4944,N_4019,N_4243);
nor U4945 (N_4945,N_3795,N_3898);
and U4946 (N_4946,N_3785,N_4156);
xor U4947 (N_4947,N_4098,N_3791);
nor U4948 (N_4948,N_4345,N_4219);
xor U4949 (N_4949,N_3862,N_3924);
nand U4950 (N_4950,N_3902,N_3792);
and U4951 (N_4951,N_4185,N_3818);
nor U4952 (N_4952,N_4346,N_3865);
xnor U4953 (N_4953,N_4132,N_4312);
nor U4954 (N_4954,N_4058,N_3966);
nand U4955 (N_4955,N_3948,N_3819);
nand U4956 (N_4956,N_3865,N_4288);
nor U4957 (N_4957,N_4142,N_4202);
nor U4958 (N_4958,N_3766,N_3761);
nor U4959 (N_4959,N_4209,N_4317);
nor U4960 (N_4960,N_4308,N_4204);
and U4961 (N_4961,N_3916,N_4288);
or U4962 (N_4962,N_4351,N_4273);
or U4963 (N_4963,N_3782,N_4282);
nand U4964 (N_4964,N_3926,N_4069);
or U4965 (N_4965,N_4336,N_4051);
and U4966 (N_4966,N_3822,N_4225);
nand U4967 (N_4967,N_4307,N_4227);
or U4968 (N_4968,N_4099,N_3987);
nand U4969 (N_4969,N_4244,N_4342);
nand U4970 (N_4970,N_3779,N_4037);
nand U4971 (N_4971,N_3925,N_4112);
and U4972 (N_4972,N_3820,N_4167);
nand U4973 (N_4973,N_4370,N_4343);
nand U4974 (N_4974,N_3891,N_4144);
nor U4975 (N_4975,N_4372,N_4036);
nand U4976 (N_4976,N_4291,N_4015);
and U4977 (N_4977,N_4108,N_4052);
nor U4978 (N_4978,N_3763,N_3887);
or U4979 (N_4979,N_3932,N_4124);
nor U4980 (N_4980,N_4211,N_4013);
or U4981 (N_4981,N_4247,N_3975);
nor U4982 (N_4982,N_3878,N_3805);
nor U4983 (N_4983,N_4006,N_3759);
or U4984 (N_4984,N_3792,N_4151);
and U4985 (N_4985,N_4267,N_3792);
and U4986 (N_4986,N_3831,N_3779);
or U4987 (N_4987,N_4167,N_3901);
or U4988 (N_4988,N_3869,N_4132);
and U4989 (N_4989,N_4242,N_3858);
and U4990 (N_4990,N_4034,N_4299);
or U4991 (N_4991,N_4161,N_3966);
or U4992 (N_4992,N_4319,N_4077);
or U4993 (N_4993,N_4187,N_3885);
or U4994 (N_4994,N_4290,N_4313);
and U4995 (N_4995,N_4208,N_4236);
nor U4996 (N_4996,N_4372,N_3836);
nand U4997 (N_4997,N_3818,N_3949);
or U4998 (N_4998,N_3897,N_4245);
and U4999 (N_4999,N_3785,N_3951);
nand U5000 (N_5000,N_4717,N_4952);
or U5001 (N_5001,N_4713,N_4913);
and U5002 (N_5002,N_4848,N_4571);
and U5003 (N_5003,N_4435,N_4694);
and U5004 (N_5004,N_4586,N_4668);
nor U5005 (N_5005,N_4776,N_4474);
nor U5006 (N_5006,N_4595,N_4819);
nor U5007 (N_5007,N_4930,N_4481);
nor U5008 (N_5008,N_4487,N_4866);
nor U5009 (N_5009,N_4786,N_4378);
nand U5010 (N_5010,N_4746,N_4661);
nand U5011 (N_5011,N_4999,N_4592);
nor U5012 (N_5012,N_4415,N_4889);
and U5013 (N_5013,N_4546,N_4430);
and U5014 (N_5014,N_4590,N_4949);
and U5015 (N_5015,N_4589,N_4750);
nand U5016 (N_5016,N_4491,N_4985);
nor U5017 (N_5017,N_4795,N_4633);
or U5018 (N_5018,N_4961,N_4472);
nand U5019 (N_5019,N_4700,N_4376);
and U5020 (N_5020,N_4662,N_4901);
or U5021 (N_5021,N_4760,N_4802);
nand U5022 (N_5022,N_4607,N_4422);
nor U5023 (N_5023,N_4704,N_4890);
nor U5024 (N_5024,N_4835,N_4955);
nor U5025 (N_5025,N_4693,N_4622);
nor U5026 (N_5026,N_4723,N_4730);
nor U5027 (N_5027,N_4868,N_4648);
and U5028 (N_5028,N_4917,N_4807);
and U5029 (N_5029,N_4732,N_4426);
nor U5030 (N_5030,N_4878,N_4900);
nor U5031 (N_5031,N_4851,N_4941);
nand U5032 (N_5032,N_4519,N_4569);
nor U5033 (N_5033,N_4852,N_4530);
nand U5034 (N_5034,N_4888,N_4715);
and U5035 (N_5035,N_4790,N_4991);
nor U5036 (N_5036,N_4635,N_4950);
nand U5037 (N_5037,N_4480,N_4636);
and U5038 (N_5038,N_4869,N_4936);
or U5039 (N_5039,N_4860,N_4740);
xnor U5040 (N_5040,N_4755,N_4624);
nand U5041 (N_5041,N_4560,N_4849);
nor U5042 (N_5042,N_4965,N_4432);
xor U5043 (N_5043,N_4984,N_4401);
nor U5044 (N_5044,N_4391,N_4399);
and U5045 (N_5045,N_4864,N_4392);
nand U5046 (N_5046,N_4911,N_4412);
or U5047 (N_5047,N_4741,N_4854);
nand U5048 (N_5048,N_4921,N_4644);
nor U5049 (N_5049,N_4594,N_4669);
or U5050 (N_5050,N_4600,N_4800);
and U5051 (N_5051,N_4440,N_4791);
nor U5052 (N_5052,N_4642,N_4645);
nor U5053 (N_5053,N_4989,N_4827);
xor U5054 (N_5054,N_4583,N_4824);
nand U5055 (N_5055,N_4489,N_4983);
and U5056 (N_5056,N_4409,N_4541);
nor U5057 (N_5057,N_4681,N_4502);
nand U5058 (N_5058,N_4724,N_4982);
or U5059 (N_5059,N_4483,N_4626);
or U5060 (N_5060,N_4512,N_4783);
xor U5061 (N_5061,N_4988,N_4943);
or U5062 (N_5062,N_4695,N_4804);
nor U5063 (N_5063,N_4523,N_4809);
xor U5064 (N_5064,N_4551,N_4833);
nor U5065 (N_5065,N_4752,N_4815);
and U5066 (N_5066,N_4773,N_4553);
or U5067 (N_5067,N_4850,N_4380);
or U5068 (N_5068,N_4812,N_4844);
and U5069 (N_5069,N_4862,N_4924);
nor U5070 (N_5070,N_4920,N_4969);
and U5071 (N_5071,N_4896,N_4504);
or U5072 (N_5072,N_4979,N_4618);
nor U5073 (N_5073,N_4801,N_4431);
nor U5074 (N_5074,N_4674,N_4805);
xnor U5075 (N_5075,N_4613,N_4408);
nand U5076 (N_5076,N_4904,N_4582);
or U5077 (N_5077,N_4987,N_4863);
nand U5078 (N_5078,N_4505,N_4667);
nand U5079 (N_5079,N_4492,N_4992);
and U5080 (N_5080,N_4777,N_4775);
nand U5081 (N_5081,N_4436,N_4909);
nor U5082 (N_5082,N_4535,N_4459);
or U5083 (N_5083,N_4885,N_4526);
or U5084 (N_5084,N_4830,N_4528);
xnor U5085 (N_5085,N_4735,N_4689);
nor U5086 (N_5086,N_4679,N_4394);
nor U5087 (N_5087,N_4388,N_4811);
or U5088 (N_5088,N_4685,N_4767);
nand U5089 (N_5089,N_4453,N_4705);
nor U5090 (N_5090,N_4711,N_4963);
nor U5091 (N_5091,N_4437,N_4718);
xor U5092 (N_5092,N_4840,N_4722);
or U5093 (N_5093,N_4923,N_4657);
or U5094 (N_5094,N_4927,N_4813);
nor U5095 (N_5095,N_4397,N_4585);
nand U5096 (N_5096,N_4736,N_4641);
nand U5097 (N_5097,N_4816,N_4877);
nand U5098 (N_5098,N_4671,N_4602);
nor U5099 (N_5099,N_4699,N_4446);
nor U5100 (N_5100,N_4400,N_4785);
or U5101 (N_5101,N_4879,N_4688);
xnor U5102 (N_5102,N_4486,N_4566);
or U5103 (N_5103,N_4696,N_4509);
or U5104 (N_5104,N_4751,N_4886);
nand U5105 (N_5105,N_4534,N_4993);
nand U5106 (N_5106,N_4788,N_4654);
or U5107 (N_5107,N_4419,N_4429);
nor U5108 (N_5108,N_4899,N_4832);
nor U5109 (N_5109,N_4609,N_4898);
nor U5110 (N_5110,N_4908,N_4957);
and U5111 (N_5111,N_4568,N_4540);
nor U5112 (N_5112,N_4496,N_4384);
and U5113 (N_5113,N_4729,N_4847);
or U5114 (N_5114,N_4880,N_4698);
nand U5115 (N_5115,N_4421,N_4604);
or U5116 (N_5116,N_4576,N_4464);
xor U5117 (N_5117,N_4906,N_4787);
or U5118 (N_5118,N_4856,N_4570);
or U5119 (N_5119,N_4411,N_4445);
or U5120 (N_5120,N_4458,N_4960);
or U5121 (N_5121,N_4475,N_4720);
nand U5122 (N_5122,N_4587,N_4895);
nor U5123 (N_5123,N_4710,N_4647);
nor U5124 (N_5124,N_4441,N_4998);
nand U5125 (N_5125,N_4452,N_4652);
nor U5126 (N_5126,N_4454,N_4680);
or U5127 (N_5127,N_4617,N_4769);
and U5128 (N_5128,N_4874,N_4975);
or U5129 (N_5129,N_4511,N_4867);
or U5130 (N_5130,N_4948,N_4402);
or U5131 (N_5131,N_4842,N_4544);
and U5132 (N_5132,N_4754,N_4702);
or U5133 (N_5133,N_4499,N_4770);
nand U5134 (N_5134,N_4784,N_4545);
xnor U5135 (N_5135,N_4381,N_4758);
nand U5136 (N_5136,N_4498,N_4527);
xnor U5137 (N_5137,N_4905,N_4947);
nor U5138 (N_5138,N_4858,N_4573);
nor U5139 (N_5139,N_4966,N_4559);
and U5140 (N_5140,N_4806,N_4581);
nand U5141 (N_5141,N_4942,N_4606);
nand U5142 (N_5142,N_4390,N_4956);
and U5143 (N_5143,N_4731,N_4470);
nor U5144 (N_5144,N_4638,N_4780);
nor U5145 (N_5145,N_4759,N_4514);
nand U5146 (N_5146,N_4771,N_4692);
and U5147 (N_5147,N_4630,N_4574);
nand U5148 (N_5148,N_4931,N_4513);
nor U5149 (N_5149,N_4403,N_4970);
or U5150 (N_5150,N_4643,N_4876);
or U5151 (N_5151,N_4621,N_4684);
xnor U5152 (N_5152,N_4423,N_4404);
and U5153 (N_5153,N_4873,N_4855);
or U5154 (N_5154,N_4623,N_4593);
and U5155 (N_5155,N_4597,N_4424);
nand U5156 (N_5156,N_4477,N_4524);
and U5157 (N_5157,N_4719,N_4831);
or U5158 (N_5158,N_4548,N_4996);
nor U5159 (N_5159,N_4610,N_4588);
or U5160 (N_5160,N_4549,N_4825);
nand U5161 (N_5161,N_4980,N_4990);
and U5162 (N_5162,N_4427,N_4425);
nor U5163 (N_5163,N_4637,N_4789);
or U5164 (N_5164,N_4656,N_4745);
or U5165 (N_5165,N_4479,N_4646);
and U5166 (N_5166,N_4473,N_4940);
and U5167 (N_5167,N_4557,N_4605);
and U5168 (N_5168,N_4884,N_4768);
nand U5169 (N_5169,N_4914,N_4572);
nand U5170 (N_5170,N_4976,N_4389);
or U5171 (N_5171,N_4902,N_4525);
nor U5172 (N_5172,N_4547,N_4981);
nand U5173 (N_5173,N_4838,N_4728);
nand U5174 (N_5174,N_4725,N_4537);
nor U5175 (N_5175,N_4515,N_4666);
nor U5176 (N_5176,N_4821,N_4640);
nand U5177 (N_5177,N_4714,N_4978);
nand U5178 (N_5178,N_4968,N_4678);
or U5179 (N_5179,N_4781,N_4385);
nor U5180 (N_5180,N_4916,N_4872);
nor U5181 (N_5181,N_4716,N_4834);
or U5182 (N_5182,N_4531,N_4443);
and U5183 (N_5183,N_4686,N_4887);
xor U5184 (N_5184,N_4794,N_4659);
nor U5185 (N_5185,N_4861,N_4562);
and U5186 (N_5186,N_4461,N_4665);
and U5187 (N_5187,N_4550,N_4871);
nor U5188 (N_5188,N_4683,N_4539);
nand U5189 (N_5189,N_4973,N_4447);
nor U5190 (N_5190,N_4747,N_4500);
nand U5191 (N_5191,N_4967,N_4912);
or U5192 (N_5192,N_4817,N_4929);
nor U5193 (N_5193,N_4706,N_4469);
nand U5194 (N_5194,N_4954,N_4383);
nor U5195 (N_5195,N_4934,N_4619);
xor U5196 (N_5196,N_4631,N_4455);
and U5197 (N_5197,N_4691,N_4893);
or U5198 (N_5198,N_4762,N_4598);
or U5199 (N_5199,N_4709,N_4485);
or U5200 (N_5200,N_4939,N_4456);
nor U5201 (N_5201,N_4612,N_4945);
and U5202 (N_5202,N_4467,N_4922);
or U5203 (N_5203,N_4687,N_4563);
nand U5204 (N_5204,N_4761,N_4529);
nor U5205 (N_5205,N_4958,N_4375);
and U5206 (N_5206,N_4558,N_4386);
nor U5207 (N_5207,N_4907,N_4655);
nand U5208 (N_5208,N_4629,N_4843);
and U5209 (N_5209,N_4416,N_4915);
and U5210 (N_5210,N_4584,N_4828);
nand U5211 (N_5211,N_4442,N_4933);
xor U5212 (N_5212,N_4733,N_4853);
nand U5213 (N_5213,N_4796,N_4903);
nor U5214 (N_5214,N_4532,N_4875);
or U5215 (N_5215,N_4554,N_4379);
xnor U5216 (N_5216,N_4742,N_4756);
nor U5217 (N_5217,N_4995,N_4937);
nand U5218 (N_5218,N_4542,N_4490);
and U5219 (N_5219,N_4977,N_4507);
nor U5220 (N_5220,N_4508,N_4651);
and U5221 (N_5221,N_4739,N_4677);
nor U5222 (N_5222,N_4596,N_4676);
or U5223 (N_5223,N_4797,N_4766);
or U5224 (N_5224,N_4611,N_4919);
and U5225 (N_5225,N_4748,N_4701);
xnor U5226 (N_5226,N_4712,N_4463);
nor U5227 (N_5227,N_4845,N_4497);
or U5228 (N_5228,N_4660,N_4634);
or U5229 (N_5229,N_4520,N_4407);
and U5230 (N_5230,N_4841,N_4543);
or U5231 (N_5231,N_4798,N_4932);
nor U5232 (N_5232,N_4410,N_4418);
nor U5233 (N_5233,N_4959,N_4823);
nor U5234 (N_5234,N_4870,N_4764);
nor U5235 (N_5235,N_4744,N_4727);
nor U5236 (N_5236,N_4910,N_4925);
nor U5237 (N_5237,N_4387,N_4536);
nand U5238 (N_5238,N_4580,N_4449);
nor U5239 (N_5239,N_4820,N_4836);
or U5240 (N_5240,N_4433,N_4413);
and U5241 (N_5241,N_4894,N_4632);
nand U5242 (N_5242,N_4482,N_4757);
or U5243 (N_5243,N_4438,N_4672);
xor U5244 (N_5244,N_4457,N_4974);
nand U5245 (N_5245,N_4420,N_4721);
nand U5246 (N_5246,N_4518,N_4774);
or U5247 (N_5247,N_4649,N_4938);
and U5248 (N_5248,N_4556,N_4564);
and U5249 (N_5249,N_4603,N_4708);
or U5250 (N_5250,N_4510,N_4478);
and U5251 (N_5251,N_4944,N_4753);
or U5252 (N_5252,N_4664,N_4964);
and U5253 (N_5253,N_4778,N_4434);
xnor U5254 (N_5254,N_4468,N_4926);
nor U5255 (N_5255,N_4465,N_4928);
nand U5256 (N_5256,N_4743,N_4591);
and U5257 (N_5257,N_4451,N_4448);
or U5258 (N_5258,N_4897,N_4865);
nor U5259 (N_5259,N_4707,N_4690);
xnor U5260 (N_5260,N_4428,N_4803);
and U5261 (N_5261,N_4565,N_4555);
and U5262 (N_5262,N_4673,N_4857);
or U5263 (N_5263,N_4738,N_4663);
and U5264 (N_5264,N_4882,N_4488);
nand U5265 (N_5265,N_4578,N_4810);
nand U5266 (N_5266,N_4883,N_4814);
or U5267 (N_5267,N_4881,N_4406);
or U5268 (N_5268,N_4396,N_4749);
or U5269 (N_5269,N_4972,N_4615);
or U5270 (N_5270,N_4675,N_4951);
nand U5271 (N_5271,N_4414,N_4627);
and U5272 (N_5272,N_4986,N_4994);
nor U5273 (N_5273,N_4501,N_4765);
and U5274 (N_5274,N_4620,N_4601);
and U5275 (N_5275,N_4639,N_4953);
xor U5276 (N_5276,N_4503,N_4650);
and U5277 (N_5277,N_4826,N_4599);
or U5278 (N_5278,N_4628,N_4891);
and U5279 (N_5279,N_4493,N_4444);
or U5280 (N_5280,N_4625,N_4484);
or U5281 (N_5281,N_4918,N_4538);
or U5282 (N_5282,N_4439,N_4552);
or U5283 (N_5283,N_4417,N_4799);
nor U5284 (N_5284,N_4614,N_4521);
and U5285 (N_5285,N_4567,N_4460);
nor U5286 (N_5286,N_4772,N_4782);
and U5287 (N_5287,N_4808,N_4494);
or U5288 (N_5288,N_4495,N_4462);
nor U5289 (N_5289,N_4395,N_4726);
xor U5290 (N_5290,N_4971,N_4377);
or U5291 (N_5291,N_4393,N_4839);
and U5292 (N_5292,N_4608,N_4575);
or U5293 (N_5293,N_4405,N_4829);
xnor U5294 (N_5294,N_4779,N_4793);
nor U5295 (N_5295,N_4892,N_4703);
and U5296 (N_5296,N_4476,N_4737);
xnor U5297 (N_5297,N_4653,N_4763);
and U5298 (N_5298,N_4506,N_4533);
nand U5299 (N_5299,N_4734,N_4579);
and U5300 (N_5300,N_4658,N_4818);
nand U5301 (N_5301,N_4670,N_4577);
nand U5302 (N_5302,N_4962,N_4517);
nor U5303 (N_5303,N_4682,N_4616);
nor U5304 (N_5304,N_4792,N_4561);
and U5305 (N_5305,N_4471,N_4382);
xnor U5306 (N_5306,N_4837,N_4946);
nor U5307 (N_5307,N_4466,N_4859);
nand U5308 (N_5308,N_4450,N_4822);
nor U5309 (N_5309,N_4398,N_4516);
nor U5310 (N_5310,N_4935,N_4997);
nand U5311 (N_5311,N_4522,N_4846);
or U5312 (N_5312,N_4697,N_4669);
xnor U5313 (N_5313,N_4584,N_4618);
xnor U5314 (N_5314,N_4896,N_4590);
or U5315 (N_5315,N_4600,N_4968);
nor U5316 (N_5316,N_4925,N_4703);
nor U5317 (N_5317,N_4754,N_4957);
nand U5318 (N_5318,N_4949,N_4599);
and U5319 (N_5319,N_4962,N_4822);
nor U5320 (N_5320,N_4650,N_4427);
and U5321 (N_5321,N_4823,N_4776);
nand U5322 (N_5322,N_4891,N_4929);
nor U5323 (N_5323,N_4524,N_4433);
and U5324 (N_5324,N_4490,N_4992);
and U5325 (N_5325,N_4402,N_4565);
nand U5326 (N_5326,N_4680,N_4912);
nand U5327 (N_5327,N_4714,N_4853);
nand U5328 (N_5328,N_4549,N_4397);
and U5329 (N_5329,N_4501,N_4520);
and U5330 (N_5330,N_4976,N_4774);
and U5331 (N_5331,N_4448,N_4584);
nand U5332 (N_5332,N_4655,N_4778);
or U5333 (N_5333,N_4962,N_4873);
or U5334 (N_5334,N_4508,N_4412);
and U5335 (N_5335,N_4795,N_4648);
or U5336 (N_5336,N_4965,N_4420);
nand U5337 (N_5337,N_4793,N_4796);
and U5338 (N_5338,N_4471,N_4625);
or U5339 (N_5339,N_4781,N_4839);
or U5340 (N_5340,N_4516,N_4409);
xor U5341 (N_5341,N_4786,N_4878);
and U5342 (N_5342,N_4682,N_4381);
nor U5343 (N_5343,N_4423,N_4681);
and U5344 (N_5344,N_4470,N_4656);
xnor U5345 (N_5345,N_4628,N_4390);
or U5346 (N_5346,N_4969,N_4818);
and U5347 (N_5347,N_4375,N_4528);
nor U5348 (N_5348,N_4505,N_4561);
nand U5349 (N_5349,N_4861,N_4416);
and U5350 (N_5350,N_4776,N_4970);
or U5351 (N_5351,N_4716,N_4546);
and U5352 (N_5352,N_4676,N_4506);
and U5353 (N_5353,N_4639,N_4618);
nor U5354 (N_5354,N_4567,N_4830);
or U5355 (N_5355,N_4786,N_4915);
nand U5356 (N_5356,N_4703,N_4469);
nor U5357 (N_5357,N_4444,N_4384);
or U5358 (N_5358,N_4920,N_4696);
or U5359 (N_5359,N_4771,N_4554);
or U5360 (N_5360,N_4557,N_4865);
nor U5361 (N_5361,N_4968,N_4931);
and U5362 (N_5362,N_4870,N_4844);
xor U5363 (N_5363,N_4751,N_4581);
nand U5364 (N_5364,N_4867,N_4497);
or U5365 (N_5365,N_4550,N_4606);
or U5366 (N_5366,N_4835,N_4557);
nor U5367 (N_5367,N_4855,N_4417);
or U5368 (N_5368,N_4425,N_4693);
or U5369 (N_5369,N_4578,N_4447);
and U5370 (N_5370,N_4861,N_4654);
nor U5371 (N_5371,N_4751,N_4950);
xnor U5372 (N_5372,N_4919,N_4447);
nand U5373 (N_5373,N_4571,N_4376);
xor U5374 (N_5374,N_4727,N_4436);
nor U5375 (N_5375,N_4595,N_4778);
and U5376 (N_5376,N_4721,N_4685);
nand U5377 (N_5377,N_4469,N_4547);
or U5378 (N_5378,N_4772,N_4860);
and U5379 (N_5379,N_4930,N_4468);
and U5380 (N_5380,N_4784,N_4993);
nor U5381 (N_5381,N_4657,N_4993);
nor U5382 (N_5382,N_4992,N_4999);
nor U5383 (N_5383,N_4381,N_4771);
nor U5384 (N_5384,N_4541,N_4943);
nor U5385 (N_5385,N_4725,N_4496);
nand U5386 (N_5386,N_4665,N_4704);
nand U5387 (N_5387,N_4830,N_4887);
or U5388 (N_5388,N_4777,N_4801);
nor U5389 (N_5389,N_4610,N_4431);
nand U5390 (N_5390,N_4685,N_4939);
nor U5391 (N_5391,N_4565,N_4786);
and U5392 (N_5392,N_4688,N_4953);
or U5393 (N_5393,N_4691,N_4953);
nand U5394 (N_5394,N_4642,N_4585);
or U5395 (N_5395,N_4376,N_4908);
xnor U5396 (N_5396,N_4961,N_4992);
nor U5397 (N_5397,N_4599,N_4501);
nor U5398 (N_5398,N_4568,N_4613);
nor U5399 (N_5399,N_4912,N_4738);
or U5400 (N_5400,N_4565,N_4806);
and U5401 (N_5401,N_4532,N_4504);
nor U5402 (N_5402,N_4687,N_4747);
nor U5403 (N_5403,N_4669,N_4929);
and U5404 (N_5404,N_4703,N_4383);
nand U5405 (N_5405,N_4949,N_4934);
nor U5406 (N_5406,N_4664,N_4987);
and U5407 (N_5407,N_4996,N_4874);
nor U5408 (N_5408,N_4396,N_4712);
nand U5409 (N_5409,N_4557,N_4979);
nand U5410 (N_5410,N_4787,N_4811);
nand U5411 (N_5411,N_4981,N_4785);
and U5412 (N_5412,N_4834,N_4393);
nand U5413 (N_5413,N_4753,N_4477);
nor U5414 (N_5414,N_4506,N_4974);
or U5415 (N_5415,N_4598,N_4574);
and U5416 (N_5416,N_4847,N_4565);
nand U5417 (N_5417,N_4815,N_4821);
or U5418 (N_5418,N_4539,N_4859);
nor U5419 (N_5419,N_4620,N_4459);
nor U5420 (N_5420,N_4419,N_4388);
nor U5421 (N_5421,N_4739,N_4755);
or U5422 (N_5422,N_4906,N_4924);
nand U5423 (N_5423,N_4548,N_4584);
or U5424 (N_5424,N_4785,N_4740);
xor U5425 (N_5425,N_4703,N_4965);
or U5426 (N_5426,N_4859,N_4732);
nor U5427 (N_5427,N_4854,N_4944);
or U5428 (N_5428,N_4661,N_4815);
or U5429 (N_5429,N_4805,N_4816);
nand U5430 (N_5430,N_4410,N_4938);
and U5431 (N_5431,N_4778,N_4846);
xor U5432 (N_5432,N_4411,N_4498);
or U5433 (N_5433,N_4978,N_4726);
nand U5434 (N_5434,N_4824,N_4480);
xnor U5435 (N_5435,N_4954,N_4544);
xnor U5436 (N_5436,N_4751,N_4511);
or U5437 (N_5437,N_4493,N_4661);
or U5438 (N_5438,N_4884,N_4626);
nor U5439 (N_5439,N_4996,N_4650);
nand U5440 (N_5440,N_4758,N_4679);
xor U5441 (N_5441,N_4986,N_4444);
nand U5442 (N_5442,N_4548,N_4636);
and U5443 (N_5443,N_4792,N_4848);
and U5444 (N_5444,N_4641,N_4981);
or U5445 (N_5445,N_4472,N_4434);
nand U5446 (N_5446,N_4823,N_4714);
nor U5447 (N_5447,N_4409,N_4964);
and U5448 (N_5448,N_4955,N_4919);
or U5449 (N_5449,N_4724,N_4605);
nor U5450 (N_5450,N_4674,N_4566);
and U5451 (N_5451,N_4858,N_4574);
nand U5452 (N_5452,N_4621,N_4696);
nor U5453 (N_5453,N_4854,N_4464);
nand U5454 (N_5454,N_4894,N_4926);
nor U5455 (N_5455,N_4419,N_4465);
nand U5456 (N_5456,N_4865,N_4547);
and U5457 (N_5457,N_4470,N_4527);
or U5458 (N_5458,N_4851,N_4685);
and U5459 (N_5459,N_4796,N_4471);
and U5460 (N_5460,N_4899,N_4788);
nor U5461 (N_5461,N_4816,N_4699);
nor U5462 (N_5462,N_4823,N_4547);
nand U5463 (N_5463,N_4858,N_4802);
nor U5464 (N_5464,N_4560,N_4703);
and U5465 (N_5465,N_4528,N_4983);
nand U5466 (N_5466,N_4548,N_4797);
nor U5467 (N_5467,N_4739,N_4806);
and U5468 (N_5468,N_4686,N_4479);
nor U5469 (N_5469,N_4396,N_4629);
or U5470 (N_5470,N_4660,N_4587);
nand U5471 (N_5471,N_4801,N_4659);
and U5472 (N_5472,N_4580,N_4463);
nor U5473 (N_5473,N_4912,N_4944);
or U5474 (N_5474,N_4862,N_4981);
or U5475 (N_5475,N_4932,N_4966);
nand U5476 (N_5476,N_4459,N_4780);
or U5477 (N_5477,N_4930,N_4994);
and U5478 (N_5478,N_4923,N_4691);
nor U5479 (N_5479,N_4679,N_4545);
and U5480 (N_5480,N_4419,N_4949);
or U5481 (N_5481,N_4438,N_4656);
xor U5482 (N_5482,N_4398,N_4601);
and U5483 (N_5483,N_4831,N_4788);
or U5484 (N_5484,N_4380,N_4829);
and U5485 (N_5485,N_4922,N_4481);
nor U5486 (N_5486,N_4667,N_4579);
and U5487 (N_5487,N_4811,N_4800);
nand U5488 (N_5488,N_4375,N_4959);
or U5489 (N_5489,N_4521,N_4555);
or U5490 (N_5490,N_4966,N_4549);
nor U5491 (N_5491,N_4835,N_4617);
or U5492 (N_5492,N_4753,N_4796);
nand U5493 (N_5493,N_4755,N_4809);
nand U5494 (N_5494,N_4815,N_4487);
nand U5495 (N_5495,N_4562,N_4620);
nand U5496 (N_5496,N_4607,N_4527);
nand U5497 (N_5497,N_4440,N_4971);
and U5498 (N_5498,N_4706,N_4440);
or U5499 (N_5499,N_4772,N_4600);
and U5500 (N_5500,N_4732,N_4972);
nor U5501 (N_5501,N_4383,N_4650);
and U5502 (N_5502,N_4376,N_4893);
xnor U5503 (N_5503,N_4819,N_4827);
nor U5504 (N_5504,N_4755,N_4614);
and U5505 (N_5505,N_4934,N_4798);
nand U5506 (N_5506,N_4697,N_4505);
or U5507 (N_5507,N_4474,N_4997);
nor U5508 (N_5508,N_4973,N_4682);
or U5509 (N_5509,N_4619,N_4942);
nand U5510 (N_5510,N_4787,N_4702);
nor U5511 (N_5511,N_4898,N_4974);
xor U5512 (N_5512,N_4668,N_4637);
and U5513 (N_5513,N_4457,N_4631);
nand U5514 (N_5514,N_4823,N_4426);
or U5515 (N_5515,N_4968,N_4506);
nand U5516 (N_5516,N_4727,N_4665);
and U5517 (N_5517,N_4856,N_4499);
nand U5518 (N_5518,N_4886,N_4889);
nand U5519 (N_5519,N_4864,N_4394);
and U5520 (N_5520,N_4492,N_4859);
and U5521 (N_5521,N_4495,N_4676);
nor U5522 (N_5522,N_4633,N_4575);
nand U5523 (N_5523,N_4545,N_4682);
xor U5524 (N_5524,N_4478,N_4412);
or U5525 (N_5525,N_4628,N_4421);
nand U5526 (N_5526,N_4767,N_4807);
xor U5527 (N_5527,N_4899,N_4848);
nor U5528 (N_5528,N_4880,N_4583);
and U5529 (N_5529,N_4754,N_4634);
xnor U5530 (N_5530,N_4566,N_4773);
nand U5531 (N_5531,N_4508,N_4940);
nand U5532 (N_5532,N_4652,N_4968);
nor U5533 (N_5533,N_4559,N_4907);
nor U5534 (N_5534,N_4690,N_4502);
nand U5535 (N_5535,N_4483,N_4878);
or U5536 (N_5536,N_4463,N_4902);
and U5537 (N_5537,N_4561,N_4875);
xor U5538 (N_5538,N_4550,N_4992);
nand U5539 (N_5539,N_4699,N_4390);
or U5540 (N_5540,N_4730,N_4918);
nor U5541 (N_5541,N_4556,N_4691);
or U5542 (N_5542,N_4885,N_4812);
nand U5543 (N_5543,N_4442,N_4505);
nor U5544 (N_5544,N_4600,N_4557);
or U5545 (N_5545,N_4978,N_4815);
or U5546 (N_5546,N_4398,N_4747);
and U5547 (N_5547,N_4396,N_4943);
nor U5548 (N_5548,N_4535,N_4745);
nor U5549 (N_5549,N_4747,N_4998);
nor U5550 (N_5550,N_4945,N_4499);
nand U5551 (N_5551,N_4840,N_4588);
nand U5552 (N_5552,N_4787,N_4583);
nor U5553 (N_5553,N_4392,N_4420);
nor U5554 (N_5554,N_4642,N_4617);
nor U5555 (N_5555,N_4786,N_4837);
nand U5556 (N_5556,N_4924,N_4389);
and U5557 (N_5557,N_4633,N_4643);
nand U5558 (N_5558,N_4713,N_4585);
nand U5559 (N_5559,N_4484,N_4712);
nand U5560 (N_5560,N_4904,N_4823);
or U5561 (N_5561,N_4721,N_4782);
nor U5562 (N_5562,N_4567,N_4668);
nor U5563 (N_5563,N_4660,N_4433);
and U5564 (N_5564,N_4759,N_4492);
and U5565 (N_5565,N_4655,N_4723);
or U5566 (N_5566,N_4837,N_4677);
nand U5567 (N_5567,N_4840,N_4563);
xor U5568 (N_5568,N_4850,N_4471);
nand U5569 (N_5569,N_4532,N_4460);
or U5570 (N_5570,N_4934,N_4379);
xor U5571 (N_5571,N_4968,N_4829);
nor U5572 (N_5572,N_4386,N_4816);
or U5573 (N_5573,N_4749,N_4847);
nor U5574 (N_5574,N_4400,N_4613);
and U5575 (N_5575,N_4759,N_4508);
and U5576 (N_5576,N_4490,N_4963);
xor U5577 (N_5577,N_4849,N_4750);
nand U5578 (N_5578,N_4879,N_4746);
nor U5579 (N_5579,N_4523,N_4697);
nor U5580 (N_5580,N_4920,N_4933);
nor U5581 (N_5581,N_4667,N_4586);
or U5582 (N_5582,N_4875,N_4956);
or U5583 (N_5583,N_4765,N_4874);
and U5584 (N_5584,N_4890,N_4377);
and U5585 (N_5585,N_4496,N_4939);
nor U5586 (N_5586,N_4639,N_4390);
and U5587 (N_5587,N_4815,N_4692);
xnor U5588 (N_5588,N_4796,N_4880);
or U5589 (N_5589,N_4974,N_4692);
and U5590 (N_5590,N_4395,N_4906);
or U5591 (N_5591,N_4487,N_4466);
and U5592 (N_5592,N_4849,N_4789);
nand U5593 (N_5593,N_4825,N_4470);
nor U5594 (N_5594,N_4751,N_4599);
nand U5595 (N_5595,N_4883,N_4989);
and U5596 (N_5596,N_4635,N_4581);
and U5597 (N_5597,N_4642,N_4513);
nor U5598 (N_5598,N_4868,N_4791);
and U5599 (N_5599,N_4621,N_4813);
nor U5600 (N_5600,N_4520,N_4720);
and U5601 (N_5601,N_4639,N_4920);
or U5602 (N_5602,N_4697,N_4813);
nand U5603 (N_5603,N_4569,N_4586);
nand U5604 (N_5604,N_4980,N_4692);
or U5605 (N_5605,N_4763,N_4975);
nand U5606 (N_5606,N_4969,N_4975);
nor U5607 (N_5607,N_4630,N_4797);
or U5608 (N_5608,N_4569,N_4724);
nor U5609 (N_5609,N_4818,N_4636);
or U5610 (N_5610,N_4660,N_4771);
nor U5611 (N_5611,N_4689,N_4526);
and U5612 (N_5612,N_4655,N_4453);
or U5613 (N_5613,N_4500,N_4741);
and U5614 (N_5614,N_4967,N_4406);
xor U5615 (N_5615,N_4556,N_4393);
nor U5616 (N_5616,N_4773,N_4823);
and U5617 (N_5617,N_4622,N_4376);
nand U5618 (N_5618,N_4888,N_4781);
or U5619 (N_5619,N_4555,N_4473);
nor U5620 (N_5620,N_4978,N_4736);
or U5621 (N_5621,N_4991,N_4570);
or U5622 (N_5622,N_4643,N_4420);
nor U5623 (N_5623,N_4495,N_4881);
nand U5624 (N_5624,N_4978,N_4588);
nand U5625 (N_5625,N_5441,N_5267);
nor U5626 (N_5626,N_5133,N_5611);
nand U5627 (N_5627,N_5180,N_5140);
and U5628 (N_5628,N_5597,N_5598);
nor U5629 (N_5629,N_5258,N_5376);
nand U5630 (N_5630,N_5016,N_5237);
or U5631 (N_5631,N_5322,N_5354);
and U5632 (N_5632,N_5141,N_5038);
nand U5633 (N_5633,N_5327,N_5533);
and U5634 (N_5634,N_5348,N_5394);
nand U5635 (N_5635,N_5340,N_5112);
and U5636 (N_5636,N_5577,N_5343);
xor U5637 (N_5637,N_5036,N_5539);
and U5638 (N_5638,N_5251,N_5253);
nand U5639 (N_5639,N_5266,N_5483);
nand U5640 (N_5640,N_5099,N_5560);
nand U5641 (N_5641,N_5186,N_5513);
and U5642 (N_5642,N_5072,N_5586);
xor U5643 (N_5643,N_5044,N_5238);
nor U5644 (N_5644,N_5110,N_5457);
or U5645 (N_5645,N_5402,N_5025);
and U5646 (N_5646,N_5175,N_5462);
nand U5647 (N_5647,N_5042,N_5329);
or U5648 (N_5648,N_5285,N_5056);
nand U5649 (N_5649,N_5459,N_5417);
nand U5650 (N_5650,N_5595,N_5135);
or U5651 (N_5651,N_5078,N_5603);
or U5652 (N_5652,N_5245,N_5410);
nor U5653 (N_5653,N_5588,N_5308);
xor U5654 (N_5654,N_5614,N_5107);
nand U5655 (N_5655,N_5204,N_5510);
nor U5656 (N_5656,N_5451,N_5464);
xnor U5657 (N_5657,N_5511,N_5275);
xor U5658 (N_5658,N_5054,N_5557);
nand U5659 (N_5659,N_5368,N_5012);
or U5660 (N_5660,N_5249,N_5129);
and U5661 (N_5661,N_5288,N_5125);
and U5662 (N_5662,N_5567,N_5356);
nand U5663 (N_5663,N_5490,N_5066);
nor U5664 (N_5664,N_5010,N_5550);
nor U5665 (N_5665,N_5532,N_5353);
and U5666 (N_5666,N_5516,N_5091);
or U5667 (N_5667,N_5440,N_5254);
or U5668 (N_5668,N_5471,N_5137);
or U5669 (N_5669,N_5362,N_5435);
nand U5670 (N_5670,N_5583,N_5017);
or U5671 (N_5671,N_5081,N_5324);
nand U5672 (N_5672,N_5339,N_5478);
or U5673 (N_5673,N_5261,N_5423);
and U5674 (N_5674,N_5127,N_5194);
nand U5675 (N_5675,N_5525,N_5024);
and U5676 (N_5676,N_5517,N_5108);
nor U5677 (N_5677,N_5281,N_5386);
nand U5678 (N_5678,N_5475,N_5156);
xor U5679 (N_5679,N_5096,N_5172);
nand U5680 (N_5680,N_5079,N_5013);
nand U5681 (N_5681,N_5334,N_5346);
nand U5682 (N_5682,N_5551,N_5111);
or U5683 (N_5683,N_5458,N_5278);
and U5684 (N_5684,N_5549,N_5591);
or U5685 (N_5685,N_5450,N_5231);
or U5686 (N_5686,N_5241,N_5542);
and U5687 (N_5687,N_5120,N_5564);
or U5688 (N_5688,N_5100,N_5105);
nand U5689 (N_5689,N_5074,N_5320);
and U5690 (N_5690,N_5561,N_5065);
nor U5691 (N_5691,N_5401,N_5495);
nor U5692 (N_5692,N_5094,N_5239);
or U5693 (N_5693,N_5021,N_5090);
and U5694 (N_5694,N_5286,N_5150);
and U5695 (N_5695,N_5480,N_5287);
and U5696 (N_5696,N_5470,N_5338);
nor U5697 (N_5697,N_5585,N_5520);
nor U5698 (N_5698,N_5443,N_5500);
nor U5699 (N_5699,N_5344,N_5210);
or U5700 (N_5700,N_5311,N_5041);
or U5701 (N_5701,N_5143,N_5230);
or U5702 (N_5702,N_5104,N_5089);
or U5703 (N_5703,N_5055,N_5144);
xor U5704 (N_5704,N_5412,N_5566);
xnor U5705 (N_5705,N_5122,N_5448);
nor U5706 (N_5706,N_5255,N_5164);
and U5707 (N_5707,N_5121,N_5103);
nand U5708 (N_5708,N_5463,N_5272);
nor U5709 (N_5709,N_5438,N_5227);
and U5710 (N_5710,N_5191,N_5233);
nand U5711 (N_5711,N_5449,N_5498);
nand U5712 (N_5712,N_5360,N_5620);
and U5713 (N_5713,N_5390,N_5414);
or U5714 (N_5714,N_5163,N_5000);
nor U5715 (N_5715,N_5070,N_5298);
nand U5716 (N_5716,N_5431,N_5575);
and U5717 (N_5717,N_5240,N_5305);
or U5718 (N_5718,N_5436,N_5373);
nor U5719 (N_5719,N_5211,N_5445);
and U5720 (N_5720,N_5162,N_5206);
nor U5721 (N_5721,N_5479,N_5170);
or U5722 (N_5722,N_5043,N_5052);
nor U5723 (N_5723,N_5359,N_5142);
nand U5724 (N_5724,N_5357,N_5008);
and U5725 (N_5725,N_5282,N_5126);
xnor U5726 (N_5726,N_5195,N_5118);
or U5727 (N_5727,N_5321,N_5248);
or U5728 (N_5728,N_5493,N_5166);
or U5729 (N_5729,N_5481,N_5005);
nand U5730 (N_5730,N_5297,N_5623);
and U5731 (N_5731,N_5377,N_5291);
and U5732 (N_5732,N_5274,N_5155);
nor U5733 (N_5733,N_5073,N_5454);
or U5734 (N_5734,N_5028,N_5224);
xnor U5735 (N_5735,N_5153,N_5439);
and U5736 (N_5736,N_5192,N_5243);
nand U5737 (N_5737,N_5011,N_5086);
and U5738 (N_5738,N_5388,N_5095);
xor U5739 (N_5739,N_5515,N_5296);
or U5740 (N_5740,N_5235,N_5313);
nand U5741 (N_5741,N_5152,N_5007);
nor U5742 (N_5742,N_5037,N_5289);
or U5743 (N_5743,N_5059,N_5543);
or U5744 (N_5744,N_5113,N_5189);
and U5745 (N_5745,N_5124,N_5209);
nand U5746 (N_5746,N_5429,N_5491);
or U5747 (N_5747,N_5381,N_5606);
nor U5748 (N_5748,N_5290,N_5472);
nor U5749 (N_5749,N_5115,N_5187);
nor U5750 (N_5750,N_5370,N_5398);
or U5751 (N_5751,N_5212,N_5051);
and U5752 (N_5752,N_5453,N_5484);
nand U5753 (N_5753,N_5461,N_5380);
nand U5754 (N_5754,N_5342,N_5465);
nor U5755 (N_5755,N_5148,N_5214);
nand U5756 (N_5756,N_5263,N_5364);
nand U5757 (N_5757,N_5367,N_5404);
nor U5758 (N_5758,N_5507,N_5622);
nand U5759 (N_5759,N_5246,N_5486);
xnor U5760 (N_5760,N_5310,N_5087);
nor U5761 (N_5761,N_5345,N_5060);
nor U5762 (N_5762,N_5396,N_5279);
xor U5763 (N_5763,N_5216,N_5312);
xnor U5764 (N_5764,N_5161,N_5361);
and U5765 (N_5765,N_5492,N_5268);
nand U5766 (N_5766,N_5589,N_5477);
nand U5767 (N_5767,N_5185,N_5046);
and U5768 (N_5768,N_5080,N_5208);
nand U5769 (N_5769,N_5145,N_5555);
and U5770 (N_5770,N_5468,N_5392);
nor U5771 (N_5771,N_5040,N_5247);
or U5772 (N_5772,N_5193,N_5607);
nand U5773 (N_5773,N_5363,N_5420);
nor U5774 (N_5774,N_5389,N_5416);
nor U5775 (N_5775,N_5505,N_5176);
and U5776 (N_5776,N_5428,N_5573);
nor U5777 (N_5777,N_5425,N_5183);
nand U5778 (N_5778,N_5252,N_5265);
nor U5779 (N_5779,N_5190,N_5590);
nor U5780 (N_5780,N_5154,N_5415);
and U5781 (N_5781,N_5613,N_5277);
nor U5782 (N_5782,N_5092,N_5022);
or U5783 (N_5783,N_5053,N_5222);
nand U5784 (N_5784,N_5535,N_5581);
nor U5785 (N_5785,N_5335,N_5242);
and U5786 (N_5786,N_5605,N_5504);
nand U5787 (N_5787,N_5349,N_5547);
nor U5788 (N_5788,N_5418,N_5084);
and U5789 (N_5789,N_5494,N_5294);
nor U5790 (N_5790,N_5201,N_5226);
and U5791 (N_5791,N_5196,N_5456);
nand U5792 (N_5792,N_5221,N_5050);
nand U5793 (N_5793,N_5026,N_5615);
and U5794 (N_5794,N_5485,N_5558);
nand U5795 (N_5795,N_5552,N_5366);
nor U5796 (N_5796,N_5341,N_5333);
and U5797 (N_5797,N_5548,N_5553);
xnor U5798 (N_5798,N_5382,N_5609);
or U5799 (N_5799,N_5378,N_5093);
and U5800 (N_5800,N_5136,N_5064);
nor U5801 (N_5801,N_5101,N_5114);
nor U5802 (N_5802,N_5442,N_5444);
or U5803 (N_5803,N_5077,N_5057);
xor U5804 (N_5804,N_5406,N_5318);
and U5805 (N_5805,N_5569,N_5503);
nor U5806 (N_5806,N_5217,N_5088);
xnor U5807 (N_5807,N_5047,N_5128);
nand U5808 (N_5808,N_5098,N_5232);
xor U5809 (N_5809,N_5119,N_5352);
or U5810 (N_5810,N_5168,N_5476);
or U5811 (N_5811,N_5534,N_5582);
and U5812 (N_5812,N_5139,N_5403);
or U5813 (N_5813,N_5301,N_5521);
or U5814 (N_5814,N_5049,N_5034);
nand U5815 (N_5815,N_5328,N_5565);
and U5816 (N_5816,N_5169,N_5528);
or U5817 (N_5817,N_5085,N_5365);
and U5818 (N_5818,N_5244,N_5508);
and U5819 (N_5819,N_5446,N_5570);
nor U5820 (N_5820,N_5307,N_5537);
nor U5821 (N_5821,N_5250,N_5541);
and U5822 (N_5822,N_5123,N_5134);
or U5823 (N_5823,N_5132,N_5213);
nand U5824 (N_5824,N_5184,N_5271);
nor U5825 (N_5825,N_5374,N_5576);
or U5826 (N_5826,N_5413,N_5023);
nor U5827 (N_5827,N_5422,N_5600);
or U5828 (N_5828,N_5536,N_5526);
nor U5829 (N_5829,N_5447,N_5020);
or U5830 (N_5830,N_5197,N_5351);
nand U5831 (N_5831,N_5002,N_5578);
nor U5832 (N_5832,N_5225,N_5391);
or U5833 (N_5833,N_5397,N_5496);
and U5834 (N_5834,N_5579,N_5350);
nor U5835 (N_5835,N_5106,N_5218);
nand U5836 (N_5836,N_5531,N_5358);
or U5837 (N_5837,N_5280,N_5229);
or U5838 (N_5838,N_5174,N_5015);
xnor U5839 (N_5839,N_5260,N_5336);
nor U5840 (N_5840,N_5068,N_5167);
or U5841 (N_5841,N_5610,N_5262);
nor U5842 (N_5842,N_5482,N_5177);
nor U5843 (N_5843,N_5562,N_5316);
nor U5844 (N_5844,N_5604,N_5116);
xnor U5845 (N_5845,N_5506,N_5393);
and U5846 (N_5846,N_5599,N_5179);
and U5847 (N_5847,N_5487,N_5337);
nor U5848 (N_5848,N_5408,N_5432);
xor U5849 (N_5849,N_5545,N_5130);
or U5850 (N_5850,N_5497,N_5509);
nand U5851 (N_5851,N_5347,N_5467);
and U5852 (N_5852,N_5502,N_5473);
or U5853 (N_5853,N_5512,N_5295);
or U5854 (N_5854,N_5489,N_5198);
nand U5855 (N_5855,N_5157,N_5131);
and U5856 (N_5856,N_5069,N_5058);
nand U5857 (N_5857,N_5385,N_5460);
nor U5858 (N_5858,N_5306,N_5315);
nor U5859 (N_5859,N_5384,N_5514);
and U5860 (N_5860,N_5371,N_5452);
or U5861 (N_5861,N_5223,N_5538);
xnor U5862 (N_5862,N_5003,N_5149);
and U5863 (N_5863,N_5014,N_5045);
or U5864 (N_5864,N_5524,N_5199);
nand U5865 (N_5865,N_5083,N_5203);
nor U5866 (N_5866,N_5499,N_5317);
nand U5867 (N_5867,N_5303,N_5031);
xor U5868 (N_5868,N_5147,N_5182);
and U5869 (N_5869,N_5608,N_5372);
or U5870 (N_5870,N_5027,N_5039);
nand U5871 (N_5871,N_5563,N_5618);
nand U5872 (N_5872,N_5421,N_5427);
and U5873 (N_5873,N_5592,N_5236);
xor U5874 (N_5874,N_5293,N_5593);
xnor U5875 (N_5875,N_5009,N_5257);
or U5876 (N_5876,N_5171,N_5319);
nor U5877 (N_5877,N_5379,N_5256);
or U5878 (N_5878,N_5304,N_5202);
nand U5879 (N_5879,N_5076,N_5544);
nor U5880 (N_5880,N_5331,N_5207);
xor U5881 (N_5881,N_5138,N_5369);
or U5882 (N_5882,N_5309,N_5574);
nand U5883 (N_5883,N_5375,N_5523);
nand U5884 (N_5884,N_5082,N_5571);
xor U5885 (N_5885,N_5424,N_5075);
nor U5886 (N_5886,N_5300,N_5234);
nor U5887 (N_5887,N_5205,N_5325);
and U5888 (N_5888,N_5621,N_5181);
nor U5889 (N_5889,N_5332,N_5160);
nand U5890 (N_5890,N_5159,N_5151);
or U5891 (N_5891,N_5061,N_5276);
and U5892 (N_5892,N_5434,N_5006);
nand U5893 (N_5893,N_5063,N_5580);
nand U5894 (N_5894,N_5488,N_5559);
xnor U5895 (N_5895,N_5117,N_5522);
nor U5896 (N_5896,N_5097,N_5302);
xnor U5897 (N_5897,N_5409,N_5527);
or U5898 (N_5898,N_5387,N_5395);
nor U5899 (N_5899,N_5109,N_5330);
or U5900 (N_5900,N_5018,N_5572);
nor U5901 (N_5901,N_5624,N_5264);
nand U5902 (N_5902,N_5430,N_5228);
xor U5903 (N_5903,N_5568,N_5146);
nand U5904 (N_5904,N_5029,N_5102);
and U5905 (N_5905,N_5518,N_5178);
nand U5906 (N_5906,N_5215,N_5399);
or U5907 (N_5907,N_5411,N_5032);
xor U5908 (N_5908,N_5437,N_5405);
nand U5909 (N_5909,N_5619,N_5469);
and U5910 (N_5910,N_5259,N_5556);
and U5911 (N_5911,N_5546,N_5220);
nor U5912 (N_5912,N_5270,N_5612);
xnor U5913 (N_5913,N_5314,N_5173);
nand U5914 (N_5914,N_5035,N_5601);
and U5915 (N_5915,N_5284,N_5466);
nor U5916 (N_5916,N_5584,N_5587);
nor U5917 (N_5917,N_5323,N_5596);
nor U5918 (N_5918,N_5273,N_5501);
nor U5919 (N_5919,N_5530,N_5326);
xnor U5920 (N_5920,N_5407,N_5617);
nand U5921 (N_5921,N_5019,N_5048);
nand U5922 (N_5922,N_5426,N_5355);
nor U5923 (N_5923,N_5455,N_5062);
nand U5924 (N_5924,N_5033,N_5540);
nor U5925 (N_5925,N_5383,N_5004);
or U5926 (N_5926,N_5400,N_5067);
and U5927 (N_5927,N_5269,N_5474);
nand U5928 (N_5928,N_5001,N_5554);
nor U5929 (N_5929,N_5219,N_5030);
nand U5930 (N_5930,N_5283,N_5529);
nand U5931 (N_5931,N_5616,N_5433);
xnor U5932 (N_5932,N_5165,N_5071);
or U5933 (N_5933,N_5299,N_5200);
and U5934 (N_5934,N_5519,N_5188);
or U5935 (N_5935,N_5419,N_5594);
nor U5936 (N_5936,N_5292,N_5158);
and U5937 (N_5937,N_5602,N_5082);
nand U5938 (N_5938,N_5050,N_5607);
or U5939 (N_5939,N_5342,N_5152);
xnor U5940 (N_5940,N_5534,N_5484);
nor U5941 (N_5941,N_5546,N_5610);
or U5942 (N_5942,N_5441,N_5305);
nand U5943 (N_5943,N_5240,N_5144);
nand U5944 (N_5944,N_5440,N_5250);
or U5945 (N_5945,N_5357,N_5235);
and U5946 (N_5946,N_5522,N_5600);
or U5947 (N_5947,N_5372,N_5585);
or U5948 (N_5948,N_5466,N_5193);
nand U5949 (N_5949,N_5018,N_5071);
xor U5950 (N_5950,N_5251,N_5237);
nand U5951 (N_5951,N_5186,N_5479);
nand U5952 (N_5952,N_5324,N_5399);
nand U5953 (N_5953,N_5468,N_5010);
nand U5954 (N_5954,N_5092,N_5017);
nor U5955 (N_5955,N_5011,N_5315);
xnor U5956 (N_5956,N_5452,N_5420);
and U5957 (N_5957,N_5429,N_5076);
nand U5958 (N_5958,N_5160,N_5500);
nor U5959 (N_5959,N_5269,N_5376);
or U5960 (N_5960,N_5428,N_5442);
nor U5961 (N_5961,N_5518,N_5357);
xor U5962 (N_5962,N_5239,N_5211);
xnor U5963 (N_5963,N_5304,N_5454);
nand U5964 (N_5964,N_5501,N_5271);
nor U5965 (N_5965,N_5082,N_5091);
nor U5966 (N_5966,N_5477,N_5479);
nand U5967 (N_5967,N_5077,N_5461);
and U5968 (N_5968,N_5177,N_5509);
or U5969 (N_5969,N_5437,N_5581);
or U5970 (N_5970,N_5407,N_5485);
or U5971 (N_5971,N_5549,N_5562);
nor U5972 (N_5972,N_5305,N_5433);
or U5973 (N_5973,N_5029,N_5129);
and U5974 (N_5974,N_5016,N_5260);
nand U5975 (N_5975,N_5037,N_5086);
or U5976 (N_5976,N_5528,N_5033);
and U5977 (N_5977,N_5221,N_5381);
or U5978 (N_5978,N_5549,N_5434);
nand U5979 (N_5979,N_5039,N_5257);
and U5980 (N_5980,N_5275,N_5467);
nor U5981 (N_5981,N_5280,N_5497);
nor U5982 (N_5982,N_5447,N_5151);
nand U5983 (N_5983,N_5390,N_5267);
or U5984 (N_5984,N_5566,N_5180);
xnor U5985 (N_5985,N_5245,N_5073);
nand U5986 (N_5986,N_5269,N_5215);
nand U5987 (N_5987,N_5163,N_5301);
or U5988 (N_5988,N_5072,N_5054);
nand U5989 (N_5989,N_5237,N_5479);
or U5990 (N_5990,N_5318,N_5476);
and U5991 (N_5991,N_5606,N_5168);
xnor U5992 (N_5992,N_5345,N_5087);
or U5993 (N_5993,N_5395,N_5334);
or U5994 (N_5994,N_5522,N_5170);
nand U5995 (N_5995,N_5351,N_5231);
or U5996 (N_5996,N_5569,N_5235);
nand U5997 (N_5997,N_5394,N_5355);
nand U5998 (N_5998,N_5198,N_5602);
or U5999 (N_5999,N_5252,N_5103);
and U6000 (N_6000,N_5378,N_5196);
nand U6001 (N_6001,N_5461,N_5331);
or U6002 (N_6002,N_5086,N_5163);
xor U6003 (N_6003,N_5117,N_5490);
nand U6004 (N_6004,N_5480,N_5177);
or U6005 (N_6005,N_5107,N_5234);
nand U6006 (N_6006,N_5285,N_5471);
and U6007 (N_6007,N_5539,N_5549);
nor U6008 (N_6008,N_5104,N_5503);
and U6009 (N_6009,N_5423,N_5026);
xnor U6010 (N_6010,N_5387,N_5231);
nand U6011 (N_6011,N_5572,N_5217);
or U6012 (N_6012,N_5332,N_5107);
nand U6013 (N_6013,N_5434,N_5150);
nand U6014 (N_6014,N_5514,N_5038);
and U6015 (N_6015,N_5302,N_5133);
nand U6016 (N_6016,N_5063,N_5537);
nand U6017 (N_6017,N_5281,N_5432);
or U6018 (N_6018,N_5554,N_5170);
and U6019 (N_6019,N_5428,N_5450);
nor U6020 (N_6020,N_5060,N_5113);
nor U6021 (N_6021,N_5014,N_5150);
or U6022 (N_6022,N_5198,N_5233);
or U6023 (N_6023,N_5155,N_5080);
or U6024 (N_6024,N_5128,N_5461);
or U6025 (N_6025,N_5277,N_5249);
nor U6026 (N_6026,N_5026,N_5249);
nor U6027 (N_6027,N_5507,N_5131);
xnor U6028 (N_6028,N_5093,N_5096);
and U6029 (N_6029,N_5574,N_5037);
and U6030 (N_6030,N_5584,N_5087);
nor U6031 (N_6031,N_5023,N_5114);
or U6032 (N_6032,N_5280,N_5138);
nand U6033 (N_6033,N_5497,N_5158);
nor U6034 (N_6034,N_5050,N_5269);
and U6035 (N_6035,N_5138,N_5359);
nor U6036 (N_6036,N_5164,N_5320);
nor U6037 (N_6037,N_5359,N_5211);
nand U6038 (N_6038,N_5618,N_5028);
nand U6039 (N_6039,N_5318,N_5192);
nor U6040 (N_6040,N_5388,N_5528);
nand U6041 (N_6041,N_5047,N_5414);
nand U6042 (N_6042,N_5141,N_5305);
and U6043 (N_6043,N_5585,N_5341);
nor U6044 (N_6044,N_5019,N_5589);
or U6045 (N_6045,N_5609,N_5273);
nor U6046 (N_6046,N_5174,N_5371);
nor U6047 (N_6047,N_5302,N_5469);
nand U6048 (N_6048,N_5033,N_5373);
xnor U6049 (N_6049,N_5623,N_5620);
and U6050 (N_6050,N_5108,N_5120);
and U6051 (N_6051,N_5468,N_5524);
xnor U6052 (N_6052,N_5169,N_5092);
and U6053 (N_6053,N_5547,N_5139);
or U6054 (N_6054,N_5389,N_5211);
nand U6055 (N_6055,N_5130,N_5350);
nor U6056 (N_6056,N_5569,N_5246);
nand U6057 (N_6057,N_5311,N_5088);
or U6058 (N_6058,N_5063,N_5185);
nor U6059 (N_6059,N_5233,N_5532);
or U6060 (N_6060,N_5006,N_5098);
nor U6061 (N_6061,N_5382,N_5251);
or U6062 (N_6062,N_5133,N_5155);
and U6063 (N_6063,N_5120,N_5144);
nand U6064 (N_6064,N_5110,N_5616);
nand U6065 (N_6065,N_5424,N_5018);
and U6066 (N_6066,N_5443,N_5536);
nor U6067 (N_6067,N_5068,N_5135);
xor U6068 (N_6068,N_5056,N_5304);
nand U6069 (N_6069,N_5437,N_5076);
nand U6070 (N_6070,N_5047,N_5438);
nor U6071 (N_6071,N_5460,N_5454);
nand U6072 (N_6072,N_5553,N_5514);
and U6073 (N_6073,N_5450,N_5321);
and U6074 (N_6074,N_5126,N_5082);
or U6075 (N_6075,N_5569,N_5254);
nand U6076 (N_6076,N_5615,N_5387);
and U6077 (N_6077,N_5437,N_5577);
nand U6078 (N_6078,N_5437,N_5332);
nor U6079 (N_6079,N_5127,N_5613);
nand U6080 (N_6080,N_5586,N_5574);
or U6081 (N_6081,N_5287,N_5482);
and U6082 (N_6082,N_5160,N_5348);
nor U6083 (N_6083,N_5213,N_5182);
or U6084 (N_6084,N_5340,N_5350);
nor U6085 (N_6085,N_5147,N_5383);
or U6086 (N_6086,N_5539,N_5485);
and U6087 (N_6087,N_5519,N_5190);
nand U6088 (N_6088,N_5187,N_5604);
and U6089 (N_6089,N_5418,N_5247);
nor U6090 (N_6090,N_5126,N_5509);
and U6091 (N_6091,N_5240,N_5254);
or U6092 (N_6092,N_5504,N_5067);
or U6093 (N_6093,N_5280,N_5604);
or U6094 (N_6094,N_5039,N_5552);
xnor U6095 (N_6095,N_5033,N_5091);
nand U6096 (N_6096,N_5041,N_5544);
or U6097 (N_6097,N_5227,N_5105);
nand U6098 (N_6098,N_5188,N_5403);
nand U6099 (N_6099,N_5235,N_5040);
and U6100 (N_6100,N_5507,N_5422);
nor U6101 (N_6101,N_5254,N_5601);
and U6102 (N_6102,N_5428,N_5508);
nor U6103 (N_6103,N_5367,N_5529);
and U6104 (N_6104,N_5545,N_5240);
or U6105 (N_6105,N_5313,N_5289);
or U6106 (N_6106,N_5153,N_5235);
nand U6107 (N_6107,N_5465,N_5623);
nor U6108 (N_6108,N_5518,N_5145);
and U6109 (N_6109,N_5115,N_5382);
or U6110 (N_6110,N_5148,N_5438);
nor U6111 (N_6111,N_5344,N_5307);
and U6112 (N_6112,N_5494,N_5623);
or U6113 (N_6113,N_5004,N_5018);
nor U6114 (N_6114,N_5294,N_5220);
or U6115 (N_6115,N_5468,N_5509);
or U6116 (N_6116,N_5355,N_5442);
and U6117 (N_6117,N_5138,N_5433);
or U6118 (N_6118,N_5454,N_5622);
nor U6119 (N_6119,N_5036,N_5556);
nor U6120 (N_6120,N_5502,N_5147);
or U6121 (N_6121,N_5198,N_5620);
nor U6122 (N_6122,N_5283,N_5190);
nand U6123 (N_6123,N_5200,N_5263);
xor U6124 (N_6124,N_5086,N_5077);
or U6125 (N_6125,N_5145,N_5035);
xor U6126 (N_6126,N_5034,N_5590);
nand U6127 (N_6127,N_5496,N_5394);
or U6128 (N_6128,N_5128,N_5433);
and U6129 (N_6129,N_5447,N_5398);
and U6130 (N_6130,N_5500,N_5051);
and U6131 (N_6131,N_5190,N_5011);
or U6132 (N_6132,N_5311,N_5017);
nor U6133 (N_6133,N_5117,N_5404);
or U6134 (N_6134,N_5037,N_5454);
nand U6135 (N_6135,N_5336,N_5404);
nor U6136 (N_6136,N_5067,N_5198);
and U6137 (N_6137,N_5323,N_5273);
nor U6138 (N_6138,N_5444,N_5342);
nand U6139 (N_6139,N_5184,N_5415);
nand U6140 (N_6140,N_5192,N_5555);
nor U6141 (N_6141,N_5189,N_5177);
and U6142 (N_6142,N_5420,N_5036);
and U6143 (N_6143,N_5061,N_5144);
nor U6144 (N_6144,N_5508,N_5530);
xor U6145 (N_6145,N_5460,N_5443);
or U6146 (N_6146,N_5579,N_5233);
nand U6147 (N_6147,N_5337,N_5343);
nand U6148 (N_6148,N_5423,N_5257);
and U6149 (N_6149,N_5381,N_5576);
or U6150 (N_6150,N_5343,N_5314);
or U6151 (N_6151,N_5223,N_5298);
and U6152 (N_6152,N_5204,N_5263);
and U6153 (N_6153,N_5495,N_5374);
nand U6154 (N_6154,N_5412,N_5503);
nand U6155 (N_6155,N_5458,N_5289);
and U6156 (N_6156,N_5537,N_5367);
nand U6157 (N_6157,N_5032,N_5007);
and U6158 (N_6158,N_5297,N_5528);
and U6159 (N_6159,N_5009,N_5311);
nor U6160 (N_6160,N_5545,N_5181);
and U6161 (N_6161,N_5080,N_5288);
nand U6162 (N_6162,N_5157,N_5039);
nand U6163 (N_6163,N_5047,N_5297);
and U6164 (N_6164,N_5087,N_5095);
nor U6165 (N_6165,N_5605,N_5167);
or U6166 (N_6166,N_5134,N_5200);
xor U6167 (N_6167,N_5601,N_5507);
and U6168 (N_6168,N_5272,N_5015);
or U6169 (N_6169,N_5527,N_5525);
nand U6170 (N_6170,N_5293,N_5589);
or U6171 (N_6171,N_5423,N_5471);
nand U6172 (N_6172,N_5178,N_5420);
nor U6173 (N_6173,N_5306,N_5327);
or U6174 (N_6174,N_5091,N_5403);
nand U6175 (N_6175,N_5145,N_5433);
nor U6176 (N_6176,N_5038,N_5113);
and U6177 (N_6177,N_5590,N_5493);
nor U6178 (N_6178,N_5284,N_5401);
nor U6179 (N_6179,N_5346,N_5045);
xor U6180 (N_6180,N_5070,N_5231);
and U6181 (N_6181,N_5477,N_5368);
nor U6182 (N_6182,N_5015,N_5341);
xor U6183 (N_6183,N_5512,N_5317);
nand U6184 (N_6184,N_5437,N_5116);
xnor U6185 (N_6185,N_5328,N_5178);
nor U6186 (N_6186,N_5435,N_5034);
and U6187 (N_6187,N_5375,N_5245);
nor U6188 (N_6188,N_5128,N_5398);
nor U6189 (N_6189,N_5527,N_5624);
xnor U6190 (N_6190,N_5091,N_5152);
and U6191 (N_6191,N_5020,N_5170);
nor U6192 (N_6192,N_5584,N_5311);
and U6193 (N_6193,N_5048,N_5254);
or U6194 (N_6194,N_5387,N_5448);
and U6195 (N_6195,N_5571,N_5392);
nand U6196 (N_6196,N_5277,N_5090);
and U6197 (N_6197,N_5050,N_5327);
and U6198 (N_6198,N_5327,N_5213);
nand U6199 (N_6199,N_5456,N_5122);
nor U6200 (N_6200,N_5005,N_5424);
nor U6201 (N_6201,N_5601,N_5304);
or U6202 (N_6202,N_5521,N_5192);
nand U6203 (N_6203,N_5463,N_5376);
xor U6204 (N_6204,N_5020,N_5048);
nand U6205 (N_6205,N_5423,N_5288);
nand U6206 (N_6206,N_5015,N_5101);
and U6207 (N_6207,N_5001,N_5524);
nand U6208 (N_6208,N_5069,N_5358);
and U6209 (N_6209,N_5222,N_5182);
and U6210 (N_6210,N_5113,N_5436);
nand U6211 (N_6211,N_5241,N_5297);
or U6212 (N_6212,N_5137,N_5246);
and U6213 (N_6213,N_5152,N_5349);
nand U6214 (N_6214,N_5089,N_5341);
and U6215 (N_6215,N_5113,N_5399);
and U6216 (N_6216,N_5573,N_5352);
or U6217 (N_6217,N_5527,N_5220);
nand U6218 (N_6218,N_5605,N_5533);
nand U6219 (N_6219,N_5474,N_5218);
or U6220 (N_6220,N_5554,N_5425);
and U6221 (N_6221,N_5290,N_5209);
and U6222 (N_6222,N_5360,N_5263);
nor U6223 (N_6223,N_5558,N_5006);
and U6224 (N_6224,N_5017,N_5248);
or U6225 (N_6225,N_5379,N_5001);
nor U6226 (N_6226,N_5029,N_5572);
and U6227 (N_6227,N_5514,N_5586);
or U6228 (N_6228,N_5211,N_5599);
or U6229 (N_6229,N_5355,N_5576);
or U6230 (N_6230,N_5295,N_5159);
nand U6231 (N_6231,N_5534,N_5336);
nand U6232 (N_6232,N_5242,N_5078);
nand U6233 (N_6233,N_5500,N_5338);
nor U6234 (N_6234,N_5600,N_5459);
or U6235 (N_6235,N_5255,N_5558);
and U6236 (N_6236,N_5008,N_5350);
or U6237 (N_6237,N_5198,N_5238);
and U6238 (N_6238,N_5464,N_5429);
nor U6239 (N_6239,N_5284,N_5328);
nor U6240 (N_6240,N_5144,N_5058);
or U6241 (N_6241,N_5163,N_5319);
nand U6242 (N_6242,N_5545,N_5463);
nand U6243 (N_6243,N_5074,N_5034);
and U6244 (N_6244,N_5244,N_5261);
nor U6245 (N_6245,N_5023,N_5286);
xnor U6246 (N_6246,N_5099,N_5031);
nand U6247 (N_6247,N_5335,N_5262);
nand U6248 (N_6248,N_5266,N_5165);
nand U6249 (N_6249,N_5506,N_5456);
and U6250 (N_6250,N_5743,N_6039);
nor U6251 (N_6251,N_5749,N_5922);
nand U6252 (N_6252,N_5671,N_6188);
nand U6253 (N_6253,N_6006,N_5795);
nand U6254 (N_6254,N_5694,N_5754);
or U6255 (N_6255,N_5905,N_5869);
nand U6256 (N_6256,N_5627,N_5808);
or U6257 (N_6257,N_5796,N_5681);
nand U6258 (N_6258,N_6068,N_6211);
nor U6259 (N_6259,N_5927,N_6055);
and U6260 (N_6260,N_6123,N_6005);
nor U6261 (N_6261,N_6161,N_6003);
or U6262 (N_6262,N_5937,N_6103);
nand U6263 (N_6263,N_5667,N_6173);
or U6264 (N_6264,N_6023,N_5722);
nand U6265 (N_6265,N_5732,N_5718);
and U6266 (N_6266,N_5946,N_5843);
nor U6267 (N_6267,N_5864,N_5824);
and U6268 (N_6268,N_5800,N_5821);
and U6269 (N_6269,N_5831,N_6079);
nand U6270 (N_6270,N_5952,N_6066);
xnor U6271 (N_6271,N_5924,N_5650);
or U6272 (N_6272,N_5727,N_5962);
nor U6273 (N_6273,N_6091,N_5899);
nor U6274 (N_6274,N_5882,N_5967);
and U6275 (N_6275,N_5879,N_6115);
or U6276 (N_6276,N_5992,N_5972);
nand U6277 (N_6277,N_5928,N_5780);
nor U6278 (N_6278,N_5855,N_5730);
nor U6279 (N_6279,N_6031,N_5716);
xor U6280 (N_6280,N_5707,N_6240);
or U6281 (N_6281,N_5759,N_6108);
or U6282 (N_6282,N_5936,N_6107);
or U6283 (N_6283,N_5745,N_5768);
nand U6284 (N_6284,N_6043,N_6184);
or U6285 (N_6285,N_5920,N_6025);
nand U6286 (N_6286,N_6144,N_5880);
or U6287 (N_6287,N_5932,N_5706);
and U6288 (N_6288,N_5939,N_6232);
or U6289 (N_6289,N_5947,N_5977);
xor U6290 (N_6290,N_6065,N_5642);
nand U6291 (N_6291,N_5987,N_5644);
and U6292 (N_6292,N_6122,N_5645);
nand U6293 (N_6293,N_5819,N_5945);
and U6294 (N_6294,N_5844,N_5878);
nand U6295 (N_6295,N_5704,N_6058);
nand U6296 (N_6296,N_5998,N_5929);
nand U6297 (N_6297,N_6151,N_5734);
and U6298 (N_6298,N_5841,N_6114);
and U6299 (N_6299,N_5753,N_6180);
or U6300 (N_6300,N_6170,N_5894);
nand U6301 (N_6301,N_6247,N_5807);
or U6302 (N_6302,N_5724,N_6221);
and U6303 (N_6303,N_6196,N_5755);
nor U6304 (N_6304,N_5955,N_5832);
or U6305 (N_6305,N_5735,N_5699);
xnor U6306 (N_6306,N_6044,N_6191);
and U6307 (N_6307,N_5911,N_5765);
nor U6308 (N_6308,N_5885,N_5823);
or U6309 (N_6309,N_5961,N_5877);
and U6310 (N_6310,N_5887,N_5690);
nand U6311 (N_6311,N_5784,N_5851);
and U6312 (N_6312,N_5629,N_5763);
and U6313 (N_6313,N_6027,N_5966);
and U6314 (N_6314,N_5838,N_6143);
nand U6315 (N_6315,N_5842,N_6233);
and U6316 (N_6316,N_5982,N_5711);
nand U6317 (N_6317,N_6204,N_5810);
and U6318 (N_6318,N_5640,N_6046);
and U6319 (N_6319,N_6069,N_6018);
xor U6320 (N_6320,N_6064,N_5760);
or U6321 (N_6321,N_6007,N_5981);
and U6322 (N_6322,N_6093,N_6001);
and U6323 (N_6323,N_5625,N_5863);
or U6324 (N_6324,N_5710,N_5648);
nand U6325 (N_6325,N_5781,N_6110);
nor U6326 (N_6326,N_6074,N_5989);
and U6327 (N_6327,N_6073,N_5893);
nor U6328 (N_6328,N_5676,N_5664);
nor U6329 (N_6329,N_5983,N_6036);
nor U6330 (N_6330,N_5756,N_5633);
and U6331 (N_6331,N_6217,N_6015);
nand U6332 (N_6332,N_6234,N_5926);
and U6333 (N_6333,N_6152,N_5956);
or U6334 (N_6334,N_5951,N_5779);
and U6335 (N_6335,N_6150,N_6048);
or U6336 (N_6336,N_5777,N_5752);
nand U6337 (N_6337,N_6220,N_5908);
and U6338 (N_6338,N_5918,N_5666);
and U6339 (N_6339,N_5723,N_6077);
nand U6340 (N_6340,N_5954,N_6155);
nand U6341 (N_6341,N_6212,N_5888);
and U6342 (N_6342,N_5830,N_6215);
or U6343 (N_6343,N_6059,N_5717);
and U6344 (N_6344,N_5767,N_6239);
nor U6345 (N_6345,N_5996,N_5909);
nand U6346 (N_6346,N_5991,N_5801);
nor U6347 (N_6347,N_5873,N_5836);
and U6348 (N_6348,N_6228,N_6021);
nor U6349 (N_6349,N_5653,N_6225);
or U6350 (N_6350,N_5682,N_5935);
nor U6351 (N_6351,N_6094,N_6158);
and U6352 (N_6352,N_5976,N_6100);
xor U6353 (N_6353,N_6072,N_5979);
nand U6354 (N_6354,N_5737,N_6040);
nand U6355 (N_6355,N_6186,N_6218);
nor U6356 (N_6356,N_6181,N_5636);
nand U6357 (N_6357,N_6030,N_6081);
or U6358 (N_6358,N_6208,N_5829);
or U6359 (N_6359,N_5742,N_6197);
xor U6360 (N_6360,N_6037,N_5815);
and U6361 (N_6361,N_6056,N_5845);
nor U6362 (N_6362,N_5953,N_6088);
and U6363 (N_6363,N_5654,N_5900);
or U6364 (N_6364,N_5811,N_5797);
and U6365 (N_6365,N_6060,N_6226);
and U6366 (N_6366,N_5805,N_5680);
and U6367 (N_6367,N_6095,N_6129);
nor U6368 (N_6368,N_6019,N_5974);
and U6369 (N_6369,N_5884,N_6085);
nand U6370 (N_6370,N_5867,N_5943);
nand U6371 (N_6371,N_5688,N_5798);
nor U6372 (N_6372,N_6185,N_5930);
nand U6373 (N_6373,N_5912,N_6216);
or U6374 (N_6374,N_5720,N_6131);
xor U6375 (N_6375,N_5816,N_5766);
nor U6376 (N_6376,N_6175,N_5835);
nor U6377 (N_6377,N_5631,N_5698);
nand U6378 (N_6378,N_6206,N_6138);
and U6379 (N_6379,N_6053,N_5738);
nor U6380 (N_6380,N_5751,N_5695);
or U6381 (N_6381,N_5701,N_5782);
nor U6382 (N_6382,N_6080,N_6246);
or U6383 (N_6383,N_5874,N_6016);
nor U6384 (N_6384,N_6013,N_6200);
nand U6385 (N_6385,N_6078,N_5638);
and U6386 (N_6386,N_6116,N_5837);
nand U6387 (N_6387,N_6125,N_5973);
nor U6388 (N_6388,N_5705,N_6238);
and U6389 (N_6389,N_6047,N_5702);
and U6390 (N_6390,N_5849,N_6210);
nand U6391 (N_6391,N_5794,N_5985);
or U6392 (N_6392,N_6199,N_6130);
nor U6393 (N_6393,N_5890,N_5964);
nor U6394 (N_6394,N_6194,N_5971);
and U6395 (N_6395,N_5813,N_5969);
nor U6396 (N_6396,N_6222,N_6086);
nor U6397 (N_6397,N_5856,N_5659);
or U6398 (N_6398,N_6174,N_6178);
and U6399 (N_6399,N_5881,N_6229);
nor U6400 (N_6400,N_6148,N_5689);
nor U6401 (N_6401,N_6145,N_5812);
and U6402 (N_6402,N_6169,N_6004);
xor U6403 (N_6403,N_5806,N_5906);
nor U6404 (N_6404,N_6231,N_6172);
and U6405 (N_6405,N_5921,N_6000);
nor U6406 (N_6406,N_5792,N_5628);
or U6407 (N_6407,N_5809,N_5703);
nor U6408 (N_6408,N_5957,N_5715);
nand U6409 (N_6409,N_6244,N_5630);
or U6410 (N_6410,N_5713,N_5787);
nor U6411 (N_6411,N_5822,N_5803);
or U6412 (N_6412,N_6045,N_6032);
nand U6413 (N_6413,N_6242,N_6083);
and U6414 (N_6414,N_5750,N_6248);
and U6415 (N_6415,N_5660,N_5901);
nor U6416 (N_6416,N_5891,N_5687);
nand U6417 (N_6417,N_5938,N_6024);
nand U6418 (N_6418,N_6099,N_6028);
and U6419 (N_6419,N_6219,N_5686);
or U6420 (N_6420,N_5643,N_6054);
and U6421 (N_6421,N_5775,N_5913);
nor U6422 (N_6422,N_6142,N_5649);
nand U6423 (N_6423,N_5791,N_5774);
and U6424 (N_6424,N_6163,N_6193);
or U6425 (N_6425,N_6026,N_5963);
nor U6426 (N_6426,N_6097,N_5778);
nor U6427 (N_6427,N_6136,N_5728);
nand U6428 (N_6428,N_6121,N_5761);
and U6429 (N_6429,N_6195,N_5948);
nor U6430 (N_6430,N_5871,N_5719);
nor U6431 (N_6431,N_5818,N_6230);
xnor U6432 (N_6432,N_5958,N_5865);
and U6433 (N_6433,N_5656,N_5714);
xnor U6434 (N_6434,N_5726,N_6101);
or U6435 (N_6435,N_5652,N_5684);
and U6436 (N_6436,N_5708,N_6109);
or U6437 (N_6437,N_6166,N_5731);
or U6438 (N_6438,N_5786,N_5984);
or U6439 (N_6439,N_5923,N_5839);
nor U6440 (N_6440,N_5758,N_6147);
and U6441 (N_6441,N_5739,N_5919);
and U6442 (N_6442,N_6223,N_5949);
nand U6443 (N_6443,N_6162,N_5744);
and U6444 (N_6444,N_5626,N_6192);
and U6445 (N_6445,N_6070,N_5826);
or U6446 (N_6446,N_5783,N_6017);
xnor U6447 (N_6447,N_5651,N_5675);
and U6448 (N_6448,N_5903,N_5757);
nor U6449 (N_6449,N_5902,N_6190);
and U6450 (N_6450,N_6042,N_6035);
and U6451 (N_6451,N_5910,N_6243);
or U6452 (N_6452,N_5988,N_6160);
nand U6453 (N_6453,N_6237,N_5725);
and U6454 (N_6454,N_5833,N_6057);
and U6455 (N_6455,N_6159,N_5868);
xnor U6456 (N_6456,N_5875,N_6133);
and U6457 (N_6457,N_5799,N_5931);
nand U6458 (N_6458,N_5915,N_6082);
nor U6459 (N_6459,N_6033,N_5670);
or U6460 (N_6460,N_5736,N_5933);
nor U6461 (N_6461,N_6061,N_5848);
nand U6462 (N_6462,N_6182,N_5986);
nand U6463 (N_6463,N_5916,N_5729);
nor U6464 (N_6464,N_5995,N_6168);
and U6465 (N_6465,N_5870,N_5999);
nor U6466 (N_6466,N_5662,N_6149);
nor U6467 (N_6467,N_5917,N_5944);
and U6468 (N_6468,N_5860,N_6227);
nor U6469 (N_6469,N_5857,N_6124);
or U6470 (N_6470,N_6127,N_5997);
nand U6471 (N_6471,N_5709,N_6090);
xor U6472 (N_6472,N_5655,N_5770);
or U6473 (N_6473,N_6012,N_6126);
nor U6474 (N_6474,N_6096,N_5691);
nand U6475 (N_6475,N_5960,N_6112);
nand U6476 (N_6476,N_6209,N_5748);
and U6477 (N_6477,N_5692,N_6120);
and U6478 (N_6478,N_5883,N_5771);
and U6479 (N_6479,N_6245,N_5641);
and U6480 (N_6480,N_5785,N_5892);
and U6481 (N_6481,N_5634,N_6117);
nor U6482 (N_6482,N_5980,N_5975);
xor U6483 (N_6483,N_6249,N_6213);
nand U6484 (N_6484,N_5828,N_5677);
xor U6485 (N_6485,N_6075,N_6177);
xnor U6486 (N_6486,N_5668,N_5802);
nand U6487 (N_6487,N_5789,N_5788);
and U6488 (N_6488,N_6119,N_6098);
and U6489 (N_6489,N_5862,N_5978);
or U6490 (N_6490,N_5657,N_6128);
nand U6491 (N_6491,N_6179,N_5934);
and U6492 (N_6492,N_6157,N_6171);
or U6493 (N_6493,N_5683,N_6187);
nand U6494 (N_6494,N_6153,N_5696);
nor U6495 (N_6495,N_6164,N_5853);
nor U6496 (N_6496,N_5721,N_5847);
and U6497 (N_6497,N_6076,N_5854);
and U6498 (N_6498,N_6014,N_6106);
nor U6499 (N_6499,N_6224,N_5950);
nand U6500 (N_6500,N_5994,N_5672);
nor U6501 (N_6501,N_5674,N_5876);
nand U6502 (N_6502,N_6111,N_5632);
nand U6503 (N_6503,N_5942,N_6049);
or U6504 (N_6504,N_5693,N_6029);
and U6505 (N_6505,N_5872,N_6214);
or U6506 (N_6506,N_6011,N_5740);
nor U6507 (N_6507,N_5663,N_6205);
or U6508 (N_6508,N_6137,N_6020);
and U6509 (N_6509,N_5846,N_5673);
xor U6510 (N_6510,N_6201,N_5817);
nand U6511 (N_6511,N_5793,N_5968);
nor U6512 (N_6512,N_5697,N_6102);
and U6513 (N_6513,N_5762,N_6009);
or U6514 (N_6514,N_6118,N_6235);
and U6515 (N_6515,N_5904,N_6241);
and U6516 (N_6516,N_5993,N_6135);
nand U6517 (N_6517,N_6156,N_5858);
nand U6518 (N_6518,N_6203,N_5637);
nand U6519 (N_6519,N_6050,N_6134);
and U6520 (N_6520,N_6146,N_6132);
and U6521 (N_6521,N_6105,N_5679);
nor U6522 (N_6522,N_6008,N_6198);
xor U6523 (N_6523,N_5940,N_6022);
nand U6524 (N_6524,N_6154,N_5814);
and U6525 (N_6525,N_6087,N_5685);
and U6526 (N_6526,N_6067,N_5861);
nand U6527 (N_6527,N_6071,N_6141);
nand U6528 (N_6528,N_6062,N_5866);
nand U6529 (N_6529,N_5850,N_6084);
nand U6530 (N_6530,N_5769,N_5914);
or U6531 (N_6531,N_5852,N_5635);
xor U6532 (N_6532,N_5941,N_5700);
and U6533 (N_6533,N_5907,N_5804);
nand U6534 (N_6534,N_5897,N_5790);
and U6535 (N_6535,N_6140,N_6113);
nor U6536 (N_6536,N_6236,N_6010);
and U6537 (N_6537,N_5741,N_6063);
nor U6538 (N_6538,N_6051,N_5820);
xor U6539 (N_6539,N_5639,N_6165);
or U6540 (N_6540,N_5665,N_5747);
and U6541 (N_6541,N_6041,N_5859);
and U6542 (N_6542,N_5712,N_5990);
nand U6543 (N_6543,N_5647,N_5678);
nor U6544 (N_6544,N_6002,N_5773);
and U6545 (N_6545,N_6104,N_5669);
nand U6546 (N_6546,N_6202,N_6034);
and U6547 (N_6547,N_5772,N_5746);
nand U6548 (N_6548,N_5827,N_5970);
and U6549 (N_6549,N_6176,N_5658);
or U6550 (N_6550,N_5886,N_5646);
and U6551 (N_6551,N_5834,N_5840);
and U6552 (N_6552,N_5661,N_5776);
and U6553 (N_6553,N_6183,N_5895);
nor U6554 (N_6554,N_5898,N_6038);
and U6555 (N_6555,N_6089,N_5896);
nand U6556 (N_6556,N_5764,N_5733);
nand U6557 (N_6557,N_5959,N_5925);
nor U6558 (N_6558,N_5889,N_5965);
and U6559 (N_6559,N_6189,N_6167);
and U6560 (N_6560,N_6052,N_5825);
nand U6561 (N_6561,N_6207,N_6092);
or U6562 (N_6562,N_6139,N_6090);
or U6563 (N_6563,N_6076,N_5890);
nand U6564 (N_6564,N_5888,N_5820);
nor U6565 (N_6565,N_6011,N_5625);
nor U6566 (N_6566,N_6218,N_6123);
nor U6567 (N_6567,N_5735,N_6042);
nor U6568 (N_6568,N_5803,N_6120);
and U6569 (N_6569,N_5813,N_6249);
nor U6570 (N_6570,N_6177,N_5908);
nor U6571 (N_6571,N_5636,N_5857);
nand U6572 (N_6572,N_5631,N_6026);
and U6573 (N_6573,N_6176,N_6036);
or U6574 (N_6574,N_5789,N_5667);
nor U6575 (N_6575,N_5763,N_5916);
or U6576 (N_6576,N_6018,N_5777);
and U6577 (N_6577,N_5864,N_5974);
nor U6578 (N_6578,N_5975,N_6048);
nand U6579 (N_6579,N_5911,N_5799);
or U6580 (N_6580,N_6214,N_6110);
or U6581 (N_6581,N_6085,N_6094);
and U6582 (N_6582,N_5782,N_5653);
xnor U6583 (N_6583,N_5861,N_6129);
and U6584 (N_6584,N_6226,N_5977);
and U6585 (N_6585,N_5745,N_5705);
xnor U6586 (N_6586,N_6155,N_5719);
nor U6587 (N_6587,N_5644,N_6126);
and U6588 (N_6588,N_5746,N_6150);
nand U6589 (N_6589,N_5691,N_5673);
nor U6590 (N_6590,N_6110,N_6120);
or U6591 (N_6591,N_6157,N_6016);
or U6592 (N_6592,N_5722,N_5782);
or U6593 (N_6593,N_6058,N_6147);
nand U6594 (N_6594,N_5991,N_5659);
nand U6595 (N_6595,N_6019,N_5904);
nand U6596 (N_6596,N_5644,N_5999);
or U6597 (N_6597,N_6140,N_6033);
nand U6598 (N_6598,N_5756,N_5807);
xor U6599 (N_6599,N_5686,N_5762);
or U6600 (N_6600,N_5665,N_5694);
or U6601 (N_6601,N_5639,N_5753);
or U6602 (N_6602,N_5738,N_5793);
and U6603 (N_6603,N_6222,N_6228);
and U6604 (N_6604,N_6205,N_6209);
nor U6605 (N_6605,N_5937,N_6066);
nand U6606 (N_6606,N_5650,N_5701);
or U6607 (N_6607,N_6231,N_6150);
xor U6608 (N_6608,N_5661,N_6057);
or U6609 (N_6609,N_6021,N_6026);
or U6610 (N_6610,N_6148,N_6146);
and U6611 (N_6611,N_5729,N_6024);
and U6612 (N_6612,N_5717,N_6079);
nor U6613 (N_6613,N_5756,N_6244);
xor U6614 (N_6614,N_6059,N_6184);
nor U6615 (N_6615,N_6082,N_5833);
nand U6616 (N_6616,N_6213,N_5795);
or U6617 (N_6617,N_6139,N_5782);
nand U6618 (N_6618,N_5892,N_5749);
or U6619 (N_6619,N_5808,N_5824);
and U6620 (N_6620,N_6104,N_6038);
and U6621 (N_6621,N_5902,N_6037);
and U6622 (N_6622,N_5972,N_5681);
or U6623 (N_6623,N_5806,N_5977);
or U6624 (N_6624,N_5630,N_6170);
nand U6625 (N_6625,N_6072,N_6169);
and U6626 (N_6626,N_5667,N_6234);
nand U6627 (N_6627,N_5968,N_5989);
or U6628 (N_6628,N_5865,N_5634);
or U6629 (N_6629,N_5955,N_6029);
nand U6630 (N_6630,N_5917,N_6123);
nand U6631 (N_6631,N_5785,N_5764);
or U6632 (N_6632,N_5841,N_5772);
and U6633 (N_6633,N_6131,N_5823);
nor U6634 (N_6634,N_5988,N_5983);
or U6635 (N_6635,N_5664,N_6192);
or U6636 (N_6636,N_5845,N_5902);
and U6637 (N_6637,N_5942,N_5751);
and U6638 (N_6638,N_5853,N_5733);
or U6639 (N_6639,N_5758,N_6110);
nand U6640 (N_6640,N_5885,N_5792);
nor U6641 (N_6641,N_6103,N_6026);
and U6642 (N_6642,N_6100,N_6207);
xor U6643 (N_6643,N_6088,N_5643);
nor U6644 (N_6644,N_5703,N_6127);
nor U6645 (N_6645,N_5927,N_5791);
nand U6646 (N_6646,N_5751,N_5741);
and U6647 (N_6647,N_5795,N_5697);
and U6648 (N_6648,N_5706,N_5657);
nand U6649 (N_6649,N_5637,N_5648);
and U6650 (N_6650,N_5924,N_6100);
and U6651 (N_6651,N_5645,N_5820);
and U6652 (N_6652,N_5628,N_5866);
or U6653 (N_6653,N_6072,N_5800);
or U6654 (N_6654,N_5757,N_6173);
and U6655 (N_6655,N_5952,N_6022);
or U6656 (N_6656,N_6002,N_5643);
or U6657 (N_6657,N_6184,N_6027);
nand U6658 (N_6658,N_5739,N_5716);
nor U6659 (N_6659,N_5979,N_5799);
and U6660 (N_6660,N_6021,N_5801);
or U6661 (N_6661,N_5796,N_6037);
nor U6662 (N_6662,N_6065,N_5771);
nor U6663 (N_6663,N_5903,N_5893);
nor U6664 (N_6664,N_5629,N_6105);
and U6665 (N_6665,N_6112,N_5787);
nor U6666 (N_6666,N_5765,N_5666);
xor U6667 (N_6667,N_5912,N_5865);
nor U6668 (N_6668,N_5955,N_6048);
xor U6669 (N_6669,N_5898,N_6133);
or U6670 (N_6670,N_6198,N_5655);
xnor U6671 (N_6671,N_5854,N_6052);
and U6672 (N_6672,N_5964,N_6225);
nor U6673 (N_6673,N_5692,N_5836);
xor U6674 (N_6674,N_6209,N_5848);
nor U6675 (N_6675,N_6202,N_5780);
nand U6676 (N_6676,N_6038,N_6246);
or U6677 (N_6677,N_6055,N_6123);
nor U6678 (N_6678,N_6009,N_5629);
nor U6679 (N_6679,N_5907,N_5978);
nand U6680 (N_6680,N_5732,N_5700);
and U6681 (N_6681,N_5986,N_6174);
and U6682 (N_6682,N_5733,N_5953);
nor U6683 (N_6683,N_5788,N_5912);
and U6684 (N_6684,N_6163,N_5776);
nand U6685 (N_6685,N_5831,N_5827);
nor U6686 (N_6686,N_6095,N_5905);
or U6687 (N_6687,N_6123,N_5918);
nand U6688 (N_6688,N_6106,N_5999);
or U6689 (N_6689,N_6212,N_6055);
or U6690 (N_6690,N_5786,N_5957);
or U6691 (N_6691,N_5815,N_5921);
nand U6692 (N_6692,N_6193,N_5667);
nor U6693 (N_6693,N_5888,N_6140);
nor U6694 (N_6694,N_5904,N_5985);
and U6695 (N_6695,N_5944,N_5879);
nor U6696 (N_6696,N_5765,N_6194);
and U6697 (N_6697,N_5754,N_5805);
nor U6698 (N_6698,N_5732,N_6068);
and U6699 (N_6699,N_5926,N_5990);
nor U6700 (N_6700,N_6039,N_5908);
nor U6701 (N_6701,N_5873,N_6011);
or U6702 (N_6702,N_5706,N_6209);
and U6703 (N_6703,N_5976,N_5778);
nand U6704 (N_6704,N_5848,N_5707);
nand U6705 (N_6705,N_6170,N_5875);
nor U6706 (N_6706,N_5628,N_6050);
nor U6707 (N_6707,N_5914,N_5902);
or U6708 (N_6708,N_5881,N_5902);
nand U6709 (N_6709,N_5745,N_5998);
and U6710 (N_6710,N_6124,N_5661);
or U6711 (N_6711,N_5943,N_5701);
xor U6712 (N_6712,N_6163,N_6125);
xnor U6713 (N_6713,N_6208,N_6009);
and U6714 (N_6714,N_5718,N_5670);
and U6715 (N_6715,N_6161,N_5745);
and U6716 (N_6716,N_5729,N_5978);
nor U6717 (N_6717,N_5828,N_6042);
or U6718 (N_6718,N_5799,N_5780);
and U6719 (N_6719,N_6248,N_5633);
or U6720 (N_6720,N_5951,N_5974);
nand U6721 (N_6721,N_6130,N_6150);
and U6722 (N_6722,N_5858,N_5848);
and U6723 (N_6723,N_5725,N_6092);
nand U6724 (N_6724,N_5988,N_5832);
nand U6725 (N_6725,N_5658,N_5680);
or U6726 (N_6726,N_5978,N_5934);
nand U6727 (N_6727,N_6185,N_5824);
nor U6728 (N_6728,N_5824,N_6108);
nand U6729 (N_6729,N_6010,N_5632);
nor U6730 (N_6730,N_5981,N_5906);
nand U6731 (N_6731,N_5811,N_5972);
nand U6732 (N_6732,N_5758,N_5802);
and U6733 (N_6733,N_6233,N_6044);
and U6734 (N_6734,N_6039,N_5696);
or U6735 (N_6735,N_5987,N_6172);
xor U6736 (N_6736,N_5822,N_5735);
or U6737 (N_6737,N_6098,N_5839);
and U6738 (N_6738,N_5769,N_5897);
nor U6739 (N_6739,N_5976,N_5761);
or U6740 (N_6740,N_5947,N_6208);
nor U6741 (N_6741,N_5882,N_5672);
nor U6742 (N_6742,N_5710,N_5770);
or U6743 (N_6743,N_5735,N_5640);
nand U6744 (N_6744,N_6063,N_5667);
and U6745 (N_6745,N_5745,N_5889);
or U6746 (N_6746,N_6119,N_5768);
nor U6747 (N_6747,N_5845,N_5846);
and U6748 (N_6748,N_5902,N_6047);
or U6749 (N_6749,N_5821,N_5869);
xnor U6750 (N_6750,N_5738,N_5769);
or U6751 (N_6751,N_5788,N_5792);
nor U6752 (N_6752,N_6244,N_5811);
nor U6753 (N_6753,N_6115,N_5685);
or U6754 (N_6754,N_6191,N_5801);
nand U6755 (N_6755,N_6148,N_5875);
and U6756 (N_6756,N_5987,N_5769);
nand U6757 (N_6757,N_5989,N_5813);
and U6758 (N_6758,N_5787,N_5756);
or U6759 (N_6759,N_5895,N_5633);
and U6760 (N_6760,N_6098,N_6173);
nor U6761 (N_6761,N_5645,N_6217);
nor U6762 (N_6762,N_5782,N_6115);
and U6763 (N_6763,N_6246,N_5690);
and U6764 (N_6764,N_5695,N_5881);
and U6765 (N_6765,N_5964,N_5825);
or U6766 (N_6766,N_5698,N_6104);
or U6767 (N_6767,N_5704,N_6247);
and U6768 (N_6768,N_6235,N_5958);
or U6769 (N_6769,N_5958,N_6079);
or U6770 (N_6770,N_5879,N_6093);
or U6771 (N_6771,N_6026,N_6015);
and U6772 (N_6772,N_6215,N_5928);
xor U6773 (N_6773,N_6058,N_5653);
and U6774 (N_6774,N_5730,N_5816);
nand U6775 (N_6775,N_5732,N_5751);
and U6776 (N_6776,N_6206,N_6189);
nor U6777 (N_6777,N_5644,N_5746);
and U6778 (N_6778,N_5938,N_5903);
and U6779 (N_6779,N_6100,N_5675);
and U6780 (N_6780,N_5774,N_5730);
nor U6781 (N_6781,N_5974,N_6075);
nor U6782 (N_6782,N_5979,N_5900);
and U6783 (N_6783,N_6015,N_6023);
and U6784 (N_6784,N_6138,N_6063);
nand U6785 (N_6785,N_6248,N_5713);
and U6786 (N_6786,N_5802,N_6066);
or U6787 (N_6787,N_5744,N_5709);
or U6788 (N_6788,N_5669,N_5719);
or U6789 (N_6789,N_5802,N_5751);
or U6790 (N_6790,N_6124,N_5680);
or U6791 (N_6791,N_6072,N_5766);
and U6792 (N_6792,N_6155,N_5736);
nor U6793 (N_6793,N_6015,N_6095);
nand U6794 (N_6794,N_5849,N_5694);
and U6795 (N_6795,N_6084,N_5627);
nand U6796 (N_6796,N_6183,N_5746);
nand U6797 (N_6797,N_6232,N_5802);
nand U6798 (N_6798,N_6115,N_5854);
nand U6799 (N_6799,N_5662,N_5932);
and U6800 (N_6800,N_6243,N_5836);
and U6801 (N_6801,N_5869,N_5892);
and U6802 (N_6802,N_5760,N_5951);
nor U6803 (N_6803,N_5695,N_5849);
or U6804 (N_6804,N_5704,N_5821);
or U6805 (N_6805,N_5645,N_5641);
and U6806 (N_6806,N_5748,N_6121);
nor U6807 (N_6807,N_6183,N_6026);
nand U6808 (N_6808,N_6051,N_6193);
nand U6809 (N_6809,N_5805,N_5762);
nor U6810 (N_6810,N_5687,N_6215);
nand U6811 (N_6811,N_5836,N_5888);
nor U6812 (N_6812,N_6202,N_6028);
nand U6813 (N_6813,N_5862,N_6177);
nor U6814 (N_6814,N_6211,N_6199);
and U6815 (N_6815,N_5629,N_6091);
and U6816 (N_6816,N_6065,N_5723);
and U6817 (N_6817,N_5675,N_5995);
xor U6818 (N_6818,N_6039,N_6216);
xor U6819 (N_6819,N_5687,N_5893);
nor U6820 (N_6820,N_6052,N_5938);
or U6821 (N_6821,N_5906,N_5680);
nor U6822 (N_6822,N_6226,N_5727);
or U6823 (N_6823,N_6002,N_5969);
nand U6824 (N_6824,N_5650,N_5778);
and U6825 (N_6825,N_5863,N_5744);
and U6826 (N_6826,N_6229,N_6211);
or U6827 (N_6827,N_6222,N_6016);
and U6828 (N_6828,N_5927,N_6099);
xnor U6829 (N_6829,N_6094,N_5908);
xnor U6830 (N_6830,N_6073,N_5918);
or U6831 (N_6831,N_5878,N_5871);
nand U6832 (N_6832,N_5963,N_5641);
or U6833 (N_6833,N_5734,N_5993);
nor U6834 (N_6834,N_5763,N_5737);
nor U6835 (N_6835,N_5794,N_5720);
and U6836 (N_6836,N_6090,N_6200);
and U6837 (N_6837,N_6081,N_6149);
nand U6838 (N_6838,N_5732,N_6184);
nand U6839 (N_6839,N_5650,N_5830);
xnor U6840 (N_6840,N_5865,N_6027);
nand U6841 (N_6841,N_6050,N_6233);
xnor U6842 (N_6842,N_6098,N_6120);
nor U6843 (N_6843,N_5882,N_5734);
nor U6844 (N_6844,N_5746,N_6191);
and U6845 (N_6845,N_6231,N_5738);
nand U6846 (N_6846,N_5784,N_6192);
and U6847 (N_6847,N_6047,N_6079);
and U6848 (N_6848,N_6211,N_6140);
and U6849 (N_6849,N_5917,N_5689);
nand U6850 (N_6850,N_6083,N_5776);
and U6851 (N_6851,N_6052,N_5857);
and U6852 (N_6852,N_5746,N_5990);
and U6853 (N_6853,N_6003,N_5746);
or U6854 (N_6854,N_5958,N_5997);
and U6855 (N_6855,N_5810,N_6008);
nor U6856 (N_6856,N_5830,N_6180);
nor U6857 (N_6857,N_5941,N_6211);
nor U6858 (N_6858,N_5709,N_5939);
and U6859 (N_6859,N_5858,N_5931);
nor U6860 (N_6860,N_6194,N_6001);
xnor U6861 (N_6861,N_5842,N_5629);
or U6862 (N_6862,N_5930,N_5854);
or U6863 (N_6863,N_5820,N_6193);
nand U6864 (N_6864,N_5713,N_6175);
nand U6865 (N_6865,N_5721,N_5851);
or U6866 (N_6866,N_6149,N_5926);
xor U6867 (N_6867,N_6102,N_6216);
xnor U6868 (N_6868,N_5752,N_5998);
or U6869 (N_6869,N_5751,N_5814);
or U6870 (N_6870,N_5952,N_6173);
or U6871 (N_6871,N_5790,N_6236);
nor U6872 (N_6872,N_5886,N_5896);
and U6873 (N_6873,N_6244,N_6248);
or U6874 (N_6874,N_6172,N_6041);
nand U6875 (N_6875,N_6624,N_6413);
nor U6876 (N_6876,N_6850,N_6851);
nor U6877 (N_6877,N_6581,N_6779);
and U6878 (N_6878,N_6504,N_6337);
nand U6879 (N_6879,N_6522,N_6476);
and U6880 (N_6880,N_6620,N_6398);
or U6881 (N_6881,N_6562,N_6285);
nand U6882 (N_6882,N_6558,N_6843);
and U6883 (N_6883,N_6422,N_6344);
xor U6884 (N_6884,N_6724,N_6683);
nor U6885 (N_6885,N_6467,N_6553);
xnor U6886 (N_6886,N_6689,N_6421);
or U6887 (N_6887,N_6294,N_6685);
and U6888 (N_6888,N_6286,N_6796);
or U6889 (N_6889,N_6387,N_6812);
xor U6890 (N_6890,N_6308,N_6697);
xor U6891 (N_6891,N_6717,N_6824);
or U6892 (N_6892,N_6813,N_6551);
and U6893 (N_6893,N_6384,N_6556);
nand U6894 (N_6894,N_6680,N_6486);
and U6895 (N_6895,N_6602,N_6383);
nand U6896 (N_6896,N_6479,N_6477);
nor U6897 (N_6897,N_6371,N_6858);
nand U6898 (N_6898,N_6280,N_6712);
xnor U6899 (N_6899,N_6678,N_6874);
xor U6900 (N_6900,N_6475,N_6441);
and U6901 (N_6901,N_6437,N_6676);
nor U6902 (N_6902,N_6391,N_6364);
or U6903 (N_6903,N_6764,N_6317);
nand U6904 (N_6904,N_6381,N_6834);
or U6905 (N_6905,N_6729,N_6292);
nand U6906 (N_6906,N_6456,N_6540);
nand U6907 (N_6907,N_6695,N_6320);
and U6908 (N_6908,N_6810,N_6619);
nand U6909 (N_6909,N_6284,N_6502);
nor U6910 (N_6910,N_6466,N_6866);
nor U6911 (N_6911,N_6636,N_6761);
and U6912 (N_6912,N_6762,N_6262);
xor U6913 (N_6913,N_6261,N_6301);
or U6914 (N_6914,N_6291,N_6626);
nand U6915 (N_6915,N_6559,N_6849);
and U6916 (N_6916,N_6404,N_6330);
or U6917 (N_6917,N_6640,N_6657);
nor U6918 (N_6918,N_6842,N_6472);
or U6919 (N_6919,N_6478,N_6811);
nand U6920 (N_6920,N_6591,N_6436);
nor U6921 (N_6921,N_6801,N_6679);
and U6922 (N_6922,N_6424,N_6855);
or U6923 (N_6923,N_6860,N_6726);
and U6924 (N_6924,N_6840,N_6661);
and U6925 (N_6925,N_6783,N_6411);
xnor U6926 (N_6926,N_6596,N_6463);
and U6927 (N_6927,N_6608,N_6823);
nor U6928 (N_6928,N_6854,N_6703);
nand U6929 (N_6929,N_6482,N_6484);
nor U6930 (N_6930,N_6684,N_6868);
or U6931 (N_6931,N_6838,N_6716);
nor U6932 (N_6932,N_6373,N_6848);
nand U6933 (N_6933,N_6544,N_6450);
nand U6934 (N_6934,N_6580,N_6628);
nor U6935 (N_6935,N_6749,N_6609);
xor U6936 (N_6936,N_6816,N_6741);
xnor U6937 (N_6937,N_6664,N_6377);
and U6938 (N_6938,N_6431,N_6615);
nand U6939 (N_6939,N_6417,N_6819);
nor U6940 (N_6940,N_6786,N_6535);
nand U6941 (N_6941,N_6662,N_6293);
or U6942 (N_6942,N_6362,N_6338);
or U6943 (N_6943,N_6639,N_6370);
and U6944 (N_6944,N_6673,N_6601);
and U6945 (N_6945,N_6603,N_6752);
and U6946 (N_6946,N_6407,N_6405);
nor U6947 (N_6947,N_6473,N_6587);
nand U6948 (N_6948,N_6395,N_6805);
or U6949 (N_6949,N_6412,N_6414);
nand U6950 (N_6950,N_6790,N_6550);
nand U6951 (N_6951,N_6461,N_6462);
or U6952 (N_6952,N_6598,N_6825);
or U6953 (N_6953,N_6314,N_6385);
nand U6954 (N_6954,N_6444,N_6361);
nand U6955 (N_6955,N_6375,N_6423);
nor U6956 (N_6956,N_6577,N_6382);
or U6957 (N_6957,N_6541,N_6299);
and U6958 (N_6958,N_6629,N_6600);
nand U6959 (N_6959,N_6442,N_6497);
nand U6960 (N_6960,N_6250,N_6483);
nand U6961 (N_6961,N_6465,N_6593);
and U6962 (N_6962,N_6523,N_6705);
nor U6963 (N_6963,N_6605,N_6372);
nand U6964 (N_6964,N_6429,N_6794);
or U6965 (N_6965,N_6651,N_6506);
nand U6966 (N_6966,N_6270,N_6536);
nand U6967 (N_6967,N_6799,N_6510);
nor U6968 (N_6968,N_6806,N_6710);
nand U6969 (N_6969,N_6302,N_6743);
nand U6970 (N_6970,N_6297,N_6433);
xnor U6971 (N_6971,N_6516,N_6788);
nand U6972 (N_6972,N_6348,N_6627);
nor U6973 (N_6973,N_6425,N_6784);
nor U6974 (N_6974,N_6588,N_6759);
or U6975 (N_6975,N_6457,N_6528);
nand U6976 (N_6976,N_6720,N_6833);
nor U6977 (N_6977,N_6800,N_6768);
nand U6978 (N_6978,N_6730,N_6765);
or U6979 (N_6979,N_6599,N_6458);
nand U6980 (N_6980,N_6756,N_6363);
nand U6981 (N_6981,N_6872,N_6728);
nand U6982 (N_6982,N_6649,N_6256);
or U6983 (N_6983,N_6832,N_6734);
nor U6984 (N_6984,N_6782,N_6774);
and U6985 (N_6985,N_6776,N_6744);
nor U6986 (N_6986,N_6772,N_6871);
or U6987 (N_6987,N_6392,N_6585);
nand U6988 (N_6988,N_6374,N_6579);
or U6989 (N_6989,N_6347,N_6691);
nand U6990 (N_6990,N_6586,N_6817);
nand U6991 (N_6991,N_6359,N_6519);
or U6992 (N_6992,N_6340,N_6545);
and U6993 (N_6993,N_6376,N_6512);
xor U6994 (N_6994,N_6826,N_6682);
or U6995 (N_6995,N_6408,N_6665);
nand U6996 (N_6996,N_6781,N_6342);
nand U6997 (N_6997,N_6827,N_6815);
nand U6998 (N_6998,N_6501,N_6443);
or U6999 (N_6999,N_6323,N_6856);
nand U7000 (N_7000,N_6650,N_6345);
nor U7001 (N_7001,N_6281,N_6565);
and U7002 (N_7002,N_6267,N_6500);
nor U7003 (N_7003,N_6403,N_6449);
nand U7004 (N_7004,N_6821,N_6439);
or U7005 (N_7005,N_6260,N_6265);
nand U7006 (N_7006,N_6427,N_6822);
xor U7007 (N_7007,N_6254,N_6464);
nor U7008 (N_7008,N_6637,N_6846);
and U7009 (N_7009,N_6760,N_6543);
and U7010 (N_7010,N_6733,N_6492);
nor U7011 (N_7011,N_6809,N_6757);
or U7012 (N_7012,N_6642,N_6349);
nor U7013 (N_7013,N_6334,N_6393);
nand U7014 (N_7014,N_6448,N_6566);
or U7015 (N_7015,N_6547,N_6455);
and U7016 (N_7016,N_6341,N_6613);
or U7017 (N_7017,N_6704,N_6604);
xor U7018 (N_7018,N_6268,N_6434);
or U7019 (N_7019,N_6400,N_6758);
and U7020 (N_7020,N_6746,N_6489);
nand U7021 (N_7021,N_6369,N_6367);
nor U7022 (N_7022,N_6276,N_6841);
nor U7023 (N_7023,N_6402,N_6335);
nor U7024 (N_7024,N_6635,N_6258);
nand U7025 (N_7025,N_6379,N_6701);
and U7026 (N_7026,N_6546,N_6271);
or U7027 (N_7027,N_6568,N_6513);
nand U7028 (N_7028,N_6718,N_6773);
nor U7029 (N_7029,N_6771,N_6737);
and U7030 (N_7030,N_6275,N_6791);
nor U7031 (N_7031,N_6715,N_6296);
or U7032 (N_7032,N_6618,N_6283);
or U7033 (N_7033,N_6399,N_6725);
nand U7034 (N_7034,N_6686,N_6445);
and U7035 (N_7035,N_6633,N_6406);
or U7036 (N_7036,N_6272,N_6331);
or U7037 (N_7037,N_6671,N_6750);
or U7038 (N_7038,N_6532,N_6529);
nand U7039 (N_7039,N_6742,N_6428);
nand U7040 (N_7040,N_6785,N_6675);
nor U7041 (N_7041,N_6847,N_6727);
or U7042 (N_7042,N_6329,N_6654);
and U7043 (N_7043,N_6625,N_6722);
nand U7044 (N_7044,N_6555,N_6870);
and U7045 (N_7045,N_6861,N_6867);
and U7046 (N_7046,N_6837,N_6643);
and U7047 (N_7047,N_6667,N_6355);
nor U7048 (N_7048,N_6518,N_6496);
nand U7049 (N_7049,N_6607,N_6641);
xor U7050 (N_7050,N_6611,N_6648);
xnor U7051 (N_7051,N_6714,N_6511);
nand U7052 (N_7052,N_6690,N_6658);
or U7053 (N_7053,N_6731,N_6288);
or U7054 (N_7054,N_6616,N_6251);
or U7055 (N_7055,N_6663,N_6560);
or U7056 (N_7056,N_6630,N_6515);
and U7057 (N_7057,N_6514,N_6573);
and U7058 (N_7058,N_6711,N_6346);
nor U7059 (N_7059,N_6365,N_6554);
and U7060 (N_7060,N_6582,N_6700);
nor U7061 (N_7061,N_6753,N_6839);
xor U7062 (N_7062,N_6687,N_6471);
nor U7063 (N_7063,N_6597,N_6312);
xor U7064 (N_7064,N_6487,N_6632);
nor U7065 (N_7065,N_6255,N_6336);
or U7066 (N_7066,N_6820,N_6313);
and U7067 (N_7067,N_6670,N_6505);
xor U7068 (N_7068,N_6343,N_6446);
xnor U7069 (N_7069,N_6257,N_6452);
or U7070 (N_7070,N_6557,N_6311);
or U7071 (N_7071,N_6797,N_6584);
nand U7072 (N_7072,N_6274,N_6739);
nand U7073 (N_7073,N_6539,N_6488);
xnor U7074 (N_7074,N_6304,N_6269);
nor U7075 (N_7075,N_6549,N_6378);
or U7076 (N_7076,N_6401,N_6592);
nor U7077 (N_7077,N_6316,N_6803);
nor U7078 (N_7078,N_6266,N_6315);
or U7079 (N_7079,N_6698,N_6430);
or U7080 (N_7080,N_6777,N_6321);
or U7081 (N_7081,N_6534,N_6298);
nand U7082 (N_7082,N_6495,N_6852);
and U7083 (N_7083,N_6804,N_6780);
nor U7084 (N_7084,N_6451,N_6569);
xor U7085 (N_7085,N_6357,N_6745);
and U7086 (N_7086,N_6614,N_6531);
or U7087 (N_7087,N_6831,N_6646);
and U7088 (N_7088,N_6468,N_6491);
or U7089 (N_7089,N_6793,N_6736);
or U7090 (N_7090,N_6869,N_6339);
nor U7091 (N_7091,N_6290,N_6533);
or U7092 (N_7092,N_6289,N_6578);
nor U7093 (N_7093,N_6808,N_6303);
and U7094 (N_7094,N_6590,N_6818);
nand U7095 (N_7095,N_6328,N_6416);
and U7096 (N_7096,N_6583,N_6252);
nor U7097 (N_7097,N_6672,N_6470);
and U7098 (N_7098,N_6747,N_6396);
nor U7099 (N_7099,N_6706,N_6623);
xor U7100 (N_7100,N_6828,N_6509);
or U7101 (N_7101,N_6440,N_6273);
nor U7102 (N_7102,N_6493,N_6360);
and U7103 (N_7103,N_6498,N_6807);
nor U7104 (N_7104,N_6480,N_6844);
or U7105 (N_7105,N_6305,N_6638);
and U7106 (N_7106,N_6460,N_6420);
nor U7107 (N_7107,N_6653,N_6754);
nor U7108 (N_7108,N_6525,N_6864);
nor U7109 (N_7109,N_6795,N_6333);
or U7110 (N_7110,N_6263,N_6517);
nor U7111 (N_7111,N_6287,N_6829);
nand U7112 (N_7112,N_6719,N_6469);
nor U7113 (N_7113,N_6748,N_6277);
nand U7114 (N_7114,N_6617,N_6564);
nor U7115 (N_7115,N_6612,N_6830);
and U7116 (N_7116,N_6865,N_6789);
or U7117 (N_7117,N_6537,N_6295);
or U7118 (N_7118,N_6681,N_6694);
or U7119 (N_7119,N_6571,N_6507);
nor U7120 (N_7120,N_6389,N_6520);
or U7121 (N_7121,N_6552,N_6873);
and U7122 (N_7122,N_6692,N_6576);
and U7123 (N_7123,N_6792,N_6863);
and U7124 (N_7124,N_6410,N_6350);
or U7125 (N_7125,N_6766,N_6418);
nand U7126 (N_7126,N_6660,N_6353);
nand U7127 (N_7127,N_6447,N_6259);
nor U7128 (N_7128,N_6574,N_6409);
and U7129 (N_7129,N_6769,N_6595);
and U7130 (N_7130,N_6853,N_6503);
and U7131 (N_7131,N_6666,N_6326);
nand U7132 (N_7132,N_6530,N_6570);
xnor U7133 (N_7133,N_6802,N_6356);
or U7134 (N_7134,N_6645,N_6438);
nor U7135 (N_7135,N_6508,N_6415);
nand U7136 (N_7136,N_6655,N_6419);
or U7137 (N_7137,N_6394,N_6306);
xnor U7138 (N_7138,N_6709,N_6322);
nand U7139 (N_7139,N_6358,N_6696);
and U7140 (N_7140,N_6735,N_6652);
nor U7141 (N_7141,N_6253,N_6324);
or U7142 (N_7142,N_6453,N_6327);
nand U7143 (N_7143,N_6738,N_6300);
nand U7144 (N_7144,N_6310,N_6688);
nor U7145 (N_7145,N_6567,N_6278);
or U7146 (N_7146,N_6721,N_6859);
nand U7147 (N_7147,N_6366,N_6319);
or U7148 (N_7148,N_6494,N_6572);
or U7149 (N_7149,N_6397,N_6713);
and U7150 (N_7150,N_6835,N_6542);
nand U7151 (N_7151,N_6621,N_6435);
and U7152 (N_7152,N_6561,N_6368);
nor U7153 (N_7153,N_6767,N_6390);
nor U7154 (N_7154,N_6763,N_6751);
or U7155 (N_7155,N_6380,N_6622);
nand U7156 (N_7156,N_6707,N_6857);
nor U7157 (N_7157,N_6307,N_6426);
nor U7158 (N_7158,N_6432,N_6499);
and U7159 (N_7159,N_6659,N_6647);
nor U7160 (N_7160,N_6351,N_6723);
nor U7161 (N_7161,N_6693,N_6755);
and U7162 (N_7162,N_6814,N_6770);
and U7163 (N_7163,N_6644,N_6699);
and U7164 (N_7164,N_6454,N_6354);
nand U7165 (N_7165,N_6631,N_6282);
and U7166 (N_7166,N_6481,N_6775);
or U7167 (N_7167,N_6668,N_6309);
nand U7168 (N_7168,N_6485,N_6836);
and U7169 (N_7169,N_6798,N_6708);
xor U7170 (N_7170,N_6388,N_6677);
or U7171 (N_7171,N_6594,N_6845);
and U7172 (N_7172,N_6279,N_6474);
or U7173 (N_7173,N_6325,N_6575);
nor U7174 (N_7174,N_6264,N_6669);
or U7175 (N_7175,N_6527,N_6634);
or U7176 (N_7176,N_6318,N_6589);
or U7177 (N_7177,N_6656,N_6778);
nor U7178 (N_7178,N_6521,N_6563);
and U7179 (N_7179,N_6526,N_6610);
nand U7180 (N_7180,N_6352,N_6732);
xor U7181 (N_7181,N_6538,N_6740);
nand U7182 (N_7182,N_6787,N_6674);
and U7183 (N_7183,N_6386,N_6332);
or U7184 (N_7184,N_6702,N_6490);
and U7185 (N_7185,N_6459,N_6862);
nand U7186 (N_7186,N_6524,N_6548);
nor U7187 (N_7187,N_6606,N_6572);
and U7188 (N_7188,N_6564,N_6575);
or U7189 (N_7189,N_6831,N_6632);
or U7190 (N_7190,N_6416,N_6713);
xnor U7191 (N_7191,N_6540,N_6482);
and U7192 (N_7192,N_6342,N_6474);
nor U7193 (N_7193,N_6680,N_6262);
and U7194 (N_7194,N_6515,N_6455);
nand U7195 (N_7195,N_6586,N_6396);
nor U7196 (N_7196,N_6282,N_6337);
nand U7197 (N_7197,N_6859,N_6694);
nor U7198 (N_7198,N_6650,N_6492);
nor U7199 (N_7199,N_6469,N_6413);
nor U7200 (N_7200,N_6276,N_6482);
and U7201 (N_7201,N_6340,N_6643);
and U7202 (N_7202,N_6870,N_6342);
nor U7203 (N_7203,N_6722,N_6501);
or U7204 (N_7204,N_6451,N_6701);
nand U7205 (N_7205,N_6862,N_6572);
or U7206 (N_7206,N_6798,N_6874);
nor U7207 (N_7207,N_6633,N_6287);
and U7208 (N_7208,N_6765,N_6405);
nand U7209 (N_7209,N_6311,N_6709);
and U7210 (N_7210,N_6733,N_6299);
or U7211 (N_7211,N_6404,N_6554);
xnor U7212 (N_7212,N_6572,N_6701);
and U7213 (N_7213,N_6366,N_6503);
nand U7214 (N_7214,N_6444,N_6375);
nand U7215 (N_7215,N_6497,N_6354);
nand U7216 (N_7216,N_6253,N_6659);
or U7217 (N_7217,N_6512,N_6702);
or U7218 (N_7218,N_6308,N_6803);
nor U7219 (N_7219,N_6375,N_6340);
xor U7220 (N_7220,N_6722,N_6700);
nand U7221 (N_7221,N_6461,N_6842);
xor U7222 (N_7222,N_6438,N_6774);
nand U7223 (N_7223,N_6332,N_6785);
nand U7224 (N_7224,N_6416,N_6283);
and U7225 (N_7225,N_6323,N_6397);
and U7226 (N_7226,N_6400,N_6297);
xnor U7227 (N_7227,N_6603,N_6646);
nor U7228 (N_7228,N_6615,N_6396);
xor U7229 (N_7229,N_6435,N_6678);
or U7230 (N_7230,N_6714,N_6662);
and U7231 (N_7231,N_6615,N_6456);
nand U7232 (N_7232,N_6410,N_6464);
or U7233 (N_7233,N_6785,N_6493);
or U7234 (N_7234,N_6564,N_6673);
or U7235 (N_7235,N_6478,N_6315);
or U7236 (N_7236,N_6526,N_6331);
nand U7237 (N_7237,N_6305,N_6552);
and U7238 (N_7238,N_6270,N_6274);
nand U7239 (N_7239,N_6805,N_6645);
and U7240 (N_7240,N_6356,N_6294);
or U7241 (N_7241,N_6520,N_6482);
and U7242 (N_7242,N_6632,N_6492);
and U7243 (N_7243,N_6533,N_6849);
nor U7244 (N_7244,N_6860,N_6464);
nor U7245 (N_7245,N_6322,N_6263);
nor U7246 (N_7246,N_6718,N_6363);
or U7247 (N_7247,N_6706,N_6518);
and U7248 (N_7248,N_6343,N_6768);
and U7249 (N_7249,N_6762,N_6393);
nand U7250 (N_7250,N_6703,N_6679);
or U7251 (N_7251,N_6416,N_6590);
xnor U7252 (N_7252,N_6763,N_6554);
or U7253 (N_7253,N_6705,N_6560);
nand U7254 (N_7254,N_6667,N_6579);
nand U7255 (N_7255,N_6262,N_6765);
nor U7256 (N_7256,N_6493,N_6255);
nand U7257 (N_7257,N_6284,N_6535);
or U7258 (N_7258,N_6740,N_6806);
nand U7259 (N_7259,N_6573,N_6305);
and U7260 (N_7260,N_6362,N_6593);
and U7261 (N_7261,N_6279,N_6320);
nand U7262 (N_7262,N_6857,N_6432);
nor U7263 (N_7263,N_6624,N_6668);
and U7264 (N_7264,N_6364,N_6801);
nor U7265 (N_7265,N_6312,N_6685);
or U7266 (N_7266,N_6586,N_6642);
and U7267 (N_7267,N_6338,N_6483);
nand U7268 (N_7268,N_6585,N_6501);
or U7269 (N_7269,N_6551,N_6873);
or U7270 (N_7270,N_6635,N_6774);
or U7271 (N_7271,N_6869,N_6680);
or U7272 (N_7272,N_6563,N_6537);
nor U7273 (N_7273,N_6475,N_6304);
nor U7274 (N_7274,N_6324,N_6474);
nor U7275 (N_7275,N_6465,N_6369);
nor U7276 (N_7276,N_6764,N_6830);
nand U7277 (N_7277,N_6447,N_6251);
xor U7278 (N_7278,N_6719,N_6785);
nand U7279 (N_7279,N_6350,N_6481);
and U7280 (N_7280,N_6414,N_6768);
nand U7281 (N_7281,N_6270,N_6587);
and U7282 (N_7282,N_6354,N_6343);
xor U7283 (N_7283,N_6282,N_6470);
nor U7284 (N_7284,N_6599,N_6697);
nand U7285 (N_7285,N_6332,N_6615);
and U7286 (N_7286,N_6391,N_6344);
and U7287 (N_7287,N_6537,N_6477);
or U7288 (N_7288,N_6514,N_6589);
nand U7289 (N_7289,N_6606,N_6355);
and U7290 (N_7290,N_6415,N_6466);
and U7291 (N_7291,N_6357,N_6702);
or U7292 (N_7292,N_6856,N_6769);
nand U7293 (N_7293,N_6787,N_6598);
and U7294 (N_7294,N_6684,N_6812);
or U7295 (N_7295,N_6591,N_6257);
nand U7296 (N_7296,N_6662,N_6438);
and U7297 (N_7297,N_6493,N_6782);
nand U7298 (N_7298,N_6460,N_6401);
nor U7299 (N_7299,N_6839,N_6349);
nor U7300 (N_7300,N_6676,N_6320);
nand U7301 (N_7301,N_6402,N_6844);
or U7302 (N_7302,N_6327,N_6344);
nand U7303 (N_7303,N_6529,N_6509);
and U7304 (N_7304,N_6846,N_6625);
xor U7305 (N_7305,N_6426,N_6689);
xnor U7306 (N_7306,N_6362,N_6361);
and U7307 (N_7307,N_6536,N_6645);
nor U7308 (N_7308,N_6629,N_6577);
or U7309 (N_7309,N_6731,N_6754);
or U7310 (N_7310,N_6435,N_6843);
nand U7311 (N_7311,N_6528,N_6863);
and U7312 (N_7312,N_6846,N_6482);
and U7313 (N_7313,N_6507,N_6293);
nand U7314 (N_7314,N_6639,N_6258);
nand U7315 (N_7315,N_6283,N_6257);
and U7316 (N_7316,N_6615,N_6535);
and U7317 (N_7317,N_6546,N_6286);
or U7318 (N_7318,N_6844,N_6436);
and U7319 (N_7319,N_6809,N_6694);
nor U7320 (N_7320,N_6804,N_6326);
and U7321 (N_7321,N_6750,N_6431);
and U7322 (N_7322,N_6270,N_6741);
and U7323 (N_7323,N_6336,N_6765);
and U7324 (N_7324,N_6451,N_6756);
nand U7325 (N_7325,N_6574,N_6491);
nor U7326 (N_7326,N_6691,N_6665);
nor U7327 (N_7327,N_6665,N_6378);
and U7328 (N_7328,N_6773,N_6820);
nand U7329 (N_7329,N_6463,N_6501);
and U7330 (N_7330,N_6735,N_6719);
or U7331 (N_7331,N_6767,N_6474);
and U7332 (N_7332,N_6362,N_6755);
and U7333 (N_7333,N_6665,N_6812);
nor U7334 (N_7334,N_6257,N_6763);
and U7335 (N_7335,N_6544,N_6585);
or U7336 (N_7336,N_6429,N_6829);
and U7337 (N_7337,N_6258,N_6728);
nor U7338 (N_7338,N_6838,N_6685);
nand U7339 (N_7339,N_6620,N_6636);
and U7340 (N_7340,N_6272,N_6801);
nand U7341 (N_7341,N_6814,N_6546);
nor U7342 (N_7342,N_6730,N_6724);
nor U7343 (N_7343,N_6556,N_6784);
nand U7344 (N_7344,N_6479,N_6258);
nor U7345 (N_7345,N_6313,N_6372);
or U7346 (N_7346,N_6404,N_6541);
or U7347 (N_7347,N_6323,N_6410);
and U7348 (N_7348,N_6808,N_6335);
and U7349 (N_7349,N_6403,N_6769);
or U7350 (N_7350,N_6675,N_6787);
and U7351 (N_7351,N_6493,N_6721);
nor U7352 (N_7352,N_6497,N_6464);
and U7353 (N_7353,N_6432,N_6508);
or U7354 (N_7354,N_6484,N_6632);
and U7355 (N_7355,N_6424,N_6273);
nand U7356 (N_7356,N_6630,N_6270);
nand U7357 (N_7357,N_6575,N_6338);
nand U7358 (N_7358,N_6734,N_6662);
and U7359 (N_7359,N_6255,N_6861);
nor U7360 (N_7360,N_6871,N_6689);
and U7361 (N_7361,N_6297,N_6363);
and U7362 (N_7362,N_6873,N_6496);
nor U7363 (N_7363,N_6312,N_6788);
xnor U7364 (N_7364,N_6308,N_6333);
nand U7365 (N_7365,N_6849,N_6502);
and U7366 (N_7366,N_6734,N_6810);
xnor U7367 (N_7367,N_6424,N_6760);
nor U7368 (N_7368,N_6839,N_6629);
and U7369 (N_7369,N_6470,N_6392);
nand U7370 (N_7370,N_6544,N_6286);
or U7371 (N_7371,N_6756,N_6393);
and U7372 (N_7372,N_6542,N_6848);
or U7373 (N_7373,N_6567,N_6515);
nand U7374 (N_7374,N_6770,N_6727);
xnor U7375 (N_7375,N_6820,N_6398);
nor U7376 (N_7376,N_6564,N_6672);
xnor U7377 (N_7377,N_6591,N_6575);
and U7378 (N_7378,N_6857,N_6751);
and U7379 (N_7379,N_6668,N_6416);
or U7380 (N_7380,N_6858,N_6376);
xor U7381 (N_7381,N_6870,N_6357);
and U7382 (N_7382,N_6288,N_6806);
and U7383 (N_7383,N_6261,N_6647);
and U7384 (N_7384,N_6718,N_6612);
or U7385 (N_7385,N_6706,N_6537);
xor U7386 (N_7386,N_6731,N_6561);
or U7387 (N_7387,N_6567,N_6423);
xnor U7388 (N_7388,N_6436,N_6425);
nand U7389 (N_7389,N_6513,N_6350);
nor U7390 (N_7390,N_6348,N_6522);
nand U7391 (N_7391,N_6859,N_6375);
xor U7392 (N_7392,N_6466,N_6782);
or U7393 (N_7393,N_6456,N_6380);
or U7394 (N_7394,N_6725,N_6694);
and U7395 (N_7395,N_6640,N_6567);
and U7396 (N_7396,N_6607,N_6721);
or U7397 (N_7397,N_6532,N_6333);
xnor U7398 (N_7398,N_6723,N_6718);
and U7399 (N_7399,N_6874,N_6543);
and U7400 (N_7400,N_6761,N_6815);
and U7401 (N_7401,N_6505,N_6653);
and U7402 (N_7402,N_6350,N_6401);
nor U7403 (N_7403,N_6424,N_6835);
nor U7404 (N_7404,N_6570,N_6302);
or U7405 (N_7405,N_6383,N_6346);
or U7406 (N_7406,N_6276,N_6772);
or U7407 (N_7407,N_6371,N_6574);
xor U7408 (N_7408,N_6864,N_6482);
xnor U7409 (N_7409,N_6355,N_6671);
and U7410 (N_7410,N_6313,N_6291);
nor U7411 (N_7411,N_6417,N_6778);
or U7412 (N_7412,N_6419,N_6322);
nor U7413 (N_7413,N_6827,N_6586);
or U7414 (N_7414,N_6297,N_6842);
xor U7415 (N_7415,N_6710,N_6507);
and U7416 (N_7416,N_6452,N_6555);
nor U7417 (N_7417,N_6718,N_6831);
and U7418 (N_7418,N_6602,N_6607);
and U7419 (N_7419,N_6417,N_6568);
nand U7420 (N_7420,N_6402,N_6606);
and U7421 (N_7421,N_6718,N_6293);
nand U7422 (N_7422,N_6273,N_6469);
nand U7423 (N_7423,N_6571,N_6825);
and U7424 (N_7424,N_6553,N_6856);
nand U7425 (N_7425,N_6870,N_6447);
or U7426 (N_7426,N_6365,N_6702);
nand U7427 (N_7427,N_6369,N_6355);
and U7428 (N_7428,N_6291,N_6826);
and U7429 (N_7429,N_6310,N_6465);
nand U7430 (N_7430,N_6591,N_6797);
and U7431 (N_7431,N_6374,N_6387);
and U7432 (N_7432,N_6298,N_6435);
or U7433 (N_7433,N_6805,N_6307);
and U7434 (N_7434,N_6462,N_6464);
or U7435 (N_7435,N_6736,N_6465);
nand U7436 (N_7436,N_6534,N_6632);
xor U7437 (N_7437,N_6708,N_6427);
and U7438 (N_7438,N_6659,N_6751);
nor U7439 (N_7439,N_6539,N_6532);
or U7440 (N_7440,N_6542,N_6429);
xor U7441 (N_7441,N_6560,N_6314);
and U7442 (N_7442,N_6601,N_6489);
nand U7443 (N_7443,N_6300,N_6530);
nand U7444 (N_7444,N_6393,N_6643);
and U7445 (N_7445,N_6365,N_6550);
nand U7446 (N_7446,N_6683,N_6554);
or U7447 (N_7447,N_6745,N_6818);
and U7448 (N_7448,N_6608,N_6553);
and U7449 (N_7449,N_6754,N_6347);
nor U7450 (N_7450,N_6563,N_6727);
and U7451 (N_7451,N_6659,N_6445);
and U7452 (N_7452,N_6395,N_6685);
and U7453 (N_7453,N_6545,N_6297);
and U7454 (N_7454,N_6636,N_6745);
or U7455 (N_7455,N_6845,N_6559);
and U7456 (N_7456,N_6629,N_6274);
or U7457 (N_7457,N_6678,N_6706);
or U7458 (N_7458,N_6433,N_6438);
nor U7459 (N_7459,N_6832,N_6272);
nand U7460 (N_7460,N_6712,N_6263);
or U7461 (N_7461,N_6650,N_6440);
or U7462 (N_7462,N_6638,N_6552);
nand U7463 (N_7463,N_6514,N_6731);
nand U7464 (N_7464,N_6690,N_6533);
nor U7465 (N_7465,N_6555,N_6466);
nand U7466 (N_7466,N_6563,N_6825);
nand U7467 (N_7467,N_6815,N_6331);
and U7468 (N_7468,N_6461,N_6689);
nand U7469 (N_7469,N_6388,N_6311);
xnor U7470 (N_7470,N_6577,N_6749);
and U7471 (N_7471,N_6651,N_6836);
and U7472 (N_7472,N_6661,N_6386);
nand U7473 (N_7473,N_6798,N_6619);
nand U7474 (N_7474,N_6391,N_6270);
and U7475 (N_7475,N_6346,N_6314);
and U7476 (N_7476,N_6806,N_6779);
nand U7477 (N_7477,N_6351,N_6301);
nand U7478 (N_7478,N_6555,N_6817);
or U7479 (N_7479,N_6589,N_6653);
or U7480 (N_7480,N_6369,N_6447);
nor U7481 (N_7481,N_6765,N_6686);
xnor U7482 (N_7482,N_6502,N_6733);
nand U7483 (N_7483,N_6428,N_6478);
or U7484 (N_7484,N_6835,N_6449);
or U7485 (N_7485,N_6752,N_6275);
nor U7486 (N_7486,N_6480,N_6395);
and U7487 (N_7487,N_6532,N_6686);
nor U7488 (N_7488,N_6808,N_6331);
nor U7489 (N_7489,N_6301,N_6735);
or U7490 (N_7490,N_6586,N_6629);
and U7491 (N_7491,N_6623,N_6452);
nor U7492 (N_7492,N_6349,N_6554);
or U7493 (N_7493,N_6303,N_6779);
or U7494 (N_7494,N_6395,N_6277);
or U7495 (N_7495,N_6762,N_6656);
or U7496 (N_7496,N_6363,N_6685);
nand U7497 (N_7497,N_6633,N_6300);
nand U7498 (N_7498,N_6749,N_6544);
nand U7499 (N_7499,N_6849,N_6473);
nor U7500 (N_7500,N_7485,N_6982);
nand U7501 (N_7501,N_7180,N_7320);
or U7502 (N_7502,N_6904,N_7307);
and U7503 (N_7503,N_7312,N_6993);
or U7504 (N_7504,N_7228,N_7185);
or U7505 (N_7505,N_6910,N_7483);
xnor U7506 (N_7506,N_7166,N_7018);
xnor U7507 (N_7507,N_6915,N_7126);
or U7508 (N_7508,N_7222,N_7326);
nand U7509 (N_7509,N_7127,N_6983);
and U7510 (N_7510,N_7002,N_6940);
nor U7511 (N_7511,N_7152,N_7082);
nand U7512 (N_7512,N_7003,N_7074);
and U7513 (N_7513,N_7278,N_7284);
and U7514 (N_7514,N_7100,N_7240);
xnor U7515 (N_7515,N_6912,N_7035);
nor U7516 (N_7516,N_7120,N_6970);
xor U7517 (N_7517,N_7430,N_7044);
or U7518 (N_7518,N_7433,N_7224);
and U7519 (N_7519,N_7087,N_7201);
nand U7520 (N_7520,N_7477,N_7131);
or U7521 (N_7521,N_7019,N_7210);
nor U7522 (N_7522,N_6890,N_7269);
nor U7523 (N_7523,N_7410,N_7025);
or U7524 (N_7524,N_7114,N_7459);
and U7525 (N_7525,N_7155,N_7254);
xnor U7526 (N_7526,N_7488,N_7253);
or U7527 (N_7527,N_7340,N_7496);
nand U7528 (N_7528,N_7069,N_6901);
or U7529 (N_7529,N_7215,N_7187);
or U7530 (N_7530,N_7072,N_7470);
or U7531 (N_7531,N_7255,N_7064);
xor U7532 (N_7532,N_6922,N_7411);
nand U7533 (N_7533,N_7271,N_7144);
or U7534 (N_7534,N_7342,N_6885);
nor U7535 (N_7535,N_7277,N_7175);
nor U7536 (N_7536,N_7321,N_7250);
xnor U7537 (N_7537,N_7373,N_6897);
and U7538 (N_7538,N_7153,N_7227);
xnor U7539 (N_7539,N_7372,N_7379);
nor U7540 (N_7540,N_7252,N_7350);
and U7541 (N_7541,N_7089,N_7456);
or U7542 (N_7542,N_7160,N_7409);
or U7543 (N_7543,N_7355,N_6880);
or U7544 (N_7544,N_7418,N_7038);
and U7545 (N_7545,N_7095,N_7335);
nand U7546 (N_7546,N_6989,N_7093);
and U7547 (N_7547,N_7280,N_6877);
nor U7548 (N_7548,N_7371,N_7233);
xor U7549 (N_7549,N_7241,N_7398);
nor U7550 (N_7550,N_6974,N_6914);
and U7551 (N_7551,N_7157,N_7036);
nor U7552 (N_7552,N_7384,N_7472);
nand U7553 (N_7553,N_6956,N_7107);
and U7554 (N_7554,N_7380,N_7286);
nand U7555 (N_7555,N_7086,N_7084);
nand U7556 (N_7556,N_6876,N_7042);
nand U7557 (N_7557,N_7282,N_7295);
and U7558 (N_7558,N_7464,N_7015);
nor U7559 (N_7559,N_6945,N_6881);
and U7560 (N_7560,N_6991,N_7260);
and U7561 (N_7561,N_7060,N_7300);
nor U7562 (N_7562,N_7426,N_7165);
and U7563 (N_7563,N_6959,N_6952);
and U7564 (N_7564,N_7369,N_7494);
nand U7565 (N_7565,N_7226,N_7112);
and U7566 (N_7566,N_7143,N_6967);
nor U7567 (N_7567,N_7231,N_6977);
or U7568 (N_7568,N_7119,N_7193);
or U7569 (N_7569,N_6903,N_7246);
and U7570 (N_7570,N_7251,N_6900);
nand U7571 (N_7571,N_7493,N_7479);
and U7572 (N_7572,N_7048,N_6990);
nand U7573 (N_7573,N_7396,N_7129);
and U7574 (N_7574,N_6939,N_7465);
and U7575 (N_7575,N_6963,N_7487);
or U7576 (N_7576,N_6960,N_7158);
or U7577 (N_7577,N_7417,N_7004);
or U7578 (N_7578,N_7329,N_7293);
nor U7579 (N_7579,N_7005,N_7471);
nand U7580 (N_7580,N_7162,N_7336);
nand U7581 (N_7581,N_7442,N_7415);
or U7582 (N_7582,N_7151,N_7367);
or U7583 (N_7583,N_7317,N_7128);
and U7584 (N_7584,N_7274,N_6978);
and U7585 (N_7585,N_7068,N_6971);
nand U7586 (N_7586,N_7366,N_7059);
and U7587 (N_7587,N_7209,N_7484);
or U7588 (N_7588,N_7429,N_7237);
nor U7589 (N_7589,N_7202,N_7383);
and U7590 (N_7590,N_6932,N_7436);
nor U7591 (N_7591,N_7285,N_6917);
or U7592 (N_7592,N_6919,N_7098);
nor U7593 (N_7593,N_7462,N_7109);
nor U7594 (N_7594,N_7046,N_6955);
and U7595 (N_7595,N_7186,N_7414);
xor U7596 (N_7596,N_7049,N_6961);
nor U7597 (N_7597,N_7101,N_7106);
or U7598 (N_7598,N_7424,N_7195);
nor U7599 (N_7599,N_7281,N_7198);
or U7600 (N_7600,N_7039,N_7123);
or U7601 (N_7601,N_7290,N_7389);
xnor U7602 (N_7602,N_7110,N_7408);
nor U7603 (N_7603,N_7376,N_7316);
nor U7604 (N_7604,N_7267,N_7359);
nand U7605 (N_7605,N_7451,N_7040);
xnor U7606 (N_7606,N_6891,N_7217);
and U7607 (N_7607,N_7348,N_7090);
or U7608 (N_7608,N_7346,N_7352);
nand U7609 (N_7609,N_7136,N_7268);
nor U7610 (N_7610,N_7275,N_7022);
or U7611 (N_7611,N_6921,N_7322);
and U7612 (N_7612,N_6925,N_7169);
and U7613 (N_7613,N_7297,N_7247);
or U7614 (N_7614,N_7422,N_7183);
nor U7615 (N_7615,N_7023,N_6913);
and U7616 (N_7616,N_7301,N_7117);
nand U7617 (N_7617,N_7481,N_7279);
nor U7618 (N_7618,N_7272,N_7388);
xnor U7619 (N_7619,N_6966,N_7363);
and U7620 (N_7620,N_7216,N_7306);
nand U7621 (N_7621,N_7154,N_7475);
nor U7622 (N_7622,N_7343,N_7212);
nand U7623 (N_7623,N_7052,N_7296);
nand U7624 (N_7624,N_7146,N_7031);
nand U7625 (N_7625,N_6948,N_7145);
and U7626 (N_7626,N_7189,N_6894);
nor U7627 (N_7627,N_6975,N_6949);
or U7628 (N_7628,N_7276,N_7181);
or U7629 (N_7629,N_7299,N_7016);
and U7630 (N_7630,N_7079,N_7498);
and U7631 (N_7631,N_6947,N_6965);
and U7632 (N_7632,N_7490,N_7478);
xnor U7633 (N_7633,N_7310,N_7103);
or U7634 (N_7634,N_7011,N_6893);
and U7635 (N_7635,N_7242,N_7370);
or U7636 (N_7636,N_7291,N_7327);
xnor U7637 (N_7637,N_7314,N_7446);
nor U7638 (N_7638,N_7287,N_7402);
nor U7639 (N_7639,N_6937,N_7261);
or U7640 (N_7640,N_7243,N_7266);
nor U7641 (N_7641,N_7262,N_7497);
nor U7642 (N_7642,N_7037,N_6957);
or U7643 (N_7643,N_7124,N_7063);
nor U7644 (N_7644,N_7263,N_6927);
and U7645 (N_7645,N_7458,N_6995);
nor U7646 (N_7646,N_7358,N_7425);
and U7647 (N_7647,N_7096,N_6968);
or U7648 (N_7648,N_7132,N_7309);
nand U7649 (N_7649,N_7244,N_6933);
nand U7650 (N_7650,N_6899,N_7164);
nor U7651 (N_7651,N_7029,N_6988);
nand U7652 (N_7652,N_7220,N_7403);
xor U7653 (N_7653,N_7303,N_7334);
nor U7654 (N_7654,N_6918,N_7000);
nand U7655 (N_7655,N_7194,N_7413);
or U7656 (N_7656,N_7214,N_6984);
or U7657 (N_7657,N_7159,N_7245);
nand U7658 (N_7658,N_7491,N_6994);
or U7659 (N_7659,N_6979,N_7174);
xnor U7660 (N_7660,N_7331,N_7199);
nor U7661 (N_7661,N_7184,N_7001);
xor U7662 (N_7662,N_7140,N_6907);
or U7663 (N_7663,N_7034,N_7088);
or U7664 (N_7664,N_7450,N_7339);
nand U7665 (N_7665,N_7156,N_6908);
or U7666 (N_7666,N_7030,N_7196);
or U7667 (N_7667,N_6882,N_6911);
xor U7668 (N_7668,N_7078,N_7139);
or U7669 (N_7669,N_7273,N_7292);
nor U7670 (N_7670,N_7289,N_6906);
and U7671 (N_7671,N_7454,N_7476);
or U7672 (N_7672,N_7420,N_6930);
or U7673 (N_7673,N_6972,N_7283);
or U7674 (N_7674,N_7486,N_7391);
xnor U7675 (N_7675,N_6936,N_7365);
nor U7676 (N_7676,N_7221,N_7407);
or U7677 (N_7677,N_6944,N_6875);
nand U7678 (N_7678,N_7105,N_7288);
and U7679 (N_7679,N_7377,N_7197);
nand U7680 (N_7680,N_7024,N_7045);
nor U7681 (N_7681,N_7097,N_7027);
nor U7682 (N_7682,N_7211,N_7073);
or U7683 (N_7683,N_7259,N_6964);
or U7684 (N_7684,N_7473,N_7457);
or U7685 (N_7685,N_7188,N_7173);
or U7686 (N_7686,N_6909,N_7033);
nand U7687 (N_7687,N_7364,N_7028);
nand U7688 (N_7688,N_6996,N_7091);
nor U7689 (N_7689,N_7161,N_7405);
nand U7690 (N_7690,N_7007,N_6999);
or U7691 (N_7691,N_7360,N_6958);
xnor U7692 (N_7692,N_7444,N_6943);
and U7693 (N_7693,N_7179,N_7449);
and U7694 (N_7694,N_7330,N_7431);
or U7695 (N_7695,N_6969,N_7323);
nand U7696 (N_7696,N_7495,N_7492);
or U7697 (N_7697,N_7204,N_6892);
and U7698 (N_7698,N_6883,N_7499);
or U7699 (N_7699,N_7111,N_7115);
xnor U7700 (N_7700,N_7337,N_7135);
and U7701 (N_7701,N_7239,N_6986);
nor U7702 (N_7702,N_7225,N_7397);
xor U7703 (N_7703,N_7219,N_6992);
and U7704 (N_7704,N_7230,N_7341);
nor U7705 (N_7705,N_6987,N_7445);
or U7706 (N_7706,N_7077,N_6985);
or U7707 (N_7707,N_7257,N_6934);
nor U7708 (N_7708,N_7235,N_7466);
nand U7709 (N_7709,N_7177,N_7270);
or U7710 (N_7710,N_7167,N_7248);
and U7711 (N_7711,N_7311,N_6942);
nor U7712 (N_7712,N_7094,N_7176);
nor U7713 (N_7713,N_7182,N_7264);
nand U7714 (N_7714,N_7054,N_7149);
or U7715 (N_7715,N_7349,N_7113);
and U7716 (N_7716,N_6950,N_7192);
or U7717 (N_7717,N_7050,N_7053);
and U7718 (N_7718,N_7385,N_7432);
nor U7719 (N_7719,N_7351,N_7421);
xnor U7720 (N_7720,N_6973,N_7134);
and U7721 (N_7721,N_7387,N_7062);
xor U7722 (N_7722,N_7441,N_7354);
and U7723 (N_7723,N_7067,N_7137);
xnor U7724 (N_7724,N_7386,N_7315);
nor U7725 (N_7725,N_7116,N_7147);
or U7726 (N_7726,N_7463,N_7308);
nand U7727 (N_7727,N_7006,N_7047);
nor U7728 (N_7728,N_7448,N_6896);
or U7729 (N_7729,N_7265,N_7313);
nor U7730 (N_7730,N_7428,N_7338);
nor U7731 (N_7731,N_7447,N_7014);
or U7732 (N_7732,N_7453,N_7333);
nor U7733 (N_7733,N_7443,N_7170);
and U7734 (N_7734,N_6884,N_7452);
nand U7735 (N_7735,N_7190,N_7208);
nor U7736 (N_7736,N_7344,N_6935);
and U7737 (N_7737,N_7401,N_6886);
or U7738 (N_7738,N_7083,N_7394);
or U7739 (N_7739,N_7085,N_7423);
nand U7740 (N_7740,N_7071,N_6887);
or U7741 (N_7741,N_7319,N_7104);
nand U7742 (N_7742,N_7395,N_7325);
nand U7743 (N_7743,N_7375,N_7399);
nand U7744 (N_7744,N_7076,N_7178);
and U7745 (N_7745,N_7455,N_7070);
nand U7746 (N_7746,N_6926,N_7480);
nand U7747 (N_7747,N_6981,N_7168);
nand U7748 (N_7748,N_7468,N_7361);
or U7749 (N_7749,N_7258,N_7055);
and U7750 (N_7750,N_7213,N_7304);
nand U7751 (N_7751,N_7440,N_6938);
xnor U7752 (N_7752,N_7345,N_7238);
nor U7753 (N_7753,N_7234,N_7150);
nor U7754 (N_7754,N_7061,N_7141);
and U7755 (N_7755,N_6924,N_7207);
or U7756 (N_7756,N_6946,N_7058);
xnor U7757 (N_7757,N_7256,N_6898);
nor U7758 (N_7758,N_7026,N_7368);
or U7759 (N_7759,N_7051,N_7013);
nor U7760 (N_7760,N_7482,N_7489);
and U7761 (N_7761,N_7294,N_7020);
or U7762 (N_7762,N_7066,N_6888);
or U7763 (N_7763,N_7324,N_6997);
nor U7764 (N_7764,N_7469,N_7118);
nand U7765 (N_7765,N_7008,N_7009);
or U7766 (N_7766,N_7249,N_7056);
and U7767 (N_7767,N_7434,N_6929);
or U7768 (N_7768,N_7416,N_6923);
or U7769 (N_7769,N_7017,N_7043);
or U7770 (N_7770,N_7438,N_7390);
and U7771 (N_7771,N_7353,N_7381);
nor U7772 (N_7772,N_6895,N_6878);
nand U7773 (N_7773,N_7302,N_6916);
nand U7774 (N_7774,N_7427,N_7171);
nor U7775 (N_7775,N_7400,N_7205);
nand U7776 (N_7776,N_7393,N_7437);
or U7777 (N_7777,N_7357,N_6951);
nand U7778 (N_7778,N_7138,N_7218);
and U7779 (N_7779,N_7080,N_7406);
nand U7780 (N_7780,N_7108,N_7148);
or U7781 (N_7781,N_7382,N_7460);
and U7782 (N_7782,N_7102,N_7057);
nand U7783 (N_7783,N_6980,N_6962);
nand U7784 (N_7784,N_7065,N_6902);
or U7785 (N_7785,N_7130,N_6889);
nand U7786 (N_7786,N_7474,N_7236);
nand U7787 (N_7787,N_7099,N_6928);
and U7788 (N_7788,N_6920,N_6879);
or U7789 (N_7789,N_7412,N_7461);
xnor U7790 (N_7790,N_7041,N_7200);
and U7791 (N_7791,N_6976,N_7125);
nand U7792 (N_7792,N_6998,N_6905);
nand U7793 (N_7793,N_7347,N_7010);
and U7794 (N_7794,N_7392,N_7229);
nor U7795 (N_7795,N_7203,N_7419);
nand U7796 (N_7796,N_7467,N_7012);
and U7797 (N_7797,N_7021,N_7172);
nand U7798 (N_7798,N_6941,N_7318);
or U7799 (N_7799,N_7206,N_7142);
nor U7800 (N_7800,N_7439,N_7223);
nor U7801 (N_7801,N_7298,N_7191);
nor U7802 (N_7802,N_7378,N_7122);
nand U7803 (N_7803,N_7374,N_7092);
and U7804 (N_7804,N_7435,N_7075);
xnor U7805 (N_7805,N_6931,N_7081);
nor U7806 (N_7806,N_7356,N_7404);
nand U7807 (N_7807,N_7032,N_7133);
nor U7808 (N_7808,N_7121,N_7305);
xnor U7809 (N_7809,N_7232,N_6954);
or U7810 (N_7810,N_7362,N_7328);
nor U7811 (N_7811,N_6953,N_7163);
nor U7812 (N_7812,N_7332,N_6990);
nand U7813 (N_7813,N_7033,N_7377);
nor U7814 (N_7814,N_7027,N_7481);
and U7815 (N_7815,N_7090,N_6984);
xor U7816 (N_7816,N_7138,N_7241);
and U7817 (N_7817,N_6966,N_7034);
or U7818 (N_7818,N_7067,N_7273);
nand U7819 (N_7819,N_7243,N_7121);
nand U7820 (N_7820,N_6932,N_6952);
and U7821 (N_7821,N_7243,N_7498);
or U7822 (N_7822,N_7124,N_7332);
nor U7823 (N_7823,N_7312,N_7478);
nand U7824 (N_7824,N_7198,N_6894);
and U7825 (N_7825,N_7124,N_6899);
and U7826 (N_7826,N_7390,N_7026);
or U7827 (N_7827,N_7272,N_6944);
nor U7828 (N_7828,N_7062,N_7336);
nor U7829 (N_7829,N_7153,N_7251);
and U7830 (N_7830,N_7184,N_7290);
nor U7831 (N_7831,N_7364,N_6974);
nand U7832 (N_7832,N_7480,N_7322);
xor U7833 (N_7833,N_7130,N_7381);
and U7834 (N_7834,N_7097,N_6920);
xor U7835 (N_7835,N_7275,N_6979);
nor U7836 (N_7836,N_7323,N_7044);
and U7837 (N_7837,N_7094,N_6883);
nor U7838 (N_7838,N_6931,N_7036);
nor U7839 (N_7839,N_7232,N_6962);
and U7840 (N_7840,N_6878,N_7396);
or U7841 (N_7841,N_7035,N_7372);
nand U7842 (N_7842,N_7399,N_7247);
nand U7843 (N_7843,N_7165,N_7139);
or U7844 (N_7844,N_7261,N_7288);
xor U7845 (N_7845,N_6968,N_7451);
nand U7846 (N_7846,N_7211,N_7403);
and U7847 (N_7847,N_7359,N_7277);
or U7848 (N_7848,N_7198,N_7103);
xor U7849 (N_7849,N_7408,N_7206);
nor U7850 (N_7850,N_7306,N_7146);
or U7851 (N_7851,N_7199,N_7349);
nor U7852 (N_7852,N_7482,N_7136);
or U7853 (N_7853,N_7050,N_6894);
and U7854 (N_7854,N_6994,N_7255);
or U7855 (N_7855,N_7050,N_6940);
and U7856 (N_7856,N_6875,N_6934);
nand U7857 (N_7857,N_7447,N_7024);
nor U7858 (N_7858,N_7260,N_7015);
and U7859 (N_7859,N_7076,N_7436);
or U7860 (N_7860,N_7337,N_7198);
or U7861 (N_7861,N_7160,N_7321);
xnor U7862 (N_7862,N_7495,N_7350);
nand U7863 (N_7863,N_7307,N_7211);
and U7864 (N_7864,N_7410,N_7484);
nand U7865 (N_7865,N_7056,N_7116);
nor U7866 (N_7866,N_6923,N_7425);
and U7867 (N_7867,N_7286,N_7184);
nand U7868 (N_7868,N_7036,N_7305);
or U7869 (N_7869,N_6973,N_7344);
or U7870 (N_7870,N_7260,N_7277);
or U7871 (N_7871,N_7180,N_6937);
or U7872 (N_7872,N_7401,N_7492);
nor U7873 (N_7873,N_7343,N_7185);
and U7874 (N_7874,N_7222,N_7141);
or U7875 (N_7875,N_7398,N_7384);
nand U7876 (N_7876,N_6964,N_7419);
nor U7877 (N_7877,N_7197,N_7425);
or U7878 (N_7878,N_6962,N_7112);
and U7879 (N_7879,N_7318,N_6979);
or U7880 (N_7880,N_7367,N_7084);
and U7881 (N_7881,N_7409,N_7260);
nor U7882 (N_7882,N_6883,N_7298);
or U7883 (N_7883,N_6961,N_7289);
nand U7884 (N_7884,N_6968,N_6987);
xnor U7885 (N_7885,N_7387,N_7365);
nor U7886 (N_7886,N_7174,N_7424);
or U7887 (N_7887,N_7415,N_7256);
nand U7888 (N_7888,N_7427,N_7232);
xnor U7889 (N_7889,N_7063,N_6972);
or U7890 (N_7890,N_7159,N_7327);
nor U7891 (N_7891,N_7167,N_7360);
nor U7892 (N_7892,N_7244,N_7173);
and U7893 (N_7893,N_7187,N_6937);
nor U7894 (N_7894,N_6912,N_7258);
nand U7895 (N_7895,N_6972,N_7330);
nor U7896 (N_7896,N_7383,N_7432);
xnor U7897 (N_7897,N_7317,N_7199);
and U7898 (N_7898,N_7328,N_7239);
nor U7899 (N_7899,N_7417,N_7384);
nor U7900 (N_7900,N_7390,N_6976);
nand U7901 (N_7901,N_7217,N_7450);
nand U7902 (N_7902,N_6905,N_7306);
nand U7903 (N_7903,N_6908,N_6984);
and U7904 (N_7904,N_7426,N_7223);
nand U7905 (N_7905,N_7444,N_7234);
xnor U7906 (N_7906,N_7354,N_7061);
and U7907 (N_7907,N_6957,N_7496);
xor U7908 (N_7908,N_7247,N_7354);
nand U7909 (N_7909,N_7405,N_7492);
or U7910 (N_7910,N_6941,N_7215);
nor U7911 (N_7911,N_7014,N_6887);
and U7912 (N_7912,N_7126,N_7276);
nand U7913 (N_7913,N_7320,N_7144);
xor U7914 (N_7914,N_6909,N_6903);
or U7915 (N_7915,N_6950,N_7049);
nor U7916 (N_7916,N_7230,N_7198);
nand U7917 (N_7917,N_6920,N_7461);
or U7918 (N_7918,N_7305,N_7398);
and U7919 (N_7919,N_6902,N_7166);
nand U7920 (N_7920,N_7405,N_7278);
nor U7921 (N_7921,N_6900,N_7034);
xnor U7922 (N_7922,N_7483,N_7327);
or U7923 (N_7923,N_7342,N_7017);
nand U7924 (N_7924,N_7136,N_7257);
or U7925 (N_7925,N_6992,N_7303);
or U7926 (N_7926,N_7225,N_7292);
nor U7927 (N_7927,N_7014,N_7432);
nor U7928 (N_7928,N_6899,N_7159);
nor U7929 (N_7929,N_6911,N_6921);
and U7930 (N_7930,N_7179,N_6908);
nor U7931 (N_7931,N_7172,N_7340);
nand U7932 (N_7932,N_6996,N_7227);
and U7933 (N_7933,N_7390,N_7056);
or U7934 (N_7934,N_7006,N_7274);
and U7935 (N_7935,N_7416,N_7447);
nor U7936 (N_7936,N_7201,N_7031);
and U7937 (N_7937,N_7122,N_6993);
and U7938 (N_7938,N_7441,N_7223);
nor U7939 (N_7939,N_7061,N_7180);
nor U7940 (N_7940,N_7197,N_7233);
or U7941 (N_7941,N_7309,N_7006);
nor U7942 (N_7942,N_7406,N_6964);
nor U7943 (N_7943,N_7353,N_6926);
nor U7944 (N_7944,N_7397,N_7067);
nand U7945 (N_7945,N_7177,N_6942);
nand U7946 (N_7946,N_7468,N_6926);
xnor U7947 (N_7947,N_6892,N_6978);
nand U7948 (N_7948,N_7157,N_7043);
or U7949 (N_7949,N_7183,N_7226);
or U7950 (N_7950,N_7389,N_7264);
nor U7951 (N_7951,N_7334,N_7426);
and U7952 (N_7952,N_7468,N_7451);
xor U7953 (N_7953,N_7275,N_7273);
or U7954 (N_7954,N_7456,N_7363);
xor U7955 (N_7955,N_6973,N_7086);
nand U7956 (N_7956,N_6902,N_7315);
nor U7957 (N_7957,N_7081,N_7090);
and U7958 (N_7958,N_7342,N_6904);
or U7959 (N_7959,N_7456,N_7479);
nand U7960 (N_7960,N_6993,N_7129);
nand U7961 (N_7961,N_7370,N_7277);
nor U7962 (N_7962,N_7283,N_7328);
nand U7963 (N_7963,N_7060,N_7049);
nand U7964 (N_7964,N_7367,N_7385);
xnor U7965 (N_7965,N_7237,N_7169);
or U7966 (N_7966,N_7371,N_7027);
and U7967 (N_7967,N_7426,N_7133);
nor U7968 (N_7968,N_7285,N_7128);
and U7969 (N_7969,N_6898,N_7015);
nor U7970 (N_7970,N_6877,N_7312);
nand U7971 (N_7971,N_6890,N_7358);
nand U7972 (N_7972,N_7054,N_7146);
and U7973 (N_7973,N_7053,N_7391);
or U7974 (N_7974,N_7059,N_7441);
and U7975 (N_7975,N_7117,N_7444);
and U7976 (N_7976,N_6983,N_7015);
and U7977 (N_7977,N_6888,N_7212);
nor U7978 (N_7978,N_7037,N_7145);
and U7979 (N_7979,N_7011,N_7493);
and U7980 (N_7980,N_7081,N_7334);
or U7981 (N_7981,N_7240,N_7042);
nand U7982 (N_7982,N_7133,N_7459);
nand U7983 (N_7983,N_6888,N_6876);
xnor U7984 (N_7984,N_7246,N_7059);
xnor U7985 (N_7985,N_6994,N_7055);
or U7986 (N_7986,N_7254,N_7115);
nand U7987 (N_7987,N_7105,N_7028);
nor U7988 (N_7988,N_7436,N_7332);
xnor U7989 (N_7989,N_6906,N_7293);
nand U7990 (N_7990,N_7475,N_6917);
or U7991 (N_7991,N_7271,N_7293);
and U7992 (N_7992,N_7336,N_7091);
nor U7993 (N_7993,N_6993,N_7281);
nor U7994 (N_7994,N_7188,N_7466);
and U7995 (N_7995,N_7112,N_7039);
nand U7996 (N_7996,N_7091,N_7070);
and U7997 (N_7997,N_7043,N_7288);
and U7998 (N_7998,N_7065,N_6891);
nand U7999 (N_7999,N_7242,N_7064);
and U8000 (N_8000,N_7282,N_6968);
and U8001 (N_8001,N_7373,N_7080);
nor U8002 (N_8002,N_7430,N_7063);
and U8003 (N_8003,N_7029,N_7301);
and U8004 (N_8004,N_7177,N_6880);
nor U8005 (N_8005,N_6902,N_7057);
nand U8006 (N_8006,N_7437,N_7032);
nor U8007 (N_8007,N_6887,N_7130);
or U8008 (N_8008,N_7133,N_7296);
or U8009 (N_8009,N_7084,N_7234);
or U8010 (N_8010,N_7339,N_7097);
or U8011 (N_8011,N_7062,N_7408);
xor U8012 (N_8012,N_7494,N_7414);
nor U8013 (N_8013,N_7346,N_6971);
nor U8014 (N_8014,N_7075,N_7383);
and U8015 (N_8015,N_7301,N_6904);
or U8016 (N_8016,N_7271,N_7051);
nand U8017 (N_8017,N_7462,N_6982);
and U8018 (N_8018,N_6934,N_7018);
nor U8019 (N_8019,N_7150,N_6898);
nand U8020 (N_8020,N_7149,N_7384);
nor U8021 (N_8021,N_6925,N_7376);
and U8022 (N_8022,N_7224,N_7074);
and U8023 (N_8023,N_6899,N_7429);
nand U8024 (N_8024,N_6914,N_6936);
nand U8025 (N_8025,N_6883,N_7376);
and U8026 (N_8026,N_7358,N_6914);
and U8027 (N_8027,N_7283,N_7201);
nor U8028 (N_8028,N_7220,N_7444);
nor U8029 (N_8029,N_7423,N_6891);
and U8030 (N_8030,N_7496,N_7269);
nand U8031 (N_8031,N_7447,N_6951);
nor U8032 (N_8032,N_6981,N_7071);
nor U8033 (N_8033,N_7364,N_7351);
and U8034 (N_8034,N_7142,N_7359);
or U8035 (N_8035,N_7397,N_7044);
nand U8036 (N_8036,N_7039,N_7386);
nand U8037 (N_8037,N_7084,N_7432);
nor U8038 (N_8038,N_7165,N_7234);
or U8039 (N_8039,N_7431,N_7311);
nor U8040 (N_8040,N_7249,N_6979);
or U8041 (N_8041,N_7022,N_6889);
and U8042 (N_8042,N_6950,N_7249);
xnor U8043 (N_8043,N_7244,N_7102);
nand U8044 (N_8044,N_6991,N_7297);
and U8045 (N_8045,N_7046,N_7237);
nand U8046 (N_8046,N_7026,N_7413);
nand U8047 (N_8047,N_7053,N_7462);
nand U8048 (N_8048,N_7311,N_7339);
nand U8049 (N_8049,N_6974,N_7182);
nor U8050 (N_8050,N_7259,N_6885);
xor U8051 (N_8051,N_7335,N_7471);
nand U8052 (N_8052,N_7049,N_7286);
and U8053 (N_8053,N_7095,N_7354);
nor U8054 (N_8054,N_7256,N_7471);
nand U8055 (N_8055,N_7135,N_7134);
nand U8056 (N_8056,N_7378,N_7159);
and U8057 (N_8057,N_7283,N_7213);
xor U8058 (N_8058,N_7232,N_7378);
or U8059 (N_8059,N_7403,N_6993);
or U8060 (N_8060,N_7395,N_6932);
nand U8061 (N_8061,N_6904,N_7322);
or U8062 (N_8062,N_7088,N_7251);
and U8063 (N_8063,N_7429,N_6993);
nor U8064 (N_8064,N_7459,N_7164);
and U8065 (N_8065,N_6958,N_7384);
xnor U8066 (N_8066,N_6931,N_7109);
or U8067 (N_8067,N_7307,N_7364);
nor U8068 (N_8068,N_7406,N_7149);
nand U8069 (N_8069,N_6997,N_6993);
nor U8070 (N_8070,N_7460,N_7214);
or U8071 (N_8071,N_7138,N_7115);
and U8072 (N_8072,N_7294,N_7279);
xnor U8073 (N_8073,N_7191,N_7123);
nand U8074 (N_8074,N_7237,N_7047);
nor U8075 (N_8075,N_7161,N_7427);
nor U8076 (N_8076,N_7167,N_7244);
or U8077 (N_8077,N_7127,N_7357);
nor U8078 (N_8078,N_6974,N_7396);
nor U8079 (N_8079,N_7363,N_6935);
or U8080 (N_8080,N_7122,N_7369);
nand U8081 (N_8081,N_7291,N_7486);
or U8082 (N_8082,N_7355,N_7074);
xor U8083 (N_8083,N_7441,N_7440);
nand U8084 (N_8084,N_7490,N_6959);
nand U8085 (N_8085,N_6929,N_7448);
and U8086 (N_8086,N_7265,N_7178);
xnor U8087 (N_8087,N_7313,N_7243);
xor U8088 (N_8088,N_7269,N_7315);
nor U8089 (N_8089,N_7360,N_7458);
and U8090 (N_8090,N_7304,N_7026);
and U8091 (N_8091,N_7380,N_6944);
or U8092 (N_8092,N_7119,N_7295);
nor U8093 (N_8093,N_7352,N_7326);
and U8094 (N_8094,N_7405,N_6937);
nor U8095 (N_8095,N_7455,N_7488);
or U8096 (N_8096,N_7323,N_7251);
or U8097 (N_8097,N_7308,N_6932);
nor U8098 (N_8098,N_6882,N_7063);
nor U8099 (N_8099,N_7035,N_7119);
nor U8100 (N_8100,N_7385,N_7476);
nor U8101 (N_8101,N_7021,N_7209);
nor U8102 (N_8102,N_7342,N_7414);
nor U8103 (N_8103,N_7074,N_6878);
nor U8104 (N_8104,N_6968,N_7339);
and U8105 (N_8105,N_7102,N_6902);
nand U8106 (N_8106,N_6996,N_7474);
or U8107 (N_8107,N_6881,N_6885);
nor U8108 (N_8108,N_7021,N_7264);
and U8109 (N_8109,N_7423,N_7326);
nor U8110 (N_8110,N_7406,N_7324);
and U8111 (N_8111,N_7026,N_6916);
nor U8112 (N_8112,N_6930,N_7099);
nor U8113 (N_8113,N_7091,N_7334);
and U8114 (N_8114,N_7381,N_7082);
nor U8115 (N_8115,N_7008,N_7058);
nand U8116 (N_8116,N_7341,N_6943);
nand U8117 (N_8117,N_7055,N_7323);
and U8118 (N_8118,N_6889,N_7105);
nand U8119 (N_8119,N_6893,N_7405);
and U8120 (N_8120,N_7043,N_7311);
nor U8121 (N_8121,N_7373,N_7309);
or U8122 (N_8122,N_7159,N_7365);
nand U8123 (N_8123,N_6964,N_7493);
or U8124 (N_8124,N_7382,N_7097);
or U8125 (N_8125,N_7572,N_8058);
or U8126 (N_8126,N_7776,N_7580);
and U8127 (N_8127,N_8080,N_7985);
nand U8128 (N_8128,N_8026,N_8042);
or U8129 (N_8129,N_8053,N_7745);
nor U8130 (N_8130,N_7685,N_7522);
nand U8131 (N_8131,N_7721,N_7591);
nand U8132 (N_8132,N_7559,N_7868);
nor U8133 (N_8133,N_7658,N_7708);
nor U8134 (N_8134,N_7777,N_7987);
xor U8135 (N_8135,N_8046,N_8089);
nand U8136 (N_8136,N_7983,N_7835);
nor U8137 (N_8137,N_7744,N_7806);
nand U8138 (N_8138,N_7869,N_7765);
nor U8139 (N_8139,N_7696,N_7957);
or U8140 (N_8140,N_7549,N_7668);
xnor U8141 (N_8141,N_8024,N_8102);
nand U8142 (N_8142,N_8075,N_7886);
nor U8143 (N_8143,N_7568,N_7622);
or U8144 (N_8144,N_7904,N_7948);
nor U8145 (N_8145,N_7910,N_7550);
and U8146 (N_8146,N_8039,N_7536);
nor U8147 (N_8147,N_8059,N_7773);
and U8148 (N_8148,N_7864,N_7681);
or U8149 (N_8149,N_8092,N_8040);
nor U8150 (N_8150,N_8054,N_7792);
and U8151 (N_8151,N_7863,N_7737);
nor U8152 (N_8152,N_7761,N_7822);
and U8153 (N_8153,N_7699,N_7624);
nand U8154 (N_8154,N_7933,N_7748);
or U8155 (N_8155,N_7547,N_7596);
nand U8156 (N_8156,N_7819,N_7878);
and U8157 (N_8157,N_7726,N_8067);
nand U8158 (N_8158,N_8049,N_7509);
nand U8159 (N_8159,N_7907,N_7724);
nor U8160 (N_8160,N_8068,N_7538);
nand U8161 (N_8161,N_7562,N_7995);
or U8162 (N_8162,N_7603,N_7992);
nand U8163 (N_8163,N_7990,N_7654);
nand U8164 (N_8164,N_7504,N_7779);
nand U8165 (N_8165,N_7614,N_7859);
nand U8166 (N_8166,N_8063,N_7762);
or U8167 (N_8167,N_7942,N_7648);
nor U8168 (N_8168,N_7690,N_7784);
and U8169 (N_8169,N_8016,N_7931);
nand U8170 (N_8170,N_7760,N_7586);
nand U8171 (N_8171,N_7578,N_8105);
nor U8172 (N_8172,N_8094,N_7976);
nor U8173 (N_8173,N_7857,N_8019);
and U8174 (N_8174,N_7924,N_8004);
and U8175 (N_8175,N_7974,N_7747);
and U8176 (N_8176,N_7853,N_7546);
or U8177 (N_8177,N_7601,N_7834);
nand U8178 (N_8178,N_7955,N_7970);
nor U8179 (N_8179,N_8109,N_7996);
nor U8180 (N_8180,N_8035,N_7675);
or U8181 (N_8181,N_8072,N_7653);
or U8182 (N_8182,N_8103,N_7590);
nor U8183 (N_8183,N_7854,N_8032);
nor U8184 (N_8184,N_7896,N_7585);
or U8185 (N_8185,N_8064,N_8108);
or U8186 (N_8186,N_8076,N_7769);
or U8187 (N_8187,N_8116,N_7888);
nand U8188 (N_8188,N_7557,N_7630);
nor U8189 (N_8189,N_7664,N_7791);
nor U8190 (N_8190,N_7960,N_7519);
and U8191 (N_8191,N_7718,N_7523);
nor U8192 (N_8192,N_7845,N_7553);
and U8193 (N_8193,N_7915,N_7537);
nor U8194 (N_8194,N_8115,N_7635);
xnor U8195 (N_8195,N_7707,N_7876);
xnor U8196 (N_8196,N_7608,N_7623);
and U8197 (N_8197,N_8121,N_7902);
nor U8198 (N_8198,N_7914,N_7820);
nand U8199 (N_8199,N_7821,N_7862);
and U8200 (N_8200,N_7991,N_8090);
nor U8201 (N_8201,N_7947,N_7576);
and U8202 (N_8202,N_7661,N_7583);
and U8203 (N_8203,N_7735,N_8051);
or U8204 (N_8204,N_7962,N_7803);
and U8205 (N_8205,N_7866,N_7698);
or U8206 (N_8206,N_7802,N_8088);
nor U8207 (N_8207,N_7597,N_7598);
and U8208 (N_8208,N_7612,N_8003);
nand U8209 (N_8209,N_7780,N_7582);
nand U8210 (N_8210,N_7558,N_7965);
nor U8211 (N_8211,N_7502,N_7540);
or U8212 (N_8212,N_7678,N_8030);
or U8213 (N_8213,N_7645,N_7934);
nor U8214 (N_8214,N_7741,N_7856);
nand U8215 (N_8215,N_7642,N_7611);
nand U8216 (N_8216,N_7565,N_7671);
nand U8217 (N_8217,N_7694,N_7506);
nand U8218 (N_8218,N_7793,N_7850);
nor U8219 (N_8219,N_7877,N_7579);
xnor U8220 (N_8220,N_8097,N_7534);
nor U8221 (N_8221,N_7984,N_7837);
nand U8222 (N_8222,N_7662,N_7812);
nand U8223 (N_8223,N_7552,N_7945);
nand U8224 (N_8224,N_7652,N_7840);
or U8225 (N_8225,N_7815,N_7541);
or U8226 (N_8226,N_7639,N_8005);
nor U8227 (N_8227,N_7943,N_8110);
nor U8228 (N_8228,N_7725,N_7629);
and U8229 (N_8229,N_7757,N_8056);
nor U8230 (N_8230,N_7617,N_7936);
nor U8231 (N_8231,N_7561,N_7971);
nor U8232 (N_8232,N_7796,N_8013);
and U8233 (N_8233,N_7594,N_7768);
nand U8234 (N_8234,N_7503,N_7879);
nand U8235 (N_8235,N_7829,N_7556);
or U8236 (N_8236,N_8104,N_7743);
nor U8237 (N_8237,N_7927,N_7575);
xnor U8238 (N_8238,N_7849,N_7670);
or U8239 (N_8239,N_7700,N_8044);
and U8240 (N_8240,N_8099,N_7905);
nor U8241 (N_8241,N_7695,N_8015);
and U8242 (N_8242,N_7573,N_7958);
and U8243 (N_8243,N_8098,N_7871);
nor U8244 (N_8244,N_7811,N_8123);
and U8245 (N_8245,N_7609,N_7627);
nor U8246 (N_8246,N_7750,N_7916);
nor U8247 (N_8247,N_7975,N_7649);
and U8248 (N_8248,N_7781,N_8006);
nor U8249 (N_8249,N_7595,N_7918);
and U8250 (N_8250,N_7500,N_7604);
or U8251 (N_8251,N_7589,N_7832);
and U8252 (N_8252,N_7655,N_7688);
nand U8253 (N_8253,N_7892,N_7510);
nand U8254 (N_8254,N_7511,N_7906);
nand U8255 (N_8255,N_7544,N_8107);
or U8256 (N_8256,N_7672,N_7701);
or U8257 (N_8257,N_7989,N_7571);
or U8258 (N_8258,N_7899,N_7501);
nand U8259 (N_8259,N_7938,N_7709);
nor U8260 (N_8260,N_7928,N_7794);
nand U8261 (N_8261,N_7628,N_8120);
or U8262 (N_8262,N_7646,N_7716);
and U8263 (N_8263,N_7911,N_8091);
nor U8264 (N_8264,N_7981,N_7993);
and U8265 (N_8265,N_7795,N_7980);
and U8266 (N_8266,N_8118,N_7754);
nand U8267 (N_8267,N_7706,N_7548);
or U8268 (N_8268,N_7715,N_7673);
nor U8269 (N_8269,N_7844,N_7529);
or U8270 (N_8270,N_7830,N_7873);
and U8271 (N_8271,N_7890,N_7632);
nand U8272 (N_8272,N_8047,N_7677);
nor U8273 (N_8273,N_7659,N_7946);
or U8274 (N_8274,N_7994,N_7808);
nand U8275 (N_8275,N_7533,N_8017);
nor U8276 (N_8276,N_7566,N_7770);
xor U8277 (N_8277,N_7799,N_7691);
nor U8278 (N_8278,N_7783,N_7680);
nor U8279 (N_8279,N_7817,N_7723);
nor U8280 (N_8280,N_7539,N_8029);
or U8281 (N_8281,N_7600,N_7663);
or U8282 (N_8282,N_8086,N_7900);
nor U8283 (N_8283,N_7641,N_8079);
nand U8284 (N_8284,N_7577,N_7764);
and U8285 (N_8285,N_7515,N_7626);
nand U8286 (N_8286,N_8087,N_7588);
or U8287 (N_8287,N_7521,N_7939);
xnor U8288 (N_8288,N_7814,N_8114);
nor U8289 (N_8289,N_8070,N_7887);
or U8290 (N_8290,N_7935,N_7894);
nor U8291 (N_8291,N_7593,N_7669);
and U8292 (N_8292,N_7838,N_7676);
nor U8293 (N_8293,N_7656,N_7736);
or U8294 (N_8294,N_7615,N_7508);
or U8295 (N_8295,N_7731,N_7599);
or U8296 (N_8296,N_8018,N_7711);
and U8297 (N_8297,N_8055,N_7775);
and U8298 (N_8298,N_7651,N_7686);
nor U8299 (N_8299,N_7542,N_7903);
or U8300 (N_8300,N_7967,N_7959);
xor U8301 (N_8301,N_7513,N_7941);
and U8302 (N_8302,N_7619,N_7882);
nand U8303 (N_8303,N_7751,N_7883);
nor U8304 (N_8304,N_7705,N_8010);
xnor U8305 (N_8305,N_7759,N_7875);
or U8306 (N_8306,N_7824,N_7746);
xor U8307 (N_8307,N_7518,N_7913);
and U8308 (N_8308,N_7785,N_7872);
nand U8309 (N_8309,N_8052,N_7969);
xnor U8310 (N_8310,N_7749,N_8100);
and U8311 (N_8311,N_7804,N_8020);
xor U8312 (N_8312,N_7897,N_8096);
xor U8313 (N_8313,N_7587,N_8033);
or U8314 (N_8314,N_7891,N_7940);
or U8315 (N_8315,N_7963,N_7925);
or U8316 (N_8316,N_7895,N_7885);
nand U8317 (N_8317,N_7827,N_7740);
nor U8318 (N_8318,N_7684,N_8048);
and U8319 (N_8319,N_7728,N_8007);
or U8320 (N_8320,N_8061,N_7618);
xnor U8321 (N_8321,N_7826,N_7956);
and U8322 (N_8322,N_7771,N_7836);
or U8323 (N_8323,N_7644,N_8038);
nand U8324 (N_8324,N_8111,N_7514);
nand U8325 (N_8325,N_8045,N_7638);
and U8326 (N_8326,N_7839,N_7825);
nor U8327 (N_8327,N_7666,N_8077);
or U8328 (N_8328,N_8011,N_8023);
or U8329 (N_8329,N_7606,N_8113);
nand U8330 (N_8330,N_7937,N_7909);
nor U8331 (N_8331,N_7602,N_7964);
nor U8332 (N_8332,N_8034,N_8071);
nand U8333 (N_8333,N_7616,N_8031);
or U8334 (N_8334,N_7543,N_7554);
nor U8335 (N_8335,N_7813,N_7634);
nor U8336 (N_8336,N_7852,N_8101);
nor U8337 (N_8337,N_8000,N_8106);
nor U8338 (N_8338,N_7790,N_7867);
nor U8339 (N_8339,N_7767,N_8025);
nand U8340 (N_8340,N_7530,N_7560);
nor U8341 (N_8341,N_7772,N_8085);
nand U8342 (N_8342,N_7732,N_7570);
nor U8343 (N_8343,N_8060,N_7507);
or U8344 (N_8344,N_7528,N_7756);
nor U8345 (N_8345,N_7921,N_7679);
or U8346 (N_8346,N_7823,N_7944);
nand U8347 (N_8347,N_8002,N_8037);
xor U8348 (N_8348,N_7919,N_7842);
or U8349 (N_8349,N_7692,N_7505);
and U8350 (N_8350,N_7843,N_7742);
xnor U8351 (N_8351,N_7551,N_7774);
nand U8352 (N_8352,N_7865,N_7858);
or U8353 (N_8353,N_7874,N_7532);
and U8354 (N_8354,N_7950,N_7755);
nor U8355 (N_8355,N_7810,N_8084);
and U8356 (N_8356,N_7564,N_7569);
and U8357 (N_8357,N_7647,N_7719);
nand U8358 (N_8358,N_8117,N_7930);
xnor U8359 (N_8359,N_7926,N_7636);
nand U8360 (N_8360,N_7816,N_7788);
or U8361 (N_8361,N_7516,N_7977);
nor U8362 (N_8362,N_7613,N_7870);
nor U8363 (N_8363,N_7986,N_8112);
nand U8364 (N_8364,N_7800,N_7999);
nand U8365 (N_8365,N_7951,N_7714);
nand U8366 (N_8366,N_7782,N_7801);
nor U8367 (N_8367,N_7923,N_7702);
nor U8368 (N_8368,N_7847,N_8027);
or U8369 (N_8369,N_7524,N_7643);
nand U8370 (N_8370,N_7978,N_8008);
and U8371 (N_8371,N_8065,N_7846);
nor U8372 (N_8372,N_7932,N_7683);
xnor U8373 (N_8373,N_7657,N_7966);
nand U8374 (N_8374,N_7789,N_7901);
nor U8375 (N_8375,N_7730,N_8066);
and U8376 (N_8376,N_7633,N_7833);
or U8377 (N_8377,N_7786,N_7893);
nand U8378 (N_8378,N_7739,N_7687);
or U8379 (N_8379,N_7798,N_7531);
nor U8380 (N_8380,N_7512,N_7831);
or U8381 (N_8381,N_7880,N_7778);
and U8382 (N_8382,N_7689,N_8022);
nand U8383 (N_8383,N_8074,N_7581);
nor U8384 (N_8384,N_8012,N_7605);
nand U8385 (N_8385,N_7982,N_8014);
nand U8386 (N_8386,N_7545,N_7787);
and U8387 (N_8387,N_7631,N_7860);
nand U8388 (N_8388,N_7952,N_7697);
nor U8389 (N_8389,N_7929,N_8062);
or U8390 (N_8390,N_7851,N_7908);
or U8391 (N_8391,N_7674,N_7682);
xnor U8392 (N_8392,N_7520,N_7693);
nand U8393 (N_8393,N_7574,N_7720);
and U8394 (N_8394,N_7667,N_7881);
nand U8395 (N_8395,N_8093,N_7704);
nand U8396 (N_8396,N_8050,N_7640);
nand U8397 (N_8397,N_7758,N_8082);
and U8398 (N_8398,N_7752,N_7912);
nand U8399 (N_8399,N_7650,N_8122);
and U8400 (N_8400,N_7584,N_8036);
nand U8401 (N_8401,N_7972,N_7592);
nor U8402 (N_8402,N_7861,N_7703);
or U8403 (N_8403,N_8043,N_7729);
or U8404 (N_8404,N_7734,N_8009);
and U8405 (N_8405,N_8041,N_7527);
or U8406 (N_8406,N_8001,N_8124);
nor U8407 (N_8407,N_7625,N_7525);
or U8408 (N_8408,N_8057,N_7973);
nand U8409 (N_8409,N_7563,N_7717);
and U8410 (N_8410,N_7526,N_7855);
or U8411 (N_8411,N_7898,N_8119);
nor U8412 (N_8412,N_7920,N_7998);
nor U8413 (N_8413,N_7805,N_7807);
nand U8414 (N_8414,N_7712,N_7607);
and U8415 (N_8415,N_7968,N_7818);
nand U8416 (N_8416,N_8073,N_7809);
and U8417 (N_8417,N_8069,N_7884);
nand U8418 (N_8418,N_7738,N_7665);
nor U8419 (N_8419,N_8095,N_7621);
xnor U8420 (N_8420,N_7555,N_7997);
and U8421 (N_8421,N_7535,N_8078);
nor U8422 (N_8422,N_7722,N_7922);
nand U8423 (N_8423,N_7797,N_7841);
nor U8424 (N_8424,N_7610,N_7763);
or U8425 (N_8425,N_8028,N_7753);
nor U8426 (N_8426,N_7567,N_7988);
nor U8427 (N_8427,N_7620,N_7660);
or U8428 (N_8428,N_7517,N_7766);
nor U8429 (N_8429,N_7713,N_8083);
xnor U8430 (N_8430,N_7954,N_7727);
nor U8431 (N_8431,N_7889,N_7949);
and U8432 (N_8432,N_7961,N_7733);
nand U8433 (N_8433,N_7637,N_7710);
xor U8434 (N_8434,N_7917,N_7979);
nor U8435 (N_8435,N_8021,N_8081);
or U8436 (N_8436,N_7828,N_7953);
and U8437 (N_8437,N_7848,N_7911);
nor U8438 (N_8438,N_7509,N_7802);
nand U8439 (N_8439,N_7807,N_8019);
xor U8440 (N_8440,N_7790,N_8011);
or U8441 (N_8441,N_7823,N_7934);
nand U8442 (N_8442,N_7525,N_8082);
and U8443 (N_8443,N_7654,N_7803);
and U8444 (N_8444,N_7832,N_7785);
xnor U8445 (N_8445,N_7786,N_7760);
nand U8446 (N_8446,N_7829,N_7704);
and U8447 (N_8447,N_7633,N_8060);
and U8448 (N_8448,N_7756,N_8087);
nor U8449 (N_8449,N_7810,N_8000);
or U8450 (N_8450,N_7636,N_7878);
nor U8451 (N_8451,N_7973,N_7556);
and U8452 (N_8452,N_7932,N_7665);
or U8453 (N_8453,N_8034,N_7624);
or U8454 (N_8454,N_7807,N_8099);
nor U8455 (N_8455,N_7791,N_7716);
and U8456 (N_8456,N_7718,N_7713);
nor U8457 (N_8457,N_7548,N_7958);
xnor U8458 (N_8458,N_7997,N_7505);
and U8459 (N_8459,N_7550,N_7893);
and U8460 (N_8460,N_7728,N_8015);
or U8461 (N_8461,N_7740,N_7983);
nor U8462 (N_8462,N_7731,N_8115);
nor U8463 (N_8463,N_8112,N_7680);
nand U8464 (N_8464,N_7509,N_7810);
nand U8465 (N_8465,N_7674,N_8112);
or U8466 (N_8466,N_7954,N_7675);
or U8467 (N_8467,N_7708,N_7759);
or U8468 (N_8468,N_7753,N_7654);
nand U8469 (N_8469,N_7860,N_7946);
or U8470 (N_8470,N_7901,N_7920);
and U8471 (N_8471,N_7824,N_7750);
xor U8472 (N_8472,N_8015,N_7511);
nor U8473 (N_8473,N_7771,N_7846);
and U8474 (N_8474,N_8007,N_7952);
nand U8475 (N_8475,N_7913,N_7878);
nand U8476 (N_8476,N_7813,N_7524);
nand U8477 (N_8477,N_8051,N_7913);
nand U8478 (N_8478,N_7831,N_7676);
nand U8479 (N_8479,N_7753,N_7915);
xnor U8480 (N_8480,N_7773,N_8005);
and U8481 (N_8481,N_7963,N_7720);
or U8482 (N_8482,N_7855,N_7622);
or U8483 (N_8483,N_7720,N_7768);
nand U8484 (N_8484,N_7542,N_7673);
nor U8485 (N_8485,N_7618,N_7864);
nor U8486 (N_8486,N_7732,N_7745);
nand U8487 (N_8487,N_8080,N_8081);
nand U8488 (N_8488,N_8095,N_8116);
or U8489 (N_8489,N_7867,N_7573);
nand U8490 (N_8490,N_7563,N_8060);
nand U8491 (N_8491,N_7905,N_7944);
and U8492 (N_8492,N_8115,N_7898);
xor U8493 (N_8493,N_7820,N_7722);
nand U8494 (N_8494,N_7569,N_7623);
nor U8495 (N_8495,N_7950,N_7553);
nor U8496 (N_8496,N_7953,N_7839);
and U8497 (N_8497,N_7777,N_8018);
or U8498 (N_8498,N_7612,N_8014);
nand U8499 (N_8499,N_8067,N_7551);
nor U8500 (N_8500,N_8000,N_7582);
nor U8501 (N_8501,N_7930,N_7767);
nor U8502 (N_8502,N_7607,N_8086);
and U8503 (N_8503,N_7864,N_7952);
nor U8504 (N_8504,N_7769,N_7645);
or U8505 (N_8505,N_7557,N_8108);
xor U8506 (N_8506,N_7924,N_7703);
nor U8507 (N_8507,N_8117,N_8087);
or U8508 (N_8508,N_8121,N_7815);
nor U8509 (N_8509,N_8119,N_7669);
xor U8510 (N_8510,N_7741,N_8016);
and U8511 (N_8511,N_7650,N_8076);
nor U8512 (N_8512,N_8101,N_7521);
nor U8513 (N_8513,N_7770,N_7585);
or U8514 (N_8514,N_7657,N_7861);
xnor U8515 (N_8515,N_8084,N_7595);
or U8516 (N_8516,N_7829,N_7939);
nand U8517 (N_8517,N_7827,N_7942);
or U8518 (N_8518,N_7558,N_7778);
or U8519 (N_8519,N_7606,N_7517);
xor U8520 (N_8520,N_8029,N_7817);
or U8521 (N_8521,N_8098,N_7577);
and U8522 (N_8522,N_8113,N_7918);
nor U8523 (N_8523,N_7633,N_7907);
or U8524 (N_8524,N_7766,N_7568);
or U8525 (N_8525,N_8080,N_7611);
and U8526 (N_8526,N_7526,N_7555);
nand U8527 (N_8527,N_7502,N_7913);
or U8528 (N_8528,N_7878,N_7599);
or U8529 (N_8529,N_7644,N_7733);
nand U8530 (N_8530,N_7751,N_7729);
and U8531 (N_8531,N_7802,N_8118);
or U8532 (N_8532,N_7842,N_7566);
and U8533 (N_8533,N_7723,N_7782);
nand U8534 (N_8534,N_7639,N_7818);
xnor U8535 (N_8535,N_7936,N_7774);
nor U8536 (N_8536,N_8054,N_7834);
or U8537 (N_8537,N_7984,N_7786);
nand U8538 (N_8538,N_7888,N_7774);
nand U8539 (N_8539,N_7917,N_7949);
nand U8540 (N_8540,N_7509,N_7611);
xor U8541 (N_8541,N_7574,N_7567);
and U8542 (N_8542,N_8107,N_7605);
xor U8543 (N_8543,N_7609,N_7691);
nor U8544 (N_8544,N_7793,N_8037);
nand U8545 (N_8545,N_7641,N_7611);
nand U8546 (N_8546,N_7902,N_8000);
nand U8547 (N_8547,N_7760,N_7516);
or U8548 (N_8548,N_7568,N_7759);
or U8549 (N_8549,N_7502,N_7769);
nand U8550 (N_8550,N_8077,N_8110);
and U8551 (N_8551,N_8030,N_7666);
or U8552 (N_8552,N_7736,N_7507);
nand U8553 (N_8553,N_7655,N_7979);
nor U8554 (N_8554,N_7998,N_7526);
nor U8555 (N_8555,N_7930,N_7661);
and U8556 (N_8556,N_7854,N_7718);
and U8557 (N_8557,N_7536,N_8061);
or U8558 (N_8558,N_7905,N_7872);
nor U8559 (N_8559,N_7991,N_7655);
nor U8560 (N_8560,N_7545,N_7650);
and U8561 (N_8561,N_8096,N_7536);
nand U8562 (N_8562,N_8054,N_7712);
and U8563 (N_8563,N_7750,N_7857);
and U8564 (N_8564,N_7654,N_7623);
nand U8565 (N_8565,N_7905,N_8060);
nand U8566 (N_8566,N_7793,N_8123);
nor U8567 (N_8567,N_8113,N_7839);
nor U8568 (N_8568,N_7834,N_8011);
and U8569 (N_8569,N_7988,N_7645);
or U8570 (N_8570,N_7923,N_7575);
xor U8571 (N_8571,N_7691,N_8022);
or U8572 (N_8572,N_7673,N_7617);
or U8573 (N_8573,N_8109,N_7774);
and U8574 (N_8574,N_7903,N_7595);
nand U8575 (N_8575,N_8037,N_8014);
nand U8576 (N_8576,N_7661,N_7671);
or U8577 (N_8577,N_8020,N_8108);
and U8578 (N_8578,N_7950,N_7630);
or U8579 (N_8579,N_7944,N_7718);
nor U8580 (N_8580,N_7828,N_7740);
nor U8581 (N_8581,N_8068,N_7972);
nand U8582 (N_8582,N_8056,N_7872);
or U8583 (N_8583,N_7968,N_7950);
xnor U8584 (N_8584,N_7873,N_7737);
and U8585 (N_8585,N_7942,N_7646);
or U8586 (N_8586,N_7579,N_7643);
nor U8587 (N_8587,N_7791,N_7518);
nand U8588 (N_8588,N_7747,N_8120);
nand U8589 (N_8589,N_8037,N_7580);
nor U8590 (N_8590,N_7970,N_7584);
nor U8591 (N_8591,N_7585,N_7861);
nand U8592 (N_8592,N_8095,N_7988);
xor U8593 (N_8593,N_8029,N_7624);
or U8594 (N_8594,N_7633,N_8097);
and U8595 (N_8595,N_7523,N_7783);
nor U8596 (N_8596,N_7879,N_8051);
nand U8597 (N_8597,N_7742,N_7751);
and U8598 (N_8598,N_7707,N_8058);
nand U8599 (N_8599,N_7731,N_7868);
xnor U8600 (N_8600,N_7580,N_7782);
nand U8601 (N_8601,N_7522,N_7870);
or U8602 (N_8602,N_8057,N_7805);
and U8603 (N_8603,N_7828,N_7925);
or U8604 (N_8604,N_8072,N_8107);
nor U8605 (N_8605,N_7615,N_7929);
nand U8606 (N_8606,N_8118,N_8057);
nand U8607 (N_8607,N_7626,N_7930);
nor U8608 (N_8608,N_8030,N_8082);
or U8609 (N_8609,N_8077,N_7863);
xnor U8610 (N_8610,N_7554,N_7599);
or U8611 (N_8611,N_7730,N_7503);
or U8612 (N_8612,N_8113,N_7719);
nand U8613 (N_8613,N_7947,N_7979);
or U8614 (N_8614,N_7622,N_7683);
nand U8615 (N_8615,N_7662,N_7589);
or U8616 (N_8616,N_7629,N_7617);
and U8617 (N_8617,N_8015,N_7769);
and U8618 (N_8618,N_7505,N_7985);
and U8619 (N_8619,N_7541,N_7527);
nor U8620 (N_8620,N_7720,N_8102);
nor U8621 (N_8621,N_8025,N_7742);
nor U8622 (N_8622,N_8116,N_7606);
nor U8623 (N_8623,N_7839,N_8062);
xor U8624 (N_8624,N_7874,N_7756);
xor U8625 (N_8625,N_7515,N_7637);
or U8626 (N_8626,N_7664,N_7666);
xnor U8627 (N_8627,N_7612,N_7625);
xor U8628 (N_8628,N_7924,N_7587);
nand U8629 (N_8629,N_7953,N_7866);
nand U8630 (N_8630,N_7565,N_8009);
nor U8631 (N_8631,N_7826,N_8008);
nand U8632 (N_8632,N_7520,N_7998);
nor U8633 (N_8633,N_7994,N_7719);
nor U8634 (N_8634,N_7937,N_7819);
nor U8635 (N_8635,N_7885,N_7658);
or U8636 (N_8636,N_7754,N_8116);
and U8637 (N_8637,N_7660,N_7694);
nor U8638 (N_8638,N_7752,N_7681);
and U8639 (N_8639,N_7539,N_7914);
nand U8640 (N_8640,N_8025,N_8102);
or U8641 (N_8641,N_7920,N_7697);
nand U8642 (N_8642,N_8084,N_8014);
or U8643 (N_8643,N_8078,N_7949);
xor U8644 (N_8644,N_7977,N_8083);
nor U8645 (N_8645,N_7528,N_7884);
nor U8646 (N_8646,N_7556,N_7546);
nand U8647 (N_8647,N_7775,N_7770);
and U8648 (N_8648,N_8018,N_8069);
xor U8649 (N_8649,N_7538,N_8108);
xor U8650 (N_8650,N_8066,N_7995);
nor U8651 (N_8651,N_8024,N_8039);
or U8652 (N_8652,N_7957,N_7860);
nand U8653 (N_8653,N_7524,N_8047);
xnor U8654 (N_8654,N_7837,N_7816);
nor U8655 (N_8655,N_8039,N_7605);
nand U8656 (N_8656,N_7821,N_7536);
nand U8657 (N_8657,N_8035,N_7665);
or U8658 (N_8658,N_7677,N_7865);
and U8659 (N_8659,N_7989,N_8046);
and U8660 (N_8660,N_7629,N_7520);
xnor U8661 (N_8661,N_7608,N_7546);
nand U8662 (N_8662,N_8036,N_7605);
nand U8663 (N_8663,N_7631,N_8067);
nand U8664 (N_8664,N_7698,N_7719);
or U8665 (N_8665,N_7650,N_7896);
and U8666 (N_8666,N_7971,N_7816);
nand U8667 (N_8667,N_7878,N_7723);
xor U8668 (N_8668,N_7894,N_7770);
or U8669 (N_8669,N_7985,N_7600);
nand U8670 (N_8670,N_7803,N_7713);
nand U8671 (N_8671,N_7522,N_8020);
nand U8672 (N_8672,N_7559,N_7927);
and U8673 (N_8673,N_7757,N_7917);
nand U8674 (N_8674,N_7989,N_7966);
xor U8675 (N_8675,N_7603,N_7793);
or U8676 (N_8676,N_7620,N_7834);
or U8677 (N_8677,N_8074,N_7627);
nor U8678 (N_8678,N_7623,N_7680);
nor U8679 (N_8679,N_7984,N_7606);
or U8680 (N_8680,N_7684,N_7553);
nor U8681 (N_8681,N_7874,N_7565);
nor U8682 (N_8682,N_8115,N_7645);
xnor U8683 (N_8683,N_7884,N_7734);
nand U8684 (N_8684,N_7687,N_8083);
and U8685 (N_8685,N_7512,N_8008);
or U8686 (N_8686,N_7696,N_7823);
or U8687 (N_8687,N_8087,N_7596);
nor U8688 (N_8688,N_7743,N_7822);
nor U8689 (N_8689,N_7982,N_7611);
nor U8690 (N_8690,N_7667,N_7546);
nand U8691 (N_8691,N_7935,N_7907);
and U8692 (N_8692,N_7506,N_7557);
nor U8693 (N_8693,N_7783,N_8107);
nor U8694 (N_8694,N_7601,N_7964);
nor U8695 (N_8695,N_8061,N_7973);
nor U8696 (N_8696,N_8015,N_7547);
nand U8697 (N_8697,N_7576,N_7760);
and U8698 (N_8698,N_7729,N_7843);
and U8699 (N_8699,N_7648,N_7609);
or U8700 (N_8700,N_7746,N_7889);
nand U8701 (N_8701,N_7903,N_8096);
or U8702 (N_8702,N_7775,N_7727);
nor U8703 (N_8703,N_7746,N_7953);
and U8704 (N_8704,N_7945,N_7592);
nand U8705 (N_8705,N_7935,N_8118);
nand U8706 (N_8706,N_7590,N_7817);
nor U8707 (N_8707,N_7837,N_7924);
and U8708 (N_8708,N_7870,N_7664);
xnor U8709 (N_8709,N_8011,N_7624);
nor U8710 (N_8710,N_7852,N_7779);
nand U8711 (N_8711,N_7639,N_7791);
or U8712 (N_8712,N_7520,N_7600);
and U8713 (N_8713,N_7698,N_7580);
nand U8714 (N_8714,N_7886,N_7715);
nand U8715 (N_8715,N_7719,N_7960);
nor U8716 (N_8716,N_7742,N_7766);
nor U8717 (N_8717,N_8039,N_7620);
nand U8718 (N_8718,N_7871,N_8071);
xor U8719 (N_8719,N_7605,N_7507);
and U8720 (N_8720,N_7761,N_7575);
and U8721 (N_8721,N_7851,N_7713);
nand U8722 (N_8722,N_7537,N_7721);
xor U8723 (N_8723,N_7598,N_7727);
nor U8724 (N_8724,N_7736,N_7564);
nor U8725 (N_8725,N_8114,N_7867);
or U8726 (N_8726,N_7663,N_7536);
xor U8727 (N_8727,N_7608,N_7837);
nor U8728 (N_8728,N_7598,N_7899);
and U8729 (N_8729,N_7506,N_7673);
nor U8730 (N_8730,N_7921,N_7972);
or U8731 (N_8731,N_7875,N_7891);
nor U8732 (N_8732,N_7533,N_8030);
or U8733 (N_8733,N_7542,N_7545);
nor U8734 (N_8734,N_7935,N_7699);
nand U8735 (N_8735,N_7596,N_7852);
nand U8736 (N_8736,N_7920,N_7937);
nor U8737 (N_8737,N_7554,N_7592);
nand U8738 (N_8738,N_7788,N_8073);
or U8739 (N_8739,N_7754,N_8002);
or U8740 (N_8740,N_7532,N_7935);
xnor U8741 (N_8741,N_7905,N_7547);
nor U8742 (N_8742,N_7849,N_7544);
and U8743 (N_8743,N_7615,N_7700);
nor U8744 (N_8744,N_7643,N_7749);
nand U8745 (N_8745,N_7664,N_7845);
and U8746 (N_8746,N_7643,N_8112);
nor U8747 (N_8747,N_7535,N_7875);
xnor U8748 (N_8748,N_7850,N_7761);
nand U8749 (N_8749,N_7861,N_7826);
nand U8750 (N_8750,N_8539,N_8168);
and U8751 (N_8751,N_8308,N_8190);
nand U8752 (N_8752,N_8321,N_8603);
or U8753 (N_8753,N_8716,N_8303);
or U8754 (N_8754,N_8326,N_8710);
and U8755 (N_8755,N_8183,N_8137);
nor U8756 (N_8756,N_8745,N_8648);
or U8757 (N_8757,N_8417,N_8240);
nor U8758 (N_8758,N_8675,N_8467);
or U8759 (N_8759,N_8257,N_8234);
or U8760 (N_8760,N_8709,N_8747);
or U8761 (N_8761,N_8211,N_8705);
nor U8762 (N_8762,N_8311,N_8480);
xnor U8763 (N_8763,N_8496,N_8582);
or U8764 (N_8764,N_8169,N_8746);
xnor U8765 (N_8765,N_8590,N_8387);
nor U8766 (N_8766,N_8152,N_8577);
or U8767 (N_8767,N_8452,N_8679);
nor U8768 (N_8768,N_8196,N_8701);
nand U8769 (N_8769,N_8600,N_8427);
nand U8770 (N_8770,N_8663,N_8409);
nand U8771 (N_8771,N_8278,N_8424);
nand U8772 (N_8772,N_8639,N_8213);
xnor U8773 (N_8773,N_8397,N_8544);
or U8774 (N_8774,N_8718,N_8394);
and U8775 (N_8775,N_8229,N_8699);
nor U8776 (N_8776,N_8595,N_8160);
nor U8777 (N_8777,N_8349,N_8332);
and U8778 (N_8778,N_8301,N_8594);
nor U8779 (N_8779,N_8127,N_8529);
nor U8780 (N_8780,N_8602,N_8445);
nor U8781 (N_8781,N_8414,N_8475);
nor U8782 (N_8782,N_8202,N_8545);
nand U8783 (N_8783,N_8572,N_8620);
and U8784 (N_8784,N_8179,N_8531);
and U8785 (N_8785,N_8191,N_8651);
nand U8786 (N_8786,N_8739,N_8297);
nand U8787 (N_8787,N_8265,N_8574);
nor U8788 (N_8788,N_8540,N_8376);
nor U8789 (N_8789,N_8547,N_8158);
and U8790 (N_8790,N_8333,N_8631);
xnor U8791 (N_8791,N_8453,N_8722);
and U8792 (N_8792,N_8459,N_8309);
nand U8793 (N_8793,N_8177,N_8432);
or U8794 (N_8794,N_8134,N_8686);
and U8795 (N_8795,N_8707,N_8357);
and U8796 (N_8796,N_8729,N_8398);
or U8797 (N_8797,N_8306,N_8528);
or U8798 (N_8798,N_8492,N_8624);
and U8799 (N_8799,N_8388,N_8222);
xnor U8800 (N_8800,N_8233,N_8421);
or U8801 (N_8801,N_8552,N_8367);
and U8802 (N_8802,N_8411,N_8185);
xor U8803 (N_8803,N_8198,N_8246);
nand U8804 (N_8804,N_8247,N_8142);
or U8805 (N_8805,N_8659,N_8541);
xor U8806 (N_8806,N_8714,N_8462);
nor U8807 (N_8807,N_8228,N_8484);
or U8808 (N_8808,N_8738,N_8132);
or U8809 (N_8809,N_8640,N_8438);
and U8810 (N_8810,N_8319,N_8342);
nor U8811 (N_8811,N_8323,N_8749);
xor U8812 (N_8812,N_8621,N_8192);
or U8813 (N_8813,N_8283,N_8286);
and U8814 (N_8814,N_8573,N_8609);
or U8815 (N_8815,N_8214,N_8643);
xor U8816 (N_8816,N_8386,N_8696);
nor U8817 (N_8817,N_8382,N_8684);
and U8818 (N_8818,N_8607,N_8506);
and U8819 (N_8819,N_8435,N_8472);
or U8820 (N_8820,N_8448,N_8622);
xor U8821 (N_8821,N_8526,N_8673);
and U8822 (N_8822,N_8530,N_8685);
nand U8823 (N_8823,N_8338,N_8290);
or U8824 (N_8824,N_8189,N_8688);
nand U8825 (N_8825,N_8500,N_8608);
nor U8826 (N_8826,N_8724,N_8721);
or U8827 (N_8827,N_8180,N_8592);
nand U8828 (N_8828,N_8549,N_8460);
and U8829 (N_8829,N_8351,N_8300);
and U8830 (N_8830,N_8741,N_8428);
and U8831 (N_8831,N_8470,N_8429);
or U8832 (N_8832,N_8310,N_8404);
nor U8833 (N_8833,N_8125,N_8511);
nor U8834 (N_8834,N_8578,N_8454);
and U8835 (N_8835,N_8706,N_8412);
nand U8836 (N_8836,N_8599,N_8258);
and U8837 (N_8837,N_8383,N_8426);
or U8838 (N_8838,N_8525,N_8261);
and U8839 (N_8839,N_8584,N_8456);
or U8840 (N_8840,N_8365,N_8353);
nor U8841 (N_8841,N_8564,N_8654);
nand U8842 (N_8842,N_8458,N_8711);
nor U8843 (N_8843,N_8556,N_8419);
xor U8844 (N_8844,N_8227,N_8245);
xor U8845 (N_8845,N_8166,N_8400);
xnor U8846 (N_8846,N_8702,N_8256);
xor U8847 (N_8847,N_8270,N_8476);
nand U8848 (N_8848,N_8512,N_8662);
and U8849 (N_8849,N_8508,N_8363);
and U8850 (N_8850,N_8567,N_8217);
nand U8851 (N_8851,N_8474,N_8399);
and U8852 (N_8852,N_8146,N_8489);
nor U8853 (N_8853,N_8153,N_8628);
nor U8854 (N_8854,N_8220,N_8587);
or U8855 (N_8855,N_8532,N_8149);
and U8856 (N_8856,N_8644,N_8155);
nand U8857 (N_8857,N_8219,N_8361);
or U8858 (N_8858,N_8681,N_8523);
nor U8859 (N_8859,N_8486,N_8505);
nor U8860 (N_8860,N_8524,N_8436);
and U8861 (N_8861,N_8369,N_8348);
and U8862 (N_8862,N_8471,N_8566);
nor U8863 (N_8863,N_8625,N_8322);
and U8864 (N_8864,N_8561,N_8188);
and U8865 (N_8865,N_8700,N_8372);
nand U8866 (N_8866,N_8284,N_8144);
nor U8867 (N_8867,N_8507,N_8554);
nand U8868 (N_8868,N_8380,N_8744);
or U8869 (N_8869,N_8271,N_8172);
or U8870 (N_8870,N_8329,N_8510);
nor U8871 (N_8871,N_8726,N_8285);
or U8872 (N_8872,N_8277,N_8226);
xnor U8873 (N_8873,N_8619,N_8280);
and U8874 (N_8874,N_8162,N_8295);
and U8875 (N_8875,N_8324,N_8645);
nand U8876 (N_8876,N_8208,N_8403);
nand U8877 (N_8877,N_8641,N_8230);
nand U8878 (N_8878,N_8586,N_8425);
or U8879 (N_8879,N_8199,N_8274);
nor U8880 (N_8880,N_8598,N_8255);
nor U8881 (N_8881,N_8359,N_8678);
and U8882 (N_8882,N_8689,N_8159);
nand U8883 (N_8883,N_8498,N_8235);
or U8884 (N_8884,N_8336,N_8184);
and U8885 (N_8885,N_8708,N_8579);
nand U8886 (N_8886,N_8494,N_8206);
or U8887 (N_8887,N_8431,N_8151);
nor U8888 (N_8888,N_8734,N_8653);
xor U8889 (N_8889,N_8518,N_8682);
nand U8890 (N_8890,N_8727,N_8455);
or U8891 (N_8891,N_8366,N_8368);
xnor U8892 (N_8892,N_8479,N_8262);
nor U8893 (N_8893,N_8165,N_8692);
nor U8894 (N_8894,N_8560,N_8656);
nand U8895 (N_8895,N_8450,N_8517);
or U8896 (N_8896,N_8610,N_8373);
nor U8897 (N_8897,N_8408,N_8420);
xor U8898 (N_8898,N_8259,N_8331);
or U8899 (N_8899,N_8447,N_8392);
xor U8900 (N_8900,N_8728,N_8221);
and U8901 (N_8901,N_8527,N_8558);
and U8902 (N_8902,N_8371,N_8439);
or U8903 (N_8903,N_8553,N_8407);
and U8904 (N_8904,N_8337,N_8279);
or U8905 (N_8905,N_8281,N_8215);
and U8906 (N_8906,N_8434,N_8635);
xnor U8907 (N_8907,N_8437,N_8642);
nor U8908 (N_8908,N_8181,N_8694);
or U8909 (N_8909,N_8464,N_8597);
and U8910 (N_8910,N_8630,N_8314);
nand U8911 (N_8911,N_8328,N_8268);
nand U8912 (N_8912,N_8223,N_8360);
xnor U8913 (N_8913,N_8187,N_8612);
nor U8914 (N_8914,N_8720,N_8473);
nand U8915 (N_8915,N_8263,N_8715);
nor U8916 (N_8916,N_8288,N_8589);
or U8917 (N_8917,N_8154,N_8242);
or U8918 (N_8918,N_8266,N_8717);
nand U8919 (N_8919,N_8478,N_8136);
or U8920 (N_8920,N_8356,N_8740);
nand U8921 (N_8921,N_8658,N_8730);
and U8922 (N_8922,N_8535,N_8588);
nand U8923 (N_8923,N_8676,N_8502);
nand U8924 (N_8924,N_8345,N_8352);
and U8925 (N_8925,N_8377,N_8563);
xor U8926 (N_8926,N_8704,N_8254);
or U8927 (N_8927,N_8156,N_8680);
or U8928 (N_8928,N_8634,N_8355);
and U8929 (N_8929,N_8731,N_8251);
nand U8930 (N_8930,N_8736,N_8719);
or U8931 (N_8931,N_8304,N_8148);
and U8932 (N_8932,N_8742,N_8646);
nand U8933 (N_8933,N_8241,N_8385);
or U8934 (N_8934,N_8157,N_8354);
nor U8935 (N_8935,N_8343,N_8495);
and U8936 (N_8936,N_8362,N_8186);
nor U8937 (N_8937,N_8315,N_8690);
and U8938 (N_8938,N_8591,N_8231);
or U8939 (N_8939,N_8389,N_8629);
xnor U8940 (N_8940,N_8509,N_8633);
nand U8941 (N_8941,N_8147,N_8287);
nor U8942 (N_8942,N_8444,N_8606);
nand U8943 (N_8943,N_8520,N_8664);
and U8944 (N_8944,N_8207,N_8391);
and U8945 (N_8945,N_8465,N_8195);
and U8946 (N_8946,N_8440,N_8374);
nand U8947 (N_8947,N_8243,N_8264);
xor U8948 (N_8948,N_8442,N_8536);
or U8949 (N_8949,N_8253,N_8743);
xnor U8950 (N_8950,N_8501,N_8167);
nor U8951 (N_8951,N_8513,N_8293);
nand U8952 (N_8952,N_8335,N_8216);
xnor U8953 (N_8953,N_8514,N_8239);
nand U8954 (N_8954,N_8693,N_8302);
or U8955 (N_8955,N_8364,N_8193);
and U8956 (N_8956,N_8164,N_8316);
or U8957 (N_8957,N_8204,N_8232);
nor U8958 (N_8958,N_8583,N_8522);
and U8959 (N_8959,N_8209,N_8441);
or U8960 (N_8960,N_8516,N_8555);
nor U8961 (N_8961,N_8171,N_8515);
nor U8962 (N_8962,N_8203,N_8406);
nor U8963 (N_8963,N_8497,N_8379);
or U8964 (N_8964,N_8212,N_8299);
nor U8965 (N_8965,N_8683,N_8519);
nand U8966 (N_8966,N_8415,N_8669);
nand U8967 (N_8967,N_8320,N_8210);
nand U8968 (N_8968,N_8568,N_8457);
or U8969 (N_8969,N_8225,N_8238);
and U8970 (N_8970,N_8416,N_8546);
xor U8971 (N_8971,N_8350,N_8305);
nand U8972 (N_8972,N_8126,N_8627);
nor U8973 (N_8973,N_8418,N_8668);
nor U8974 (N_8974,N_8143,N_8735);
or U8975 (N_8975,N_8135,N_8657);
and U8976 (N_8976,N_8252,N_8655);
xor U8977 (N_8977,N_8559,N_8666);
xor U8978 (N_8978,N_8378,N_8384);
nor U8979 (N_8979,N_8626,N_8248);
xor U8980 (N_8980,N_8182,N_8638);
xor U8981 (N_8981,N_8613,N_8712);
nand U8982 (N_8982,N_8405,N_8347);
and U8983 (N_8983,N_8201,N_8580);
and U8984 (N_8984,N_8468,N_8581);
nor U8985 (N_8985,N_8557,N_8260);
and U8986 (N_8986,N_8576,N_8298);
or U8987 (N_8987,N_8732,N_8466);
nand U8988 (N_8988,N_8481,N_8194);
nor U8989 (N_8989,N_8623,N_8542);
or U8990 (N_8990,N_8748,N_8341);
xor U8991 (N_8991,N_8237,N_8325);
nor U8992 (N_8992,N_8477,N_8490);
and U8993 (N_8993,N_8487,N_8339);
or U8994 (N_8994,N_8163,N_8636);
nand U8995 (N_8995,N_8430,N_8601);
and U8996 (N_8996,N_8174,N_8537);
or U8997 (N_8997,N_8585,N_8618);
nor U8998 (N_8998,N_8596,N_8723);
nand U8999 (N_8999,N_8401,N_8485);
xor U9000 (N_9000,N_8200,N_8313);
nand U9001 (N_9001,N_8538,N_8503);
nand U9002 (N_9002,N_8504,N_8317);
or U9003 (N_9003,N_8340,N_8282);
xnor U9004 (N_9004,N_8605,N_8649);
and U9005 (N_9005,N_8346,N_8521);
nand U9006 (N_9006,N_8691,N_8150);
nand U9007 (N_9007,N_8493,N_8615);
nand U9008 (N_9008,N_8616,N_8661);
xor U9009 (N_9009,N_8604,N_8614);
and U9010 (N_9010,N_8334,N_8677);
nor U9011 (N_9011,N_8449,N_8272);
and U9012 (N_9012,N_8176,N_8197);
or U9013 (N_9013,N_8296,N_8652);
xnor U9014 (N_9014,N_8697,N_8451);
or U9015 (N_9015,N_8393,N_8491);
or U9016 (N_9016,N_8413,N_8130);
or U9017 (N_9017,N_8703,N_8562);
and U9018 (N_9018,N_8291,N_8632);
nand U9019 (N_9019,N_8698,N_8443);
and U9020 (N_9020,N_8330,N_8611);
and U9021 (N_9021,N_8218,N_8236);
or U9022 (N_9022,N_8402,N_8733);
nand U9023 (N_9023,N_8617,N_8395);
nand U9024 (N_9024,N_8381,N_8175);
and U9025 (N_9025,N_8570,N_8224);
nor U9026 (N_9026,N_8390,N_8307);
nor U9027 (N_9027,N_8267,N_8575);
and U9028 (N_9028,N_8671,N_8461);
nand U9029 (N_9029,N_8318,N_8141);
and U9030 (N_9030,N_8672,N_8273);
xor U9031 (N_9031,N_8128,N_8647);
xor U9032 (N_9032,N_8548,N_8469);
xnor U9033 (N_9033,N_8138,N_8375);
or U9034 (N_9034,N_8131,N_8275);
or U9035 (N_9035,N_8483,N_8423);
and U9036 (N_9036,N_8593,N_8269);
or U9037 (N_9037,N_8396,N_8482);
or U9038 (N_9038,N_8422,N_8670);
nand U9039 (N_9039,N_8250,N_8565);
or U9040 (N_9040,N_8674,N_8725);
and U9041 (N_9041,N_8433,N_8660);
and U9042 (N_9042,N_8550,N_8249);
and U9043 (N_9043,N_8129,N_8463);
or U9044 (N_9044,N_8687,N_8140);
or U9045 (N_9045,N_8139,N_8667);
and U9046 (N_9046,N_8488,N_8244);
or U9047 (N_9047,N_8170,N_8292);
and U9048 (N_9048,N_8173,N_8737);
xnor U9049 (N_9049,N_8178,N_8294);
and U9050 (N_9050,N_8499,N_8534);
nand U9051 (N_9051,N_8312,N_8446);
and U9052 (N_9052,N_8695,N_8713);
nand U9053 (N_9053,N_8276,N_8571);
nor U9054 (N_9054,N_8637,N_8551);
nand U9055 (N_9055,N_8543,N_8665);
nand U9056 (N_9056,N_8650,N_8133);
and U9057 (N_9057,N_8410,N_8358);
nand U9058 (N_9058,N_8533,N_8370);
or U9059 (N_9059,N_8327,N_8161);
and U9060 (N_9060,N_8289,N_8344);
nand U9061 (N_9061,N_8569,N_8145);
nor U9062 (N_9062,N_8205,N_8708);
and U9063 (N_9063,N_8481,N_8177);
nor U9064 (N_9064,N_8156,N_8234);
or U9065 (N_9065,N_8513,N_8248);
and U9066 (N_9066,N_8636,N_8332);
and U9067 (N_9067,N_8667,N_8584);
nand U9068 (N_9068,N_8201,N_8502);
nor U9069 (N_9069,N_8497,N_8676);
nand U9070 (N_9070,N_8232,N_8596);
nor U9071 (N_9071,N_8615,N_8672);
nand U9072 (N_9072,N_8183,N_8421);
nor U9073 (N_9073,N_8470,N_8374);
nor U9074 (N_9074,N_8327,N_8741);
and U9075 (N_9075,N_8553,N_8294);
nand U9076 (N_9076,N_8303,N_8199);
xnor U9077 (N_9077,N_8621,N_8324);
or U9078 (N_9078,N_8305,N_8671);
nand U9079 (N_9079,N_8683,N_8559);
xnor U9080 (N_9080,N_8295,N_8358);
nor U9081 (N_9081,N_8551,N_8511);
or U9082 (N_9082,N_8235,N_8747);
nand U9083 (N_9083,N_8194,N_8276);
or U9084 (N_9084,N_8425,N_8346);
and U9085 (N_9085,N_8644,N_8191);
nor U9086 (N_9086,N_8725,N_8147);
nor U9087 (N_9087,N_8143,N_8464);
or U9088 (N_9088,N_8283,N_8492);
nor U9089 (N_9089,N_8294,N_8618);
nor U9090 (N_9090,N_8727,N_8146);
nand U9091 (N_9091,N_8548,N_8309);
nor U9092 (N_9092,N_8711,N_8459);
nor U9093 (N_9093,N_8310,N_8210);
or U9094 (N_9094,N_8545,N_8252);
or U9095 (N_9095,N_8630,N_8666);
nand U9096 (N_9096,N_8141,N_8591);
nand U9097 (N_9097,N_8171,N_8373);
or U9098 (N_9098,N_8522,N_8596);
nand U9099 (N_9099,N_8253,N_8538);
or U9100 (N_9100,N_8526,N_8564);
and U9101 (N_9101,N_8529,N_8505);
xor U9102 (N_9102,N_8589,N_8664);
nand U9103 (N_9103,N_8260,N_8510);
or U9104 (N_9104,N_8372,N_8344);
nor U9105 (N_9105,N_8275,N_8304);
nor U9106 (N_9106,N_8471,N_8505);
nand U9107 (N_9107,N_8516,N_8389);
and U9108 (N_9108,N_8707,N_8169);
nand U9109 (N_9109,N_8203,N_8459);
or U9110 (N_9110,N_8254,N_8703);
nor U9111 (N_9111,N_8508,N_8288);
and U9112 (N_9112,N_8238,N_8408);
nand U9113 (N_9113,N_8203,N_8187);
nor U9114 (N_9114,N_8581,N_8143);
and U9115 (N_9115,N_8443,N_8139);
and U9116 (N_9116,N_8473,N_8353);
or U9117 (N_9117,N_8303,N_8532);
and U9118 (N_9118,N_8514,N_8364);
or U9119 (N_9119,N_8375,N_8211);
or U9120 (N_9120,N_8490,N_8562);
nor U9121 (N_9121,N_8680,N_8139);
nor U9122 (N_9122,N_8531,N_8592);
nand U9123 (N_9123,N_8156,N_8393);
or U9124 (N_9124,N_8557,N_8425);
nor U9125 (N_9125,N_8536,N_8448);
xor U9126 (N_9126,N_8377,N_8126);
and U9127 (N_9127,N_8159,N_8697);
nand U9128 (N_9128,N_8403,N_8280);
or U9129 (N_9129,N_8145,N_8549);
nor U9130 (N_9130,N_8465,N_8574);
or U9131 (N_9131,N_8638,N_8617);
nor U9132 (N_9132,N_8687,N_8328);
and U9133 (N_9133,N_8240,N_8350);
nand U9134 (N_9134,N_8235,N_8374);
nor U9135 (N_9135,N_8322,N_8702);
or U9136 (N_9136,N_8604,N_8277);
and U9137 (N_9137,N_8132,N_8639);
and U9138 (N_9138,N_8428,N_8612);
nor U9139 (N_9139,N_8136,N_8214);
nand U9140 (N_9140,N_8738,N_8441);
nand U9141 (N_9141,N_8658,N_8483);
nor U9142 (N_9142,N_8329,N_8682);
nor U9143 (N_9143,N_8234,N_8273);
or U9144 (N_9144,N_8591,N_8610);
nor U9145 (N_9145,N_8645,N_8184);
and U9146 (N_9146,N_8453,N_8497);
nand U9147 (N_9147,N_8570,N_8365);
or U9148 (N_9148,N_8619,N_8636);
and U9149 (N_9149,N_8646,N_8354);
or U9150 (N_9150,N_8272,N_8171);
nand U9151 (N_9151,N_8212,N_8159);
nand U9152 (N_9152,N_8433,N_8454);
and U9153 (N_9153,N_8692,N_8404);
and U9154 (N_9154,N_8165,N_8490);
nand U9155 (N_9155,N_8171,N_8488);
and U9156 (N_9156,N_8454,N_8303);
or U9157 (N_9157,N_8569,N_8150);
and U9158 (N_9158,N_8617,N_8336);
nand U9159 (N_9159,N_8482,N_8730);
nor U9160 (N_9160,N_8552,N_8293);
xnor U9161 (N_9161,N_8545,N_8300);
and U9162 (N_9162,N_8501,N_8151);
or U9163 (N_9163,N_8336,N_8681);
nand U9164 (N_9164,N_8296,N_8232);
and U9165 (N_9165,N_8312,N_8541);
and U9166 (N_9166,N_8742,N_8550);
xor U9167 (N_9167,N_8271,N_8207);
and U9168 (N_9168,N_8588,N_8735);
or U9169 (N_9169,N_8200,N_8319);
and U9170 (N_9170,N_8265,N_8533);
or U9171 (N_9171,N_8334,N_8390);
xor U9172 (N_9172,N_8342,N_8284);
nor U9173 (N_9173,N_8505,N_8601);
nor U9174 (N_9174,N_8572,N_8419);
or U9175 (N_9175,N_8281,N_8259);
nor U9176 (N_9176,N_8573,N_8527);
or U9177 (N_9177,N_8191,N_8173);
nor U9178 (N_9178,N_8584,N_8307);
nor U9179 (N_9179,N_8748,N_8317);
or U9180 (N_9180,N_8129,N_8229);
nand U9181 (N_9181,N_8308,N_8632);
nand U9182 (N_9182,N_8480,N_8701);
xnor U9183 (N_9183,N_8269,N_8438);
or U9184 (N_9184,N_8164,N_8499);
or U9185 (N_9185,N_8401,N_8242);
or U9186 (N_9186,N_8470,N_8507);
and U9187 (N_9187,N_8643,N_8736);
and U9188 (N_9188,N_8228,N_8679);
nand U9189 (N_9189,N_8272,N_8346);
or U9190 (N_9190,N_8523,N_8746);
nand U9191 (N_9191,N_8543,N_8291);
nor U9192 (N_9192,N_8704,N_8236);
nand U9193 (N_9193,N_8233,N_8250);
and U9194 (N_9194,N_8586,N_8551);
and U9195 (N_9195,N_8667,N_8348);
nand U9196 (N_9196,N_8669,N_8238);
nand U9197 (N_9197,N_8595,N_8257);
and U9198 (N_9198,N_8155,N_8235);
nand U9199 (N_9199,N_8318,N_8137);
nand U9200 (N_9200,N_8270,N_8547);
nor U9201 (N_9201,N_8328,N_8499);
or U9202 (N_9202,N_8635,N_8681);
or U9203 (N_9203,N_8162,N_8158);
nor U9204 (N_9204,N_8337,N_8508);
and U9205 (N_9205,N_8149,N_8655);
nand U9206 (N_9206,N_8432,N_8333);
xnor U9207 (N_9207,N_8576,N_8442);
and U9208 (N_9208,N_8172,N_8735);
nand U9209 (N_9209,N_8448,N_8608);
nor U9210 (N_9210,N_8483,N_8574);
or U9211 (N_9211,N_8193,N_8711);
and U9212 (N_9212,N_8546,N_8314);
nor U9213 (N_9213,N_8643,N_8747);
nor U9214 (N_9214,N_8153,N_8162);
and U9215 (N_9215,N_8659,N_8374);
nand U9216 (N_9216,N_8595,N_8645);
or U9217 (N_9217,N_8411,N_8253);
nor U9218 (N_9218,N_8154,N_8410);
nor U9219 (N_9219,N_8138,N_8290);
nand U9220 (N_9220,N_8628,N_8315);
or U9221 (N_9221,N_8654,N_8576);
nor U9222 (N_9222,N_8409,N_8375);
nand U9223 (N_9223,N_8256,N_8630);
nor U9224 (N_9224,N_8141,N_8200);
nand U9225 (N_9225,N_8242,N_8402);
nor U9226 (N_9226,N_8502,N_8377);
nor U9227 (N_9227,N_8663,N_8332);
and U9228 (N_9228,N_8565,N_8661);
nand U9229 (N_9229,N_8710,N_8543);
and U9230 (N_9230,N_8618,N_8407);
nor U9231 (N_9231,N_8452,N_8531);
nand U9232 (N_9232,N_8217,N_8246);
or U9233 (N_9233,N_8572,N_8177);
xor U9234 (N_9234,N_8582,N_8383);
nor U9235 (N_9235,N_8541,N_8654);
nor U9236 (N_9236,N_8710,N_8261);
nand U9237 (N_9237,N_8225,N_8349);
or U9238 (N_9238,N_8359,N_8625);
nor U9239 (N_9239,N_8632,N_8341);
or U9240 (N_9240,N_8351,N_8349);
or U9241 (N_9241,N_8405,N_8535);
xnor U9242 (N_9242,N_8420,N_8663);
or U9243 (N_9243,N_8260,N_8342);
xor U9244 (N_9244,N_8716,N_8655);
xnor U9245 (N_9245,N_8146,N_8743);
and U9246 (N_9246,N_8622,N_8537);
nand U9247 (N_9247,N_8275,N_8319);
nor U9248 (N_9248,N_8439,N_8622);
and U9249 (N_9249,N_8142,N_8587);
and U9250 (N_9250,N_8712,N_8621);
nor U9251 (N_9251,N_8140,N_8603);
or U9252 (N_9252,N_8559,N_8526);
nor U9253 (N_9253,N_8707,N_8284);
and U9254 (N_9254,N_8577,N_8636);
nor U9255 (N_9255,N_8438,N_8239);
and U9256 (N_9256,N_8273,N_8231);
or U9257 (N_9257,N_8386,N_8667);
nand U9258 (N_9258,N_8242,N_8525);
and U9259 (N_9259,N_8451,N_8596);
nand U9260 (N_9260,N_8683,N_8552);
nand U9261 (N_9261,N_8726,N_8471);
nand U9262 (N_9262,N_8275,N_8246);
or U9263 (N_9263,N_8664,N_8542);
and U9264 (N_9264,N_8569,N_8568);
xor U9265 (N_9265,N_8413,N_8551);
xor U9266 (N_9266,N_8606,N_8306);
nor U9267 (N_9267,N_8214,N_8228);
and U9268 (N_9268,N_8528,N_8339);
and U9269 (N_9269,N_8154,N_8277);
and U9270 (N_9270,N_8344,N_8512);
and U9271 (N_9271,N_8677,N_8384);
and U9272 (N_9272,N_8646,N_8455);
nand U9273 (N_9273,N_8580,N_8354);
or U9274 (N_9274,N_8137,N_8616);
xnor U9275 (N_9275,N_8671,N_8203);
nand U9276 (N_9276,N_8169,N_8563);
nor U9277 (N_9277,N_8681,N_8685);
xnor U9278 (N_9278,N_8330,N_8631);
nor U9279 (N_9279,N_8650,N_8506);
or U9280 (N_9280,N_8405,N_8645);
nor U9281 (N_9281,N_8652,N_8745);
and U9282 (N_9282,N_8219,N_8394);
nand U9283 (N_9283,N_8662,N_8366);
and U9284 (N_9284,N_8563,N_8243);
nand U9285 (N_9285,N_8723,N_8558);
nand U9286 (N_9286,N_8343,N_8681);
and U9287 (N_9287,N_8336,N_8723);
nand U9288 (N_9288,N_8525,N_8721);
xor U9289 (N_9289,N_8442,N_8395);
nand U9290 (N_9290,N_8742,N_8521);
or U9291 (N_9291,N_8384,N_8729);
nor U9292 (N_9292,N_8609,N_8579);
and U9293 (N_9293,N_8175,N_8200);
and U9294 (N_9294,N_8721,N_8303);
nand U9295 (N_9295,N_8163,N_8558);
nand U9296 (N_9296,N_8366,N_8694);
or U9297 (N_9297,N_8213,N_8597);
and U9298 (N_9298,N_8546,N_8383);
xnor U9299 (N_9299,N_8624,N_8258);
and U9300 (N_9300,N_8352,N_8254);
nor U9301 (N_9301,N_8305,N_8417);
or U9302 (N_9302,N_8328,N_8300);
xor U9303 (N_9303,N_8519,N_8280);
xnor U9304 (N_9304,N_8416,N_8362);
nor U9305 (N_9305,N_8629,N_8523);
or U9306 (N_9306,N_8653,N_8126);
nand U9307 (N_9307,N_8694,N_8251);
or U9308 (N_9308,N_8412,N_8546);
and U9309 (N_9309,N_8618,N_8366);
and U9310 (N_9310,N_8430,N_8676);
nor U9311 (N_9311,N_8700,N_8621);
or U9312 (N_9312,N_8557,N_8673);
or U9313 (N_9313,N_8691,N_8576);
and U9314 (N_9314,N_8717,N_8599);
and U9315 (N_9315,N_8588,N_8365);
and U9316 (N_9316,N_8391,N_8698);
or U9317 (N_9317,N_8456,N_8227);
xnor U9318 (N_9318,N_8531,N_8676);
nand U9319 (N_9319,N_8472,N_8668);
or U9320 (N_9320,N_8413,N_8155);
nand U9321 (N_9321,N_8526,N_8348);
or U9322 (N_9322,N_8668,N_8290);
nand U9323 (N_9323,N_8224,N_8647);
nor U9324 (N_9324,N_8408,N_8653);
and U9325 (N_9325,N_8173,N_8697);
and U9326 (N_9326,N_8555,N_8317);
nor U9327 (N_9327,N_8703,N_8575);
or U9328 (N_9328,N_8726,N_8522);
nand U9329 (N_9329,N_8562,N_8559);
nand U9330 (N_9330,N_8332,N_8210);
nand U9331 (N_9331,N_8477,N_8471);
and U9332 (N_9332,N_8705,N_8301);
or U9333 (N_9333,N_8496,N_8498);
nor U9334 (N_9334,N_8603,N_8157);
nand U9335 (N_9335,N_8537,N_8528);
nor U9336 (N_9336,N_8502,N_8215);
xnor U9337 (N_9337,N_8642,N_8697);
nor U9338 (N_9338,N_8255,N_8446);
nor U9339 (N_9339,N_8339,N_8394);
nor U9340 (N_9340,N_8703,N_8381);
nor U9341 (N_9341,N_8300,N_8315);
nor U9342 (N_9342,N_8249,N_8657);
nor U9343 (N_9343,N_8209,N_8530);
nor U9344 (N_9344,N_8741,N_8284);
and U9345 (N_9345,N_8575,N_8589);
nand U9346 (N_9346,N_8560,N_8715);
nand U9347 (N_9347,N_8200,N_8473);
and U9348 (N_9348,N_8634,N_8465);
or U9349 (N_9349,N_8580,N_8500);
or U9350 (N_9350,N_8333,N_8327);
and U9351 (N_9351,N_8129,N_8137);
nand U9352 (N_9352,N_8357,N_8443);
or U9353 (N_9353,N_8559,N_8339);
or U9354 (N_9354,N_8405,N_8716);
xor U9355 (N_9355,N_8743,N_8243);
nand U9356 (N_9356,N_8535,N_8621);
xnor U9357 (N_9357,N_8698,N_8664);
or U9358 (N_9358,N_8135,N_8491);
xnor U9359 (N_9359,N_8425,N_8332);
nor U9360 (N_9360,N_8336,N_8249);
xor U9361 (N_9361,N_8219,N_8602);
or U9362 (N_9362,N_8210,N_8493);
and U9363 (N_9363,N_8145,N_8504);
nand U9364 (N_9364,N_8414,N_8712);
nand U9365 (N_9365,N_8488,N_8608);
or U9366 (N_9366,N_8211,N_8565);
nor U9367 (N_9367,N_8494,N_8731);
xnor U9368 (N_9368,N_8498,N_8221);
or U9369 (N_9369,N_8533,N_8595);
and U9370 (N_9370,N_8216,N_8222);
nor U9371 (N_9371,N_8128,N_8480);
and U9372 (N_9372,N_8507,N_8149);
and U9373 (N_9373,N_8663,N_8317);
and U9374 (N_9374,N_8359,N_8537);
xor U9375 (N_9375,N_9271,N_8932);
nor U9376 (N_9376,N_9213,N_8806);
and U9377 (N_9377,N_8789,N_8922);
or U9378 (N_9378,N_8909,N_8763);
or U9379 (N_9379,N_9114,N_8965);
and U9380 (N_9380,N_8813,N_8814);
and U9381 (N_9381,N_8920,N_9055);
nor U9382 (N_9382,N_8793,N_9319);
and U9383 (N_9383,N_9341,N_9149);
nor U9384 (N_9384,N_9002,N_9069);
nand U9385 (N_9385,N_8956,N_8948);
nor U9386 (N_9386,N_9192,N_8846);
or U9387 (N_9387,N_9245,N_9193);
nor U9388 (N_9388,N_9008,N_9117);
xnor U9389 (N_9389,N_9065,N_8809);
or U9390 (N_9390,N_8874,N_9130);
and U9391 (N_9391,N_8780,N_8761);
or U9392 (N_9392,N_9095,N_9359);
nor U9393 (N_9393,N_9247,N_8759);
or U9394 (N_9394,N_9040,N_8785);
and U9395 (N_9395,N_8801,N_8981);
nand U9396 (N_9396,N_9294,N_8770);
and U9397 (N_9397,N_9177,N_8990);
nand U9398 (N_9398,N_8910,N_8894);
nand U9399 (N_9399,N_8849,N_9041);
nor U9400 (N_9400,N_8861,N_9332);
nand U9401 (N_9401,N_8886,N_8876);
nand U9402 (N_9402,N_9310,N_8980);
nand U9403 (N_9403,N_9198,N_9288);
nand U9404 (N_9404,N_8805,N_9035);
and U9405 (N_9405,N_8788,N_9089);
and U9406 (N_9406,N_9141,N_9331);
nor U9407 (N_9407,N_9307,N_9034);
or U9408 (N_9408,N_8816,N_9268);
and U9409 (N_9409,N_8888,N_9273);
nor U9410 (N_9410,N_8885,N_9090);
nand U9411 (N_9411,N_9142,N_9060);
and U9412 (N_9412,N_8783,N_9074);
or U9413 (N_9413,N_9256,N_9044);
xnor U9414 (N_9414,N_9314,N_9150);
nor U9415 (N_9415,N_8891,N_9143);
nand U9416 (N_9416,N_9299,N_8945);
and U9417 (N_9417,N_8799,N_9165);
nand U9418 (N_9418,N_9099,N_9262);
nand U9419 (N_9419,N_8898,N_8796);
and U9420 (N_9420,N_9230,N_9160);
and U9421 (N_9421,N_8957,N_9364);
xor U9422 (N_9422,N_9270,N_9047);
nand U9423 (N_9423,N_9349,N_8850);
xnor U9424 (N_9424,N_9012,N_9087);
and U9425 (N_9425,N_8929,N_9077);
nand U9426 (N_9426,N_9138,N_8978);
nand U9427 (N_9427,N_9145,N_8810);
or U9428 (N_9428,N_9227,N_9258);
nor U9429 (N_9429,N_9333,N_9133);
nor U9430 (N_9430,N_8998,N_8947);
and U9431 (N_9431,N_8881,N_9123);
or U9432 (N_9432,N_9257,N_9368);
or U9433 (N_9433,N_9067,N_9309);
nor U9434 (N_9434,N_8933,N_8811);
and U9435 (N_9435,N_9315,N_9119);
or U9436 (N_9436,N_9101,N_9110);
xnor U9437 (N_9437,N_9174,N_8870);
or U9438 (N_9438,N_9023,N_9369);
nand U9439 (N_9439,N_8952,N_9269);
or U9440 (N_9440,N_9007,N_8994);
or U9441 (N_9441,N_9300,N_8988);
xnor U9442 (N_9442,N_8830,N_8837);
nand U9443 (N_9443,N_9313,N_8913);
nor U9444 (N_9444,N_9266,N_9249);
nor U9445 (N_9445,N_8977,N_9237);
nor U9446 (N_9446,N_9281,N_8890);
nor U9447 (N_9447,N_9337,N_8840);
nand U9448 (N_9448,N_8835,N_9136);
nand U9449 (N_9449,N_9267,N_8751);
or U9450 (N_9450,N_9124,N_8960);
nand U9451 (N_9451,N_9120,N_8868);
nor U9452 (N_9452,N_8872,N_9043);
or U9453 (N_9453,N_8856,N_9372);
nor U9454 (N_9454,N_9205,N_8845);
nand U9455 (N_9455,N_9081,N_9216);
xnor U9456 (N_9456,N_8962,N_8836);
or U9457 (N_9457,N_9080,N_9220);
and U9458 (N_9458,N_8865,N_9292);
and U9459 (N_9459,N_8991,N_9347);
nand U9460 (N_9460,N_9360,N_9304);
or U9461 (N_9461,N_8807,N_9062);
nor U9462 (N_9462,N_9179,N_8989);
or U9463 (N_9463,N_9021,N_9355);
or U9464 (N_9464,N_8824,N_9063);
or U9465 (N_9465,N_9203,N_9032);
and U9466 (N_9466,N_8887,N_8794);
nor U9467 (N_9467,N_9030,N_8862);
and U9468 (N_9468,N_9358,N_8867);
nand U9469 (N_9469,N_8971,N_9061);
or U9470 (N_9470,N_8982,N_9286);
nand U9471 (N_9471,N_8790,N_9056);
and U9472 (N_9472,N_9224,N_8866);
and U9473 (N_9473,N_8879,N_9251);
nor U9474 (N_9474,N_8847,N_9215);
and U9475 (N_9475,N_9340,N_8934);
or U9476 (N_9476,N_9261,N_8848);
and U9477 (N_9477,N_9017,N_9018);
or U9478 (N_9478,N_9076,N_9167);
nand U9479 (N_9479,N_9152,N_8926);
xnor U9480 (N_9480,N_9155,N_9202);
nand U9481 (N_9481,N_9161,N_8985);
nand U9482 (N_9482,N_8963,N_9362);
and U9483 (N_9483,N_9235,N_8882);
nand U9484 (N_9484,N_8765,N_9107);
and U9485 (N_9485,N_9000,N_9222);
and U9486 (N_9486,N_8827,N_9036);
or U9487 (N_9487,N_8775,N_8970);
or U9488 (N_9488,N_8939,N_8996);
nor U9489 (N_9489,N_8859,N_8976);
and U9490 (N_9490,N_9070,N_9318);
and U9491 (N_9491,N_9115,N_8777);
or U9492 (N_9492,N_8966,N_9255);
and U9493 (N_9493,N_8961,N_9186);
nor U9494 (N_9494,N_9301,N_9264);
and U9495 (N_9495,N_9113,N_9345);
nand U9496 (N_9496,N_9206,N_9118);
nand U9497 (N_9497,N_9144,N_9352);
nor U9498 (N_9498,N_8758,N_8974);
nand U9499 (N_9499,N_9293,N_8900);
and U9500 (N_9500,N_9091,N_9019);
or U9501 (N_9501,N_8906,N_8903);
and U9502 (N_9502,N_9011,N_8875);
and U9503 (N_9503,N_9045,N_9014);
nor U9504 (N_9504,N_8987,N_8917);
nand U9505 (N_9505,N_9285,N_9033);
or U9506 (N_9506,N_9151,N_8930);
or U9507 (N_9507,N_9088,N_9284);
or U9508 (N_9508,N_8787,N_9025);
nand U9509 (N_9509,N_8967,N_9325);
or U9510 (N_9510,N_8969,N_8949);
nand U9511 (N_9511,N_9001,N_8833);
nor U9512 (N_9512,N_8832,N_8858);
or U9513 (N_9513,N_9210,N_8893);
nor U9514 (N_9514,N_9280,N_9024);
nor U9515 (N_9515,N_8778,N_8774);
and U9516 (N_9516,N_8826,N_9079);
and U9517 (N_9517,N_8800,N_9243);
nand U9518 (N_9518,N_9135,N_9199);
and U9519 (N_9519,N_8973,N_9194);
and U9520 (N_9520,N_8841,N_8750);
nand U9521 (N_9521,N_8820,N_9181);
nor U9522 (N_9522,N_9189,N_8907);
and U9523 (N_9523,N_9351,N_9013);
and U9524 (N_9524,N_8822,N_8781);
nand U9525 (N_9525,N_8912,N_9201);
or U9526 (N_9526,N_9121,N_8823);
and U9527 (N_9527,N_9098,N_9291);
nand U9528 (N_9528,N_8842,N_8880);
or U9529 (N_9529,N_9365,N_9188);
and U9530 (N_9530,N_9336,N_8851);
nor U9531 (N_9531,N_9207,N_9042);
xor U9532 (N_9532,N_9038,N_9112);
nand U9533 (N_9533,N_8938,N_8899);
and U9534 (N_9534,N_8937,N_9086);
nand U9535 (N_9535,N_9197,N_9373);
and U9536 (N_9536,N_9232,N_8767);
xor U9537 (N_9537,N_9219,N_8869);
nand U9538 (N_9538,N_8828,N_9078);
nor U9539 (N_9539,N_8803,N_9240);
nor U9540 (N_9540,N_8911,N_8776);
nand U9541 (N_9541,N_9083,N_9236);
nand U9542 (N_9542,N_8935,N_8942);
nand U9543 (N_9543,N_8915,N_9354);
nand U9544 (N_9544,N_9111,N_9277);
and U9545 (N_9545,N_8769,N_9298);
nand U9546 (N_9546,N_9027,N_8863);
nand U9547 (N_9547,N_8795,N_8844);
and U9548 (N_9548,N_9330,N_9051);
or U9549 (N_9549,N_8757,N_9159);
nor U9550 (N_9550,N_8958,N_8916);
xor U9551 (N_9551,N_9005,N_9289);
xnor U9552 (N_9552,N_9191,N_9326);
or U9553 (N_9553,N_9353,N_9295);
or U9554 (N_9554,N_8755,N_8772);
or U9555 (N_9555,N_9185,N_8928);
nor U9556 (N_9556,N_9085,N_9126);
and U9557 (N_9557,N_8897,N_8895);
or U9558 (N_9558,N_9075,N_9272);
and U9559 (N_9559,N_8798,N_8908);
or U9560 (N_9560,N_9335,N_9217);
and U9561 (N_9561,N_9253,N_8838);
nor U9562 (N_9562,N_9153,N_9073);
and U9563 (N_9563,N_9239,N_8771);
or U9564 (N_9564,N_9342,N_9163);
nand U9565 (N_9565,N_8979,N_9031);
nand U9566 (N_9566,N_8839,N_8852);
and U9567 (N_9567,N_9297,N_9103);
or U9568 (N_9568,N_8764,N_9246);
xor U9569 (N_9569,N_9046,N_9172);
or U9570 (N_9570,N_9139,N_8864);
nand U9571 (N_9571,N_8878,N_8766);
nor U9572 (N_9572,N_9290,N_9148);
nor U9573 (N_9573,N_9279,N_9164);
and U9574 (N_9574,N_8901,N_9241);
nor U9575 (N_9575,N_8918,N_8786);
nor U9576 (N_9576,N_8924,N_8923);
nand U9577 (N_9577,N_8817,N_9221);
or U9578 (N_9578,N_9250,N_9020);
nor U9579 (N_9579,N_8964,N_9204);
nand U9580 (N_9580,N_9180,N_8931);
and U9581 (N_9581,N_9068,N_8992);
and U9582 (N_9582,N_8914,N_8756);
and U9583 (N_9583,N_9209,N_8940);
nor U9584 (N_9584,N_8853,N_9312);
and U9585 (N_9585,N_8802,N_9305);
nor U9586 (N_9586,N_9190,N_9134);
and U9587 (N_9587,N_8941,N_9223);
or U9588 (N_9588,N_9228,N_8904);
nand U9589 (N_9589,N_9225,N_8871);
nand U9590 (N_9590,N_9178,N_8784);
and U9591 (N_9591,N_8854,N_8925);
or U9592 (N_9592,N_9328,N_9324);
xor U9593 (N_9593,N_8762,N_9233);
or U9594 (N_9594,N_8855,N_9109);
xor U9595 (N_9595,N_9053,N_9361);
or U9596 (N_9596,N_9374,N_8773);
and U9597 (N_9597,N_8997,N_8953);
nand U9598 (N_9598,N_9003,N_9238);
or U9599 (N_9599,N_8821,N_9057);
nor U9600 (N_9600,N_8752,N_9029);
and U9601 (N_9601,N_9339,N_9367);
nand U9602 (N_9602,N_9263,N_8829);
and U9603 (N_9603,N_9321,N_9350);
nand U9604 (N_9604,N_9125,N_9175);
nand U9605 (N_9605,N_9231,N_8943);
and U9606 (N_9606,N_8843,N_8753);
nand U9607 (N_9607,N_9287,N_9183);
nor U9608 (N_9608,N_8818,N_9108);
nand U9609 (N_9609,N_9059,N_8984);
nand U9610 (N_9610,N_9212,N_9100);
nor U9611 (N_9611,N_8768,N_9218);
nor U9612 (N_9612,N_8825,N_9158);
nand U9613 (N_9613,N_9296,N_8819);
nand U9614 (N_9614,N_9173,N_8905);
nor U9615 (N_9615,N_9259,N_9327);
or U9616 (N_9616,N_9348,N_9015);
or U9617 (N_9617,N_9370,N_9275);
or U9618 (N_9618,N_9058,N_9137);
or U9619 (N_9619,N_9276,N_9343);
or U9620 (N_9620,N_8936,N_8999);
and U9621 (N_9621,N_9208,N_9322);
nand U9622 (N_9622,N_8873,N_8877);
nor U9623 (N_9623,N_9072,N_9157);
nor U9624 (N_9624,N_8782,N_9127);
nand U9625 (N_9625,N_9092,N_8995);
nand U9626 (N_9626,N_8959,N_8889);
nand U9627 (N_9627,N_8831,N_9122);
and U9628 (N_9628,N_9010,N_9363);
or U9629 (N_9629,N_9084,N_8944);
nand U9630 (N_9630,N_9054,N_8857);
and U9631 (N_9631,N_9323,N_9140);
and U9632 (N_9632,N_9316,N_8834);
nor U9633 (N_9633,N_9195,N_9156);
and U9634 (N_9634,N_9200,N_9106);
nand U9635 (N_9635,N_8950,N_9317);
nand U9636 (N_9636,N_9366,N_9039);
xor U9637 (N_9637,N_9182,N_9356);
and U9638 (N_9638,N_8792,N_8946);
or U9639 (N_9639,N_9082,N_9244);
nor U9640 (N_9640,N_8779,N_9129);
nor U9641 (N_9641,N_9128,N_9154);
and U9642 (N_9642,N_9311,N_9334);
or U9643 (N_9643,N_9283,N_8812);
xor U9644 (N_9644,N_8797,N_9096);
and U9645 (N_9645,N_8804,N_9162);
or U9646 (N_9646,N_9049,N_8815);
and U9647 (N_9647,N_8892,N_9248);
nor U9648 (N_9648,N_8883,N_9064);
nand U9649 (N_9649,N_9196,N_9097);
or U9650 (N_9650,N_9252,N_8921);
or U9651 (N_9651,N_8902,N_9306);
and U9652 (N_9652,N_9371,N_8975);
or U9653 (N_9653,N_9242,N_8896);
nor U9654 (N_9654,N_9357,N_9116);
or U9655 (N_9655,N_9176,N_9066);
or U9656 (N_9656,N_8754,N_9308);
and U9657 (N_9657,N_9226,N_8993);
nand U9658 (N_9658,N_9016,N_8884);
nor U9659 (N_9659,N_8972,N_9254);
or U9660 (N_9660,N_9009,N_9303);
or U9661 (N_9661,N_9274,N_9260);
and U9662 (N_9662,N_9320,N_9168);
nor U9663 (N_9663,N_9037,N_9234);
xor U9664 (N_9664,N_8927,N_9052);
and U9665 (N_9665,N_9170,N_9282);
xnor U9666 (N_9666,N_9302,N_8791);
nor U9667 (N_9667,N_9093,N_8919);
or U9668 (N_9668,N_9184,N_9229);
or U9669 (N_9669,N_9146,N_9171);
nand U9670 (N_9670,N_9344,N_8955);
xor U9671 (N_9671,N_9105,N_8954);
and U9672 (N_9672,N_9166,N_9048);
nand U9673 (N_9673,N_9211,N_9346);
or U9674 (N_9674,N_9187,N_9028);
nor U9675 (N_9675,N_9050,N_8760);
nor U9676 (N_9676,N_9071,N_9278);
or U9677 (N_9677,N_9214,N_9026);
or U9678 (N_9678,N_9132,N_9102);
nand U9679 (N_9679,N_9094,N_9006);
nor U9680 (N_9680,N_9147,N_8983);
nand U9681 (N_9681,N_8968,N_8808);
nand U9682 (N_9682,N_8986,N_9131);
nor U9683 (N_9683,N_9329,N_8860);
and U9684 (N_9684,N_8951,N_9338);
and U9685 (N_9685,N_9265,N_9004);
xnor U9686 (N_9686,N_9104,N_9022);
nand U9687 (N_9687,N_9169,N_8883);
and U9688 (N_9688,N_9178,N_9083);
nor U9689 (N_9689,N_8768,N_8976);
and U9690 (N_9690,N_9327,N_9278);
or U9691 (N_9691,N_8760,N_9305);
or U9692 (N_9692,N_9007,N_8894);
or U9693 (N_9693,N_9059,N_8895);
nor U9694 (N_9694,N_9168,N_9121);
or U9695 (N_9695,N_8944,N_8894);
and U9696 (N_9696,N_9167,N_9289);
xnor U9697 (N_9697,N_9197,N_8811);
or U9698 (N_9698,N_9145,N_9330);
and U9699 (N_9699,N_9013,N_9287);
nand U9700 (N_9700,N_9046,N_9335);
xor U9701 (N_9701,N_8816,N_9273);
or U9702 (N_9702,N_9064,N_8950);
xnor U9703 (N_9703,N_9011,N_9043);
nor U9704 (N_9704,N_9219,N_8970);
and U9705 (N_9705,N_8879,N_9237);
or U9706 (N_9706,N_9229,N_8757);
xor U9707 (N_9707,N_9081,N_8873);
nor U9708 (N_9708,N_8796,N_9165);
nor U9709 (N_9709,N_8913,N_9002);
and U9710 (N_9710,N_9128,N_8928);
nor U9711 (N_9711,N_8998,N_9187);
nand U9712 (N_9712,N_9066,N_9347);
nor U9713 (N_9713,N_9101,N_9300);
and U9714 (N_9714,N_9348,N_9240);
or U9715 (N_9715,N_9251,N_8821);
and U9716 (N_9716,N_9224,N_9088);
nor U9717 (N_9717,N_8907,N_9328);
nor U9718 (N_9718,N_9327,N_9249);
xnor U9719 (N_9719,N_8850,N_8834);
nand U9720 (N_9720,N_9238,N_9075);
xnor U9721 (N_9721,N_8916,N_9172);
or U9722 (N_9722,N_8931,N_9161);
or U9723 (N_9723,N_8790,N_8813);
nor U9724 (N_9724,N_9244,N_9072);
and U9725 (N_9725,N_8954,N_9299);
nand U9726 (N_9726,N_9098,N_9042);
nand U9727 (N_9727,N_9160,N_8827);
and U9728 (N_9728,N_8861,N_8953);
or U9729 (N_9729,N_9270,N_8779);
or U9730 (N_9730,N_8905,N_8777);
or U9731 (N_9731,N_8829,N_9033);
and U9732 (N_9732,N_9031,N_8846);
xnor U9733 (N_9733,N_9344,N_9145);
or U9734 (N_9734,N_9169,N_8946);
and U9735 (N_9735,N_9255,N_9139);
nand U9736 (N_9736,N_9057,N_9133);
or U9737 (N_9737,N_9161,N_8954);
and U9738 (N_9738,N_9363,N_9325);
nor U9739 (N_9739,N_8915,N_8755);
nor U9740 (N_9740,N_8917,N_9309);
nand U9741 (N_9741,N_9359,N_9174);
nand U9742 (N_9742,N_8909,N_9076);
nand U9743 (N_9743,N_9262,N_9137);
and U9744 (N_9744,N_8813,N_9103);
nor U9745 (N_9745,N_8833,N_9293);
and U9746 (N_9746,N_8847,N_9035);
xnor U9747 (N_9747,N_9046,N_9054);
or U9748 (N_9748,N_9126,N_9123);
or U9749 (N_9749,N_8984,N_9190);
or U9750 (N_9750,N_9057,N_9331);
or U9751 (N_9751,N_9019,N_9148);
nand U9752 (N_9752,N_9079,N_9142);
nand U9753 (N_9753,N_9127,N_9279);
nand U9754 (N_9754,N_9179,N_9283);
xor U9755 (N_9755,N_8961,N_9180);
and U9756 (N_9756,N_9275,N_9152);
or U9757 (N_9757,N_9259,N_9185);
nor U9758 (N_9758,N_8848,N_8785);
nor U9759 (N_9759,N_9176,N_9161);
and U9760 (N_9760,N_9277,N_9335);
and U9761 (N_9761,N_9295,N_9322);
nand U9762 (N_9762,N_8809,N_8897);
nand U9763 (N_9763,N_8789,N_8988);
xor U9764 (N_9764,N_8804,N_8884);
nor U9765 (N_9765,N_8970,N_9363);
nor U9766 (N_9766,N_9216,N_9327);
or U9767 (N_9767,N_9236,N_9086);
nand U9768 (N_9768,N_9171,N_8877);
or U9769 (N_9769,N_9249,N_9105);
or U9770 (N_9770,N_9229,N_9114);
or U9771 (N_9771,N_8800,N_9269);
nand U9772 (N_9772,N_9116,N_8866);
and U9773 (N_9773,N_8900,N_9223);
and U9774 (N_9774,N_9268,N_9287);
and U9775 (N_9775,N_8825,N_9335);
or U9776 (N_9776,N_8880,N_9132);
nand U9777 (N_9777,N_8787,N_8849);
or U9778 (N_9778,N_8851,N_9319);
xnor U9779 (N_9779,N_8891,N_9226);
and U9780 (N_9780,N_9092,N_9333);
or U9781 (N_9781,N_9314,N_9052);
and U9782 (N_9782,N_9329,N_8914);
nor U9783 (N_9783,N_9009,N_8841);
or U9784 (N_9784,N_9339,N_9039);
nor U9785 (N_9785,N_8808,N_8819);
nand U9786 (N_9786,N_8934,N_9070);
or U9787 (N_9787,N_9013,N_9054);
or U9788 (N_9788,N_9330,N_9192);
and U9789 (N_9789,N_9000,N_9232);
nor U9790 (N_9790,N_9195,N_9257);
nor U9791 (N_9791,N_8823,N_8864);
nand U9792 (N_9792,N_9186,N_9016);
nor U9793 (N_9793,N_9069,N_9163);
or U9794 (N_9794,N_8893,N_8832);
nand U9795 (N_9795,N_9046,N_9011);
xor U9796 (N_9796,N_8886,N_9076);
or U9797 (N_9797,N_9202,N_9327);
nor U9798 (N_9798,N_9372,N_9277);
xnor U9799 (N_9799,N_8802,N_8893);
and U9800 (N_9800,N_8804,N_8984);
nand U9801 (N_9801,N_9136,N_9079);
xor U9802 (N_9802,N_9096,N_9118);
and U9803 (N_9803,N_8993,N_9178);
nand U9804 (N_9804,N_8832,N_9106);
nand U9805 (N_9805,N_8827,N_9354);
nand U9806 (N_9806,N_9100,N_8838);
nand U9807 (N_9807,N_9171,N_9272);
or U9808 (N_9808,N_8812,N_8950);
and U9809 (N_9809,N_9290,N_9019);
nor U9810 (N_9810,N_9147,N_8995);
and U9811 (N_9811,N_9290,N_8959);
nor U9812 (N_9812,N_9218,N_8764);
nor U9813 (N_9813,N_9251,N_9102);
or U9814 (N_9814,N_8847,N_9367);
nand U9815 (N_9815,N_9197,N_8995);
or U9816 (N_9816,N_8941,N_8881);
xor U9817 (N_9817,N_9122,N_8822);
or U9818 (N_9818,N_9122,N_9288);
nand U9819 (N_9819,N_8829,N_9106);
nor U9820 (N_9820,N_8955,N_8873);
nor U9821 (N_9821,N_9309,N_9226);
or U9822 (N_9822,N_8837,N_8800);
nand U9823 (N_9823,N_8953,N_8787);
nor U9824 (N_9824,N_9055,N_9041);
xor U9825 (N_9825,N_9208,N_9326);
or U9826 (N_9826,N_9173,N_9010);
and U9827 (N_9827,N_8884,N_9017);
xor U9828 (N_9828,N_8865,N_8750);
and U9829 (N_9829,N_9364,N_9051);
nor U9830 (N_9830,N_9168,N_9013);
nand U9831 (N_9831,N_8774,N_8837);
nand U9832 (N_9832,N_8917,N_8998);
and U9833 (N_9833,N_9241,N_9246);
nor U9834 (N_9834,N_9333,N_8951);
nor U9835 (N_9835,N_9307,N_8863);
nand U9836 (N_9836,N_9242,N_9120);
or U9837 (N_9837,N_8781,N_9311);
nor U9838 (N_9838,N_9274,N_8910);
nand U9839 (N_9839,N_9348,N_9268);
nand U9840 (N_9840,N_9326,N_9017);
or U9841 (N_9841,N_9006,N_9007);
nor U9842 (N_9842,N_8889,N_9184);
or U9843 (N_9843,N_9208,N_9198);
xnor U9844 (N_9844,N_9242,N_9062);
nor U9845 (N_9845,N_8902,N_9086);
nor U9846 (N_9846,N_9055,N_9225);
nor U9847 (N_9847,N_9269,N_9131);
nor U9848 (N_9848,N_8827,N_9303);
or U9849 (N_9849,N_9154,N_9012);
xor U9850 (N_9850,N_9370,N_9341);
nor U9851 (N_9851,N_8797,N_8879);
and U9852 (N_9852,N_8929,N_9362);
and U9853 (N_9853,N_8921,N_8991);
xor U9854 (N_9854,N_9361,N_9080);
or U9855 (N_9855,N_8857,N_9251);
nor U9856 (N_9856,N_8756,N_8906);
xor U9857 (N_9857,N_8894,N_9289);
nor U9858 (N_9858,N_9202,N_8812);
or U9859 (N_9859,N_8975,N_9227);
or U9860 (N_9860,N_8922,N_8787);
or U9861 (N_9861,N_8785,N_8929);
nand U9862 (N_9862,N_9055,N_8872);
or U9863 (N_9863,N_9162,N_9351);
or U9864 (N_9864,N_9342,N_8985);
nand U9865 (N_9865,N_9357,N_9267);
and U9866 (N_9866,N_9225,N_9028);
nand U9867 (N_9867,N_9235,N_8887);
or U9868 (N_9868,N_8941,N_8905);
or U9869 (N_9869,N_8901,N_9330);
nor U9870 (N_9870,N_9178,N_8971);
or U9871 (N_9871,N_8829,N_9223);
or U9872 (N_9872,N_9368,N_9193);
nand U9873 (N_9873,N_9348,N_9017);
xnor U9874 (N_9874,N_8791,N_8837);
nor U9875 (N_9875,N_8959,N_9064);
xnor U9876 (N_9876,N_8932,N_9256);
and U9877 (N_9877,N_8757,N_9048);
and U9878 (N_9878,N_9025,N_9012);
or U9879 (N_9879,N_9139,N_9243);
nor U9880 (N_9880,N_8824,N_9331);
xnor U9881 (N_9881,N_9323,N_8980);
nand U9882 (N_9882,N_8774,N_9191);
nor U9883 (N_9883,N_9118,N_9164);
nor U9884 (N_9884,N_9260,N_9206);
and U9885 (N_9885,N_9308,N_8820);
nand U9886 (N_9886,N_9113,N_9081);
xnor U9887 (N_9887,N_9364,N_9274);
nand U9888 (N_9888,N_9187,N_9160);
nand U9889 (N_9889,N_9291,N_9268);
or U9890 (N_9890,N_9350,N_8890);
nor U9891 (N_9891,N_8961,N_9239);
nor U9892 (N_9892,N_9366,N_8843);
or U9893 (N_9893,N_8758,N_8988);
nand U9894 (N_9894,N_8926,N_8757);
nor U9895 (N_9895,N_8885,N_9362);
nand U9896 (N_9896,N_8780,N_9273);
or U9897 (N_9897,N_9037,N_8972);
nor U9898 (N_9898,N_9245,N_9218);
nor U9899 (N_9899,N_9202,N_8971);
nand U9900 (N_9900,N_9147,N_9037);
or U9901 (N_9901,N_9222,N_9306);
nand U9902 (N_9902,N_8823,N_8752);
nor U9903 (N_9903,N_9331,N_9228);
and U9904 (N_9904,N_8898,N_9179);
nor U9905 (N_9905,N_9260,N_9304);
nand U9906 (N_9906,N_9362,N_8892);
and U9907 (N_9907,N_8978,N_9216);
or U9908 (N_9908,N_9097,N_8851);
nand U9909 (N_9909,N_8799,N_8853);
or U9910 (N_9910,N_9293,N_9072);
nand U9911 (N_9911,N_8999,N_8956);
nor U9912 (N_9912,N_9088,N_8932);
and U9913 (N_9913,N_9360,N_9284);
xor U9914 (N_9914,N_9054,N_9348);
nand U9915 (N_9915,N_9178,N_8772);
nand U9916 (N_9916,N_8783,N_8938);
nand U9917 (N_9917,N_8975,N_8764);
or U9918 (N_9918,N_8937,N_9134);
xor U9919 (N_9919,N_9365,N_8810);
or U9920 (N_9920,N_9114,N_8946);
nand U9921 (N_9921,N_8879,N_8752);
nand U9922 (N_9922,N_8946,N_8885);
xor U9923 (N_9923,N_8778,N_9096);
xnor U9924 (N_9924,N_8981,N_8754);
nand U9925 (N_9925,N_9043,N_9245);
nand U9926 (N_9926,N_9371,N_8919);
or U9927 (N_9927,N_8784,N_8914);
and U9928 (N_9928,N_9193,N_9165);
or U9929 (N_9929,N_9348,N_9163);
and U9930 (N_9930,N_8833,N_8863);
or U9931 (N_9931,N_8971,N_9262);
nand U9932 (N_9932,N_9202,N_8775);
nand U9933 (N_9933,N_9211,N_8831);
and U9934 (N_9934,N_8973,N_9103);
and U9935 (N_9935,N_8796,N_9195);
nor U9936 (N_9936,N_8774,N_8930);
nand U9937 (N_9937,N_9309,N_9103);
or U9938 (N_9938,N_9075,N_9197);
nor U9939 (N_9939,N_9016,N_8908);
and U9940 (N_9940,N_8944,N_9245);
nor U9941 (N_9941,N_9142,N_8848);
nor U9942 (N_9942,N_8918,N_8933);
and U9943 (N_9943,N_9229,N_8932);
nand U9944 (N_9944,N_8942,N_9143);
and U9945 (N_9945,N_9172,N_9194);
and U9946 (N_9946,N_8804,N_9191);
and U9947 (N_9947,N_9315,N_8974);
or U9948 (N_9948,N_9341,N_9013);
nand U9949 (N_9949,N_9006,N_8980);
xnor U9950 (N_9950,N_9070,N_9289);
or U9951 (N_9951,N_8858,N_9180);
xor U9952 (N_9952,N_9318,N_9184);
and U9953 (N_9953,N_9025,N_9201);
nor U9954 (N_9954,N_8883,N_9047);
xor U9955 (N_9955,N_9121,N_8805);
nand U9956 (N_9956,N_8983,N_8841);
or U9957 (N_9957,N_9305,N_9212);
or U9958 (N_9958,N_9008,N_9151);
and U9959 (N_9959,N_8878,N_9287);
and U9960 (N_9960,N_9331,N_9289);
nand U9961 (N_9961,N_8797,N_8835);
and U9962 (N_9962,N_9097,N_9045);
or U9963 (N_9963,N_9297,N_9001);
and U9964 (N_9964,N_9327,N_9234);
and U9965 (N_9965,N_9124,N_8891);
xor U9966 (N_9966,N_9069,N_8942);
xor U9967 (N_9967,N_9266,N_9145);
and U9968 (N_9968,N_9291,N_8798);
or U9969 (N_9969,N_8834,N_8780);
and U9970 (N_9970,N_9295,N_9235);
or U9971 (N_9971,N_8794,N_9085);
or U9972 (N_9972,N_8884,N_8842);
nand U9973 (N_9973,N_8811,N_8770);
and U9974 (N_9974,N_8751,N_8750);
nor U9975 (N_9975,N_9143,N_9280);
nand U9976 (N_9976,N_9055,N_9372);
or U9977 (N_9977,N_9202,N_9167);
or U9978 (N_9978,N_9148,N_9036);
nor U9979 (N_9979,N_9030,N_8841);
and U9980 (N_9980,N_9289,N_9355);
and U9981 (N_9981,N_9253,N_9176);
nand U9982 (N_9982,N_9283,N_8960);
and U9983 (N_9983,N_9340,N_8952);
and U9984 (N_9984,N_9094,N_9300);
and U9985 (N_9985,N_9027,N_9153);
and U9986 (N_9986,N_9325,N_9008);
nand U9987 (N_9987,N_9013,N_8880);
or U9988 (N_9988,N_8890,N_9209);
nor U9989 (N_9989,N_8883,N_8836);
xor U9990 (N_9990,N_8765,N_9054);
nand U9991 (N_9991,N_9250,N_8838);
and U9992 (N_9992,N_8897,N_9155);
and U9993 (N_9993,N_8941,N_9012);
nor U9994 (N_9994,N_8820,N_8827);
or U9995 (N_9995,N_9115,N_8789);
nand U9996 (N_9996,N_9318,N_9095);
nor U9997 (N_9997,N_9369,N_8820);
xnor U9998 (N_9998,N_8996,N_9241);
nor U9999 (N_9999,N_9044,N_9356);
or U10000 (N_10000,N_9950,N_9517);
or U10001 (N_10001,N_9658,N_9702);
or U10002 (N_10002,N_9894,N_9890);
and U10003 (N_10003,N_9997,N_9735);
nor U10004 (N_10004,N_9657,N_9472);
nor U10005 (N_10005,N_9972,N_9577);
nor U10006 (N_10006,N_9454,N_9486);
nand U10007 (N_10007,N_9740,N_9378);
xor U10008 (N_10008,N_9551,N_9791);
nor U10009 (N_10009,N_9613,N_9408);
nand U10010 (N_10010,N_9560,N_9929);
nor U10011 (N_10011,N_9622,N_9803);
xor U10012 (N_10012,N_9700,N_9415);
nand U10013 (N_10013,N_9855,N_9970);
nor U10014 (N_10014,N_9790,N_9401);
xor U10015 (N_10015,N_9967,N_9646);
or U10016 (N_10016,N_9960,N_9532);
or U10017 (N_10017,N_9647,N_9919);
xor U10018 (N_10018,N_9417,N_9456);
nand U10019 (N_10019,N_9439,N_9769);
or U10020 (N_10020,N_9474,N_9722);
nor U10021 (N_10021,N_9597,N_9768);
or U10022 (N_10022,N_9980,N_9930);
and U10023 (N_10023,N_9839,N_9781);
nand U10024 (N_10024,N_9953,N_9822);
and U10025 (N_10025,N_9745,N_9868);
nor U10026 (N_10026,N_9631,N_9734);
and U10027 (N_10027,N_9978,N_9833);
nand U10028 (N_10028,N_9796,N_9695);
or U10029 (N_10029,N_9873,N_9874);
nor U10030 (N_10030,N_9507,N_9836);
nand U10031 (N_10031,N_9653,N_9850);
nor U10032 (N_10032,N_9393,N_9825);
and U10033 (N_10033,N_9721,N_9819);
or U10034 (N_10034,N_9608,N_9792);
xor U10035 (N_10035,N_9485,N_9901);
and U10036 (N_10036,N_9804,N_9824);
xnor U10037 (N_10037,N_9982,N_9905);
xor U10038 (N_10038,N_9893,N_9815);
nand U10039 (N_10039,N_9958,N_9459);
nand U10040 (N_10040,N_9879,N_9934);
or U10041 (N_10041,N_9420,N_9491);
or U10042 (N_10042,N_9724,N_9433);
nor U10043 (N_10043,N_9466,N_9959);
nand U10044 (N_10044,N_9998,N_9654);
or U10045 (N_10045,N_9442,N_9552);
xnor U10046 (N_10046,N_9392,N_9526);
xnor U10047 (N_10047,N_9849,N_9559);
or U10048 (N_10048,N_9891,N_9451);
or U10049 (N_10049,N_9523,N_9388);
nand U10050 (N_10050,N_9522,N_9536);
nand U10051 (N_10051,N_9616,N_9685);
and U10052 (N_10052,N_9535,N_9663);
nor U10053 (N_10053,N_9460,N_9640);
nand U10054 (N_10054,N_9828,N_9394);
xor U10055 (N_10055,N_9540,N_9587);
and U10056 (N_10056,N_9714,N_9924);
xnor U10057 (N_10057,N_9549,N_9948);
nor U10058 (N_10058,N_9962,N_9497);
nor U10059 (N_10059,N_9407,N_9773);
nor U10060 (N_10060,N_9807,N_9945);
and U10061 (N_10061,N_9519,N_9525);
nor U10062 (N_10062,N_9854,N_9410);
or U10063 (N_10063,N_9453,N_9776);
or U10064 (N_10064,N_9794,N_9397);
and U10065 (N_10065,N_9690,N_9999);
nand U10066 (N_10066,N_9539,N_9876);
or U10067 (N_10067,N_9675,N_9593);
xnor U10068 (N_10068,N_9437,N_9742);
or U10069 (N_10069,N_9676,N_9767);
nor U10070 (N_10070,N_9500,N_9949);
nor U10071 (N_10071,N_9966,N_9503);
nor U10072 (N_10072,N_9600,N_9389);
or U10073 (N_10073,N_9412,N_9431);
nor U10074 (N_10074,N_9404,N_9521);
xnor U10075 (N_10075,N_9462,N_9856);
and U10076 (N_10076,N_9859,N_9565);
nand U10077 (N_10077,N_9708,N_9886);
or U10078 (N_10078,N_9508,N_9479);
nand U10079 (N_10079,N_9902,N_9584);
nand U10080 (N_10080,N_9943,N_9892);
xnor U10081 (N_10081,N_9778,N_9384);
nand U10082 (N_10082,N_9435,N_9835);
and U10083 (N_10083,N_9968,N_9871);
xnor U10084 (N_10084,N_9994,N_9770);
nand U10085 (N_10085,N_9727,N_9779);
nor U10086 (N_10086,N_9684,N_9492);
or U10087 (N_10087,N_9862,N_9649);
nand U10088 (N_10088,N_9406,N_9940);
and U10089 (N_10089,N_9538,N_9820);
and U10090 (N_10090,N_9464,N_9562);
or U10091 (N_10091,N_9624,N_9467);
and U10092 (N_10092,N_9784,N_9841);
and U10093 (N_10093,N_9547,N_9751);
nand U10094 (N_10094,N_9422,N_9645);
or U10095 (N_10095,N_9911,N_9793);
nor U10096 (N_10096,N_9601,N_9897);
nor U10097 (N_10097,N_9711,N_9556);
or U10098 (N_10098,N_9561,N_9888);
nand U10099 (N_10099,N_9843,N_9704);
nor U10100 (N_10100,N_9444,N_9816);
and U10101 (N_10101,N_9746,N_9615);
or U10102 (N_10102,N_9964,N_9564);
nand U10103 (N_10103,N_9916,N_9910);
nor U10104 (N_10104,N_9477,N_9840);
and U10105 (N_10105,N_9754,N_9527);
and U10106 (N_10106,N_9848,N_9920);
nor U10107 (N_10107,N_9883,N_9687);
nand U10108 (N_10108,N_9917,N_9563);
and U10109 (N_10109,N_9443,N_9788);
nand U10110 (N_10110,N_9635,N_9718);
or U10111 (N_10111,N_9900,N_9634);
nand U10112 (N_10112,N_9866,N_9814);
or U10113 (N_10113,N_9733,N_9895);
or U10114 (N_10114,N_9381,N_9887);
nand U10115 (N_10115,N_9568,N_9595);
or U10116 (N_10116,N_9495,N_9937);
nand U10117 (N_10117,N_9989,N_9800);
xor U10118 (N_10118,N_9637,N_9683);
nand U10119 (N_10119,N_9400,N_9489);
nand U10120 (N_10120,N_9723,N_9992);
and U10121 (N_10121,N_9534,N_9674);
nor U10122 (N_10122,N_9611,N_9694);
nor U10123 (N_10123,N_9604,N_9743);
xnor U10124 (N_10124,N_9932,N_9870);
nand U10125 (N_10125,N_9596,N_9882);
nand U10126 (N_10126,N_9598,N_9537);
and U10127 (N_10127,N_9944,N_9529);
nor U10128 (N_10128,N_9679,N_9504);
nand U10129 (N_10129,N_9505,N_9681);
and U10130 (N_10130,N_9956,N_9402);
nand U10131 (N_10131,N_9789,N_9570);
nand U10132 (N_10132,N_9963,N_9955);
nor U10133 (N_10133,N_9682,N_9703);
nor U10134 (N_10134,N_9386,N_9864);
or U10135 (N_10135,N_9880,N_9461);
xor U10136 (N_10136,N_9627,N_9785);
nand U10137 (N_10137,N_9419,N_9603);
nor U10138 (N_10138,N_9729,N_9667);
or U10139 (N_10139,N_9558,N_9628);
or U10140 (N_10140,N_9455,N_9736);
or U10141 (N_10141,N_9512,N_9625);
nor U10142 (N_10142,N_9531,N_9403);
or U10143 (N_10143,N_9632,N_9383);
or U10144 (N_10144,N_9725,N_9445);
nor U10145 (N_10145,N_9813,N_9530);
and U10146 (N_10146,N_9590,N_9385);
nor U10147 (N_10147,N_9481,N_9990);
nand U10148 (N_10148,N_9993,N_9376);
nand U10149 (N_10149,N_9612,N_9720);
nand U10150 (N_10150,N_9837,N_9541);
nor U10151 (N_10151,N_9428,N_9669);
nand U10152 (N_10152,N_9973,N_9983);
or U10153 (N_10153,N_9728,N_9984);
or U10154 (N_10154,N_9701,N_9954);
and U10155 (N_10155,N_9639,N_9899);
or U10156 (N_10156,N_9752,N_9758);
or U10157 (N_10157,N_9626,N_9961);
or U10158 (N_10158,N_9591,N_9812);
or U10159 (N_10159,N_9971,N_9688);
nor U10160 (N_10160,N_9737,N_9851);
nand U10161 (N_10161,N_9436,N_9642);
and U10162 (N_10162,N_9847,N_9914);
nor U10163 (N_10163,N_9660,N_9429);
or U10164 (N_10164,N_9896,N_9689);
nand U10165 (N_10165,N_9898,N_9434);
and U10166 (N_10166,N_9748,N_9418);
and U10167 (N_10167,N_9757,N_9903);
or U10168 (N_10168,N_9520,N_9764);
nor U10169 (N_10169,N_9375,N_9524);
and U10170 (N_10170,N_9922,N_9926);
nor U10171 (N_10171,N_9699,N_9712);
nor U10172 (N_10172,N_9574,N_9648);
or U10173 (N_10173,N_9799,N_9448);
and U10174 (N_10174,N_9877,N_9935);
or U10175 (N_10175,N_9957,N_9923);
or U10176 (N_10176,N_9787,N_9567);
and U10177 (N_10177,N_9502,N_9450);
nor U10178 (N_10178,N_9475,N_9672);
or U10179 (N_10179,N_9831,N_9452);
nor U10180 (N_10180,N_9775,N_9875);
or U10181 (N_10181,N_9629,N_9513);
or U10182 (N_10182,N_9469,N_9952);
nand U10183 (N_10183,N_9986,N_9795);
or U10184 (N_10184,N_9878,N_9661);
or U10185 (N_10185,N_9542,N_9906);
nand U10186 (N_10186,N_9490,N_9630);
or U10187 (N_10187,N_9655,N_9947);
nor U10188 (N_10188,N_9827,N_9579);
nand U10189 (N_10189,N_9907,N_9623);
nor U10190 (N_10190,N_9426,N_9755);
and U10191 (N_10191,N_9802,N_9692);
and U10192 (N_10192,N_9446,N_9395);
nand U10193 (N_10193,N_9965,N_9582);
and U10194 (N_10194,N_9656,N_9548);
or U10195 (N_10195,N_9913,N_9636);
or U10196 (N_10196,N_9761,N_9414);
nor U10197 (N_10197,N_9697,N_9664);
xor U10198 (N_10198,N_9808,N_9942);
and U10199 (N_10199,N_9749,N_9643);
or U10200 (N_10200,N_9573,N_9921);
or U10201 (N_10201,N_9777,N_9605);
nor U10202 (N_10202,N_9763,N_9946);
and U10203 (N_10203,N_9482,N_9838);
or U10204 (N_10204,N_9380,N_9610);
nand U10205 (N_10205,N_9939,N_9713);
or U10206 (N_10206,N_9387,N_9666);
nor U10207 (N_10207,N_9470,N_9382);
nor U10208 (N_10208,N_9377,N_9543);
nand U10209 (N_10209,N_9863,N_9379);
and U10210 (N_10210,N_9438,N_9731);
nor U10211 (N_10211,N_9818,N_9915);
or U10212 (N_10212,N_9717,N_9480);
or U10213 (N_10213,N_9421,N_9979);
nor U10214 (N_10214,N_9473,N_9869);
or U10215 (N_10215,N_9976,N_9427);
and U10216 (N_10216,N_9602,N_9941);
nor U10217 (N_10217,N_9677,N_9756);
or U10218 (N_10218,N_9747,N_9908);
nor U10219 (N_10219,N_9588,N_9889);
xnor U10220 (N_10220,N_9730,N_9545);
and U10221 (N_10221,N_9498,N_9811);
nor U10222 (N_10222,N_9705,N_9586);
and U10223 (N_10223,N_9478,N_9884);
or U10224 (N_10224,N_9494,N_9912);
or U10225 (N_10225,N_9995,N_9707);
nand U10226 (N_10226,N_9652,N_9861);
nor U10227 (N_10227,N_9762,N_9578);
and U10228 (N_10228,N_9499,N_9391);
nor U10229 (N_10229,N_9798,N_9571);
nor U10230 (N_10230,N_9441,N_9390);
nor U10231 (N_10231,N_9881,N_9413);
or U10232 (N_10232,N_9846,N_9659);
or U10233 (N_10233,N_9774,N_9741);
nand U10234 (N_10234,N_9739,N_9619);
and U10235 (N_10235,N_9447,N_9987);
or U10236 (N_10236,N_9546,N_9396);
nor U10237 (N_10237,N_9671,N_9618);
nand U10238 (N_10238,N_9398,N_9693);
or U10239 (N_10239,N_9858,N_9553);
nand U10240 (N_10240,N_9511,N_9569);
nor U10241 (N_10241,N_9853,N_9715);
nor U10242 (N_10242,N_9834,N_9592);
nand U10243 (N_10243,N_9555,N_9471);
nor U10244 (N_10244,N_9969,N_9641);
and U10245 (N_10245,N_9583,N_9865);
or U10246 (N_10246,N_9449,N_9432);
nor U10247 (N_10247,N_9409,N_9440);
nor U10248 (N_10248,N_9501,N_9996);
nand U10249 (N_10249,N_9716,N_9829);
nand U10250 (N_10250,N_9585,N_9533);
and U10251 (N_10251,N_9621,N_9977);
nor U10252 (N_10252,N_9732,N_9726);
or U10253 (N_10253,N_9510,N_9801);
nand U10254 (N_10254,N_9665,N_9809);
and U10255 (N_10255,N_9744,N_9772);
and U10256 (N_10256,N_9830,N_9782);
and U10257 (N_10257,N_9430,N_9975);
and U10258 (N_10258,N_9515,N_9575);
and U10259 (N_10259,N_9668,N_9867);
or U10260 (N_10260,N_9670,N_9810);
or U10261 (N_10261,N_9780,N_9783);
nand U10262 (N_10262,N_9925,N_9416);
or U10263 (N_10263,N_9759,N_9885);
and U10264 (N_10264,N_9576,N_9857);
nor U10265 (N_10265,N_9753,N_9826);
nor U10266 (N_10266,N_9860,N_9719);
or U10267 (N_10267,N_9765,N_9918);
and U10268 (N_10268,N_9518,N_9844);
nor U10269 (N_10269,N_9845,N_9933);
or U10270 (N_10270,N_9706,N_9496);
nor U10271 (N_10271,N_9817,N_9594);
or U10272 (N_10272,N_9488,N_9806);
nand U10273 (N_10273,N_9691,N_9581);
and U10274 (N_10274,N_9617,N_9457);
nor U10275 (N_10275,N_9424,N_9673);
and U10276 (N_10276,N_9928,N_9936);
xor U10277 (N_10277,N_9938,N_9484);
and U10278 (N_10278,N_9832,N_9606);
nor U10279 (N_10279,N_9589,N_9493);
and U10280 (N_10280,N_9750,N_9738);
and U10281 (N_10281,N_9468,N_9872);
nor U10282 (N_10282,N_9516,N_9425);
and U10283 (N_10283,N_9458,N_9476);
nor U10284 (N_10284,N_9662,N_9483);
nor U10285 (N_10285,N_9686,N_9599);
nand U10286 (N_10286,N_9580,N_9985);
or U10287 (N_10287,N_9550,N_9698);
and U10288 (N_10288,N_9554,N_9696);
nand U10289 (N_10289,N_9678,N_9544);
nand U10290 (N_10290,N_9709,N_9852);
and U10291 (N_10291,N_9607,N_9644);
nand U10292 (N_10292,N_9760,N_9951);
nand U10293 (N_10293,N_9909,N_9465);
and U10294 (N_10294,N_9931,N_9710);
and U10295 (N_10295,N_9506,N_9620);
xnor U10296 (N_10296,N_9988,N_9411);
or U10297 (N_10297,N_9399,N_9633);
xor U10298 (N_10298,N_9766,N_9638);
nor U10299 (N_10299,N_9566,N_9528);
nand U10300 (N_10300,N_9974,N_9487);
nand U10301 (N_10301,N_9927,N_9771);
and U10302 (N_10302,N_9651,N_9650);
or U10303 (N_10303,N_9797,N_9805);
xnor U10304 (N_10304,N_9786,N_9981);
or U10305 (N_10305,N_9614,N_9991);
nor U10306 (N_10306,N_9904,N_9423);
nand U10307 (N_10307,N_9405,N_9463);
xnor U10308 (N_10308,N_9509,N_9823);
or U10309 (N_10309,N_9680,N_9572);
nor U10310 (N_10310,N_9557,N_9842);
nor U10311 (N_10311,N_9514,N_9609);
nand U10312 (N_10312,N_9821,N_9491);
or U10313 (N_10313,N_9923,N_9920);
nand U10314 (N_10314,N_9784,N_9515);
nor U10315 (N_10315,N_9696,N_9694);
or U10316 (N_10316,N_9674,N_9870);
or U10317 (N_10317,N_9726,N_9485);
xnor U10318 (N_10318,N_9571,N_9508);
or U10319 (N_10319,N_9944,N_9792);
nor U10320 (N_10320,N_9760,N_9566);
nor U10321 (N_10321,N_9773,N_9903);
nand U10322 (N_10322,N_9763,N_9923);
and U10323 (N_10323,N_9576,N_9867);
or U10324 (N_10324,N_9439,N_9797);
xor U10325 (N_10325,N_9495,N_9585);
and U10326 (N_10326,N_9725,N_9775);
nor U10327 (N_10327,N_9502,N_9727);
nand U10328 (N_10328,N_9669,N_9457);
nor U10329 (N_10329,N_9953,N_9870);
nor U10330 (N_10330,N_9705,N_9758);
nor U10331 (N_10331,N_9994,N_9577);
nor U10332 (N_10332,N_9471,N_9874);
nand U10333 (N_10333,N_9809,N_9528);
nand U10334 (N_10334,N_9602,N_9922);
and U10335 (N_10335,N_9461,N_9579);
nor U10336 (N_10336,N_9939,N_9606);
nand U10337 (N_10337,N_9909,N_9623);
nand U10338 (N_10338,N_9707,N_9451);
and U10339 (N_10339,N_9468,N_9733);
nand U10340 (N_10340,N_9640,N_9415);
and U10341 (N_10341,N_9960,N_9874);
xnor U10342 (N_10342,N_9525,N_9822);
nand U10343 (N_10343,N_9464,N_9512);
nand U10344 (N_10344,N_9593,N_9955);
nand U10345 (N_10345,N_9728,N_9523);
nand U10346 (N_10346,N_9979,N_9907);
nand U10347 (N_10347,N_9487,N_9779);
or U10348 (N_10348,N_9747,N_9402);
or U10349 (N_10349,N_9470,N_9608);
or U10350 (N_10350,N_9607,N_9892);
or U10351 (N_10351,N_9637,N_9615);
and U10352 (N_10352,N_9956,N_9815);
and U10353 (N_10353,N_9889,N_9557);
and U10354 (N_10354,N_9979,N_9476);
or U10355 (N_10355,N_9852,N_9870);
xor U10356 (N_10356,N_9475,N_9376);
xnor U10357 (N_10357,N_9776,N_9941);
and U10358 (N_10358,N_9986,N_9783);
or U10359 (N_10359,N_9962,N_9629);
nand U10360 (N_10360,N_9380,N_9865);
and U10361 (N_10361,N_9878,N_9879);
nand U10362 (N_10362,N_9453,N_9583);
or U10363 (N_10363,N_9512,N_9413);
nor U10364 (N_10364,N_9729,N_9419);
and U10365 (N_10365,N_9526,N_9664);
xor U10366 (N_10366,N_9779,N_9534);
or U10367 (N_10367,N_9967,N_9387);
or U10368 (N_10368,N_9403,N_9954);
nand U10369 (N_10369,N_9860,N_9657);
and U10370 (N_10370,N_9387,N_9884);
or U10371 (N_10371,N_9632,N_9873);
or U10372 (N_10372,N_9576,N_9407);
xor U10373 (N_10373,N_9630,N_9688);
nand U10374 (N_10374,N_9718,N_9763);
nand U10375 (N_10375,N_9959,N_9398);
or U10376 (N_10376,N_9681,N_9694);
or U10377 (N_10377,N_9811,N_9776);
or U10378 (N_10378,N_9722,N_9860);
nor U10379 (N_10379,N_9866,N_9512);
nand U10380 (N_10380,N_9837,N_9610);
or U10381 (N_10381,N_9414,N_9594);
and U10382 (N_10382,N_9412,N_9778);
and U10383 (N_10383,N_9529,N_9816);
nand U10384 (N_10384,N_9929,N_9621);
and U10385 (N_10385,N_9690,N_9553);
nor U10386 (N_10386,N_9498,N_9527);
and U10387 (N_10387,N_9792,N_9670);
nor U10388 (N_10388,N_9797,N_9523);
or U10389 (N_10389,N_9815,N_9393);
nor U10390 (N_10390,N_9390,N_9834);
nand U10391 (N_10391,N_9810,N_9659);
nor U10392 (N_10392,N_9862,N_9723);
and U10393 (N_10393,N_9566,N_9544);
or U10394 (N_10394,N_9493,N_9554);
xnor U10395 (N_10395,N_9685,N_9527);
nand U10396 (N_10396,N_9729,N_9654);
or U10397 (N_10397,N_9978,N_9747);
nor U10398 (N_10398,N_9886,N_9936);
and U10399 (N_10399,N_9911,N_9743);
or U10400 (N_10400,N_9888,N_9715);
and U10401 (N_10401,N_9704,N_9936);
or U10402 (N_10402,N_9422,N_9758);
nand U10403 (N_10403,N_9646,N_9845);
or U10404 (N_10404,N_9530,N_9671);
nor U10405 (N_10405,N_9473,N_9641);
or U10406 (N_10406,N_9803,N_9904);
nor U10407 (N_10407,N_9811,N_9443);
and U10408 (N_10408,N_9827,N_9591);
nand U10409 (N_10409,N_9699,N_9413);
and U10410 (N_10410,N_9414,N_9671);
or U10411 (N_10411,N_9548,N_9641);
and U10412 (N_10412,N_9401,N_9932);
and U10413 (N_10413,N_9398,N_9579);
nor U10414 (N_10414,N_9661,N_9916);
or U10415 (N_10415,N_9416,N_9498);
nor U10416 (N_10416,N_9996,N_9738);
nand U10417 (N_10417,N_9501,N_9787);
or U10418 (N_10418,N_9759,N_9679);
and U10419 (N_10419,N_9786,N_9961);
or U10420 (N_10420,N_9850,N_9405);
or U10421 (N_10421,N_9579,N_9733);
nand U10422 (N_10422,N_9867,N_9944);
nand U10423 (N_10423,N_9968,N_9548);
nor U10424 (N_10424,N_9486,N_9861);
and U10425 (N_10425,N_9461,N_9682);
nand U10426 (N_10426,N_9909,N_9550);
nor U10427 (N_10427,N_9680,N_9426);
nor U10428 (N_10428,N_9592,N_9698);
and U10429 (N_10429,N_9620,N_9966);
or U10430 (N_10430,N_9443,N_9604);
nor U10431 (N_10431,N_9843,N_9594);
nand U10432 (N_10432,N_9697,N_9786);
nor U10433 (N_10433,N_9601,N_9554);
or U10434 (N_10434,N_9861,N_9808);
or U10435 (N_10435,N_9553,N_9834);
nor U10436 (N_10436,N_9924,N_9537);
and U10437 (N_10437,N_9935,N_9773);
and U10438 (N_10438,N_9537,N_9706);
nand U10439 (N_10439,N_9911,N_9784);
nand U10440 (N_10440,N_9581,N_9667);
nand U10441 (N_10441,N_9857,N_9648);
or U10442 (N_10442,N_9415,N_9388);
and U10443 (N_10443,N_9433,N_9592);
or U10444 (N_10444,N_9563,N_9850);
and U10445 (N_10445,N_9847,N_9469);
and U10446 (N_10446,N_9770,N_9765);
nand U10447 (N_10447,N_9472,N_9735);
or U10448 (N_10448,N_9441,N_9716);
nor U10449 (N_10449,N_9902,N_9401);
nor U10450 (N_10450,N_9637,N_9961);
nand U10451 (N_10451,N_9660,N_9512);
xnor U10452 (N_10452,N_9621,N_9459);
and U10453 (N_10453,N_9949,N_9808);
nor U10454 (N_10454,N_9982,N_9929);
and U10455 (N_10455,N_9622,N_9651);
nand U10456 (N_10456,N_9486,N_9685);
nand U10457 (N_10457,N_9560,N_9652);
or U10458 (N_10458,N_9420,N_9852);
nand U10459 (N_10459,N_9908,N_9958);
nand U10460 (N_10460,N_9659,N_9486);
nand U10461 (N_10461,N_9512,N_9817);
and U10462 (N_10462,N_9429,N_9742);
and U10463 (N_10463,N_9884,N_9594);
nor U10464 (N_10464,N_9451,N_9821);
and U10465 (N_10465,N_9814,N_9587);
and U10466 (N_10466,N_9838,N_9993);
and U10467 (N_10467,N_9965,N_9943);
nor U10468 (N_10468,N_9556,N_9919);
or U10469 (N_10469,N_9512,N_9722);
or U10470 (N_10470,N_9483,N_9586);
and U10471 (N_10471,N_9784,N_9464);
nor U10472 (N_10472,N_9539,N_9545);
nor U10473 (N_10473,N_9855,N_9663);
nor U10474 (N_10474,N_9743,N_9778);
or U10475 (N_10475,N_9824,N_9868);
nor U10476 (N_10476,N_9904,N_9519);
nor U10477 (N_10477,N_9816,N_9452);
or U10478 (N_10478,N_9883,N_9770);
nor U10479 (N_10479,N_9405,N_9564);
and U10480 (N_10480,N_9808,N_9566);
nor U10481 (N_10481,N_9552,N_9758);
or U10482 (N_10482,N_9422,N_9736);
and U10483 (N_10483,N_9398,N_9479);
nor U10484 (N_10484,N_9567,N_9988);
or U10485 (N_10485,N_9421,N_9803);
and U10486 (N_10486,N_9686,N_9854);
nand U10487 (N_10487,N_9885,N_9459);
and U10488 (N_10488,N_9788,N_9719);
nand U10489 (N_10489,N_9739,N_9979);
nor U10490 (N_10490,N_9863,N_9631);
nor U10491 (N_10491,N_9877,N_9816);
nor U10492 (N_10492,N_9693,N_9484);
or U10493 (N_10493,N_9484,N_9972);
nor U10494 (N_10494,N_9750,N_9448);
nor U10495 (N_10495,N_9798,N_9727);
nor U10496 (N_10496,N_9918,N_9809);
nor U10497 (N_10497,N_9763,N_9741);
nand U10498 (N_10498,N_9666,N_9827);
and U10499 (N_10499,N_9885,N_9986);
nor U10500 (N_10500,N_9668,N_9614);
or U10501 (N_10501,N_9969,N_9468);
nor U10502 (N_10502,N_9560,N_9646);
and U10503 (N_10503,N_9900,N_9757);
nor U10504 (N_10504,N_9968,N_9855);
and U10505 (N_10505,N_9950,N_9864);
nor U10506 (N_10506,N_9571,N_9377);
or U10507 (N_10507,N_9900,N_9672);
xor U10508 (N_10508,N_9413,N_9709);
or U10509 (N_10509,N_9802,N_9549);
nor U10510 (N_10510,N_9954,N_9495);
and U10511 (N_10511,N_9865,N_9636);
nor U10512 (N_10512,N_9973,N_9376);
and U10513 (N_10513,N_9794,N_9710);
or U10514 (N_10514,N_9564,N_9804);
nor U10515 (N_10515,N_9814,N_9382);
xnor U10516 (N_10516,N_9426,N_9769);
and U10517 (N_10517,N_9686,N_9978);
and U10518 (N_10518,N_9891,N_9483);
nand U10519 (N_10519,N_9888,N_9624);
nand U10520 (N_10520,N_9436,N_9410);
xor U10521 (N_10521,N_9793,N_9978);
nand U10522 (N_10522,N_9535,N_9920);
nand U10523 (N_10523,N_9687,N_9762);
nor U10524 (N_10524,N_9633,N_9966);
and U10525 (N_10525,N_9762,N_9651);
or U10526 (N_10526,N_9954,N_9492);
and U10527 (N_10527,N_9780,N_9390);
or U10528 (N_10528,N_9822,N_9389);
or U10529 (N_10529,N_9604,N_9421);
or U10530 (N_10530,N_9738,N_9575);
nand U10531 (N_10531,N_9427,N_9567);
and U10532 (N_10532,N_9748,N_9839);
and U10533 (N_10533,N_9860,N_9948);
nand U10534 (N_10534,N_9515,N_9990);
or U10535 (N_10535,N_9565,N_9533);
and U10536 (N_10536,N_9828,N_9625);
or U10537 (N_10537,N_9615,N_9929);
nand U10538 (N_10538,N_9837,N_9592);
or U10539 (N_10539,N_9773,N_9836);
and U10540 (N_10540,N_9993,N_9624);
or U10541 (N_10541,N_9512,N_9535);
nor U10542 (N_10542,N_9730,N_9657);
nor U10543 (N_10543,N_9693,N_9979);
and U10544 (N_10544,N_9806,N_9864);
or U10545 (N_10545,N_9693,N_9825);
and U10546 (N_10546,N_9693,N_9447);
or U10547 (N_10547,N_9681,N_9959);
nand U10548 (N_10548,N_9634,N_9501);
and U10549 (N_10549,N_9738,N_9782);
and U10550 (N_10550,N_9861,N_9624);
nor U10551 (N_10551,N_9788,N_9799);
nor U10552 (N_10552,N_9424,N_9689);
nor U10553 (N_10553,N_9540,N_9390);
xor U10554 (N_10554,N_9515,N_9720);
nand U10555 (N_10555,N_9820,N_9489);
nand U10556 (N_10556,N_9916,N_9418);
and U10557 (N_10557,N_9817,N_9996);
xor U10558 (N_10558,N_9384,N_9936);
or U10559 (N_10559,N_9870,N_9767);
or U10560 (N_10560,N_9480,N_9746);
or U10561 (N_10561,N_9570,N_9904);
nand U10562 (N_10562,N_9739,N_9456);
or U10563 (N_10563,N_9817,N_9618);
and U10564 (N_10564,N_9500,N_9653);
nand U10565 (N_10565,N_9637,N_9627);
and U10566 (N_10566,N_9496,N_9648);
nor U10567 (N_10567,N_9445,N_9970);
or U10568 (N_10568,N_9498,N_9810);
nand U10569 (N_10569,N_9882,N_9412);
or U10570 (N_10570,N_9724,N_9425);
xor U10571 (N_10571,N_9648,N_9699);
nor U10572 (N_10572,N_9444,N_9612);
and U10573 (N_10573,N_9393,N_9666);
xor U10574 (N_10574,N_9466,N_9660);
or U10575 (N_10575,N_9843,N_9859);
nor U10576 (N_10576,N_9597,N_9398);
and U10577 (N_10577,N_9389,N_9854);
or U10578 (N_10578,N_9809,N_9808);
nor U10579 (N_10579,N_9475,N_9784);
or U10580 (N_10580,N_9958,N_9547);
nor U10581 (N_10581,N_9467,N_9758);
nor U10582 (N_10582,N_9431,N_9545);
nand U10583 (N_10583,N_9483,N_9620);
nor U10584 (N_10584,N_9539,N_9950);
or U10585 (N_10585,N_9687,N_9926);
xnor U10586 (N_10586,N_9536,N_9614);
and U10587 (N_10587,N_9777,N_9713);
and U10588 (N_10588,N_9806,N_9934);
nor U10589 (N_10589,N_9720,N_9451);
nand U10590 (N_10590,N_9816,N_9758);
and U10591 (N_10591,N_9866,N_9659);
or U10592 (N_10592,N_9809,N_9515);
nand U10593 (N_10593,N_9936,N_9557);
xnor U10594 (N_10594,N_9935,N_9576);
nand U10595 (N_10595,N_9918,N_9873);
or U10596 (N_10596,N_9872,N_9902);
nand U10597 (N_10597,N_9461,N_9504);
nand U10598 (N_10598,N_9687,N_9747);
and U10599 (N_10599,N_9930,N_9766);
nand U10600 (N_10600,N_9411,N_9603);
and U10601 (N_10601,N_9376,N_9817);
or U10602 (N_10602,N_9856,N_9647);
nor U10603 (N_10603,N_9834,N_9423);
and U10604 (N_10604,N_9894,N_9690);
or U10605 (N_10605,N_9557,N_9536);
nand U10606 (N_10606,N_9637,N_9784);
nor U10607 (N_10607,N_9931,N_9415);
xnor U10608 (N_10608,N_9633,N_9429);
or U10609 (N_10609,N_9560,N_9607);
nor U10610 (N_10610,N_9418,N_9493);
or U10611 (N_10611,N_9746,N_9624);
or U10612 (N_10612,N_9781,N_9624);
nand U10613 (N_10613,N_9601,N_9430);
nand U10614 (N_10614,N_9805,N_9473);
nand U10615 (N_10615,N_9787,N_9537);
or U10616 (N_10616,N_9590,N_9383);
nor U10617 (N_10617,N_9988,N_9575);
xnor U10618 (N_10618,N_9501,N_9516);
nand U10619 (N_10619,N_9382,N_9650);
nor U10620 (N_10620,N_9639,N_9396);
or U10621 (N_10621,N_9883,N_9504);
nor U10622 (N_10622,N_9385,N_9856);
or U10623 (N_10623,N_9421,N_9779);
or U10624 (N_10624,N_9980,N_9863);
nor U10625 (N_10625,N_10337,N_10156);
nand U10626 (N_10626,N_10619,N_10004);
nand U10627 (N_10627,N_10584,N_10184);
nor U10628 (N_10628,N_10226,N_10217);
nor U10629 (N_10629,N_10081,N_10115);
and U10630 (N_10630,N_10215,N_10512);
and U10631 (N_10631,N_10548,N_10363);
nand U10632 (N_10632,N_10261,N_10014);
or U10633 (N_10633,N_10154,N_10442);
nand U10634 (N_10634,N_10188,N_10069);
xnor U10635 (N_10635,N_10331,N_10136);
and U10636 (N_10636,N_10408,N_10611);
nand U10637 (N_10637,N_10364,N_10622);
nor U10638 (N_10638,N_10453,N_10600);
and U10639 (N_10639,N_10484,N_10545);
nand U10640 (N_10640,N_10507,N_10464);
nand U10641 (N_10641,N_10557,N_10320);
nor U10642 (N_10642,N_10079,N_10111);
or U10643 (N_10643,N_10509,N_10387);
nor U10644 (N_10644,N_10056,N_10492);
nor U10645 (N_10645,N_10301,N_10284);
and U10646 (N_10646,N_10050,N_10286);
or U10647 (N_10647,N_10046,N_10245);
or U10648 (N_10648,N_10202,N_10349);
nand U10649 (N_10649,N_10422,N_10103);
xor U10650 (N_10650,N_10410,N_10065);
nor U10651 (N_10651,N_10501,N_10098);
and U10652 (N_10652,N_10062,N_10610);
nor U10653 (N_10653,N_10585,N_10102);
and U10654 (N_10654,N_10414,N_10182);
or U10655 (N_10655,N_10447,N_10294);
xor U10656 (N_10656,N_10391,N_10126);
or U10657 (N_10657,N_10045,N_10469);
and U10658 (N_10658,N_10339,N_10171);
nand U10659 (N_10659,N_10093,N_10083);
nand U10660 (N_10660,N_10415,N_10236);
nand U10661 (N_10661,N_10072,N_10165);
and U10662 (N_10662,N_10299,N_10609);
and U10663 (N_10663,N_10169,N_10031);
and U10664 (N_10664,N_10411,N_10057);
and U10665 (N_10665,N_10225,N_10187);
xnor U10666 (N_10666,N_10563,N_10402);
and U10667 (N_10667,N_10445,N_10581);
or U10668 (N_10668,N_10227,N_10077);
xnor U10669 (N_10669,N_10303,N_10369);
or U10670 (N_10670,N_10597,N_10157);
nor U10671 (N_10671,N_10325,N_10434);
and U10672 (N_10672,N_10405,N_10210);
and U10673 (N_10673,N_10107,N_10515);
nand U10674 (N_10674,N_10094,N_10003);
or U10675 (N_10675,N_10592,N_10174);
or U10676 (N_10676,N_10511,N_10181);
and U10677 (N_10677,N_10234,N_10257);
and U10678 (N_10678,N_10263,N_10375);
and U10679 (N_10679,N_10139,N_10362);
or U10680 (N_10680,N_10420,N_10233);
or U10681 (N_10681,N_10209,N_10019);
nand U10682 (N_10682,N_10218,N_10617);
xnor U10683 (N_10683,N_10394,N_10016);
nor U10684 (N_10684,N_10404,N_10467);
or U10685 (N_10685,N_10444,N_10385);
nand U10686 (N_10686,N_10288,N_10354);
or U10687 (N_10687,N_10172,N_10163);
nor U10688 (N_10688,N_10043,N_10570);
or U10689 (N_10689,N_10473,N_10523);
xor U10690 (N_10690,N_10477,N_10560);
and U10691 (N_10691,N_10435,N_10238);
or U10692 (N_10692,N_10589,N_10266);
and U10693 (N_10693,N_10521,N_10092);
and U10694 (N_10694,N_10490,N_10503);
nand U10695 (N_10695,N_10471,N_10378);
or U10696 (N_10696,N_10390,N_10309);
nand U10697 (N_10697,N_10571,N_10252);
nor U10698 (N_10698,N_10265,N_10012);
or U10699 (N_10699,N_10293,N_10470);
xor U10700 (N_10700,N_10542,N_10175);
xor U10701 (N_10701,N_10430,N_10397);
nor U10702 (N_10702,N_10192,N_10432);
nand U10703 (N_10703,N_10123,N_10051);
nand U10704 (N_10704,N_10207,N_10134);
and U10705 (N_10705,N_10025,N_10601);
xnor U10706 (N_10706,N_10472,N_10335);
nand U10707 (N_10707,N_10311,N_10374);
and U10708 (N_10708,N_10168,N_10321);
nor U10709 (N_10709,N_10359,N_10119);
xor U10710 (N_10710,N_10305,N_10504);
and U10711 (N_10711,N_10147,N_10495);
or U10712 (N_10712,N_10277,N_10555);
nand U10713 (N_10713,N_10304,N_10269);
and U10714 (N_10714,N_10344,N_10044);
nand U10715 (N_10715,N_10067,N_10358);
or U10716 (N_10716,N_10070,N_10195);
or U10717 (N_10717,N_10528,N_10379);
and U10718 (N_10718,N_10275,N_10376);
and U10719 (N_10719,N_10384,N_10075);
nand U10720 (N_10720,N_10491,N_10087);
nand U10721 (N_10721,N_10440,N_10080);
nor U10722 (N_10722,N_10539,N_10010);
or U10723 (N_10723,N_10499,N_10537);
nand U10724 (N_10724,N_10149,N_10034);
and U10725 (N_10725,N_10498,N_10201);
and U10726 (N_10726,N_10148,N_10343);
xor U10727 (N_10727,N_10413,N_10302);
or U10728 (N_10728,N_10052,N_10315);
and U10729 (N_10729,N_10316,N_10439);
nand U10730 (N_10730,N_10524,N_10530);
or U10731 (N_10731,N_10232,N_10222);
xnor U10732 (N_10732,N_10108,N_10575);
nand U10733 (N_10733,N_10382,N_10566);
nand U10734 (N_10734,N_10508,N_10287);
xnor U10735 (N_10735,N_10451,N_10392);
or U10736 (N_10736,N_10536,N_10255);
xor U10737 (N_10737,N_10357,N_10582);
nand U10738 (N_10738,N_10620,N_10170);
and U10739 (N_10739,N_10086,N_10596);
nor U10740 (N_10740,N_10160,N_10099);
nand U10741 (N_10741,N_10406,N_10527);
and U10742 (N_10742,N_10254,N_10048);
nand U10743 (N_10743,N_10480,N_10036);
nor U10744 (N_10744,N_10403,N_10023);
and U10745 (N_10745,N_10438,N_10591);
nor U10746 (N_10746,N_10030,N_10476);
nand U10747 (N_10747,N_10588,N_10317);
or U10748 (N_10748,N_10289,N_10206);
nor U10749 (N_10749,N_10423,N_10334);
and U10750 (N_10750,N_10142,N_10367);
and U10751 (N_10751,N_10310,N_10214);
nor U10752 (N_10752,N_10543,N_10053);
xor U10753 (N_10753,N_10113,N_10455);
nor U10754 (N_10754,N_10264,N_10616);
and U10755 (N_10755,N_10389,N_10308);
nand U10756 (N_10756,N_10039,N_10203);
nand U10757 (N_10757,N_10475,N_10118);
and U10758 (N_10758,N_10361,N_10606);
and U10759 (N_10759,N_10505,N_10164);
nor U10760 (N_10760,N_10292,N_10493);
or U10761 (N_10761,N_10298,N_10368);
nand U10762 (N_10762,N_10055,N_10054);
or U10763 (N_10763,N_10130,N_10248);
and U10764 (N_10764,N_10431,N_10561);
or U10765 (N_10765,N_10267,N_10327);
or U10766 (N_10766,N_10541,N_10395);
nand U10767 (N_10767,N_10572,N_10027);
or U10768 (N_10768,N_10330,N_10525);
nand U10769 (N_10769,N_10351,N_10485);
or U10770 (N_10770,N_10185,N_10300);
nand U10771 (N_10771,N_10441,N_10198);
or U10772 (N_10772,N_10239,N_10017);
nor U10773 (N_10773,N_10574,N_10290);
nor U10774 (N_10774,N_10388,N_10262);
nor U10775 (N_10775,N_10338,N_10604);
xor U10776 (N_10776,N_10244,N_10373);
xor U10777 (N_10777,N_10583,N_10573);
and U10778 (N_10778,N_10285,N_10488);
and U10779 (N_10779,N_10449,N_10613);
or U10780 (N_10780,N_10409,N_10028);
nand U10781 (N_10781,N_10328,N_10450);
nand U10782 (N_10782,N_10220,N_10106);
nor U10783 (N_10783,N_10496,N_10313);
xor U10784 (N_10784,N_10460,N_10461);
or U10785 (N_10785,N_10546,N_10112);
nand U10786 (N_10786,N_10618,N_10569);
or U10787 (N_10787,N_10005,N_10173);
and U10788 (N_10788,N_10614,N_10346);
nand U10789 (N_10789,N_10319,N_10114);
xor U10790 (N_10790,N_10270,N_10249);
nand U10791 (N_10791,N_10224,N_10058);
and U10792 (N_10792,N_10006,N_10129);
and U10793 (N_10793,N_10417,N_10526);
nand U10794 (N_10794,N_10268,N_10061);
xor U10795 (N_10795,N_10347,N_10193);
nor U10796 (N_10796,N_10602,N_10448);
and U10797 (N_10797,N_10196,N_10533);
nand U10798 (N_10798,N_10011,N_10466);
nand U10799 (N_10799,N_10191,N_10159);
nand U10800 (N_10800,N_10020,N_10314);
and U10801 (N_10801,N_10326,N_10318);
and U10802 (N_10802,N_10151,N_10518);
nand U10803 (N_10803,N_10568,N_10117);
nor U10804 (N_10804,N_10009,N_10177);
nand U10805 (N_10805,N_10615,N_10135);
nand U10806 (N_10806,N_10138,N_10603);
nand U10807 (N_10807,N_10356,N_10260);
nand U10808 (N_10808,N_10026,N_10399);
nor U10809 (N_10809,N_10088,N_10340);
or U10810 (N_10810,N_10580,N_10258);
or U10811 (N_10811,N_10576,N_10183);
and U10812 (N_10812,N_10105,N_10279);
nand U10813 (N_10813,N_10153,N_10089);
and U10814 (N_10814,N_10186,N_10586);
or U10815 (N_10815,N_10221,N_10500);
and U10816 (N_10816,N_10551,N_10535);
nand U10817 (N_10817,N_10071,N_10213);
nand U10818 (N_10818,N_10137,N_10481);
or U10819 (N_10819,N_10001,N_10428);
or U10820 (N_10820,N_10018,N_10125);
nor U10821 (N_10821,N_10021,N_10110);
nand U10822 (N_10822,N_10529,N_10068);
or U10823 (N_10823,N_10295,N_10345);
or U10824 (N_10824,N_10109,N_10587);
nor U10825 (N_10825,N_10366,N_10312);
nor U10826 (N_10826,N_10540,N_10152);
nor U10827 (N_10827,N_10097,N_10324);
nor U10828 (N_10828,N_10443,N_10166);
nand U10829 (N_10829,N_10228,N_10231);
or U10830 (N_10830,N_10229,N_10256);
nor U10831 (N_10831,N_10468,N_10037);
or U10832 (N_10832,N_10066,N_10082);
nand U10833 (N_10833,N_10425,N_10063);
and U10834 (N_10834,N_10623,N_10280);
nor U10835 (N_10835,N_10281,N_10096);
and U10836 (N_10836,N_10237,N_10143);
nand U10837 (N_10837,N_10372,N_10534);
nand U10838 (N_10838,N_10246,N_10033);
and U10839 (N_10839,N_10205,N_10607);
or U10840 (N_10840,N_10038,N_10132);
and U10841 (N_10841,N_10190,N_10452);
or U10842 (N_10842,N_10155,N_10283);
nor U10843 (N_10843,N_10598,N_10296);
and U10844 (N_10844,N_10178,N_10116);
nand U10845 (N_10845,N_10241,N_10095);
nor U10846 (N_10846,N_10519,N_10352);
or U10847 (N_10847,N_10538,N_10078);
and U10848 (N_10848,N_10595,N_10380);
nand U10849 (N_10849,N_10276,N_10590);
nand U10850 (N_10850,N_10074,N_10612);
and U10851 (N_10851,N_10180,N_10424);
nor U10852 (N_10852,N_10144,N_10307);
nand U10853 (N_10853,N_10559,N_10042);
xor U10854 (N_10854,N_10336,N_10085);
nor U10855 (N_10855,N_10520,N_10024);
or U10856 (N_10856,N_10479,N_10162);
and U10857 (N_10857,N_10482,N_10446);
or U10858 (N_10858,N_10383,N_10274);
nor U10859 (N_10859,N_10032,N_10015);
or U10860 (N_10860,N_10579,N_10386);
nor U10861 (N_10861,N_10553,N_10250);
or U10862 (N_10862,N_10421,N_10407);
nor U10863 (N_10863,N_10040,N_10333);
or U10864 (N_10864,N_10341,N_10516);
nand U10865 (N_10865,N_10483,N_10002);
xnor U10866 (N_10866,N_10348,N_10532);
or U10867 (N_10867,N_10008,N_10223);
and U10868 (N_10868,N_10059,N_10377);
nor U10869 (N_10869,N_10510,N_10567);
nand U10870 (N_10870,N_10306,N_10605);
nand U10871 (N_10871,N_10454,N_10427);
or U10872 (N_10872,N_10517,N_10272);
and U10873 (N_10873,N_10122,N_10577);
and U10874 (N_10874,N_10350,N_10199);
or U10875 (N_10875,N_10370,N_10259);
or U10876 (N_10876,N_10506,N_10360);
or U10877 (N_10877,N_10329,N_10035);
nand U10878 (N_10878,N_10456,N_10041);
nor U10879 (N_10879,N_10297,N_10242);
nor U10880 (N_10880,N_10558,N_10131);
and U10881 (N_10881,N_10593,N_10127);
or U10882 (N_10882,N_10437,N_10353);
nor U10883 (N_10883,N_10278,N_10418);
nand U10884 (N_10884,N_10552,N_10502);
or U10885 (N_10885,N_10465,N_10060);
nor U10886 (N_10886,N_10578,N_10064);
or U10887 (N_10887,N_10145,N_10179);
nand U10888 (N_10888,N_10150,N_10556);
nor U10889 (N_10889,N_10489,N_10478);
nor U10890 (N_10890,N_10342,N_10121);
or U10891 (N_10891,N_10211,N_10426);
nor U10892 (N_10892,N_10522,N_10282);
or U10893 (N_10893,N_10141,N_10176);
xor U10894 (N_10894,N_10291,N_10167);
nand U10895 (N_10895,N_10084,N_10189);
or U10896 (N_10896,N_10400,N_10457);
or U10897 (N_10897,N_10158,N_10599);
and U10898 (N_10898,N_10412,N_10416);
or U10899 (N_10899,N_10251,N_10429);
or U10900 (N_10900,N_10271,N_10100);
and U10901 (N_10901,N_10513,N_10104);
nand U10902 (N_10902,N_10029,N_10544);
nor U10903 (N_10903,N_10487,N_10140);
or U10904 (N_10904,N_10076,N_10243);
nor U10905 (N_10905,N_10090,N_10419);
xnor U10906 (N_10906,N_10401,N_10549);
xnor U10907 (N_10907,N_10514,N_10000);
or U10908 (N_10908,N_10197,N_10124);
and U10909 (N_10909,N_10355,N_10101);
and U10910 (N_10910,N_10565,N_10247);
and U10911 (N_10911,N_10273,N_10494);
nor U10912 (N_10912,N_10091,N_10398);
nor U10913 (N_10913,N_10128,N_10235);
xnor U10914 (N_10914,N_10459,N_10462);
nand U10915 (N_10915,N_10073,N_10547);
and U10916 (N_10916,N_10562,N_10049);
nor U10917 (N_10917,N_10624,N_10463);
xor U10918 (N_10918,N_10322,N_10204);
and U10919 (N_10919,N_10393,N_10194);
and U10920 (N_10920,N_10120,N_10200);
or U10921 (N_10921,N_10212,N_10146);
and U10922 (N_10922,N_10486,N_10022);
nor U10923 (N_10923,N_10531,N_10608);
or U10924 (N_10924,N_10381,N_10219);
nor U10925 (N_10925,N_10013,N_10554);
nor U10926 (N_10926,N_10133,N_10550);
or U10927 (N_10927,N_10208,N_10240);
xnor U10928 (N_10928,N_10458,N_10216);
xnor U10929 (N_10929,N_10161,N_10497);
and U10930 (N_10930,N_10433,N_10230);
xor U10931 (N_10931,N_10474,N_10365);
and U10932 (N_10932,N_10621,N_10323);
or U10933 (N_10933,N_10396,N_10436);
and U10934 (N_10934,N_10253,N_10594);
nand U10935 (N_10935,N_10564,N_10371);
nor U10936 (N_10936,N_10007,N_10047);
xnor U10937 (N_10937,N_10332,N_10331);
xor U10938 (N_10938,N_10083,N_10213);
nand U10939 (N_10939,N_10540,N_10459);
and U10940 (N_10940,N_10356,N_10202);
nor U10941 (N_10941,N_10119,N_10132);
nand U10942 (N_10942,N_10256,N_10086);
nor U10943 (N_10943,N_10083,N_10024);
and U10944 (N_10944,N_10567,N_10533);
nor U10945 (N_10945,N_10219,N_10128);
and U10946 (N_10946,N_10330,N_10238);
and U10947 (N_10947,N_10218,N_10147);
xor U10948 (N_10948,N_10425,N_10041);
nor U10949 (N_10949,N_10213,N_10485);
nor U10950 (N_10950,N_10437,N_10081);
and U10951 (N_10951,N_10256,N_10187);
nand U10952 (N_10952,N_10039,N_10393);
or U10953 (N_10953,N_10020,N_10053);
and U10954 (N_10954,N_10471,N_10466);
or U10955 (N_10955,N_10485,N_10118);
xnor U10956 (N_10956,N_10599,N_10131);
and U10957 (N_10957,N_10198,N_10359);
nand U10958 (N_10958,N_10273,N_10555);
or U10959 (N_10959,N_10158,N_10004);
nor U10960 (N_10960,N_10361,N_10507);
or U10961 (N_10961,N_10058,N_10558);
nand U10962 (N_10962,N_10590,N_10293);
and U10963 (N_10963,N_10347,N_10600);
nor U10964 (N_10964,N_10507,N_10248);
nand U10965 (N_10965,N_10216,N_10046);
nand U10966 (N_10966,N_10209,N_10433);
nor U10967 (N_10967,N_10133,N_10156);
xnor U10968 (N_10968,N_10000,N_10240);
xor U10969 (N_10969,N_10170,N_10496);
xnor U10970 (N_10970,N_10350,N_10017);
nor U10971 (N_10971,N_10068,N_10185);
nand U10972 (N_10972,N_10330,N_10353);
xnor U10973 (N_10973,N_10100,N_10469);
nor U10974 (N_10974,N_10134,N_10192);
xnor U10975 (N_10975,N_10201,N_10513);
nand U10976 (N_10976,N_10351,N_10583);
and U10977 (N_10977,N_10367,N_10049);
and U10978 (N_10978,N_10029,N_10215);
xnor U10979 (N_10979,N_10282,N_10275);
xor U10980 (N_10980,N_10579,N_10116);
or U10981 (N_10981,N_10329,N_10454);
nand U10982 (N_10982,N_10541,N_10523);
or U10983 (N_10983,N_10329,N_10379);
nand U10984 (N_10984,N_10578,N_10147);
or U10985 (N_10985,N_10585,N_10583);
and U10986 (N_10986,N_10520,N_10173);
and U10987 (N_10987,N_10243,N_10390);
nor U10988 (N_10988,N_10171,N_10123);
xnor U10989 (N_10989,N_10009,N_10318);
nor U10990 (N_10990,N_10073,N_10455);
or U10991 (N_10991,N_10537,N_10005);
xnor U10992 (N_10992,N_10367,N_10101);
xnor U10993 (N_10993,N_10552,N_10493);
xnor U10994 (N_10994,N_10299,N_10375);
or U10995 (N_10995,N_10260,N_10083);
nand U10996 (N_10996,N_10579,N_10155);
and U10997 (N_10997,N_10176,N_10227);
or U10998 (N_10998,N_10375,N_10168);
or U10999 (N_10999,N_10573,N_10466);
or U11000 (N_11000,N_10248,N_10317);
or U11001 (N_11001,N_10466,N_10369);
nor U11002 (N_11002,N_10134,N_10406);
xor U11003 (N_11003,N_10532,N_10356);
nand U11004 (N_11004,N_10275,N_10208);
and U11005 (N_11005,N_10221,N_10048);
nor U11006 (N_11006,N_10123,N_10486);
nor U11007 (N_11007,N_10299,N_10246);
or U11008 (N_11008,N_10266,N_10516);
nand U11009 (N_11009,N_10413,N_10612);
nand U11010 (N_11010,N_10528,N_10485);
nand U11011 (N_11011,N_10003,N_10077);
nand U11012 (N_11012,N_10327,N_10395);
and U11013 (N_11013,N_10128,N_10426);
nand U11014 (N_11014,N_10361,N_10436);
nand U11015 (N_11015,N_10288,N_10215);
or U11016 (N_11016,N_10538,N_10442);
and U11017 (N_11017,N_10534,N_10303);
and U11018 (N_11018,N_10459,N_10294);
and U11019 (N_11019,N_10347,N_10461);
or U11020 (N_11020,N_10583,N_10611);
nand U11021 (N_11021,N_10120,N_10610);
nor U11022 (N_11022,N_10067,N_10066);
xor U11023 (N_11023,N_10009,N_10106);
and U11024 (N_11024,N_10241,N_10480);
nor U11025 (N_11025,N_10136,N_10237);
nor U11026 (N_11026,N_10176,N_10242);
and U11027 (N_11027,N_10326,N_10153);
nor U11028 (N_11028,N_10114,N_10224);
or U11029 (N_11029,N_10544,N_10052);
nor U11030 (N_11030,N_10244,N_10232);
xnor U11031 (N_11031,N_10205,N_10540);
or U11032 (N_11032,N_10349,N_10087);
and U11033 (N_11033,N_10038,N_10349);
nand U11034 (N_11034,N_10178,N_10262);
nand U11035 (N_11035,N_10186,N_10263);
nor U11036 (N_11036,N_10483,N_10168);
and U11037 (N_11037,N_10006,N_10208);
or U11038 (N_11038,N_10029,N_10420);
nor U11039 (N_11039,N_10066,N_10493);
nand U11040 (N_11040,N_10560,N_10259);
or U11041 (N_11041,N_10522,N_10341);
nand U11042 (N_11042,N_10086,N_10388);
nor U11043 (N_11043,N_10101,N_10437);
and U11044 (N_11044,N_10574,N_10365);
nand U11045 (N_11045,N_10163,N_10607);
nor U11046 (N_11046,N_10378,N_10178);
nor U11047 (N_11047,N_10138,N_10214);
nor U11048 (N_11048,N_10110,N_10415);
and U11049 (N_11049,N_10606,N_10036);
nand U11050 (N_11050,N_10293,N_10519);
nand U11051 (N_11051,N_10610,N_10244);
or U11052 (N_11052,N_10401,N_10094);
nor U11053 (N_11053,N_10144,N_10261);
nor U11054 (N_11054,N_10230,N_10455);
and U11055 (N_11055,N_10595,N_10501);
xnor U11056 (N_11056,N_10451,N_10161);
nor U11057 (N_11057,N_10492,N_10139);
and U11058 (N_11058,N_10100,N_10506);
nand U11059 (N_11059,N_10560,N_10293);
or U11060 (N_11060,N_10516,N_10053);
nor U11061 (N_11061,N_10528,N_10365);
nor U11062 (N_11062,N_10261,N_10420);
xor U11063 (N_11063,N_10227,N_10229);
nand U11064 (N_11064,N_10203,N_10572);
nor U11065 (N_11065,N_10291,N_10136);
or U11066 (N_11066,N_10086,N_10029);
xor U11067 (N_11067,N_10103,N_10034);
nor U11068 (N_11068,N_10549,N_10009);
xnor U11069 (N_11069,N_10277,N_10511);
xnor U11070 (N_11070,N_10164,N_10180);
or U11071 (N_11071,N_10555,N_10602);
and U11072 (N_11072,N_10196,N_10034);
nor U11073 (N_11073,N_10535,N_10446);
nand U11074 (N_11074,N_10466,N_10576);
or U11075 (N_11075,N_10296,N_10286);
nor U11076 (N_11076,N_10254,N_10093);
and U11077 (N_11077,N_10234,N_10378);
or U11078 (N_11078,N_10606,N_10230);
nor U11079 (N_11079,N_10255,N_10597);
nand U11080 (N_11080,N_10152,N_10436);
nor U11081 (N_11081,N_10465,N_10207);
nand U11082 (N_11082,N_10291,N_10250);
nor U11083 (N_11083,N_10368,N_10048);
nor U11084 (N_11084,N_10610,N_10011);
nor U11085 (N_11085,N_10324,N_10279);
and U11086 (N_11086,N_10603,N_10393);
nand U11087 (N_11087,N_10525,N_10138);
nor U11088 (N_11088,N_10298,N_10055);
nor U11089 (N_11089,N_10438,N_10200);
and U11090 (N_11090,N_10082,N_10276);
nand U11091 (N_11091,N_10088,N_10470);
nand U11092 (N_11092,N_10359,N_10138);
nor U11093 (N_11093,N_10386,N_10033);
nand U11094 (N_11094,N_10434,N_10541);
nor U11095 (N_11095,N_10270,N_10083);
nand U11096 (N_11096,N_10245,N_10586);
nor U11097 (N_11097,N_10386,N_10507);
nand U11098 (N_11098,N_10590,N_10185);
and U11099 (N_11099,N_10505,N_10479);
xnor U11100 (N_11100,N_10376,N_10271);
nand U11101 (N_11101,N_10027,N_10154);
nand U11102 (N_11102,N_10340,N_10215);
or U11103 (N_11103,N_10566,N_10500);
nand U11104 (N_11104,N_10522,N_10144);
nor U11105 (N_11105,N_10010,N_10576);
and U11106 (N_11106,N_10173,N_10261);
nand U11107 (N_11107,N_10162,N_10315);
and U11108 (N_11108,N_10124,N_10260);
nand U11109 (N_11109,N_10527,N_10084);
and U11110 (N_11110,N_10487,N_10563);
xnor U11111 (N_11111,N_10542,N_10477);
nor U11112 (N_11112,N_10182,N_10355);
nor U11113 (N_11113,N_10129,N_10067);
or U11114 (N_11114,N_10483,N_10491);
nor U11115 (N_11115,N_10007,N_10387);
nand U11116 (N_11116,N_10484,N_10389);
or U11117 (N_11117,N_10000,N_10017);
nor U11118 (N_11118,N_10221,N_10180);
or U11119 (N_11119,N_10528,N_10533);
and U11120 (N_11120,N_10275,N_10256);
and U11121 (N_11121,N_10249,N_10387);
nor U11122 (N_11122,N_10111,N_10320);
and U11123 (N_11123,N_10294,N_10402);
or U11124 (N_11124,N_10471,N_10358);
or U11125 (N_11125,N_10412,N_10521);
or U11126 (N_11126,N_10220,N_10623);
nor U11127 (N_11127,N_10046,N_10550);
nor U11128 (N_11128,N_10529,N_10463);
and U11129 (N_11129,N_10397,N_10147);
or U11130 (N_11130,N_10186,N_10447);
nor U11131 (N_11131,N_10355,N_10320);
and U11132 (N_11132,N_10304,N_10077);
xor U11133 (N_11133,N_10083,N_10140);
nor U11134 (N_11134,N_10375,N_10526);
xnor U11135 (N_11135,N_10097,N_10445);
nand U11136 (N_11136,N_10429,N_10557);
nor U11137 (N_11137,N_10533,N_10606);
or U11138 (N_11138,N_10062,N_10161);
xor U11139 (N_11139,N_10224,N_10593);
nand U11140 (N_11140,N_10021,N_10350);
nand U11141 (N_11141,N_10209,N_10385);
nor U11142 (N_11142,N_10129,N_10179);
nor U11143 (N_11143,N_10447,N_10030);
and U11144 (N_11144,N_10426,N_10467);
nand U11145 (N_11145,N_10541,N_10514);
and U11146 (N_11146,N_10037,N_10081);
nor U11147 (N_11147,N_10178,N_10182);
nor U11148 (N_11148,N_10319,N_10312);
nor U11149 (N_11149,N_10389,N_10375);
nor U11150 (N_11150,N_10260,N_10111);
or U11151 (N_11151,N_10489,N_10407);
nand U11152 (N_11152,N_10293,N_10004);
nand U11153 (N_11153,N_10245,N_10047);
or U11154 (N_11154,N_10087,N_10100);
nand U11155 (N_11155,N_10351,N_10507);
and U11156 (N_11156,N_10157,N_10154);
nor U11157 (N_11157,N_10291,N_10173);
xnor U11158 (N_11158,N_10337,N_10181);
xnor U11159 (N_11159,N_10065,N_10288);
nand U11160 (N_11160,N_10522,N_10115);
nand U11161 (N_11161,N_10068,N_10338);
or U11162 (N_11162,N_10567,N_10031);
or U11163 (N_11163,N_10525,N_10570);
nor U11164 (N_11164,N_10035,N_10179);
and U11165 (N_11165,N_10301,N_10113);
and U11166 (N_11166,N_10046,N_10558);
and U11167 (N_11167,N_10254,N_10252);
and U11168 (N_11168,N_10104,N_10113);
nand U11169 (N_11169,N_10566,N_10419);
and U11170 (N_11170,N_10259,N_10497);
and U11171 (N_11171,N_10174,N_10589);
or U11172 (N_11172,N_10427,N_10041);
nand U11173 (N_11173,N_10274,N_10130);
nand U11174 (N_11174,N_10254,N_10277);
nor U11175 (N_11175,N_10020,N_10315);
and U11176 (N_11176,N_10383,N_10155);
or U11177 (N_11177,N_10050,N_10153);
nor U11178 (N_11178,N_10360,N_10179);
nor U11179 (N_11179,N_10376,N_10339);
or U11180 (N_11180,N_10496,N_10295);
xor U11181 (N_11181,N_10368,N_10424);
xor U11182 (N_11182,N_10228,N_10201);
xor U11183 (N_11183,N_10215,N_10473);
nor U11184 (N_11184,N_10321,N_10420);
or U11185 (N_11185,N_10434,N_10483);
nor U11186 (N_11186,N_10474,N_10312);
nand U11187 (N_11187,N_10258,N_10377);
and U11188 (N_11188,N_10587,N_10277);
nor U11189 (N_11189,N_10236,N_10118);
nand U11190 (N_11190,N_10541,N_10613);
nor U11191 (N_11191,N_10427,N_10036);
xnor U11192 (N_11192,N_10550,N_10075);
nor U11193 (N_11193,N_10413,N_10229);
xor U11194 (N_11194,N_10497,N_10457);
or U11195 (N_11195,N_10520,N_10010);
nor U11196 (N_11196,N_10528,N_10396);
and U11197 (N_11197,N_10242,N_10000);
nand U11198 (N_11198,N_10537,N_10032);
and U11199 (N_11199,N_10279,N_10357);
or U11200 (N_11200,N_10548,N_10503);
or U11201 (N_11201,N_10334,N_10489);
xnor U11202 (N_11202,N_10000,N_10511);
nand U11203 (N_11203,N_10120,N_10250);
and U11204 (N_11204,N_10408,N_10454);
and U11205 (N_11205,N_10306,N_10554);
and U11206 (N_11206,N_10263,N_10162);
xnor U11207 (N_11207,N_10617,N_10141);
nand U11208 (N_11208,N_10274,N_10225);
or U11209 (N_11209,N_10590,N_10209);
xor U11210 (N_11210,N_10370,N_10267);
nand U11211 (N_11211,N_10149,N_10394);
and U11212 (N_11212,N_10385,N_10461);
nand U11213 (N_11213,N_10578,N_10305);
nand U11214 (N_11214,N_10447,N_10014);
nand U11215 (N_11215,N_10395,N_10169);
and U11216 (N_11216,N_10167,N_10467);
or U11217 (N_11217,N_10553,N_10485);
nor U11218 (N_11218,N_10165,N_10018);
or U11219 (N_11219,N_10526,N_10466);
or U11220 (N_11220,N_10238,N_10068);
nand U11221 (N_11221,N_10231,N_10230);
and U11222 (N_11222,N_10362,N_10452);
or U11223 (N_11223,N_10214,N_10272);
nand U11224 (N_11224,N_10350,N_10165);
xnor U11225 (N_11225,N_10122,N_10206);
or U11226 (N_11226,N_10066,N_10540);
and U11227 (N_11227,N_10579,N_10499);
xnor U11228 (N_11228,N_10397,N_10132);
nor U11229 (N_11229,N_10162,N_10179);
nor U11230 (N_11230,N_10368,N_10596);
and U11231 (N_11231,N_10177,N_10349);
nor U11232 (N_11232,N_10060,N_10618);
and U11233 (N_11233,N_10476,N_10247);
and U11234 (N_11234,N_10611,N_10318);
or U11235 (N_11235,N_10053,N_10357);
nor U11236 (N_11236,N_10412,N_10143);
nand U11237 (N_11237,N_10348,N_10323);
nor U11238 (N_11238,N_10543,N_10068);
and U11239 (N_11239,N_10360,N_10171);
nor U11240 (N_11240,N_10595,N_10351);
nor U11241 (N_11241,N_10281,N_10301);
or U11242 (N_11242,N_10119,N_10252);
and U11243 (N_11243,N_10160,N_10492);
and U11244 (N_11244,N_10340,N_10099);
xor U11245 (N_11245,N_10326,N_10613);
and U11246 (N_11246,N_10037,N_10547);
or U11247 (N_11247,N_10057,N_10131);
nand U11248 (N_11248,N_10241,N_10304);
and U11249 (N_11249,N_10424,N_10105);
or U11250 (N_11250,N_11169,N_10971);
and U11251 (N_11251,N_11181,N_10640);
and U11252 (N_11252,N_11249,N_10933);
and U11253 (N_11253,N_11224,N_11212);
nor U11254 (N_11254,N_11242,N_11168);
or U11255 (N_11255,N_11209,N_10848);
xnor U11256 (N_11256,N_10880,N_10730);
and U11257 (N_11257,N_10712,N_10901);
nor U11258 (N_11258,N_11077,N_10815);
xor U11259 (N_11259,N_11115,N_10791);
nand U11260 (N_11260,N_10708,N_11175);
or U11261 (N_11261,N_11172,N_10960);
and U11262 (N_11262,N_10654,N_11014);
nor U11263 (N_11263,N_11098,N_11106);
and U11264 (N_11264,N_10914,N_10800);
nand U11265 (N_11265,N_10842,N_10784);
nand U11266 (N_11266,N_11017,N_11201);
or U11267 (N_11267,N_10911,N_10824);
nor U11268 (N_11268,N_11157,N_10736);
nor U11269 (N_11269,N_10707,N_10838);
xor U11270 (N_11270,N_10790,N_10811);
or U11271 (N_11271,N_11192,N_10644);
and U11272 (N_11272,N_10785,N_10775);
and U11273 (N_11273,N_10667,N_10752);
nor U11274 (N_11274,N_10856,N_10998);
nor U11275 (N_11275,N_10836,N_10809);
nand U11276 (N_11276,N_10695,N_10897);
nor U11277 (N_11277,N_10637,N_10955);
nand U11278 (N_11278,N_11103,N_10686);
nand U11279 (N_11279,N_10777,N_10858);
xor U11280 (N_11280,N_11178,N_11237);
or U11281 (N_11281,N_11033,N_10700);
and U11282 (N_11282,N_10680,N_10756);
nand U11283 (N_11283,N_10761,N_10731);
and U11284 (N_11284,N_10670,N_10857);
nor U11285 (N_11285,N_11185,N_10678);
and U11286 (N_11286,N_10814,N_10884);
nand U11287 (N_11287,N_11117,N_10662);
nor U11288 (N_11288,N_11223,N_10930);
xor U11289 (N_11289,N_11045,N_10772);
nand U11290 (N_11290,N_11174,N_10816);
and U11291 (N_11291,N_10821,N_10636);
and U11292 (N_11292,N_10988,N_11068);
and U11293 (N_11293,N_11005,N_10905);
nand U11294 (N_11294,N_10656,N_10675);
nor U11295 (N_11295,N_11134,N_10684);
nand U11296 (N_11296,N_10668,N_10826);
nand U11297 (N_11297,N_11198,N_11111);
nand U11298 (N_11298,N_11137,N_10889);
xor U11299 (N_11299,N_11167,N_11161);
xnor U11300 (N_11300,N_10688,N_10628);
nor U11301 (N_11301,N_11021,N_11200);
nor U11302 (N_11302,N_11015,N_10883);
and U11303 (N_11303,N_11081,N_11136);
nand U11304 (N_11304,N_11009,N_10788);
nor U11305 (N_11305,N_10633,N_11228);
nand U11306 (N_11306,N_11022,N_11207);
xor U11307 (N_11307,N_11101,N_10794);
and U11308 (N_11308,N_10732,N_10839);
nand U11309 (N_11309,N_11218,N_11058);
nor U11310 (N_11310,N_11165,N_10725);
and U11311 (N_11311,N_11202,N_10854);
nor U11312 (N_11312,N_10750,N_10822);
or U11313 (N_11313,N_10912,N_10807);
xor U11314 (N_11314,N_11247,N_11113);
and U11315 (N_11315,N_11144,N_10647);
and U11316 (N_11316,N_10990,N_10944);
and U11317 (N_11317,N_11231,N_10724);
nand U11318 (N_11318,N_10710,N_11196);
and U11319 (N_11319,N_11019,N_10849);
nand U11320 (N_11320,N_11076,N_11075);
or U11321 (N_11321,N_10954,N_11149);
and U11322 (N_11322,N_11065,N_10973);
and U11323 (N_11323,N_10949,N_11164);
nor U11324 (N_11324,N_10748,N_11159);
and U11325 (N_11325,N_11063,N_11160);
and U11326 (N_11326,N_11083,N_10653);
nand U11327 (N_11327,N_11084,N_10735);
and U11328 (N_11328,N_10673,N_10650);
nand U11329 (N_11329,N_10845,N_10904);
or U11330 (N_11330,N_10760,N_11107);
or U11331 (N_11331,N_10886,N_10629);
nor U11332 (N_11332,N_10950,N_11069);
or U11333 (N_11333,N_10694,N_10701);
or U11334 (N_11334,N_11012,N_10726);
nand U11335 (N_11335,N_11238,N_10728);
nand U11336 (N_11336,N_10702,N_10658);
nor U11337 (N_11337,N_10632,N_10691);
nor U11338 (N_11338,N_11131,N_10820);
nor U11339 (N_11339,N_11124,N_10803);
or U11340 (N_11340,N_10698,N_11094);
xor U11341 (N_11341,N_11085,N_11186);
nor U11342 (N_11342,N_10676,N_10948);
and U11343 (N_11343,N_11146,N_10720);
nor U11344 (N_11344,N_11156,N_10639);
xnor U11345 (N_11345,N_10672,N_11116);
nand U11346 (N_11346,N_10934,N_11195);
nand U11347 (N_11347,N_10951,N_11214);
nor U11348 (N_11348,N_10837,N_10751);
or U11349 (N_11349,N_10817,N_10829);
nand U11350 (N_11350,N_11206,N_11010);
nor U11351 (N_11351,N_10742,N_11204);
xnor U11352 (N_11352,N_10903,N_10825);
nand U11353 (N_11353,N_11229,N_10759);
nand U11354 (N_11354,N_10733,N_10850);
and U11355 (N_11355,N_10655,N_11064);
nand U11356 (N_11356,N_10860,N_10652);
and U11357 (N_11357,N_10866,N_11138);
xnor U11358 (N_11358,N_11087,N_11180);
nor U11359 (N_11359,N_10873,N_11034);
and U11360 (N_11360,N_11147,N_10746);
or U11361 (N_11361,N_10771,N_10666);
xnor U11362 (N_11362,N_11028,N_10669);
nand U11363 (N_11363,N_11176,N_10718);
nor U11364 (N_11364,N_10875,N_11199);
xnor U11365 (N_11365,N_11143,N_11150);
nand U11366 (N_11366,N_10919,N_10705);
xor U11367 (N_11367,N_11193,N_11004);
and U11368 (N_11368,N_10872,N_10876);
nand U11369 (N_11369,N_10709,N_10677);
or U11370 (N_11370,N_11226,N_11213);
nor U11371 (N_11371,N_11197,N_10774);
and U11372 (N_11372,N_11114,N_10645);
and U11373 (N_11373,N_11244,N_10982);
and U11374 (N_11374,N_11050,N_10687);
nand U11375 (N_11375,N_11091,N_10643);
nor U11376 (N_11376,N_10964,N_10841);
nand U11377 (N_11377,N_11099,N_10874);
and U11378 (N_11378,N_10810,N_11062);
and U11379 (N_11379,N_10766,N_10734);
nand U11380 (N_11380,N_11179,N_10943);
or U11381 (N_11381,N_10781,N_10945);
nor U11382 (N_11382,N_11024,N_11188);
nor U11383 (N_11383,N_10987,N_10906);
nor U11384 (N_11384,N_10974,N_10902);
xor U11385 (N_11385,N_11027,N_10681);
nand U11386 (N_11386,N_10717,N_10986);
or U11387 (N_11387,N_10635,N_11026);
and U11388 (N_11388,N_10855,N_10900);
xor U11389 (N_11389,N_10755,N_10864);
nor U11390 (N_11390,N_10882,N_10690);
nand U11391 (N_11391,N_10992,N_11108);
nor U11392 (N_11392,N_10846,N_10721);
xor U11393 (N_11393,N_10868,N_11217);
nor U11394 (N_11394,N_10630,N_10641);
nand U11395 (N_11395,N_11073,N_10932);
and U11396 (N_11396,N_10852,N_11215);
or U11397 (N_11397,N_10835,N_11040);
xor U11398 (N_11398,N_10898,N_10862);
nand U11399 (N_11399,N_10685,N_10867);
nor U11400 (N_11400,N_10881,N_10744);
nor U11401 (N_11401,N_11233,N_10719);
xnor U11402 (N_11402,N_10834,N_10989);
or U11403 (N_11403,N_10741,N_10887);
nor U11404 (N_11404,N_10661,N_11007);
nand U11405 (N_11405,N_10963,N_11049);
nand U11406 (N_11406,N_11070,N_10967);
nor U11407 (N_11407,N_10722,N_11236);
or U11408 (N_11408,N_10830,N_10715);
and U11409 (N_11409,N_10778,N_10793);
nor U11410 (N_11410,N_11052,N_10627);
and U11411 (N_11411,N_10847,N_10958);
nor U11412 (N_11412,N_11235,N_10940);
nand U11413 (N_11413,N_11125,N_10657);
nand U11414 (N_11414,N_10663,N_10659);
nor U11415 (N_11415,N_11000,N_11151);
or U11416 (N_11416,N_10828,N_10928);
xnor U11417 (N_11417,N_10994,N_10783);
or U11418 (N_11418,N_10798,N_10851);
and U11419 (N_11419,N_10697,N_10865);
or U11420 (N_11420,N_10863,N_10878);
or U11421 (N_11421,N_11030,N_10767);
nor U11422 (N_11422,N_11042,N_11239);
nor U11423 (N_11423,N_10885,N_10787);
or U11424 (N_11424,N_11142,N_10626);
xnor U11425 (N_11425,N_11211,N_11055);
nor U11426 (N_11426,N_10981,N_11182);
or U11427 (N_11427,N_10634,N_10923);
and U11428 (N_11428,N_11126,N_10983);
nor U11429 (N_11429,N_10980,N_10764);
nand U11430 (N_11430,N_11123,N_10638);
nand U11431 (N_11431,N_10713,N_10704);
nand U11432 (N_11432,N_11232,N_11047);
nand U11433 (N_11433,N_11067,N_11153);
and U11434 (N_11434,N_10966,N_10985);
or U11435 (N_11435,N_11095,N_10765);
nor U11436 (N_11436,N_11121,N_10913);
nor U11437 (N_11437,N_10792,N_10871);
nand U11438 (N_11438,N_10796,N_11219);
or U11439 (N_11439,N_10740,N_11130);
xnor U11440 (N_11440,N_11139,N_10795);
and U11441 (N_11441,N_10780,N_11170);
and U11442 (N_11442,N_11129,N_10674);
nor U11443 (N_11443,N_10642,N_10808);
nand U11444 (N_11444,N_11002,N_11035);
nor U11445 (N_11445,N_11023,N_10819);
nor U11446 (N_11446,N_10925,N_11003);
and U11447 (N_11447,N_11020,N_11135);
nand U11448 (N_11448,N_10893,N_11194);
xor U11449 (N_11449,N_11145,N_10916);
nor U11450 (N_11450,N_11205,N_10693);
and U11451 (N_11451,N_11248,N_10679);
xor U11452 (N_11452,N_10692,N_11088);
nand U11453 (N_11453,N_11006,N_11241);
nor U11454 (N_11454,N_10786,N_10976);
and U11455 (N_11455,N_10706,N_10696);
and U11456 (N_11456,N_10975,N_10869);
xnor U11457 (N_11457,N_10776,N_10757);
or U11458 (N_11458,N_10918,N_11025);
nand U11459 (N_11459,N_11041,N_11054);
and U11460 (N_11460,N_10861,N_11029);
nor U11461 (N_11461,N_11013,N_10888);
and U11462 (N_11462,N_10961,N_10813);
xnor U11463 (N_11463,N_10631,N_10683);
and U11464 (N_11464,N_10921,N_11148);
nor U11465 (N_11465,N_11122,N_11246);
nand U11466 (N_11466,N_11191,N_10799);
nand U11467 (N_11467,N_10664,N_10859);
nand U11468 (N_11468,N_11066,N_11105);
or U11469 (N_11469,N_10779,N_10969);
nor U11470 (N_11470,N_10823,N_10953);
nand U11471 (N_11471,N_10754,N_11089);
nor U11472 (N_11472,N_10927,N_10952);
nand U11473 (N_11473,N_10625,N_11184);
nor U11474 (N_11474,N_11187,N_10716);
xor U11475 (N_11475,N_11039,N_10737);
or U11476 (N_11476,N_10753,N_10711);
nand U11477 (N_11477,N_10999,N_10995);
xnor U11478 (N_11478,N_10763,N_11018);
nor U11479 (N_11479,N_10832,N_10979);
and U11480 (N_11480,N_11234,N_11109);
or U11481 (N_11481,N_11220,N_10942);
or U11482 (N_11482,N_10649,N_11080);
or U11483 (N_11483,N_11189,N_10915);
and U11484 (N_11484,N_11036,N_10833);
or U11485 (N_11485,N_10939,N_10965);
and U11486 (N_11486,N_11078,N_11163);
and U11487 (N_11487,N_10896,N_10745);
and U11488 (N_11488,N_11093,N_10827);
or U11489 (N_11489,N_11128,N_11120);
and U11490 (N_11490,N_11037,N_11221);
xor U11491 (N_11491,N_11031,N_10671);
nand U11492 (N_11492,N_11210,N_11059);
nor U11493 (N_11493,N_11071,N_10773);
nor U11494 (N_11494,N_10899,N_10972);
nor U11495 (N_11495,N_11177,N_11008);
or U11496 (N_11496,N_10970,N_10879);
or U11497 (N_11497,N_10747,N_11051);
nor U11498 (N_11498,N_11046,N_11072);
or U11499 (N_11499,N_10908,N_10937);
nor U11500 (N_11500,N_11227,N_11141);
nand U11501 (N_11501,N_10959,N_11102);
xnor U11502 (N_11502,N_10714,N_10907);
xnor U11503 (N_11503,N_11011,N_10891);
nand U11504 (N_11504,N_10922,N_10910);
and U11505 (N_11505,N_10660,N_11090);
nand U11506 (N_11506,N_10931,N_11243);
xnor U11507 (N_11507,N_11016,N_11057);
nand U11508 (N_11508,N_10789,N_10739);
nand U11509 (N_11509,N_10895,N_11082);
and U11510 (N_11510,N_10993,N_11171);
nor U11511 (N_11511,N_11060,N_11096);
or U11512 (N_11512,N_10743,N_10727);
and U11513 (N_11513,N_11092,N_10917);
or U11514 (N_11514,N_10996,N_10812);
and U11515 (N_11515,N_11043,N_11166);
or U11516 (N_11516,N_10646,N_10729);
nand U11517 (N_11517,N_10804,N_10997);
xor U11518 (N_11518,N_11240,N_10769);
xnor U11519 (N_11519,N_10762,N_10818);
xor U11520 (N_11520,N_10877,N_10749);
or U11521 (N_11521,N_10797,N_10894);
nor U11522 (N_11522,N_11110,N_10723);
nor U11523 (N_11523,N_11162,N_10651);
nor U11524 (N_11524,N_11086,N_11001);
and U11525 (N_11525,N_10978,N_11152);
nand U11526 (N_11526,N_11053,N_11158);
nor U11527 (N_11527,N_11203,N_11183);
and U11528 (N_11528,N_10689,N_11154);
or U11529 (N_11529,N_11112,N_10956);
or U11530 (N_11530,N_10840,N_11119);
nor U11531 (N_11531,N_10768,N_10892);
or U11532 (N_11532,N_11155,N_10968);
nor U11533 (N_11533,N_10844,N_10782);
and U11534 (N_11534,N_11132,N_10738);
nand U11535 (N_11535,N_11038,N_11173);
xnor U11536 (N_11536,N_10890,N_11032);
and U11537 (N_11537,N_10831,N_10991);
and U11538 (N_11538,N_10957,N_10665);
nand U11539 (N_11539,N_11118,N_10929);
nor U11540 (N_11540,N_10682,N_10843);
nor U11541 (N_11541,N_11079,N_10648);
and U11542 (N_11542,N_11056,N_10853);
nand U11543 (N_11543,N_11074,N_10870);
nand U11544 (N_11544,N_10936,N_11230);
nor U11545 (N_11545,N_10758,N_10938);
or U11546 (N_11546,N_10941,N_10935);
and U11547 (N_11547,N_11140,N_10924);
or U11548 (N_11548,N_11208,N_11048);
xnor U11549 (N_11549,N_11127,N_11216);
nand U11550 (N_11550,N_10920,N_10962);
nand U11551 (N_11551,N_10703,N_11104);
nand U11552 (N_11552,N_10802,N_10806);
nand U11553 (N_11553,N_11190,N_10801);
and U11554 (N_11554,N_11133,N_10770);
and U11555 (N_11555,N_10699,N_11222);
nor U11556 (N_11556,N_11061,N_11097);
nand U11557 (N_11557,N_11100,N_10946);
and U11558 (N_11558,N_11225,N_11044);
or U11559 (N_11559,N_11245,N_10909);
nor U11560 (N_11560,N_10947,N_10984);
or U11561 (N_11561,N_10805,N_10926);
xor U11562 (N_11562,N_10977,N_11072);
nand U11563 (N_11563,N_10966,N_10634);
and U11564 (N_11564,N_10638,N_10830);
nor U11565 (N_11565,N_10899,N_10821);
xnor U11566 (N_11566,N_10659,N_11096);
or U11567 (N_11567,N_10946,N_10713);
or U11568 (N_11568,N_11125,N_10972);
or U11569 (N_11569,N_10953,N_10826);
nand U11570 (N_11570,N_10984,N_10671);
or U11571 (N_11571,N_10814,N_10859);
nor U11572 (N_11572,N_10953,N_10930);
or U11573 (N_11573,N_10698,N_11237);
nor U11574 (N_11574,N_10740,N_10637);
or U11575 (N_11575,N_10715,N_10784);
and U11576 (N_11576,N_10890,N_11204);
nand U11577 (N_11577,N_10973,N_11109);
nand U11578 (N_11578,N_11061,N_10996);
or U11579 (N_11579,N_11076,N_10977);
nor U11580 (N_11580,N_10731,N_11165);
nor U11581 (N_11581,N_11248,N_10819);
and U11582 (N_11582,N_11205,N_11232);
nand U11583 (N_11583,N_10756,N_11028);
xnor U11584 (N_11584,N_10743,N_10676);
nor U11585 (N_11585,N_10715,N_10964);
nor U11586 (N_11586,N_10801,N_10885);
or U11587 (N_11587,N_10881,N_11142);
xnor U11588 (N_11588,N_11168,N_11059);
nor U11589 (N_11589,N_10639,N_10732);
and U11590 (N_11590,N_10868,N_11204);
nor U11591 (N_11591,N_10957,N_10871);
xor U11592 (N_11592,N_11083,N_11075);
and U11593 (N_11593,N_10938,N_10648);
nor U11594 (N_11594,N_10688,N_11209);
nand U11595 (N_11595,N_10781,N_11219);
nor U11596 (N_11596,N_11205,N_10759);
nor U11597 (N_11597,N_10625,N_11215);
or U11598 (N_11598,N_11239,N_10815);
and U11599 (N_11599,N_11211,N_10946);
nor U11600 (N_11600,N_10740,N_10909);
or U11601 (N_11601,N_11165,N_11153);
nor U11602 (N_11602,N_10686,N_10790);
and U11603 (N_11603,N_10862,N_10809);
nor U11604 (N_11604,N_10849,N_11203);
and U11605 (N_11605,N_10968,N_10668);
nand U11606 (N_11606,N_10722,N_11140);
nand U11607 (N_11607,N_10854,N_11065);
and U11608 (N_11608,N_10777,N_11002);
nand U11609 (N_11609,N_10810,N_10978);
and U11610 (N_11610,N_11230,N_10754);
nor U11611 (N_11611,N_11224,N_11080);
nor U11612 (N_11612,N_10974,N_11246);
or U11613 (N_11613,N_10808,N_10877);
xor U11614 (N_11614,N_10761,N_10962);
nand U11615 (N_11615,N_10857,N_11047);
and U11616 (N_11616,N_10880,N_11152);
or U11617 (N_11617,N_10967,N_11153);
and U11618 (N_11618,N_10677,N_10818);
and U11619 (N_11619,N_10731,N_10920);
nand U11620 (N_11620,N_11226,N_11243);
nor U11621 (N_11621,N_10894,N_10779);
or U11622 (N_11622,N_11184,N_10753);
and U11623 (N_11623,N_10663,N_11039);
xor U11624 (N_11624,N_10772,N_11206);
and U11625 (N_11625,N_11209,N_11173);
nor U11626 (N_11626,N_11212,N_11249);
or U11627 (N_11627,N_10841,N_11216);
nand U11628 (N_11628,N_10629,N_11194);
and U11629 (N_11629,N_11072,N_10843);
and U11630 (N_11630,N_10643,N_11108);
nand U11631 (N_11631,N_10822,N_10962);
and U11632 (N_11632,N_10929,N_11214);
nor U11633 (N_11633,N_10887,N_10974);
or U11634 (N_11634,N_10743,N_10736);
nor U11635 (N_11635,N_10737,N_10913);
or U11636 (N_11636,N_11149,N_10928);
or U11637 (N_11637,N_11174,N_11191);
xnor U11638 (N_11638,N_10930,N_10867);
and U11639 (N_11639,N_11241,N_11054);
nor U11640 (N_11640,N_11225,N_10647);
or U11641 (N_11641,N_11034,N_10745);
nand U11642 (N_11642,N_10973,N_10990);
nand U11643 (N_11643,N_10885,N_11130);
nand U11644 (N_11644,N_11177,N_10641);
or U11645 (N_11645,N_10851,N_10970);
or U11646 (N_11646,N_10641,N_10792);
or U11647 (N_11647,N_10851,N_11008);
or U11648 (N_11648,N_11179,N_10840);
nand U11649 (N_11649,N_11049,N_10937);
and U11650 (N_11650,N_11155,N_11022);
or U11651 (N_11651,N_11009,N_10685);
or U11652 (N_11652,N_10639,N_10946);
and U11653 (N_11653,N_10741,N_10971);
nor U11654 (N_11654,N_10867,N_11051);
nor U11655 (N_11655,N_11151,N_10950);
nor U11656 (N_11656,N_11161,N_10992);
nand U11657 (N_11657,N_11224,N_10699);
and U11658 (N_11658,N_10999,N_11186);
nand U11659 (N_11659,N_11000,N_11005);
and U11660 (N_11660,N_11034,N_10664);
and U11661 (N_11661,N_10874,N_10640);
nand U11662 (N_11662,N_11116,N_10767);
xnor U11663 (N_11663,N_10853,N_10899);
and U11664 (N_11664,N_10999,N_11214);
nor U11665 (N_11665,N_11002,N_11082);
xor U11666 (N_11666,N_10829,N_11223);
nor U11667 (N_11667,N_10957,N_11106);
nor U11668 (N_11668,N_10853,N_11004);
nand U11669 (N_11669,N_11147,N_11068);
and U11670 (N_11670,N_10828,N_10705);
nor U11671 (N_11671,N_11059,N_10835);
and U11672 (N_11672,N_10635,N_10955);
nand U11673 (N_11673,N_10769,N_10899);
or U11674 (N_11674,N_10662,N_10969);
nand U11675 (N_11675,N_11004,N_10912);
nand U11676 (N_11676,N_10880,N_11088);
xor U11677 (N_11677,N_10763,N_10860);
nand U11678 (N_11678,N_11165,N_11015);
or U11679 (N_11679,N_11127,N_10743);
xor U11680 (N_11680,N_10898,N_11169);
nor U11681 (N_11681,N_11093,N_10944);
and U11682 (N_11682,N_10784,N_10819);
xnor U11683 (N_11683,N_11191,N_10759);
nand U11684 (N_11684,N_11164,N_10668);
and U11685 (N_11685,N_10797,N_11166);
or U11686 (N_11686,N_11039,N_10865);
or U11687 (N_11687,N_11161,N_10861);
nand U11688 (N_11688,N_10921,N_10891);
nand U11689 (N_11689,N_11147,N_11132);
nor U11690 (N_11690,N_11088,N_11097);
or U11691 (N_11691,N_10925,N_10710);
or U11692 (N_11692,N_10994,N_11179);
and U11693 (N_11693,N_11087,N_10747);
or U11694 (N_11694,N_10846,N_10763);
nand U11695 (N_11695,N_10969,N_11094);
or U11696 (N_11696,N_11139,N_10816);
nor U11697 (N_11697,N_11211,N_10978);
nor U11698 (N_11698,N_11151,N_11063);
and U11699 (N_11699,N_10855,N_11050);
nor U11700 (N_11700,N_11021,N_10834);
nor U11701 (N_11701,N_10871,N_10714);
nor U11702 (N_11702,N_10709,N_10883);
nand U11703 (N_11703,N_11163,N_11002);
and U11704 (N_11704,N_11188,N_10667);
nand U11705 (N_11705,N_10846,N_10958);
nand U11706 (N_11706,N_11071,N_10877);
nor U11707 (N_11707,N_10701,N_11135);
or U11708 (N_11708,N_10924,N_10742);
nor U11709 (N_11709,N_10740,N_10888);
and U11710 (N_11710,N_10921,N_11224);
nor U11711 (N_11711,N_10680,N_10778);
or U11712 (N_11712,N_10880,N_10977);
and U11713 (N_11713,N_11099,N_11120);
nand U11714 (N_11714,N_11226,N_10784);
nand U11715 (N_11715,N_10852,N_10821);
and U11716 (N_11716,N_11197,N_10785);
xor U11717 (N_11717,N_10691,N_11063);
or U11718 (N_11718,N_10689,N_10758);
nand U11719 (N_11719,N_10676,N_11208);
nor U11720 (N_11720,N_10893,N_10768);
and U11721 (N_11721,N_11013,N_11240);
or U11722 (N_11722,N_11219,N_10841);
and U11723 (N_11723,N_11008,N_10630);
or U11724 (N_11724,N_11160,N_10786);
and U11725 (N_11725,N_11114,N_10849);
or U11726 (N_11726,N_10980,N_10859);
nor U11727 (N_11727,N_11181,N_10744);
nand U11728 (N_11728,N_11086,N_10757);
nor U11729 (N_11729,N_10637,N_11094);
and U11730 (N_11730,N_10739,N_11078);
or U11731 (N_11731,N_11160,N_10782);
or U11732 (N_11732,N_10975,N_11199);
or U11733 (N_11733,N_10696,N_11009);
nor U11734 (N_11734,N_10791,N_11025);
or U11735 (N_11735,N_10807,N_11176);
and U11736 (N_11736,N_11198,N_10745);
nand U11737 (N_11737,N_10693,N_10647);
or U11738 (N_11738,N_10788,N_10702);
and U11739 (N_11739,N_10646,N_10971);
and U11740 (N_11740,N_10925,N_11083);
or U11741 (N_11741,N_11049,N_10930);
or U11742 (N_11742,N_11087,N_10754);
nor U11743 (N_11743,N_10900,N_11086);
nand U11744 (N_11744,N_10917,N_11059);
or U11745 (N_11745,N_10955,N_10826);
xor U11746 (N_11746,N_10830,N_11143);
nor U11747 (N_11747,N_10677,N_10701);
nand U11748 (N_11748,N_10952,N_10795);
xnor U11749 (N_11749,N_11247,N_10637);
and U11750 (N_11750,N_11187,N_11186);
nor U11751 (N_11751,N_11080,N_11217);
xor U11752 (N_11752,N_10879,N_11158);
nand U11753 (N_11753,N_11030,N_10843);
and U11754 (N_11754,N_11192,N_11017);
and U11755 (N_11755,N_11048,N_10783);
and U11756 (N_11756,N_10940,N_10842);
nor U11757 (N_11757,N_11157,N_11220);
nand U11758 (N_11758,N_11229,N_10653);
or U11759 (N_11759,N_11234,N_10626);
nand U11760 (N_11760,N_11050,N_10829);
nor U11761 (N_11761,N_10729,N_11189);
and U11762 (N_11762,N_11157,N_10959);
or U11763 (N_11763,N_11190,N_10707);
xnor U11764 (N_11764,N_10821,N_10894);
and U11765 (N_11765,N_11021,N_10664);
and U11766 (N_11766,N_10650,N_10964);
nand U11767 (N_11767,N_10975,N_11172);
and U11768 (N_11768,N_10991,N_11133);
and U11769 (N_11769,N_11004,N_11104);
nor U11770 (N_11770,N_10923,N_10790);
xor U11771 (N_11771,N_11151,N_11132);
nand U11772 (N_11772,N_10877,N_10816);
and U11773 (N_11773,N_10646,N_11243);
nor U11774 (N_11774,N_10827,N_10703);
nor U11775 (N_11775,N_10975,N_10974);
or U11776 (N_11776,N_10817,N_10816);
or U11777 (N_11777,N_10871,N_10874);
nand U11778 (N_11778,N_11191,N_11009);
or U11779 (N_11779,N_10752,N_11239);
xor U11780 (N_11780,N_10798,N_11180);
nor U11781 (N_11781,N_10705,N_10762);
and U11782 (N_11782,N_11135,N_11006);
and U11783 (N_11783,N_10893,N_11237);
or U11784 (N_11784,N_11232,N_10817);
or U11785 (N_11785,N_11047,N_10659);
nand U11786 (N_11786,N_11173,N_11211);
and U11787 (N_11787,N_11021,N_10768);
xor U11788 (N_11788,N_10982,N_11245);
nand U11789 (N_11789,N_11207,N_11114);
nand U11790 (N_11790,N_10809,N_11246);
nor U11791 (N_11791,N_10650,N_11147);
or U11792 (N_11792,N_10651,N_11152);
and U11793 (N_11793,N_10884,N_10815);
nand U11794 (N_11794,N_11228,N_11003);
or U11795 (N_11795,N_10980,N_11203);
nand U11796 (N_11796,N_10815,N_10716);
and U11797 (N_11797,N_10680,N_11208);
nor U11798 (N_11798,N_10975,N_11037);
nor U11799 (N_11799,N_11115,N_11019);
xor U11800 (N_11800,N_11228,N_10859);
nor U11801 (N_11801,N_11198,N_11234);
or U11802 (N_11802,N_10933,N_10763);
or U11803 (N_11803,N_10916,N_10995);
nor U11804 (N_11804,N_11068,N_10985);
and U11805 (N_11805,N_11126,N_10895);
nor U11806 (N_11806,N_10675,N_11014);
nor U11807 (N_11807,N_11021,N_10690);
nor U11808 (N_11808,N_11160,N_10636);
xor U11809 (N_11809,N_11007,N_10814);
nor U11810 (N_11810,N_11194,N_10821);
or U11811 (N_11811,N_10843,N_11100);
nor U11812 (N_11812,N_10846,N_11031);
or U11813 (N_11813,N_11190,N_11100);
nand U11814 (N_11814,N_10898,N_10670);
xor U11815 (N_11815,N_10882,N_11104);
xnor U11816 (N_11816,N_10985,N_10844);
nand U11817 (N_11817,N_10883,N_10811);
nor U11818 (N_11818,N_10642,N_11145);
and U11819 (N_11819,N_10655,N_11155);
xor U11820 (N_11820,N_11045,N_10948);
nand U11821 (N_11821,N_11018,N_10648);
and U11822 (N_11822,N_10836,N_10923);
and U11823 (N_11823,N_10625,N_11192);
nand U11824 (N_11824,N_11114,N_11079);
nand U11825 (N_11825,N_10848,N_11170);
nor U11826 (N_11826,N_11032,N_10741);
or U11827 (N_11827,N_11192,N_10694);
xnor U11828 (N_11828,N_10996,N_11152);
nand U11829 (N_11829,N_11232,N_10677);
xor U11830 (N_11830,N_10882,N_11068);
xor U11831 (N_11831,N_10846,N_10966);
and U11832 (N_11832,N_10914,N_10846);
nand U11833 (N_11833,N_11201,N_11223);
xnor U11834 (N_11834,N_10924,N_11196);
nand U11835 (N_11835,N_11001,N_11038);
or U11836 (N_11836,N_11199,N_10656);
nand U11837 (N_11837,N_11202,N_11148);
and U11838 (N_11838,N_11034,N_11093);
nand U11839 (N_11839,N_11189,N_10931);
nor U11840 (N_11840,N_10946,N_10826);
xnor U11841 (N_11841,N_11056,N_11071);
nand U11842 (N_11842,N_10969,N_11141);
xnor U11843 (N_11843,N_10738,N_11118);
nor U11844 (N_11844,N_10702,N_10913);
or U11845 (N_11845,N_10983,N_10733);
and U11846 (N_11846,N_11152,N_11203);
or U11847 (N_11847,N_11003,N_11154);
nor U11848 (N_11848,N_10782,N_10976);
or U11849 (N_11849,N_10700,N_11213);
or U11850 (N_11850,N_10824,N_10967);
nand U11851 (N_11851,N_10786,N_11137);
nor U11852 (N_11852,N_10855,N_10935);
and U11853 (N_11853,N_11192,N_11129);
or U11854 (N_11854,N_11017,N_11085);
and U11855 (N_11855,N_10941,N_11127);
nor U11856 (N_11856,N_10947,N_11241);
and U11857 (N_11857,N_10937,N_11122);
nand U11858 (N_11858,N_10873,N_10867);
nor U11859 (N_11859,N_11029,N_11169);
or U11860 (N_11860,N_10792,N_11235);
or U11861 (N_11861,N_10685,N_10662);
or U11862 (N_11862,N_10760,N_10767);
nand U11863 (N_11863,N_10778,N_10760);
and U11864 (N_11864,N_10939,N_10644);
and U11865 (N_11865,N_10814,N_10983);
nand U11866 (N_11866,N_11036,N_11237);
or U11867 (N_11867,N_11139,N_11018);
nand U11868 (N_11868,N_11062,N_11079);
nor U11869 (N_11869,N_10630,N_10672);
or U11870 (N_11870,N_11066,N_10999);
and U11871 (N_11871,N_10848,N_10919);
nand U11872 (N_11872,N_11140,N_11055);
nand U11873 (N_11873,N_10820,N_10661);
or U11874 (N_11874,N_11210,N_11061);
and U11875 (N_11875,N_11851,N_11375);
nor U11876 (N_11876,N_11287,N_11489);
and U11877 (N_11877,N_11609,N_11474);
or U11878 (N_11878,N_11591,N_11271);
or U11879 (N_11879,N_11267,N_11488);
and U11880 (N_11880,N_11771,N_11722);
xnor U11881 (N_11881,N_11266,N_11505);
nand U11882 (N_11882,N_11671,N_11509);
and U11883 (N_11883,N_11466,N_11377);
xnor U11884 (N_11884,N_11842,N_11286);
nand U11885 (N_11885,N_11443,N_11477);
xnor U11886 (N_11886,N_11476,N_11741);
and U11887 (N_11887,N_11858,N_11732);
and U11888 (N_11888,N_11371,N_11284);
or U11889 (N_11889,N_11696,N_11648);
and U11890 (N_11890,N_11690,N_11360);
nor U11891 (N_11891,N_11574,N_11770);
or U11892 (N_11892,N_11810,N_11265);
nand U11893 (N_11893,N_11593,N_11407);
nand U11894 (N_11894,N_11320,N_11816);
nand U11895 (N_11895,N_11758,N_11781);
and U11896 (N_11896,N_11366,N_11429);
or U11897 (N_11897,N_11381,N_11277);
and U11898 (N_11898,N_11307,N_11874);
xnor U11899 (N_11899,N_11420,N_11693);
nor U11900 (N_11900,N_11340,N_11829);
nor U11901 (N_11901,N_11677,N_11409);
or U11902 (N_11902,N_11512,N_11386);
nand U11903 (N_11903,N_11322,N_11864);
nand U11904 (N_11904,N_11520,N_11497);
or U11905 (N_11905,N_11753,N_11662);
nand U11906 (N_11906,N_11706,N_11581);
nor U11907 (N_11907,N_11463,N_11451);
nand U11908 (N_11908,N_11805,N_11659);
xor U11909 (N_11909,N_11744,N_11608);
nand U11910 (N_11910,N_11362,N_11657);
and U11911 (N_11911,N_11844,N_11332);
nand U11912 (N_11912,N_11660,N_11329);
nor U11913 (N_11913,N_11542,N_11632);
and U11914 (N_11914,N_11395,N_11708);
nand U11915 (N_11915,N_11786,N_11513);
and U11916 (N_11916,N_11623,N_11754);
nand U11917 (N_11917,N_11470,N_11298);
xnor U11918 (N_11918,N_11646,N_11358);
nor U11919 (N_11919,N_11638,N_11764);
nand U11920 (N_11920,N_11427,N_11567);
nor U11921 (N_11921,N_11725,N_11557);
and U11922 (N_11922,N_11485,N_11288);
nor U11923 (N_11923,N_11578,N_11422);
nand U11924 (N_11924,N_11746,N_11825);
or U11925 (N_11925,N_11668,N_11596);
or U11926 (N_11926,N_11674,N_11773);
nand U11927 (N_11927,N_11647,N_11406);
nand U11928 (N_11928,N_11599,N_11262);
and U11929 (N_11929,N_11572,N_11683);
and U11930 (N_11930,N_11432,N_11280);
and U11931 (N_11931,N_11584,N_11803);
xor U11932 (N_11932,N_11317,N_11516);
or U11933 (N_11933,N_11496,N_11855);
and U11934 (N_11934,N_11819,N_11873);
nand U11935 (N_11935,N_11761,N_11694);
nand U11936 (N_11936,N_11795,N_11532);
nand U11937 (N_11937,N_11510,N_11425);
nor U11938 (N_11938,N_11491,N_11800);
nor U11939 (N_11939,N_11270,N_11653);
nor U11940 (N_11940,N_11272,N_11282);
or U11941 (N_11941,N_11484,N_11459);
and U11942 (N_11942,N_11724,N_11335);
nor U11943 (N_11943,N_11498,N_11762);
nand U11944 (N_11944,N_11734,N_11403);
nor U11945 (N_11945,N_11467,N_11791);
nand U11946 (N_11946,N_11643,N_11811);
or U11947 (N_11947,N_11849,N_11723);
or U11948 (N_11948,N_11837,N_11388);
nor U11949 (N_11949,N_11796,N_11302);
xnor U11950 (N_11950,N_11251,N_11555);
xor U11951 (N_11951,N_11530,N_11794);
and U11952 (N_11952,N_11279,N_11590);
nor U11953 (N_11953,N_11308,N_11504);
and U11954 (N_11954,N_11768,N_11718);
and U11955 (N_11955,N_11319,N_11334);
and U11956 (N_11956,N_11374,N_11503);
xor U11957 (N_11957,N_11323,N_11644);
xor U11958 (N_11958,N_11424,N_11614);
and U11959 (N_11959,N_11861,N_11268);
or U11960 (N_11960,N_11621,N_11398);
xor U11961 (N_11961,N_11444,N_11742);
nor U11962 (N_11962,N_11801,N_11835);
and U11963 (N_11963,N_11804,N_11856);
nor U11964 (N_11964,N_11448,N_11564);
or U11965 (N_11965,N_11872,N_11667);
nor U11966 (N_11966,N_11352,N_11684);
nor U11967 (N_11967,N_11600,N_11393);
nand U11968 (N_11968,N_11691,N_11511);
nand U11969 (N_11969,N_11613,N_11766);
nor U11970 (N_11970,N_11397,N_11812);
xnor U11971 (N_11971,N_11309,N_11547);
or U11972 (N_11972,N_11365,N_11688);
nand U11973 (N_11973,N_11654,N_11678);
nor U11974 (N_11974,N_11501,N_11556);
and U11975 (N_11975,N_11651,N_11533);
and U11976 (N_11976,N_11412,N_11281);
and U11977 (N_11977,N_11713,N_11839);
nor U11978 (N_11978,N_11767,N_11487);
xnor U11979 (N_11979,N_11740,N_11345);
nand U11980 (N_11980,N_11418,N_11853);
and U11981 (N_11981,N_11588,N_11356);
and U11982 (N_11982,N_11363,N_11624);
nand U11983 (N_11983,N_11612,N_11344);
or U11984 (N_11984,N_11346,N_11670);
xnor U11985 (N_11985,N_11528,N_11703);
nand U11986 (N_11986,N_11715,N_11756);
or U11987 (N_11987,N_11454,N_11868);
nand U11988 (N_11988,N_11757,N_11685);
nand U11989 (N_11989,N_11622,N_11414);
or U11990 (N_11990,N_11431,N_11628);
and U11991 (N_11991,N_11481,N_11539);
nand U11992 (N_11992,N_11502,N_11368);
nor U11993 (N_11993,N_11438,N_11442);
and U11994 (N_11994,N_11604,N_11351);
nand U11995 (N_11995,N_11680,N_11494);
nand U11996 (N_11996,N_11765,N_11404);
and U11997 (N_11997,N_11847,N_11790);
nor U11998 (N_11998,N_11821,N_11536);
xor U11999 (N_11999,N_11348,N_11626);
or U12000 (N_12000,N_11370,N_11682);
and U12001 (N_12001,N_11373,N_11832);
or U12002 (N_12002,N_11413,N_11769);
xnor U12003 (N_12003,N_11276,N_11618);
or U12004 (N_12004,N_11752,N_11263);
nor U12005 (N_12005,N_11552,N_11645);
and U12006 (N_12006,N_11392,N_11433);
nand U12007 (N_12007,N_11633,N_11695);
or U12008 (N_12008,N_11866,N_11824);
nor U12009 (N_12009,N_11782,N_11382);
and U12010 (N_12010,N_11702,N_11293);
xnor U12011 (N_12011,N_11699,N_11558);
xor U12012 (N_12012,N_11750,N_11522);
nand U12013 (N_12013,N_11828,N_11390);
and U12014 (N_12014,N_11355,N_11321);
nor U12015 (N_12015,N_11598,N_11294);
or U12016 (N_12016,N_11384,N_11871);
nor U12017 (N_12017,N_11610,N_11870);
and U12018 (N_12018,N_11391,N_11629);
and U12019 (N_12019,N_11326,N_11303);
or U12020 (N_12020,N_11549,N_11434);
and U12021 (N_12021,N_11834,N_11807);
nand U12022 (N_12022,N_11748,N_11527);
nand U12023 (N_12023,N_11721,N_11486);
nand U12024 (N_12024,N_11772,N_11299);
nor U12025 (N_12025,N_11405,N_11252);
and U12026 (N_12026,N_11324,N_11450);
nand U12027 (N_12027,N_11843,N_11692);
and U12028 (N_12028,N_11712,N_11378);
nor U12029 (N_12029,N_11551,N_11447);
or U12030 (N_12030,N_11714,N_11305);
nor U12031 (N_12031,N_11274,N_11430);
or U12032 (N_12032,N_11658,N_11594);
and U12033 (N_12033,N_11777,N_11827);
xor U12034 (N_12034,N_11636,N_11455);
nor U12035 (N_12035,N_11561,N_11639);
and U12036 (N_12036,N_11697,N_11473);
and U12037 (N_12037,N_11865,N_11353);
xor U12038 (N_12038,N_11469,N_11701);
or U12039 (N_12039,N_11291,N_11440);
nand U12040 (N_12040,N_11642,N_11793);
nor U12041 (N_12041,N_11717,N_11707);
nor U12042 (N_12042,N_11566,N_11415);
or U12043 (N_12043,N_11784,N_11426);
nand U12044 (N_12044,N_11495,N_11820);
or U12045 (N_12045,N_11656,N_11799);
nand U12046 (N_12046,N_11774,N_11526);
or U12047 (N_12047,N_11649,N_11400);
or U12048 (N_12048,N_11738,N_11797);
and U12049 (N_12049,N_11508,N_11806);
or U12050 (N_12050,N_11710,N_11479);
nor U12051 (N_12051,N_11840,N_11327);
and U12052 (N_12052,N_11285,N_11576);
xnor U12053 (N_12053,N_11676,N_11802);
or U12054 (N_12054,N_11269,N_11411);
nand U12055 (N_12055,N_11437,N_11537);
nor U12056 (N_12056,N_11318,N_11541);
nor U12057 (N_12057,N_11260,N_11417);
nor U12058 (N_12058,N_11261,N_11739);
nor U12059 (N_12059,N_11822,N_11419);
or U12060 (N_12060,N_11401,N_11544);
and U12061 (N_12061,N_11607,N_11337);
and U12062 (N_12062,N_11585,N_11376);
or U12063 (N_12063,N_11867,N_11300);
nand U12064 (N_12064,N_11283,N_11312);
nor U12065 (N_12065,N_11850,N_11663);
nor U12066 (N_12066,N_11689,N_11705);
and U12067 (N_12067,N_11780,N_11304);
nand U12068 (N_12068,N_11273,N_11749);
nor U12069 (N_12069,N_11665,N_11361);
and U12070 (N_12070,N_11809,N_11783);
nand U12071 (N_12071,N_11728,N_11854);
nor U12072 (N_12072,N_11775,N_11357);
nor U12073 (N_12073,N_11367,N_11347);
nor U12074 (N_12074,N_11529,N_11760);
xor U12075 (N_12075,N_11331,N_11635);
and U12076 (N_12076,N_11278,N_11560);
nor U12077 (N_12077,N_11387,N_11258);
nor U12078 (N_12078,N_11457,N_11500);
nor U12079 (N_12079,N_11545,N_11606);
nand U12080 (N_12080,N_11571,N_11255);
or U12081 (N_12081,N_11468,N_11506);
nor U12082 (N_12082,N_11313,N_11860);
and U12083 (N_12083,N_11583,N_11364);
and U12084 (N_12084,N_11634,N_11751);
nand U12085 (N_12085,N_11446,N_11369);
or U12086 (N_12086,N_11640,N_11380);
nand U12087 (N_12087,N_11836,N_11435);
and U12088 (N_12088,N_11314,N_11253);
and U12089 (N_12089,N_11589,N_11823);
and U12090 (N_12090,N_11514,N_11681);
xor U12091 (N_12091,N_11465,N_11471);
nand U12092 (N_12092,N_11808,N_11499);
and U12093 (N_12093,N_11845,N_11521);
nor U12094 (N_12094,N_11436,N_11568);
nand U12095 (N_12095,N_11815,N_11306);
xnor U12096 (N_12096,N_11254,N_11587);
and U12097 (N_12097,N_11830,N_11661);
or U12098 (N_12098,N_11534,N_11492);
xnor U12099 (N_12099,N_11630,N_11517);
and U12100 (N_12100,N_11582,N_11833);
or U12101 (N_12101,N_11727,N_11814);
or U12102 (N_12102,N_11538,N_11655);
or U12103 (N_12103,N_11563,N_11577);
and U12104 (N_12104,N_11535,N_11562);
nor U12105 (N_12105,N_11666,N_11720);
and U12106 (N_12106,N_11453,N_11264);
and U12107 (N_12107,N_11846,N_11817);
and U12108 (N_12108,N_11421,N_11402);
xnor U12109 (N_12109,N_11379,N_11863);
nor U12110 (N_12110,N_11259,N_11523);
or U12111 (N_12111,N_11704,N_11579);
nand U12112 (N_12112,N_11428,N_11316);
nor U12113 (N_12113,N_11755,N_11831);
xnor U12114 (N_12114,N_11519,N_11342);
nor U12115 (N_12115,N_11543,N_11698);
or U12116 (N_12116,N_11275,N_11869);
nor U12117 (N_12117,N_11441,N_11333);
nand U12118 (N_12118,N_11611,N_11826);
or U12119 (N_12119,N_11852,N_11383);
or U12120 (N_12120,N_11838,N_11625);
or U12121 (N_12121,N_11290,N_11615);
xor U12122 (N_12122,N_11711,N_11408);
or U12123 (N_12123,N_11452,N_11857);
xnor U12124 (N_12124,N_11641,N_11546);
or U12125 (N_12125,N_11396,N_11592);
nor U12126 (N_12126,N_11788,N_11730);
xnor U12127 (N_12127,N_11296,N_11595);
nand U12128 (N_12128,N_11672,N_11743);
nand U12129 (N_12129,N_11605,N_11480);
or U12130 (N_12130,N_11862,N_11439);
and U12131 (N_12131,N_11664,N_11416);
nor U12132 (N_12132,N_11779,N_11601);
and U12133 (N_12133,N_11462,N_11673);
and U12134 (N_12134,N_11620,N_11548);
nor U12135 (N_12135,N_11464,N_11341);
and U12136 (N_12136,N_11531,N_11745);
or U12137 (N_12137,N_11616,N_11603);
or U12138 (N_12138,N_11569,N_11445);
or U12139 (N_12139,N_11540,N_11733);
nand U12140 (N_12140,N_11716,N_11559);
or U12141 (N_12141,N_11686,N_11841);
and U12142 (N_12142,N_11385,N_11349);
and U12143 (N_12143,N_11478,N_11483);
and U12144 (N_12144,N_11336,N_11257);
xnor U12145 (N_12145,N_11410,N_11289);
nor U12146 (N_12146,N_11325,N_11787);
nor U12147 (N_12147,N_11778,N_11525);
nand U12148 (N_12148,N_11679,N_11565);
nor U12149 (N_12149,N_11737,N_11652);
nand U12150 (N_12150,N_11399,N_11729);
nand U12151 (N_12151,N_11493,N_11354);
nor U12152 (N_12152,N_11458,N_11315);
nor U12153 (N_12153,N_11575,N_11461);
xnor U12154 (N_12154,N_11389,N_11338);
or U12155 (N_12155,N_11292,N_11339);
and U12156 (N_12156,N_11586,N_11343);
and U12157 (N_12157,N_11394,N_11818);
nor U12158 (N_12158,N_11813,N_11515);
and U12159 (N_12159,N_11310,N_11763);
nor U12160 (N_12160,N_11627,N_11669);
nor U12161 (N_12161,N_11848,N_11460);
nor U12162 (N_12162,N_11518,N_11709);
or U12163 (N_12163,N_11554,N_11580);
nor U12164 (N_12164,N_11726,N_11785);
nor U12165 (N_12165,N_11619,N_11687);
nand U12166 (N_12166,N_11482,N_11731);
nor U12167 (N_12167,N_11789,N_11256);
nor U12168 (N_12168,N_11637,N_11759);
nor U12169 (N_12169,N_11297,N_11301);
and U12170 (N_12170,N_11859,N_11350);
nand U12171 (N_12171,N_11736,N_11330);
nor U12172 (N_12172,N_11311,N_11423);
nand U12173 (N_12173,N_11372,N_11449);
nand U12174 (N_12174,N_11295,N_11456);
and U12175 (N_12175,N_11719,N_11553);
and U12176 (N_12176,N_11631,N_11602);
or U12177 (N_12177,N_11747,N_11792);
and U12178 (N_12178,N_11617,N_11359);
nor U12179 (N_12179,N_11675,N_11597);
or U12180 (N_12180,N_11475,N_11570);
xor U12181 (N_12181,N_11573,N_11250);
and U12182 (N_12182,N_11798,N_11550);
nor U12183 (N_12183,N_11700,N_11735);
or U12184 (N_12184,N_11507,N_11776);
nand U12185 (N_12185,N_11472,N_11524);
and U12186 (N_12186,N_11650,N_11490);
xor U12187 (N_12187,N_11328,N_11830);
nand U12188 (N_12188,N_11820,N_11795);
nor U12189 (N_12189,N_11334,N_11496);
nor U12190 (N_12190,N_11353,N_11789);
nor U12191 (N_12191,N_11494,N_11767);
nand U12192 (N_12192,N_11812,N_11850);
or U12193 (N_12193,N_11757,N_11714);
and U12194 (N_12194,N_11660,N_11483);
nand U12195 (N_12195,N_11715,N_11377);
xnor U12196 (N_12196,N_11781,N_11302);
and U12197 (N_12197,N_11751,N_11345);
nor U12198 (N_12198,N_11649,N_11658);
or U12199 (N_12199,N_11734,N_11473);
or U12200 (N_12200,N_11711,N_11614);
and U12201 (N_12201,N_11832,N_11663);
xor U12202 (N_12202,N_11465,N_11435);
and U12203 (N_12203,N_11501,N_11271);
or U12204 (N_12204,N_11629,N_11811);
xor U12205 (N_12205,N_11344,N_11734);
or U12206 (N_12206,N_11830,N_11583);
or U12207 (N_12207,N_11502,N_11632);
or U12208 (N_12208,N_11449,N_11691);
or U12209 (N_12209,N_11271,N_11338);
nand U12210 (N_12210,N_11255,N_11368);
nand U12211 (N_12211,N_11453,N_11405);
and U12212 (N_12212,N_11393,N_11789);
xnor U12213 (N_12213,N_11506,N_11446);
nand U12214 (N_12214,N_11824,N_11622);
nand U12215 (N_12215,N_11812,N_11590);
and U12216 (N_12216,N_11561,N_11515);
or U12217 (N_12217,N_11562,N_11799);
xor U12218 (N_12218,N_11856,N_11264);
xnor U12219 (N_12219,N_11258,N_11271);
nand U12220 (N_12220,N_11392,N_11645);
nor U12221 (N_12221,N_11736,N_11597);
or U12222 (N_12222,N_11280,N_11299);
nand U12223 (N_12223,N_11350,N_11795);
and U12224 (N_12224,N_11710,N_11260);
nand U12225 (N_12225,N_11340,N_11498);
or U12226 (N_12226,N_11835,N_11341);
and U12227 (N_12227,N_11526,N_11563);
nand U12228 (N_12228,N_11513,N_11685);
and U12229 (N_12229,N_11351,N_11358);
nor U12230 (N_12230,N_11588,N_11726);
nand U12231 (N_12231,N_11274,N_11489);
xnor U12232 (N_12232,N_11716,N_11597);
xnor U12233 (N_12233,N_11290,N_11462);
or U12234 (N_12234,N_11539,N_11823);
nand U12235 (N_12235,N_11840,N_11743);
and U12236 (N_12236,N_11391,N_11308);
nand U12237 (N_12237,N_11302,N_11715);
nor U12238 (N_12238,N_11727,N_11355);
xnor U12239 (N_12239,N_11435,N_11401);
nand U12240 (N_12240,N_11676,N_11738);
nand U12241 (N_12241,N_11686,N_11821);
or U12242 (N_12242,N_11550,N_11790);
xnor U12243 (N_12243,N_11380,N_11613);
and U12244 (N_12244,N_11485,N_11750);
or U12245 (N_12245,N_11392,N_11432);
nor U12246 (N_12246,N_11320,N_11506);
and U12247 (N_12247,N_11301,N_11313);
nor U12248 (N_12248,N_11291,N_11870);
or U12249 (N_12249,N_11832,N_11324);
nand U12250 (N_12250,N_11275,N_11485);
nor U12251 (N_12251,N_11495,N_11677);
and U12252 (N_12252,N_11455,N_11545);
nand U12253 (N_12253,N_11690,N_11664);
nand U12254 (N_12254,N_11635,N_11753);
nand U12255 (N_12255,N_11742,N_11379);
nor U12256 (N_12256,N_11784,N_11477);
or U12257 (N_12257,N_11441,N_11309);
nor U12258 (N_12258,N_11508,N_11285);
and U12259 (N_12259,N_11281,N_11478);
nor U12260 (N_12260,N_11866,N_11258);
nand U12261 (N_12261,N_11467,N_11437);
and U12262 (N_12262,N_11635,N_11547);
nor U12263 (N_12263,N_11799,N_11261);
nand U12264 (N_12264,N_11803,N_11871);
nand U12265 (N_12265,N_11664,N_11397);
or U12266 (N_12266,N_11808,N_11550);
nand U12267 (N_12267,N_11737,N_11755);
nor U12268 (N_12268,N_11639,N_11345);
or U12269 (N_12269,N_11674,N_11702);
and U12270 (N_12270,N_11261,N_11854);
and U12271 (N_12271,N_11610,N_11622);
and U12272 (N_12272,N_11637,N_11803);
nor U12273 (N_12273,N_11367,N_11520);
xnor U12274 (N_12274,N_11343,N_11848);
and U12275 (N_12275,N_11510,N_11542);
or U12276 (N_12276,N_11780,N_11510);
or U12277 (N_12277,N_11677,N_11645);
and U12278 (N_12278,N_11816,N_11786);
and U12279 (N_12279,N_11713,N_11266);
nand U12280 (N_12280,N_11388,N_11464);
nand U12281 (N_12281,N_11385,N_11443);
nand U12282 (N_12282,N_11606,N_11442);
or U12283 (N_12283,N_11440,N_11773);
nor U12284 (N_12284,N_11670,N_11642);
nand U12285 (N_12285,N_11731,N_11376);
xor U12286 (N_12286,N_11793,N_11395);
or U12287 (N_12287,N_11310,N_11250);
nand U12288 (N_12288,N_11498,N_11356);
and U12289 (N_12289,N_11594,N_11730);
nor U12290 (N_12290,N_11592,N_11530);
nand U12291 (N_12291,N_11624,N_11749);
and U12292 (N_12292,N_11276,N_11333);
xnor U12293 (N_12293,N_11279,N_11677);
nor U12294 (N_12294,N_11454,N_11775);
nor U12295 (N_12295,N_11324,N_11724);
or U12296 (N_12296,N_11477,N_11271);
and U12297 (N_12297,N_11714,N_11273);
and U12298 (N_12298,N_11357,N_11536);
or U12299 (N_12299,N_11616,N_11332);
and U12300 (N_12300,N_11622,N_11547);
nand U12301 (N_12301,N_11579,N_11745);
and U12302 (N_12302,N_11404,N_11468);
nor U12303 (N_12303,N_11695,N_11416);
nand U12304 (N_12304,N_11674,N_11836);
nor U12305 (N_12305,N_11548,N_11788);
nand U12306 (N_12306,N_11569,N_11460);
xnor U12307 (N_12307,N_11629,N_11356);
or U12308 (N_12308,N_11522,N_11340);
or U12309 (N_12309,N_11828,N_11486);
nor U12310 (N_12310,N_11479,N_11771);
or U12311 (N_12311,N_11565,N_11646);
and U12312 (N_12312,N_11862,N_11615);
nand U12313 (N_12313,N_11674,N_11514);
nor U12314 (N_12314,N_11514,N_11759);
or U12315 (N_12315,N_11559,N_11653);
nand U12316 (N_12316,N_11463,N_11257);
nor U12317 (N_12317,N_11393,N_11386);
and U12318 (N_12318,N_11353,N_11541);
nor U12319 (N_12319,N_11367,N_11831);
nor U12320 (N_12320,N_11841,N_11728);
and U12321 (N_12321,N_11813,N_11406);
and U12322 (N_12322,N_11256,N_11491);
nand U12323 (N_12323,N_11725,N_11727);
nand U12324 (N_12324,N_11303,N_11808);
nor U12325 (N_12325,N_11273,N_11857);
or U12326 (N_12326,N_11738,N_11638);
nand U12327 (N_12327,N_11500,N_11849);
nor U12328 (N_12328,N_11735,N_11697);
or U12329 (N_12329,N_11797,N_11464);
or U12330 (N_12330,N_11847,N_11446);
nor U12331 (N_12331,N_11815,N_11327);
and U12332 (N_12332,N_11519,N_11641);
or U12333 (N_12333,N_11527,N_11530);
or U12334 (N_12334,N_11369,N_11729);
nand U12335 (N_12335,N_11504,N_11284);
xor U12336 (N_12336,N_11815,N_11840);
or U12337 (N_12337,N_11255,N_11281);
and U12338 (N_12338,N_11587,N_11499);
or U12339 (N_12339,N_11856,N_11373);
and U12340 (N_12340,N_11687,N_11507);
xnor U12341 (N_12341,N_11534,N_11814);
or U12342 (N_12342,N_11420,N_11767);
nor U12343 (N_12343,N_11444,N_11864);
nor U12344 (N_12344,N_11555,N_11315);
or U12345 (N_12345,N_11323,N_11482);
nor U12346 (N_12346,N_11266,N_11340);
nor U12347 (N_12347,N_11767,N_11465);
xnor U12348 (N_12348,N_11648,N_11263);
nor U12349 (N_12349,N_11798,N_11659);
nand U12350 (N_12350,N_11352,N_11268);
or U12351 (N_12351,N_11729,N_11289);
nor U12352 (N_12352,N_11721,N_11286);
nor U12353 (N_12353,N_11258,N_11707);
or U12354 (N_12354,N_11756,N_11817);
nor U12355 (N_12355,N_11310,N_11808);
and U12356 (N_12356,N_11524,N_11598);
or U12357 (N_12357,N_11743,N_11371);
nor U12358 (N_12358,N_11648,N_11301);
and U12359 (N_12359,N_11384,N_11290);
nand U12360 (N_12360,N_11679,N_11510);
nand U12361 (N_12361,N_11715,N_11730);
nor U12362 (N_12362,N_11498,N_11354);
or U12363 (N_12363,N_11834,N_11541);
nand U12364 (N_12364,N_11859,N_11807);
xor U12365 (N_12365,N_11475,N_11683);
xnor U12366 (N_12366,N_11316,N_11740);
nor U12367 (N_12367,N_11812,N_11620);
nand U12368 (N_12368,N_11379,N_11628);
nor U12369 (N_12369,N_11571,N_11622);
and U12370 (N_12370,N_11708,N_11537);
and U12371 (N_12371,N_11797,N_11583);
nand U12372 (N_12372,N_11468,N_11612);
nand U12373 (N_12373,N_11651,N_11633);
nand U12374 (N_12374,N_11840,N_11780);
nand U12375 (N_12375,N_11456,N_11736);
and U12376 (N_12376,N_11612,N_11345);
or U12377 (N_12377,N_11662,N_11490);
nand U12378 (N_12378,N_11856,N_11512);
and U12379 (N_12379,N_11598,N_11350);
nor U12380 (N_12380,N_11825,N_11335);
nand U12381 (N_12381,N_11762,N_11626);
nand U12382 (N_12382,N_11502,N_11433);
or U12383 (N_12383,N_11739,N_11318);
or U12384 (N_12384,N_11707,N_11552);
and U12385 (N_12385,N_11284,N_11589);
or U12386 (N_12386,N_11761,N_11302);
nor U12387 (N_12387,N_11399,N_11489);
or U12388 (N_12388,N_11264,N_11381);
nand U12389 (N_12389,N_11688,N_11687);
nand U12390 (N_12390,N_11250,N_11818);
or U12391 (N_12391,N_11477,N_11733);
or U12392 (N_12392,N_11474,N_11360);
xor U12393 (N_12393,N_11822,N_11728);
and U12394 (N_12394,N_11625,N_11291);
xnor U12395 (N_12395,N_11843,N_11343);
xor U12396 (N_12396,N_11357,N_11320);
nand U12397 (N_12397,N_11707,N_11354);
or U12398 (N_12398,N_11491,N_11558);
nand U12399 (N_12399,N_11355,N_11700);
or U12400 (N_12400,N_11689,N_11809);
and U12401 (N_12401,N_11687,N_11586);
or U12402 (N_12402,N_11651,N_11632);
xor U12403 (N_12403,N_11481,N_11662);
or U12404 (N_12404,N_11676,N_11719);
nand U12405 (N_12405,N_11574,N_11702);
or U12406 (N_12406,N_11751,N_11355);
or U12407 (N_12407,N_11699,N_11868);
or U12408 (N_12408,N_11855,N_11312);
nand U12409 (N_12409,N_11431,N_11596);
xnor U12410 (N_12410,N_11329,N_11661);
and U12411 (N_12411,N_11689,N_11413);
or U12412 (N_12412,N_11433,N_11683);
xor U12413 (N_12413,N_11285,N_11873);
and U12414 (N_12414,N_11680,N_11331);
and U12415 (N_12415,N_11681,N_11592);
nand U12416 (N_12416,N_11784,N_11814);
nand U12417 (N_12417,N_11562,N_11707);
and U12418 (N_12418,N_11496,N_11460);
nand U12419 (N_12419,N_11482,N_11254);
nor U12420 (N_12420,N_11370,N_11720);
nand U12421 (N_12421,N_11514,N_11600);
or U12422 (N_12422,N_11377,N_11300);
and U12423 (N_12423,N_11658,N_11788);
xor U12424 (N_12424,N_11702,N_11790);
or U12425 (N_12425,N_11660,N_11699);
nor U12426 (N_12426,N_11342,N_11707);
nand U12427 (N_12427,N_11719,N_11635);
nor U12428 (N_12428,N_11776,N_11856);
and U12429 (N_12429,N_11814,N_11440);
or U12430 (N_12430,N_11281,N_11257);
and U12431 (N_12431,N_11529,N_11767);
or U12432 (N_12432,N_11597,N_11729);
or U12433 (N_12433,N_11524,N_11663);
nand U12434 (N_12434,N_11453,N_11280);
or U12435 (N_12435,N_11728,N_11348);
nor U12436 (N_12436,N_11869,N_11343);
and U12437 (N_12437,N_11770,N_11728);
and U12438 (N_12438,N_11548,N_11799);
or U12439 (N_12439,N_11829,N_11305);
and U12440 (N_12440,N_11715,N_11467);
and U12441 (N_12441,N_11649,N_11496);
nor U12442 (N_12442,N_11291,N_11278);
nor U12443 (N_12443,N_11451,N_11383);
and U12444 (N_12444,N_11722,N_11550);
and U12445 (N_12445,N_11753,N_11540);
nor U12446 (N_12446,N_11854,N_11301);
xor U12447 (N_12447,N_11782,N_11305);
nor U12448 (N_12448,N_11350,N_11353);
and U12449 (N_12449,N_11722,N_11660);
nand U12450 (N_12450,N_11420,N_11298);
and U12451 (N_12451,N_11633,N_11510);
nor U12452 (N_12452,N_11382,N_11593);
nand U12453 (N_12453,N_11523,N_11409);
nand U12454 (N_12454,N_11449,N_11333);
nor U12455 (N_12455,N_11307,N_11835);
and U12456 (N_12456,N_11694,N_11849);
and U12457 (N_12457,N_11667,N_11602);
nor U12458 (N_12458,N_11332,N_11251);
nor U12459 (N_12459,N_11557,N_11606);
nand U12460 (N_12460,N_11407,N_11820);
nor U12461 (N_12461,N_11381,N_11640);
and U12462 (N_12462,N_11730,N_11377);
nand U12463 (N_12463,N_11458,N_11601);
or U12464 (N_12464,N_11734,N_11828);
and U12465 (N_12465,N_11804,N_11819);
or U12466 (N_12466,N_11847,N_11259);
nand U12467 (N_12467,N_11857,N_11340);
or U12468 (N_12468,N_11769,N_11765);
xnor U12469 (N_12469,N_11590,N_11336);
and U12470 (N_12470,N_11266,N_11267);
or U12471 (N_12471,N_11815,N_11672);
and U12472 (N_12472,N_11732,N_11871);
or U12473 (N_12473,N_11578,N_11523);
nor U12474 (N_12474,N_11785,N_11491);
nor U12475 (N_12475,N_11334,N_11874);
and U12476 (N_12476,N_11334,N_11822);
nand U12477 (N_12477,N_11548,N_11680);
nor U12478 (N_12478,N_11374,N_11280);
nand U12479 (N_12479,N_11600,N_11344);
nand U12480 (N_12480,N_11607,N_11857);
nand U12481 (N_12481,N_11538,N_11758);
nand U12482 (N_12482,N_11853,N_11280);
nand U12483 (N_12483,N_11661,N_11255);
and U12484 (N_12484,N_11645,N_11289);
and U12485 (N_12485,N_11297,N_11485);
nor U12486 (N_12486,N_11819,N_11587);
or U12487 (N_12487,N_11516,N_11832);
or U12488 (N_12488,N_11783,N_11361);
xor U12489 (N_12489,N_11854,N_11367);
or U12490 (N_12490,N_11298,N_11474);
or U12491 (N_12491,N_11485,N_11782);
nor U12492 (N_12492,N_11528,N_11474);
and U12493 (N_12493,N_11661,N_11376);
nand U12494 (N_12494,N_11637,N_11406);
nand U12495 (N_12495,N_11765,N_11717);
and U12496 (N_12496,N_11296,N_11337);
nand U12497 (N_12497,N_11818,N_11607);
nor U12498 (N_12498,N_11585,N_11419);
or U12499 (N_12499,N_11745,N_11503);
nand U12500 (N_12500,N_12440,N_12225);
nand U12501 (N_12501,N_12330,N_12165);
or U12502 (N_12502,N_11977,N_12294);
nand U12503 (N_12503,N_11989,N_12305);
nor U12504 (N_12504,N_12361,N_12350);
xnor U12505 (N_12505,N_12406,N_12214);
and U12506 (N_12506,N_11879,N_12342);
and U12507 (N_12507,N_12327,N_12306);
nand U12508 (N_12508,N_12090,N_12289);
and U12509 (N_12509,N_12016,N_11928);
xnor U12510 (N_12510,N_12161,N_12270);
nand U12511 (N_12511,N_12021,N_12379);
xor U12512 (N_12512,N_12220,N_12099);
xor U12513 (N_12513,N_12065,N_11986);
nand U12514 (N_12514,N_11950,N_11880);
nand U12515 (N_12515,N_12474,N_11885);
and U12516 (N_12516,N_12337,N_12320);
nor U12517 (N_12517,N_12239,N_12167);
nor U12518 (N_12518,N_12496,N_12045);
xnor U12519 (N_12519,N_12345,N_11980);
and U12520 (N_12520,N_12101,N_12378);
nor U12521 (N_12521,N_12138,N_12024);
nor U12522 (N_12522,N_12190,N_12250);
nand U12523 (N_12523,N_12124,N_12051);
nor U12524 (N_12524,N_12210,N_12006);
xor U12525 (N_12525,N_12187,N_12418);
or U12526 (N_12526,N_12475,N_12300);
nand U12527 (N_12527,N_11907,N_12113);
nor U12528 (N_12528,N_12422,N_12233);
and U12529 (N_12529,N_12019,N_12228);
xnor U12530 (N_12530,N_12389,N_12380);
and U12531 (N_12531,N_12287,N_12344);
or U12532 (N_12532,N_12176,N_12472);
or U12533 (N_12533,N_12175,N_11942);
nor U12534 (N_12534,N_12148,N_12497);
nor U12535 (N_12535,N_12286,N_12430);
nor U12536 (N_12536,N_12458,N_12209);
nor U12537 (N_12537,N_12074,N_12040);
and U12538 (N_12538,N_12159,N_12353);
and U12539 (N_12539,N_12028,N_12256);
nor U12540 (N_12540,N_12078,N_12011);
and U12541 (N_12541,N_12243,N_12485);
nor U12542 (N_12542,N_12034,N_12089);
xor U12543 (N_12543,N_12298,N_11965);
nand U12544 (N_12544,N_12399,N_12408);
or U12545 (N_12545,N_12193,N_11915);
or U12546 (N_12546,N_12046,N_11946);
xor U12547 (N_12547,N_12030,N_11964);
or U12548 (N_12548,N_12396,N_12236);
nor U12549 (N_12549,N_12272,N_12010);
nor U12550 (N_12550,N_12255,N_12318);
or U12551 (N_12551,N_12237,N_11932);
xor U12552 (N_12552,N_11967,N_12087);
xor U12553 (N_12553,N_12299,N_12035);
nor U12554 (N_12554,N_12240,N_12271);
xnor U12555 (N_12555,N_12116,N_12448);
xor U12556 (N_12556,N_12111,N_12400);
nand U12557 (N_12557,N_11900,N_12156);
nor U12558 (N_12558,N_12230,N_12316);
or U12559 (N_12559,N_11890,N_11975);
nor U12560 (N_12560,N_12080,N_12266);
or U12561 (N_12561,N_11884,N_11926);
nand U12562 (N_12562,N_12032,N_12431);
and U12563 (N_12563,N_12085,N_12164);
or U12564 (N_12564,N_12137,N_12076);
or U12565 (N_12565,N_11990,N_11944);
and U12566 (N_12566,N_12288,N_12425);
and U12567 (N_12567,N_12459,N_12366);
xor U12568 (N_12568,N_12309,N_12246);
nand U12569 (N_12569,N_12208,N_12296);
and U12570 (N_12570,N_11888,N_12359);
or U12571 (N_12571,N_12126,N_11902);
nor U12572 (N_12572,N_12248,N_12231);
xnor U12573 (N_12573,N_12033,N_12154);
and U12574 (N_12574,N_11922,N_12093);
and U12575 (N_12575,N_12144,N_11937);
xnor U12576 (N_12576,N_12435,N_12451);
and U12577 (N_12577,N_11881,N_11887);
nand U12578 (N_12578,N_11914,N_11991);
nand U12579 (N_12579,N_12323,N_12377);
nor U12580 (N_12580,N_12216,N_12002);
and U12581 (N_12581,N_12104,N_12281);
nor U12582 (N_12582,N_12026,N_12499);
or U12583 (N_12583,N_12110,N_12264);
nand U12584 (N_12584,N_12205,N_12455);
nor U12585 (N_12585,N_11886,N_12061);
nand U12586 (N_12586,N_12207,N_12311);
nand U12587 (N_12587,N_12415,N_12487);
nand U12588 (N_12588,N_12212,N_11906);
and U12589 (N_12589,N_12338,N_12120);
or U12590 (N_12590,N_12491,N_12457);
xnor U12591 (N_12591,N_11903,N_12232);
and U12592 (N_12592,N_12064,N_11925);
xor U12593 (N_12593,N_12493,N_12155);
nor U12594 (N_12594,N_12001,N_11909);
xnor U12595 (N_12595,N_12115,N_12362);
or U12596 (N_12596,N_12343,N_12424);
nand U12597 (N_12597,N_11939,N_12194);
nor U12598 (N_12598,N_12371,N_12461);
or U12599 (N_12599,N_12473,N_12058);
nand U12600 (N_12600,N_11883,N_12160);
xor U12601 (N_12601,N_11954,N_12139);
or U12602 (N_12602,N_12284,N_12152);
nor U12603 (N_12603,N_12317,N_12008);
and U12604 (N_12604,N_11904,N_12339);
or U12605 (N_12605,N_11882,N_11996);
and U12606 (N_12606,N_12123,N_12218);
and U12607 (N_12607,N_12304,N_12322);
or U12608 (N_12608,N_12267,N_12276);
or U12609 (N_12609,N_12128,N_12245);
or U12610 (N_12610,N_11987,N_11878);
nand U12611 (N_12611,N_12285,N_12042);
and U12612 (N_12612,N_11994,N_12199);
nand U12613 (N_12613,N_11945,N_11963);
nand U12614 (N_12614,N_12050,N_11971);
nand U12615 (N_12615,N_11962,N_11889);
nor U12616 (N_12616,N_12150,N_11912);
nor U12617 (N_12617,N_11921,N_12314);
or U12618 (N_12618,N_12188,N_12013);
and U12619 (N_12619,N_12278,N_11985);
and U12620 (N_12620,N_11927,N_12054);
and U12621 (N_12621,N_11898,N_12127);
and U12622 (N_12622,N_11958,N_12022);
nand U12623 (N_12623,N_12395,N_11913);
nand U12624 (N_12624,N_11984,N_11919);
or U12625 (N_12625,N_12492,N_12037);
and U12626 (N_12626,N_12202,N_12125);
or U12627 (N_12627,N_11899,N_12464);
xnor U12628 (N_12628,N_12201,N_12004);
or U12629 (N_12629,N_12373,N_12094);
nand U12630 (N_12630,N_12081,N_12067);
or U12631 (N_12631,N_12049,N_11875);
nor U12632 (N_12632,N_12335,N_12169);
or U12633 (N_12633,N_12153,N_12069);
and U12634 (N_12634,N_11997,N_12387);
nand U12635 (N_12635,N_11955,N_12372);
xor U12636 (N_12636,N_12402,N_11988);
and U12637 (N_12637,N_12162,N_12141);
nand U12638 (N_12638,N_12119,N_12062);
or U12639 (N_12639,N_12073,N_12357);
or U12640 (N_12640,N_12157,N_11935);
nand U12641 (N_12641,N_12319,N_12177);
or U12642 (N_12642,N_12439,N_12244);
nor U12643 (N_12643,N_12135,N_12003);
and U12644 (N_12644,N_12109,N_12047);
xnor U12645 (N_12645,N_12180,N_12018);
or U12646 (N_12646,N_12409,N_12252);
nor U12647 (N_12647,N_11976,N_12191);
nand U12648 (N_12648,N_12363,N_12453);
nor U12649 (N_12649,N_12433,N_12333);
nor U12650 (N_12650,N_12025,N_12358);
nor U12651 (N_12651,N_12254,N_12027);
xnor U12652 (N_12652,N_11923,N_12163);
nand U12653 (N_12653,N_12189,N_12436);
nand U12654 (N_12654,N_12105,N_12465);
and U12655 (N_12655,N_12057,N_12039);
and U12656 (N_12656,N_12347,N_12390);
nor U12657 (N_12657,N_11970,N_12068);
or U12658 (N_12658,N_12481,N_12421);
or U12659 (N_12659,N_12426,N_12211);
nor U12660 (N_12660,N_12172,N_12122);
xnor U12661 (N_12661,N_12313,N_11893);
or U12662 (N_12662,N_12303,N_12134);
or U12663 (N_12663,N_12083,N_12352);
xor U12664 (N_12664,N_12416,N_12417);
or U12665 (N_12665,N_12235,N_12412);
xor U12666 (N_12666,N_12301,N_12381);
nor U12667 (N_12667,N_11960,N_12098);
and U12668 (N_12668,N_12055,N_12171);
and U12669 (N_12669,N_12223,N_12114);
nand U12670 (N_12670,N_11891,N_12149);
or U12671 (N_12671,N_11981,N_12392);
xnor U12672 (N_12672,N_12000,N_11924);
and U12673 (N_12673,N_12364,N_12495);
and U12674 (N_12674,N_12437,N_12498);
and U12675 (N_12675,N_12029,N_12043);
nor U12676 (N_12676,N_12484,N_12106);
and U12677 (N_12677,N_11993,N_12091);
nor U12678 (N_12678,N_12118,N_12178);
and U12679 (N_12679,N_12325,N_12082);
nand U12680 (N_12680,N_12321,N_11876);
nor U12681 (N_12681,N_11877,N_11974);
nor U12682 (N_12682,N_12397,N_11978);
or U12683 (N_12683,N_12195,N_11892);
nor U12684 (N_12684,N_11949,N_12290);
nor U12685 (N_12685,N_12183,N_12253);
or U12686 (N_12686,N_12203,N_12401);
xor U12687 (N_12687,N_12048,N_12053);
nor U12688 (N_12688,N_12251,N_12247);
and U12689 (N_12689,N_12132,N_11930);
and U12690 (N_12690,N_12197,N_12088);
nor U12691 (N_12691,N_11896,N_12385);
or U12692 (N_12692,N_12258,N_12075);
nor U12693 (N_12693,N_12249,N_12428);
nand U12694 (N_12694,N_12147,N_11934);
or U12695 (N_12695,N_12221,N_11933);
and U12696 (N_12696,N_12012,N_12117);
and U12697 (N_12697,N_12151,N_12419);
nor U12698 (N_12698,N_12066,N_11968);
nand U12699 (N_12699,N_12370,N_12384);
xnor U12700 (N_12700,N_12447,N_12476);
and U12701 (N_12701,N_12349,N_12173);
xnor U12702 (N_12702,N_12023,N_12222);
and U12703 (N_12703,N_12332,N_11901);
xor U12704 (N_12704,N_12365,N_12086);
and U12705 (N_12705,N_12463,N_12097);
xnor U12706 (N_12706,N_12382,N_12336);
nor U12707 (N_12707,N_12063,N_12443);
and U12708 (N_12708,N_12427,N_12291);
or U12709 (N_12709,N_12226,N_12326);
nand U12710 (N_12710,N_12077,N_12174);
or U12711 (N_12711,N_12185,N_12471);
or U12712 (N_12712,N_12297,N_12467);
and U12713 (N_12713,N_12410,N_12444);
or U12714 (N_12714,N_12488,N_11953);
nor U12715 (N_12715,N_12072,N_12005);
or U12716 (N_12716,N_12224,N_11951);
nor U12717 (N_12717,N_12130,N_12438);
and U12718 (N_12718,N_12292,N_12182);
nand U12719 (N_12719,N_12140,N_12413);
xor U12720 (N_12720,N_11895,N_11947);
xnor U12721 (N_12721,N_12103,N_12307);
nand U12722 (N_12722,N_12015,N_12059);
or U12723 (N_12723,N_12340,N_12121);
and U12724 (N_12724,N_12096,N_11943);
nor U12725 (N_12725,N_12462,N_11966);
and U12726 (N_12726,N_11973,N_12478);
nor U12727 (N_12727,N_11910,N_12084);
nor U12728 (N_12728,N_12060,N_12456);
or U12729 (N_12729,N_12108,N_11916);
or U12730 (N_12730,N_12441,N_12295);
nor U12731 (N_12731,N_12391,N_11948);
or U12732 (N_12732,N_11979,N_12079);
nand U12733 (N_12733,N_12198,N_12265);
and U12734 (N_12734,N_12192,N_12329);
xor U12735 (N_12735,N_11940,N_12056);
or U12736 (N_12736,N_12031,N_12275);
and U12737 (N_12737,N_11905,N_12494);
and U12738 (N_12738,N_12394,N_12442);
nor U12739 (N_12739,N_12449,N_12466);
or U12740 (N_12740,N_12383,N_12489);
nand U12741 (N_12741,N_12181,N_12129);
nand U12742 (N_12742,N_12007,N_12386);
and U12743 (N_12743,N_11938,N_12405);
or U12744 (N_12744,N_12367,N_12274);
xnor U12745 (N_12745,N_12268,N_12241);
and U12746 (N_12746,N_12186,N_12092);
nor U12747 (N_12747,N_12469,N_12238);
nor U12748 (N_12748,N_12277,N_12213);
nor U12749 (N_12749,N_12020,N_12486);
and U12750 (N_12750,N_12215,N_12269);
or U12751 (N_12751,N_12460,N_12470);
and U12752 (N_12752,N_12483,N_12302);
and U12753 (N_12753,N_12143,N_12346);
and U12754 (N_12754,N_12229,N_11995);
nand U12755 (N_12755,N_12477,N_12328);
and U12756 (N_12756,N_11917,N_12388);
or U12757 (N_12757,N_12200,N_12411);
and U12758 (N_12758,N_12142,N_11956);
nand U12759 (N_12759,N_11897,N_12432);
and U12760 (N_12760,N_12310,N_12324);
nand U12761 (N_12761,N_12044,N_12354);
nand U12762 (N_12762,N_12423,N_12017);
nor U12763 (N_12763,N_12070,N_12312);
or U12764 (N_12764,N_12052,N_12434);
and U12765 (N_12765,N_12334,N_12100);
nor U12766 (N_12766,N_12273,N_12014);
and U12767 (N_12767,N_11918,N_12398);
and U12768 (N_12768,N_12450,N_12360);
nor U12769 (N_12769,N_11920,N_12260);
and U12770 (N_12770,N_12204,N_12036);
xor U12771 (N_12771,N_12331,N_12445);
nor U12772 (N_12772,N_12482,N_12158);
or U12773 (N_12773,N_12403,N_11961);
and U12774 (N_12774,N_12166,N_12170);
xor U12775 (N_12775,N_11908,N_12280);
nor U12776 (N_12776,N_12257,N_12420);
xnor U12777 (N_12777,N_12480,N_12242);
or U12778 (N_12778,N_12206,N_11999);
or U12779 (N_12779,N_12452,N_12009);
nor U12780 (N_12780,N_12145,N_12095);
or U12781 (N_12781,N_12038,N_12356);
nor U12782 (N_12782,N_11992,N_11982);
or U12783 (N_12783,N_11931,N_11929);
or U12784 (N_12784,N_11969,N_12468);
and U12785 (N_12785,N_12263,N_12102);
nand U12786 (N_12786,N_11911,N_12234);
xnor U12787 (N_12787,N_12351,N_12393);
nand U12788 (N_12788,N_12184,N_12374);
nand U12789 (N_12789,N_11894,N_11936);
and U12790 (N_12790,N_11941,N_12131);
xor U12791 (N_12791,N_12293,N_12315);
nand U12792 (N_12792,N_12369,N_11959);
and U12793 (N_12793,N_12490,N_12308);
xnor U12794 (N_12794,N_12376,N_12136);
nand U12795 (N_12795,N_12404,N_12107);
or U12796 (N_12796,N_12446,N_12355);
nor U12797 (N_12797,N_12219,N_12071);
nand U12798 (N_12798,N_11983,N_12261);
nor U12799 (N_12799,N_12041,N_12429);
and U12800 (N_12800,N_11998,N_12217);
nor U12801 (N_12801,N_12146,N_12179);
xor U12802 (N_12802,N_11972,N_12262);
or U12803 (N_12803,N_12112,N_12133);
or U12804 (N_12804,N_12414,N_12375);
and U12805 (N_12805,N_12348,N_12196);
or U12806 (N_12806,N_11952,N_12259);
nor U12807 (N_12807,N_12407,N_12282);
xnor U12808 (N_12808,N_12279,N_12168);
or U12809 (N_12809,N_12283,N_12368);
or U12810 (N_12810,N_12479,N_12341);
nand U12811 (N_12811,N_11957,N_12454);
nor U12812 (N_12812,N_12227,N_12092);
or U12813 (N_12813,N_12286,N_11891);
and U12814 (N_12814,N_11888,N_12003);
or U12815 (N_12815,N_11928,N_12216);
xnor U12816 (N_12816,N_12112,N_12345);
and U12817 (N_12817,N_12033,N_11881);
and U12818 (N_12818,N_12422,N_12227);
nor U12819 (N_12819,N_11887,N_12141);
nand U12820 (N_12820,N_11928,N_12030);
xor U12821 (N_12821,N_12188,N_12448);
or U12822 (N_12822,N_12232,N_12221);
xnor U12823 (N_12823,N_12242,N_12285);
nor U12824 (N_12824,N_12246,N_12234);
and U12825 (N_12825,N_12143,N_12362);
and U12826 (N_12826,N_11901,N_12246);
xor U12827 (N_12827,N_12237,N_12052);
and U12828 (N_12828,N_11935,N_11940);
xnor U12829 (N_12829,N_12219,N_12257);
and U12830 (N_12830,N_11891,N_11995);
nand U12831 (N_12831,N_11964,N_11929);
nor U12832 (N_12832,N_11981,N_11943);
nand U12833 (N_12833,N_12128,N_12472);
nand U12834 (N_12834,N_12155,N_12399);
and U12835 (N_12835,N_12210,N_12062);
nand U12836 (N_12836,N_11936,N_11899);
nor U12837 (N_12837,N_12203,N_12409);
nor U12838 (N_12838,N_12263,N_11976);
and U12839 (N_12839,N_12089,N_12126);
nor U12840 (N_12840,N_12267,N_11969);
xor U12841 (N_12841,N_11921,N_11982);
and U12842 (N_12842,N_11970,N_11888);
and U12843 (N_12843,N_11884,N_12413);
nand U12844 (N_12844,N_12236,N_12016);
nor U12845 (N_12845,N_11941,N_12251);
nand U12846 (N_12846,N_12234,N_12378);
or U12847 (N_12847,N_12436,N_12307);
and U12848 (N_12848,N_12400,N_12020);
nor U12849 (N_12849,N_12362,N_12319);
or U12850 (N_12850,N_12461,N_12036);
xor U12851 (N_12851,N_12176,N_12495);
nor U12852 (N_12852,N_12089,N_12109);
and U12853 (N_12853,N_12105,N_11939);
and U12854 (N_12854,N_11953,N_11903);
nor U12855 (N_12855,N_11902,N_12392);
nand U12856 (N_12856,N_11979,N_12378);
nand U12857 (N_12857,N_12397,N_11900);
or U12858 (N_12858,N_12290,N_12329);
nand U12859 (N_12859,N_11880,N_12057);
nor U12860 (N_12860,N_12211,N_11889);
and U12861 (N_12861,N_12007,N_12443);
or U12862 (N_12862,N_11979,N_12083);
and U12863 (N_12863,N_12133,N_12292);
or U12864 (N_12864,N_12454,N_12242);
nor U12865 (N_12865,N_12053,N_12000);
and U12866 (N_12866,N_12020,N_12309);
and U12867 (N_12867,N_12058,N_12292);
or U12868 (N_12868,N_12198,N_11882);
nand U12869 (N_12869,N_12434,N_12475);
xnor U12870 (N_12870,N_11981,N_11986);
and U12871 (N_12871,N_12430,N_12237);
or U12872 (N_12872,N_11947,N_12106);
nor U12873 (N_12873,N_12291,N_12335);
nor U12874 (N_12874,N_11987,N_12298);
or U12875 (N_12875,N_11953,N_12418);
nor U12876 (N_12876,N_12163,N_12456);
xor U12877 (N_12877,N_12298,N_12235);
and U12878 (N_12878,N_12417,N_12050);
nor U12879 (N_12879,N_11883,N_11992);
nand U12880 (N_12880,N_12084,N_12241);
nor U12881 (N_12881,N_12003,N_12164);
xor U12882 (N_12882,N_12200,N_12375);
nor U12883 (N_12883,N_12025,N_12498);
nor U12884 (N_12884,N_12069,N_12215);
and U12885 (N_12885,N_12138,N_11932);
nand U12886 (N_12886,N_12290,N_11955);
nor U12887 (N_12887,N_12075,N_11891);
and U12888 (N_12888,N_12128,N_11893);
and U12889 (N_12889,N_12063,N_12053);
nand U12890 (N_12890,N_11957,N_11904);
nand U12891 (N_12891,N_11888,N_11989);
xor U12892 (N_12892,N_12258,N_12106);
xnor U12893 (N_12893,N_12432,N_12140);
and U12894 (N_12894,N_11910,N_11900);
nor U12895 (N_12895,N_11881,N_12132);
and U12896 (N_12896,N_12287,N_12296);
nor U12897 (N_12897,N_12177,N_12472);
nor U12898 (N_12898,N_12307,N_12140);
or U12899 (N_12899,N_11922,N_12091);
and U12900 (N_12900,N_12471,N_11879);
and U12901 (N_12901,N_11884,N_12302);
nor U12902 (N_12902,N_12408,N_12343);
and U12903 (N_12903,N_12320,N_12195);
nor U12904 (N_12904,N_11933,N_12276);
and U12905 (N_12905,N_11990,N_11919);
or U12906 (N_12906,N_12472,N_12244);
xor U12907 (N_12907,N_12043,N_11923);
and U12908 (N_12908,N_12010,N_12091);
nand U12909 (N_12909,N_11941,N_12495);
xnor U12910 (N_12910,N_12316,N_12195);
or U12911 (N_12911,N_12295,N_12381);
xor U12912 (N_12912,N_12022,N_12217);
nor U12913 (N_12913,N_12255,N_12007);
and U12914 (N_12914,N_12060,N_12107);
and U12915 (N_12915,N_12307,N_12069);
nor U12916 (N_12916,N_12232,N_12418);
nand U12917 (N_12917,N_12478,N_11994);
nand U12918 (N_12918,N_12100,N_12201);
nand U12919 (N_12919,N_12028,N_12375);
nand U12920 (N_12920,N_12280,N_11998);
and U12921 (N_12921,N_12000,N_12222);
nor U12922 (N_12922,N_12321,N_12016);
or U12923 (N_12923,N_12335,N_12097);
and U12924 (N_12924,N_12140,N_11902);
nor U12925 (N_12925,N_12446,N_12038);
nand U12926 (N_12926,N_12416,N_12442);
and U12927 (N_12927,N_12323,N_12019);
nand U12928 (N_12928,N_12112,N_11895);
and U12929 (N_12929,N_12277,N_11936);
xor U12930 (N_12930,N_11922,N_12023);
and U12931 (N_12931,N_12354,N_12184);
or U12932 (N_12932,N_12342,N_12090);
nor U12933 (N_12933,N_12213,N_12420);
or U12934 (N_12934,N_12319,N_12192);
nand U12935 (N_12935,N_12148,N_12056);
and U12936 (N_12936,N_12296,N_12105);
nor U12937 (N_12937,N_11977,N_12318);
nand U12938 (N_12938,N_12383,N_12089);
nor U12939 (N_12939,N_12247,N_12036);
or U12940 (N_12940,N_12445,N_12218);
nand U12941 (N_12941,N_12135,N_12061);
nand U12942 (N_12942,N_11898,N_12217);
nor U12943 (N_12943,N_12291,N_11991);
or U12944 (N_12944,N_12267,N_12403);
nand U12945 (N_12945,N_12085,N_12436);
xnor U12946 (N_12946,N_12470,N_12480);
nor U12947 (N_12947,N_12359,N_12068);
or U12948 (N_12948,N_12330,N_12468);
nand U12949 (N_12949,N_12239,N_12295);
nor U12950 (N_12950,N_12012,N_11976);
nand U12951 (N_12951,N_12155,N_12022);
and U12952 (N_12952,N_12229,N_12131);
or U12953 (N_12953,N_12286,N_12273);
or U12954 (N_12954,N_11906,N_12439);
nand U12955 (N_12955,N_12278,N_12162);
nor U12956 (N_12956,N_12485,N_11947);
and U12957 (N_12957,N_12087,N_12243);
nand U12958 (N_12958,N_11941,N_12025);
xnor U12959 (N_12959,N_11876,N_12180);
nand U12960 (N_12960,N_12246,N_11920);
xnor U12961 (N_12961,N_12100,N_12269);
nand U12962 (N_12962,N_11923,N_12411);
or U12963 (N_12963,N_11921,N_11928);
and U12964 (N_12964,N_12176,N_12379);
nor U12965 (N_12965,N_12498,N_12233);
and U12966 (N_12966,N_12268,N_12493);
and U12967 (N_12967,N_12266,N_12420);
nand U12968 (N_12968,N_12274,N_12059);
or U12969 (N_12969,N_12196,N_12263);
nor U12970 (N_12970,N_11969,N_12167);
xor U12971 (N_12971,N_12491,N_11963);
xnor U12972 (N_12972,N_11995,N_12281);
xnor U12973 (N_12973,N_12476,N_12175);
or U12974 (N_12974,N_12469,N_12308);
nor U12975 (N_12975,N_11943,N_11914);
and U12976 (N_12976,N_11929,N_12085);
and U12977 (N_12977,N_12122,N_12232);
xnor U12978 (N_12978,N_12303,N_12359);
and U12979 (N_12979,N_12434,N_12437);
nand U12980 (N_12980,N_12273,N_12242);
nor U12981 (N_12981,N_12449,N_11912);
or U12982 (N_12982,N_12041,N_12199);
or U12983 (N_12983,N_12311,N_12167);
and U12984 (N_12984,N_12401,N_12391);
nand U12985 (N_12985,N_11948,N_12059);
xnor U12986 (N_12986,N_12359,N_12013);
and U12987 (N_12987,N_12215,N_11908);
nor U12988 (N_12988,N_12215,N_12083);
nor U12989 (N_12989,N_12367,N_12010);
nand U12990 (N_12990,N_11923,N_12285);
nor U12991 (N_12991,N_12314,N_12312);
and U12992 (N_12992,N_12199,N_12451);
and U12993 (N_12993,N_12252,N_12168);
nor U12994 (N_12994,N_12277,N_12456);
or U12995 (N_12995,N_12070,N_11940);
xnor U12996 (N_12996,N_12384,N_12311);
and U12997 (N_12997,N_11963,N_12494);
nand U12998 (N_12998,N_12338,N_12265);
nor U12999 (N_12999,N_12366,N_12194);
or U13000 (N_13000,N_12255,N_12352);
nor U13001 (N_13001,N_12435,N_12432);
and U13002 (N_13002,N_12465,N_12106);
nor U13003 (N_13003,N_12425,N_12155);
nor U13004 (N_13004,N_12041,N_12121);
xor U13005 (N_13005,N_12374,N_12057);
and U13006 (N_13006,N_12260,N_11934);
nand U13007 (N_13007,N_12159,N_12237);
nand U13008 (N_13008,N_12255,N_12245);
and U13009 (N_13009,N_12114,N_12219);
and U13010 (N_13010,N_12174,N_12139);
nand U13011 (N_13011,N_12174,N_11962);
or U13012 (N_13012,N_12053,N_12006);
nand U13013 (N_13013,N_12294,N_12353);
and U13014 (N_13014,N_12210,N_11904);
or U13015 (N_13015,N_12317,N_12254);
xnor U13016 (N_13016,N_11903,N_12041);
nor U13017 (N_13017,N_11985,N_12321);
nor U13018 (N_13018,N_12109,N_12074);
nor U13019 (N_13019,N_11890,N_12403);
nor U13020 (N_13020,N_11941,N_12252);
and U13021 (N_13021,N_12075,N_12436);
or U13022 (N_13022,N_12009,N_12462);
and U13023 (N_13023,N_12304,N_12315);
nor U13024 (N_13024,N_12487,N_12479);
and U13025 (N_13025,N_12240,N_12043);
xor U13026 (N_13026,N_11876,N_12201);
nor U13027 (N_13027,N_12153,N_12224);
or U13028 (N_13028,N_12077,N_12135);
xor U13029 (N_13029,N_12400,N_12227);
nor U13030 (N_13030,N_12224,N_12051);
nor U13031 (N_13031,N_11905,N_12072);
and U13032 (N_13032,N_12288,N_11990);
nand U13033 (N_13033,N_12400,N_12059);
nand U13034 (N_13034,N_11984,N_12364);
and U13035 (N_13035,N_12426,N_12197);
and U13036 (N_13036,N_12109,N_12277);
nand U13037 (N_13037,N_12147,N_12430);
xnor U13038 (N_13038,N_12033,N_12286);
nand U13039 (N_13039,N_12102,N_12250);
and U13040 (N_13040,N_12330,N_12043);
nor U13041 (N_13041,N_12096,N_11925);
or U13042 (N_13042,N_12009,N_12330);
and U13043 (N_13043,N_12243,N_11875);
or U13044 (N_13044,N_12248,N_12337);
nor U13045 (N_13045,N_12019,N_12149);
and U13046 (N_13046,N_12378,N_12163);
xnor U13047 (N_13047,N_12479,N_12336);
nand U13048 (N_13048,N_12339,N_12010);
nor U13049 (N_13049,N_11936,N_12004);
or U13050 (N_13050,N_12483,N_12176);
nor U13051 (N_13051,N_12207,N_12164);
and U13052 (N_13052,N_11954,N_11974);
nand U13053 (N_13053,N_12018,N_12187);
xnor U13054 (N_13054,N_11935,N_11931);
nand U13055 (N_13055,N_12073,N_12486);
and U13056 (N_13056,N_11930,N_11917);
and U13057 (N_13057,N_12338,N_12401);
nor U13058 (N_13058,N_12436,N_12096);
nor U13059 (N_13059,N_12160,N_12101);
and U13060 (N_13060,N_12002,N_12303);
nand U13061 (N_13061,N_12342,N_12167);
and U13062 (N_13062,N_12215,N_12078);
and U13063 (N_13063,N_11876,N_12249);
nand U13064 (N_13064,N_12135,N_11925);
and U13065 (N_13065,N_12372,N_12155);
and U13066 (N_13066,N_12285,N_11941);
and U13067 (N_13067,N_11966,N_11990);
nor U13068 (N_13068,N_12405,N_12302);
and U13069 (N_13069,N_12319,N_12393);
nor U13070 (N_13070,N_11994,N_12279);
and U13071 (N_13071,N_12467,N_12116);
nor U13072 (N_13072,N_11929,N_12125);
and U13073 (N_13073,N_12227,N_12249);
nand U13074 (N_13074,N_11889,N_12151);
or U13075 (N_13075,N_11959,N_12007);
nor U13076 (N_13076,N_11918,N_11904);
or U13077 (N_13077,N_11914,N_12364);
nor U13078 (N_13078,N_12007,N_12353);
and U13079 (N_13079,N_12447,N_12404);
and U13080 (N_13080,N_12406,N_11974);
xnor U13081 (N_13081,N_12399,N_12081);
or U13082 (N_13082,N_12291,N_11951);
xor U13083 (N_13083,N_11925,N_11955);
and U13084 (N_13084,N_12391,N_12472);
and U13085 (N_13085,N_11967,N_12491);
nor U13086 (N_13086,N_11975,N_12057);
or U13087 (N_13087,N_12333,N_12358);
nand U13088 (N_13088,N_12444,N_11954);
nor U13089 (N_13089,N_12152,N_12317);
or U13090 (N_13090,N_12396,N_12262);
and U13091 (N_13091,N_12455,N_12173);
and U13092 (N_13092,N_12072,N_11963);
and U13093 (N_13093,N_12245,N_12318);
or U13094 (N_13094,N_12341,N_11985);
xnor U13095 (N_13095,N_11985,N_11940);
xnor U13096 (N_13096,N_12236,N_12144);
or U13097 (N_13097,N_12287,N_11933);
xor U13098 (N_13098,N_12448,N_12274);
nand U13099 (N_13099,N_12311,N_12072);
and U13100 (N_13100,N_12077,N_12372);
or U13101 (N_13101,N_12007,N_11941);
nor U13102 (N_13102,N_12157,N_12281);
xor U13103 (N_13103,N_12025,N_12023);
and U13104 (N_13104,N_12366,N_12445);
nand U13105 (N_13105,N_12183,N_11958);
and U13106 (N_13106,N_12410,N_11969);
nor U13107 (N_13107,N_11976,N_12123);
nor U13108 (N_13108,N_12138,N_11901);
and U13109 (N_13109,N_12172,N_12200);
or U13110 (N_13110,N_12487,N_12199);
and U13111 (N_13111,N_12167,N_12473);
and U13112 (N_13112,N_11909,N_12297);
or U13113 (N_13113,N_12372,N_12475);
or U13114 (N_13114,N_12115,N_12306);
or U13115 (N_13115,N_12418,N_12499);
nand U13116 (N_13116,N_12121,N_12332);
or U13117 (N_13117,N_12395,N_12376);
and U13118 (N_13118,N_12024,N_11883);
nand U13119 (N_13119,N_11907,N_12082);
nor U13120 (N_13120,N_12302,N_12499);
and U13121 (N_13121,N_12376,N_12034);
nand U13122 (N_13122,N_12268,N_11981);
or U13123 (N_13123,N_11875,N_12194);
or U13124 (N_13124,N_12380,N_12429);
and U13125 (N_13125,N_12835,N_12867);
nand U13126 (N_13126,N_12989,N_12902);
nor U13127 (N_13127,N_12759,N_13014);
nand U13128 (N_13128,N_12695,N_13005);
or U13129 (N_13129,N_12528,N_13039);
xor U13130 (N_13130,N_12676,N_12859);
or U13131 (N_13131,N_12871,N_12948);
nor U13132 (N_13132,N_12925,N_12951);
nor U13133 (N_13133,N_13070,N_12693);
and U13134 (N_13134,N_12936,N_13058);
nor U13135 (N_13135,N_12796,N_12612);
nor U13136 (N_13136,N_13104,N_12656);
nand U13137 (N_13137,N_12526,N_12779);
nor U13138 (N_13138,N_12884,N_12513);
xor U13139 (N_13139,N_13032,N_13027);
and U13140 (N_13140,N_12511,N_13031);
xor U13141 (N_13141,N_12714,N_12651);
and U13142 (N_13142,N_12805,N_12574);
nand U13143 (N_13143,N_12850,N_12893);
or U13144 (N_13144,N_12719,N_12502);
nor U13145 (N_13145,N_12957,N_12556);
and U13146 (N_13146,N_12545,N_12735);
nand U13147 (N_13147,N_12768,N_13007);
xnor U13148 (N_13148,N_13022,N_12953);
nor U13149 (N_13149,N_12572,N_12892);
and U13150 (N_13150,N_12648,N_12637);
or U13151 (N_13151,N_12803,N_12840);
and U13152 (N_13152,N_12692,N_12827);
and U13153 (N_13153,N_12826,N_12844);
or U13154 (N_13154,N_13048,N_12913);
nand U13155 (N_13155,N_12677,N_12882);
or U13156 (N_13156,N_12602,N_12622);
and U13157 (N_13157,N_12928,N_12865);
nand U13158 (N_13158,N_12571,N_12744);
nand U13159 (N_13159,N_12771,N_13068);
and U13160 (N_13160,N_12565,N_12646);
or U13161 (N_13161,N_13077,N_13119);
nor U13162 (N_13162,N_12518,N_12749);
nor U13163 (N_13163,N_12944,N_12943);
nor U13164 (N_13164,N_13100,N_12649);
and U13165 (N_13165,N_12527,N_12914);
or U13166 (N_13166,N_13090,N_13021);
nand U13167 (N_13167,N_13105,N_12972);
nand U13168 (N_13168,N_12950,N_12689);
or U13169 (N_13169,N_12736,N_12672);
and U13170 (N_13170,N_13061,N_12998);
nor U13171 (N_13171,N_12631,N_12849);
nand U13172 (N_13172,N_12642,N_12561);
or U13173 (N_13173,N_13049,N_12721);
and U13174 (N_13174,N_12563,N_13086);
or U13175 (N_13175,N_13001,N_12924);
nand U13176 (N_13176,N_12723,N_12675);
xnor U13177 (N_13177,N_12878,N_13097);
and U13178 (N_13178,N_12541,N_12600);
nor U13179 (N_13179,N_12916,N_12533);
nor U13180 (N_13180,N_12985,N_12831);
and U13181 (N_13181,N_12746,N_13000);
and U13182 (N_13182,N_12906,N_12911);
nor U13183 (N_13183,N_12555,N_12852);
xnor U13184 (N_13184,N_12727,N_12512);
and U13185 (N_13185,N_13115,N_12806);
nor U13186 (N_13186,N_13095,N_13034);
xnor U13187 (N_13187,N_13063,N_12659);
or U13188 (N_13188,N_13059,N_12996);
nand U13189 (N_13189,N_13121,N_12529);
nand U13190 (N_13190,N_12857,N_12931);
nor U13191 (N_13191,N_12903,N_12783);
or U13192 (N_13192,N_12841,N_12991);
nand U13193 (N_13193,N_13028,N_13062);
and U13194 (N_13194,N_12918,N_12738);
or U13195 (N_13195,N_12596,N_13044);
and U13196 (N_13196,N_12794,N_12980);
and U13197 (N_13197,N_12772,N_13055);
nor U13198 (N_13198,N_13013,N_12769);
nand U13199 (N_13199,N_12807,N_12725);
nand U13200 (N_13200,N_12828,N_12983);
or U13201 (N_13201,N_12718,N_13054);
or U13202 (N_13202,N_12536,N_12897);
or U13203 (N_13203,N_12975,N_13113);
and U13204 (N_13204,N_12605,N_13064);
nand U13205 (N_13205,N_12955,N_12886);
nand U13206 (N_13206,N_13053,N_12930);
xor U13207 (N_13207,N_13025,N_12587);
nand U13208 (N_13208,N_12908,N_12509);
xnor U13209 (N_13209,N_13057,N_12595);
xor U13210 (N_13210,N_12594,N_12653);
xnor U13211 (N_13211,N_12818,N_12926);
and U13212 (N_13212,N_12824,N_13009);
xnor U13213 (N_13213,N_12506,N_12781);
nand U13214 (N_13214,N_13046,N_12687);
and U13215 (N_13215,N_12979,N_13091);
nand U13216 (N_13216,N_12685,N_12822);
or U13217 (N_13217,N_12650,N_13019);
nand U13218 (N_13218,N_12866,N_12701);
and U13219 (N_13219,N_12755,N_12553);
or U13220 (N_13220,N_12775,N_12583);
and U13221 (N_13221,N_12760,N_13037);
and U13222 (N_13222,N_12833,N_12724);
and U13223 (N_13223,N_12858,N_12734);
or U13224 (N_13224,N_12669,N_12907);
or U13225 (N_13225,N_12896,N_13035);
and U13226 (N_13226,N_12811,N_12668);
nor U13227 (N_13227,N_12643,N_12542);
nand U13228 (N_13228,N_12804,N_12728);
nor U13229 (N_13229,N_12793,N_12591);
and U13230 (N_13230,N_12615,N_12764);
nand U13231 (N_13231,N_12638,N_13060);
nand U13232 (N_13232,N_12960,N_12514);
and U13233 (N_13233,N_13082,N_12971);
and U13234 (N_13234,N_12641,N_13109);
and U13235 (N_13235,N_12703,N_13102);
or U13236 (N_13236,N_12750,N_12862);
nor U13237 (N_13237,N_13041,N_12860);
nor U13238 (N_13238,N_12500,N_12854);
and U13239 (N_13239,N_12997,N_12543);
nand U13240 (N_13240,N_12674,N_13067);
and U13241 (N_13241,N_12901,N_12635);
xor U13242 (N_13242,N_12883,N_12763);
nor U13243 (N_13243,N_12654,N_12503);
or U13244 (N_13244,N_12964,N_13008);
nand U13245 (N_13245,N_12510,N_12743);
or U13246 (N_13246,N_12973,N_12851);
and U13247 (N_13247,N_12785,N_13096);
or U13248 (N_13248,N_13020,N_12624);
or U13249 (N_13249,N_12834,N_12620);
or U13250 (N_13250,N_12933,N_12888);
nand U13251 (N_13251,N_13106,N_12832);
nor U13252 (N_13252,N_12993,N_12917);
and U13253 (N_13253,N_12531,N_12702);
nor U13254 (N_13254,N_12715,N_12525);
or U13255 (N_13255,N_12522,N_12956);
xnor U13256 (N_13256,N_13124,N_12912);
or U13257 (N_13257,N_13029,N_13114);
nor U13258 (N_13258,N_12977,N_12532);
xnor U13259 (N_13259,N_13103,N_12778);
nand U13260 (N_13260,N_12853,N_12877);
nand U13261 (N_13261,N_12586,N_12639);
nor U13262 (N_13262,N_12868,N_12552);
nand U13263 (N_13263,N_12966,N_13006);
nand U13264 (N_13264,N_12657,N_12717);
or U13265 (N_13265,N_12589,N_12515);
nand U13266 (N_13266,N_12745,N_12660);
nor U13267 (N_13267,N_12754,N_13072);
or U13268 (N_13268,N_12969,N_13089);
nand U13269 (N_13269,N_12968,N_12699);
nand U13270 (N_13270,N_12776,N_13026);
xor U13271 (N_13271,N_12680,N_12787);
or U13272 (N_13272,N_12588,N_12567);
nor U13273 (N_13273,N_12644,N_12797);
or U13274 (N_13274,N_12710,N_12626);
or U13275 (N_13275,N_13076,N_12974);
nand U13276 (N_13276,N_12756,N_12619);
or U13277 (N_13277,N_12630,N_13112);
nand U13278 (N_13278,N_12726,N_12982);
xor U13279 (N_13279,N_12921,N_12898);
and U13280 (N_13280,N_12945,N_12632);
and U13281 (N_13281,N_12959,N_12821);
or U13282 (N_13282,N_12523,N_12986);
or U13283 (N_13283,N_12863,N_12837);
or U13284 (N_13284,N_12815,N_12549);
nor U13285 (N_13285,N_12946,N_12829);
and U13286 (N_13286,N_12740,N_12795);
or U13287 (N_13287,N_12994,N_12576);
nand U13288 (N_13288,N_12618,N_12729);
nand U13289 (N_13289,N_12873,N_13052);
nand U13290 (N_13290,N_12627,N_13042);
or U13291 (N_13291,N_12904,N_12999);
and U13292 (N_13292,N_12938,N_12604);
and U13293 (N_13293,N_12570,N_12568);
or U13294 (N_13294,N_12560,N_12846);
nor U13295 (N_13295,N_12838,N_13080);
xnor U13296 (N_13296,N_12655,N_12663);
nor U13297 (N_13297,N_13024,N_13123);
nor U13298 (N_13298,N_12872,N_12590);
nor U13299 (N_13299,N_12874,N_12739);
nor U13300 (N_13300,N_12575,N_12582);
nor U13301 (N_13301,N_12603,N_12988);
or U13302 (N_13302,N_12876,N_12616);
or U13303 (N_13303,N_13098,N_12516);
nand U13304 (N_13304,N_12730,N_12580);
and U13305 (N_13305,N_12579,N_12690);
and U13306 (N_13306,N_12606,N_12520);
and U13307 (N_13307,N_12909,N_12667);
nor U13308 (N_13308,N_12809,N_13040);
nand U13309 (N_13309,N_12830,N_12504);
and U13310 (N_13310,N_12934,N_12737);
nor U13311 (N_13311,N_12823,N_12698);
and U13312 (N_13312,N_12847,N_13107);
nand U13313 (N_13313,N_12915,N_12708);
and U13314 (N_13314,N_12961,N_12608);
and U13315 (N_13315,N_12770,N_13081);
or U13316 (N_13316,N_12538,N_13084);
or U13317 (N_13317,N_12990,N_12684);
nand U13318 (N_13318,N_13078,N_13110);
and U13319 (N_13319,N_12890,N_12870);
nand U13320 (N_13320,N_13045,N_12780);
or U13321 (N_13321,N_12885,N_12662);
nor U13322 (N_13322,N_12731,N_12636);
or U13323 (N_13323,N_12761,N_12505);
nor U13324 (N_13324,N_12569,N_13074);
nand U13325 (N_13325,N_12788,N_12798);
or U13326 (N_13326,N_12577,N_13117);
and U13327 (N_13327,N_12601,N_13099);
nor U13328 (N_13328,N_12713,N_13092);
or U13329 (N_13329,N_12962,N_13018);
nor U13330 (N_13330,N_13108,N_13036);
nand U13331 (N_13331,N_12843,N_12941);
nand U13332 (N_13332,N_12634,N_12585);
nor U13333 (N_13333,N_12609,N_12696);
and U13334 (N_13334,N_12704,N_12611);
or U13335 (N_13335,N_12564,N_12810);
nand U13336 (N_13336,N_12597,N_12899);
nand U13337 (N_13337,N_12679,N_12976);
or U13338 (N_13338,N_12774,N_12958);
nand U13339 (N_13339,N_12932,N_12610);
or U13340 (N_13340,N_12645,N_13073);
nor U13341 (N_13341,N_12978,N_13038);
xnor U13342 (N_13342,N_12664,N_12848);
nand U13343 (N_13343,N_13050,N_12963);
xor U13344 (N_13344,N_12995,N_12673);
and U13345 (N_13345,N_12517,N_12939);
nor U13346 (N_13346,N_12954,N_12891);
nor U13347 (N_13347,N_12875,N_13094);
xor U13348 (N_13348,N_12686,N_12540);
and U13349 (N_13349,N_12856,N_12741);
nor U13350 (N_13350,N_12633,N_12666);
nor U13351 (N_13351,N_12598,N_12519);
and U13352 (N_13352,N_12881,N_13016);
or U13353 (N_13353,N_12947,N_12566);
nor U13354 (N_13354,N_12621,N_12905);
or U13355 (N_13355,N_12765,N_12593);
nor U13356 (N_13356,N_12766,N_12927);
nor U13357 (N_13357,N_12919,N_12521);
nor U13358 (N_13358,N_12573,N_13010);
or U13359 (N_13359,N_12751,N_12813);
or U13360 (N_13360,N_12762,N_13023);
or U13361 (N_13361,N_12508,N_12599);
nor U13362 (N_13362,N_12940,N_13030);
nor U13363 (N_13363,N_12697,N_12530);
xnor U13364 (N_13364,N_12551,N_12861);
nand U13365 (N_13365,N_12732,N_12880);
nor U13366 (N_13366,N_12923,N_12709);
and U13367 (N_13367,N_12613,N_12784);
nand U13368 (N_13368,N_12789,N_12691);
xnor U13369 (N_13369,N_13003,N_13051);
xor U13370 (N_13370,N_12681,N_12808);
and U13371 (N_13371,N_12757,N_12665);
nand U13372 (N_13372,N_12711,N_13118);
nand U13373 (N_13373,N_13075,N_12501);
nor U13374 (N_13374,N_12887,N_12817);
or U13375 (N_13375,N_12700,N_12825);
nand U13376 (N_13376,N_12777,N_12836);
or U13377 (N_13377,N_13056,N_12792);
and U13378 (N_13378,N_12922,N_12937);
nand U13379 (N_13379,N_12753,N_12706);
nand U13380 (N_13380,N_12800,N_12790);
nor U13381 (N_13381,N_12658,N_12889);
nor U13382 (N_13382,N_12628,N_13002);
nand U13383 (N_13383,N_12712,N_13111);
and U13384 (N_13384,N_12820,N_13079);
nor U13385 (N_13385,N_12965,N_12647);
and U13386 (N_13386,N_12678,N_12814);
or U13387 (N_13387,N_12623,N_12683);
nor U13388 (N_13388,N_12767,N_12910);
nor U13389 (N_13389,N_12535,N_12537);
or U13390 (N_13390,N_12929,N_12984);
or U13391 (N_13391,N_12949,N_12987);
nand U13392 (N_13392,N_12707,N_12640);
nand U13393 (N_13393,N_12625,N_13120);
and U13394 (N_13394,N_12720,N_12864);
and U13395 (N_13395,N_12970,N_13101);
nand U13396 (N_13396,N_12722,N_12607);
xor U13397 (N_13397,N_12548,N_12845);
or U13398 (N_13398,N_12661,N_12812);
or U13399 (N_13399,N_13116,N_12559);
nand U13400 (N_13400,N_12799,N_12581);
xnor U13401 (N_13401,N_12791,N_12842);
xnor U13402 (N_13402,N_12524,N_13069);
and U13403 (N_13403,N_12747,N_13066);
nand U13404 (N_13404,N_12688,N_12935);
nor U13405 (N_13405,N_12802,N_13085);
or U13406 (N_13406,N_13122,N_12554);
or U13407 (N_13407,N_12748,N_12879);
and U13408 (N_13408,N_13015,N_12546);
xnor U13409 (N_13409,N_12816,N_12562);
nor U13410 (N_13410,N_12952,N_12981);
nor U13411 (N_13411,N_12507,N_12716);
xnor U13412 (N_13412,N_13065,N_12550);
nand U13413 (N_13413,N_12855,N_12705);
or U13414 (N_13414,N_12967,N_12742);
nand U13415 (N_13415,N_12534,N_13033);
and U13416 (N_13416,N_12652,N_12614);
xnor U13417 (N_13417,N_13017,N_12670);
nor U13418 (N_13418,N_12782,N_12682);
nand U13419 (N_13419,N_12592,N_12869);
xnor U13420 (N_13420,N_12629,N_13083);
or U13421 (N_13421,N_12558,N_12773);
and U13422 (N_13422,N_12992,N_13012);
and U13423 (N_13423,N_13093,N_12900);
xnor U13424 (N_13424,N_13087,N_12694);
and U13425 (N_13425,N_12584,N_12557);
or U13426 (N_13426,N_12819,N_13088);
nor U13427 (N_13427,N_12894,N_12578);
nand U13428 (N_13428,N_12617,N_12752);
nand U13429 (N_13429,N_12671,N_12733);
nand U13430 (N_13430,N_13011,N_12786);
nand U13431 (N_13431,N_13047,N_12920);
and U13432 (N_13432,N_12801,N_12839);
or U13433 (N_13433,N_13043,N_12547);
or U13434 (N_13434,N_12758,N_13004);
nand U13435 (N_13435,N_12895,N_13071);
nor U13436 (N_13436,N_12539,N_12942);
and U13437 (N_13437,N_12544,N_12689);
nand U13438 (N_13438,N_13024,N_12597);
and U13439 (N_13439,N_12796,N_12519);
nand U13440 (N_13440,N_12778,N_12643);
or U13441 (N_13441,N_12951,N_12725);
nor U13442 (N_13442,N_12524,N_12541);
nand U13443 (N_13443,N_12595,N_12662);
xnor U13444 (N_13444,N_13038,N_12865);
and U13445 (N_13445,N_12831,N_12774);
and U13446 (N_13446,N_12947,N_12811);
nand U13447 (N_13447,N_12500,N_13088);
xor U13448 (N_13448,N_12600,N_12694);
or U13449 (N_13449,N_12673,N_12778);
nor U13450 (N_13450,N_12835,N_12860);
or U13451 (N_13451,N_12516,N_12746);
nor U13452 (N_13452,N_12689,N_12818);
nand U13453 (N_13453,N_12640,N_13071);
nor U13454 (N_13454,N_12978,N_12921);
or U13455 (N_13455,N_12756,N_12701);
and U13456 (N_13456,N_13040,N_12991);
nand U13457 (N_13457,N_12524,N_12819);
or U13458 (N_13458,N_12618,N_13033);
xnor U13459 (N_13459,N_13009,N_13019);
xnor U13460 (N_13460,N_12588,N_12561);
or U13461 (N_13461,N_12610,N_13006);
nand U13462 (N_13462,N_12502,N_12644);
and U13463 (N_13463,N_12763,N_12884);
nand U13464 (N_13464,N_12938,N_12937);
xnor U13465 (N_13465,N_12837,N_12750);
and U13466 (N_13466,N_12921,N_12764);
and U13467 (N_13467,N_12876,N_12765);
nor U13468 (N_13468,N_12696,N_12695);
nor U13469 (N_13469,N_12758,N_12605);
nand U13470 (N_13470,N_12622,N_12551);
nor U13471 (N_13471,N_13022,N_12513);
nor U13472 (N_13472,N_13056,N_12702);
nand U13473 (N_13473,N_12869,N_12767);
nor U13474 (N_13474,N_12727,N_12809);
nor U13475 (N_13475,N_12756,N_12609);
nand U13476 (N_13476,N_12944,N_13117);
and U13477 (N_13477,N_12900,N_12585);
nand U13478 (N_13478,N_13093,N_12815);
and U13479 (N_13479,N_12587,N_12987);
nor U13480 (N_13480,N_13026,N_13091);
and U13481 (N_13481,N_12707,N_12976);
nand U13482 (N_13482,N_12679,N_12739);
nor U13483 (N_13483,N_12674,N_13042);
or U13484 (N_13484,N_12730,N_13021);
nor U13485 (N_13485,N_13093,N_12813);
xor U13486 (N_13486,N_12985,N_12939);
or U13487 (N_13487,N_12871,N_12587);
nand U13488 (N_13488,N_12585,N_12545);
and U13489 (N_13489,N_12720,N_13092);
nor U13490 (N_13490,N_12890,N_12599);
or U13491 (N_13491,N_12755,N_12551);
or U13492 (N_13492,N_12901,N_12932);
nor U13493 (N_13493,N_12738,N_12519);
or U13494 (N_13494,N_13073,N_12602);
nor U13495 (N_13495,N_12524,N_12555);
or U13496 (N_13496,N_13068,N_12746);
nor U13497 (N_13497,N_13031,N_12747);
xnor U13498 (N_13498,N_12684,N_13053);
or U13499 (N_13499,N_12828,N_13046);
or U13500 (N_13500,N_13037,N_13090);
and U13501 (N_13501,N_12521,N_13027);
nand U13502 (N_13502,N_13009,N_12980);
and U13503 (N_13503,N_12781,N_12852);
and U13504 (N_13504,N_12586,N_13050);
nor U13505 (N_13505,N_12845,N_13033);
nor U13506 (N_13506,N_12956,N_12750);
or U13507 (N_13507,N_12965,N_12663);
or U13508 (N_13508,N_12889,N_13050);
nor U13509 (N_13509,N_13078,N_12529);
and U13510 (N_13510,N_13048,N_12881);
nor U13511 (N_13511,N_13101,N_12643);
and U13512 (N_13512,N_12839,N_12919);
or U13513 (N_13513,N_12955,N_12758);
and U13514 (N_13514,N_12998,N_12895);
or U13515 (N_13515,N_12586,N_12823);
and U13516 (N_13516,N_12970,N_12764);
nor U13517 (N_13517,N_13043,N_12609);
nor U13518 (N_13518,N_12996,N_12879);
nand U13519 (N_13519,N_12645,N_13101);
and U13520 (N_13520,N_12943,N_12903);
and U13521 (N_13521,N_12695,N_13104);
or U13522 (N_13522,N_12848,N_12856);
or U13523 (N_13523,N_12620,N_13028);
and U13524 (N_13524,N_12868,N_12657);
or U13525 (N_13525,N_12675,N_12545);
nor U13526 (N_13526,N_12666,N_12734);
or U13527 (N_13527,N_12723,N_12950);
or U13528 (N_13528,N_12510,N_13022);
nor U13529 (N_13529,N_12819,N_12713);
nand U13530 (N_13530,N_13111,N_12968);
or U13531 (N_13531,N_12757,N_13072);
nand U13532 (N_13532,N_12760,N_12990);
and U13533 (N_13533,N_12938,N_12854);
nor U13534 (N_13534,N_12641,N_12561);
nor U13535 (N_13535,N_12673,N_12833);
nand U13536 (N_13536,N_12584,N_12924);
and U13537 (N_13537,N_12645,N_12656);
nor U13538 (N_13538,N_12943,N_12588);
nand U13539 (N_13539,N_12638,N_12668);
nand U13540 (N_13540,N_12596,N_12873);
nand U13541 (N_13541,N_12561,N_12535);
nand U13542 (N_13542,N_12665,N_12628);
or U13543 (N_13543,N_12586,N_13107);
and U13544 (N_13544,N_12737,N_12663);
nand U13545 (N_13545,N_12504,N_12852);
nand U13546 (N_13546,N_12856,N_12621);
nand U13547 (N_13547,N_12616,N_13058);
and U13548 (N_13548,N_12675,N_12829);
and U13549 (N_13549,N_12991,N_12650);
nor U13550 (N_13550,N_13098,N_12825);
or U13551 (N_13551,N_12547,N_12650);
nand U13552 (N_13552,N_12561,N_12680);
nand U13553 (N_13553,N_13054,N_12674);
or U13554 (N_13554,N_12945,N_12562);
nand U13555 (N_13555,N_12997,N_12763);
nor U13556 (N_13556,N_12899,N_12961);
or U13557 (N_13557,N_12537,N_13049);
or U13558 (N_13558,N_12674,N_12914);
or U13559 (N_13559,N_12767,N_12582);
and U13560 (N_13560,N_12543,N_13038);
and U13561 (N_13561,N_12647,N_12574);
nand U13562 (N_13562,N_13073,N_12899);
or U13563 (N_13563,N_13006,N_13102);
and U13564 (N_13564,N_12639,N_12764);
and U13565 (N_13565,N_12974,N_12773);
nor U13566 (N_13566,N_12719,N_13021);
nand U13567 (N_13567,N_12549,N_13056);
nand U13568 (N_13568,N_12585,N_12626);
nor U13569 (N_13569,N_12591,N_12821);
and U13570 (N_13570,N_12981,N_12734);
nand U13571 (N_13571,N_12977,N_13091);
nand U13572 (N_13572,N_12533,N_12596);
xnor U13573 (N_13573,N_12704,N_13090);
or U13574 (N_13574,N_12842,N_12711);
nand U13575 (N_13575,N_12992,N_12539);
nand U13576 (N_13576,N_13013,N_12844);
or U13577 (N_13577,N_12598,N_13038);
or U13578 (N_13578,N_12768,N_12764);
nor U13579 (N_13579,N_12960,N_12821);
nand U13580 (N_13580,N_12906,N_12927);
nand U13581 (N_13581,N_12551,N_12862);
or U13582 (N_13582,N_12822,N_13038);
nand U13583 (N_13583,N_12759,N_12703);
and U13584 (N_13584,N_13072,N_12758);
nor U13585 (N_13585,N_12723,N_12667);
xor U13586 (N_13586,N_12561,N_12639);
nand U13587 (N_13587,N_12592,N_12657);
and U13588 (N_13588,N_12565,N_13033);
nor U13589 (N_13589,N_12938,N_12987);
nand U13590 (N_13590,N_13005,N_13016);
nand U13591 (N_13591,N_12752,N_13072);
and U13592 (N_13592,N_12506,N_13056);
nor U13593 (N_13593,N_12610,N_12689);
nand U13594 (N_13594,N_12771,N_12651);
and U13595 (N_13595,N_13003,N_12602);
or U13596 (N_13596,N_12501,N_12975);
and U13597 (N_13597,N_12690,N_12824);
or U13598 (N_13598,N_12537,N_12640);
or U13599 (N_13599,N_12983,N_12694);
nand U13600 (N_13600,N_13021,N_12977);
nand U13601 (N_13601,N_12909,N_12638);
nand U13602 (N_13602,N_12632,N_12823);
and U13603 (N_13603,N_13119,N_12952);
or U13604 (N_13604,N_13083,N_12864);
nand U13605 (N_13605,N_12752,N_12887);
or U13606 (N_13606,N_13062,N_12784);
or U13607 (N_13607,N_12518,N_12907);
or U13608 (N_13608,N_12534,N_13042);
nor U13609 (N_13609,N_13071,N_13045);
nor U13610 (N_13610,N_12875,N_12728);
nor U13611 (N_13611,N_12532,N_12825);
nor U13612 (N_13612,N_12642,N_12931);
nor U13613 (N_13613,N_12721,N_12576);
xor U13614 (N_13614,N_12511,N_13068);
or U13615 (N_13615,N_12789,N_12546);
and U13616 (N_13616,N_13032,N_12652);
and U13617 (N_13617,N_12596,N_12599);
and U13618 (N_13618,N_13086,N_12810);
and U13619 (N_13619,N_12626,N_12644);
xor U13620 (N_13620,N_12795,N_12709);
or U13621 (N_13621,N_12723,N_12988);
xnor U13622 (N_13622,N_12615,N_12544);
or U13623 (N_13623,N_12816,N_12995);
xor U13624 (N_13624,N_13038,N_12616);
xnor U13625 (N_13625,N_12735,N_12885);
nor U13626 (N_13626,N_13041,N_12587);
nand U13627 (N_13627,N_13013,N_12569);
or U13628 (N_13628,N_12881,N_12969);
or U13629 (N_13629,N_13105,N_12977);
nor U13630 (N_13630,N_12580,N_12917);
nand U13631 (N_13631,N_12629,N_13108);
and U13632 (N_13632,N_13095,N_13012);
and U13633 (N_13633,N_12868,N_13099);
nor U13634 (N_13634,N_12766,N_12599);
xor U13635 (N_13635,N_13028,N_12534);
xnor U13636 (N_13636,N_12657,N_12826);
and U13637 (N_13637,N_12846,N_12863);
nand U13638 (N_13638,N_12824,N_12513);
nand U13639 (N_13639,N_12758,N_12525);
or U13640 (N_13640,N_12942,N_13077);
nor U13641 (N_13641,N_12832,N_12730);
or U13642 (N_13642,N_12601,N_13117);
nand U13643 (N_13643,N_12738,N_12954);
and U13644 (N_13644,N_13033,N_12874);
and U13645 (N_13645,N_12904,N_12931);
nand U13646 (N_13646,N_12566,N_12941);
or U13647 (N_13647,N_12709,N_12637);
or U13648 (N_13648,N_12762,N_13103);
or U13649 (N_13649,N_12870,N_12852);
nor U13650 (N_13650,N_12588,N_13016);
and U13651 (N_13651,N_12672,N_13014);
or U13652 (N_13652,N_12510,N_12854);
nor U13653 (N_13653,N_13092,N_13004);
nand U13654 (N_13654,N_12574,N_12794);
nand U13655 (N_13655,N_12564,N_12604);
or U13656 (N_13656,N_12801,N_12527);
nand U13657 (N_13657,N_12532,N_12949);
nand U13658 (N_13658,N_12996,N_13047);
nor U13659 (N_13659,N_12995,N_13048);
xnor U13660 (N_13660,N_12755,N_12739);
or U13661 (N_13661,N_13039,N_12943);
nand U13662 (N_13662,N_12562,N_12669);
and U13663 (N_13663,N_12692,N_13044);
or U13664 (N_13664,N_12739,N_12684);
nand U13665 (N_13665,N_12872,N_12798);
or U13666 (N_13666,N_12687,N_12530);
nand U13667 (N_13667,N_12658,N_12849);
nor U13668 (N_13668,N_13056,N_13055);
nor U13669 (N_13669,N_12661,N_12995);
xor U13670 (N_13670,N_13046,N_12775);
or U13671 (N_13671,N_13078,N_12940);
or U13672 (N_13672,N_12733,N_12634);
and U13673 (N_13673,N_12846,N_12592);
or U13674 (N_13674,N_12870,N_12736);
and U13675 (N_13675,N_12840,N_12765);
nand U13676 (N_13676,N_12647,N_12695);
or U13677 (N_13677,N_12966,N_12960);
or U13678 (N_13678,N_12786,N_13100);
nand U13679 (N_13679,N_12554,N_12919);
xnor U13680 (N_13680,N_12779,N_12991);
or U13681 (N_13681,N_12777,N_12870);
and U13682 (N_13682,N_13006,N_12781);
nor U13683 (N_13683,N_12708,N_12552);
nor U13684 (N_13684,N_12955,N_13112);
or U13685 (N_13685,N_13029,N_12604);
xnor U13686 (N_13686,N_12959,N_12624);
xor U13687 (N_13687,N_12918,N_13066);
or U13688 (N_13688,N_12944,N_12680);
and U13689 (N_13689,N_12840,N_12931);
nor U13690 (N_13690,N_12534,N_12727);
or U13691 (N_13691,N_12582,N_12568);
or U13692 (N_13692,N_12741,N_13081);
or U13693 (N_13693,N_12658,N_12546);
and U13694 (N_13694,N_13067,N_13007);
nand U13695 (N_13695,N_13118,N_12907);
or U13696 (N_13696,N_12577,N_12993);
nand U13697 (N_13697,N_12647,N_13071);
nor U13698 (N_13698,N_12823,N_13107);
and U13699 (N_13699,N_12503,N_12878);
or U13700 (N_13700,N_12622,N_12862);
or U13701 (N_13701,N_12968,N_12824);
nand U13702 (N_13702,N_13049,N_12852);
nor U13703 (N_13703,N_12712,N_13115);
or U13704 (N_13704,N_12836,N_12690);
xnor U13705 (N_13705,N_13028,N_12550);
and U13706 (N_13706,N_12896,N_12647);
nand U13707 (N_13707,N_12940,N_13100);
or U13708 (N_13708,N_12843,N_12624);
and U13709 (N_13709,N_12905,N_12573);
and U13710 (N_13710,N_12707,N_12722);
or U13711 (N_13711,N_12995,N_12699);
nand U13712 (N_13712,N_13044,N_13030);
or U13713 (N_13713,N_12812,N_12939);
nor U13714 (N_13714,N_12983,N_13017);
nor U13715 (N_13715,N_12718,N_12592);
and U13716 (N_13716,N_12549,N_12744);
and U13717 (N_13717,N_12514,N_12948);
nand U13718 (N_13718,N_12864,N_13121);
xnor U13719 (N_13719,N_12957,N_12639);
nand U13720 (N_13720,N_12682,N_12633);
nor U13721 (N_13721,N_12950,N_13066);
nor U13722 (N_13722,N_12562,N_13103);
and U13723 (N_13723,N_12640,N_12567);
xnor U13724 (N_13724,N_12775,N_12542);
xnor U13725 (N_13725,N_12841,N_12581);
and U13726 (N_13726,N_12578,N_12823);
xor U13727 (N_13727,N_12582,N_12632);
and U13728 (N_13728,N_12676,N_12758);
and U13729 (N_13729,N_12852,N_12693);
nand U13730 (N_13730,N_13044,N_12748);
nor U13731 (N_13731,N_12510,N_12965);
or U13732 (N_13732,N_12778,N_12541);
nand U13733 (N_13733,N_12775,N_12777);
nand U13734 (N_13734,N_12713,N_12695);
and U13735 (N_13735,N_12948,N_12710);
nor U13736 (N_13736,N_12883,N_12739);
xor U13737 (N_13737,N_12735,N_12911);
nor U13738 (N_13738,N_12829,N_13084);
or U13739 (N_13739,N_12640,N_12626);
and U13740 (N_13740,N_13056,N_12747);
and U13741 (N_13741,N_13062,N_12810);
and U13742 (N_13742,N_12866,N_12811);
or U13743 (N_13743,N_12885,N_13087);
nand U13744 (N_13744,N_12622,N_12505);
nand U13745 (N_13745,N_13044,N_12632);
and U13746 (N_13746,N_12552,N_12659);
nor U13747 (N_13747,N_12975,N_12854);
nor U13748 (N_13748,N_12799,N_12891);
and U13749 (N_13749,N_12531,N_12542);
nor U13750 (N_13750,N_13271,N_13699);
nor U13751 (N_13751,N_13673,N_13608);
or U13752 (N_13752,N_13712,N_13331);
xor U13753 (N_13753,N_13586,N_13596);
and U13754 (N_13754,N_13411,N_13487);
nor U13755 (N_13755,N_13383,N_13664);
xor U13756 (N_13756,N_13474,N_13234);
and U13757 (N_13757,N_13501,N_13626);
nor U13758 (N_13758,N_13523,N_13723);
or U13759 (N_13759,N_13389,N_13578);
nor U13760 (N_13760,N_13283,N_13440);
xor U13761 (N_13761,N_13486,N_13278);
nor U13762 (N_13762,N_13714,N_13306);
and U13763 (N_13763,N_13311,N_13293);
or U13764 (N_13764,N_13679,N_13238);
nor U13765 (N_13765,N_13345,N_13576);
nand U13766 (N_13766,N_13162,N_13453);
or U13767 (N_13767,N_13659,N_13263);
nor U13768 (N_13768,N_13669,N_13320);
xor U13769 (N_13769,N_13400,N_13211);
nor U13770 (N_13770,N_13177,N_13294);
and U13771 (N_13771,N_13488,N_13197);
or U13772 (N_13772,N_13549,N_13734);
xnor U13773 (N_13773,N_13393,N_13359);
or U13774 (N_13774,N_13404,N_13392);
nor U13775 (N_13775,N_13468,N_13705);
nand U13776 (N_13776,N_13460,N_13715);
nand U13777 (N_13777,N_13507,N_13192);
nand U13778 (N_13778,N_13451,N_13250);
or U13779 (N_13779,N_13713,N_13328);
or U13780 (N_13780,N_13581,N_13567);
or U13781 (N_13781,N_13701,N_13377);
nand U13782 (N_13782,N_13461,N_13255);
or U13783 (N_13783,N_13550,N_13357);
or U13784 (N_13784,N_13738,N_13204);
and U13785 (N_13785,N_13671,N_13195);
nand U13786 (N_13786,N_13351,N_13735);
xor U13787 (N_13787,N_13141,N_13387);
and U13788 (N_13788,N_13744,N_13539);
and U13789 (N_13789,N_13399,N_13401);
nor U13790 (N_13790,N_13741,N_13180);
nor U13791 (N_13791,N_13533,N_13483);
or U13792 (N_13792,N_13277,N_13171);
nor U13793 (N_13793,N_13559,N_13482);
nand U13794 (N_13794,N_13538,N_13260);
nand U13795 (N_13795,N_13508,N_13134);
and U13796 (N_13796,N_13707,N_13161);
or U13797 (N_13797,N_13290,N_13506);
nor U13798 (N_13798,N_13609,N_13340);
xor U13799 (N_13799,N_13259,N_13163);
or U13800 (N_13800,N_13139,N_13412);
nor U13801 (N_13801,N_13381,N_13360);
and U13802 (N_13802,N_13146,N_13144);
nor U13803 (N_13803,N_13739,N_13223);
nand U13804 (N_13804,N_13464,N_13716);
and U13805 (N_13805,N_13480,N_13656);
or U13806 (N_13806,N_13267,N_13555);
or U13807 (N_13807,N_13519,N_13406);
nor U13808 (N_13808,N_13184,N_13225);
nor U13809 (N_13809,N_13649,N_13643);
and U13810 (N_13810,N_13354,N_13529);
nand U13811 (N_13811,N_13231,N_13502);
nor U13812 (N_13812,N_13339,N_13660);
and U13813 (N_13813,N_13215,N_13648);
or U13814 (N_13814,N_13245,N_13428);
xor U13815 (N_13815,N_13446,N_13179);
and U13816 (N_13816,N_13720,N_13711);
nand U13817 (N_13817,N_13235,N_13496);
xor U13818 (N_13818,N_13583,N_13205);
nand U13819 (N_13819,N_13347,N_13686);
nand U13820 (N_13820,N_13329,N_13477);
nand U13821 (N_13821,N_13319,N_13206);
nand U13822 (N_13822,N_13422,N_13418);
and U13823 (N_13823,N_13173,N_13433);
nand U13824 (N_13824,N_13305,N_13587);
or U13825 (N_13825,N_13237,N_13233);
and U13826 (N_13826,N_13644,N_13394);
nand U13827 (N_13827,N_13154,N_13719);
nor U13828 (N_13828,N_13372,N_13749);
nand U13829 (N_13829,N_13532,N_13547);
or U13830 (N_13830,N_13537,N_13491);
nor U13831 (N_13831,N_13125,N_13458);
or U13832 (N_13832,N_13315,N_13288);
and U13833 (N_13833,N_13697,N_13414);
nand U13834 (N_13834,N_13333,N_13456);
nand U13835 (N_13835,N_13261,N_13429);
or U13836 (N_13836,N_13415,N_13694);
nand U13837 (N_13837,N_13747,N_13657);
nor U13838 (N_13838,N_13338,N_13455);
nor U13839 (N_13839,N_13527,N_13438);
and U13840 (N_13840,N_13216,N_13265);
xnor U13841 (N_13841,N_13242,N_13427);
and U13842 (N_13842,N_13217,N_13128);
and U13843 (N_13843,N_13661,N_13654);
nor U13844 (N_13844,N_13615,N_13700);
or U13845 (N_13845,N_13379,N_13236);
xor U13846 (N_13846,N_13187,N_13513);
or U13847 (N_13847,N_13585,N_13356);
nand U13848 (N_13848,N_13280,N_13708);
or U13849 (N_13849,N_13241,N_13680);
or U13850 (N_13850,N_13308,N_13743);
nor U13851 (N_13851,N_13362,N_13317);
and U13852 (N_13852,N_13476,N_13722);
and U13853 (N_13853,N_13639,N_13499);
or U13854 (N_13854,N_13454,N_13425);
nor U13855 (N_13855,N_13510,N_13598);
and U13856 (N_13856,N_13201,N_13678);
or U13857 (N_13857,N_13515,N_13193);
or U13858 (N_13858,N_13129,N_13160);
nand U13859 (N_13859,N_13498,N_13682);
or U13860 (N_13860,N_13588,N_13616);
xnor U13861 (N_13861,N_13405,N_13301);
nand U13862 (N_13862,N_13692,N_13624);
nor U13863 (N_13863,N_13239,N_13191);
nor U13864 (N_13864,N_13419,N_13321);
nand U13865 (N_13865,N_13632,N_13470);
and U13866 (N_13866,N_13565,N_13168);
xor U13867 (N_13867,N_13208,N_13158);
and U13868 (N_13868,N_13542,N_13164);
nand U13869 (N_13869,N_13732,N_13324);
nand U13870 (N_13870,N_13552,N_13346);
nand U13871 (N_13871,N_13309,N_13218);
and U13872 (N_13872,N_13582,N_13509);
nor U13873 (N_13873,N_13426,N_13731);
and U13874 (N_13874,N_13175,N_13230);
and U13875 (N_13875,N_13384,N_13603);
nand U13876 (N_13876,N_13504,N_13570);
and U13877 (N_13877,N_13612,N_13640);
xor U13878 (N_13878,N_13232,N_13316);
or U13879 (N_13879,N_13676,N_13220);
or U13880 (N_13880,N_13485,N_13687);
and U13881 (N_13881,N_13631,N_13558);
nand U13882 (N_13882,N_13449,N_13222);
and U13883 (N_13883,N_13448,N_13652);
nand U13884 (N_13884,N_13181,N_13672);
or U13885 (N_13885,N_13416,N_13326);
nand U13886 (N_13886,N_13209,N_13376);
nand U13887 (N_13887,N_13736,N_13580);
nor U13888 (N_13888,N_13430,N_13363);
nand U13889 (N_13889,N_13170,N_13172);
and U13890 (N_13890,N_13268,N_13295);
nor U13891 (N_13891,N_13467,N_13619);
and U13892 (N_13892,N_13681,N_13138);
and U13893 (N_13893,N_13266,N_13614);
nor U13894 (N_13894,N_13437,N_13473);
nor U13895 (N_13895,N_13133,N_13590);
or U13896 (N_13896,N_13410,N_13688);
xnor U13897 (N_13897,N_13248,N_13584);
nor U13898 (N_13898,N_13421,N_13490);
nor U13899 (N_13899,N_13434,N_13322);
or U13900 (N_13900,N_13489,N_13365);
and U13901 (N_13901,N_13221,N_13505);
nand U13902 (N_13902,N_13579,N_13332);
nor U13903 (N_13903,N_13252,N_13691);
and U13904 (N_13904,N_13748,N_13742);
or U13905 (N_13905,N_13435,N_13469);
and U13906 (N_13906,N_13127,N_13155);
nand U13907 (N_13907,N_13622,N_13495);
or U13908 (N_13908,N_13167,N_13314);
nand U13909 (N_13909,N_13207,N_13174);
xnor U13910 (N_13910,N_13642,N_13497);
nand U13911 (N_13911,N_13257,N_13641);
and U13912 (N_13912,N_13546,N_13471);
nand U13913 (N_13913,N_13289,N_13541);
nor U13914 (N_13914,N_13229,N_13663);
nor U13915 (N_13915,N_13169,N_13465);
and U13916 (N_13916,N_13459,N_13685);
and U13917 (N_13917,N_13275,N_13299);
and U13918 (N_13918,N_13287,N_13284);
nor U13919 (N_13919,N_13307,N_13620);
and U13920 (N_13920,N_13249,N_13545);
or U13921 (N_13921,N_13408,N_13402);
nand U13922 (N_13922,N_13272,N_13517);
nor U13923 (N_13923,N_13264,N_13397);
or U13924 (N_13924,N_13452,N_13516);
nor U13925 (N_13925,N_13373,N_13247);
nor U13926 (N_13926,N_13156,N_13244);
and U13927 (N_13927,N_13636,N_13481);
and U13928 (N_13928,N_13746,N_13591);
nand U13929 (N_13929,N_13251,N_13343);
and U13930 (N_13930,N_13296,N_13457);
and U13931 (N_13931,N_13226,N_13213);
nor U13932 (N_13932,N_13728,N_13466);
or U13933 (N_13933,N_13274,N_13514);
xnor U13934 (N_13934,N_13613,N_13536);
nand U13935 (N_13935,N_13605,N_13361);
nor U13936 (N_13936,N_13599,N_13703);
and U13937 (N_13937,N_13634,N_13382);
or U13938 (N_13938,N_13186,N_13441);
nor U13939 (N_13939,N_13159,N_13553);
xnor U13940 (N_13940,N_13395,N_13745);
nand U13941 (N_13941,N_13407,N_13646);
and U13942 (N_13942,N_13183,N_13548);
xnor U13943 (N_13943,N_13135,N_13645);
nor U13944 (N_13944,N_13291,N_13302);
or U13945 (N_13945,N_13534,N_13610);
nor U13946 (N_13946,N_13655,N_13704);
nor U13947 (N_13947,N_13653,N_13721);
nor U13948 (N_13948,N_13531,N_13572);
or U13949 (N_13949,N_13262,N_13604);
or U13950 (N_13950,N_13729,N_13358);
and U13951 (N_13951,N_13203,N_13413);
nand U13952 (N_13952,N_13386,N_13684);
or U13953 (N_13953,N_13355,N_13352);
nand U13954 (N_13954,N_13151,N_13409);
xor U13955 (N_13955,N_13518,N_13442);
or U13956 (N_13956,N_13450,N_13554);
nor U13957 (N_13957,N_13285,N_13371);
or U13958 (N_13958,N_13182,N_13601);
or U13959 (N_13959,N_13630,N_13512);
nor U13960 (N_13960,N_13668,N_13142);
nand U13961 (N_13961,N_13188,N_13165);
xor U13962 (N_13962,N_13327,N_13618);
xnor U13963 (N_13963,N_13369,N_13617);
and U13964 (N_13964,N_13540,N_13677);
nand U13965 (N_13965,N_13606,N_13132);
and U13966 (N_13966,N_13424,N_13330);
and U13967 (N_13967,N_13258,N_13185);
xnor U13968 (N_13968,N_13143,N_13313);
nor U13969 (N_13969,N_13312,N_13297);
nor U13970 (N_13970,N_13562,N_13420);
nand U13971 (N_13971,N_13349,N_13417);
and U13972 (N_13972,N_13292,N_13628);
and U13973 (N_13973,N_13256,N_13202);
and U13974 (N_13974,N_13350,N_13157);
and U13975 (N_13975,N_13544,N_13635);
or U13976 (N_13976,N_13318,N_13368);
and U13977 (N_13977,N_13398,N_13600);
or U13978 (N_13978,N_13166,N_13637);
xnor U13979 (N_13979,N_13503,N_13569);
xnor U13980 (N_13980,N_13666,N_13693);
xnor U13981 (N_13981,N_13432,N_13131);
or U13982 (N_13982,N_13323,N_13335);
and U13983 (N_13983,N_13623,N_13589);
and U13984 (N_13984,N_13214,N_13391);
nand U13985 (N_13985,N_13243,N_13575);
and U13986 (N_13986,N_13269,N_13445);
nand U13987 (N_13987,N_13560,N_13147);
and U13988 (N_13988,N_13650,N_13690);
or U13989 (N_13989,N_13303,N_13484);
xnor U13990 (N_13990,N_13136,N_13336);
nor U13991 (N_13991,N_13279,N_13710);
and U13992 (N_13992,N_13520,N_13210);
or U13993 (N_13993,N_13726,N_13334);
nand U13994 (N_13994,N_13190,N_13563);
and U13995 (N_13995,N_13629,N_13219);
and U13996 (N_13996,N_13689,N_13246);
or U13997 (N_13997,N_13494,N_13447);
nand U13998 (N_13998,N_13436,N_13281);
nand U13999 (N_13999,N_13557,N_13286);
nor U14000 (N_14000,N_13196,N_13390);
xnor U14001 (N_14001,N_13150,N_13730);
and U14002 (N_14002,N_13276,N_13385);
xor U14003 (N_14003,N_13727,N_13638);
xnor U14004 (N_14004,N_13152,N_13592);
and U14005 (N_14005,N_13176,N_13633);
and U14006 (N_14006,N_13366,N_13444);
xnor U14007 (N_14007,N_13702,N_13594);
and U14008 (N_14008,N_13198,N_13607);
or U14009 (N_14009,N_13149,N_13667);
nor U14010 (N_14010,N_13725,N_13200);
and U14011 (N_14011,N_13602,N_13556);
nand U14012 (N_14012,N_13240,N_13577);
nand U14013 (N_14013,N_13228,N_13621);
and U14014 (N_14014,N_13479,N_13227);
nor U14015 (N_14015,N_13528,N_13443);
or U14016 (N_14016,N_13337,N_13270);
or U14017 (N_14017,N_13310,N_13611);
nand U14018 (N_14018,N_13493,N_13137);
or U14019 (N_14019,N_13593,N_13140);
nand U14020 (N_14020,N_13717,N_13380);
nand U14021 (N_14021,N_13737,N_13375);
or U14022 (N_14022,N_13253,N_13472);
xor U14023 (N_14023,N_13574,N_13478);
or U14024 (N_14024,N_13683,N_13378);
and U14025 (N_14025,N_13463,N_13665);
xor U14026 (N_14026,N_13199,N_13696);
or U14027 (N_14027,N_13733,N_13595);
and U14028 (N_14028,N_13530,N_13396);
xnor U14029 (N_14029,N_13740,N_13364);
and U14030 (N_14030,N_13282,N_13462);
or U14031 (N_14031,N_13662,N_13526);
or U14032 (N_14032,N_13706,N_13675);
nor U14033 (N_14033,N_13153,N_13625);
and U14034 (N_14034,N_13194,N_13178);
nand U14035 (N_14035,N_13423,N_13130);
nor U14036 (N_14036,N_13374,N_13148);
or U14037 (N_14037,N_13254,N_13370);
nor U14038 (N_14038,N_13658,N_13597);
or U14039 (N_14039,N_13348,N_13670);
xnor U14040 (N_14040,N_13524,N_13525);
or U14041 (N_14041,N_13189,N_13145);
nor U14042 (N_14042,N_13627,N_13431);
or U14043 (N_14043,N_13300,N_13344);
nand U14044 (N_14044,N_13475,N_13561);
and U14045 (N_14045,N_13212,N_13367);
nand U14046 (N_14046,N_13724,N_13353);
xnor U14047 (N_14047,N_13674,N_13325);
or U14048 (N_14048,N_13573,N_13388);
and U14049 (N_14049,N_13224,N_13298);
xnor U14050 (N_14050,N_13566,N_13511);
nor U14051 (N_14051,N_13718,N_13304);
or U14052 (N_14052,N_13651,N_13695);
or U14053 (N_14053,N_13709,N_13342);
nor U14054 (N_14054,N_13698,N_13551);
or U14055 (N_14055,N_13341,N_13126);
nor U14056 (N_14056,N_13273,N_13535);
nand U14057 (N_14057,N_13500,N_13492);
nor U14058 (N_14058,N_13543,N_13439);
and U14059 (N_14059,N_13571,N_13647);
nand U14060 (N_14060,N_13521,N_13564);
nor U14061 (N_14061,N_13568,N_13403);
nand U14062 (N_14062,N_13522,N_13697);
nor U14063 (N_14063,N_13342,N_13546);
or U14064 (N_14064,N_13714,N_13330);
nor U14065 (N_14065,N_13708,N_13149);
and U14066 (N_14066,N_13664,N_13330);
nand U14067 (N_14067,N_13359,N_13152);
xor U14068 (N_14068,N_13422,N_13467);
nand U14069 (N_14069,N_13501,N_13668);
nor U14070 (N_14070,N_13369,N_13142);
xnor U14071 (N_14071,N_13374,N_13462);
and U14072 (N_14072,N_13706,N_13352);
or U14073 (N_14073,N_13708,N_13524);
xnor U14074 (N_14074,N_13144,N_13467);
and U14075 (N_14075,N_13694,N_13609);
xnor U14076 (N_14076,N_13471,N_13658);
xor U14077 (N_14077,N_13503,N_13222);
and U14078 (N_14078,N_13191,N_13746);
nand U14079 (N_14079,N_13604,N_13531);
or U14080 (N_14080,N_13444,N_13159);
and U14081 (N_14081,N_13137,N_13685);
nor U14082 (N_14082,N_13731,N_13727);
and U14083 (N_14083,N_13355,N_13532);
xnor U14084 (N_14084,N_13512,N_13473);
xnor U14085 (N_14085,N_13724,N_13537);
nor U14086 (N_14086,N_13554,N_13491);
or U14087 (N_14087,N_13165,N_13417);
nand U14088 (N_14088,N_13173,N_13693);
or U14089 (N_14089,N_13357,N_13254);
and U14090 (N_14090,N_13333,N_13519);
and U14091 (N_14091,N_13243,N_13326);
nor U14092 (N_14092,N_13310,N_13671);
and U14093 (N_14093,N_13249,N_13207);
or U14094 (N_14094,N_13357,N_13470);
or U14095 (N_14095,N_13456,N_13509);
nor U14096 (N_14096,N_13256,N_13406);
nand U14097 (N_14097,N_13475,N_13298);
or U14098 (N_14098,N_13465,N_13636);
or U14099 (N_14099,N_13417,N_13521);
nand U14100 (N_14100,N_13177,N_13292);
nor U14101 (N_14101,N_13396,N_13333);
xnor U14102 (N_14102,N_13611,N_13276);
and U14103 (N_14103,N_13262,N_13636);
nor U14104 (N_14104,N_13258,N_13409);
nor U14105 (N_14105,N_13257,N_13561);
and U14106 (N_14106,N_13660,N_13727);
nor U14107 (N_14107,N_13462,N_13243);
or U14108 (N_14108,N_13263,N_13702);
or U14109 (N_14109,N_13290,N_13648);
or U14110 (N_14110,N_13165,N_13344);
nor U14111 (N_14111,N_13199,N_13608);
nand U14112 (N_14112,N_13672,N_13681);
nand U14113 (N_14113,N_13224,N_13288);
xor U14114 (N_14114,N_13567,N_13473);
nor U14115 (N_14115,N_13291,N_13283);
nor U14116 (N_14116,N_13274,N_13496);
or U14117 (N_14117,N_13296,N_13577);
or U14118 (N_14118,N_13174,N_13435);
nand U14119 (N_14119,N_13378,N_13423);
nand U14120 (N_14120,N_13450,N_13725);
nand U14121 (N_14121,N_13491,N_13161);
and U14122 (N_14122,N_13660,N_13502);
nand U14123 (N_14123,N_13316,N_13508);
and U14124 (N_14124,N_13492,N_13364);
xor U14125 (N_14125,N_13519,N_13459);
or U14126 (N_14126,N_13347,N_13240);
xnor U14127 (N_14127,N_13342,N_13656);
and U14128 (N_14128,N_13527,N_13672);
or U14129 (N_14129,N_13601,N_13230);
or U14130 (N_14130,N_13135,N_13339);
or U14131 (N_14131,N_13529,N_13553);
nand U14132 (N_14132,N_13603,N_13249);
nor U14133 (N_14133,N_13611,N_13443);
nand U14134 (N_14134,N_13310,N_13677);
nand U14135 (N_14135,N_13419,N_13341);
or U14136 (N_14136,N_13707,N_13594);
and U14137 (N_14137,N_13375,N_13480);
or U14138 (N_14138,N_13642,N_13354);
nor U14139 (N_14139,N_13670,N_13564);
or U14140 (N_14140,N_13465,N_13407);
nand U14141 (N_14141,N_13711,N_13144);
and U14142 (N_14142,N_13330,N_13677);
or U14143 (N_14143,N_13338,N_13221);
nand U14144 (N_14144,N_13636,N_13634);
and U14145 (N_14145,N_13242,N_13637);
or U14146 (N_14146,N_13221,N_13268);
nor U14147 (N_14147,N_13275,N_13623);
or U14148 (N_14148,N_13502,N_13229);
and U14149 (N_14149,N_13383,N_13316);
and U14150 (N_14150,N_13367,N_13257);
and U14151 (N_14151,N_13669,N_13160);
nor U14152 (N_14152,N_13535,N_13209);
and U14153 (N_14153,N_13726,N_13292);
and U14154 (N_14154,N_13132,N_13430);
nor U14155 (N_14155,N_13440,N_13712);
nor U14156 (N_14156,N_13320,N_13175);
and U14157 (N_14157,N_13561,N_13588);
nor U14158 (N_14158,N_13636,N_13496);
nand U14159 (N_14159,N_13516,N_13618);
nand U14160 (N_14160,N_13608,N_13485);
or U14161 (N_14161,N_13136,N_13285);
and U14162 (N_14162,N_13450,N_13356);
or U14163 (N_14163,N_13140,N_13314);
or U14164 (N_14164,N_13569,N_13689);
and U14165 (N_14165,N_13661,N_13552);
and U14166 (N_14166,N_13611,N_13724);
nand U14167 (N_14167,N_13367,N_13396);
or U14168 (N_14168,N_13229,N_13749);
nor U14169 (N_14169,N_13479,N_13689);
nor U14170 (N_14170,N_13344,N_13353);
nand U14171 (N_14171,N_13422,N_13463);
nor U14172 (N_14172,N_13129,N_13282);
nor U14173 (N_14173,N_13705,N_13561);
or U14174 (N_14174,N_13544,N_13626);
nor U14175 (N_14175,N_13224,N_13688);
or U14176 (N_14176,N_13468,N_13405);
nand U14177 (N_14177,N_13141,N_13205);
nand U14178 (N_14178,N_13593,N_13735);
nor U14179 (N_14179,N_13635,N_13455);
or U14180 (N_14180,N_13144,N_13276);
nand U14181 (N_14181,N_13356,N_13289);
and U14182 (N_14182,N_13311,N_13152);
nor U14183 (N_14183,N_13148,N_13549);
and U14184 (N_14184,N_13343,N_13148);
or U14185 (N_14185,N_13386,N_13625);
nor U14186 (N_14186,N_13553,N_13311);
or U14187 (N_14187,N_13543,N_13731);
and U14188 (N_14188,N_13683,N_13277);
and U14189 (N_14189,N_13304,N_13477);
xor U14190 (N_14190,N_13347,N_13700);
xor U14191 (N_14191,N_13331,N_13404);
or U14192 (N_14192,N_13685,N_13213);
nand U14193 (N_14193,N_13391,N_13553);
nand U14194 (N_14194,N_13679,N_13229);
nand U14195 (N_14195,N_13496,N_13507);
nor U14196 (N_14196,N_13503,N_13397);
nor U14197 (N_14197,N_13512,N_13671);
nor U14198 (N_14198,N_13304,N_13714);
and U14199 (N_14199,N_13553,N_13449);
nor U14200 (N_14200,N_13357,N_13647);
and U14201 (N_14201,N_13336,N_13530);
and U14202 (N_14202,N_13549,N_13687);
nor U14203 (N_14203,N_13604,N_13455);
or U14204 (N_14204,N_13206,N_13463);
xor U14205 (N_14205,N_13311,N_13654);
or U14206 (N_14206,N_13237,N_13677);
nor U14207 (N_14207,N_13391,N_13541);
or U14208 (N_14208,N_13248,N_13140);
nor U14209 (N_14209,N_13622,N_13224);
nand U14210 (N_14210,N_13222,N_13152);
nor U14211 (N_14211,N_13676,N_13210);
nand U14212 (N_14212,N_13556,N_13481);
or U14213 (N_14213,N_13621,N_13327);
or U14214 (N_14214,N_13537,N_13308);
or U14215 (N_14215,N_13393,N_13541);
nand U14216 (N_14216,N_13541,N_13162);
nand U14217 (N_14217,N_13486,N_13287);
nor U14218 (N_14218,N_13447,N_13545);
and U14219 (N_14219,N_13390,N_13537);
nand U14220 (N_14220,N_13660,N_13478);
nor U14221 (N_14221,N_13514,N_13270);
or U14222 (N_14222,N_13592,N_13739);
nand U14223 (N_14223,N_13234,N_13502);
nand U14224 (N_14224,N_13450,N_13713);
nand U14225 (N_14225,N_13171,N_13499);
and U14226 (N_14226,N_13144,N_13507);
or U14227 (N_14227,N_13209,N_13379);
nand U14228 (N_14228,N_13168,N_13194);
or U14229 (N_14229,N_13265,N_13321);
nand U14230 (N_14230,N_13504,N_13466);
and U14231 (N_14231,N_13480,N_13400);
xor U14232 (N_14232,N_13457,N_13420);
or U14233 (N_14233,N_13454,N_13377);
and U14234 (N_14234,N_13454,N_13215);
or U14235 (N_14235,N_13486,N_13243);
nor U14236 (N_14236,N_13349,N_13318);
nor U14237 (N_14237,N_13726,N_13675);
nand U14238 (N_14238,N_13660,N_13151);
nor U14239 (N_14239,N_13189,N_13417);
nand U14240 (N_14240,N_13647,N_13329);
nor U14241 (N_14241,N_13496,N_13564);
nand U14242 (N_14242,N_13713,N_13250);
nand U14243 (N_14243,N_13467,N_13615);
nand U14244 (N_14244,N_13558,N_13563);
nand U14245 (N_14245,N_13259,N_13555);
and U14246 (N_14246,N_13323,N_13724);
and U14247 (N_14247,N_13454,N_13135);
nand U14248 (N_14248,N_13566,N_13573);
or U14249 (N_14249,N_13148,N_13617);
and U14250 (N_14250,N_13381,N_13341);
or U14251 (N_14251,N_13609,N_13581);
nand U14252 (N_14252,N_13672,N_13336);
and U14253 (N_14253,N_13714,N_13205);
xor U14254 (N_14254,N_13164,N_13697);
nor U14255 (N_14255,N_13682,N_13415);
and U14256 (N_14256,N_13341,N_13539);
nand U14257 (N_14257,N_13747,N_13592);
and U14258 (N_14258,N_13566,N_13248);
nor U14259 (N_14259,N_13472,N_13250);
nor U14260 (N_14260,N_13607,N_13171);
and U14261 (N_14261,N_13518,N_13176);
nand U14262 (N_14262,N_13544,N_13481);
or U14263 (N_14263,N_13619,N_13351);
xor U14264 (N_14264,N_13286,N_13281);
and U14265 (N_14265,N_13557,N_13283);
and U14266 (N_14266,N_13454,N_13132);
nor U14267 (N_14267,N_13484,N_13537);
or U14268 (N_14268,N_13560,N_13463);
nor U14269 (N_14269,N_13591,N_13477);
nor U14270 (N_14270,N_13745,N_13310);
and U14271 (N_14271,N_13312,N_13651);
nand U14272 (N_14272,N_13471,N_13140);
nor U14273 (N_14273,N_13324,N_13499);
nor U14274 (N_14274,N_13364,N_13731);
xor U14275 (N_14275,N_13175,N_13227);
nand U14276 (N_14276,N_13233,N_13410);
nor U14277 (N_14277,N_13720,N_13658);
nand U14278 (N_14278,N_13354,N_13356);
nand U14279 (N_14279,N_13209,N_13519);
nor U14280 (N_14280,N_13290,N_13694);
and U14281 (N_14281,N_13466,N_13266);
nor U14282 (N_14282,N_13196,N_13655);
or U14283 (N_14283,N_13742,N_13712);
nand U14284 (N_14284,N_13317,N_13623);
or U14285 (N_14285,N_13407,N_13517);
nand U14286 (N_14286,N_13305,N_13169);
or U14287 (N_14287,N_13243,N_13312);
or U14288 (N_14288,N_13644,N_13652);
nor U14289 (N_14289,N_13201,N_13168);
nor U14290 (N_14290,N_13495,N_13505);
or U14291 (N_14291,N_13581,N_13511);
nand U14292 (N_14292,N_13365,N_13291);
or U14293 (N_14293,N_13294,N_13530);
nand U14294 (N_14294,N_13414,N_13458);
and U14295 (N_14295,N_13357,N_13599);
nor U14296 (N_14296,N_13691,N_13587);
and U14297 (N_14297,N_13525,N_13535);
nor U14298 (N_14298,N_13351,N_13241);
and U14299 (N_14299,N_13523,N_13636);
nand U14300 (N_14300,N_13199,N_13746);
or U14301 (N_14301,N_13162,N_13468);
nand U14302 (N_14302,N_13516,N_13226);
and U14303 (N_14303,N_13522,N_13604);
or U14304 (N_14304,N_13600,N_13743);
or U14305 (N_14305,N_13259,N_13338);
and U14306 (N_14306,N_13635,N_13403);
nor U14307 (N_14307,N_13212,N_13738);
or U14308 (N_14308,N_13575,N_13239);
and U14309 (N_14309,N_13174,N_13635);
and U14310 (N_14310,N_13623,N_13746);
nand U14311 (N_14311,N_13410,N_13513);
nand U14312 (N_14312,N_13278,N_13329);
or U14313 (N_14313,N_13465,N_13389);
nand U14314 (N_14314,N_13718,N_13138);
nand U14315 (N_14315,N_13273,N_13356);
and U14316 (N_14316,N_13193,N_13629);
xor U14317 (N_14317,N_13345,N_13481);
or U14318 (N_14318,N_13256,N_13213);
or U14319 (N_14319,N_13619,N_13605);
nand U14320 (N_14320,N_13429,N_13710);
nand U14321 (N_14321,N_13139,N_13645);
and U14322 (N_14322,N_13690,N_13631);
nand U14323 (N_14323,N_13238,N_13349);
and U14324 (N_14324,N_13167,N_13285);
nor U14325 (N_14325,N_13324,N_13431);
nor U14326 (N_14326,N_13134,N_13519);
nand U14327 (N_14327,N_13228,N_13609);
or U14328 (N_14328,N_13217,N_13483);
or U14329 (N_14329,N_13690,N_13614);
xor U14330 (N_14330,N_13169,N_13463);
nor U14331 (N_14331,N_13394,N_13339);
nand U14332 (N_14332,N_13566,N_13366);
nor U14333 (N_14333,N_13718,N_13539);
xor U14334 (N_14334,N_13608,N_13394);
nor U14335 (N_14335,N_13600,N_13428);
nor U14336 (N_14336,N_13545,N_13312);
xnor U14337 (N_14337,N_13178,N_13343);
or U14338 (N_14338,N_13160,N_13748);
nand U14339 (N_14339,N_13561,N_13638);
nand U14340 (N_14340,N_13180,N_13482);
nand U14341 (N_14341,N_13722,N_13132);
nand U14342 (N_14342,N_13549,N_13407);
nand U14343 (N_14343,N_13249,N_13399);
nor U14344 (N_14344,N_13148,N_13652);
or U14345 (N_14345,N_13344,N_13748);
nand U14346 (N_14346,N_13377,N_13745);
or U14347 (N_14347,N_13580,N_13126);
or U14348 (N_14348,N_13440,N_13344);
nor U14349 (N_14349,N_13492,N_13344);
or U14350 (N_14350,N_13336,N_13231);
nand U14351 (N_14351,N_13477,N_13640);
and U14352 (N_14352,N_13614,N_13681);
or U14353 (N_14353,N_13141,N_13349);
or U14354 (N_14354,N_13241,N_13712);
nor U14355 (N_14355,N_13409,N_13350);
xnor U14356 (N_14356,N_13461,N_13627);
nor U14357 (N_14357,N_13531,N_13221);
xor U14358 (N_14358,N_13316,N_13166);
or U14359 (N_14359,N_13182,N_13448);
or U14360 (N_14360,N_13355,N_13370);
nor U14361 (N_14361,N_13461,N_13396);
xor U14362 (N_14362,N_13291,N_13158);
and U14363 (N_14363,N_13642,N_13237);
or U14364 (N_14364,N_13138,N_13528);
and U14365 (N_14365,N_13678,N_13241);
or U14366 (N_14366,N_13478,N_13654);
nor U14367 (N_14367,N_13703,N_13501);
nor U14368 (N_14368,N_13131,N_13609);
nor U14369 (N_14369,N_13309,N_13281);
nor U14370 (N_14370,N_13251,N_13701);
and U14371 (N_14371,N_13171,N_13461);
nand U14372 (N_14372,N_13412,N_13385);
or U14373 (N_14373,N_13628,N_13726);
nand U14374 (N_14374,N_13288,N_13386);
nor U14375 (N_14375,N_13987,N_14321);
and U14376 (N_14376,N_14334,N_14074);
nor U14377 (N_14377,N_13783,N_14245);
xor U14378 (N_14378,N_14311,N_14136);
or U14379 (N_14379,N_13939,N_13902);
nand U14380 (N_14380,N_14046,N_13839);
and U14381 (N_14381,N_13972,N_14243);
and U14382 (N_14382,N_14331,N_13834);
nor U14383 (N_14383,N_14244,N_13798);
nand U14384 (N_14384,N_14220,N_14366);
nand U14385 (N_14385,N_14352,N_14358);
nor U14386 (N_14386,N_13836,N_14310);
nand U14387 (N_14387,N_14037,N_13921);
nand U14388 (N_14388,N_14284,N_14052);
or U14389 (N_14389,N_13952,N_14302);
nand U14390 (N_14390,N_14105,N_13837);
nor U14391 (N_14391,N_14189,N_13945);
or U14392 (N_14392,N_13754,N_13845);
or U14393 (N_14393,N_13769,N_14278);
and U14394 (N_14394,N_13790,N_14180);
or U14395 (N_14395,N_14003,N_13853);
and U14396 (N_14396,N_14240,N_13793);
or U14397 (N_14397,N_13843,N_13881);
and U14398 (N_14398,N_13991,N_14222);
nand U14399 (N_14399,N_14024,N_14230);
nand U14400 (N_14400,N_14301,N_14210);
and U14401 (N_14401,N_13930,N_14038);
or U14402 (N_14402,N_13918,N_13849);
xnor U14403 (N_14403,N_13944,N_13847);
and U14404 (N_14404,N_14285,N_14147);
nor U14405 (N_14405,N_13878,N_13951);
nor U14406 (N_14406,N_13931,N_14277);
nor U14407 (N_14407,N_14149,N_14354);
nor U14408 (N_14408,N_13919,N_13774);
nor U14409 (N_14409,N_14169,N_13992);
nand U14410 (N_14410,N_14096,N_14257);
nand U14411 (N_14411,N_14344,N_13971);
and U14412 (N_14412,N_14281,N_14077);
or U14413 (N_14413,N_13863,N_14112);
and U14414 (N_14414,N_14247,N_14050);
nor U14415 (N_14415,N_13984,N_14200);
or U14416 (N_14416,N_13810,N_13941);
and U14417 (N_14417,N_14069,N_14282);
xor U14418 (N_14418,N_13994,N_14110);
nor U14419 (N_14419,N_14241,N_14129);
and U14420 (N_14420,N_14097,N_14056);
or U14421 (N_14421,N_13841,N_14261);
and U14422 (N_14422,N_13786,N_13903);
nor U14423 (N_14423,N_13985,N_14005);
nand U14424 (N_14424,N_14330,N_13832);
or U14425 (N_14425,N_14373,N_13755);
and U14426 (N_14426,N_13791,N_13840);
and U14427 (N_14427,N_13990,N_13970);
nor U14428 (N_14428,N_14288,N_14060);
nand U14429 (N_14429,N_13821,N_14130);
nor U14430 (N_14430,N_13898,N_13765);
nand U14431 (N_14431,N_14342,N_14201);
xnor U14432 (N_14432,N_14124,N_13880);
nor U14433 (N_14433,N_14059,N_13823);
or U14434 (N_14434,N_14058,N_14007);
or U14435 (N_14435,N_14323,N_14203);
nor U14436 (N_14436,N_14094,N_13969);
nand U14437 (N_14437,N_14369,N_13768);
xor U14438 (N_14438,N_13901,N_14365);
or U14439 (N_14439,N_14020,N_13956);
nand U14440 (N_14440,N_14175,N_14320);
nor U14441 (N_14441,N_13884,N_14335);
and U14442 (N_14442,N_14192,N_14254);
nor U14443 (N_14443,N_14080,N_14066);
or U14444 (N_14444,N_14085,N_13852);
nand U14445 (N_14445,N_13792,N_14166);
nor U14446 (N_14446,N_13759,N_14049);
xor U14447 (N_14447,N_14040,N_13908);
nor U14448 (N_14448,N_13846,N_14206);
and U14449 (N_14449,N_13982,N_13831);
xnor U14450 (N_14450,N_13996,N_13955);
or U14451 (N_14451,N_14296,N_13932);
and U14452 (N_14452,N_14078,N_14054);
nand U14453 (N_14453,N_14034,N_14100);
or U14454 (N_14454,N_13867,N_13829);
or U14455 (N_14455,N_13789,N_14116);
nor U14456 (N_14456,N_14167,N_14174);
nand U14457 (N_14457,N_14178,N_14044);
or U14458 (N_14458,N_14216,N_14063);
nand U14459 (N_14459,N_14157,N_14231);
or U14460 (N_14460,N_14179,N_14252);
or U14461 (N_14461,N_13914,N_14265);
nor U14462 (N_14462,N_13889,N_14140);
and U14463 (N_14463,N_13804,N_13796);
and U14464 (N_14464,N_14029,N_14120);
or U14465 (N_14465,N_14011,N_13965);
nor U14466 (N_14466,N_14146,N_14099);
or U14467 (N_14467,N_14215,N_14165);
and U14468 (N_14468,N_14187,N_13819);
nand U14469 (N_14469,N_14086,N_14004);
and U14470 (N_14470,N_13865,N_14090);
nor U14471 (N_14471,N_14031,N_14359);
or U14472 (N_14472,N_14304,N_13808);
xor U14473 (N_14473,N_13770,N_13876);
and U14474 (N_14474,N_14164,N_14308);
or U14475 (N_14475,N_14188,N_14101);
nand U14476 (N_14476,N_14028,N_14131);
nand U14477 (N_14477,N_14273,N_13771);
nor U14478 (N_14478,N_14204,N_13983);
nand U14479 (N_14479,N_13882,N_13803);
xor U14480 (N_14480,N_14234,N_14137);
xor U14481 (N_14481,N_14082,N_13957);
nand U14482 (N_14482,N_14324,N_13953);
nor U14483 (N_14483,N_14275,N_13851);
nor U14484 (N_14484,N_13822,N_14111);
nor U14485 (N_14485,N_14009,N_14139);
or U14486 (N_14486,N_14163,N_14289);
nand U14487 (N_14487,N_14306,N_14212);
nor U14488 (N_14488,N_13778,N_14032);
and U14489 (N_14489,N_13784,N_13854);
and U14490 (N_14490,N_14336,N_13864);
nor U14491 (N_14491,N_13871,N_14238);
nand U14492 (N_14492,N_14221,N_14119);
nand U14493 (N_14493,N_13926,N_14318);
nand U14494 (N_14494,N_13891,N_14042);
nand U14495 (N_14495,N_13968,N_13979);
or U14496 (N_14496,N_14012,N_14266);
nor U14497 (N_14497,N_14209,N_14368);
or U14498 (N_14498,N_13824,N_13772);
nor U14499 (N_14499,N_14084,N_13906);
nor U14500 (N_14500,N_13856,N_14154);
nand U14501 (N_14501,N_14195,N_13811);
and U14502 (N_14502,N_14303,N_14172);
or U14503 (N_14503,N_13860,N_14207);
nor U14504 (N_14504,N_14041,N_13937);
nand U14505 (N_14505,N_14083,N_13873);
and U14506 (N_14506,N_14143,N_14186);
or U14507 (N_14507,N_14317,N_14271);
nand U14508 (N_14508,N_13758,N_13756);
nand U14509 (N_14509,N_13900,N_14073);
nor U14510 (N_14510,N_14185,N_13927);
and U14511 (N_14511,N_13963,N_14319);
and U14512 (N_14512,N_14098,N_13933);
and U14513 (N_14513,N_14177,N_13869);
nand U14514 (N_14514,N_13879,N_13795);
or U14515 (N_14515,N_14045,N_14332);
and U14516 (N_14516,N_14339,N_13801);
nand U14517 (N_14517,N_14030,N_14064);
nand U14518 (N_14518,N_14333,N_14249);
or U14519 (N_14519,N_13935,N_13805);
nand U14520 (N_14520,N_13775,N_14263);
nor U14521 (N_14521,N_13844,N_14113);
or U14522 (N_14522,N_14162,N_14291);
nor U14523 (N_14523,N_14297,N_14160);
or U14524 (N_14524,N_14269,N_14126);
or U14525 (N_14525,N_14087,N_13830);
nand U14526 (N_14526,N_13895,N_13961);
nand U14527 (N_14527,N_14347,N_13850);
or U14528 (N_14528,N_13875,N_14292);
xnor U14529 (N_14529,N_14251,N_14076);
nand U14530 (N_14530,N_13960,N_14246);
nand U14531 (N_14531,N_14295,N_14202);
and U14532 (N_14532,N_14279,N_13916);
and U14533 (N_14533,N_14138,N_13974);
nor U14534 (N_14534,N_14360,N_14355);
nor U14535 (N_14535,N_14345,N_14115);
or U14536 (N_14536,N_14010,N_13782);
nor U14537 (N_14537,N_13777,N_14190);
nor U14538 (N_14538,N_14270,N_14170);
nor U14539 (N_14539,N_14367,N_14362);
or U14540 (N_14540,N_14351,N_14079);
and U14541 (N_14541,N_13975,N_13998);
and U14542 (N_14542,N_13904,N_13966);
and U14543 (N_14543,N_13973,N_14144);
nand U14544 (N_14544,N_13842,N_14371);
xor U14545 (N_14545,N_13780,N_14218);
nand U14546 (N_14546,N_13807,N_13928);
nand U14547 (N_14547,N_13787,N_14205);
or U14548 (N_14548,N_13802,N_13760);
and U14549 (N_14549,N_13897,N_13870);
nand U14550 (N_14550,N_13779,N_13866);
nor U14551 (N_14551,N_13977,N_14299);
nor U14552 (N_14552,N_14276,N_14305);
or U14553 (N_14553,N_14260,N_14312);
nor U14554 (N_14554,N_14298,N_13936);
and U14555 (N_14555,N_13767,N_13762);
and U14556 (N_14556,N_14196,N_13924);
and U14557 (N_14557,N_13911,N_13923);
or U14558 (N_14558,N_14000,N_13997);
nand U14559 (N_14559,N_14250,N_14316);
or U14560 (N_14560,N_14338,N_13958);
and U14561 (N_14561,N_14280,N_14242);
or U14562 (N_14562,N_14227,N_14017);
nor U14563 (N_14563,N_13999,N_14062);
or U14564 (N_14564,N_14008,N_13828);
or U14565 (N_14565,N_13761,N_13892);
and U14566 (N_14566,N_14364,N_14194);
xor U14567 (N_14567,N_14300,N_13989);
nor U14568 (N_14568,N_14237,N_14363);
nand U14569 (N_14569,N_14264,N_14072);
or U14570 (N_14570,N_14075,N_14141);
xor U14571 (N_14571,N_14307,N_13763);
or U14572 (N_14572,N_13883,N_14026);
or U14573 (N_14573,N_13896,N_13948);
and U14574 (N_14574,N_13964,N_13855);
or U14575 (N_14575,N_14340,N_14152);
nor U14576 (N_14576,N_14006,N_13934);
nand U14577 (N_14577,N_14081,N_14224);
nor U14578 (N_14578,N_13910,N_14374);
nor U14579 (N_14579,N_14106,N_14193);
nand U14580 (N_14580,N_14173,N_13899);
nand U14581 (N_14581,N_13827,N_13885);
or U14582 (N_14582,N_14211,N_14103);
nor U14583 (N_14583,N_13800,N_14095);
and U14584 (N_14584,N_14039,N_13912);
and U14585 (N_14585,N_14102,N_13886);
and U14586 (N_14586,N_13814,N_13981);
or U14587 (N_14587,N_13909,N_14290);
and U14588 (N_14588,N_13753,N_14315);
or U14589 (N_14589,N_13797,N_14197);
nand U14590 (N_14590,N_13818,N_14055);
or U14591 (N_14591,N_14132,N_13835);
or U14592 (N_14592,N_14134,N_14047);
nand U14593 (N_14593,N_14327,N_14255);
and U14594 (N_14594,N_13806,N_14309);
and U14595 (N_14595,N_14208,N_14036);
nor U14596 (N_14596,N_14349,N_14070);
nand U14597 (N_14597,N_14122,N_14150);
nor U14598 (N_14598,N_13757,N_13781);
and U14599 (N_14599,N_13799,N_14191);
and U14600 (N_14600,N_13862,N_13813);
or U14601 (N_14601,N_14343,N_14329);
and U14602 (N_14602,N_14114,N_13874);
or U14603 (N_14603,N_14161,N_13817);
nand U14604 (N_14604,N_14065,N_14027);
nand U14605 (N_14605,N_13894,N_14226);
nor U14606 (N_14606,N_13967,N_14214);
nor U14607 (N_14607,N_14348,N_13888);
or U14608 (N_14608,N_13868,N_14287);
and U14609 (N_14609,N_14341,N_14235);
and U14610 (N_14610,N_14213,N_14014);
xnor U14611 (N_14611,N_14313,N_14176);
nor U14612 (N_14612,N_14043,N_14217);
or U14613 (N_14613,N_14361,N_14322);
and U14614 (N_14614,N_14233,N_14283);
or U14615 (N_14615,N_14155,N_14328);
and U14616 (N_14616,N_14089,N_13858);
nand U14617 (N_14617,N_13764,N_13922);
and U14618 (N_14618,N_14325,N_14128);
or U14619 (N_14619,N_13859,N_13943);
nand U14620 (N_14620,N_13750,N_14093);
xnor U14621 (N_14621,N_14256,N_14356);
and U14622 (N_14622,N_13986,N_14002);
and U14623 (N_14623,N_13788,N_13890);
nand U14624 (N_14624,N_13978,N_14286);
or U14625 (N_14625,N_14326,N_14127);
nor U14626 (N_14626,N_14357,N_14021);
and U14627 (N_14627,N_14183,N_14171);
xnor U14628 (N_14628,N_13949,N_13920);
and U14629 (N_14629,N_13929,N_13752);
nor U14630 (N_14630,N_14199,N_14259);
nor U14631 (N_14631,N_14294,N_14225);
xor U14632 (N_14632,N_14314,N_14001);
nor U14633 (N_14633,N_13773,N_13938);
nand U14634 (N_14634,N_14135,N_14274);
or U14635 (N_14635,N_13976,N_13857);
nor U14636 (N_14636,N_14148,N_14346);
and U14637 (N_14637,N_14158,N_13913);
nand U14638 (N_14638,N_14145,N_14268);
or U14639 (N_14639,N_13872,N_14258);
or U14640 (N_14640,N_14372,N_13794);
nand U14641 (N_14641,N_14091,N_14293);
nor U14642 (N_14642,N_14109,N_13947);
nor U14643 (N_14643,N_14019,N_13826);
nand U14644 (N_14644,N_14181,N_14168);
and U14645 (N_14645,N_13766,N_14025);
nor U14646 (N_14646,N_14118,N_13861);
nand U14647 (N_14647,N_13809,N_13988);
nand U14648 (N_14648,N_14013,N_13751);
nand U14649 (N_14649,N_14133,N_14153);
and U14650 (N_14650,N_13848,N_13980);
or U14651 (N_14651,N_13940,N_13942);
or U14652 (N_14652,N_14184,N_13995);
nor U14653 (N_14653,N_14125,N_13776);
nand U14654 (N_14654,N_14267,N_13915);
and U14655 (N_14655,N_14219,N_14051);
and U14656 (N_14656,N_14107,N_14232);
xnor U14657 (N_14657,N_14198,N_13925);
or U14658 (N_14658,N_14253,N_14337);
nand U14659 (N_14659,N_14182,N_13838);
xnor U14660 (N_14660,N_14016,N_14057);
and U14661 (N_14661,N_14370,N_14022);
or U14662 (N_14662,N_13877,N_14121);
nor U14663 (N_14663,N_13946,N_13833);
nand U14664 (N_14664,N_13905,N_14092);
nand U14665 (N_14665,N_14071,N_14015);
nand U14666 (N_14666,N_14350,N_14023);
or U14667 (N_14667,N_14123,N_14156);
and U14668 (N_14668,N_13962,N_13954);
xor U14669 (N_14669,N_14228,N_14053);
nand U14670 (N_14670,N_13993,N_14236);
nand U14671 (N_14671,N_13907,N_13959);
nor U14672 (N_14672,N_14353,N_14048);
nand U14673 (N_14673,N_13917,N_14151);
nor U14674 (N_14674,N_14239,N_13825);
and U14675 (N_14675,N_14104,N_14117);
xor U14676 (N_14676,N_14033,N_14088);
xnor U14677 (N_14677,N_14142,N_14272);
and U14678 (N_14678,N_14229,N_14108);
nand U14679 (N_14679,N_14223,N_14035);
nand U14680 (N_14680,N_14159,N_14061);
nor U14681 (N_14681,N_14068,N_13812);
or U14682 (N_14682,N_13893,N_13815);
and U14683 (N_14683,N_13785,N_13950);
nor U14684 (N_14684,N_14018,N_14262);
nand U14685 (N_14685,N_14248,N_13887);
or U14686 (N_14686,N_13820,N_14067);
and U14687 (N_14687,N_13816,N_13754);
nand U14688 (N_14688,N_14097,N_14065);
and U14689 (N_14689,N_13913,N_13815);
or U14690 (N_14690,N_13799,N_14264);
nor U14691 (N_14691,N_13820,N_14114);
xnor U14692 (N_14692,N_14266,N_13885);
or U14693 (N_14693,N_13990,N_14372);
nand U14694 (N_14694,N_14323,N_13786);
nand U14695 (N_14695,N_14060,N_14141);
xnor U14696 (N_14696,N_14316,N_14165);
nand U14697 (N_14697,N_13880,N_13815);
or U14698 (N_14698,N_13881,N_13856);
nor U14699 (N_14699,N_13841,N_14316);
or U14700 (N_14700,N_14099,N_13963);
or U14701 (N_14701,N_14093,N_13800);
or U14702 (N_14702,N_13782,N_13959);
or U14703 (N_14703,N_14287,N_13911);
nand U14704 (N_14704,N_13954,N_13760);
and U14705 (N_14705,N_14132,N_13791);
nor U14706 (N_14706,N_14010,N_14102);
or U14707 (N_14707,N_14005,N_14279);
nand U14708 (N_14708,N_14009,N_14344);
and U14709 (N_14709,N_14125,N_14070);
nand U14710 (N_14710,N_14249,N_13874);
nor U14711 (N_14711,N_13954,N_13942);
nor U14712 (N_14712,N_14262,N_14328);
nor U14713 (N_14713,N_14178,N_14010);
or U14714 (N_14714,N_14121,N_14091);
nor U14715 (N_14715,N_14363,N_14264);
nor U14716 (N_14716,N_13789,N_13855);
or U14717 (N_14717,N_14142,N_14091);
nand U14718 (N_14718,N_13783,N_14306);
or U14719 (N_14719,N_13872,N_14277);
nand U14720 (N_14720,N_14370,N_14084);
and U14721 (N_14721,N_13785,N_14240);
and U14722 (N_14722,N_14075,N_14070);
and U14723 (N_14723,N_13804,N_14365);
xnor U14724 (N_14724,N_14022,N_14023);
nor U14725 (N_14725,N_14211,N_14286);
or U14726 (N_14726,N_13787,N_14099);
nand U14727 (N_14727,N_14025,N_14240);
nor U14728 (N_14728,N_14029,N_14322);
nor U14729 (N_14729,N_14188,N_13822);
nand U14730 (N_14730,N_14371,N_14200);
nand U14731 (N_14731,N_14021,N_13783);
nor U14732 (N_14732,N_14169,N_14309);
nand U14733 (N_14733,N_14274,N_14193);
or U14734 (N_14734,N_14352,N_13915);
or U14735 (N_14735,N_14321,N_14048);
or U14736 (N_14736,N_14153,N_14332);
and U14737 (N_14737,N_14183,N_13858);
or U14738 (N_14738,N_13945,N_14105);
nor U14739 (N_14739,N_14338,N_14265);
or U14740 (N_14740,N_13875,N_14080);
nor U14741 (N_14741,N_14009,N_14227);
or U14742 (N_14742,N_13769,N_13878);
or U14743 (N_14743,N_14114,N_13998);
nand U14744 (N_14744,N_13807,N_14358);
and U14745 (N_14745,N_13902,N_13770);
nor U14746 (N_14746,N_13806,N_13893);
or U14747 (N_14747,N_13868,N_14033);
nand U14748 (N_14748,N_14076,N_14042);
xor U14749 (N_14749,N_14210,N_14014);
and U14750 (N_14750,N_14192,N_13826);
nand U14751 (N_14751,N_13750,N_13874);
or U14752 (N_14752,N_13906,N_14059);
or U14753 (N_14753,N_14299,N_14224);
nand U14754 (N_14754,N_13786,N_14015);
and U14755 (N_14755,N_14264,N_14328);
nand U14756 (N_14756,N_14282,N_13827);
and U14757 (N_14757,N_14274,N_14323);
nand U14758 (N_14758,N_14167,N_13976);
nand U14759 (N_14759,N_14173,N_14116);
or U14760 (N_14760,N_13836,N_13831);
and U14761 (N_14761,N_13891,N_13884);
and U14762 (N_14762,N_14350,N_14091);
nor U14763 (N_14763,N_13944,N_13774);
and U14764 (N_14764,N_14132,N_14327);
and U14765 (N_14765,N_13953,N_13982);
or U14766 (N_14766,N_13984,N_14199);
nor U14767 (N_14767,N_14259,N_13930);
or U14768 (N_14768,N_14063,N_14234);
or U14769 (N_14769,N_13912,N_14356);
nand U14770 (N_14770,N_14274,N_14260);
xor U14771 (N_14771,N_14235,N_13805);
and U14772 (N_14772,N_14144,N_14328);
or U14773 (N_14773,N_14182,N_13872);
and U14774 (N_14774,N_13896,N_13980);
nor U14775 (N_14775,N_14296,N_13840);
nor U14776 (N_14776,N_14027,N_14208);
nand U14777 (N_14777,N_14011,N_13931);
or U14778 (N_14778,N_13979,N_14256);
nand U14779 (N_14779,N_14219,N_13821);
nand U14780 (N_14780,N_13939,N_13847);
nor U14781 (N_14781,N_14229,N_14073);
and U14782 (N_14782,N_14029,N_14024);
nor U14783 (N_14783,N_13960,N_14242);
nand U14784 (N_14784,N_14304,N_13804);
and U14785 (N_14785,N_13841,N_13769);
or U14786 (N_14786,N_14236,N_13757);
nand U14787 (N_14787,N_13805,N_13840);
nand U14788 (N_14788,N_14335,N_13772);
nand U14789 (N_14789,N_14211,N_14089);
and U14790 (N_14790,N_14321,N_14340);
and U14791 (N_14791,N_14124,N_14178);
nand U14792 (N_14792,N_14271,N_13944);
nor U14793 (N_14793,N_14052,N_13891);
nand U14794 (N_14794,N_13812,N_14218);
nor U14795 (N_14795,N_13848,N_13933);
nor U14796 (N_14796,N_13973,N_14217);
nand U14797 (N_14797,N_14216,N_14076);
or U14798 (N_14798,N_13919,N_14111);
nand U14799 (N_14799,N_14200,N_13764);
and U14800 (N_14800,N_14340,N_13971);
and U14801 (N_14801,N_14044,N_14337);
nor U14802 (N_14802,N_14035,N_13825);
or U14803 (N_14803,N_13849,N_14355);
nand U14804 (N_14804,N_13754,N_14043);
nor U14805 (N_14805,N_13812,N_14026);
nand U14806 (N_14806,N_14143,N_14071);
nand U14807 (N_14807,N_14341,N_13890);
and U14808 (N_14808,N_13928,N_14159);
nand U14809 (N_14809,N_13871,N_13954);
nand U14810 (N_14810,N_13971,N_14368);
and U14811 (N_14811,N_13805,N_14057);
or U14812 (N_14812,N_14136,N_14123);
nand U14813 (N_14813,N_14251,N_14168);
and U14814 (N_14814,N_14138,N_13849);
nand U14815 (N_14815,N_13881,N_14205);
nand U14816 (N_14816,N_13936,N_13750);
and U14817 (N_14817,N_13931,N_13956);
or U14818 (N_14818,N_14118,N_13958);
or U14819 (N_14819,N_14084,N_13847);
nand U14820 (N_14820,N_14329,N_14148);
or U14821 (N_14821,N_14364,N_13988);
nor U14822 (N_14822,N_13934,N_14115);
xor U14823 (N_14823,N_13832,N_13941);
and U14824 (N_14824,N_14113,N_14045);
or U14825 (N_14825,N_14268,N_13833);
or U14826 (N_14826,N_14341,N_13814);
xnor U14827 (N_14827,N_14191,N_14008);
nor U14828 (N_14828,N_14119,N_14266);
xnor U14829 (N_14829,N_14367,N_13841);
nor U14830 (N_14830,N_14180,N_14012);
and U14831 (N_14831,N_14250,N_13968);
nor U14832 (N_14832,N_13829,N_13957);
or U14833 (N_14833,N_13750,N_13908);
xor U14834 (N_14834,N_14225,N_14027);
nor U14835 (N_14835,N_13999,N_14208);
xor U14836 (N_14836,N_13900,N_14096);
nand U14837 (N_14837,N_13963,N_14051);
or U14838 (N_14838,N_14373,N_14152);
and U14839 (N_14839,N_14018,N_13964);
nand U14840 (N_14840,N_14253,N_14119);
xnor U14841 (N_14841,N_13944,N_14013);
xnor U14842 (N_14842,N_14015,N_13813);
and U14843 (N_14843,N_13811,N_14044);
nor U14844 (N_14844,N_13974,N_13976);
nand U14845 (N_14845,N_14143,N_14144);
nand U14846 (N_14846,N_13840,N_14270);
and U14847 (N_14847,N_13876,N_14264);
and U14848 (N_14848,N_13813,N_13997);
nand U14849 (N_14849,N_14287,N_14272);
nand U14850 (N_14850,N_13894,N_14041);
and U14851 (N_14851,N_14237,N_14151);
xnor U14852 (N_14852,N_14374,N_14150);
nor U14853 (N_14853,N_14163,N_14155);
and U14854 (N_14854,N_13907,N_13855);
nand U14855 (N_14855,N_14097,N_13902);
nor U14856 (N_14856,N_14241,N_14344);
or U14857 (N_14857,N_14181,N_14238);
and U14858 (N_14858,N_14220,N_13805);
and U14859 (N_14859,N_14257,N_14286);
nor U14860 (N_14860,N_14083,N_13984);
nor U14861 (N_14861,N_14028,N_14013);
xnor U14862 (N_14862,N_14277,N_13903);
nand U14863 (N_14863,N_14158,N_14371);
nor U14864 (N_14864,N_14097,N_14281);
xnor U14865 (N_14865,N_14035,N_13810);
or U14866 (N_14866,N_14197,N_13841);
nor U14867 (N_14867,N_14233,N_13792);
and U14868 (N_14868,N_14009,N_13962);
nand U14869 (N_14869,N_14297,N_14081);
and U14870 (N_14870,N_14061,N_13813);
or U14871 (N_14871,N_13843,N_14284);
and U14872 (N_14872,N_14051,N_14112);
and U14873 (N_14873,N_13896,N_14183);
nand U14874 (N_14874,N_14119,N_14209);
or U14875 (N_14875,N_13913,N_14118);
or U14876 (N_14876,N_14165,N_14056);
xnor U14877 (N_14877,N_14009,N_13960);
nor U14878 (N_14878,N_14330,N_13990);
or U14879 (N_14879,N_13868,N_13853);
and U14880 (N_14880,N_13803,N_13798);
or U14881 (N_14881,N_14057,N_13981);
nor U14882 (N_14882,N_13847,N_14106);
and U14883 (N_14883,N_13974,N_13752);
nand U14884 (N_14884,N_13847,N_14115);
nand U14885 (N_14885,N_13876,N_14333);
and U14886 (N_14886,N_13950,N_13786);
or U14887 (N_14887,N_14098,N_14334);
and U14888 (N_14888,N_13968,N_14199);
or U14889 (N_14889,N_14325,N_13812);
or U14890 (N_14890,N_14369,N_13971);
and U14891 (N_14891,N_13988,N_13879);
nand U14892 (N_14892,N_13936,N_14013);
and U14893 (N_14893,N_14084,N_14303);
or U14894 (N_14894,N_14137,N_14246);
and U14895 (N_14895,N_14253,N_14313);
or U14896 (N_14896,N_14053,N_13990);
nand U14897 (N_14897,N_13786,N_14176);
nor U14898 (N_14898,N_14128,N_13895);
and U14899 (N_14899,N_13872,N_13785);
or U14900 (N_14900,N_14070,N_13822);
and U14901 (N_14901,N_14342,N_14267);
nand U14902 (N_14902,N_14116,N_14243);
nand U14903 (N_14903,N_13786,N_13905);
and U14904 (N_14904,N_13764,N_14199);
or U14905 (N_14905,N_13757,N_14292);
or U14906 (N_14906,N_14002,N_14095);
nand U14907 (N_14907,N_14194,N_13888);
and U14908 (N_14908,N_14016,N_14026);
nor U14909 (N_14909,N_13832,N_13826);
or U14910 (N_14910,N_14282,N_14253);
or U14911 (N_14911,N_14169,N_14256);
nand U14912 (N_14912,N_14018,N_14350);
or U14913 (N_14913,N_14293,N_14296);
and U14914 (N_14914,N_14089,N_14218);
nor U14915 (N_14915,N_14224,N_13771);
nand U14916 (N_14916,N_13864,N_14160);
nand U14917 (N_14917,N_14200,N_13854);
or U14918 (N_14918,N_14245,N_13886);
nor U14919 (N_14919,N_13861,N_14163);
nor U14920 (N_14920,N_14215,N_14227);
or U14921 (N_14921,N_14204,N_14096);
nand U14922 (N_14922,N_13783,N_14049);
nand U14923 (N_14923,N_13905,N_14228);
or U14924 (N_14924,N_14178,N_14363);
or U14925 (N_14925,N_14181,N_13797);
and U14926 (N_14926,N_13882,N_14336);
nand U14927 (N_14927,N_13962,N_14175);
nor U14928 (N_14928,N_13787,N_13835);
nor U14929 (N_14929,N_14015,N_14023);
or U14930 (N_14930,N_14016,N_14070);
and U14931 (N_14931,N_13759,N_14086);
or U14932 (N_14932,N_14285,N_14011);
and U14933 (N_14933,N_14338,N_14192);
nor U14934 (N_14934,N_13869,N_13983);
and U14935 (N_14935,N_13849,N_14373);
nor U14936 (N_14936,N_14230,N_13864);
nor U14937 (N_14937,N_13843,N_13761);
nand U14938 (N_14938,N_13952,N_13823);
nor U14939 (N_14939,N_14008,N_14040);
and U14940 (N_14940,N_14282,N_14000);
and U14941 (N_14941,N_13934,N_14001);
nand U14942 (N_14942,N_14070,N_14292);
or U14943 (N_14943,N_13754,N_13896);
or U14944 (N_14944,N_14162,N_14265);
xor U14945 (N_14945,N_13774,N_13976);
and U14946 (N_14946,N_14373,N_13970);
or U14947 (N_14947,N_13981,N_14085);
nor U14948 (N_14948,N_14049,N_14077);
xnor U14949 (N_14949,N_13879,N_13758);
and U14950 (N_14950,N_13865,N_13982);
or U14951 (N_14951,N_13780,N_14162);
and U14952 (N_14952,N_14136,N_13826);
nor U14953 (N_14953,N_14078,N_13784);
and U14954 (N_14954,N_14335,N_14296);
xor U14955 (N_14955,N_14254,N_14233);
and U14956 (N_14956,N_14074,N_14351);
or U14957 (N_14957,N_13903,N_14248);
or U14958 (N_14958,N_13804,N_13977);
or U14959 (N_14959,N_14217,N_13860);
and U14960 (N_14960,N_13952,N_13771);
nand U14961 (N_14961,N_13958,N_13884);
nand U14962 (N_14962,N_13895,N_14209);
and U14963 (N_14963,N_14115,N_14068);
and U14964 (N_14964,N_14127,N_14322);
and U14965 (N_14965,N_14301,N_13819);
or U14966 (N_14966,N_14354,N_14285);
nand U14967 (N_14967,N_14173,N_13873);
nor U14968 (N_14968,N_14136,N_14279);
xor U14969 (N_14969,N_14125,N_13866);
and U14970 (N_14970,N_13944,N_14177);
and U14971 (N_14971,N_13879,N_13826);
and U14972 (N_14972,N_13973,N_14300);
and U14973 (N_14973,N_14273,N_14026);
or U14974 (N_14974,N_14065,N_14188);
and U14975 (N_14975,N_13935,N_14162);
and U14976 (N_14976,N_13915,N_14223);
and U14977 (N_14977,N_13980,N_13893);
or U14978 (N_14978,N_13897,N_13833);
and U14979 (N_14979,N_14368,N_14202);
or U14980 (N_14980,N_14021,N_13987);
or U14981 (N_14981,N_13869,N_14156);
and U14982 (N_14982,N_13978,N_13903);
or U14983 (N_14983,N_14247,N_13914);
and U14984 (N_14984,N_14199,N_14127);
and U14985 (N_14985,N_13979,N_14097);
nor U14986 (N_14986,N_14197,N_14357);
xor U14987 (N_14987,N_13842,N_13766);
nor U14988 (N_14988,N_13884,N_14068);
or U14989 (N_14989,N_13955,N_13922);
and U14990 (N_14990,N_13835,N_13776);
or U14991 (N_14991,N_14018,N_13866);
nand U14992 (N_14992,N_14241,N_14150);
or U14993 (N_14993,N_13979,N_13921);
or U14994 (N_14994,N_14059,N_13806);
xnor U14995 (N_14995,N_14004,N_14269);
nor U14996 (N_14996,N_13954,N_14194);
nor U14997 (N_14997,N_13897,N_14135);
nor U14998 (N_14998,N_13841,N_14238);
or U14999 (N_14999,N_14095,N_13923);
nor U15000 (N_15000,N_14498,N_14402);
and U15001 (N_15001,N_14787,N_14490);
or U15002 (N_15002,N_14509,N_14837);
nor U15003 (N_15003,N_14992,N_14618);
nand U15004 (N_15004,N_14758,N_14974);
and U15005 (N_15005,N_14803,N_14864);
nand U15006 (N_15006,N_14685,N_14907);
nand U15007 (N_15007,N_14869,N_14957);
and U15008 (N_15008,N_14559,N_14538);
nor U15009 (N_15009,N_14886,N_14772);
or U15010 (N_15010,N_14451,N_14844);
nor U15011 (N_15011,N_14825,N_14578);
and U15012 (N_15012,N_14983,N_14676);
nor U15013 (N_15013,N_14699,N_14583);
or U15014 (N_15014,N_14857,N_14807);
nor U15015 (N_15015,N_14884,N_14475);
and U15016 (N_15016,N_14880,N_14591);
nor U15017 (N_15017,N_14963,N_14673);
nor U15018 (N_15018,N_14980,N_14926);
and U15019 (N_15019,N_14437,N_14505);
nand U15020 (N_15020,N_14532,N_14744);
nand U15021 (N_15021,N_14416,N_14650);
xnor U15022 (N_15022,N_14883,N_14707);
nor U15023 (N_15023,N_14608,N_14683);
xor U15024 (N_15024,N_14541,N_14670);
xor U15025 (N_15025,N_14860,N_14562);
xor U15026 (N_15026,N_14548,N_14750);
or U15027 (N_15027,N_14652,N_14634);
xnor U15028 (N_15028,N_14503,N_14477);
xor U15029 (N_15029,N_14898,N_14522);
nor U15030 (N_15030,N_14692,N_14735);
or U15031 (N_15031,N_14891,N_14823);
and U15032 (N_15032,N_14977,N_14757);
xor U15033 (N_15033,N_14688,N_14812);
xnor U15034 (N_15034,N_14700,N_14798);
xnor U15035 (N_15035,N_14593,N_14553);
nor U15036 (N_15036,N_14403,N_14910);
or U15037 (N_15037,N_14877,N_14656);
nand U15038 (N_15038,N_14472,N_14784);
or U15039 (N_15039,N_14419,N_14939);
and U15040 (N_15040,N_14946,N_14818);
or U15041 (N_15041,N_14681,N_14494);
or U15042 (N_15042,N_14894,N_14870);
nor U15043 (N_15043,N_14485,N_14441);
or U15044 (N_15044,N_14762,N_14956);
nand U15045 (N_15045,N_14783,N_14835);
nand U15046 (N_15046,N_14727,N_14380);
nand U15047 (N_15047,N_14628,N_14631);
and U15048 (N_15048,N_14840,N_14551);
nand U15049 (N_15049,N_14533,N_14520);
nand U15050 (N_15050,N_14516,N_14859);
nor U15051 (N_15051,N_14941,N_14932);
nand U15052 (N_15052,N_14693,N_14420);
nand U15053 (N_15053,N_14666,N_14464);
and U15054 (N_15054,N_14550,N_14756);
nor U15055 (N_15055,N_14904,N_14597);
or U15056 (N_15056,N_14760,N_14721);
and U15057 (N_15057,N_14995,N_14810);
or U15058 (N_15058,N_14947,N_14426);
nand U15059 (N_15059,N_14718,N_14919);
or U15060 (N_15060,N_14920,N_14937);
nor U15061 (N_15061,N_14796,N_14465);
nor U15062 (N_15062,N_14715,N_14610);
or U15063 (N_15063,N_14741,N_14852);
xor U15064 (N_15064,N_14714,N_14861);
or U15065 (N_15065,N_14515,N_14854);
nor U15066 (N_15066,N_14511,N_14876);
xnor U15067 (N_15067,N_14710,N_14701);
and U15068 (N_15068,N_14731,N_14950);
nor U15069 (N_15069,N_14755,N_14887);
nor U15070 (N_15070,N_14739,N_14406);
or U15071 (N_15071,N_14577,N_14815);
nand U15072 (N_15072,N_14708,N_14620);
and U15073 (N_15073,N_14568,N_14691);
or U15074 (N_15074,N_14732,N_14982);
and U15075 (N_15075,N_14563,N_14952);
or U15076 (N_15076,N_14381,N_14421);
and U15077 (N_15077,N_14927,N_14418);
or U15078 (N_15078,N_14549,N_14613);
nand U15079 (N_15079,N_14508,N_14863);
and U15080 (N_15080,N_14543,N_14930);
nand U15081 (N_15081,N_14761,N_14448);
and U15082 (N_15082,N_14990,N_14445);
and U15083 (N_15083,N_14399,N_14745);
nand U15084 (N_15084,N_14817,N_14734);
and U15085 (N_15085,N_14949,N_14822);
nand U15086 (N_15086,N_14793,N_14425);
or U15087 (N_15087,N_14879,N_14856);
or U15088 (N_15088,N_14836,N_14914);
xnor U15089 (N_15089,N_14985,N_14853);
nand U15090 (N_15090,N_14888,N_14737);
nand U15091 (N_15091,N_14530,N_14604);
xnor U15092 (N_15092,N_14609,N_14924);
nor U15093 (N_15093,N_14386,N_14393);
xnor U15094 (N_15094,N_14599,N_14633);
nor U15095 (N_15095,N_14696,N_14684);
nor U15096 (N_15096,N_14596,N_14991);
nor U15097 (N_15097,N_14637,N_14571);
or U15098 (N_15098,N_14720,N_14875);
nand U15099 (N_15099,N_14482,N_14849);
or U15100 (N_15100,N_14736,N_14642);
nand U15101 (N_15101,N_14502,N_14753);
nand U15102 (N_15102,N_14407,N_14943);
nand U15103 (N_15103,N_14558,N_14646);
nand U15104 (N_15104,N_14722,N_14889);
xnor U15105 (N_15105,N_14975,N_14858);
nor U15106 (N_15106,N_14627,N_14713);
and U15107 (N_15107,N_14899,N_14453);
nor U15108 (N_15108,N_14662,N_14851);
or U15109 (N_15109,N_14717,N_14581);
or U15110 (N_15110,N_14987,N_14589);
xor U15111 (N_15111,N_14679,N_14751);
nand U15112 (N_15112,N_14424,N_14590);
and U15113 (N_15113,N_14725,N_14917);
or U15114 (N_15114,N_14377,N_14706);
nor U15115 (N_15115,N_14774,N_14617);
or U15116 (N_15116,N_14436,N_14458);
or U15117 (N_15117,N_14896,N_14481);
and U15118 (N_15118,N_14624,N_14671);
and U15119 (N_15119,N_14978,N_14566);
nor U15120 (N_15120,N_14561,N_14697);
nand U15121 (N_15121,N_14848,N_14728);
xnor U15122 (N_15122,N_14970,N_14915);
nand U15123 (N_15123,N_14964,N_14387);
nor U15124 (N_15124,N_14669,N_14874);
nor U15125 (N_15125,N_14430,N_14546);
or U15126 (N_15126,N_14459,N_14576);
xor U15127 (N_15127,N_14592,N_14933);
or U15128 (N_15128,N_14612,N_14973);
and U15129 (N_15129,N_14994,N_14544);
nor U15130 (N_15130,N_14616,N_14658);
nor U15131 (N_15131,N_14567,N_14655);
or U15132 (N_15132,N_14890,N_14529);
and U15133 (N_15133,N_14800,N_14828);
nor U15134 (N_15134,N_14906,N_14623);
nor U15135 (N_15135,N_14893,N_14855);
nor U15136 (N_15136,N_14841,N_14411);
and U15137 (N_15137,N_14659,N_14555);
nand U15138 (N_15138,N_14526,N_14582);
or U15139 (N_15139,N_14928,N_14640);
nor U15140 (N_15140,N_14375,N_14382);
or U15141 (N_15141,N_14663,N_14376);
xnor U15142 (N_15142,N_14677,N_14452);
or U15143 (N_15143,N_14913,N_14469);
and U15144 (N_15144,N_14766,N_14535);
or U15145 (N_15145,N_14958,N_14759);
and U15146 (N_15146,N_14971,N_14776);
or U15147 (N_15147,N_14791,N_14686);
nor U15148 (N_15148,N_14705,N_14556);
nand U15149 (N_15149,N_14903,N_14622);
nor U15150 (N_15150,N_14711,N_14528);
nor U15151 (N_15151,N_14976,N_14940);
or U15152 (N_15152,N_14444,N_14545);
and U15153 (N_15153,N_14636,N_14769);
nand U15154 (N_15154,N_14394,N_14443);
xnor U15155 (N_15155,N_14629,N_14385);
or U15156 (N_15156,N_14547,N_14694);
nor U15157 (N_15157,N_14584,N_14554);
nor U15158 (N_15158,N_14476,N_14461);
nor U15159 (N_15159,N_14743,N_14492);
nand U15160 (N_15160,N_14569,N_14999);
or U15161 (N_15161,N_14621,N_14954);
nand U15162 (N_15162,N_14905,N_14434);
xor U15163 (N_15163,N_14519,N_14586);
and U15164 (N_15164,N_14647,N_14724);
xnor U15165 (N_15165,N_14965,N_14517);
nor U15166 (N_15166,N_14850,N_14872);
or U15167 (N_15167,N_14979,N_14829);
nor U15168 (N_15168,N_14495,N_14786);
and U15169 (N_15169,N_14768,N_14531);
or U15170 (N_15170,N_14955,N_14908);
or U15171 (N_15171,N_14439,N_14902);
and U15172 (N_15172,N_14948,N_14487);
and U15173 (N_15173,N_14767,N_14660);
or U15174 (N_15174,N_14748,N_14493);
or U15175 (N_15175,N_14468,N_14514);
xnor U15176 (N_15176,N_14625,N_14912);
or U15177 (N_15177,N_14518,N_14614);
nor U15178 (N_15178,N_14993,N_14833);
xor U15179 (N_15179,N_14805,N_14579);
and U15180 (N_15180,N_14703,N_14478);
and U15181 (N_15181,N_14474,N_14649);
and U15182 (N_15182,N_14824,N_14934);
or U15183 (N_15183,N_14820,N_14830);
or U15184 (N_15184,N_14540,N_14704);
and U15185 (N_15185,N_14921,N_14777);
nand U15186 (N_15186,N_14638,N_14813);
nor U15187 (N_15187,N_14395,N_14689);
or U15188 (N_15188,N_14542,N_14998);
and U15189 (N_15189,N_14454,N_14587);
or U15190 (N_15190,N_14456,N_14537);
and U15191 (N_15191,N_14429,N_14945);
and U15192 (N_15192,N_14497,N_14414);
or U15193 (N_15193,N_14484,N_14674);
or U15194 (N_15194,N_14878,N_14698);
and U15195 (N_15195,N_14885,N_14962);
nor U15196 (N_15196,N_14450,N_14966);
and U15197 (N_15197,N_14968,N_14738);
or U15198 (N_15198,N_14440,N_14400);
nor U15199 (N_15199,N_14862,N_14832);
nor U15200 (N_15200,N_14644,N_14560);
and U15201 (N_15201,N_14672,N_14521);
and U15202 (N_15202,N_14778,N_14695);
or U15203 (N_15203,N_14570,N_14539);
nor U15204 (N_15204,N_14630,N_14846);
xor U15205 (N_15205,N_14938,N_14588);
and U15206 (N_15206,N_14463,N_14389);
nand U15207 (N_15207,N_14496,N_14447);
nor U15208 (N_15208,N_14808,N_14657);
and U15209 (N_15209,N_14398,N_14981);
nand U15210 (N_15210,N_14873,N_14733);
nand U15211 (N_15211,N_14392,N_14564);
xnor U15212 (N_15212,N_14749,N_14557);
nand U15213 (N_15213,N_14504,N_14600);
and U15214 (N_15214,N_14536,N_14967);
and U15215 (N_15215,N_14687,N_14422);
or U15216 (N_15216,N_14635,N_14712);
and U15217 (N_15217,N_14431,N_14388);
or U15218 (N_15218,N_14782,N_14961);
and U15219 (N_15219,N_14845,N_14918);
or U15220 (N_15220,N_14802,N_14811);
xnor U15221 (N_15221,N_14653,N_14868);
xnor U15222 (N_15222,N_14740,N_14794);
nand U15223 (N_15223,N_14892,N_14729);
or U15224 (N_15224,N_14648,N_14479);
or U15225 (N_15225,N_14882,N_14931);
nand U15226 (N_15226,N_14726,N_14922);
or U15227 (N_15227,N_14865,N_14702);
and U15228 (N_15228,N_14916,N_14489);
and U15229 (N_15229,N_14816,N_14988);
nor U15230 (N_15230,N_14680,N_14598);
and U15231 (N_15231,N_14483,N_14942);
nor U15232 (N_15232,N_14754,N_14801);
xnor U15233 (N_15233,N_14821,N_14763);
and U15234 (N_15234,N_14747,N_14843);
and U15235 (N_15235,N_14442,N_14661);
or U15236 (N_15236,N_14771,N_14765);
xor U15237 (N_15237,N_14510,N_14410);
or U15238 (N_15238,N_14675,N_14523);
xor U15239 (N_15239,N_14378,N_14969);
nand U15240 (N_15240,N_14491,N_14925);
xor U15241 (N_15241,N_14460,N_14455);
nor U15242 (N_15242,N_14607,N_14651);
or U15243 (N_15243,N_14831,N_14842);
and U15244 (N_15244,N_14997,N_14895);
or U15245 (N_15245,N_14433,N_14795);
nor U15246 (N_15246,N_14716,N_14960);
and U15247 (N_15247,N_14742,N_14524);
and U15248 (N_15248,N_14838,N_14923);
xnor U15249 (N_15249,N_14789,N_14580);
or U15250 (N_15250,N_14471,N_14639);
nor U15251 (N_15251,N_14413,N_14814);
or U15252 (N_15252,N_14396,N_14682);
nand U15253 (N_15253,N_14909,N_14435);
xnor U15254 (N_15254,N_14438,N_14575);
nor U15255 (N_15255,N_14601,N_14780);
nor U15256 (N_15256,N_14500,N_14900);
or U15257 (N_15257,N_14984,N_14645);
and U15258 (N_15258,N_14897,N_14866);
or U15259 (N_15259,N_14664,N_14573);
or U15260 (N_15260,N_14781,N_14643);
and U15261 (N_15261,N_14797,N_14488);
nor U15262 (N_15262,N_14462,N_14901);
xor U15263 (N_15263,N_14507,N_14391);
nand U15264 (N_15264,N_14944,N_14972);
nand U15265 (N_15265,N_14552,N_14480);
and U15266 (N_15266,N_14951,N_14632);
or U15267 (N_15267,N_14412,N_14626);
nand U15268 (N_15268,N_14585,N_14752);
nor U15269 (N_15269,N_14779,N_14595);
and U15270 (N_15270,N_14486,N_14594);
nor U15271 (N_15271,N_14408,N_14428);
nor U15272 (N_15272,N_14723,N_14574);
and U15273 (N_15273,N_14678,N_14506);
nor U15274 (N_15274,N_14788,N_14775);
or U15275 (N_15275,N_14525,N_14953);
and U15276 (N_15276,N_14415,N_14665);
or U15277 (N_15277,N_14404,N_14989);
and U15278 (N_15278,N_14534,N_14565);
nor U15279 (N_15279,N_14809,N_14605);
or U15280 (N_15280,N_14512,N_14615);
xnor U15281 (N_15281,N_14513,N_14603);
and U15282 (N_15282,N_14467,N_14826);
and U15283 (N_15283,N_14770,N_14785);
or U15284 (N_15284,N_14446,N_14709);
nand U15285 (N_15285,N_14384,N_14959);
or U15286 (N_15286,N_14936,N_14834);
nor U15287 (N_15287,N_14881,N_14572);
or U15288 (N_15288,N_14690,N_14449);
or U15289 (N_15289,N_14606,N_14827);
xnor U15290 (N_15290,N_14667,N_14929);
nor U15291 (N_15291,N_14804,N_14602);
nand U15292 (N_15292,N_14501,N_14473);
or U15293 (N_15293,N_14867,N_14383);
nand U15294 (N_15294,N_14427,N_14417);
or U15295 (N_15295,N_14466,N_14730);
and U15296 (N_15296,N_14819,N_14871);
or U15297 (N_15297,N_14470,N_14379);
and U15298 (N_15298,N_14764,N_14935);
nor U15299 (N_15299,N_14996,N_14847);
or U15300 (N_15300,N_14499,N_14401);
or U15301 (N_15301,N_14654,N_14619);
or U15302 (N_15302,N_14806,N_14397);
and U15303 (N_15303,N_14799,N_14390);
and U15304 (N_15304,N_14527,N_14911);
and U15305 (N_15305,N_14409,N_14668);
or U15306 (N_15306,N_14405,N_14790);
nor U15307 (N_15307,N_14986,N_14611);
xor U15308 (N_15308,N_14746,N_14719);
nor U15309 (N_15309,N_14641,N_14792);
nor U15310 (N_15310,N_14839,N_14432);
or U15311 (N_15311,N_14773,N_14423);
nor U15312 (N_15312,N_14457,N_14497);
or U15313 (N_15313,N_14427,N_14706);
nor U15314 (N_15314,N_14404,N_14709);
xnor U15315 (N_15315,N_14655,N_14812);
nand U15316 (N_15316,N_14381,N_14547);
and U15317 (N_15317,N_14798,N_14624);
xnor U15318 (N_15318,N_14945,N_14672);
nand U15319 (N_15319,N_14616,N_14656);
xnor U15320 (N_15320,N_14688,N_14724);
or U15321 (N_15321,N_14625,N_14968);
or U15322 (N_15322,N_14717,N_14798);
nand U15323 (N_15323,N_14534,N_14869);
and U15324 (N_15324,N_14579,N_14983);
nand U15325 (N_15325,N_14418,N_14555);
and U15326 (N_15326,N_14697,N_14707);
and U15327 (N_15327,N_14881,N_14846);
nor U15328 (N_15328,N_14664,N_14527);
or U15329 (N_15329,N_14595,N_14386);
and U15330 (N_15330,N_14633,N_14857);
nand U15331 (N_15331,N_14831,N_14395);
xor U15332 (N_15332,N_14767,N_14473);
and U15333 (N_15333,N_14818,N_14517);
and U15334 (N_15334,N_14748,N_14772);
and U15335 (N_15335,N_14663,N_14552);
nand U15336 (N_15336,N_14745,N_14902);
and U15337 (N_15337,N_14708,N_14933);
and U15338 (N_15338,N_14566,N_14679);
and U15339 (N_15339,N_14588,N_14414);
and U15340 (N_15340,N_14906,N_14960);
and U15341 (N_15341,N_14583,N_14707);
nor U15342 (N_15342,N_14941,N_14420);
and U15343 (N_15343,N_14655,N_14423);
nand U15344 (N_15344,N_14859,N_14596);
or U15345 (N_15345,N_14653,N_14610);
nand U15346 (N_15346,N_14900,N_14436);
nor U15347 (N_15347,N_14467,N_14510);
and U15348 (N_15348,N_14494,N_14680);
xor U15349 (N_15349,N_14827,N_14964);
or U15350 (N_15350,N_14587,N_14624);
nand U15351 (N_15351,N_14698,N_14641);
nand U15352 (N_15352,N_14610,N_14890);
nor U15353 (N_15353,N_14562,N_14850);
xor U15354 (N_15354,N_14670,N_14445);
nand U15355 (N_15355,N_14841,N_14679);
and U15356 (N_15356,N_14745,N_14777);
xnor U15357 (N_15357,N_14397,N_14797);
nand U15358 (N_15358,N_14669,N_14711);
or U15359 (N_15359,N_14957,N_14566);
nor U15360 (N_15360,N_14979,N_14476);
nor U15361 (N_15361,N_14759,N_14741);
or U15362 (N_15362,N_14389,N_14559);
or U15363 (N_15363,N_14984,N_14443);
or U15364 (N_15364,N_14628,N_14911);
nor U15365 (N_15365,N_14577,N_14412);
and U15366 (N_15366,N_14787,N_14652);
nor U15367 (N_15367,N_14385,N_14449);
nor U15368 (N_15368,N_14591,N_14619);
and U15369 (N_15369,N_14533,N_14767);
xor U15370 (N_15370,N_14747,N_14444);
nor U15371 (N_15371,N_14767,N_14653);
nand U15372 (N_15372,N_14911,N_14988);
nor U15373 (N_15373,N_14484,N_14418);
and U15374 (N_15374,N_14870,N_14796);
and U15375 (N_15375,N_14484,N_14535);
xor U15376 (N_15376,N_14740,N_14604);
and U15377 (N_15377,N_14401,N_14820);
nor U15378 (N_15378,N_14849,N_14477);
nand U15379 (N_15379,N_14557,N_14809);
and U15380 (N_15380,N_14470,N_14671);
and U15381 (N_15381,N_14448,N_14474);
or U15382 (N_15382,N_14557,N_14968);
nor U15383 (N_15383,N_14543,N_14489);
nand U15384 (N_15384,N_14410,N_14945);
or U15385 (N_15385,N_14876,N_14776);
nor U15386 (N_15386,N_14919,N_14514);
nor U15387 (N_15387,N_14701,N_14675);
nor U15388 (N_15388,N_14680,N_14686);
or U15389 (N_15389,N_14502,N_14420);
nor U15390 (N_15390,N_14591,N_14636);
nor U15391 (N_15391,N_14627,N_14646);
and U15392 (N_15392,N_14810,N_14624);
xnor U15393 (N_15393,N_14418,N_14929);
xnor U15394 (N_15394,N_14747,N_14637);
xor U15395 (N_15395,N_14859,N_14384);
and U15396 (N_15396,N_14503,N_14731);
nor U15397 (N_15397,N_14928,N_14634);
nand U15398 (N_15398,N_14927,N_14883);
nor U15399 (N_15399,N_14877,N_14469);
and U15400 (N_15400,N_14425,N_14807);
or U15401 (N_15401,N_14558,N_14427);
and U15402 (N_15402,N_14930,N_14864);
nor U15403 (N_15403,N_14472,N_14629);
and U15404 (N_15404,N_14743,N_14456);
or U15405 (N_15405,N_14695,N_14559);
xor U15406 (N_15406,N_14614,N_14774);
or U15407 (N_15407,N_14778,N_14656);
and U15408 (N_15408,N_14865,N_14560);
and U15409 (N_15409,N_14956,N_14754);
and U15410 (N_15410,N_14408,N_14520);
nor U15411 (N_15411,N_14389,N_14629);
nor U15412 (N_15412,N_14549,N_14800);
nor U15413 (N_15413,N_14400,N_14964);
and U15414 (N_15414,N_14778,N_14798);
nor U15415 (N_15415,N_14426,N_14925);
or U15416 (N_15416,N_14820,N_14520);
nor U15417 (N_15417,N_14954,N_14806);
or U15418 (N_15418,N_14859,N_14754);
xnor U15419 (N_15419,N_14750,N_14518);
nor U15420 (N_15420,N_14928,N_14725);
and U15421 (N_15421,N_14984,N_14902);
or U15422 (N_15422,N_14715,N_14697);
and U15423 (N_15423,N_14833,N_14567);
nand U15424 (N_15424,N_14392,N_14621);
or U15425 (N_15425,N_14518,N_14869);
nand U15426 (N_15426,N_14850,N_14650);
nand U15427 (N_15427,N_14389,N_14486);
or U15428 (N_15428,N_14579,N_14802);
and U15429 (N_15429,N_14984,N_14436);
and U15430 (N_15430,N_14565,N_14753);
or U15431 (N_15431,N_14932,N_14497);
and U15432 (N_15432,N_14751,N_14782);
or U15433 (N_15433,N_14701,N_14385);
nand U15434 (N_15434,N_14642,N_14592);
nand U15435 (N_15435,N_14489,N_14569);
and U15436 (N_15436,N_14754,N_14734);
nand U15437 (N_15437,N_14437,N_14905);
or U15438 (N_15438,N_14600,N_14920);
nor U15439 (N_15439,N_14964,N_14457);
nand U15440 (N_15440,N_14387,N_14982);
or U15441 (N_15441,N_14633,N_14466);
or U15442 (N_15442,N_14675,N_14759);
nand U15443 (N_15443,N_14767,N_14912);
nor U15444 (N_15444,N_14978,N_14525);
or U15445 (N_15445,N_14630,N_14855);
nor U15446 (N_15446,N_14389,N_14912);
nand U15447 (N_15447,N_14943,N_14771);
or U15448 (N_15448,N_14819,N_14751);
and U15449 (N_15449,N_14815,N_14873);
nand U15450 (N_15450,N_14501,N_14656);
or U15451 (N_15451,N_14508,N_14579);
nand U15452 (N_15452,N_14426,N_14837);
or U15453 (N_15453,N_14769,N_14544);
nor U15454 (N_15454,N_14738,N_14501);
or U15455 (N_15455,N_14512,N_14883);
nor U15456 (N_15456,N_14884,N_14873);
or U15457 (N_15457,N_14504,N_14921);
and U15458 (N_15458,N_14552,N_14855);
nor U15459 (N_15459,N_14788,N_14512);
nor U15460 (N_15460,N_14560,N_14627);
nor U15461 (N_15461,N_14757,N_14468);
nand U15462 (N_15462,N_14559,N_14512);
nor U15463 (N_15463,N_14486,N_14425);
and U15464 (N_15464,N_14994,N_14477);
or U15465 (N_15465,N_14740,N_14802);
xnor U15466 (N_15466,N_14977,N_14776);
and U15467 (N_15467,N_14735,N_14380);
and U15468 (N_15468,N_14396,N_14928);
nand U15469 (N_15469,N_14402,N_14734);
nor U15470 (N_15470,N_14832,N_14874);
nand U15471 (N_15471,N_14877,N_14889);
and U15472 (N_15472,N_14475,N_14508);
or U15473 (N_15473,N_14493,N_14604);
and U15474 (N_15474,N_14745,N_14840);
xnor U15475 (N_15475,N_14967,N_14704);
nor U15476 (N_15476,N_14948,N_14575);
nor U15477 (N_15477,N_14397,N_14973);
nor U15478 (N_15478,N_14390,N_14512);
nand U15479 (N_15479,N_14406,N_14967);
xor U15480 (N_15480,N_14831,N_14805);
nand U15481 (N_15481,N_14526,N_14568);
or U15482 (N_15482,N_14987,N_14812);
or U15483 (N_15483,N_14439,N_14932);
and U15484 (N_15484,N_14772,N_14798);
nor U15485 (N_15485,N_14644,N_14427);
nor U15486 (N_15486,N_14787,N_14744);
nand U15487 (N_15487,N_14640,N_14618);
or U15488 (N_15488,N_14500,N_14820);
nand U15489 (N_15489,N_14417,N_14453);
or U15490 (N_15490,N_14450,N_14650);
nand U15491 (N_15491,N_14546,N_14859);
nand U15492 (N_15492,N_14971,N_14613);
or U15493 (N_15493,N_14737,N_14493);
nor U15494 (N_15494,N_14760,N_14950);
nand U15495 (N_15495,N_14826,N_14375);
nor U15496 (N_15496,N_14939,N_14748);
and U15497 (N_15497,N_14603,N_14731);
and U15498 (N_15498,N_14965,N_14798);
nor U15499 (N_15499,N_14735,N_14425);
nand U15500 (N_15500,N_14491,N_14551);
and U15501 (N_15501,N_14502,N_14556);
nand U15502 (N_15502,N_14509,N_14673);
and U15503 (N_15503,N_14873,N_14858);
or U15504 (N_15504,N_14390,N_14590);
and U15505 (N_15505,N_14567,N_14777);
xor U15506 (N_15506,N_14904,N_14434);
and U15507 (N_15507,N_14958,N_14418);
nor U15508 (N_15508,N_14764,N_14595);
nand U15509 (N_15509,N_14767,N_14664);
nor U15510 (N_15510,N_14466,N_14506);
nor U15511 (N_15511,N_14738,N_14558);
nand U15512 (N_15512,N_14849,N_14916);
nor U15513 (N_15513,N_14514,N_14761);
or U15514 (N_15514,N_14416,N_14553);
and U15515 (N_15515,N_14463,N_14961);
and U15516 (N_15516,N_14528,N_14977);
nor U15517 (N_15517,N_14869,N_14445);
nor U15518 (N_15518,N_14646,N_14671);
nand U15519 (N_15519,N_14380,N_14647);
nand U15520 (N_15520,N_14646,N_14635);
nand U15521 (N_15521,N_14881,N_14702);
nand U15522 (N_15522,N_14986,N_14631);
xnor U15523 (N_15523,N_14790,N_14715);
and U15524 (N_15524,N_14653,N_14758);
xnor U15525 (N_15525,N_14827,N_14815);
and U15526 (N_15526,N_14825,N_14748);
nor U15527 (N_15527,N_14432,N_14936);
nor U15528 (N_15528,N_14804,N_14415);
nand U15529 (N_15529,N_14678,N_14849);
and U15530 (N_15530,N_14879,N_14933);
nor U15531 (N_15531,N_14807,N_14808);
nor U15532 (N_15532,N_14574,N_14771);
nor U15533 (N_15533,N_14456,N_14896);
nor U15534 (N_15534,N_14889,N_14617);
xor U15535 (N_15535,N_14507,N_14680);
and U15536 (N_15536,N_14941,N_14812);
and U15537 (N_15537,N_14889,N_14958);
or U15538 (N_15538,N_14395,N_14975);
xor U15539 (N_15539,N_14718,N_14695);
or U15540 (N_15540,N_14419,N_14998);
nand U15541 (N_15541,N_14955,N_14423);
and U15542 (N_15542,N_14412,N_14557);
nor U15543 (N_15543,N_14596,N_14375);
nand U15544 (N_15544,N_14679,N_14913);
or U15545 (N_15545,N_14672,N_14919);
xnor U15546 (N_15546,N_14710,N_14706);
nand U15547 (N_15547,N_14763,N_14554);
nor U15548 (N_15548,N_14504,N_14639);
nand U15549 (N_15549,N_14597,N_14449);
or U15550 (N_15550,N_14846,N_14929);
and U15551 (N_15551,N_14556,N_14465);
nor U15552 (N_15552,N_14597,N_14887);
nand U15553 (N_15553,N_14795,N_14728);
nand U15554 (N_15554,N_14422,N_14916);
and U15555 (N_15555,N_14729,N_14747);
nor U15556 (N_15556,N_14427,N_14430);
nor U15557 (N_15557,N_14906,N_14603);
nand U15558 (N_15558,N_14681,N_14878);
and U15559 (N_15559,N_14560,N_14866);
nand U15560 (N_15560,N_14376,N_14485);
nor U15561 (N_15561,N_14808,N_14843);
nor U15562 (N_15562,N_14462,N_14649);
nand U15563 (N_15563,N_14573,N_14988);
nor U15564 (N_15564,N_14910,N_14540);
nor U15565 (N_15565,N_14699,N_14627);
nand U15566 (N_15566,N_14461,N_14530);
nand U15567 (N_15567,N_14565,N_14911);
or U15568 (N_15568,N_14679,N_14966);
xor U15569 (N_15569,N_14612,N_14881);
nand U15570 (N_15570,N_14749,N_14673);
or U15571 (N_15571,N_14731,N_14610);
or U15572 (N_15572,N_14995,N_14702);
or U15573 (N_15573,N_14984,N_14611);
nor U15574 (N_15574,N_14859,N_14381);
and U15575 (N_15575,N_14837,N_14600);
nand U15576 (N_15576,N_14530,N_14980);
nand U15577 (N_15577,N_14577,N_14575);
nor U15578 (N_15578,N_14938,N_14778);
or U15579 (N_15579,N_14381,N_14928);
xor U15580 (N_15580,N_14705,N_14471);
nand U15581 (N_15581,N_14613,N_14502);
nor U15582 (N_15582,N_14894,N_14711);
or U15583 (N_15583,N_14535,N_14695);
nand U15584 (N_15584,N_14678,N_14508);
nand U15585 (N_15585,N_14590,N_14974);
nand U15586 (N_15586,N_14747,N_14712);
nor U15587 (N_15587,N_14567,N_14614);
and U15588 (N_15588,N_14593,N_14420);
nand U15589 (N_15589,N_14536,N_14886);
xor U15590 (N_15590,N_14703,N_14525);
nor U15591 (N_15591,N_14473,N_14859);
nand U15592 (N_15592,N_14746,N_14540);
nor U15593 (N_15593,N_14736,N_14548);
nor U15594 (N_15594,N_14858,N_14741);
nand U15595 (N_15595,N_14688,N_14888);
or U15596 (N_15596,N_14485,N_14551);
nand U15597 (N_15597,N_14713,N_14945);
or U15598 (N_15598,N_14838,N_14942);
or U15599 (N_15599,N_14946,N_14713);
and U15600 (N_15600,N_14412,N_14584);
nor U15601 (N_15601,N_14579,N_14694);
xnor U15602 (N_15602,N_14798,N_14776);
nand U15603 (N_15603,N_14699,N_14537);
or U15604 (N_15604,N_14473,N_14780);
and U15605 (N_15605,N_14583,N_14667);
nor U15606 (N_15606,N_14541,N_14500);
and U15607 (N_15607,N_14989,N_14780);
or U15608 (N_15608,N_14783,N_14538);
nand U15609 (N_15609,N_14844,N_14840);
nor U15610 (N_15610,N_14626,N_14893);
nand U15611 (N_15611,N_14453,N_14521);
nor U15612 (N_15612,N_14669,N_14848);
nand U15613 (N_15613,N_14687,N_14991);
xnor U15614 (N_15614,N_14561,N_14868);
or U15615 (N_15615,N_14379,N_14592);
xor U15616 (N_15616,N_14705,N_14893);
nor U15617 (N_15617,N_14839,N_14843);
nand U15618 (N_15618,N_14876,N_14787);
nand U15619 (N_15619,N_14642,N_14514);
or U15620 (N_15620,N_14410,N_14942);
nor U15621 (N_15621,N_14409,N_14553);
or U15622 (N_15622,N_14743,N_14864);
xnor U15623 (N_15623,N_14733,N_14966);
nand U15624 (N_15624,N_14860,N_14990);
or U15625 (N_15625,N_15287,N_15544);
nand U15626 (N_15626,N_15087,N_15161);
or U15627 (N_15627,N_15591,N_15204);
xor U15628 (N_15628,N_15130,N_15072);
nor U15629 (N_15629,N_15488,N_15564);
or U15630 (N_15630,N_15592,N_15430);
or U15631 (N_15631,N_15189,N_15498);
nand U15632 (N_15632,N_15390,N_15433);
or U15633 (N_15633,N_15469,N_15594);
or U15634 (N_15634,N_15445,N_15090);
or U15635 (N_15635,N_15079,N_15292);
nand U15636 (N_15636,N_15303,N_15426);
nand U15637 (N_15637,N_15493,N_15370);
or U15638 (N_15638,N_15552,N_15455);
or U15639 (N_15639,N_15463,N_15240);
nor U15640 (N_15640,N_15320,N_15521);
and U15641 (N_15641,N_15329,N_15360);
nor U15642 (N_15642,N_15295,N_15143);
nor U15643 (N_15643,N_15378,N_15182);
xor U15644 (N_15644,N_15089,N_15050);
nor U15645 (N_15645,N_15271,N_15096);
xor U15646 (N_15646,N_15480,N_15407);
and U15647 (N_15647,N_15137,N_15416);
or U15648 (N_15648,N_15155,N_15487);
and U15649 (N_15649,N_15436,N_15230);
xnor U15650 (N_15650,N_15044,N_15525);
nand U15651 (N_15651,N_15421,N_15032);
nor U15652 (N_15652,N_15123,N_15315);
xnor U15653 (N_15653,N_15457,N_15034);
nand U15654 (N_15654,N_15492,N_15502);
or U15655 (N_15655,N_15567,N_15250);
and U15656 (N_15656,N_15424,N_15356);
nor U15657 (N_15657,N_15105,N_15289);
and U15658 (N_15658,N_15254,N_15031);
or U15659 (N_15659,N_15337,N_15039);
nand U15660 (N_15660,N_15414,N_15067);
and U15661 (N_15661,N_15185,N_15569);
xnor U15662 (N_15662,N_15226,N_15372);
and U15663 (N_15663,N_15474,N_15222);
nand U15664 (N_15664,N_15456,N_15175);
and U15665 (N_15665,N_15037,N_15194);
and U15666 (N_15666,N_15348,N_15125);
xnor U15667 (N_15667,N_15396,N_15177);
nand U15668 (N_15668,N_15410,N_15604);
or U15669 (N_15669,N_15460,N_15237);
or U15670 (N_15670,N_15003,N_15023);
or U15671 (N_15671,N_15092,N_15326);
nand U15672 (N_15672,N_15160,N_15363);
and U15673 (N_15673,N_15409,N_15027);
and U15674 (N_15674,N_15179,N_15305);
xnor U15675 (N_15675,N_15539,N_15425);
and U15676 (N_15676,N_15111,N_15076);
xor U15677 (N_15677,N_15002,N_15614);
xnor U15678 (N_15678,N_15412,N_15556);
nand U15679 (N_15679,N_15098,N_15064);
nand U15680 (N_15680,N_15586,N_15578);
nand U15681 (N_15681,N_15309,N_15188);
or U15682 (N_15682,N_15281,N_15499);
nand U15683 (N_15683,N_15324,N_15013);
nand U15684 (N_15684,N_15475,N_15359);
or U15685 (N_15685,N_15261,N_15559);
nand U15686 (N_15686,N_15308,N_15503);
or U15687 (N_15687,N_15572,N_15550);
nor U15688 (N_15688,N_15065,N_15181);
xnor U15689 (N_15689,N_15357,N_15236);
nor U15690 (N_15690,N_15104,N_15202);
xnor U15691 (N_15691,N_15134,N_15273);
xnor U15692 (N_15692,N_15267,N_15015);
xnor U15693 (N_15693,N_15443,N_15132);
and U15694 (N_15694,N_15114,N_15333);
nor U15695 (N_15695,N_15063,N_15220);
nor U15696 (N_15696,N_15611,N_15485);
nand U15697 (N_15697,N_15570,N_15477);
xnor U15698 (N_15698,N_15163,N_15514);
and U15699 (N_15699,N_15352,N_15124);
and U15700 (N_15700,N_15468,N_15355);
and U15701 (N_15701,N_15540,N_15330);
nand U15702 (N_15702,N_15444,N_15447);
nor U15703 (N_15703,N_15579,N_15035);
or U15704 (N_15704,N_15523,N_15342);
xor U15705 (N_15705,N_15047,N_15112);
nor U15706 (N_15706,N_15500,N_15393);
or U15707 (N_15707,N_15555,N_15347);
xnor U15708 (N_15708,N_15619,N_15154);
xor U15709 (N_15709,N_15312,N_15235);
nand U15710 (N_15710,N_15127,N_15209);
or U15711 (N_15711,N_15613,N_15253);
xnor U15712 (N_15712,N_15007,N_15541);
nor U15713 (N_15713,N_15300,N_15077);
and U15714 (N_15714,N_15429,N_15590);
and U15715 (N_15715,N_15319,N_15120);
nand U15716 (N_15716,N_15562,N_15070);
or U15717 (N_15717,N_15138,N_15263);
or U15718 (N_15718,N_15233,N_15068);
or U15719 (N_15719,N_15511,N_15528);
nand U15720 (N_15720,N_15054,N_15207);
nand U15721 (N_15721,N_15394,N_15078);
and U15722 (N_15722,N_15301,N_15546);
nand U15723 (N_15723,N_15479,N_15509);
xnor U15724 (N_15724,N_15024,N_15071);
or U15725 (N_15725,N_15527,N_15100);
and U15726 (N_15726,N_15505,N_15400);
nor U15727 (N_15727,N_15561,N_15009);
nor U15728 (N_15728,N_15616,N_15317);
nor U15729 (N_15729,N_15219,N_15141);
and U15730 (N_15730,N_15291,N_15368);
nor U15731 (N_15731,N_15200,N_15019);
and U15732 (N_15732,N_15199,N_15406);
nor U15733 (N_15733,N_15156,N_15458);
or U15734 (N_15734,N_15473,N_15507);
or U15735 (N_15735,N_15489,N_15413);
nand U15736 (N_15736,N_15148,N_15187);
nor U15737 (N_15737,N_15059,N_15515);
nand U15738 (N_15738,N_15290,N_15530);
and U15739 (N_15739,N_15587,N_15345);
xor U15740 (N_15740,N_15617,N_15165);
nand U15741 (N_15741,N_15375,N_15022);
and U15742 (N_15742,N_15113,N_15248);
xor U15743 (N_15743,N_15102,N_15470);
nor U15744 (N_15744,N_15581,N_15296);
and U15745 (N_15745,N_15203,N_15069);
and U15746 (N_15746,N_15461,N_15385);
and U15747 (N_15747,N_15029,N_15106);
nand U15748 (N_15748,N_15325,N_15398);
nor U15749 (N_15749,N_15603,N_15331);
nand U15750 (N_15750,N_15323,N_15536);
nand U15751 (N_15751,N_15180,N_15510);
and U15752 (N_15752,N_15361,N_15216);
nor U15753 (N_15753,N_15268,N_15431);
nand U15754 (N_15754,N_15129,N_15252);
xor U15755 (N_15755,N_15304,N_15408);
nor U15756 (N_15756,N_15109,N_15198);
and U15757 (N_15757,N_15516,N_15451);
and U15758 (N_15758,N_15086,N_15467);
or U15759 (N_15759,N_15588,N_15388);
and U15760 (N_15760,N_15454,N_15103);
xor U15761 (N_15761,N_15214,N_15526);
xnor U15762 (N_15762,N_15549,N_15081);
or U15763 (N_15763,N_15051,N_15285);
nor U15764 (N_15764,N_15184,N_15450);
or U15765 (N_15765,N_15589,N_15327);
and U15766 (N_15766,N_15223,N_15508);
and U15767 (N_15767,N_15075,N_15448);
and U15768 (N_15768,N_15150,N_15313);
nand U15769 (N_15769,N_15045,N_15049);
or U15770 (N_15770,N_15293,N_15021);
nand U15771 (N_15771,N_15173,N_15597);
nand U15772 (N_15772,N_15598,N_15115);
and U15773 (N_15773,N_15418,N_15183);
nor U15774 (N_15774,N_15101,N_15332);
nor U15775 (N_15775,N_15381,N_15225);
and U15776 (N_15776,N_15575,N_15367);
or U15777 (N_15777,N_15294,N_15212);
and U15778 (N_15778,N_15191,N_15117);
nand U15779 (N_15779,N_15052,N_15283);
or U15780 (N_15780,N_15382,N_15542);
and U15781 (N_15781,N_15119,N_15437);
and U15782 (N_15782,N_15012,N_15014);
xnor U15783 (N_15783,N_15010,N_15277);
and U15784 (N_15784,N_15386,N_15001);
and U15785 (N_15785,N_15441,N_15558);
and U15786 (N_15786,N_15142,N_15284);
nand U15787 (N_15787,N_15419,N_15464);
nor U15788 (N_15788,N_15146,N_15095);
and U15789 (N_15789,N_15517,N_15380);
or U15790 (N_15790,N_15274,N_15334);
and U15791 (N_15791,N_15153,N_15335);
and U15792 (N_15792,N_15478,N_15582);
nor U15793 (N_15793,N_15311,N_15172);
or U15794 (N_15794,N_15405,N_15440);
or U15795 (N_15795,N_15073,N_15196);
nand U15796 (N_15796,N_15270,N_15205);
xor U15797 (N_15797,N_15126,N_15318);
nand U15798 (N_15798,N_15251,N_15577);
nor U15799 (N_15799,N_15535,N_15118);
xnor U15800 (N_15800,N_15099,N_15157);
and U15801 (N_15801,N_15116,N_15135);
nand U15802 (N_15802,N_15053,N_15080);
nand U15803 (N_15803,N_15612,N_15244);
xnor U15804 (N_15804,N_15434,N_15538);
xor U15805 (N_15805,N_15583,N_15066);
and U15806 (N_15806,N_15446,N_15260);
nor U15807 (N_15807,N_15600,N_15084);
nor U15808 (N_15808,N_15545,N_15322);
or U15809 (N_15809,N_15030,N_15082);
or U15810 (N_15810,N_15085,N_15046);
nand U15811 (N_15811,N_15234,N_15346);
nand U15812 (N_15812,N_15178,N_15306);
nor U15813 (N_15813,N_15238,N_15055);
or U15814 (N_15814,N_15415,N_15159);
nand U15815 (N_15815,N_15504,N_15056);
and U15816 (N_15816,N_15403,N_15497);
and U15817 (N_15817,N_15008,N_15288);
and U15818 (N_15818,N_15245,N_15350);
and U15819 (N_15819,N_15195,N_15602);
nand U15820 (N_15820,N_15547,N_15224);
nand U15821 (N_15821,N_15481,N_15266);
nand U15822 (N_15822,N_15354,N_15610);
nand U15823 (N_15823,N_15036,N_15383);
or U15824 (N_15824,N_15227,N_15608);
nor U15825 (N_15825,N_15341,N_15307);
or U15826 (N_15826,N_15269,N_15422);
nor U15827 (N_15827,N_15338,N_15091);
or U15828 (N_15828,N_15484,N_15491);
or U15829 (N_15829,N_15279,N_15162);
and U15830 (N_15830,N_15495,N_15038);
or U15831 (N_15831,N_15190,N_15276);
and U15832 (N_15832,N_15232,N_15620);
nand U15833 (N_15833,N_15147,N_15192);
and U15834 (N_15834,N_15257,N_15262);
or U15835 (N_15835,N_15272,N_15171);
and U15836 (N_15836,N_15229,N_15353);
or U15837 (N_15837,N_15011,N_15041);
nor U15838 (N_15838,N_15374,N_15373);
and U15839 (N_15839,N_15060,N_15551);
xor U15840 (N_15840,N_15197,N_15623);
or U15841 (N_15841,N_15399,N_15524);
and U15842 (N_15842,N_15483,N_15122);
nand U15843 (N_15843,N_15040,N_15417);
nand U15844 (N_15844,N_15379,N_15439);
nor U15845 (N_15845,N_15151,N_15404);
nor U15846 (N_15846,N_15449,N_15074);
or U15847 (N_15847,N_15249,N_15108);
nand U15848 (N_15848,N_15553,N_15364);
nand U15849 (N_15849,N_15210,N_15618);
or U15850 (N_15850,N_15343,N_15482);
nor U15851 (N_15851,N_15606,N_15573);
and U15852 (N_15852,N_15624,N_15533);
nor U15853 (N_15853,N_15365,N_15256);
or U15854 (N_15854,N_15158,N_15043);
nor U15855 (N_15855,N_15377,N_15278);
nor U15856 (N_15856,N_15133,N_15593);
and U15857 (N_15857,N_15371,N_15428);
xor U15858 (N_15858,N_15000,N_15366);
nor U15859 (N_15859,N_15453,N_15004);
xnor U15860 (N_15860,N_15174,N_15208);
and U15861 (N_15861,N_15088,N_15358);
or U15862 (N_15862,N_15144,N_15241);
or U15863 (N_15863,N_15369,N_15391);
nand U15864 (N_15864,N_15297,N_15136);
or U15865 (N_15865,N_15420,N_15093);
nand U15866 (N_15866,N_15411,N_15595);
nor U15867 (N_15867,N_15152,N_15242);
nand U15868 (N_15868,N_15615,N_15452);
and U15869 (N_15869,N_15519,N_15494);
or U15870 (N_15870,N_15310,N_15435);
and U15871 (N_15871,N_15344,N_15282);
nand U15872 (N_15872,N_15228,N_15264);
and U15873 (N_15873,N_15258,N_15275);
and U15874 (N_15874,N_15490,N_15328);
or U15875 (N_15875,N_15472,N_15042);
and U15876 (N_15876,N_15048,N_15255);
nor U15877 (N_15877,N_15609,N_15351);
and U15878 (N_15878,N_15402,N_15299);
xnor U15879 (N_15879,N_15164,N_15548);
nor U15880 (N_15880,N_15336,N_15231);
xnor U15881 (N_15881,N_15427,N_15557);
xor U15882 (N_15882,N_15221,N_15362);
nor U15883 (N_15883,N_15585,N_15496);
nor U15884 (N_15884,N_15280,N_15574);
xnor U15885 (N_15885,N_15518,N_15286);
nor U15886 (N_15886,N_15442,N_15349);
and U15887 (N_15887,N_15168,N_15061);
or U15888 (N_15888,N_15601,N_15128);
and U15889 (N_15889,N_15563,N_15139);
nor U15890 (N_15890,N_15599,N_15376);
and U15891 (N_15891,N_15097,N_15094);
or U15892 (N_15892,N_15395,N_15176);
nor U15893 (N_15893,N_15018,N_15576);
nand U15894 (N_15894,N_15016,N_15321);
and U15895 (N_15895,N_15083,N_15476);
nor U15896 (N_15896,N_15387,N_15466);
nor U15897 (N_15897,N_15543,N_15215);
and U15898 (N_15898,N_15607,N_15513);
and U15899 (N_15899,N_15298,N_15392);
nor U15900 (N_15900,N_15217,N_15584);
or U15901 (N_15901,N_15486,N_15167);
and U15902 (N_15902,N_15314,N_15622);
and U15903 (N_15903,N_15020,N_15246);
nor U15904 (N_15904,N_15057,N_15501);
nand U15905 (N_15905,N_15512,N_15140);
and U15906 (N_15906,N_15537,N_15397);
nand U15907 (N_15907,N_15432,N_15520);
nand U15908 (N_15908,N_15531,N_15529);
nand U15909 (N_15909,N_15423,N_15596);
nand U15910 (N_15910,N_15121,N_15149);
nor U15911 (N_15911,N_15028,N_15033);
and U15912 (N_15912,N_15206,N_15005);
nor U15913 (N_15913,N_15170,N_15247);
nand U15914 (N_15914,N_15568,N_15239);
nand U15915 (N_15915,N_15384,N_15107);
nor U15916 (N_15916,N_15259,N_15302);
nand U15917 (N_15917,N_15459,N_15506);
nand U15918 (N_15918,N_15218,N_15131);
or U15919 (N_15919,N_15465,N_15438);
nand U15920 (N_15920,N_15605,N_15339);
nand U15921 (N_15921,N_15213,N_15389);
and U15922 (N_15922,N_15571,N_15265);
or U15923 (N_15923,N_15062,N_15462);
nand U15924 (N_15924,N_15560,N_15166);
and U15925 (N_15925,N_15169,N_15058);
or U15926 (N_15926,N_15186,N_15017);
and U15927 (N_15927,N_15401,N_15193);
xor U15928 (N_15928,N_15534,N_15243);
nor U15929 (N_15929,N_15145,N_15211);
xnor U15930 (N_15930,N_15110,N_15025);
nand U15931 (N_15931,N_15532,N_15554);
and U15932 (N_15932,N_15621,N_15316);
or U15933 (N_15933,N_15580,N_15026);
nand U15934 (N_15934,N_15471,N_15522);
xnor U15935 (N_15935,N_15565,N_15566);
and U15936 (N_15936,N_15340,N_15006);
and U15937 (N_15937,N_15201,N_15430);
xnor U15938 (N_15938,N_15347,N_15093);
nand U15939 (N_15939,N_15239,N_15023);
nor U15940 (N_15940,N_15250,N_15031);
nand U15941 (N_15941,N_15525,N_15556);
and U15942 (N_15942,N_15062,N_15105);
and U15943 (N_15943,N_15561,N_15057);
nor U15944 (N_15944,N_15484,N_15312);
nand U15945 (N_15945,N_15437,N_15201);
and U15946 (N_15946,N_15386,N_15547);
and U15947 (N_15947,N_15121,N_15131);
or U15948 (N_15948,N_15126,N_15117);
nor U15949 (N_15949,N_15613,N_15086);
nor U15950 (N_15950,N_15497,N_15104);
nor U15951 (N_15951,N_15139,N_15069);
xor U15952 (N_15952,N_15298,N_15487);
xnor U15953 (N_15953,N_15577,N_15111);
or U15954 (N_15954,N_15569,N_15032);
nand U15955 (N_15955,N_15296,N_15183);
and U15956 (N_15956,N_15210,N_15584);
xnor U15957 (N_15957,N_15242,N_15416);
and U15958 (N_15958,N_15293,N_15471);
and U15959 (N_15959,N_15048,N_15240);
nor U15960 (N_15960,N_15140,N_15195);
nor U15961 (N_15961,N_15147,N_15156);
nor U15962 (N_15962,N_15298,N_15386);
and U15963 (N_15963,N_15114,N_15010);
or U15964 (N_15964,N_15279,N_15252);
and U15965 (N_15965,N_15351,N_15369);
or U15966 (N_15966,N_15082,N_15305);
nor U15967 (N_15967,N_15620,N_15303);
nand U15968 (N_15968,N_15051,N_15289);
and U15969 (N_15969,N_15138,N_15542);
or U15970 (N_15970,N_15060,N_15316);
nor U15971 (N_15971,N_15015,N_15377);
nand U15972 (N_15972,N_15192,N_15361);
xnor U15973 (N_15973,N_15390,N_15499);
xor U15974 (N_15974,N_15230,N_15548);
nor U15975 (N_15975,N_15493,N_15099);
or U15976 (N_15976,N_15610,N_15301);
or U15977 (N_15977,N_15094,N_15082);
nand U15978 (N_15978,N_15288,N_15440);
and U15979 (N_15979,N_15075,N_15109);
and U15980 (N_15980,N_15278,N_15417);
or U15981 (N_15981,N_15595,N_15120);
or U15982 (N_15982,N_15035,N_15117);
nand U15983 (N_15983,N_15151,N_15181);
xnor U15984 (N_15984,N_15014,N_15441);
xnor U15985 (N_15985,N_15103,N_15374);
and U15986 (N_15986,N_15370,N_15469);
and U15987 (N_15987,N_15167,N_15120);
nand U15988 (N_15988,N_15608,N_15581);
or U15989 (N_15989,N_15075,N_15500);
xor U15990 (N_15990,N_15534,N_15558);
nand U15991 (N_15991,N_15059,N_15353);
or U15992 (N_15992,N_15469,N_15106);
or U15993 (N_15993,N_15071,N_15240);
nand U15994 (N_15994,N_15357,N_15561);
nor U15995 (N_15995,N_15239,N_15612);
nor U15996 (N_15996,N_15184,N_15051);
xor U15997 (N_15997,N_15488,N_15618);
or U15998 (N_15998,N_15312,N_15491);
nand U15999 (N_15999,N_15484,N_15128);
or U16000 (N_16000,N_15558,N_15492);
nor U16001 (N_16001,N_15168,N_15592);
nor U16002 (N_16002,N_15179,N_15531);
or U16003 (N_16003,N_15370,N_15169);
nor U16004 (N_16004,N_15304,N_15425);
nor U16005 (N_16005,N_15515,N_15098);
and U16006 (N_16006,N_15449,N_15183);
nor U16007 (N_16007,N_15255,N_15383);
or U16008 (N_16008,N_15280,N_15468);
xor U16009 (N_16009,N_15006,N_15594);
nor U16010 (N_16010,N_15200,N_15110);
and U16011 (N_16011,N_15263,N_15594);
and U16012 (N_16012,N_15221,N_15584);
nor U16013 (N_16013,N_15270,N_15524);
and U16014 (N_16014,N_15151,N_15613);
or U16015 (N_16015,N_15591,N_15134);
or U16016 (N_16016,N_15372,N_15604);
and U16017 (N_16017,N_15114,N_15495);
and U16018 (N_16018,N_15612,N_15387);
and U16019 (N_16019,N_15083,N_15070);
or U16020 (N_16020,N_15099,N_15215);
or U16021 (N_16021,N_15382,N_15393);
xnor U16022 (N_16022,N_15304,N_15017);
nand U16023 (N_16023,N_15322,N_15195);
xnor U16024 (N_16024,N_15546,N_15023);
nor U16025 (N_16025,N_15557,N_15114);
xnor U16026 (N_16026,N_15514,N_15087);
nand U16027 (N_16027,N_15380,N_15559);
nand U16028 (N_16028,N_15169,N_15570);
xor U16029 (N_16029,N_15443,N_15010);
xnor U16030 (N_16030,N_15461,N_15263);
nor U16031 (N_16031,N_15620,N_15375);
nor U16032 (N_16032,N_15420,N_15098);
and U16033 (N_16033,N_15240,N_15622);
and U16034 (N_16034,N_15157,N_15228);
and U16035 (N_16035,N_15009,N_15323);
and U16036 (N_16036,N_15182,N_15415);
and U16037 (N_16037,N_15298,N_15186);
and U16038 (N_16038,N_15222,N_15076);
and U16039 (N_16039,N_15344,N_15186);
or U16040 (N_16040,N_15580,N_15418);
nor U16041 (N_16041,N_15188,N_15493);
or U16042 (N_16042,N_15213,N_15545);
or U16043 (N_16043,N_15589,N_15366);
nor U16044 (N_16044,N_15111,N_15037);
nand U16045 (N_16045,N_15135,N_15281);
xnor U16046 (N_16046,N_15367,N_15401);
or U16047 (N_16047,N_15367,N_15072);
and U16048 (N_16048,N_15558,N_15509);
or U16049 (N_16049,N_15144,N_15253);
and U16050 (N_16050,N_15563,N_15451);
nand U16051 (N_16051,N_15528,N_15212);
xor U16052 (N_16052,N_15439,N_15497);
or U16053 (N_16053,N_15136,N_15010);
and U16054 (N_16054,N_15094,N_15297);
and U16055 (N_16055,N_15624,N_15431);
nor U16056 (N_16056,N_15157,N_15246);
nor U16057 (N_16057,N_15164,N_15157);
nand U16058 (N_16058,N_15319,N_15122);
xor U16059 (N_16059,N_15046,N_15144);
or U16060 (N_16060,N_15138,N_15360);
or U16061 (N_16061,N_15442,N_15200);
and U16062 (N_16062,N_15467,N_15620);
nor U16063 (N_16063,N_15089,N_15422);
or U16064 (N_16064,N_15309,N_15146);
and U16065 (N_16065,N_15158,N_15324);
nand U16066 (N_16066,N_15320,N_15080);
or U16067 (N_16067,N_15440,N_15497);
and U16068 (N_16068,N_15529,N_15098);
and U16069 (N_16069,N_15103,N_15110);
and U16070 (N_16070,N_15550,N_15500);
nor U16071 (N_16071,N_15076,N_15034);
xnor U16072 (N_16072,N_15084,N_15023);
nand U16073 (N_16073,N_15347,N_15203);
xnor U16074 (N_16074,N_15339,N_15189);
xnor U16075 (N_16075,N_15044,N_15062);
nand U16076 (N_16076,N_15503,N_15445);
xnor U16077 (N_16077,N_15109,N_15471);
nor U16078 (N_16078,N_15292,N_15003);
xnor U16079 (N_16079,N_15539,N_15485);
xnor U16080 (N_16080,N_15419,N_15093);
nand U16081 (N_16081,N_15422,N_15081);
nor U16082 (N_16082,N_15146,N_15247);
or U16083 (N_16083,N_15566,N_15403);
nand U16084 (N_16084,N_15527,N_15128);
or U16085 (N_16085,N_15361,N_15512);
nand U16086 (N_16086,N_15118,N_15487);
or U16087 (N_16087,N_15235,N_15515);
nor U16088 (N_16088,N_15489,N_15171);
and U16089 (N_16089,N_15266,N_15001);
nor U16090 (N_16090,N_15308,N_15556);
nand U16091 (N_16091,N_15605,N_15341);
or U16092 (N_16092,N_15251,N_15229);
nor U16093 (N_16093,N_15377,N_15539);
nor U16094 (N_16094,N_15449,N_15222);
xnor U16095 (N_16095,N_15549,N_15250);
and U16096 (N_16096,N_15301,N_15519);
nor U16097 (N_16097,N_15227,N_15059);
nor U16098 (N_16098,N_15076,N_15472);
and U16099 (N_16099,N_15284,N_15365);
nor U16100 (N_16100,N_15238,N_15466);
nand U16101 (N_16101,N_15230,N_15190);
and U16102 (N_16102,N_15538,N_15052);
nor U16103 (N_16103,N_15004,N_15581);
xnor U16104 (N_16104,N_15511,N_15055);
xnor U16105 (N_16105,N_15031,N_15052);
and U16106 (N_16106,N_15564,N_15451);
nand U16107 (N_16107,N_15101,N_15127);
and U16108 (N_16108,N_15372,N_15488);
nor U16109 (N_16109,N_15289,N_15452);
and U16110 (N_16110,N_15037,N_15383);
or U16111 (N_16111,N_15104,N_15053);
nand U16112 (N_16112,N_15033,N_15094);
nor U16113 (N_16113,N_15137,N_15211);
and U16114 (N_16114,N_15033,N_15153);
or U16115 (N_16115,N_15262,N_15496);
nor U16116 (N_16116,N_15225,N_15396);
nand U16117 (N_16117,N_15393,N_15620);
nand U16118 (N_16118,N_15557,N_15172);
nand U16119 (N_16119,N_15575,N_15002);
nor U16120 (N_16120,N_15463,N_15522);
xor U16121 (N_16121,N_15333,N_15244);
nand U16122 (N_16122,N_15212,N_15154);
or U16123 (N_16123,N_15211,N_15193);
xnor U16124 (N_16124,N_15111,N_15192);
nor U16125 (N_16125,N_15175,N_15255);
nor U16126 (N_16126,N_15176,N_15040);
nand U16127 (N_16127,N_15142,N_15513);
or U16128 (N_16128,N_15258,N_15333);
or U16129 (N_16129,N_15369,N_15567);
or U16130 (N_16130,N_15244,N_15437);
nand U16131 (N_16131,N_15586,N_15470);
or U16132 (N_16132,N_15197,N_15527);
nand U16133 (N_16133,N_15483,N_15352);
nand U16134 (N_16134,N_15605,N_15007);
and U16135 (N_16135,N_15353,N_15369);
nand U16136 (N_16136,N_15231,N_15437);
nor U16137 (N_16137,N_15551,N_15439);
or U16138 (N_16138,N_15375,N_15569);
or U16139 (N_16139,N_15374,N_15229);
or U16140 (N_16140,N_15191,N_15545);
nor U16141 (N_16141,N_15427,N_15376);
nand U16142 (N_16142,N_15582,N_15555);
and U16143 (N_16143,N_15209,N_15151);
and U16144 (N_16144,N_15069,N_15386);
or U16145 (N_16145,N_15384,N_15414);
and U16146 (N_16146,N_15394,N_15087);
nand U16147 (N_16147,N_15339,N_15350);
or U16148 (N_16148,N_15413,N_15605);
and U16149 (N_16149,N_15479,N_15578);
or U16150 (N_16150,N_15240,N_15103);
nand U16151 (N_16151,N_15517,N_15459);
and U16152 (N_16152,N_15405,N_15076);
xnor U16153 (N_16153,N_15430,N_15519);
nor U16154 (N_16154,N_15066,N_15429);
and U16155 (N_16155,N_15543,N_15161);
and U16156 (N_16156,N_15606,N_15604);
nand U16157 (N_16157,N_15284,N_15250);
and U16158 (N_16158,N_15001,N_15623);
nand U16159 (N_16159,N_15071,N_15574);
and U16160 (N_16160,N_15219,N_15602);
nand U16161 (N_16161,N_15314,N_15075);
nand U16162 (N_16162,N_15341,N_15087);
and U16163 (N_16163,N_15379,N_15246);
and U16164 (N_16164,N_15259,N_15112);
nor U16165 (N_16165,N_15304,N_15215);
and U16166 (N_16166,N_15229,N_15009);
nand U16167 (N_16167,N_15623,N_15268);
nand U16168 (N_16168,N_15025,N_15315);
and U16169 (N_16169,N_15546,N_15551);
or U16170 (N_16170,N_15278,N_15594);
and U16171 (N_16171,N_15134,N_15586);
or U16172 (N_16172,N_15536,N_15437);
nor U16173 (N_16173,N_15083,N_15571);
xor U16174 (N_16174,N_15101,N_15590);
or U16175 (N_16175,N_15550,N_15142);
nand U16176 (N_16176,N_15402,N_15134);
nor U16177 (N_16177,N_15308,N_15363);
xnor U16178 (N_16178,N_15009,N_15091);
nand U16179 (N_16179,N_15120,N_15402);
or U16180 (N_16180,N_15467,N_15122);
or U16181 (N_16181,N_15034,N_15242);
nand U16182 (N_16182,N_15530,N_15043);
nand U16183 (N_16183,N_15447,N_15187);
or U16184 (N_16184,N_15154,N_15181);
nor U16185 (N_16185,N_15121,N_15383);
or U16186 (N_16186,N_15102,N_15589);
or U16187 (N_16187,N_15574,N_15257);
and U16188 (N_16188,N_15200,N_15409);
nand U16189 (N_16189,N_15568,N_15248);
and U16190 (N_16190,N_15482,N_15336);
nand U16191 (N_16191,N_15532,N_15363);
nand U16192 (N_16192,N_15451,N_15200);
or U16193 (N_16193,N_15504,N_15539);
and U16194 (N_16194,N_15047,N_15045);
and U16195 (N_16195,N_15399,N_15241);
and U16196 (N_16196,N_15190,N_15605);
nand U16197 (N_16197,N_15015,N_15276);
nand U16198 (N_16198,N_15062,N_15270);
nor U16199 (N_16199,N_15582,N_15122);
or U16200 (N_16200,N_15198,N_15489);
and U16201 (N_16201,N_15502,N_15032);
nand U16202 (N_16202,N_15531,N_15514);
nand U16203 (N_16203,N_15176,N_15164);
xnor U16204 (N_16204,N_15349,N_15275);
nor U16205 (N_16205,N_15246,N_15023);
or U16206 (N_16206,N_15203,N_15578);
nand U16207 (N_16207,N_15357,N_15504);
xnor U16208 (N_16208,N_15526,N_15148);
or U16209 (N_16209,N_15465,N_15065);
or U16210 (N_16210,N_15120,N_15448);
xnor U16211 (N_16211,N_15030,N_15557);
or U16212 (N_16212,N_15168,N_15608);
or U16213 (N_16213,N_15292,N_15170);
nand U16214 (N_16214,N_15420,N_15176);
nor U16215 (N_16215,N_15527,N_15328);
or U16216 (N_16216,N_15528,N_15268);
and U16217 (N_16217,N_15371,N_15433);
or U16218 (N_16218,N_15443,N_15327);
or U16219 (N_16219,N_15114,N_15210);
and U16220 (N_16220,N_15487,N_15449);
nor U16221 (N_16221,N_15249,N_15202);
and U16222 (N_16222,N_15348,N_15182);
and U16223 (N_16223,N_15209,N_15376);
nor U16224 (N_16224,N_15122,N_15267);
or U16225 (N_16225,N_15051,N_15178);
xor U16226 (N_16226,N_15539,N_15505);
nand U16227 (N_16227,N_15299,N_15416);
nor U16228 (N_16228,N_15285,N_15128);
nor U16229 (N_16229,N_15589,N_15360);
and U16230 (N_16230,N_15228,N_15386);
xnor U16231 (N_16231,N_15193,N_15346);
and U16232 (N_16232,N_15388,N_15408);
nor U16233 (N_16233,N_15087,N_15177);
nand U16234 (N_16234,N_15393,N_15314);
or U16235 (N_16235,N_15192,N_15454);
nand U16236 (N_16236,N_15286,N_15526);
or U16237 (N_16237,N_15552,N_15469);
nor U16238 (N_16238,N_15499,N_15065);
nor U16239 (N_16239,N_15080,N_15334);
nor U16240 (N_16240,N_15261,N_15381);
and U16241 (N_16241,N_15593,N_15002);
nor U16242 (N_16242,N_15362,N_15206);
or U16243 (N_16243,N_15234,N_15404);
or U16244 (N_16244,N_15005,N_15214);
xnor U16245 (N_16245,N_15229,N_15100);
and U16246 (N_16246,N_15153,N_15232);
xor U16247 (N_16247,N_15378,N_15030);
and U16248 (N_16248,N_15116,N_15261);
nand U16249 (N_16249,N_15046,N_15302);
nand U16250 (N_16250,N_16126,N_15649);
or U16251 (N_16251,N_16005,N_16145);
nand U16252 (N_16252,N_15996,N_15703);
nor U16253 (N_16253,N_16090,N_15732);
nand U16254 (N_16254,N_15652,N_16172);
nor U16255 (N_16255,N_16021,N_15745);
or U16256 (N_16256,N_15672,N_15923);
or U16257 (N_16257,N_15846,N_15844);
and U16258 (N_16258,N_15637,N_16201);
nor U16259 (N_16259,N_16100,N_15630);
nand U16260 (N_16260,N_15779,N_15663);
nand U16261 (N_16261,N_15651,N_15734);
nor U16262 (N_16262,N_15836,N_15816);
or U16263 (N_16263,N_16178,N_16241);
nor U16264 (N_16264,N_15876,N_15763);
xor U16265 (N_16265,N_15939,N_16124);
nor U16266 (N_16266,N_15947,N_15889);
or U16267 (N_16267,N_15688,N_15853);
nor U16268 (N_16268,N_15720,N_16117);
nand U16269 (N_16269,N_16052,N_15883);
nand U16270 (N_16270,N_16046,N_16038);
nand U16271 (N_16271,N_15848,N_15767);
nor U16272 (N_16272,N_16107,N_16239);
nand U16273 (N_16273,N_16249,N_15809);
nand U16274 (N_16274,N_15694,N_15768);
nand U16275 (N_16275,N_16141,N_15792);
nand U16276 (N_16276,N_15906,N_15729);
or U16277 (N_16277,N_15631,N_16160);
nand U16278 (N_16278,N_15686,N_16111);
nand U16279 (N_16279,N_16012,N_16237);
nor U16280 (N_16280,N_16133,N_15925);
xor U16281 (N_16281,N_15834,N_15981);
and U16282 (N_16282,N_15892,N_16045);
nor U16283 (N_16283,N_15695,N_15949);
nand U16284 (N_16284,N_16135,N_15691);
and U16285 (N_16285,N_16170,N_16235);
or U16286 (N_16286,N_16244,N_16054);
and U16287 (N_16287,N_16115,N_16169);
nor U16288 (N_16288,N_15887,N_15682);
or U16289 (N_16289,N_15955,N_15668);
and U16290 (N_16290,N_16043,N_15976);
nor U16291 (N_16291,N_16214,N_15904);
nor U16292 (N_16292,N_16007,N_16087);
nand U16293 (N_16293,N_15960,N_15969);
and U16294 (N_16294,N_16119,N_16068);
or U16295 (N_16295,N_15773,N_15916);
or U16296 (N_16296,N_16030,N_15967);
or U16297 (N_16297,N_15849,N_15986);
xnor U16298 (N_16298,N_15736,N_15852);
or U16299 (N_16299,N_15693,N_16226);
or U16300 (N_16300,N_15895,N_15817);
nand U16301 (N_16301,N_16089,N_15951);
nand U16302 (N_16302,N_16193,N_16158);
nand U16303 (N_16303,N_15988,N_15657);
and U16304 (N_16304,N_16078,N_16136);
or U16305 (N_16305,N_15719,N_15933);
and U16306 (N_16306,N_16002,N_16081);
and U16307 (N_16307,N_15716,N_16138);
or U16308 (N_16308,N_16173,N_16157);
nor U16309 (N_16309,N_15759,N_16000);
and U16310 (N_16310,N_16096,N_15774);
xor U16311 (N_16311,N_15869,N_15722);
or U16312 (N_16312,N_15635,N_16229);
nor U16313 (N_16313,N_15858,N_16099);
nand U16314 (N_16314,N_16001,N_15833);
and U16315 (N_16315,N_15808,N_15692);
xnor U16316 (N_16316,N_16047,N_15805);
nor U16317 (N_16317,N_16074,N_16112);
and U16318 (N_16318,N_15702,N_16025);
xor U16319 (N_16319,N_16246,N_15678);
nor U16320 (N_16320,N_15704,N_15888);
nand U16321 (N_16321,N_15675,N_15891);
or U16322 (N_16322,N_15897,N_15807);
xnor U16323 (N_16323,N_15977,N_15874);
nand U16324 (N_16324,N_15748,N_16049);
and U16325 (N_16325,N_15919,N_16220);
or U16326 (N_16326,N_15881,N_15825);
nand U16327 (N_16327,N_15655,N_15915);
or U16328 (N_16328,N_15928,N_16248);
or U16329 (N_16329,N_16080,N_15994);
nand U16330 (N_16330,N_15829,N_16195);
nor U16331 (N_16331,N_16143,N_16211);
or U16332 (N_16332,N_15903,N_16153);
nor U16333 (N_16333,N_15761,N_16148);
nand U16334 (N_16334,N_15991,N_16215);
and U16335 (N_16335,N_15721,N_15879);
nand U16336 (N_16336,N_16034,N_15975);
nor U16337 (N_16337,N_15932,N_16171);
xor U16338 (N_16338,N_15856,N_15850);
or U16339 (N_16339,N_16156,N_16183);
nor U16340 (N_16340,N_15819,N_15735);
nand U16341 (N_16341,N_16233,N_15777);
and U16342 (N_16342,N_15937,N_15868);
nor U16343 (N_16343,N_16146,N_15677);
and U16344 (N_16344,N_15841,N_15796);
and U16345 (N_16345,N_15769,N_16155);
nor U16346 (N_16346,N_16161,N_15633);
and U16347 (N_16347,N_15926,N_15942);
or U16348 (N_16348,N_15963,N_15646);
xnor U16349 (N_16349,N_15835,N_15689);
and U16350 (N_16350,N_16010,N_16026);
or U16351 (N_16351,N_16077,N_15629);
nand U16352 (N_16352,N_16037,N_15886);
and U16353 (N_16353,N_16167,N_16031);
and U16354 (N_16354,N_15627,N_15697);
nor U16355 (N_16355,N_15823,N_15950);
nor U16356 (N_16356,N_15914,N_15786);
and U16357 (N_16357,N_15638,N_15990);
or U16358 (N_16358,N_16044,N_15810);
nand U16359 (N_16359,N_15799,N_15917);
and U16360 (N_16360,N_16018,N_16088);
nand U16361 (N_16361,N_15987,N_16221);
or U16362 (N_16362,N_15860,N_15642);
and U16363 (N_16363,N_16091,N_15982);
or U16364 (N_16364,N_16102,N_15877);
nor U16365 (N_16365,N_15709,N_15656);
or U16366 (N_16366,N_16182,N_15920);
or U16367 (N_16367,N_15857,N_15793);
or U16368 (N_16368,N_15782,N_15648);
or U16369 (N_16369,N_15902,N_16056);
nand U16370 (N_16370,N_15864,N_15958);
nor U16371 (N_16371,N_15861,N_15690);
and U16372 (N_16372,N_15815,N_15780);
nor U16373 (N_16373,N_16234,N_15896);
and U16374 (N_16374,N_15900,N_16060);
and U16375 (N_16375,N_16175,N_15806);
or U16376 (N_16376,N_16042,N_15725);
nand U16377 (N_16377,N_16150,N_16217);
or U16378 (N_16378,N_15867,N_16101);
or U16379 (N_16379,N_16085,N_16152);
or U16380 (N_16380,N_15787,N_16048);
and U16381 (N_16381,N_15968,N_16216);
and U16382 (N_16382,N_16238,N_16154);
nor U16383 (N_16383,N_15760,N_16166);
nor U16384 (N_16384,N_16097,N_15973);
xnor U16385 (N_16385,N_15666,N_16165);
and U16386 (N_16386,N_15749,N_15873);
or U16387 (N_16387,N_15894,N_15643);
nor U16388 (N_16388,N_15827,N_15739);
nand U16389 (N_16389,N_15685,N_16013);
or U16390 (N_16390,N_15855,N_16128);
or U16391 (N_16391,N_16186,N_15843);
nor U16392 (N_16392,N_16140,N_16086);
xor U16393 (N_16393,N_16106,N_16011);
nand U16394 (N_16394,N_15775,N_15706);
or U16395 (N_16395,N_16240,N_15756);
or U16396 (N_16396,N_15712,N_15870);
and U16397 (N_16397,N_15899,N_16200);
and U16398 (N_16398,N_15847,N_15681);
xnor U16399 (N_16399,N_15974,N_16230);
nor U16400 (N_16400,N_16036,N_15698);
and U16401 (N_16401,N_15885,N_16118);
nand U16402 (N_16402,N_15670,N_15674);
or U16403 (N_16403,N_15845,N_15821);
nor U16404 (N_16404,N_16041,N_16016);
and U16405 (N_16405,N_15884,N_15660);
and U16406 (N_16406,N_15730,N_16070);
nand U16407 (N_16407,N_16050,N_15893);
and U16408 (N_16408,N_16065,N_15784);
nand U16409 (N_16409,N_15755,N_15764);
nand U16410 (N_16410,N_15766,N_15737);
nor U16411 (N_16411,N_16108,N_16071);
nor U16412 (N_16412,N_15723,N_16008);
nor U16413 (N_16413,N_16162,N_15872);
xor U16414 (N_16414,N_15934,N_16219);
or U16415 (N_16415,N_15828,N_16185);
xnor U16416 (N_16416,N_16123,N_15993);
and U16417 (N_16417,N_15908,N_16197);
nor U16418 (N_16418,N_15758,N_15907);
xnor U16419 (N_16419,N_15653,N_16144);
nor U16420 (N_16420,N_15992,N_15980);
or U16421 (N_16421,N_15989,N_16066);
nor U16422 (N_16422,N_15783,N_15812);
nand U16423 (N_16423,N_16192,N_16208);
or U16424 (N_16424,N_15740,N_15880);
nor U16425 (N_16425,N_15842,N_15744);
and U16426 (N_16426,N_15957,N_16039);
nor U16427 (N_16427,N_15979,N_15707);
nor U16428 (N_16428,N_16067,N_15813);
or U16429 (N_16429,N_15832,N_15822);
nand U16430 (N_16430,N_16242,N_15770);
or U16431 (N_16431,N_15634,N_15781);
nor U16432 (N_16432,N_15776,N_16130);
or U16433 (N_16433,N_15650,N_15983);
nor U16434 (N_16434,N_16147,N_16032);
and U16435 (N_16435,N_15664,N_15826);
and U16436 (N_16436,N_15927,N_15683);
or U16437 (N_16437,N_15636,N_16176);
nor U16438 (N_16438,N_16006,N_15964);
or U16439 (N_16439,N_15995,N_15715);
xnor U16440 (N_16440,N_16121,N_16062);
or U16441 (N_16441,N_15661,N_15978);
nor U16442 (N_16442,N_16209,N_16142);
nor U16443 (N_16443,N_16084,N_16207);
nand U16444 (N_16444,N_16210,N_16196);
nand U16445 (N_16445,N_16024,N_15930);
and U16446 (N_16446,N_15854,N_15938);
or U16447 (N_16447,N_15998,N_15658);
xnor U16448 (N_16448,N_15713,N_15632);
xor U16449 (N_16449,N_15999,N_16022);
and U16450 (N_16450,N_15830,N_15667);
or U16451 (N_16451,N_15862,N_16213);
nor U16452 (N_16452,N_16129,N_16203);
or U16453 (N_16453,N_16212,N_16095);
nor U16454 (N_16454,N_16190,N_15728);
or U16455 (N_16455,N_15803,N_15708);
and U16456 (N_16456,N_15785,N_15639);
and U16457 (N_16457,N_15757,N_15790);
nor U16458 (N_16458,N_15910,N_15865);
nor U16459 (N_16459,N_16028,N_15800);
and U16460 (N_16460,N_16231,N_15741);
nor U16461 (N_16461,N_16224,N_16204);
or U16462 (N_16462,N_15831,N_15673);
nand U16463 (N_16463,N_16104,N_16191);
xnor U16464 (N_16464,N_15641,N_15714);
nor U16465 (N_16465,N_16202,N_16082);
nor U16466 (N_16466,N_15985,N_16094);
xor U16467 (N_16467,N_15838,N_15724);
nor U16468 (N_16468,N_15954,N_15935);
and U16469 (N_16469,N_15727,N_16132);
xor U16470 (N_16470,N_16177,N_15762);
or U16471 (N_16471,N_15751,N_16053);
nand U16472 (N_16472,N_15645,N_16180);
nor U16473 (N_16473,N_16113,N_15753);
or U16474 (N_16474,N_15625,N_16164);
nand U16475 (N_16475,N_15684,N_15909);
nand U16476 (N_16476,N_15801,N_16227);
nor U16477 (N_16477,N_16174,N_15943);
and U16478 (N_16478,N_15898,N_16009);
or U16479 (N_16479,N_16149,N_15804);
nor U16480 (N_16480,N_15918,N_15972);
xor U16481 (N_16481,N_15901,N_16199);
or U16482 (N_16482,N_16168,N_16003);
nor U16483 (N_16483,N_16187,N_15859);
nor U16484 (N_16484,N_16223,N_15687);
nand U16485 (N_16485,N_15905,N_16073);
nor U16486 (N_16486,N_16051,N_16076);
and U16487 (N_16487,N_15788,N_15956);
xnor U16488 (N_16488,N_16232,N_15626);
nor U16489 (N_16489,N_16131,N_15659);
and U16490 (N_16490,N_16222,N_15811);
and U16491 (N_16491,N_15944,N_16063);
nor U16492 (N_16492,N_16093,N_16109);
and U16493 (N_16493,N_15948,N_16137);
nor U16494 (N_16494,N_16079,N_15738);
nor U16495 (N_16495,N_15733,N_15705);
or U16496 (N_16496,N_15699,N_15941);
nand U16497 (N_16497,N_16035,N_15802);
xor U16498 (N_16498,N_16188,N_15717);
nor U16499 (N_16499,N_16218,N_16139);
and U16500 (N_16500,N_15961,N_15746);
and U16501 (N_16501,N_15965,N_15840);
nor U16502 (N_16502,N_16134,N_15839);
xnor U16503 (N_16503,N_15742,N_15662);
and U16504 (N_16504,N_16033,N_15665);
nand U16505 (N_16505,N_16236,N_15953);
and U16506 (N_16506,N_16059,N_16055);
nor U16507 (N_16507,N_15671,N_15946);
nor U16508 (N_16508,N_15936,N_15797);
xnor U16509 (N_16509,N_15647,N_15824);
or U16510 (N_16510,N_15754,N_16075);
and U16511 (N_16511,N_15701,N_15710);
and U16512 (N_16512,N_15669,N_16098);
and U16513 (N_16513,N_15731,N_15750);
nor U16514 (N_16514,N_15747,N_16194);
nand U16515 (N_16515,N_16064,N_16092);
nand U16516 (N_16516,N_16245,N_16205);
nand U16517 (N_16517,N_15778,N_15970);
nor U16518 (N_16518,N_15743,N_15921);
xor U16519 (N_16519,N_15890,N_16083);
and U16520 (N_16520,N_16116,N_16029);
and U16521 (N_16521,N_15818,N_16184);
nand U16522 (N_16522,N_16159,N_16004);
nand U16523 (N_16523,N_16243,N_16027);
xor U16524 (N_16524,N_16179,N_15676);
nor U16525 (N_16525,N_16058,N_15640);
nor U16526 (N_16526,N_15794,N_15711);
nor U16527 (N_16527,N_16247,N_16189);
or U16528 (N_16528,N_15644,N_15795);
xnor U16529 (N_16529,N_16105,N_16069);
and U16530 (N_16530,N_16040,N_15680);
or U16531 (N_16531,N_16017,N_15851);
xnor U16532 (N_16532,N_15726,N_16015);
nand U16533 (N_16533,N_16163,N_16151);
nor U16534 (N_16534,N_16114,N_15654);
nor U16535 (N_16535,N_16206,N_15765);
or U16536 (N_16536,N_15820,N_15913);
or U16537 (N_16537,N_15882,N_15789);
xnor U16538 (N_16538,N_16023,N_15814);
nand U16539 (N_16539,N_15878,N_15752);
nor U16540 (N_16540,N_15912,N_15922);
and U16541 (N_16541,N_15962,N_15871);
or U16542 (N_16542,N_15952,N_15700);
nor U16543 (N_16543,N_15837,N_16122);
nor U16544 (N_16544,N_16072,N_15679);
nor U16545 (N_16545,N_15966,N_15911);
and U16546 (N_16546,N_16057,N_15771);
nand U16547 (N_16547,N_15959,N_16225);
or U16548 (N_16548,N_15984,N_16014);
nor U16549 (N_16549,N_16120,N_16228);
nor U16550 (N_16550,N_15945,N_16198);
nor U16551 (N_16551,N_15718,N_15940);
nand U16552 (N_16552,N_16127,N_15924);
xor U16553 (N_16553,N_15931,N_16103);
and U16554 (N_16554,N_15628,N_16125);
and U16555 (N_16555,N_16181,N_15696);
or U16556 (N_16556,N_15772,N_15875);
xor U16557 (N_16557,N_15971,N_15863);
and U16558 (N_16558,N_16020,N_15866);
or U16559 (N_16559,N_16061,N_15791);
and U16560 (N_16560,N_15997,N_15929);
and U16561 (N_16561,N_16110,N_15798);
nand U16562 (N_16562,N_16019,N_15695);
nor U16563 (N_16563,N_16087,N_15963);
and U16564 (N_16564,N_15817,N_15645);
and U16565 (N_16565,N_15631,N_16036);
and U16566 (N_16566,N_15837,N_16013);
nand U16567 (N_16567,N_15820,N_16170);
nor U16568 (N_16568,N_15958,N_15780);
nand U16569 (N_16569,N_16137,N_15861);
nand U16570 (N_16570,N_16186,N_16231);
and U16571 (N_16571,N_15654,N_16016);
or U16572 (N_16572,N_16040,N_16164);
or U16573 (N_16573,N_16156,N_15782);
nand U16574 (N_16574,N_15961,N_15726);
or U16575 (N_16575,N_15886,N_16241);
nand U16576 (N_16576,N_16075,N_15627);
nor U16577 (N_16577,N_16068,N_16077);
or U16578 (N_16578,N_15987,N_15652);
and U16579 (N_16579,N_15883,N_15993);
nor U16580 (N_16580,N_15862,N_16199);
nand U16581 (N_16581,N_16054,N_16139);
and U16582 (N_16582,N_15938,N_15728);
and U16583 (N_16583,N_16021,N_15988);
nor U16584 (N_16584,N_16100,N_15701);
and U16585 (N_16585,N_16061,N_16012);
or U16586 (N_16586,N_15711,N_16090);
nand U16587 (N_16587,N_15643,N_15999);
xnor U16588 (N_16588,N_16201,N_16127);
nand U16589 (N_16589,N_15693,N_16116);
nand U16590 (N_16590,N_15652,N_15835);
nor U16591 (N_16591,N_16089,N_15969);
or U16592 (N_16592,N_15940,N_15909);
or U16593 (N_16593,N_15912,N_16214);
or U16594 (N_16594,N_16024,N_16231);
nand U16595 (N_16595,N_16082,N_16095);
and U16596 (N_16596,N_16081,N_15855);
nand U16597 (N_16597,N_15749,N_15662);
xnor U16598 (N_16598,N_16118,N_15926);
nor U16599 (N_16599,N_15989,N_15693);
nand U16600 (N_16600,N_15747,N_16118);
nand U16601 (N_16601,N_16199,N_16191);
nor U16602 (N_16602,N_16011,N_15999);
or U16603 (N_16603,N_15863,N_15648);
or U16604 (N_16604,N_15930,N_16016);
or U16605 (N_16605,N_16037,N_15725);
or U16606 (N_16606,N_15946,N_15641);
nor U16607 (N_16607,N_16115,N_16049);
nand U16608 (N_16608,N_15739,N_15861);
and U16609 (N_16609,N_15653,N_15990);
and U16610 (N_16610,N_15801,N_15786);
nand U16611 (N_16611,N_15763,N_15709);
nor U16612 (N_16612,N_16074,N_15762);
nand U16613 (N_16613,N_16238,N_15828);
nor U16614 (N_16614,N_16041,N_15899);
and U16615 (N_16615,N_15937,N_15803);
and U16616 (N_16616,N_15767,N_15693);
nor U16617 (N_16617,N_15880,N_16242);
and U16618 (N_16618,N_16087,N_15731);
nand U16619 (N_16619,N_16197,N_15852);
or U16620 (N_16620,N_15878,N_16195);
and U16621 (N_16621,N_16223,N_15856);
or U16622 (N_16622,N_16215,N_15712);
nor U16623 (N_16623,N_15880,N_15670);
or U16624 (N_16624,N_16048,N_15743);
nand U16625 (N_16625,N_16217,N_15651);
nand U16626 (N_16626,N_15665,N_15995);
nor U16627 (N_16627,N_15877,N_15863);
nand U16628 (N_16628,N_15811,N_15915);
nand U16629 (N_16629,N_15934,N_16050);
nand U16630 (N_16630,N_15934,N_16084);
and U16631 (N_16631,N_15674,N_16230);
nor U16632 (N_16632,N_16219,N_15872);
nand U16633 (N_16633,N_15722,N_15749);
and U16634 (N_16634,N_15711,N_15716);
xor U16635 (N_16635,N_15790,N_15763);
nand U16636 (N_16636,N_15945,N_15853);
nor U16637 (N_16637,N_16026,N_15635);
nor U16638 (N_16638,N_16020,N_15976);
nand U16639 (N_16639,N_16083,N_15938);
nor U16640 (N_16640,N_15806,N_15911);
or U16641 (N_16641,N_15747,N_15974);
and U16642 (N_16642,N_15857,N_16053);
and U16643 (N_16643,N_16154,N_16045);
and U16644 (N_16644,N_15676,N_15827);
xnor U16645 (N_16645,N_16070,N_15982);
and U16646 (N_16646,N_15734,N_15897);
nand U16647 (N_16647,N_16057,N_16135);
nand U16648 (N_16648,N_16207,N_16126);
nor U16649 (N_16649,N_15633,N_16017);
or U16650 (N_16650,N_16199,N_15671);
nand U16651 (N_16651,N_16209,N_16222);
nand U16652 (N_16652,N_15819,N_15860);
nand U16653 (N_16653,N_15865,N_15889);
and U16654 (N_16654,N_15929,N_16054);
nand U16655 (N_16655,N_15662,N_16143);
and U16656 (N_16656,N_15821,N_16214);
or U16657 (N_16657,N_16149,N_15818);
xnor U16658 (N_16658,N_15960,N_16204);
or U16659 (N_16659,N_15830,N_15695);
and U16660 (N_16660,N_15652,N_16171);
nor U16661 (N_16661,N_15686,N_15919);
or U16662 (N_16662,N_16028,N_15646);
and U16663 (N_16663,N_15717,N_15716);
and U16664 (N_16664,N_15760,N_15820);
and U16665 (N_16665,N_15854,N_16177);
or U16666 (N_16666,N_16025,N_15761);
nand U16667 (N_16667,N_15738,N_15972);
nor U16668 (N_16668,N_15640,N_16082);
or U16669 (N_16669,N_16065,N_15666);
nand U16670 (N_16670,N_16137,N_15758);
nor U16671 (N_16671,N_15757,N_15734);
nor U16672 (N_16672,N_16113,N_15968);
or U16673 (N_16673,N_15769,N_15647);
or U16674 (N_16674,N_15636,N_16105);
nor U16675 (N_16675,N_16097,N_15915);
nor U16676 (N_16676,N_16188,N_16043);
nand U16677 (N_16677,N_16192,N_15730);
nor U16678 (N_16678,N_15913,N_16097);
nor U16679 (N_16679,N_16174,N_16249);
nand U16680 (N_16680,N_16042,N_16101);
or U16681 (N_16681,N_16217,N_15964);
nand U16682 (N_16682,N_15837,N_15789);
and U16683 (N_16683,N_16137,N_16087);
nand U16684 (N_16684,N_16195,N_15963);
nand U16685 (N_16685,N_15832,N_15930);
and U16686 (N_16686,N_15789,N_15872);
nor U16687 (N_16687,N_16089,N_15735);
nand U16688 (N_16688,N_15873,N_15823);
or U16689 (N_16689,N_16186,N_15811);
xnor U16690 (N_16690,N_16108,N_15794);
nor U16691 (N_16691,N_15857,N_15881);
and U16692 (N_16692,N_15784,N_15854);
nor U16693 (N_16693,N_16135,N_15971);
nor U16694 (N_16694,N_16173,N_16039);
or U16695 (N_16695,N_15947,N_16167);
and U16696 (N_16696,N_16216,N_15954);
or U16697 (N_16697,N_15994,N_15973);
xnor U16698 (N_16698,N_15635,N_15895);
and U16699 (N_16699,N_15973,N_15862);
and U16700 (N_16700,N_15708,N_15890);
or U16701 (N_16701,N_15779,N_16175);
or U16702 (N_16702,N_16167,N_16028);
xnor U16703 (N_16703,N_16082,N_15670);
nand U16704 (N_16704,N_15853,N_16195);
nand U16705 (N_16705,N_15994,N_16099);
xnor U16706 (N_16706,N_15876,N_15794);
nand U16707 (N_16707,N_15831,N_15933);
nand U16708 (N_16708,N_15815,N_16197);
nand U16709 (N_16709,N_15876,N_15761);
and U16710 (N_16710,N_15705,N_15744);
or U16711 (N_16711,N_15947,N_16125);
nor U16712 (N_16712,N_16033,N_15633);
nand U16713 (N_16713,N_15966,N_15906);
or U16714 (N_16714,N_16150,N_15902);
or U16715 (N_16715,N_15658,N_15843);
or U16716 (N_16716,N_16187,N_16226);
nand U16717 (N_16717,N_15767,N_16065);
and U16718 (N_16718,N_15775,N_16131);
nor U16719 (N_16719,N_15855,N_16215);
or U16720 (N_16720,N_16219,N_16136);
nor U16721 (N_16721,N_15699,N_15944);
nand U16722 (N_16722,N_16181,N_15993);
nand U16723 (N_16723,N_16065,N_15706);
nor U16724 (N_16724,N_15778,N_15934);
nand U16725 (N_16725,N_15722,N_15664);
or U16726 (N_16726,N_15734,N_15694);
nor U16727 (N_16727,N_15743,N_16052);
and U16728 (N_16728,N_16153,N_16030);
nor U16729 (N_16729,N_15943,N_15810);
nand U16730 (N_16730,N_16097,N_16104);
nor U16731 (N_16731,N_16031,N_15637);
or U16732 (N_16732,N_16094,N_15752);
or U16733 (N_16733,N_16004,N_16207);
or U16734 (N_16734,N_16236,N_15940);
and U16735 (N_16735,N_15930,N_16006);
or U16736 (N_16736,N_15796,N_16046);
and U16737 (N_16737,N_16100,N_15734);
nand U16738 (N_16738,N_15665,N_15795);
and U16739 (N_16739,N_16024,N_15959);
or U16740 (N_16740,N_16231,N_15965);
and U16741 (N_16741,N_15912,N_15885);
or U16742 (N_16742,N_15701,N_15881);
and U16743 (N_16743,N_15673,N_15675);
nor U16744 (N_16744,N_15706,N_15806);
xor U16745 (N_16745,N_15778,N_15627);
nand U16746 (N_16746,N_15977,N_15657);
nand U16747 (N_16747,N_16012,N_15664);
xor U16748 (N_16748,N_15678,N_16008);
nor U16749 (N_16749,N_15939,N_16161);
xnor U16750 (N_16750,N_15774,N_15836);
and U16751 (N_16751,N_15638,N_16056);
or U16752 (N_16752,N_15971,N_15761);
nand U16753 (N_16753,N_16205,N_16123);
nand U16754 (N_16754,N_16193,N_15655);
and U16755 (N_16755,N_16164,N_15758);
xor U16756 (N_16756,N_15950,N_16227);
nor U16757 (N_16757,N_16181,N_15739);
or U16758 (N_16758,N_16094,N_16114);
or U16759 (N_16759,N_15671,N_15886);
and U16760 (N_16760,N_15868,N_15652);
or U16761 (N_16761,N_15711,N_15966);
nand U16762 (N_16762,N_15824,N_16170);
nor U16763 (N_16763,N_16165,N_16137);
nor U16764 (N_16764,N_15839,N_16076);
and U16765 (N_16765,N_15897,N_15735);
nor U16766 (N_16766,N_15731,N_15843);
and U16767 (N_16767,N_15698,N_15842);
nand U16768 (N_16768,N_16021,N_15780);
nor U16769 (N_16769,N_16074,N_15679);
and U16770 (N_16770,N_16243,N_15690);
nor U16771 (N_16771,N_15932,N_15965);
and U16772 (N_16772,N_15798,N_15914);
nor U16773 (N_16773,N_16052,N_16131);
nor U16774 (N_16774,N_15655,N_15930);
nor U16775 (N_16775,N_15644,N_15730);
nor U16776 (N_16776,N_16044,N_15887);
nand U16777 (N_16777,N_15975,N_16225);
or U16778 (N_16778,N_15954,N_16112);
or U16779 (N_16779,N_16244,N_15736);
xor U16780 (N_16780,N_16232,N_15777);
and U16781 (N_16781,N_15943,N_15907);
xor U16782 (N_16782,N_16101,N_15994);
nor U16783 (N_16783,N_16106,N_16092);
nand U16784 (N_16784,N_16024,N_16033);
nor U16785 (N_16785,N_16167,N_15694);
xnor U16786 (N_16786,N_16183,N_16191);
and U16787 (N_16787,N_15923,N_15946);
nand U16788 (N_16788,N_16126,N_15824);
xor U16789 (N_16789,N_15741,N_15909);
nand U16790 (N_16790,N_15690,N_16118);
and U16791 (N_16791,N_15883,N_15728);
or U16792 (N_16792,N_15935,N_16150);
nor U16793 (N_16793,N_16080,N_15682);
nand U16794 (N_16794,N_15833,N_15668);
or U16795 (N_16795,N_15671,N_15717);
nor U16796 (N_16796,N_16177,N_16201);
xnor U16797 (N_16797,N_16106,N_16000);
nor U16798 (N_16798,N_16187,N_15949);
nor U16799 (N_16799,N_16182,N_15689);
or U16800 (N_16800,N_15783,N_16200);
nand U16801 (N_16801,N_15870,N_15768);
nand U16802 (N_16802,N_15818,N_16218);
xor U16803 (N_16803,N_15824,N_15668);
nand U16804 (N_16804,N_15750,N_15721);
or U16805 (N_16805,N_15625,N_16087);
nand U16806 (N_16806,N_15844,N_16102);
and U16807 (N_16807,N_15954,N_15850);
xor U16808 (N_16808,N_16162,N_15811);
xor U16809 (N_16809,N_15693,N_16076);
nand U16810 (N_16810,N_15877,N_15999);
nor U16811 (N_16811,N_15638,N_15835);
or U16812 (N_16812,N_15880,N_15772);
nand U16813 (N_16813,N_15812,N_16060);
or U16814 (N_16814,N_15917,N_15862);
nor U16815 (N_16815,N_15708,N_16240);
and U16816 (N_16816,N_15681,N_15912);
nor U16817 (N_16817,N_15722,N_15629);
and U16818 (N_16818,N_16046,N_16129);
nor U16819 (N_16819,N_15772,N_15852);
or U16820 (N_16820,N_15679,N_15799);
and U16821 (N_16821,N_15980,N_15865);
and U16822 (N_16822,N_15819,N_15702);
or U16823 (N_16823,N_15658,N_15700);
or U16824 (N_16824,N_16234,N_15778);
xor U16825 (N_16825,N_16216,N_15681);
nand U16826 (N_16826,N_15989,N_15889);
or U16827 (N_16827,N_16087,N_16004);
nand U16828 (N_16828,N_16062,N_16065);
nand U16829 (N_16829,N_16169,N_15996);
nand U16830 (N_16830,N_15986,N_15843);
nor U16831 (N_16831,N_15723,N_15645);
xor U16832 (N_16832,N_16183,N_15646);
nor U16833 (N_16833,N_15903,N_15700);
nor U16834 (N_16834,N_15701,N_15865);
or U16835 (N_16835,N_15910,N_15631);
nand U16836 (N_16836,N_15696,N_15653);
nor U16837 (N_16837,N_15706,N_15666);
or U16838 (N_16838,N_16113,N_15820);
nor U16839 (N_16839,N_15716,N_15817);
and U16840 (N_16840,N_16096,N_16220);
and U16841 (N_16841,N_16172,N_15750);
or U16842 (N_16842,N_15649,N_15658);
and U16843 (N_16843,N_15832,N_15677);
and U16844 (N_16844,N_16129,N_16056);
and U16845 (N_16845,N_15914,N_15950);
and U16846 (N_16846,N_16136,N_15896);
nand U16847 (N_16847,N_15967,N_16098);
or U16848 (N_16848,N_16236,N_15765);
nor U16849 (N_16849,N_16106,N_16014);
or U16850 (N_16850,N_16225,N_15926);
nand U16851 (N_16851,N_16229,N_16125);
xnor U16852 (N_16852,N_15729,N_16121);
nand U16853 (N_16853,N_16156,N_15627);
and U16854 (N_16854,N_15850,N_16183);
nand U16855 (N_16855,N_15669,N_15635);
nor U16856 (N_16856,N_15697,N_15984);
xnor U16857 (N_16857,N_16075,N_15650);
nand U16858 (N_16858,N_15698,N_15646);
and U16859 (N_16859,N_16092,N_16008);
or U16860 (N_16860,N_15976,N_16165);
nor U16861 (N_16861,N_16039,N_15676);
or U16862 (N_16862,N_16194,N_15958);
nand U16863 (N_16863,N_16145,N_16046);
nand U16864 (N_16864,N_15959,N_16053);
nand U16865 (N_16865,N_15973,N_16239);
xnor U16866 (N_16866,N_15906,N_16001);
xor U16867 (N_16867,N_15944,N_16170);
nand U16868 (N_16868,N_15933,N_15967);
nor U16869 (N_16869,N_15825,N_16184);
or U16870 (N_16870,N_15911,N_15848);
nand U16871 (N_16871,N_15872,N_15829);
or U16872 (N_16872,N_15829,N_16176);
and U16873 (N_16873,N_16060,N_15847);
nand U16874 (N_16874,N_16175,N_15837);
xnor U16875 (N_16875,N_16584,N_16841);
and U16876 (N_16876,N_16270,N_16349);
or U16877 (N_16877,N_16641,N_16374);
nand U16878 (N_16878,N_16520,N_16373);
or U16879 (N_16879,N_16649,N_16709);
nor U16880 (N_16880,N_16341,N_16323);
or U16881 (N_16881,N_16747,N_16253);
or U16882 (N_16882,N_16823,N_16330);
nand U16883 (N_16883,N_16770,N_16665);
nor U16884 (N_16884,N_16833,N_16704);
nor U16885 (N_16885,N_16441,N_16369);
or U16886 (N_16886,N_16459,N_16815);
or U16887 (N_16887,N_16456,N_16435);
or U16888 (N_16888,N_16557,N_16596);
or U16889 (N_16889,N_16254,N_16511);
nor U16890 (N_16890,N_16866,N_16480);
nand U16891 (N_16891,N_16411,N_16637);
or U16892 (N_16892,N_16263,N_16422);
nand U16893 (N_16893,N_16793,N_16769);
nand U16894 (N_16894,N_16262,N_16491);
xnor U16895 (N_16895,N_16636,N_16711);
and U16896 (N_16896,N_16790,N_16261);
nor U16897 (N_16897,N_16608,N_16701);
nor U16898 (N_16898,N_16489,N_16756);
and U16899 (N_16899,N_16697,N_16388);
and U16900 (N_16900,N_16648,N_16558);
nor U16901 (N_16901,N_16306,N_16796);
and U16902 (N_16902,N_16541,N_16327);
nor U16903 (N_16903,N_16255,N_16296);
or U16904 (N_16904,N_16300,N_16407);
nor U16905 (N_16905,N_16612,N_16809);
nand U16906 (N_16906,N_16700,N_16761);
or U16907 (N_16907,N_16408,N_16817);
nand U16908 (N_16908,N_16366,N_16475);
and U16909 (N_16909,N_16370,N_16376);
nor U16910 (N_16910,N_16763,N_16331);
nor U16911 (N_16911,N_16774,N_16414);
nor U16912 (N_16912,N_16400,N_16324);
or U16913 (N_16913,N_16500,N_16871);
nor U16914 (N_16914,N_16614,N_16333);
nor U16915 (N_16915,N_16867,N_16791);
nand U16916 (N_16916,N_16322,N_16404);
nor U16917 (N_16917,N_16444,N_16730);
or U16918 (N_16918,N_16865,N_16736);
nor U16919 (N_16919,N_16348,N_16452);
nor U16920 (N_16920,N_16372,N_16529);
and U16921 (N_16921,N_16788,N_16874);
nand U16922 (N_16922,N_16543,N_16757);
nor U16923 (N_16923,N_16492,N_16299);
or U16924 (N_16924,N_16470,N_16304);
nand U16925 (N_16925,N_16783,N_16628);
nand U16926 (N_16926,N_16506,N_16463);
or U16927 (N_16927,N_16275,N_16749);
or U16928 (N_16928,N_16743,N_16420);
xor U16929 (N_16929,N_16447,N_16576);
nor U16930 (N_16930,N_16250,N_16273);
nor U16931 (N_16931,N_16825,N_16502);
nor U16932 (N_16932,N_16283,N_16691);
nor U16933 (N_16933,N_16504,N_16313);
or U16934 (N_16934,N_16851,N_16395);
and U16935 (N_16935,N_16803,N_16510);
nor U16936 (N_16936,N_16741,N_16703);
nor U16937 (N_16937,N_16496,N_16610);
nor U16938 (N_16938,N_16339,N_16605);
and U16939 (N_16939,N_16818,N_16325);
or U16940 (N_16940,N_16434,N_16364);
nor U16941 (N_16941,N_16337,N_16617);
or U16942 (N_16942,N_16772,N_16735);
nor U16943 (N_16943,N_16354,N_16282);
and U16944 (N_16944,N_16514,N_16632);
or U16945 (N_16945,N_16314,N_16352);
and U16946 (N_16946,N_16827,N_16657);
and U16947 (N_16947,N_16271,N_16615);
or U16948 (N_16948,N_16289,N_16269);
xnor U16949 (N_16949,N_16578,N_16454);
and U16950 (N_16950,N_16564,N_16278);
and U16951 (N_16951,N_16288,N_16748);
nor U16952 (N_16952,N_16845,N_16525);
nor U16953 (N_16953,N_16868,N_16347);
nor U16954 (N_16954,N_16277,N_16509);
or U16955 (N_16955,N_16426,N_16534);
nor U16956 (N_16956,N_16490,N_16478);
nand U16957 (N_16957,N_16599,N_16622);
or U16958 (N_16958,N_16837,N_16860);
or U16959 (N_16959,N_16381,N_16401);
nor U16960 (N_16960,N_16448,N_16355);
and U16961 (N_16961,N_16814,N_16428);
nand U16962 (N_16962,N_16762,N_16379);
xor U16963 (N_16963,N_16450,N_16806);
nand U16964 (N_16964,N_16684,N_16621);
nand U16965 (N_16965,N_16471,N_16712);
or U16966 (N_16966,N_16659,N_16503);
nand U16967 (N_16967,N_16579,N_16753);
nor U16968 (N_16968,N_16451,N_16780);
and U16969 (N_16969,N_16591,N_16284);
nand U16970 (N_16970,N_16781,N_16530);
and U16971 (N_16971,N_16731,N_16309);
nor U16972 (N_16972,N_16722,N_16830);
nand U16973 (N_16973,N_16673,N_16638);
nor U16974 (N_16974,N_16732,N_16424);
or U16975 (N_16975,N_16553,N_16350);
and U16976 (N_16976,N_16853,N_16716);
nor U16977 (N_16977,N_16516,N_16662);
xnor U16978 (N_16978,N_16586,N_16702);
nand U16979 (N_16979,N_16755,N_16842);
and U16980 (N_16980,N_16685,N_16816);
nand U16981 (N_16981,N_16760,N_16670);
xnor U16982 (N_16982,N_16678,N_16391);
nor U16983 (N_16983,N_16546,N_16680);
or U16984 (N_16984,N_16519,N_16583);
or U16985 (N_16985,N_16433,N_16455);
or U16986 (N_16986,N_16256,N_16316);
nor U16987 (N_16987,N_16409,N_16291);
nor U16988 (N_16988,N_16522,N_16719);
or U16989 (N_16989,N_16779,N_16695);
nor U16990 (N_16990,N_16494,N_16368);
nand U16991 (N_16991,N_16402,N_16524);
or U16992 (N_16992,N_16764,N_16645);
nor U16993 (N_16993,N_16359,N_16416);
nor U16994 (N_16994,N_16619,N_16329);
nand U16995 (N_16995,N_16826,N_16353);
nand U16996 (N_16996,N_16260,N_16848);
or U16997 (N_16997,N_16595,N_16307);
or U16998 (N_16998,N_16873,N_16436);
xor U16999 (N_16999,N_16340,N_16536);
and U17000 (N_17000,N_16676,N_16824);
or U17001 (N_17001,N_16639,N_16765);
nand U17002 (N_17002,N_16518,N_16412);
and U17003 (N_17003,N_16854,N_16342);
xor U17004 (N_17004,N_16857,N_16752);
or U17005 (N_17005,N_16335,N_16281);
and U17006 (N_17006,N_16446,N_16423);
nand U17007 (N_17007,N_16419,N_16259);
nor U17008 (N_17008,N_16643,N_16499);
or U17009 (N_17009,N_16425,N_16287);
or U17010 (N_17010,N_16336,N_16512);
or U17011 (N_17011,N_16677,N_16603);
or U17012 (N_17012,N_16802,N_16303);
nor U17013 (N_17013,N_16551,N_16718);
nor U17014 (N_17014,N_16733,N_16767);
or U17015 (N_17015,N_16721,N_16737);
nor U17016 (N_17016,N_16526,N_16367);
and U17017 (N_17017,N_16759,N_16686);
and U17018 (N_17018,N_16290,N_16710);
nand U17019 (N_17019,N_16547,N_16357);
nor U17020 (N_17020,N_16656,N_16394);
nor U17021 (N_17021,N_16807,N_16417);
and U17022 (N_17022,N_16723,N_16318);
or U17023 (N_17023,N_16786,N_16298);
nand U17024 (N_17024,N_16870,N_16351);
xor U17025 (N_17025,N_16675,N_16286);
xor U17026 (N_17026,N_16655,N_16646);
and U17027 (N_17027,N_16515,N_16631);
and U17028 (N_17028,N_16540,N_16497);
or U17029 (N_17029,N_16822,N_16594);
or U17030 (N_17030,N_16819,N_16482);
nor U17031 (N_17031,N_16787,N_16474);
nand U17032 (N_17032,N_16627,N_16427);
and U17033 (N_17033,N_16629,N_16485);
or U17034 (N_17034,N_16604,N_16580);
or U17035 (N_17035,N_16738,N_16344);
or U17036 (N_17036,N_16593,N_16460);
nand U17037 (N_17037,N_16384,N_16835);
or U17038 (N_17038,N_16863,N_16794);
nand U17039 (N_17039,N_16831,N_16634);
nor U17040 (N_17040,N_16398,N_16377);
nand U17041 (N_17041,N_16663,N_16795);
nor U17042 (N_17042,N_16708,N_16577);
and U17043 (N_17043,N_16305,N_16727);
or U17044 (N_17044,N_16389,N_16371);
and U17045 (N_17045,N_16467,N_16266);
nor U17046 (N_17046,N_16862,N_16828);
nand U17047 (N_17047,N_16544,N_16539);
nand U17048 (N_17048,N_16751,N_16265);
or U17049 (N_17049,N_16674,N_16799);
nor U17050 (N_17050,N_16633,N_16321);
or U17051 (N_17051,N_16664,N_16714);
and U17052 (N_17052,N_16575,N_16838);
nor U17053 (N_17053,N_16533,N_16295);
or U17054 (N_17054,N_16505,N_16778);
or U17055 (N_17055,N_16517,N_16545);
nand U17056 (N_17056,N_16375,N_16813);
xor U17057 (N_17057,N_16279,N_16561);
xnor U17058 (N_17058,N_16683,N_16562);
nor U17059 (N_17059,N_16776,N_16466);
nor U17060 (N_17060,N_16570,N_16443);
nor U17061 (N_17061,N_16654,N_16742);
and U17062 (N_17062,N_16625,N_16805);
nor U17063 (N_17063,N_16720,N_16672);
xor U17064 (N_17064,N_16481,N_16442);
nand U17065 (N_17065,N_16623,N_16559);
nor U17066 (N_17066,N_16811,N_16264);
nand U17067 (N_17067,N_16521,N_16272);
and U17068 (N_17068,N_16768,N_16725);
or U17069 (N_17069,N_16859,N_16403);
and U17070 (N_17070,N_16439,N_16458);
and U17071 (N_17071,N_16651,N_16315);
nand U17072 (N_17072,N_16461,N_16410);
nand U17073 (N_17073,N_16589,N_16650);
nand U17074 (N_17074,N_16810,N_16782);
xnor U17075 (N_17075,N_16479,N_16687);
or U17076 (N_17076,N_16556,N_16465);
or U17077 (N_17077,N_16592,N_16319);
and U17078 (N_17078,N_16808,N_16574);
and U17079 (N_17079,N_16498,N_16563);
nor U17080 (N_17080,N_16274,N_16869);
or U17081 (N_17081,N_16387,N_16385);
or U17082 (N_17082,N_16724,N_16523);
and U17083 (N_17083,N_16844,N_16413);
nor U17084 (N_17084,N_16600,N_16390);
and U17085 (N_17085,N_16542,N_16280);
and U17086 (N_17086,N_16396,N_16715);
and U17087 (N_17087,N_16847,N_16858);
and U17088 (N_17088,N_16820,N_16658);
xor U17089 (N_17089,N_16483,N_16754);
nor U17090 (N_17090,N_16785,N_16453);
nor U17091 (N_17091,N_16251,N_16493);
and U17092 (N_17092,N_16294,N_16642);
or U17093 (N_17093,N_16438,N_16804);
and U17094 (N_17094,N_16362,N_16484);
nand U17095 (N_17095,N_16569,N_16766);
and U17096 (N_17096,N_16597,N_16365);
nor U17097 (N_17097,N_16849,N_16573);
nand U17098 (N_17098,N_16468,N_16777);
xnor U17099 (N_17099,N_16568,N_16552);
nor U17100 (N_17100,N_16635,N_16801);
or U17101 (N_17101,N_16343,N_16549);
nand U17102 (N_17102,N_16449,N_16445);
nor U17103 (N_17103,N_16571,N_16689);
nand U17104 (N_17104,N_16363,N_16332);
nor U17105 (N_17105,N_16588,N_16268);
and U17106 (N_17106,N_16285,N_16399);
and U17107 (N_17107,N_16688,N_16630);
and U17108 (N_17108,N_16361,N_16378);
xnor U17109 (N_17109,N_16666,N_16829);
nor U17110 (N_17110,N_16430,N_16554);
nor U17111 (N_17111,N_16745,N_16626);
nor U17112 (N_17112,N_16537,N_16528);
nor U17113 (N_17113,N_16538,N_16383);
nand U17114 (N_17114,N_16356,N_16640);
and U17115 (N_17115,N_16258,N_16840);
or U17116 (N_17116,N_16740,N_16616);
and U17117 (N_17117,N_16405,N_16821);
nor U17118 (N_17118,N_16699,N_16611);
and U17119 (N_17119,N_16647,N_16620);
and U17120 (N_17120,N_16836,N_16784);
or U17121 (N_17121,N_16293,N_16346);
or U17122 (N_17122,N_16746,N_16861);
nand U17123 (N_17123,N_16598,N_16706);
or U17124 (N_17124,N_16513,N_16679);
nand U17125 (N_17125,N_16358,N_16415);
or U17126 (N_17126,N_16846,N_16527);
xor U17127 (N_17127,N_16477,N_16582);
xor U17128 (N_17128,N_16850,N_16393);
nand U17129 (N_17129,N_16326,N_16773);
or U17130 (N_17130,N_16276,N_16713);
or U17131 (N_17131,N_16797,N_16566);
and U17132 (N_17132,N_16567,N_16690);
or U17133 (N_17133,N_16328,N_16345);
xnor U17134 (N_17134,N_16535,N_16440);
nor U17135 (N_17135,N_16800,N_16590);
and U17136 (N_17136,N_16437,N_16682);
or U17137 (N_17137,N_16602,N_16812);
and U17138 (N_17138,N_16421,N_16855);
nand U17139 (N_17139,N_16508,N_16667);
and U17140 (N_17140,N_16717,N_16798);
nor U17141 (N_17141,N_16301,N_16864);
nor U17142 (N_17142,N_16694,N_16432);
nor U17143 (N_17143,N_16312,N_16693);
or U17144 (N_17144,N_16302,N_16473);
nor U17145 (N_17145,N_16607,N_16681);
nand U17146 (N_17146,N_16429,N_16572);
or U17147 (N_17147,N_16320,N_16472);
or U17148 (N_17148,N_16486,N_16555);
nor U17149 (N_17149,N_16476,N_16792);
nand U17150 (N_17150,N_16671,N_16652);
nor U17151 (N_17151,N_16668,N_16488);
and U17152 (N_17152,N_16310,N_16734);
and U17153 (N_17153,N_16338,N_16257);
and U17154 (N_17154,N_16392,N_16660);
and U17155 (N_17155,N_16669,N_16744);
and U17156 (N_17156,N_16661,N_16462);
nor U17157 (N_17157,N_16618,N_16334);
nor U17158 (N_17158,N_16750,N_16729);
nand U17159 (N_17159,N_16609,N_16728);
nor U17160 (N_17160,N_16501,N_16771);
xnor U17161 (N_17161,N_16856,N_16581);
and U17162 (N_17162,N_16606,N_16531);
nand U17163 (N_17163,N_16252,N_16507);
and U17164 (N_17164,N_16267,N_16560);
nand U17165 (N_17165,N_16431,N_16565);
nand U17166 (N_17166,N_16308,N_16380);
and U17167 (N_17167,N_16726,N_16601);
and U17168 (N_17168,N_16532,N_16292);
and U17169 (N_17169,N_16843,N_16397);
or U17170 (N_17170,N_16775,N_16418);
or U17171 (N_17171,N_16758,N_16382);
nand U17172 (N_17172,N_16739,N_16872);
nor U17173 (N_17173,N_16832,N_16624);
and U17174 (N_17174,N_16692,N_16696);
nor U17175 (N_17175,N_16548,N_16587);
nor U17176 (N_17176,N_16487,N_16550);
and U17177 (N_17177,N_16705,N_16317);
and U17178 (N_17178,N_16653,N_16406);
nand U17179 (N_17179,N_16852,N_16707);
and U17180 (N_17180,N_16834,N_16469);
and U17181 (N_17181,N_16457,N_16297);
and U17182 (N_17182,N_16360,N_16464);
or U17183 (N_17183,N_16613,N_16386);
nor U17184 (N_17184,N_16495,N_16311);
nor U17185 (N_17185,N_16644,N_16789);
and U17186 (N_17186,N_16839,N_16585);
nand U17187 (N_17187,N_16698,N_16691);
xor U17188 (N_17188,N_16258,N_16568);
nand U17189 (N_17189,N_16683,N_16723);
xor U17190 (N_17190,N_16317,N_16292);
or U17191 (N_17191,N_16416,N_16406);
nor U17192 (N_17192,N_16728,N_16604);
nor U17193 (N_17193,N_16353,N_16380);
xor U17194 (N_17194,N_16767,N_16622);
nor U17195 (N_17195,N_16392,N_16356);
or U17196 (N_17196,N_16557,N_16266);
nor U17197 (N_17197,N_16761,N_16443);
nand U17198 (N_17198,N_16793,N_16489);
and U17199 (N_17199,N_16543,N_16333);
and U17200 (N_17200,N_16309,N_16848);
nand U17201 (N_17201,N_16265,N_16789);
and U17202 (N_17202,N_16289,N_16272);
or U17203 (N_17203,N_16573,N_16506);
and U17204 (N_17204,N_16304,N_16303);
and U17205 (N_17205,N_16642,N_16755);
or U17206 (N_17206,N_16574,N_16719);
and U17207 (N_17207,N_16377,N_16607);
nor U17208 (N_17208,N_16561,N_16640);
or U17209 (N_17209,N_16288,N_16662);
and U17210 (N_17210,N_16259,N_16567);
and U17211 (N_17211,N_16356,N_16258);
nor U17212 (N_17212,N_16513,N_16817);
and U17213 (N_17213,N_16581,N_16738);
nor U17214 (N_17214,N_16576,N_16284);
or U17215 (N_17215,N_16558,N_16512);
nand U17216 (N_17216,N_16726,N_16816);
xnor U17217 (N_17217,N_16835,N_16360);
and U17218 (N_17218,N_16546,N_16335);
and U17219 (N_17219,N_16508,N_16429);
or U17220 (N_17220,N_16428,N_16589);
nor U17221 (N_17221,N_16645,N_16449);
and U17222 (N_17222,N_16351,N_16333);
nand U17223 (N_17223,N_16707,N_16277);
nor U17224 (N_17224,N_16821,N_16732);
or U17225 (N_17225,N_16728,N_16306);
or U17226 (N_17226,N_16362,N_16383);
or U17227 (N_17227,N_16559,N_16849);
and U17228 (N_17228,N_16378,N_16661);
nand U17229 (N_17229,N_16762,N_16698);
nor U17230 (N_17230,N_16656,N_16787);
and U17231 (N_17231,N_16487,N_16533);
or U17232 (N_17232,N_16486,N_16341);
or U17233 (N_17233,N_16701,N_16780);
nor U17234 (N_17234,N_16549,N_16424);
and U17235 (N_17235,N_16570,N_16465);
nand U17236 (N_17236,N_16743,N_16298);
nand U17237 (N_17237,N_16377,N_16628);
nor U17238 (N_17238,N_16671,N_16684);
nor U17239 (N_17239,N_16842,N_16400);
and U17240 (N_17240,N_16426,N_16463);
nor U17241 (N_17241,N_16814,N_16688);
nor U17242 (N_17242,N_16718,N_16327);
nand U17243 (N_17243,N_16499,N_16874);
or U17244 (N_17244,N_16874,N_16340);
nand U17245 (N_17245,N_16672,N_16485);
nand U17246 (N_17246,N_16761,N_16413);
xnor U17247 (N_17247,N_16262,N_16484);
nor U17248 (N_17248,N_16308,N_16624);
and U17249 (N_17249,N_16304,N_16822);
or U17250 (N_17250,N_16678,N_16540);
nand U17251 (N_17251,N_16335,N_16524);
or U17252 (N_17252,N_16665,N_16463);
nand U17253 (N_17253,N_16532,N_16481);
or U17254 (N_17254,N_16844,N_16799);
nor U17255 (N_17255,N_16750,N_16400);
nor U17256 (N_17256,N_16729,N_16466);
or U17257 (N_17257,N_16595,N_16605);
nor U17258 (N_17258,N_16545,N_16455);
xnor U17259 (N_17259,N_16307,N_16717);
or U17260 (N_17260,N_16517,N_16571);
nand U17261 (N_17261,N_16575,N_16268);
nor U17262 (N_17262,N_16591,N_16254);
and U17263 (N_17263,N_16618,N_16487);
nand U17264 (N_17264,N_16784,N_16354);
nor U17265 (N_17265,N_16771,N_16292);
nor U17266 (N_17266,N_16630,N_16342);
nor U17267 (N_17267,N_16774,N_16575);
and U17268 (N_17268,N_16763,N_16282);
or U17269 (N_17269,N_16382,N_16265);
nand U17270 (N_17270,N_16780,N_16481);
and U17271 (N_17271,N_16485,N_16846);
nor U17272 (N_17272,N_16463,N_16858);
nor U17273 (N_17273,N_16363,N_16645);
or U17274 (N_17274,N_16776,N_16542);
xor U17275 (N_17275,N_16609,N_16766);
or U17276 (N_17276,N_16467,N_16412);
xnor U17277 (N_17277,N_16526,N_16348);
nor U17278 (N_17278,N_16369,N_16860);
or U17279 (N_17279,N_16262,N_16429);
and U17280 (N_17280,N_16749,N_16555);
nand U17281 (N_17281,N_16258,N_16502);
xor U17282 (N_17282,N_16838,N_16786);
and U17283 (N_17283,N_16799,N_16497);
and U17284 (N_17284,N_16559,N_16571);
nand U17285 (N_17285,N_16760,N_16616);
and U17286 (N_17286,N_16271,N_16592);
nand U17287 (N_17287,N_16617,N_16640);
or U17288 (N_17288,N_16498,N_16382);
or U17289 (N_17289,N_16300,N_16413);
nand U17290 (N_17290,N_16588,N_16723);
xnor U17291 (N_17291,N_16302,N_16603);
and U17292 (N_17292,N_16429,N_16828);
and U17293 (N_17293,N_16444,N_16696);
nand U17294 (N_17294,N_16661,N_16763);
or U17295 (N_17295,N_16708,N_16697);
nand U17296 (N_17296,N_16708,N_16650);
or U17297 (N_17297,N_16864,N_16668);
nor U17298 (N_17298,N_16586,N_16476);
nand U17299 (N_17299,N_16473,N_16760);
nand U17300 (N_17300,N_16527,N_16659);
or U17301 (N_17301,N_16521,N_16464);
or U17302 (N_17302,N_16780,N_16721);
xnor U17303 (N_17303,N_16390,N_16339);
or U17304 (N_17304,N_16828,N_16340);
xnor U17305 (N_17305,N_16762,N_16385);
nand U17306 (N_17306,N_16522,N_16528);
nand U17307 (N_17307,N_16345,N_16489);
nand U17308 (N_17308,N_16725,N_16304);
and U17309 (N_17309,N_16365,N_16732);
or U17310 (N_17310,N_16592,N_16309);
nor U17311 (N_17311,N_16300,N_16614);
nand U17312 (N_17312,N_16711,N_16317);
nor U17313 (N_17313,N_16379,N_16536);
nand U17314 (N_17314,N_16625,N_16694);
nand U17315 (N_17315,N_16571,N_16748);
nand U17316 (N_17316,N_16381,N_16531);
nor U17317 (N_17317,N_16741,N_16721);
nand U17318 (N_17318,N_16557,N_16722);
nand U17319 (N_17319,N_16808,N_16765);
nand U17320 (N_17320,N_16297,N_16713);
and U17321 (N_17321,N_16469,N_16338);
nor U17322 (N_17322,N_16257,N_16424);
xor U17323 (N_17323,N_16334,N_16801);
and U17324 (N_17324,N_16825,N_16657);
nor U17325 (N_17325,N_16295,N_16686);
or U17326 (N_17326,N_16338,N_16663);
and U17327 (N_17327,N_16769,N_16389);
nand U17328 (N_17328,N_16493,N_16365);
nor U17329 (N_17329,N_16682,N_16612);
nand U17330 (N_17330,N_16451,N_16680);
and U17331 (N_17331,N_16570,N_16368);
nor U17332 (N_17332,N_16371,N_16295);
nand U17333 (N_17333,N_16555,N_16661);
or U17334 (N_17334,N_16799,N_16456);
and U17335 (N_17335,N_16415,N_16694);
nor U17336 (N_17336,N_16430,N_16464);
and U17337 (N_17337,N_16288,N_16772);
or U17338 (N_17338,N_16758,N_16380);
or U17339 (N_17339,N_16478,N_16291);
or U17340 (N_17340,N_16860,N_16773);
or U17341 (N_17341,N_16552,N_16851);
or U17342 (N_17342,N_16822,N_16526);
and U17343 (N_17343,N_16391,N_16538);
nand U17344 (N_17344,N_16342,N_16681);
or U17345 (N_17345,N_16585,N_16469);
nand U17346 (N_17346,N_16832,N_16775);
nor U17347 (N_17347,N_16551,N_16539);
xor U17348 (N_17348,N_16840,N_16283);
and U17349 (N_17349,N_16453,N_16726);
or U17350 (N_17350,N_16428,N_16621);
or U17351 (N_17351,N_16428,N_16333);
and U17352 (N_17352,N_16379,N_16501);
nor U17353 (N_17353,N_16276,N_16868);
and U17354 (N_17354,N_16370,N_16407);
nor U17355 (N_17355,N_16431,N_16350);
and U17356 (N_17356,N_16456,N_16399);
nand U17357 (N_17357,N_16810,N_16353);
and U17358 (N_17358,N_16313,N_16416);
nand U17359 (N_17359,N_16842,N_16658);
nor U17360 (N_17360,N_16413,N_16739);
or U17361 (N_17361,N_16522,N_16290);
xor U17362 (N_17362,N_16856,N_16543);
nor U17363 (N_17363,N_16352,N_16748);
nand U17364 (N_17364,N_16351,N_16869);
xnor U17365 (N_17365,N_16502,N_16327);
and U17366 (N_17366,N_16511,N_16735);
and U17367 (N_17367,N_16320,N_16851);
nand U17368 (N_17368,N_16571,N_16514);
or U17369 (N_17369,N_16390,N_16630);
or U17370 (N_17370,N_16365,N_16794);
and U17371 (N_17371,N_16579,N_16826);
nand U17372 (N_17372,N_16465,N_16730);
or U17373 (N_17373,N_16686,N_16370);
nand U17374 (N_17374,N_16766,N_16460);
or U17375 (N_17375,N_16277,N_16478);
nor U17376 (N_17376,N_16554,N_16583);
nor U17377 (N_17377,N_16573,N_16660);
nor U17378 (N_17378,N_16579,N_16385);
or U17379 (N_17379,N_16452,N_16331);
nor U17380 (N_17380,N_16465,N_16663);
or U17381 (N_17381,N_16752,N_16263);
xnor U17382 (N_17382,N_16304,N_16735);
or U17383 (N_17383,N_16316,N_16505);
and U17384 (N_17384,N_16360,N_16506);
nand U17385 (N_17385,N_16565,N_16552);
or U17386 (N_17386,N_16272,N_16684);
and U17387 (N_17387,N_16493,N_16865);
nand U17388 (N_17388,N_16419,N_16573);
nor U17389 (N_17389,N_16321,N_16599);
nor U17390 (N_17390,N_16558,N_16689);
nand U17391 (N_17391,N_16408,N_16585);
nand U17392 (N_17392,N_16421,N_16763);
nand U17393 (N_17393,N_16460,N_16289);
and U17394 (N_17394,N_16493,N_16492);
or U17395 (N_17395,N_16864,N_16822);
nand U17396 (N_17396,N_16324,N_16389);
and U17397 (N_17397,N_16683,N_16494);
and U17398 (N_17398,N_16530,N_16665);
nor U17399 (N_17399,N_16828,N_16651);
nand U17400 (N_17400,N_16305,N_16766);
or U17401 (N_17401,N_16545,N_16512);
and U17402 (N_17402,N_16811,N_16468);
and U17403 (N_17403,N_16868,N_16656);
xor U17404 (N_17404,N_16771,N_16475);
nand U17405 (N_17405,N_16672,N_16779);
nor U17406 (N_17406,N_16466,N_16586);
xor U17407 (N_17407,N_16264,N_16311);
nor U17408 (N_17408,N_16675,N_16679);
xnor U17409 (N_17409,N_16355,N_16534);
xnor U17410 (N_17410,N_16250,N_16564);
or U17411 (N_17411,N_16765,N_16786);
and U17412 (N_17412,N_16380,N_16535);
nand U17413 (N_17413,N_16780,N_16532);
nand U17414 (N_17414,N_16493,N_16518);
xnor U17415 (N_17415,N_16856,N_16669);
nand U17416 (N_17416,N_16756,N_16513);
nor U17417 (N_17417,N_16340,N_16795);
xnor U17418 (N_17418,N_16563,N_16710);
nor U17419 (N_17419,N_16581,N_16673);
or U17420 (N_17420,N_16833,N_16398);
nand U17421 (N_17421,N_16834,N_16400);
nor U17422 (N_17422,N_16533,N_16747);
or U17423 (N_17423,N_16598,N_16596);
nor U17424 (N_17424,N_16356,N_16490);
xor U17425 (N_17425,N_16328,N_16841);
or U17426 (N_17426,N_16771,N_16355);
and U17427 (N_17427,N_16786,N_16354);
nor U17428 (N_17428,N_16695,N_16413);
xnor U17429 (N_17429,N_16371,N_16570);
or U17430 (N_17430,N_16587,N_16416);
or U17431 (N_17431,N_16869,N_16811);
or U17432 (N_17432,N_16313,N_16303);
nor U17433 (N_17433,N_16264,N_16401);
nor U17434 (N_17434,N_16469,N_16437);
and U17435 (N_17435,N_16518,N_16439);
nand U17436 (N_17436,N_16281,N_16422);
and U17437 (N_17437,N_16829,N_16504);
and U17438 (N_17438,N_16438,N_16687);
nor U17439 (N_17439,N_16833,N_16469);
or U17440 (N_17440,N_16352,N_16412);
nor U17441 (N_17441,N_16313,N_16508);
nor U17442 (N_17442,N_16491,N_16438);
nand U17443 (N_17443,N_16257,N_16382);
xor U17444 (N_17444,N_16535,N_16297);
nor U17445 (N_17445,N_16570,N_16822);
nor U17446 (N_17446,N_16732,N_16421);
or U17447 (N_17447,N_16707,N_16528);
nor U17448 (N_17448,N_16674,N_16276);
nand U17449 (N_17449,N_16415,N_16863);
and U17450 (N_17450,N_16742,N_16724);
xor U17451 (N_17451,N_16356,N_16839);
nand U17452 (N_17452,N_16428,N_16401);
and U17453 (N_17453,N_16862,N_16839);
and U17454 (N_17454,N_16828,N_16290);
or U17455 (N_17455,N_16275,N_16761);
and U17456 (N_17456,N_16858,N_16495);
or U17457 (N_17457,N_16256,N_16476);
nor U17458 (N_17458,N_16474,N_16396);
nand U17459 (N_17459,N_16866,N_16431);
nor U17460 (N_17460,N_16316,N_16374);
nand U17461 (N_17461,N_16504,N_16291);
or U17462 (N_17462,N_16469,N_16581);
nand U17463 (N_17463,N_16343,N_16612);
and U17464 (N_17464,N_16374,N_16312);
nor U17465 (N_17465,N_16487,N_16252);
nor U17466 (N_17466,N_16746,N_16405);
nor U17467 (N_17467,N_16361,N_16693);
nor U17468 (N_17468,N_16816,N_16494);
nor U17469 (N_17469,N_16710,N_16498);
nand U17470 (N_17470,N_16250,N_16552);
nand U17471 (N_17471,N_16339,N_16333);
xnor U17472 (N_17472,N_16510,N_16643);
or U17473 (N_17473,N_16718,N_16761);
and U17474 (N_17474,N_16811,N_16614);
and U17475 (N_17475,N_16306,N_16826);
nand U17476 (N_17476,N_16619,N_16836);
nand U17477 (N_17477,N_16783,N_16389);
nor U17478 (N_17478,N_16605,N_16525);
nand U17479 (N_17479,N_16600,N_16442);
xnor U17480 (N_17480,N_16358,N_16359);
or U17481 (N_17481,N_16299,N_16659);
nand U17482 (N_17482,N_16797,N_16507);
nor U17483 (N_17483,N_16530,N_16279);
or U17484 (N_17484,N_16668,N_16257);
xnor U17485 (N_17485,N_16345,N_16403);
xnor U17486 (N_17486,N_16380,N_16558);
nand U17487 (N_17487,N_16577,N_16405);
xor U17488 (N_17488,N_16417,N_16669);
and U17489 (N_17489,N_16714,N_16340);
or U17490 (N_17490,N_16495,N_16659);
and U17491 (N_17491,N_16278,N_16536);
and U17492 (N_17492,N_16561,N_16283);
nand U17493 (N_17493,N_16611,N_16489);
nor U17494 (N_17494,N_16709,N_16698);
nand U17495 (N_17495,N_16569,N_16777);
nand U17496 (N_17496,N_16291,N_16775);
and U17497 (N_17497,N_16679,N_16418);
and U17498 (N_17498,N_16705,N_16668);
nand U17499 (N_17499,N_16265,N_16576);
and U17500 (N_17500,N_17433,N_16901);
nand U17501 (N_17501,N_16982,N_17334);
nand U17502 (N_17502,N_17317,N_17206);
or U17503 (N_17503,N_17204,N_17238);
nor U17504 (N_17504,N_16911,N_17213);
nand U17505 (N_17505,N_17114,N_17190);
nor U17506 (N_17506,N_17001,N_17093);
nand U17507 (N_17507,N_17233,N_17025);
and U17508 (N_17508,N_17182,N_16960);
nor U17509 (N_17509,N_17031,N_17336);
nor U17510 (N_17510,N_17309,N_17036);
nor U17511 (N_17511,N_17045,N_17287);
xor U17512 (N_17512,N_17485,N_16900);
nand U17513 (N_17513,N_17434,N_16884);
nand U17514 (N_17514,N_17062,N_17320);
nor U17515 (N_17515,N_17063,N_17165);
nor U17516 (N_17516,N_17117,N_17370);
xor U17517 (N_17517,N_16997,N_17424);
nor U17518 (N_17518,N_17030,N_17157);
xor U17519 (N_17519,N_17222,N_17112);
and U17520 (N_17520,N_17430,N_16895);
or U17521 (N_17521,N_17316,N_17197);
nor U17522 (N_17522,N_17249,N_17059);
or U17523 (N_17523,N_17286,N_17250);
or U17524 (N_17524,N_17361,N_17089);
nand U17525 (N_17525,N_17337,N_17200);
nor U17526 (N_17526,N_17472,N_17408);
nor U17527 (N_17527,N_17111,N_17259);
nor U17528 (N_17528,N_17094,N_17037);
and U17529 (N_17529,N_17479,N_17209);
nor U17530 (N_17530,N_17137,N_17332);
nor U17531 (N_17531,N_16959,N_17052);
xnor U17532 (N_17532,N_17470,N_17443);
nor U17533 (N_17533,N_17178,N_17431);
nand U17534 (N_17534,N_17151,N_17203);
and U17535 (N_17535,N_16938,N_17453);
and U17536 (N_17536,N_17406,N_16937);
or U17537 (N_17537,N_17444,N_17235);
nand U17538 (N_17538,N_17474,N_17409);
nor U17539 (N_17539,N_16880,N_17116);
nand U17540 (N_17540,N_17418,N_17065);
nor U17541 (N_17541,N_17283,N_16913);
xor U17542 (N_17542,N_17401,N_17263);
or U17543 (N_17543,N_17324,N_17016);
or U17544 (N_17544,N_17279,N_17303);
and U17545 (N_17545,N_17278,N_17145);
nand U17546 (N_17546,N_16886,N_17131);
or U17547 (N_17547,N_17373,N_17179);
nand U17548 (N_17548,N_16882,N_16973);
xnor U17549 (N_17549,N_16894,N_17271);
or U17550 (N_17550,N_17080,N_17244);
and U17551 (N_17551,N_16939,N_16955);
or U17552 (N_17552,N_17207,N_17374);
nor U17553 (N_17553,N_16970,N_16907);
and U17554 (N_17554,N_16898,N_17274);
nor U17555 (N_17555,N_17471,N_17293);
or U17556 (N_17556,N_16916,N_17099);
and U17557 (N_17557,N_17127,N_16885);
nand U17558 (N_17558,N_17139,N_17446);
nor U17559 (N_17559,N_16891,N_17422);
or U17560 (N_17560,N_17428,N_17024);
and U17561 (N_17561,N_16928,N_17218);
or U17562 (N_17562,N_17215,N_16931);
xor U17563 (N_17563,N_17224,N_17352);
and U17564 (N_17564,N_17199,N_17467);
xnor U17565 (N_17565,N_17393,N_17288);
and U17566 (N_17566,N_17313,N_17277);
xnor U17567 (N_17567,N_17386,N_17429);
nand U17568 (N_17568,N_17118,N_17040);
nor U17569 (N_17569,N_17009,N_17113);
or U17570 (N_17570,N_17342,N_17214);
and U17571 (N_17571,N_17410,N_17018);
and U17572 (N_17572,N_16947,N_17201);
or U17573 (N_17573,N_17302,N_17143);
and U17574 (N_17574,N_17110,N_17308);
and U17575 (N_17575,N_17000,N_17133);
nor U17576 (N_17576,N_16954,N_17395);
or U17577 (N_17577,N_17478,N_17101);
nor U17578 (N_17578,N_16967,N_16932);
nor U17579 (N_17579,N_17241,N_16943);
nor U17580 (N_17580,N_17448,N_17109);
or U17581 (N_17581,N_17482,N_17298);
nor U17582 (N_17582,N_16953,N_17069);
nand U17583 (N_17583,N_17384,N_17217);
xor U17584 (N_17584,N_17172,N_17311);
and U17585 (N_17585,N_17144,N_17276);
xnor U17586 (N_17586,N_17236,N_17362);
and U17587 (N_17587,N_17107,N_17003);
nand U17588 (N_17588,N_16879,N_17483);
or U17589 (N_17589,N_17439,N_16990);
and U17590 (N_17590,N_16989,N_17231);
xnor U17591 (N_17591,N_16996,N_17256);
nand U17592 (N_17592,N_16909,N_17310);
and U17593 (N_17593,N_17416,N_16976);
nand U17594 (N_17594,N_17380,N_17042);
or U17595 (N_17595,N_17141,N_17022);
nor U17596 (N_17596,N_17346,N_17437);
xor U17597 (N_17597,N_16889,N_17355);
and U17598 (N_17598,N_17152,N_17053);
and U17599 (N_17599,N_17035,N_17447);
nand U17600 (N_17600,N_17289,N_17198);
or U17601 (N_17601,N_17377,N_16887);
and U17602 (N_17602,N_17162,N_17125);
nand U17603 (N_17603,N_17014,N_17230);
or U17604 (N_17604,N_17449,N_17008);
and U17605 (N_17605,N_17385,N_16961);
nor U17606 (N_17606,N_17104,N_17105);
nor U17607 (N_17607,N_17375,N_17358);
and U17608 (N_17608,N_16966,N_17396);
nor U17609 (N_17609,N_17299,N_17173);
nor U17610 (N_17610,N_17387,N_16915);
and U17611 (N_17611,N_17294,N_17464);
and U17612 (N_17612,N_17079,N_17134);
nand U17613 (N_17613,N_17155,N_16919);
and U17614 (N_17614,N_17291,N_17329);
nor U17615 (N_17615,N_17028,N_17388);
nand U17616 (N_17616,N_17304,N_16994);
and U17617 (N_17617,N_17477,N_17347);
xnor U17618 (N_17618,N_17366,N_17120);
or U17619 (N_17619,N_17160,N_16899);
nor U17620 (N_17620,N_17136,N_17058);
nand U17621 (N_17621,N_17086,N_17297);
nand U17622 (N_17622,N_17247,N_17315);
or U17623 (N_17623,N_17475,N_17458);
xor U17624 (N_17624,N_17466,N_17026);
and U17625 (N_17625,N_17457,N_17212);
nor U17626 (N_17626,N_16925,N_16923);
or U17627 (N_17627,N_17252,N_16983);
nand U17628 (N_17628,N_16935,N_17002);
or U17629 (N_17629,N_17228,N_17184);
and U17630 (N_17630,N_17096,N_17415);
xnor U17631 (N_17631,N_17270,N_17229);
or U17632 (N_17632,N_17068,N_17378);
nand U17633 (N_17633,N_17195,N_17495);
xnor U17634 (N_17634,N_17340,N_17073);
nand U17635 (N_17635,N_17174,N_16974);
and U17636 (N_17636,N_17364,N_17292);
and U17637 (N_17637,N_17345,N_17454);
or U17638 (N_17638,N_17460,N_17142);
nand U17639 (N_17639,N_17463,N_16965);
and U17640 (N_17640,N_17436,N_17493);
nand U17641 (N_17641,N_16890,N_17285);
or U17642 (N_17642,N_17208,N_17435);
or U17643 (N_17643,N_16936,N_17284);
xnor U17644 (N_17644,N_17211,N_16948);
and U17645 (N_17645,N_17383,N_17216);
nand U17646 (N_17646,N_17234,N_17083);
nand U17647 (N_17647,N_17177,N_17491);
xnor U17648 (N_17648,N_16914,N_17459);
xnor U17649 (N_17649,N_16963,N_17456);
nand U17650 (N_17650,N_17124,N_17248);
nand U17651 (N_17651,N_16946,N_17156);
and U17652 (N_17652,N_17108,N_17426);
nor U17653 (N_17653,N_17027,N_17397);
nand U17654 (N_17654,N_17057,N_17251);
nand U17655 (N_17655,N_17402,N_16920);
or U17656 (N_17656,N_17067,N_17392);
nor U17657 (N_17657,N_16904,N_16888);
nand U17658 (N_17658,N_17264,N_17398);
nand U17659 (N_17659,N_17064,N_17044);
nand U17660 (N_17660,N_16940,N_17189);
nand U17661 (N_17661,N_17322,N_17084);
and U17662 (N_17662,N_17245,N_17029);
xor U17663 (N_17663,N_17301,N_17092);
xnor U17664 (N_17664,N_17305,N_17382);
and U17665 (N_17665,N_17066,N_17300);
and U17666 (N_17666,N_17074,N_17181);
nand U17667 (N_17667,N_17013,N_17462);
xor U17668 (N_17668,N_17452,N_17072);
nor U17669 (N_17669,N_16903,N_17306);
nand U17670 (N_17670,N_17441,N_17242);
nand U17671 (N_17671,N_17357,N_16942);
xor U17672 (N_17672,N_17328,N_17129);
nand U17673 (N_17673,N_17360,N_17330);
nor U17674 (N_17674,N_17489,N_17295);
nor U17675 (N_17675,N_17038,N_17379);
xnor U17676 (N_17676,N_17338,N_17090);
or U17677 (N_17677,N_17188,N_16881);
and U17678 (N_17678,N_17060,N_17240);
nand U17679 (N_17679,N_17411,N_17239);
nand U17680 (N_17680,N_17048,N_17150);
nor U17681 (N_17681,N_17341,N_17017);
nand U17682 (N_17682,N_17451,N_17255);
nand U17683 (N_17683,N_17275,N_16995);
nand U17684 (N_17684,N_16978,N_16896);
or U17685 (N_17685,N_16941,N_17423);
or U17686 (N_17686,N_16952,N_17220);
nor U17687 (N_17687,N_17266,N_17394);
nand U17688 (N_17688,N_17221,N_17047);
nand U17689 (N_17689,N_17497,N_17153);
and U17690 (N_17690,N_17268,N_17171);
and U17691 (N_17691,N_17267,N_17319);
nand U17692 (N_17692,N_17280,N_17243);
nor U17693 (N_17693,N_16972,N_17254);
and U17694 (N_17694,N_17138,N_17356);
and U17695 (N_17695,N_17161,N_17205);
and U17696 (N_17696,N_17186,N_17390);
or U17697 (N_17697,N_17168,N_17265);
or U17698 (N_17698,N_16992,N_16975);
and U17699 (N_17699,N_17095,N_17135);
nor U17700 (N_17700,N_16968,N_17175);
nor U17701 (N_17701,N_17253,N_17227);
and U17702 (N_17702,N_17365,N_16883);
or U17703 (N_17703,N_17326,N_17425);
nand U17704 (N_17704,N_17369,N_17032);
nor U17705 (N_17705,N_16918,N_17010);
xor U17706 (N_17706,N_17461,N_17055);
and U17707 (N_17707,N_17078,N_17331);
nand U17708 (N_17708,N_17445,N_16984);
nor U17709 (N_17709,N_17043,N_17158);
nand U17710 (N_17710,N_17166,N_17440);
nand U17711 (N_17711,N_17147,N_16964);
and U17712 (N_17712,N_17262,N_17033);
nor U17713 (N_17713,N_16988,N_17007);
nand U17714 (N_17714,N_17307,N_17019);
nor U17715 (N_17715,N_17046,N_17354);
nor U17716 (N_17716,N_17359,N_17498);
nand U17717 (N_17717,N_17149,N_17011);
and U17718 (N_17718,N_17473,N_16893);
xnor U17719 (N_17719,N_16957,N_17496);
and U17720 (N_17720,N_17403,N_17187);
and U17721 (N_17721,N_17076,N_17363);
nand U17722 (N_17722,N_17050,N_16922);
and U17723 (N_17723,N_16912,N_17061);
and U17724 (N_17724,N_17075,N_17194);
nor U17725 (N_17725,N_17494,N_17100);
nand U17726 (N_17726,N_16986,N_17492);
xor U17727 (N_17727,N_17081,N_17327);
or U17728 (N_17728,N_16956,N_16958);
nand U17729 (N_17729,N_16908,N_17469);
and U17730 (N_17730,N_17480,N_16991);
or U17731 (N_17731,N_17119,N_17097);
nand U17732 (N_17732,N_16921,N_17367);
nor U17733 (N_17733,N_17039,N_17071);
or U17734 (N_17734,N_17414,N_17413);
nand U17735 (N_17735,N_17232,N_17106);
or U17736 (N_17736,N_17407,N_17088);
xor U17737 (N_17737,N_17481,N_17132);
and U17738 (N_17738,N_17169,N_17091);
nand U17739 (N_17739,N_17349,N_17054);
nor U17740 (N_17740,N_17128,N_17077);
or U17741 (N_17741,N_16934,N_17223);
or U17742 (N_17742,N_17389,N_16878);
nand U17743 (N_17743,N_17368,N_17023);
and U17744 (N_17744,N_17318,N_17296);
and U17745 (N_17745,N_17183,N_17468);
or U17746 (N_17746,N_17126,N_17321);
nor U17747 (N_17747,N_17412,N_17432);
and U17748 (N_17748,N_16977,N_17314);
or U17749 (N_17749,N_17115,N_17202);
and U17750 (N_17750,N_17405,N_17034);
nor U17751 (N_17751,N_16924,N_16910);
nor U17752 (N_17752,N_17192,N_17176);
nand U17753 (N_17753,N_17348,N_17122);
or U17754 (N_17754,N_17005,N_17258);
or U17755 (N_17755,N_17420,N_17419);
nand U17756 (N_17756,N_17159,N_17015);
or U17757 (N_17757,N_17269,N_17281);
nand U17758 (N_17758,N_17323,N_16906);
and U17759 (N_17759,N_17465,N_17140);
nand U17760 (N_17760,N_16917,N_17021);
nand U17761 (N_17761,N_17372,N_17056);
or U17762 (N_17762,N_17487,N_16930);
nand U17763 (N_17763,N_17051,N_17103);
and U17764 (N_17764,N_17381,N_17376);
nand U17765 (N_17765,N_17391,N_17225);
or U17766 (N_17766,N_17148,N_17226);
and U17767 (N_17767,N_17098,N_16980);
xnor U17768 (N_17768,N_17164,N_17163);
nor U17769 (N_17769,N_17070,N_17421);
xnor U17770 (N_17770,N_16950,N_17012);
nand U17771 (N_17771,N_17427,N_17082);
xnor U17772 (N_17772,N_17351,N_16987);
and U17773 (N_17773,N_17325,N_16897);
or U17774 (N_17774,N_17261,N_17438);
and U17775 (N_17775,N_17353,N_17130);
nand U17776 (N_17776,N_16979,N_17237);
xnor U17777 (N_17777,N_17154,N_17490);
or U17778 (N_17778,N_16985,N_17146);
or U17779 (N_17779,N_16927,N_16999);
or U17780 (N_17780,N_17087,N_17180);
and U17781 (N_17781,N_17219,N_17085);
nand U17782 (N_17782,N_17484,N_17335);
or U17783 (N_17783,N_17006,N_17196);
xnor U17784 (N_17784,N_17041,N_17020);
or U17785 (N_17785,N_17350,N_17123);
and U17786 (N_17786,N_16981,N_17442);
or U17787 (N_17787,N_16933,N_17312);
xnor U17788 (N_17788,N_17246,N_17450);
xor U17789 (N_17789,N_16875,N_17339);
or U17790 (N_17790,N_17404,N_16945);
nand U17791 (N_17791,N_17400,N_16877);
and U17792 (N_17792,N_17399,N_17290);
nor U17793 (N_17793,N_16993,N_17185);
and U17794 (N_17794,N_17371,N_17121);
or U17795 (N_17795,N_17488,N_17343);
and U17796 (N_17796,N_16944,N_17282);
nand U17797 (N_17797,N_16892,N_17167);
xor U17798 (N_17798,N_17260,N_16876);
nor U17799 (N_17799,N_16902,N_16951);
nand U17800 (N_17800,N_17210,N_17333);
or U17801 (N_17801,N_16905,N_17344);
nand U17802 (N_17802,N_16949,N_17191);
and U17803 (N_17803,N_17476,N_17170);
nand U17804 (N_17804,N_17272,N_16926);
or U17805 (N_17805,N_17455,N_16962);
nand U17806 (N_17806,N_17257,N_17004);
or U17807 (N_17807,N_16998,N_17273);
and U17808 (N_17808,N_17486,N_17049);
nand U17809 (N_17809,N_17102,N_17193);
xor U17810 (N_17810,N_16969,N_16971);
or U17811 (N_17811,N_17499,N_17417);
nor U17812 (N_17812,N_16929,N_17185);
and U17813 (N_17813,N_17089,N_16962);
or U17814 (N_17814,N_17215,N_16959);
or U17815 (N_17815,N_17288,N_17203);
nand U17816 (N_17816,N_17099,N_17169);
or U17817 (N_17817,N_17352,N_17054);
or U17818 (N_17818,N_17121,N_16943);
and U17819 (N_17819,N_17099,N_16992);
nand U17820 (N_17820,N_17079,N_17059);
or U17821 (N_17821,N_17271,N_16883);
nand U17822 (N_17822,N_17074,N_17086);
or U17823 (N_17823,N_16931,N_17268);
nor U17824 (N_17824,N_17018,N_17295);
nor U17825 (N_17825,N_17203,N_17397);
nor U17826 (N_17826,N_17362,N_17422);
nand U17827 (N_17827,N_17382,N_17076);
xnor U17828 (N_17828,N_16896,N_17254);
xnor U17829 (N_17829,N_16974,N_17378);
nand U17830 (N_17830,N_17426,N_17114);
nor U17831 (N_17831,N_17002,N_17375);
or U17832 (N_17832,N_16938,N_17376);
and U17833 (N_17833,N_17241,N_16906);
nor U17834 (N_17834,N_17401,N_16988);
nor U17835 (N_17835,N_17461,N_17135);
and U17836 (N_17836,N_17256,N_17136);
xnor U17837 (N_17837,N_17387,N_17095);
nor U17838 (N_17838,N_16883,N_17170);
nor U17839 (N_17839,N_17098,N_17145);
nand U17840 (N_17840,N_17109,N_16907);
nand U17841 (N_17841,N_17146,N_17112);
nand U17842 (N_17842,N_17458,N_16909);
or U17843 (N_17843,N_17072,N_17495);
or U17844 (N_17844,N_17198,N_16901);
and U17845 (N_17845,N_17488,N_17332);
or U17846 (N_17846,N_17105,N_17120);
and U17847 (N_17847,N_17031,N_17473);
nor U17848 (N_17848,N_16934,N_17158);
or U17849 (N_17849,N_17179,N_17494);
or U17850 (N_17850,N_17486,N_17001);
nor U17851 (N_17851,N_16931,N_17279);
and U17852 (N_17852,N_17273,N_17365);
or U17853 (N_17853,N_17380,N_17378);
or U17854 (N_17854,N_17148,N_17213);
or U17855 (N_17855,N_16956,N_17226);
or U17856 (N_17856,N_17130,N_17387);
nand U17857 (N_17857,N_17048,N_17459);
and U17858 (N_17858,N_17225,N_17011);
and U17859 (N_17859,N_17178,N_17106);
and U17860 (N_17860,N_16967,N_17291);
nor U17861 (N_17861,N_17202,N_17058);
and U17862 (N_17862,N_16962,N_17355);
or U17863 (N_17863,N_17093,N_17309);
nand U17864 (N_17864,N_16915,N_17321);
and U17865 (N_17865,N_16905,N_17336);
xor U17866 (N_17866,N_17300,N_16908);
nand U17867 (N_17867,N_16967,N_17497);
and U17868 (N_17868,N_17111,N_17234);
nand U17869 (N_17869,N_17148,N_16889);
or U17870 (N_17870,N_17323,N_17456);
or U17871 (N_17871,N_17074,N_17459);
nor U17872 (N_17872,N_17220,N_17028);
or U17873 (N_17873,N_17168,N_17105);
nor U17874 (N_17874,N_17309,N_17029);
nand U17875 (N_17875,N_17457,N_16882);
or U17876 (N_17876,N_17048,N_17372);
and U17877 (N_17877,N_16985,N_16909);
and U17878 (N_17878,N_17072,N_16905);
and U17879 (N_17879,N_17238,N_17091);
nand U17880 (N_17880,N_17468,N_17058);
or U17881 (N_17881,N_16891,N_17168);
nor U17882 (N_17882,N_17086,N_17103);
or U17883 (N_17883,N_17357,N_17169);
nand U17884 (N_17884,N_17377,N_17472);
xnor U17885 (N_17885,N_17172,N_17134);
or U17886 (N_17886,N_17106,N_17444);
nand U17887 (N_17887,N_17084,N_17191);
nand U17888 (N_17888,N_17399,N_17284);
nand U17889 (N_17889,N_17240,N_16902);
nand U17890 (N_17890,N_16977,N_17149);
nand U17891 (N_17891,N_17245,N_17053);
and U17892 (N_17892,N_17287,N_17117);
or U17893 (N_17893,N_17244,N_17229);
or U17894 (N_17894,N_17162,N_16998);
nor U17895 (N_17895,N_17184,N_16887);
and U17896 (N_17896,N_16919,N_17317);
nand U17897 (N_17897,N_16891,N_16921);
nor U17898 (N_17898,N_16875,N_17158);
and U17899 (N_17899,N_16881,N_17295);
nand U17900 (N_17900,N_17032,N_17333);
nor U17901 (N_17901,N_16991,N_17077);
nor U17902 (N_17902,N_17209,N_16966);
xor U17903 (N_17903,N_16926,N_17410);
nand U17904 (N_17904,N_16983,N_17348);
and U17905 (N_17905,N_16929,N_17091);
or U17906 (N_17906,N_17003,N_17289);
or U17907 (N_17907,N_17143,N_17346);
and U17908 (N_17908,N_17178,N_16971);
nor U17909 (N_17909,N_16973,N_17093);
nand U17910 (N_17910,N_17482,N_17362);
or U17911 (N_17911,N_16911,N_17081);
and U17912 (N_17912,N_17123,N_17088);
xnor U17913 (N_17913,N_17123,N_17484);
nand U17914 (N_17914,N_17437,N_17491);
or U17915 (N_17915,N_17174,N_16995);
nor U17916 (N_17916,N_17192,N_17459);
nor U17917 (N_17917,N_16915,N_17055);
and U17918 (N_17918,N_16929,N_17058);
nand U17919 (N_17919,N_17358,N_17239);
nor U17920 (N_17920,N_17345,N_17415);
nand U17921 (N_17921,N_17229,N_17051);
nand U17922 (N_17922,N_17086,N_17246);
and U17923 (N_17923,N_17104,N_17134);
or U17924 (N_17924,N_17348,N_17070);
or U17925 (N_17925,N_17011,N_17260);
or U17926 (N_17926,N_16913,N_17371);
nor U17927 (N_17927,N_16887,N_17271);
nor U17928 (N_17928,N_16892,N_17339);
nor U17929 (N_17929,N_17118,N_17397);
nand U17930 (N_17930,N_17200,N_17471);
nand U17931 (N_17931,N_17429,N_17120);
xnor U17932 (N_17932,N_17049,N_17451);
nand U17933 (N_17933,N_17323,N_17230);
and U17934 (N_17934,N_17338,N_17290);
and U17935 (N_17935,N_17228,N_17203);
nor U17936 (N_17936,N_17235,N_17022);
or U17937 (N_17937,N_17301,N_16897);
and U17938 (N_17938,N_17293,N_17072);
nor U17939 (N_17939,N_17392,N_17254);
nand U17940 (N_17940,N_17279,N_17124);
nand U17941 (N_17941,N_16973,N_16889);
or U17942 (N_17942,N_17189,N_17269);
and U17943 (N_17943,N_16918,N_17200);
nand U17944 (N_17944,N_17053,N_17411);
xor U17945 (N_17945,N_17280,N_17221);
nor U17946 (N_17946,N_16890,N_17352);
xor U17947 (N_17947,N_17432,N_17227);
and U17948 (N_17948,N_17416,N_17223);
or U17949 (N_17949,N_17121,N_17061);
or U17950 (N_17950,N_17285,N_17369);
and U17951 (N_17951,N_17136,N_16876);
nand U17952 (N_17952,N_17309,N_16997);
and U17953 (N_17953,N_17344,N_17332);
nor U17954 (N_17954,N_17303,N_16921);
nor U17955 (N_17955,N_17243,N_17011);
nor U17956 (N_17956,N_17367,N_17244);
or U17957 (N_17957,N_17160,N_17407);
nor U17958 (N_17958,N_16875,N_17137);
and U17959 (N_17959,N_17385,N_17143);
or U17960 (N_17960,N_17481,N_17201);
and U17961 (N_17961,N_16961,N_17207);
and U17962 (N_17962,N_16977,N_17372);
or U17963 (N_17963,N_16950,N_17301);
or U17964 (N_17964,N_16916,N_17236);
xnor U17965 (N_17965,N_17101,N_16901);
and U17966 (N_17966,N_17045,N_17035);
nor U17967 (N_17967,N_17374,N_17215);
or U17968 (N_17968,N_16961,N_17121);
nor U17969 (N_17969,N_17012,N_17455);
nor U17970 (N_17970,N_17283,N_17050);
nor U17971 (N_17971,N_17150,N_17418);
nor U17972 (N_17972,N_17428,N_16956);
nand U17973 (N_17973,N_17111,N_16910);
xor U17974 (N_17974,N_17040,N_17025);
and U17975 (N_17975,N_16909,N_17054);
and U17976 (N_17976,N_17080,N_17121);
and U17977 (N_17977,N_17136,N_17150);
and U17978 (N_17978,N_16897,N_17142);
nand U17979 (N_17979,N_17049,N_17242);
nor U17980 (N_17980,N_16982,N_17328);
nor U17981 (N_17981,N_17012,N_17405);
nand U17982 (N_17982,N_17192,N_17479);
xnor U17983 (N_17983,N_17316,N_17262);
xnor U17984 (N_17984,N_16959,N_16914);
or U17985 (N_17985,N_16956,N_17114);
nor U17986 (N_17986,N_16878,N_16955);
xor U17987 (N_17987,N_17472,N_17447);
nor U17988 (N_17988,N_16878,N_17028);
xnor U17989 (N_17989,N_17061,N_17492);
or U17990 (N_17990,N_17452,N_17265);
nor U17991 (N_17991,N_17260,N_17161);
nand U17992 (N_17992,N_17034,N_17084);
nor U17993 (N_17993,N_17281,N_17408);
and U17994 (N_17994,N_17445,N_17329);
or U17995 (N_17995,N_17416,N_17410);
xor U17996 (N_17996,N_17407,N_17197);
nor U17997 (N_17997,N_17030,N_16916);
nor U17998 (N_17998,N_16914,N_17400);
or U17999 (N_17999,N_17003,N_17369);
nand U18000 (N_18000,N_17115,N_17298);
and U18001 (N_18001,N_17217,N_17345);
nand U18002 (N_18002,N_17385,N_17071);
and U18003 (N_18003,N_17276,N_17485);
xnor U18004 (N_18004,N_16893,N_17432);
and U18005 (N_18005,N_17415,N_16903);
nor U18006 (N_18006,N_17200,N_16987);
and U18007 (N_18007,N_17232,N_17135);
nor U18008 (N_18008,N_17316,N_17336);
and U18009 (N_18009,N_17288,N_17149);
xnor U18010 (N_18010,N_17358,N_17306);
xnor U18011 (N_18011,N_17377,N_17408);
and U18012 (N_18012,N_17385,N_16929);
nor U18013 (N_18013,N_17065,N_16906);
or U18014 (N_18014,N_17226,N_17382);
nor U18015 (N_18015,N_16957,N_17480);
xnor U18016 (N_18016,N_17017,N_17059);
nand U18017 (N_18017,N_17490,N_17092);
nor U18018 (N_18018,N_17304,N_17278);
or U18019 (N_18019,N_17019,N_16940);
or U18020 (N_18020,N_17356,N_17007);
or U18021 (N_18021,N_17275,N_16955);
nor U18022 (N_18022,N_16939,N_17381);
nand U18023 (N_18023,N_17008,N_17066);
nand U18024 (N_18024,N_17275,N_17132);
nand U18025 (N_18025,N_16945,N_17121);
or U18026 (N_18026,N_17159,N_17362);
xor U18027 (N_18027,N_17186,N_17230);
and U18028 (N_18028,N_17201,N_17416);
and U18029 (N_18029,N_17428,N_17296);
nand U18030 (N_18030,N_16958,N_17117);
xnor U18031 (N_18031,N_17034,N_17340);
or U18032 (N_18032,N_17133,N_17163);
or U18033 (N_18033,N_16962,N_17181);
nor U18034 (N_18034,N_17000,N_17313);
nand U18035 (N_18035,N_17312,N_17037);
or U18036 (N_18036,N_17305,N_17349);
and U18037 (N_18037,N_17364,N_17117);
or U18038 (N_18038,N_16965,N_16929);
xnor U18039 (N_18039,N_17060,N_17185);
and U18040 (N_18040,N_17420,N_17007);
nor U18041 (N_18041,N_17287,N_17361);
or U18042 (N_18042,N_17275,N_17192);
and U18043 (N_18043,N_17479,N_17363);
xnor U18044 (N_18044,N_17096,N_17373);
or U18045 (N_18045,N_16956,N_17149);
or U18046 (N_18046,N_17450,N_17404);
and U18047 (N_18047,N_16985,N_17322);
or U18048 (N_18048,N_17257,N_17453);
nor U18049 (N_18049,N_17271,N_17223);
or U18050 (N_18050,N_17335,N_17338);
or U18051 (N_18051,N_17254,N_17069);
nor U18052 (N_18052,N_17408,N_17265);
or U18053 (N_18053,N_17175,N_17394);
nor U18054 (N_18054,N_17056,N_16968);
or U18055 (N_18055,N_17353,N_17254);
or U18056 (N_18056,N_17257,N_17416);
or U18057 (N_18057,N_16995,N_16980);
and U18058 (N_18058,N_17402,N_17378);
nor U18059 (N_18059,N_16943,N_17354);
nor U18060 (N_18060,N_17182,N_17449);
or U18061 (N_18061,N_17261,N_17065);
nand U18062 (N_18062,N_16928,N_17465);
or U18063 (N_18063,N_17310,N_16935);
nor U18064 (N_18064,N_17475,N_17365);
nor U18065 (N_18065,N_17420,N_17164);
nand U18066 (N_18066,N_17471,N_16877);
xor U18067 (N_18067,N_16948,N_17209);
nand U18068 (N_18068,N_17193,N_17166);
nor U18069 (N_18069,N_17003,N_17225);
or U18070 (N_18070,N_17384,N_17132);
nand U18071 (N_18071,N_16961,N_17420);
nor U18072 (N_18072,N_17306,N_17444);
and U18073 (N_18073,N_17087,N_16966);
nand U18074 (N_18074,N_17089,N_17255);
or U18075 (N_18075,N_17137,N_17262);
or U18076 (N_18076,N_17055,N_16972);
and U18077 (N_18077,N_16905,N_17275);
nor U18078 (N_18078,N_17323,N_16987);
and U18079 (N_18079,N_17020,N_17216);
and U18080 (N_18080,N_17128,N_17401);
nor U18081 (N_18081,N_17315,N_17206);
nor U18082 (N_18082,N_17101,N_17383);
and U18083 (N_18083,N_17224,N_16904);
nand U18084 (N_18084,N_16922,N_17056);
nand U18085 (N_18085,N_17323,N_17130);
nor U18086 (N_18086,N_16960,N_17099);
or U18087 (N_18087,N_17403,N_17471);
xor U18088 (N_18088,N_16993,N_17012);
nor U18089 (N_18089,N_17031,N_17225);
and U18090 (N_18090,N_17266,N_16927);
or U18091 (N_18091,N_17306,N_17433);
nand U18092 (N_18092,N_17494,N_17192);
nand U18093 (N_18093,N_16910,N_16984);
nand U18094 (N_18094,N_17302,N_16955);
nand U18095 (N_18095,N_17172,N_17040);
xor U18096 (N_18096,N_16931,N_17087);
or U18097 (N_18097,N_17266,N_17213);
xor U18098 (N_18098,N_17272,N_16898);
nand U18099 (N_18099,N_17468,N_16978);
or U18100 (N_18100,N_17271,N_17225);
nor U18101 (N_18101,N_16900,N_17468);
nor U18102 (N_18102,N_17172,N_17316);
and U18103 (N_18103,N_17195,N_17385);
or U18104 (N_18104,N_16903,N_16989);
and U18105 (N_18105,N_16996,N_17064);
or U18106 (N_18106,N_17434,N_17398);
nor U18107 (N_18107,N_17388,N_17007);
and U18108 (N_18108,N_17243,N_16904);
or U18109 (N_18109,N_17313,N_17205);
or U18110 (N_18110,N_17449,N_17228);
nand U18111 (N_18111,N_16876,N_17456);
or U18112 (N_18112,N_17259,N_16964);
nor U18113 (N_18113,N_17002,N_17095);
nand U18114 (N_18114,N_17227,N_17007);
nand U18115 (N_18115,N_17040,N_17483);
and U18116 (N_18116,N_17399,N_17129);
nand U18117 (N_18117,N_17153,N_17062);
or U18118 (N_18118,N_16998,N_17047);
nor U18119 (N_18119,N_17111,N_17301);
nor U18120 (N_18120,N_17093,N_17403);
and U18121 (N_18121,N_17236,N_17330);
xnor U18122 (N_18122,N_17041,N_17094);
nor U18123 (N_18123,N_17143,N_17137);
and U18124 (N_18124,N_17130,N_17227);
or U18125 (N_18125,N_18066,N_17561);
nand U18126 (N_18126,N_17995,N_17637);
or U18127 (N_18127,N_17673,N_17866);
and U18128 (N_18128,N_17689,N_17534);
xnor U18129 (N_18129,N_17829,N_17849);
xor U18130 (N_18130,N_17724,N_17874);
xnor U18131 (N_18131,N_17973,N_17532);
and U18132 (N_18132,N_17962,N_17794);
and U18133 (N_18133,N_17654,N_18080);
or U18134 (N_18134,N_17584,N_18033);
nand U18135 (N_18135,N_17509,N_17606);
nand U18136 (N_18136,N_18096,N_17690);
and U18137 (N_18137,N_17602,N_17708);
or U18138 (N_18138,N_17862,N_17635);
xnor U18139 (N_18139,N_17957,N_17868);
nand U18140 (N_18140,N_17738,N_17744);
xnor U18141 (N_18141,N_17552,N_17861);
or U18142 (N_18142,N_17609,N_18003);
nor U18143 (N_18143,N_18043,N_17528);
and U18144 (N_18144,N_17770,N_17547);
and U18145 (N_18145,N_17853,N_17808);
and U18146 (N_18146,N_17684,N_17723);
nor U18147 (N_18147,N_18027,N_17951);
and U18148 (N_18148,N_17856,N_17508);
xor U18149 (N_18149,N_18065,N_17942);
or U18150 (N_18150,N_17809,N_17877);
nand U18151 (N_18151,N_17865,N_17860);
or U18152 (N_18152,N_18014,N_17700);
and U18153 (N_18153,N_17913,N_17638);
or U18154 (N_18154,N_17789,N_18054);
or U18155 (N_18155,N_17766,N_17823);
nand U18156 (N_18156,N_17947,N_17728);
nand U18157 (N_18157,N_17969,N_17870);
or U18158 (N_18158,N_17627,N_17767);
nor U18159 (N_18159,N_17935,N_17990);
or U18160 (N_18160,N_17880,N_18036);
nand U18161 (N_18161,N_17790,N_17979);
nor U18162 (N_18162,N_17692,N_17936);
and U18163 (N_18163,N_17573,N_17858);
and U18164 (N_18164,N_18034,N_17838);
nand U18165 (N_18165,N_17578,N_17590);
or U18166 (N_18166,N_17668,N_17907);
nand U18167 (N_18167,N_17966,N_17616);
or U18168 (N_18168,N_17650,N_17816);
nor U18169 (N_18169,N_17911,N_17575);
and U18170 (N_18170,N_17903,N_18078);
and U18171 (N_18171,N_18072,N_17747);
or U18172 (N_18172,N_17831,N_17782);
and U18173 (N_18173,N_17893,N_17642);
and U18174 (N_18174,N_17683,N_17727);
and U18175 (N_18175,N_18094,N_17956);
nor U18176 (N_18176,N_17647,N_17834);
nor U18177 (N_18177,N_17719,N_17653);
nand U18178 (N_18178,N_18093,N_17878);
nor U18179 (N_18179,N_17793,N_17639);
nor U18180 (N_18180,N_17945,N_18097);
nor U18181 (N_18181,N_17787,N_17984);
or U18182 (N_18182,N_17539,N_17546);
nand U18183 (N_18183,N_18047,N_18110);
nor U18184 (N_18184,N_17730,N_17851);
nand U18185 (N_18185,N_17614,N_17677);
xnor U18186 (N_18186,N_17693,N_18109);
nand U18187 (N_18187,N_17734,N_17769);
nand U18188 (N_18188,N_17845,N_17537);
or U18189 (N_18189,N_18042,N_18108);
nand U18190 (N_18190,N_17612,N_17622);
xor U18191 (N_18191,N_18114,N_17615);
and U18192 (N_18192,N_17895,N_17522);
and U18193 (N_18193,N_17797,N_17567);
and U18194 (N_18194,N_17970,N_17843);
or U18195 (N_18195,N_17560,N_17545);
nand U18196 (N_18196,N_18016,N_17515);
nand U18197 (N_18197,N_17520,N_17804);
nand U18198 (N_18198,N_17748,N_17523);
nor U18199 (N_18199,N_17892,N_18099);
nor U18200 (N_18200,N_17764,N_17822);
or U18201 (N_18201,N_17771,N_17781);
or U18202 (N_18202,N_17910,N_17646);
or U18203 (N_18203,N_17553,N_18051);
or U18204 (N_18204,N_17817,N_18120);
nand U18205 (N_18205,N_17691,N_18035);
nand U18206 (N_18206,N_17848,N_17811);
nand U18207 (N_18207,N_17983,N_17674);
or U18208 (N_18208,N_18061,N_18117);
nor U18209 (N_18209,N_17980,N_17830);
or U18210 (N_18210,N_18102,N_17887);
or U18211 (N_18211,N_17824,N_18083);
or U18212 (N_18212,N_17750,N_18029);
or U18213 (N_18213,N_17786,N_17967);
nor U18214 (N_18214,N_17720,N_17699);
nor U18215 (N_18215,N_17897,N_17918);
and U18216 (N_18216,N_18019,N_18113);
nand U18217 (N_18217,N_17576,N_17896);
and U18218 (N_18218,N_18067,N_18021);
nand U18219 (N_18219,N_18026,N_17976);
xnor U18220 (N_18220,N_17890,N_17605);
nand U18221 (N_18221,N_17569,N_18122);
and U18222 (N_18222,N_17931,N_17521);
nand U18223 (N_18223,N_17991,N_18062);
nor U18224 (N_18224,N_18008,N_17826);
nor U18225 (N_18225,N_17999,N_17978);
or U18226 (N_18226,N_17565,N_17755);
nand U18227 (N_18227,N_18090,N_18037);
nor U18228 (N_18228,N_17968,N_18046);
and U18229 (N_18229,N_17923,N_17617);
and U18230 (N_18230,N_17680,N_17921);
and U18231 (N_18231,N_18118,N_17675);
or U18232 (N_18232,N_17595,N_17981);
nand U18233 (N_18233,N_17618,N_17608);
nand U18234 (N_18234,N_17871,N_17721);
nand U18235 (N_18235,N_17549,N_17542);
or U18236 (N_18236,N_17846,N_17884);
or U18237 (N_18237,N_17676,N_17917);
nand U18238 (N_18238,N_18025,N_17511);
nand U18239 (N_18239,N_17555,N_17814);
or U18240 (N_18240,N_17556,N_17795);
nand U18241 (N_18241,N_17624,N_18020);
nand U18242 (N_18242,N_17570,N_17517);
xnor U18243 (N_18243,N_17807,N_17704);
and U18244 (N_18244,N_18049,N_17577);
nor U18245 (N_18245,N_17526,N_17538);
nand U18246 (N_18246,N_18100,N_18063);
and U18247 (N_18247,N_17579,N_17964);
and U18248 (N_18248,N_17827,N_17876);
nor U18249 (N_18249,N_17670,N_17792);
and U18250 (N_18250,N_18001,N_17930);
nand U18251 (N_18251,N_17732,N_18112);
nor U18252 (N_18252,N_18011,N_17953);
nand U18253 (N_18253,N_17869,N_17682);
or U18254 (N_18254,N_17788,N_17773);
nor U18255 (N_18255,N_17735,N_17941);
nand U18256 (N_18256,N_17630,N_17919);
nand U18257 (N_18257,N_17939,N_18073);
and U18258 (N_18258,N_17601,N_17714);
or U18259 (N_18259,N_17629,N_17558);
nor U18260 (N_18260,N_17658,N_17599);
or U18261 (N_18261,N_17888,N_18107);
xor U18262 (N_18262,N_17985,N_18071);
or U18263 (N_18263,N_17836,N_17971);
nand U18264 (N_18264,N_18119,N_18116);
nor U18265 (N_18265,N_17926,N_17711);
or U18266 (N_18266,N_17933,N_18024);
nor U18267 (N_18267,N_17551,N_17524);
nor U18268 (N_18268,N_17803,N_17882);
nor U18269 (N_18269,N_17841,N_17927);
and U18270 (N_18270,N_17932,N_17663);
nor U18271 (N_18271,N_17655,N_17548);
or U18272 (N_18272,N_18087,N_17864);
or U18273 (N_18273,N_17916,N_18057);
or U18274 (N_18274,N_17960,N_18088);
nor U18275 (N_18275,N_17881,N_17664);
or U18276 (N_18276,N_17800,N_17581);
or U18277 (N_18277,N_18038,N_18040);
or U18278 (N_18278,N_18064,N_18115);
nor U18279 (N_18279,N_17571,N_18053);
nor U18280 (N_18280,N_17514,N_18013);
or U18281 (N_18281,N_17610,N_17974);
and U18282 (N_18282,N_17661,N_17733);
nand U18283 (N_18283,N_18081,N_17656);
nand U18284 (N_18284,N_17925,N_17975);
nand U18285 (N_18285,N_17961,N_17889);
xor U18286 (N_18286,N_17988,N_17943);
and U18287 (N_18287,N_17937,N_17620);
xnor U18288 (N_18288,N_17996,N_17959);
xor U18289 (N_18289,N_17594,N_17710);
nor U18290 (N_18290,N_17530,N_18044);
or U18291 (N_18291,N_17867,N_17667);
nand U18292 (N_18292,N_17702,N_17543);
and U18293 (N_18293,N_17621,N_17852);
and U18294 (N_18294,N_17994,N_18074);
nor U18295 (N_18295,N_17940,N_17778);
or U18296 (N_18296,N_17885,N_18077);
xor U18297 (N_18297,N_17687,N_17593);
nor U18298 (N_18298,N_17688,N_17791);
nor U18299 (N_18299,N_18023,N_17516);
nor U18300 (N_18300,N_18085,N_17669);
nand U18301 (N_18301,N_17905,N_18068);
nand U18302 (N_18302,N_17761,N_17562);
nand U18303 (N_18303,N_17920,N_17850);
nor U18304 (N_18304,N_17540,N_18048);
nor U18305 (N_18305,N_18030,N_17706);
or U18306 (N_18306,N_17934,N_17844);
and U18307 (N_18307,N_17697,N_17740);
or U18308 (N_18308,N_17745,N_18079);
nor U18309 (N_18309,N_18000,N_17950);
nor U18310 (N_18310,N_17666,N_17652);
nor U18311 (N_18311,N_17762,N_17828);
and U18312 (N_18312,N_17802,N_18069);
and U18313 (N_18313,N_17760,N_17722);
nor U18314 (N_18314,N_17891,N_17922);
nand U18315 (N_18315,N_17908,N_17703);
or U18316 (N_18316,N_18028,N_17997);
nand U18317 (N_18317,N_17725,N_18022);
and U18318 (N_18318,N_18056,N_17554);
nand U18319 (N_18319,N_17505,N_17672);
nor U18320 (N_18320,N_17686,N_17557);
or U18321 (N_18321,N_17671,N_18050);
or U18322 (N_18322,N_18032,N_18009);
and U18323 (N_18323,N_18017,N_17883);
nand U18324 (N_18324,N_17518,N_17519);
nor U18325 (N_18325,N_18058,N_17946);
xor U18326 (N_18326,N_17712,N_17582);
or U18327 (N_18327,N_18002,N_17713);
or U18328 (N_18328,N_17863,N_18004);
nor U18329 (N_18329,N_17564,N_17963);
or U18330 (N_18330,N_17813,N_18010);
and U18331 (N_18331,N_17806,N_17758);
nor U18332 (N_18332,N_17580,N_18105);
nand U18333 (N_18333,N_17596,N_17659);
nor U18334 (N_18334,N_18055,N_17749);
nor U18335 (N_18335,N_17533,N_17815);
nand U18336 (N_18336,N_17527,N_17998);
nand U18337 (N_18337,N_17611,N_17900);
or U18338 (N_18338,N_17741,N_17801);
nand U18339 (N_18339,N_18124,N_17736);
and U18340 (N_18340,N_17625,N_18059);
and U18341 (N_18341,N_18041,N_17541);
xor U18342 (N_18342,N_17512,N_17879);
nor U18343 (N_18343,N_17717,N_17525);
and U18344 (N_18344,N_18095,N_18086);
nor U18345 (N_18345,N_17774,N_17886);
and U18346 (N_18346,N_17698,N_17949);
and U18347 (N_18347,N_17644,N_17597);
nor U18348 (N_18348,N_17757,N_17657);
nor U18349 (N_18349,N_17598,N_17914);
and U18350 (N_18350,N_17531,N_17742);
nor U18351 (N_18351,N_17909,N_17535);
and U18352 (N_18352,N_17912,N_18091);
nor U18353 (N_18353,N_17607,N_17752);
xor U18354 (N_18354,N_17948,N_17855);
xnor U18355 (N_18355,N_17501,N_17681);
nand U18356 (N_18356,N_17660,N_18089);
or U18357 (N_18357,N_17513,N_17928);
and U18358 (N_18358,N_17894,N_18082);
and U18359 (N_18359,N_17854,N_17604);
or U18360 (N_18360,N_17634,N_17768);
xor U18361 (N_18361,N_18121,N_17628);
and U18362 (N_18362,N_17759,N_17833);
nand U18363 (N_18363,N_17847,N_18012);
nor U18364 (N_18364,N_17772,N_17623);
nand U18365 (N_18365,N_18007,N_17965);
nand U18366 (N_18366,N_18060,N_17812);
and U18367 (N_18367,N_17636,N_18104);
nand U18368 (N_18368,N_17662,N_17753);
xor U18369 (N_18369,N_17583,N_17678);
or U18370 (N_18370,N_18092,N_17756);
or U18371 (N_18371,N_17777,N_18052);
nand U18372 (N_18372,N_17643,N_17987);
nor U18373 (N_18373,N_17600,N_17648);
nor U18374 (N_18374,N_17819,N_17743);
and U18375 (N_18375,N_18106,N_17603);
xnor U18376 (N_18376,N_17837,N_18084);
and U18377 (N_18377,N_17729,N_17685);
or U18378 (N_18378,N_17589,N_17776);
nand U18379 (N_18379,N_17718,N_18101);
nand U18380 (N_18380,N_17857,N_18018);
and U18381 (N_18381,N_17765,N_17779);
nand U18382 (N_18382,N_18103,N_17563);
or U18383 (N_18383,N_17825,N_17784);
nor U18384 (N_18384,N_17739,N_17754);
nand U18385 (N_18385,N_17592,N_17529);
and U18386 (N_18386,N_17641,N_17550);
nand U18387 (N_18387,N_17954,N_17679);
and U18388 (N_18388,N_17588,N_17707);
nand U18389 (N_18389,N_17559,N_17977);
nand U18390 (N_18390,N_17619,N_17986);
nor U18391 (N_18391,N_17510,N_17566);
and U18392 (N_18392,N_18123,N_17709);
or U18393 (N_18393,N_17737,N_17785);
or U18394 (N_18394,N_17839,N_17972);
nand U18395 (N_18395,N_17842,N_17536);
and U18396 (N_18396,N_17632,N_17716);
nand U18397 (N_18397,N_17915,N_17780);
and U18398 (N_18398,N_17906,N_17938);
and U18399 (N_18399,N_17901,N_17899);
and U18400 (N_18400,N_17993,N_18006);
and U18401 (N_18401,N_17587,N_17818);
xor U18402 (N_18402,N_17626,N_17502);
nor U18403 (N_18403,N_17585,N_17955);
or U18404 (N_18404,N_17775,N_17820);
or U18405 (N_18405,N_18111,N_17568);
and U18406 (N_18406,N_18045,N_17799);
nand U18407 (N_18407,N_17898,N_17924);
nand U18408 (N_18408,N_17835,N_17751);
nor U18409 (N_18409,N_17810,N_17783);
or U18410 (N_18410,N_18075,N_17705);
or U18411 (N_18411,N_17992,N_17798);
or U18412 (N_18412,N_17821,N_17696);
nor U18413 (N_18413,N_17651,N_17731);
and U18414 (N_18414,N_17746,N_17952);
nand U18415 (N_18415,N_17859,N_17904);
nor U18416 (N_18416,N_17645,N_17701);
or U18417 (N_18417,N_18098,N_17796);
or U18418 (N_18418,N_18005,N_17982);
and U18419 (N_18419,N_17665,N_17694);
nor U18420 (N_18420,N_17640,N_17989);
and U18421 (N_18421,N_18076,N_17544);
or U18422 (N_18422,N_17506,N_17944);
nor U18423 (N_18423,N_18070,N_17875);
and U18424 (N_18424,N_18015,N_17695);
or U18425 (N_18425,N_17726,N_17591);
xor U18426 (N_18426,N_18039,N_17574);
nor U18427 (N_18427,N_17586,N_17840);
nor U18428 (N_18428,N_17633,N_17763);
nand U18429 (N_18429,N_17872,N_17503);
or U18430 (N_18430,N_17929,N_17572);
nor U18431 (N_18431,N_17873,N_17902);
or U18432 (N_18432,N_17649,N_17613);
nand U18433 (N_18433,N_17504,N_17507);
nor U18434 (N_18434,N_18031,N_17805);
or U18435 (N_18435,N_17715,N_17500);
nor U18436 (N_18436,N_17631,N_17832);
nor U18437 (N_18437,N_17958,N_17831);
nand U18438 (N_18438,N_17770,N_18076);
xnor U18439 (N_18439,N_17585,N_17673);
xnor U18440 (N_18440,N_17766,N_17604);
nand U18441 (N_18441,N_17860,N_17947);
nand U18442 (N_18442,N_17961,N_17564);
or U18443 (N_18443,N_17878,N_18105);
nor U18444 (N_18444,N_17850,N_17729);
or U18445 (N_18445,N_17873,N_17849);
nor U18446 (N_18446,N_17553,N_17850);
nand U18447 (N_18447,N_17596,N_17672);
and U18448 (N_18448,N_17555,N_17784);
and U18449 (N_18449,N_17649,N_17539);
and U18450 (N_18450,N_18079,N_17656);
xor U18451 (N_18451,N_18097,N_17657);
and U18452 (N_18452,N_17761,N_17908);
nor U18453 (N_18453,N_17885,N_17745);
nor U18454 (N_18454,N_17935,N_17682);
or U18455 (N_18455,N_17845,N_17993);
nand U18456 (N_18456,N_17662,N_18019);
or U18457 (N_18457,N_17573,N_17666);
and U18458 (N_18458,N_18101,N_17703);
and U18459 (N_18459,N_17519,N_18052);
or U18460 (N_18460,N_17877,N_17568);
or U18461 (N_18461,N_17657,N_18065);
and U18462 (N_18462,N_17760,N_17871);
nor U18463 (N_18463,N_17708,N_17997);
nor U18464 (N_18464,N_17762,N_17642);
nor U18465 (N_18465,N_18005,N_17734);
or U18466 (N_18466,N_17754,N_17729);
or U18467 (N_18467,N_17877,N_17820);
nand U18468 (N_18468,N_17708,N_17845);
or U18469 (N_18469,N_17951,N_18123);
and U18470 (N_18470,N_17843,N_18033);
and U18471 (N_18471,N_18054,N_17880);
nand U18472 (N_18472,N_17860,N_17835);
and U18473 (N_18473,N_17634,N_17559);
or U18474 (N_18474,N_17954,N_17899);
nor U18475 (N_18475,N_17725,N_18084);
and U18476 (N_18476,N_17844,N_17641);
nor U18477 (N_18477,N_17958,N_17758);
or U18478 (N_18478,N_17821,N_18015);
or U18479 (N_18479,N_17565,N_17805);
nand U18480 (N_18480,N_17898,N_17710);
or U18481 (N_18481,N_17628,N_17933);
nor U18482 (N_18482,N_17611,N_17837);
or U18483 (N_18483,N_17551,N_17876);
xnor U18484 (N_18484,N_17797,N_17763);
or U18485 (N_18485,N_18024,N_17720);
nand U18486 (N_18486,N_17723,N_17977);
nor U18487 (N_18487,N_17736,N_17975);
or U18488 (N_18488,N_18031,N_17620);
or U18489 (N_18489,N_17503,N_17974);
and U18490 (N_18490,N_17910,N_18085);
nand U18491 (N_18491,N_17776,N_18086);
xnor U18492 (N_18492,N_17608,N_17784);
xor U18493 (N_18493,N_17803,N_17984);
and U18494 (N_18494,N_17863,N_17656);
or U18495 (N_18495,N_17766,N_17996);
nand U18496 (N_18496,N_17933,N_17916);
nand U18497 (N_18497,N_17863,N_17530);
and U18498 (N_18498,N_17821,N_17536);
or U18499 (N_18499,N_18074,N_18119);
nor U18500 (N_18500,N_17655,N_17521);
and U18501 (N_18501,N_17769,N_18050);
nand U18502 (N_18502,N_17834,N_17948);
and U18503 (N_18503,N_17709,N_17996);
and U18504 (N_18504,N_18058,N_17824);
xnor U18505 (N_18505,N_18008,N_17851);
nor U18506 (N_18506,N_17970,N_18091);
or U18507 (N_18507,N_17802,N_17695);
nand U18508 (N_18508,N_18017,N_17640);
or U18509 (N_18509,N_17957,N_17624);
nor U18510 (N_18510,N_17624,N_17630);
nor U18511 (N_18511,N_17868,N_17585);
nor U18512 (N_18512,N_17683,N_17641);
nand U18513 (N_18513,N_17920,N_17631);
nor U18514 (N_18514,N_17974,N_17748);
nor U18515 (N_18515,N_17760,N_17960);
nand U18516 (N_18516,N_17502,N_18042);
and U18517 (N_18517,N_17876,N_18110);
and U18518 (N_18518,N_17726,N_17559);
nor U18519 (N_18519,N_18039,N_17792);
nand U18520 (N_18520,N_17585,N_18088);
nand U18521 (N_18521,N_17542,N_17869);
and U18522 (N_18522,N_17964,N_18101);
or U18523 (N_18523,N_18073,N_17872);
xnor U18524 (N_18524,N_17939,N_17507);
and U18525 (N_18525,N_17859,N_18042);
nand U18526 (N_18526,N_17553,N_17801);
nand U18527 (N_18527,N_17501,N_17539);
nor U18528 (N_18528,N_17653,N_17759);
or U18529 (N_18529,N_18089,N_17743);
and U18530 (N_18530,N_17871,N_17819);
nand U18531 (N_18531,N_17587,N_18118);
nor U18532 (N_18532,N_17974,N_17834);
nand U18533 (N_18533,N_17959,N_17638);
nor U18534 (N_18534,N_17737,N_17848);
and U18535 (N_18535,N_17709,N_17949);
nor U18536 (N_18536,N_17998,N_17705);
nand U18537 (N_18537,N_17913,N_18080);
or U18538 (N_18538,N_17905,N_17514);
xnor U18539 (N_18539,N_17549,N_17897);
nor U18540 (N_18540,N_17594,N_17722);
nor U18541 (N_18541,N_18068,N_17707);
nand U18542 (N_18542,N_17882,N_17670);
nand U18543 (N_18543,N_17537,N_17641);
nand U18544 (N_18544,N_17578,N_17625);
or U18545 (N_18545,N_17706,N_17516);
or U18546 (N_18546,N_17943,N_17694);
and U18547 (N_18547,N_17924,N_17566);
or U18548 (N_18548,N_17595,N_17942);
nor U18549 (N_18549,N_18069,N_17708);
nor U18550 (N_18550,N_18030,N_17726);
nand U18551 (N_18551,N_17576,N_17789);
nor U18552 (N_18552,N_17699,N_17776);
or U18553 (N_18553,N_17618,N_17883);
and U18554 (N_18554,N_17536,N_17988);
xor U18555 (N_18555,N_18004,N_17991);
or U18556 (N_18556,N_17878,N_18106);
or U18557 (N_18557,N_17973,N_18013);
or U18558 (N_18558,N_17921,N_17934);
nand U18559 (N_18559,N_17677,N_17649);
or U18560 (N_18560,N_17518,N_17899);
nand U18561 (N_18561,N_17535,N_17788);
and U18562 (N_18562,N_18074,N_17977);
nor U18563 (N_18563,N_17576,N_18122);
nand U18564 (N_18564,N_18090,N_18118);
and U18565 (N_18565,N_17946,N_17539);
xor U18566 (N_18566,N_17952,N_18019);
nor U18567 (N_18567,N_17676,N_17621);
and U18568 (N_18568,N_17815,N_17772);
or U18569 (N_18569,N_17822,N_17598);
and U18570 (N_18570,N_18123,N_17966);
nand U18571 (N_18571,N_18090,N_17969);
xor U18572 (N_18572,N_17827,N_17839);
nor U18573 (N_18573,N_17503,N_17993);
and U18574 (N_18574,N_17708,N_17558);
or U18575 (N_18575,N_17632,N_17957);
xor U18576 (N_18576,N_17665,N_17670);
nand U18577 (N_18577,N_17644,N_17618);
and U18578 (N_18578,N_17706,N_17840);
nor U18579 (N_18579,N_17729,N_17974);
nand U18580 (N_18580,N_17527,N_17750);
xnor U18581 (N_18581,N_17578,N_17680);
nor U18582 (N_18582,N_18055,N_17531);
and U18583 (N_18583,N_18082,N_17817);
nand U18584 (N_18584,N_17716,N_18009);
and U18585 (N_18585,N_17953,N_17960);
nand U18586 (N_18586,N_17712,N_17650);
nand U18587 (N_18587,N_18107,N_17646);
or U18588 (N_18588,N_18076,N_17819);
xnor U18589 (N_18589,N_17891,N_18016);
and U18590 (N_18590,N_17823,N_17578);
xor U18591 (N_18591,N_17995,N_17786);
nor U18592 (N_18592,N_18040,N_18045);
or U18593 (N_18593,N_17632,N_17823);
nor U18594 (N_18594,N_17910,N_18002);
nor U18595 (N_18595,N_18080,N_17793);
xor U18596 (N_18596,N_18011,N_17745);
xor U18597 (N_18597,N_17571,N_17597);
nand U18598 (N_18598,N_18084,N_17862);
xor U18599 (N_18599,N_17825,N_17915);
nand U18600 (N_18600,N_17831,N_17994);
nor U18601 (N_18601,N_18105,N_17677);
nand U18602 (N_18602,N_17819,N_17663);
and U18603 (N_18603,N_17827,N_17577);
nor U18604 (N_18604,N_17760,N_17552);
nor U18605 (N_18605,N_18096,N_17716);
and U18606 (N_18606,N_18118,N_17998);
and U18607 (N_18607,N_17796,N_18095);
and U18608 (N_18608,N_17612,N_18001);
and U18609 (N_18609,N_17612,N_17958);
nand U18610 (N_18610,N_17534,N_17764);
and U18611 (N_18611,N_17998,N_17775);
and U18612 (N_18612,N_17725,N_17994);
nor U18613 (N_18613,N_17967,N_17535);
or U18614 (N_18614,N_17559,N_17656);
or U18615 (N_18615,N_17898,N_17643);
and U18616 (N_18616,N_17942,N_17568);
or U18617 (N_18617,N_17601,N_17611);
nand U18618 (N_18618,N_17952,N_17797);
and U18619 (N_18619,N_17599,N_17668);
and U18620 (N_18620,N_17698,N_17516);
nand U18621 (N_18621,N_17510,N_17621);
and U18622 (N_18622,N_18041,N_17586);
or U18623 (N_18623,N_17828,N_17647);
nor U18624 (N_18624,N_17652,N_17936);
and U18625 (N_18625,N_17890,N_17936);
nor U18626 (N_18626,N_17683,N_17854);
nor U18627 (N_18627,N_17884,N_17750);
and U18628 (N_18628,N_17626,N_18013);
nor U18629 (N_18629,N_18055,N_17601);
xnor U18630 (N_18630,N_17788,N_17779);
or U18631 (N_18631,N_17668,N_18085);
nor U18632 (N_18632,N_17942,N_17792);
nand U18633 (N_18633,N_18017,N_17661);
and U18634 (N_18634,N_17835,N_17729);
and U18635 (N_18635,N_17859,N_17534);
nand U18636 (N_18636,N_17865,N_17755);
nor U18637 (N_18637,N_17648,N_17530);
nand U18638 (N_18638,N_17675,N_17860);
and U18639 (N_18639,N_17674,N_17707);
and U18640 (N_18640,N_18098,N_18085);
nand U18641 (N_18641,N_17793,N_17934);
and U18642 (N_18642,N_18094,N_17525);
nand U18643 (N_18643,N_17755,N_17553);
or U18644 (N_18644,N_17627,N_17948);
nand U18645 (N_18645,N_17743,N_18037);
and U18646 (N_18646,N_17608,N_17757);
nand U18647 (N_18647,N_17601,N_17639);
and U18648 (N_18648,N_17899,N_17971);
nand U18649 (N_18649,N_17793,N_17770);
nand U18650 (N_18650,N_17942,N_18117);
xnor U18651 (N_18651,N_17868,N_18087);
and U18652 (N_18652,N_17594,N_17815);
or U18653 (N_18653,N_18034,N_17767);
and U18654 (N_18654,N_17732,N_18092);
nor U18655 (N_18655,N_18099,N_17665);
xor U18656 (N_18656,N_17791,N_17829);
xor U18657 (N_18657,N_17760,N_17531);
nor U18658 (N_18658,N_17860,N_17572);
nor U18659 (N_18659,N_17687,N_18099);
and U18660 (N_18660,N_17750,N_17522);
nor U18661 (N_18661,N_17693,N_18093);
nor U18662 (N_18662,N_17751,N_17971);
nand U18663 (N_18663,N_17529,N_17831);
nor U18664 (N_18664,N_17942,N_17943);
nor U18665 (N_18665,N_18010,N_17757);
and U18666 (N_18666,N_17831,N_17987);
nand U18667 (N_18667,N_17817,N_17664);
or U18668 (N_18668,N_17803,N_17867);
and U18669 (N_18669,N_18080,N_17803);
or U18670 (N_18670,N_18102,N_17640);
and U18671 (N_18671,N_17756,N_17621);
nand U18672 (N_18672,N_17750,N_17517);
xnor U18673 (N_18673,N_17900,N_18104);
and U18674 (N_18674,N_17532,N_17810);
or U18675 (N_18675,N_17691,N_17633);
or U18676 (N_18676,N_17918,N_17743);
nand U18677 (N_18677,N_17709,N_17561);
nor U18678 (N_18678,N_17726,N_17787);
nor U18679 (N_18679,N_17724,N_18109);
and U18680 (N_18680,N_17799,N_17594);
or U18681 (N_18681,N_17762,N_17705);
nor U18682 (N_18682,N_17830,N_17866);
nor U18683 (N_18683,N_17718,N_17661);
or U18684 (N_18684,N_17503,N_17533);
or U18685 (N_18685,N_17629,N_17615);
and U18686 (N_18686,N_17631,N_17948);
nor U18687 (N_18687,N_18033,N_17641);
xor U18688 (N_18688,N_17533,N_17600);
nand U18689 (N_18689,N_17519,N_18117);
or U18690 (N_18690,N_17868,N_17721);
and U18691 (N_18691,N_17656,N_17857);
and U18692 (N_18692,N_17849,N_17503);
nor U18693 (N_18693,N_18120,N_18099);
or U18694 (N_18694,N_17870,N_18025);
and U18695 (N_18695,N_17954,N_17696);
nor U18696 (N_18696,N_18075,N_17861);
nand U18697 (N_18697,N_18028,N_17511);
and U18698 (N_18698,N_18067,N_17690);
or U18699 (N_18699,N_17816,N_17665);
xor U18700 (N_18700,N_17889,N_17709);
nand U18701 (N_18701,N_17720,N_17607);
nor U18702 (N_18702,N_18100,N_18056);
and U18703 (N_18703,N_17788,N_17840);
and U18704 (N_18704,N_17827,N_17547);
and U18705 (N_18705,N_18076,N_18114);
and U18706 (N_18706,N_17807,N_17752);
and U18707 (N_18707,N_17665,N_17585);
and U18708 (N_18708,N_17762,N_17576);
and U18709 (N_18709,N_17890,N_18101);
nand U18710 (N_18710,N_17898,N_17988);
xnor U18711 (N_18711,N_17844,N_17625);
nand U18712 (N_18712,N_17793,N_17582);
nor U18713 (N_18713,N_17968,N_18117);
or U18714 (N_18714,N_18071,N_17581);
and U18715 (N_18715,N_18021,N_17902);
nor U18716 (N_18716,N_18059,N_17774);
and U18717 (N_18717,N_17749,N_17877);
or U18718 (N_18718,N_17764,N_17500);
and U18719 (N_18719,N_17682,N_17734);
nand U18720 (N_18720,N_17758,N_18056);
nand U18721 (N_18721,N_18040,N_18108);
nand U18722 (N_18722,N_17568,N_17584);
nand U18723 (N_18723,N_18073,N_17500);
nor U18724 (N_18724,N_17906,N_17574);
nor U18725 (N_18725,N_18123,N_17622);
and U18726 (N_18726,N_18001,N_17994);
and U18727 (N_18727,N_17867,N_18009);
nand U18728 (N_18728,N_17546,N_17766);
nand U18729 (N_18729,N_18117,N_17903);
nor U18730 (N_18730,N_17943,N_17734);
nor U18731 (N_18731,N_17599,N_18088);
or U18732 (N_18732,N_17562,N_17816);
xor U18733 (N_18733,N_17991,N_18013);
nand U18734 (N_18734,N_17982,N_17842);
or U18735 (N_18735,N_17703,N_17845);
or U18736 (N_18736,N_17988,N_17551);
nor U18737 (N_18737,N_17866,N_17732);
and U18738 (N_18738,N_17689,N_17732);
nand U18739 (N_18739,N_17694,N_17554);
nor U18740 (N_18740,N_17815,N_18077);
or U18741 (N_18741,N_17941,N_18068);
nand U18742 (N_18742,N_17972,N_17905);
nor U18743 (N_18743,N_17938,N_17865);
xnor U18744 (N_18744,N_17843,N_17551);
or U18745 (N_18745,N_18015,N_17788);
and U18746 (N_18746,N_17872,N_17947);
nor U18747 (N_18747,N_17775,N_17515);
or U18748 (N_18748,N_18089,N_17836);
and U18749 (N_18749,N_17857,N_17756);
or U18750 (N_18750,N_18231,N_18696);
and U18751 (N_18751,N_18338,N_18318);
nand U18752 (N_18752,N_18319,N_18547);
or U18753 (N_18753,N_18540,N_18498);
or U18754 (N_18754,N_18599,N_18604);
and U18755 (N_18755,N_18624,N_18437);
nor U18756 (N_18756,N_18476,N_18496);
or U18757 (N_18757,N_18595,N_18259);
nand U18758 (N_18758,N_18337,N_18233);
nor U18759 (N_18759,N_18166,N_18450);
and U18760 (N_18760,N_18683,N_18240);
or U18761 (N_18761,N_18179,N_18408);
or U18762 (N_18762,N_18130,N_18523);
and U18763 (N_18763,N_18584,N_18550);
nand U18764 (N_18764,N_18208,N_18570);
nor U18765 (N_18765,N_18325,N_18176);
or U18766 (N_18766,N_18499,N_18144);
and U18767 (N_18767,N_18341,N_18158);
and U18768 (N_18768,N_18588,N_18429);
nor U18769 (N_18769,N_18210,N_18578);
nand U18770 (N_18770,N_18185,N_18333);
or U18771 (N_18771,N_18435,N_18384);
or U18772 (N_18772,N_18258,N_18474);
xnor U18773 (N_18773,N_18676,N_18534);
or U18774 (N_18774,N_18321,N_18307);
and U18775 (N_18775,N_18261,N_18273);
nand U18776 (N_18776,N_18565,N_18665);
nor U18777 (N_18777,N_18541,N_18555);
nand U18778 (N_18778,N_18316,N_18711);
nand U18779 (N_18779,N_18682,N_18377);
and U18780 (N_18780,N_18157,N_18740);
nand U18781 (N_18781,N_18481,N_18618);
or U18782 (N_18782,N_18658,N_18277);
or U18783 (N_18783,N_18141,N_18546);
or U18784 (N_18784,N_18434,N_18440);
nand U18785 (N_18785,N_18242,N_18544);
or U18786 (N_18786,N_18661,N_18276);
nand U18787 (N_18787,N_18287,N_18553);
nand U18788 (N_18788,N_18371,N_18386);
nand U18789 (N_18789,N_18198,N_18397);
nor U18790 (N_18790,N_18416,N_18573);
and U18791 (N_18791,N_18712,N_18394);
or U18792 (N_18792,N_18274,N_18525);
and U18793 (N_18793,N_18359,N_18520);
and U18794 (N_18794,N_18691,N_18640);
nand U18795 (N_18795,N_18404,N_18267);
nor U18796 (N_18796,N_18326,N_18657);
and U18797 (N_18797,N_18485,N_18471);
and U18798 (N_18798,N_18514,N_18656);
xor U18799 (N_18799,N_18597,N_18494);
nor U18800 (N_18800,N_18497,N_18687);
and U18801 (N_18801,N_18366,N_18428);
and U18802 (N_18802,N_18165,N_18549);
xor U18803 (N_18803,N_18167,N_18625);
or U18804 (N_18804,N_18355,N_18343);
nand U18805 (N_18805,N_18344,N_18279);
nand U18806 (N_18806,N_18432,N_18635);
or U18807 (N_18807,N_18126,N_18317);
and U18808 (N_18808,N_18479,N_18666);
nor U18809 (N_18809,N_18225,N_18154);
and U18810 (N_18810,N_18306,N_18678);
nor U18811 (N_18811,N_18142,N_18655);
or U18812 (N_18812,N_18207,N_18572);
and U18813 (N_18813,N_18419,N_18327);
nand U18814 (N_18814,N_18294,N_18241);
or U18815 (N_18815,N_18293,N_18695);
nor U18816 (N_18816,N_18304,N_18168);
and U18817 (N_18817,N_18732,N_18462);
nand U18818 (N_18818,N_18405,N_18707);
nor U18819 (N_18819,N_18467,N_18155);
xor U18820 (N_18820,N_18622,N_18517);
and U18821 (N_18821,N_18455,N_18127);
and U18822 (N_18822,N_18390,N_18605);
nor U18823 (N_18823,N_18477,N_18160);
and U18824 (N_18824,N_18470,N_18391);
xor U18825 (N_18825,N_18353,N_18367);
nor U18826 (N_18826,N_18564,N_18690);
nand U18827 (N_18827,N_18634,N_18215);
nand U18828 (N_18828,N_18131,N_18576);
nand U18829 (N_18829,N_18369,N_18509);
or U18830 (N_18830,N_18269,N_18719);
and U18831 (N_18831,N_18406,N_18463);
xor U18832 (N_18832,N_18686,N_18430);
nand U18833 (N_18833,N_18177,N_18521);
and U18834 (N_18834,N_18340,N_18352);
or U18835 (N_18835,N_18164,N_18370);
or U18836 (N_18836,N_18201,N_18156);
xor U18837 (N_18837,N_18161,N_18254);
and U18838 (N_18838,N_18146,N_18381);
or U18839 (N_18839,N_18420,N_18291);
nand U18840 (N_18840,N_18645,N_18689);
nand U18841 (N_18841,N_18280,N_18680);
and U18842 (N_18842,N_18409,N_18171);
nand U18843 (N_18843,N_18735,N_18412);
nand U18844 (N_18844,N_18533,N_18720);
and U18845 (N_18845,N_18673,N_18558);
and U18846 (N_18846,N_18217,N_18646);
or U18847 (N_18847,N_18310,N_18556);
nand U18848 (N_18848,N_18378,N_18290);
nor U18849 (N_18849,N_18191,N_18539);
nor U18850 (N_18850,N_18357,N_18305);
nand U18851 (N_18851,N_18222,N_18348);
nand U18852 (N_18852,N_18422,N_18251);
nand U18853 (N_18853,N_18385,N_18328);
and U18854 (N_18854,N_18503,N_18452);
xnor U18855 (N_18855,N_18211,N_18436);
xor U18856 (N_18856,N_18180,N_18414);
nand U18857 (N_18857,N_18139,N_18322);
or U18858 (N_18858,N_18175,N_18163);
or U18859 (N_18859,N_18232,N_18528);
nand U18860 (N_18860,N_18182,N_18392);
and U18861 (N_18861,N_18728,N_18616);
nand U18862 (N_18862,N_18505,N_18739);
or U18863 (N_18863,N_18363,N_18303);
and U18864 (N_18864,N_18465,N_18302);
and U18865 (N_18865,N_18454,N_18490);
and U18866 (N_18866,N_18598,N_18609);
and U18867 (N_18867,N_18668,N_18246);
and U18868 (N_18868,N_18135,N_18698);
nand U18869 (N_18869,N_18425,N_18538);
and U18870 (N_18870,N_18608,N_18580);
or U18871 (N_18871,N_18714,N_18472);
xnor U18872 (N_18872,N_18263,N_18372);
xnor U18873 (N_18873,N_18438,N_18650);
or U18874 (N_18874,N_18250,N_18361);
and U18875 (N_18875,N_18443,N_18324);
xor U18876 (N_18876,N_18684,N_18214);
nor U18877 (N_18877,N_18330,N_18364);
and U18878 (N_18878,N_18351,N_18747);
and U18879 (N_18879,N_18284,N_18134);
xor U18880 (N_18880,N_18445,N_18563);
or U18881 (N_18881,N_18532,N_18663);
nand U18882 (N_18882,N_18143,N_18522);
nand U18883 (N_18883,N_18519,N_18295);
or U18884 (N_18884,N_18733,N_18209);
or U18885 (N_18885,N_18239,N_18213);
and U18886 (N_18886,N_18138,N_18697);
nand U18887 (N_18887,N_18268,N_18694);
or U18888 (N_18888,N_18632,N_18265);
or U18889 (N_18889,N_18526,N_18506);
nor U18890 (N_18890,N_18483,N_18568);
nand U18891 (N_18891,N_18283,N_18706);
nor U18892 (N_18892,N_18623,N_18145);
xnor U18893 (N_18893,N_18648,N_18426);
xor U18894 (N_18894,N_18196,N_18542);
or U18895 (N_18895,N_18644,N_18486);
nand U18896 (N_18896,N_18281,N_18571);
nand U18897 (N_18897,N_18466,N_18730);
nand U18898 (N_18898,N_18181,N_18475);
and U18899 (N_18899,N_18137,N_18488);
or U18900 (N_18900,N_18252,N_18199);
nand U18901 (N_18901,N_18189,N_18212);
and U18902 (N_18902,N_18688,N_18518);
or U18903 (N_18903,N_18524,N_18221);
nor U18904 (N_18904,N_18621,N_18243);
and U18905 (N_18905,N_18692,N_18413);
and U18906 (N_18906,N_18672,N_18504);
nand U18907 (N_18907,N_18551,N_18235);
nor U18908 (N_18908,N_18264,N_18626);
nor U18909 (N_18909,N_18271,N_18446);
and U18910 (N_18910,N_18654,N_18169);
and U18911 (N_18911,N_18257,N_18742);
and U18912 (N_18912,N_18734,N_18407);
and U18913 (N_18913,N_18427,N_18502);
and U18914 (N_18914,N_18671,N_18448);
or U18915 (N_18915,N_18724,N_18223);
nand U18916 (N_18916,N_18238,N_18636);
xor U18917 (N_18917,N_18537,N_18190);
and U18918 (N_18918,N_18299,N_18423);
and U18919 (N_18919,N_18587,N_18218);
nand U18920 (N_18920,N_18628,N_18285);
or U18921 (N_18921,N_18260,N_18743);
nand U18922 (N_18922,N_18469,N_18458);
and U18923 (N_18923,N_18402,N_18708);
nor U18924 (N_18924,N_18703,N_18301);
nor U18925 (N_18925,N_18721,N_18178);
or U18926 (N_18926,N_18275,N_18444);
or U18927 (N_18927,N_18399,N_18629);
nor U18928 (N_18928,N_18482,N_18334);
and U18929 (N_18929,N_18320,N_18216);
nor U18930 (N_18930,N_18748,N_18511);
nand U18931 (N_18931,N_18375,N_18585);
nor U18932 (N_18932,N_18230,N_18718);
nand U18933 (N_18933,N_18709,N_18659);
xnor U18934 (N_18934,N_18453,N_18187);
and U18935 (N_18935,N_18495,N_18675);
xnor U18936 (N_18936,N_18559,N_18569);
and U18937 (N_18937,N_18726,N_18159);
xor U18938 (N_18938,N_18693,N_18172);
or U18939 (N_18939,N_18148,N_18174);
nor U18940 (N_18940,N_18567,N_18744);
and U18941 (N_18941,N_18581,N_18312);
nor U18942 (N_18942,N_18630,N_18219);
nand U18943 (N_18943,N_18329,N_18561);
nand U18944 (N_18944,N_18677,N_18236);
nor U18945 (N_18945,N_18610,N_18459);
or U18946 (N_18946,N_18194,N_18704);
or U18947 (N_18947,N_18162,N_18237);
or U18948 (N_18948,N_18492,N_18638);
nand U18949 (N_18949,N_18323,N_18383);
nand U18950 (N_18950,N_18468,N_18746);
xor U18951 (N_18951,N_18461,N_18449);
xnor U18952 (N_18952,N_18292,N_18653);
and U18953 (N_18953,N_18373,N_18244);
or U18954 (N_18954,N_18639,N_18128);
nand U18955 (N_18955,N_18380,N_18331);
nand U18956 (N_18956,N_18620,N_18226);
and U18957 (N_18957,N_18699,N_18195);
or U18958 (N_18958,N_18335,N_18560);
nor U18959 (N_18959,N_18202,N_18360);
nor U18960 (N_18960,N_18308,N_18535);
and U18961 (N_18961,N_18667,N_18637);
nand U18962 (N_18962,N_18633,N_18229);
xnor U18963 (N_18963,N_18586,N_18149);
xor U18964 (N_18964,N_18562,N_18421);
xnor U18965 (N_18965,N_18262,N_18715);
or U18966 (N_18966,N_18593,N_18660);
nand U18967 (N_18967,N_18669,N_18702);
and U18968 (N_18968,N_18332,N_18354);
or U18969 (N_18969,N_18206,N_18342);
and U18970 (N_18970,N_18297,N_18345);
nor U18971 (N_18971,N_18200,N_18309);
nand U18972 (N_18972,N_18582,N_18140);
nor U18973 (N_18973,N_18717,N_18286);
nand U18974 (N_18974,N_18311,N_18530);
or U18975 (N_18975,N_18651,N_18515);
nand U18976 (N_18976,N_18603,N_18513);
nor U18977 (N_18977,N_18460,N_18531);
nor U18978 (N_18978,N_18220,N_18395);
or U18979 (N_18979,N_18376,N_18125);
or U18980 (N_18980,N_18374,N_18315);
nor U18981 (N_18981,N_18255,N_18478);
nand U18982 (N_18982,N_18670,N_18396);
or U18983 (N_18983,N_18431,N_18614);
and U18984 (N_18984,N_18619,N_18249);
and U18985 (N_18985,N_18288,N_18133);
and U18986 (N_18986,N_18701,N_18457);
and U18987 (N_18987,N_18184,N_18183);
nor U18988 (N_18988,N_18664,N_18188);
nand U18989 (N_18989,N_18234,N_18617);
nor U18990 (N_18990,N_18681,N_18674);
or U18991 (N_18991,N_18480,N_18282);
nor U18992 (N_18992,N_18245,N_18379);
xor U18993 (N_18993,N_18193,N_18508);
nor U18994 (N_18994,N_18596,N_18389);
nand U18995 (N_18995,N_18387,N_18347);
nand U18996 (N_18996,N_18574,N_18545);
or U18997 (N_18997,N_18170,N_18197);
or U18998 (N_18998,N_18247,N_18451);
nor U18999 (N_18999,N_18579,N_18615);
nand U19000 (N_19000,N_18132,N_18716);
nor U19001 (N_19001,N_18415,N_18649);
nand U19002 (N_19002,N_18442,N_18516);
and U19003 (N_19003,N_18253,N_18652);
nor U19004 (N_19004,N_18362,N_18749);
and U19005 (N_19005,N_18512,N_18129);
nor U19006 (N_19006,N_18152,N_18313);
xor U19007 (N_19007,N_18205,N_18662);
nor U19008 (N_19008,N_18501,N_18418);
nor U19009 (N_19009,N_18248,N_18358);
xnor U19010 (N_19010,N_18401,N_18601);
or U19011 (N_19011,N_18592,N_18685);
nand U19012 (N_19012,N_18627,N_18289);
xnor U19013 (N_19013,N_18433,N_18710);
and U19014 (N_19014,N_18613,N_18737);
xor U19015 (N_19015,N_18741,N_18487);
nor U19016 (N_19016,N_18186,N_18543);
or U19017 (N_19017,N_18228,N_18300);
and U19018 (N_19018,N_18424,N_18473);
xnor U19019 (N_19019,N_18256,N_18529);
and U19020 (N_19020,N_18705,N_18439);
and U19021 (N_19021,N_18410,N_18548);
or U19022 (N_19022,N_18566,N_18417);
nor U19023 (N_19023,N_18722,N_18602);
nor U19024 (N_19024,N_18270,N_18493);
and U19025 (N_19025,N_18679,N_18204);
nand U19026 (N_19026,N_18607,N_18552);
or U19027 (N_19027,N_18136,N_18725);
or U19028 (N_19028,N_18349,N_18278);
and U19029 (N_19029,N_18557,N_18382);
nand U19030 (N_19030,N_18575,N_18173);
and U19031 (N_19031,N_18727,N_18203);
or U19032 (N_19032,N_18510,N_18700);
and U19033 (N_19033,N_18314,N_18224);
or U19034 (N_19034,N_18729,N_18600);
or U19035 (N_19035,N_18272,N_18464);
or U19036 (N_19036,N_18356,N_18350);
or U19037 (N_19037,N_18365,N_18642);
and U19038 (N_19038,N_18456,N_18594);
nor U19039 (N_19039,N_18192,N_18398);
or U19040 (N_19040,N_18489,N_18441);
nand U19041 (N_19041,N_18536,N_18577);
nor U19042 (N_19042,N_18151,N_18411);
or U19043 (N_19043,N_18393,N_18713);
nand U19044 (N_19044,N_18336,N_18736);
and U19045 (N_19045,N_18368,N_18647);
nor U19046 (N_19046,N_18298,N_18500);
and U19047 (N_19047,N_18589,N_18346);
nand U19048 (N_19048,N_18296,N_18227);
nand U19049 (N_19049,N_18400,N_18339);
or U19050 (N_19050,N_18745,N_18723);
or U19051 (N_19051,N_18388,N_18507);
nand U19052 (N_19052,N_18591,N_18150);
and U19053 (N_19053,N_18147,N_18643);
and U19054 (N_19054,N_18527,N_18611);
nand U19055 (N_19055,N_18731,N_18153);
and U19056 (N_19056,N_18447,N_18403);
nor U19057 (N_19057,N_18641,N_18606);
nand U19058 (N_19058,N_18631,N_18590);
and U19059 (N_19059,N_18554,N_18484);
nor U19060 (N_19060,N_18738,N_18266);
xnor U19061 (N_19061,N_18583,N_18491);
or U19062 (N_19062,N_18612,N_18591);
nor U19063 (N_19063,N_18126,N_18464);
and U19064 (N_19064,N_18538,N_18464);
or U19065 (N_19065,N_18363,N_18512);
and U19066 (N_19066,N_18675,N_18139);
nand U19067 (N_19067,N_18685,N_18262);
nand U19068 (N_19068,N_18223,N_18396);
nor U19069 (N_19069,N_18285,N_18505);
or U19070 (N_19070,N_18167,N_18438);
and U19071 (N_19071,N_18567,N_18507);
or U19072 (N_19072,N_18463,N_18175);
nor U19073 (N_19073,N_18388,N_18525);
nor U19074 (N_19074,N_18571,N_18165);
and U19075 (N_19075,N_18724,N_18325);
or U19076 (N_19076,N_18144,N_18222);
nor U19077 (N_19077,N_18613,N_18410);
and U19078 (N_19078,N_18590,N_18176);
nand U19079 (N_19079,N_18548,N_18712);
nor U19080 (N_19080,N_18222,N_18426);
nor U19081 (N_19081,N_18357,N_18500);
nor U19082 (N_19082,N_18155,N_18290);
nor U19083 (N_19083,N_18532,N_18596);
or U19084 (N_19084,N_18256,N_18324);
and U19085 (N_19085,N_18590,N_18327);
nor U19086 (N_19086,N_18617,N_18337);
xor U19087 (N_19087,N_18672,N_18346);
nor U19088 (N_19088,N_18621,N_18229);
nand U19089 (N_19089,N_18187,N_18738);
or U19090 (N_19090,N_18371,N_18570);
or U19091 (N_19091,N_18135,N_18190);
and U19092 (N_19092,N_18154,N_18730);
or U19093 (N_19093,N_18539,N_18670);
nor U19094 (N_19094,N_18329,N_18510);
nor U19095 (N_19095,N_18737,N_18440);
xnor U19096 (N_19096,N_18456,N_18411);
nand U19097 (N_19097,N_18468,N_18360);
nand U19098 (N_19098,N_18524,N_18615);
nand U19099 (N_19099,N_18449,N_18148);
and U19100 (N_19100,N_18563,N_18508);
xor U19101 (N_19101,N_18125,N_18430);
nand U19102 (N_19102,N_18553,N_18444);
nor U19103 (N_19103,N_18608,N_18573);
xnor U19104 (N_19104,N_18415,N_18402);
nand U19105 (N_19105,N_18415,N_18513);
nor U19106 (N_19106,N_18392,N_18527);
nand U19107 (N_19107,N_18565,N_18574);
or U19108 (N_19108,N_18340,N_18231);
nand U19109 (N_19109,N_18694,N_18338);
and U19110 (N_19110,N_18706,N_18248);
or U19111 (N_19111,N_18243,N_18342);
or U19112 (N_19112,N_18743,N_18168);
or U19113 (N_19113,N_18191,N_18637);
and U19114 (N_19114,N_18367,N_18142);
nor U19115 (N_19115,N_18572,N_18621);
nor U19116 (N_19116,N_18129,N_18262);
xnor U19117 (N_19117,N_18458,N_18635);
nand U19118 (N_19118,N_18654,N_18401);
nor U19119 (N_19119,N_18399,N_18394);
nand U19120 (N_19120,N_18749,N_18569);
xor U19121 (N_19121,N_18326,N_18285);
nor U19122 (N_19122,N_18615,N_18277);
or U19123 (N_19123,N_18749,N_18460);
or U19124 (N_19124,N_18128,N_18720);
and U19125 (N_19125,N_18355,N_18654);
xnor U19126 (N_19126,N_18327,N_18721);
nand U19127 (N_19127,N_18541,N_18685);
nand U19128 (N_19128,N_18125,N_18178);
xnor U19129 (N_19129,N_18136,N_18149);
nor U19130 (N_19130,N_18154,N_18306);
or U19131 (N_19131,N_18593,N_18381);
or U19132 (N_19132,N_18359,N_18637);
nand U19133 (N_19133,N_18468,N_18313);
nand U19134 (N_19134,N_18628,N_18367);
xnor U19135 (N_19135,N_18445,N_18520);
and U19136 (N_19136,N_18437,N_18563);
nor U19137 (N_19137,N_18585,N_18383);
nand U19138 (N_19138,N_18700,N_18334);
or U19139 (N_19139,N_18224,N_18520);
xor U19140 (N_19140,N_18203,N_18240);
and U19141 (N_19141,N_18412,N_18451);
nor U19142 (N_19142,N_18369,N_18336);
nand U19143 (N_19143,N_18605,N_18685);
xnor U19144 (N_19144,N_18543,N_18579);
nor U19145 (N_19145,N_18491,N_18364);
and U19146 (N_19146,N_18311,N_18506);
nor U19147 (N_19147,N_18212,N_18647);
or U19148 (N_19148,N_18417,N_18213);
or U19149 (N_19149,N_18676,N_18385);
nand U19150 (N_19150,N_18640,N_18583);
or U19151 (N_19151,N_18730,N_18449);
and U19152 (N_19152,N_18624,N_18527);
or U19153 (N_19153,N_18745,N_18336);
nor U19154 (N_19154,N_18143,N_18664);
or U19155 (N_19155,N_18518,N_18465);
nand U19156 (N_19156,N_18288,N_18397);
and U19157 (N_19157,N_18140,N_18680);
nand U19158 (N_19158,N_18518,N_18682);
or U19159 (N_19159,N_18642,N_18620);
nor U19160 (N_19160,N_18595,N_18673);
xor U19161 (N_19161,N_18637,N_18663);
xnor U19162 (N_19162,N_18152,N_18469);
or U19163 (N_19163,N_18434,N_18363);
or U19164 (N_19164,N_18518,N_18632);
and U19165 (N_19165,N_18622,N_18227);
or U19166 (N_19166,N_18747,N_18570);
xnor U19167 (N_19167,N_18398,N_18681);
nor U19168 (N_19168,N_18634,N_18422);
nand U19169 (N_19169,N_18414,N_18413);
nand U19170 (N_19170,N_18313,N_18348);
nand U19171 (N_19171,N_18185,N_18499);
or U19172 (N_19172,N_18735,N_18404);
and U19173 (N_19173,N_18307,N_18453);
or U19174 (N_19174,N_18165,N_18513);
xnor U19175 (N_19175,N_18142,N_18264);
nor U19176 (N_19176,N_18578,N_18442);
and U19177 (N_19177,N_18156,N_18446);
or U19178 (N_19178,N_18189,N_18648);
and U19179 (N_19179,N_18255,N_18186);
nor U19180 (N_19180,N_18157,N_18703);
nor U19181 (N_19181,N_18567,N_18557);
nor U19182 (N_19182,N_18343,N_18239);
and U19183 (N_19183,N_18356,N_18398);
and U19184 (N_19184,N_18272,N_18240);
nor U19185 (N_19185,N_18205,N_18158);
nor U19186 (N_19186,N_18664,N_18646);
or U19187 (N_19187,N_18593,N_18310);
xnor U19188 (N_19188,N_18453,N_18543);
or U19189 (N_19189,N_18590,N_18142);
nor U19190 (N_19190,N_18313,N_18370);
and U19191 (N_19191,N_18339,N_18449);
or U19192 (N_19192,N_18136,N_18281);
and U19193 (N_19193,N_18749,N_18389);
nand U19194 (N_19194,N_18419,N_18496);
and U19195 (N_19195,N_18378,N_18587);
nor U19196 (N_19196,N_18684,N_18304);
or U19197 (N_19197,N_18220,N_18312);
nand U19198 (N_19198,N_18677,N_18747);
and U19199 (N_19199,N_18332,N_18540);
and U19200 (N_19200,N_18321,N_18527);
nand U19201 (N_19201,N_18139,N_18248);
nor U19202 (N_19202,N_18508,N_18317);
xor U19203 (N_19203,N_18150,N_18289);
or U19204 (N_19204,N_18545,N_18539);
nor U19205 (N_19205,N_18404,N_18420);
or U19206 (N_19206,N_18490,N_18166);
or U19207 (N_19207,N_18528,N_18167);
nor U19208 (N_19208,N_18371,N_18475);
nor U19209 (N_19209,N_18179,N_18329);
nor U19210 (N_19210,N_18614,N_18200);
nand U19211 (N_19211,N_18214,N_18183);
nor U19212 (N_19212,N_18145,N_18412);
nor U19213 (N_19213,N_18672,N_18220);
nor U19214 (N_19214,N_18265,N_18443);
nor U19215 (N_19215,N_18745,N_18633);
or U19216 (N_19216,N_18198,N_18245);
xor U19217 (N_19217,N_18335,N_18551);
nand U19218 (N_19218,N_18606,N_18447);
nor U19219 (N_19219,N_18193,N_18143);
nor U19220 (N_19220,N_18638,N_18446);
and U19221 (N_19221,N_18625,N_18571);
or U19222 (N_19222,N_18127,N_18232);
or U19223 (N_19223,N_18369,N_18620);
nand U19224 (N_19224,N_18515,N_18143);
or U19225 (N_19225,N_18639,N_18518);
nor U19226 (N_19226,N_18736,N_18671);
nor U19227 (N_19227,N_18211,N_18698);
and U19228 (N_19228,N_18744,N_18674);
xor U19229 (N_19229,N_18621,N_18155);
nand U19230 (N_19230,N_18412,N_18410);
nand U19231 (N_19231,N_18565,N_18294);
nor U19232 (N_19232,N_18293,N_18687);
and U19233 (N_19233,N_18529,N_18403);
or U19234 (N_19234,N_18504,N_18480);
xnor U19235 (N_19235,N_18342,N_18601);
nand U19236 (N_19236,N_18230,N_18707);
and U19237 (N_19237,N_18485,N_18663);
nor U19238 (N_19238,N_18631,N_18205);
nor U19239 (N_19239,N_18699,N_18622);
or U19240 (N_19240,N_18263,N_18578);
nor U19241 (N_19241,N_18709,N_18328);
or U19242 (N_19242,N_18371,N_18334);
nor U19243 (N_19243,N_18516,N_18642);
nand U19244 (N_19244,N_18287,N_18165);
and U19245 (N_19245,N_18502,N_18694);
nor U19246 (N_19246,N_18612,N_18635);
nand U19247 (N_19247,N_18748,N_18691);
nand U19248 (N_19248,N_18511,N_18670);
and U19249 (N_19249,N_18371,N_18262);
nand U19250 (N_19250,N_18494,N_18546);
nand U19251 (N_19251,N_18413,N_18387);
nor U19252 (N_19252,N_18411,N_18729);
or U19253 (N_19253,N_18424,N_18638);
nand U19254 (N_19254,N_18604,N_18378);
and U19255 (N_19255,N_18133,N_18175);
or U19256 (N_19256,N_18205,N_18484);
nor U19257 (N_19257,N_18404,N_18298);
or U19258 (N_19258,N_18545,N_18386);
nor U19259 (N_19259,N_18211,N_18523);
xor U19260 (N_19260,N_18184,N_18494);
nor U19261 (N_19261,N_18197,N_18126);
nor U19262 (N_19262,N_18535,N_18454);
nor U19263 (N_19263,N_18425,N_18382);
or U19264 (N_19264,N_18264,N_18373);
xnor U19265 (N_19265,N_18246,N_18571);
nand U19266 (N_19266,N_18363,N_18731);
or U19267 (N_19267,N_18402,N_18627);
nor U19268 (N_19268,N_18226,N_18738);
or U19269 (N_19269,N_18299,N_18267);
nand U19270 (N_19270,N_18348,N_18620);
nor U19271 (N_19271,N_18196,N_18390);
and U19272 (N_19272,N_18726,N_18589);
nor U19273 (N_19273,N_18453,N_18604);
nor U19274 (N_19274,N_18676,N_18245);
and U19275 (N_19275,N_18684,N_18480);
or U19276 (N_19276,N_18130,N_18559);
nor U19277 (N_19277,N_18398,N_18371);
nand U19278 (N_19278,N_18658,N_18692);
xnor U19279 (N_19279,N_18135,N_18218);
or U19280 (N_19280,N_18323,N_18738);
or U19281 (N_19281,N_18505,N_18647);
nand U19282 (N_19282,N_18200,N_18477);
or U19283 (N_19283,N_18665,N_18340);
nand U19284 (N_19284,N_18506,N_18557);
nor U19285 (N_19285,N_18181,N_18136);
or U19286 (N_19286,N_18731,N_18389);
nand U19287 (N_19287,N_18538,N_18165);
or U19288 (N_19288,N_18664,N_18170);
nor U19289 (N_19289,N_18388,N_18284);
and U19290 (N_19290,N_18518,N_18575);
nand U19291 (N_19291,N_18666,N_18272);
nand U19292 (N_19292,N_18715,N_18334);
nand U19293 (N_19293,N_18564,N_18737);
and U19294 (N_19294,N_18177,N_18297);
or U19295 (N_19295,N_18486,N_18240);
or U19296 (N_19296,N_18568,N_18579);
xnor U19297 (N_19297,N_18732,N_18580);
or U19298 (N_19298,N_18150,N_18696);
or U19299 (N_19299,N_18431,N_18613);
nand U19300 (N_19300,N_18424,N_18684);
nor U19301 (N_19301,N_18582,N_18418);
nor U19302 (N_19302,N_18553,N_18617);
or U19303 (N_19303,N_18326,N_18671);
and U19304 (N_19304,N_18622,N_18177);
or U19305 (N_19305,N_18387,N_18519);
or U19306 (N_19306,N_18437,N_18175);
nor U19307 (N_19307,N_18430,N_18298);
nor U19308 (N_19308,N_18737,N_18281);
nor U19309 (N_19309,N_18616,N_18591);
nor U19310 (N_19310,N_18473,N_18364);
nand U19311 (N_19311,N_18580,N_18636);
xor U19312 (N_19312,N_18398,N_18250);
nor U19313 (N_19313,N_18223,N_18311);
and U19314 (N_19314,N_18228,N_18308);
or U19315 (N_19315,N_18240,N_18675);
and U19316 (N_19316,N_18600,N_18365);
xor U19317 (N_19317,N_18452,N_18340);
or U19318 (N_19318,N_18474,N_18713);
and U19319 (N_19319,N_18191,N_18361);
xor U19320 (N_19320,N_18174,N_18528);
or U19321 (N_19321,N_18486,N_18135);
or U19322 (N_19322,N_18679,N_18284);
nor U19323 (N_19323,N_18399,N_18158);
xnor U19324 (N_19324,N_18458,N_18275);
nand U19325 (N_19325,N_18436,N_18143);
and U19326 (N_19326,N_18458,N_18359);
nor U19327 (N_19327,N_18715,N_18650);
nand U19328 (N_19328,N_18366,N_18198);
nor U19329 (N_19329,N_18397,N_18152);
xor U19330 (N_19330,N_18540,N_18461);
nand U19331 (N_19331,N_18420,N_18275);
or U19332 (N_19332,N_18187,N_18175);
nor U19333 (N_19333,N_18671,N_18306);
or U19334 (N_19334,N_18655,N_18430);
nand U19335 (N_19335,N_18454,N_18594);
and U19336 (N_19336,N_18584,N_18498);
or U19337 (N_19337,N_18486,N_18395);
nor U19338 (N_19338,N_18539,N_18394);
nor U19339 (N_19339,N_18174,N_18126);
and U19340 (N_19340,N_18283,N_18263);
or U19341 (N_19341,N_18333,N_18186);
and U19342 (N_19342,N_18611,N_18163);
nand U19343 (N_19343,N_18622,N_18269);
and U19344 (N_19344,N_18592,N_18554);
nor U19345 (N_19345,N_18662,N_18268);
and U19346 (N_19346,N_18468,N_18197);
and U19347 (N_19347,N_18573,N_18195);
xor U19348 (N_19348,N_18152,N_18325);
and U19349 (N_19349,N_18488,N_18335);
nand U19350 (N_19350,N_18324,N_18510);
or U19351 (N_19351,N_18718,N_18206);
or U19352 (N_19352,N_18637,N_18614);
and U19353 (N_19353,N_18442,N_18526);
nand U19354 (N_19354,N_18368,N_18514);
or U19355 (N_19355,N_18643,N_18585);
nor U19356 (N_19356,N_18613,N_18694);
or U19357 (N_19357,N_18516,N_18432);
or U19358 (N_19358,N_18491,N_18178);
or U19359 (N_19359,N_18689,N_18668);
or U19360 (N_19360,N_18516,N_18380);
and U19361 (N_19361,N_18549,N_18140);
nand U19362 (N_19362,N_18442,N_18228);
nor U19363 (N_19363,N_18342,N_18239);
or U19364 (N_19364,N_18342,N_18195);
xnor U19365 (N_19365,N_18632,N_18653);
or U19366 (N_19366,N_18149,N_18158);
nand U19367 (N_19367,N_18572,N_18604);
and U19368 (N_19368,N_18133,N_18195);
nor U19369 (N_19369,N_18158,N_18686);
or U19370 (N_19370,N_18402,N_18584);
nand U19371 (N_19371,N_18371,N_18309);
or U19372 (N_19372,N_18209,N_18334);
xor U19373 (N_19373,N_18309,N_18379);
nor U19374 (N_19374,N_18391,N_18739);
and U19375 (N_19375,N_18998,N_19081);
nor U19376 (N_19376,N_18834,N_19331);
and U19377 (N_19377,N_19260,N_19097);
nor U19378 (N_19378,N_18795,N_19007);
or U19379 (N_19379,N_19221,N_19075);
nand U19380 (N_19380,N_18776,N_18777);
nor U19381 (N_19381,N_19155,N_19215);
nand U19382 (N_19382,N_19095,N_19112);
nand U19383 (N_19383,N_18893,N_18824);
and U19384 (N_19384,N_18785,N_19094);
xor U19385 (N_19385,N_19175,N_19205);
nor U19386 (N_19386,N_19241,N_19149);
nor U19387 (N_19387,N_19143,N_19090);
and U19388 (N_19388,N_19275,N_18852);
or U19389 (N_19389,N_19104,N_18829);
nand U19390 (N_19390,N_18766,N_18842);
nor U19391 (N_19391,N_19253,N_18894);
nor U19392 (N_19392,N_18938,N_18787);
nand U19393 (N_19393,N_19005,N_18755);
or U19394 (N_19394,N_19234,N_19169);
nand U19395 (N_19395,N_18986,N_19099);
and U19396 (N_19396,N_19259,N_18942);
nand U19397 (N_19397,N_19356,N_19225);
nand U19398 (N_19398,N_19077,N_18912);
xor U19399 (N_19399,N_18906,N_19133);
nand U19400 (N_19400,N_18987,N_19011);
nor U19401 (N_19401,N_19130,N_19083);
or U19402 (N_19402,N_18979,N_19276);
and U19403 (N_19403,N_19268,N_19121);
nor U19404 (N_19404,N_19069,N_18836);
and U19405 (N_19405,N_18769,N_18761);
nand U19406 (N_19406,N_19206,N_19243);
and U19407 (N_19407,N_19118,N_19191);
nor U19408 (N_19408,N_18762,N_18873);
and U19409 (N_19409,N_19132,N_19085);
or U19410 (N_19410,N_19150,N_18818);
and U19411 (N_19411,N_19102,N_18946);
nand U19412 (N_19412,N_19328,N_19245);
and U19413 (N_19413,N_18822,N_19127);
and U19414 (N_19414,N_18870,N_18874);
or U19415 (N_19415,N_19286,N_19349);
or U19416 (N_19416,N_19046,N_19078);
and U19417 (N_19417,N_19096,N_19318);
or U19418 (N_19418,N_19001,N_18884);
or U19419 (N_19419,N_18967,N_19262);
or U19420 (N_19420,N_19354,N_19189);
nand U19421 (N_19421,N_19038,N_18910);
nor U19422 (N_19422,N_18918,N_19016);
nor U19423 (N_19423,N_19371,N_19273);
nand U19424 (N_19424,N_19314,N_19335);
nor U19425 (N_19425,N_18971,N_19255);
and U19426 (N_19426,N_18976,N_19358);
nand U19427 (N_19427,N_19157,N_19125);
nand U19428 (N_19428,N_19263,N_18974);
xnor U19429 (N_19429,N_19184,N_19084);
nand U19430 (N_19430,N_19014,N_19352);
xnor U19431 (N_19431,N_19195,N_18859);
nand U19432 (N_19432,N_19010,N_19071);
and U19433 (N_19433,N_19364,N_19154);
nor U19434 (N_19434,N_19100,N_18897);
nand U19435 (N_19435,N_18904,N_18866);
or U19436 (N_19436,N_18922,N_19338);
and U19437 (N_19437,N_19165,N_18809);
nand U19438 (N_19438,N_19110,N_19250);
nand U19439 (N_19439,N_19146,N_18936);
or U19440 (N_19440,N_19066,N_19108);
nor U19441 (N_19441,N_19185,N_18995);
nand U19442 (N_19442,N_18871,N_18768);
or U19443 (N_19443,N_19319,N_19126);
or U19444 (N_19444,N_18810,N_19171);
or U19445 (N_19445,N_19285,N_19012);
and U19446 (N_19446,N_19366,N_19117);
and U19447 (N_19447,N_19296,N_19135);
nor U19448 (N_19448,N_19030,N_18862);
and U19449 (N_19449,N_19087,N_19124);
nand U19450 (N_19450,N_19043,N_18925);
and U19451 (N_19451,N_18789,N_18933);
xnor U19452 (N_19452,N_18781,N_19049);
nor U19453 (N_19453,N_18772,N_19266);
xnor U19454 (N_19454,N_19086,N_18931);
nand U19455 (N_19455,N_19278,N_18783);
and U19456 (N_19456,N_19092,N_18790);
nor U19457 (N_19457,N_18993,N_19337);
and U19458 (N_19458,N_19256,N_18883);
xnor U19459 (N_19459,N_19339,N_19018);
and U19460 (N_19460,N_19080,N_18991);
nand U19461 (N_19461,N_19107,N_18813);
and U19462 (N_19462,N_18929,N_19194);
nand U19463 (N_19463,N_18774,N_19362);
and U19464 (N_19464,N_18955,N_18989);
or U19465 (N_19465,N_19247,N_19122);
nor U19466 (N_19466,N_18863,N_19373);
or U19467 (N_19467,N_19309,N_18764);
or U19468 (N_19468,N_19166,N_19021);
or U19469 (N_19469,N_19330,N_18850);
nor U19470 (N_19470,N_18988,N_18860);
nor U19471 (N_19471,N_19345,N_19312);
nor U19472 (N_19472,N_19004,N_19332);
nor U19473 (N_19473,N_18994,N_19105);
xnor U19474 (N_19474,N_18821,N_19131);
xnor U19475 (N_19475,N_18954,N_19246);
xnor U19476 (N_19476,N_18964,N_19272);
nor U19477 (N_19477,N_19148,N_19176);
and U19478 (N_19478,N_19288,N_19074);
or U19479 (N_19479,N_19281,N_19251);
or U19480 (N_19480,N_19200,N_18844);
or U19481 (N_19481,N_18792,N_19106);
or U19482 (N_19482,N_19289,N_19283);
nor U19483 (N_19483,N_19180,N_19182);
nand U19484 (N_19484,N_19291,N_18791);
or U19485 (N_19485,N_19152,N_19211);
and U19486 (N_19486,N_19213,N_19050);
xnor U19487 (N_19487,N_19311,N_19320);
nand U19488 (N_19488,N_18750,N_19279);
or U19489 (N_19489,N_18948,N_18984);
nor U19490 (N_19490,N_19231,N_18779);
xnor U19491 (N_19491,N_18797,N_19091);
nand U19492 (N_19492,N_19115,N_19254);
nand U19493 (N_19493,N_18962,N_18924);
or U19494 (N_19494,N_18832,N_19045);
and U19495 (N_19495,N_19026,N_18830);
and U19496 (N_19496,N_18796,N_18794);
or U19497 (N_19497,N_18996,N_18939);
nor U19498 (N_19498,N_19162,N_19218);
xnor U19499 (N_19499,N_19070,N_19370);
nor U19500 (N_19500,N_18869,N_18753);
or U19501 (N_19501,N_19039,N_18812);
or U19502 (N_19502,N_19028,N_19302);
and U19503 (N_19503,N_19212,N_19308);
or U19504 (N_19504,N_19041,N_19202);
nand U19505 (N_19505,N_19188,N_18786);
nor U19506 (N_19506,N_18978,N_18926);
and U19507 (N_19507,N_19196,N_19156);
xnor U19508 (N_19508,N_18877,N_19027);
xnor U19509 (N_19509,N_18800,N_19067);
or U19510 (N_19510,N_19164,N_18833);
nand U19511 (N_19511,N_18826,N_18950);
and U19512 (N_19512,N_19114,N_18920);
nand U19513 (N_19513,N_18778,N_19013);
nor U19514 (N_19514,N_18997,N_19161);
and U19515 (N_19515,N_19216,N_19181);
and U19516 (N_19516,N_18945,N_19151);
and U19517 (N_19517,N_19361,N_18837);
xnor U19518 (N_19518,N_19183,N_18804);
and U19519 (N_19519,N_19301,N_18798);
nor U19520 (N_19520,N_18793,N_19210);
nand U19521 (N_19521,N_18811,N_18802);
and U19522 (N_19522,N_19227,N_18903);
nand U19523 (N_19523,N_19329,N_19034);
nand U19524 (N_19524,N_19129,N_18843);
and U19525 (N_19525,N_19187,N_19303);
xnor U19526 (N_19526,N_19153,N_19101);
or U19527 (N_19527,N_19022,N_18828);
nor U19528 (N_19528,N_18803,N_19002);
or U19529 (N_19529,N_18838,N_19137);
or U19530 (N_19530,N_18973,N_19248);
and U19531 (N_19531,N_18853,N_18835);
nor U19532 (N_19532,N_19008,N_18890);
and U19533 (N_19533,N_18953,N_18868);
and U19534 (N_19534,N_19052,N_18981);
and U19535 (N_19535,N_18817,N_19280);
nor U19536 (N_19536,N_18908,N_19235);
nand U19537 (N_19537,N_19024,N_19267);
or U19538 (N_19538,N_19238,N_19119);
nand U19539 (N_19539,N_18815,N_19025);
and U19540 (N_19540,N_19140,N_18891);
or U19541 (N_19541,N_18754,N_19158);
nor U19542 (N_19542,N_18928,N_18845);
and U19543 (N_19543,N_19261,N_18858);
and U19544 (N_19544,N_19103,N_19214);
or U19545 (N_19545,N_18881,N_18864);
and U19546 (N_19546,N_18980,N_19047);
or U19547 (N_19547,N_19229,N_19368);
nor U19548 (N_19548,N_18956,N_19357);
or U19549 (N_19549,N_18900,N_19219);
and U19550 (N_19550,N_19073,N_18855);
nand U19551 (N_19551,N_18851,N_19292);
nand U19552 (N_19552,N_19051,N_19033);
or U19553 (N_19553,N_18839,N_19340);
xor U19554 (N_19554,N_18968,N_19306);
or U19555 (N_19555,N_19350,N_18782);
or U19556 (N_19556,N_19333,N_19174);
or U19557 (N_19557,N_19347,N_19003);
or U19558 (N_19558,N_19230,N_18872);
or U19559 (N_19559,N_19224,N_18935);
nand U19560 (N_19560,N_18915,N_19145);
nand U19561 (N_19561,N_19056,N_19116);
nand U19562 (N_19562,N_18889,N_19284);
nand U19563 (N_19563,N_18885,N_19277);
xor U19564 (N_19564,N_19029,N_19113);
nor U19565 (N_19565,N_19139,N_19023);
or U19566 (N_19566,N_18765,N_18959);
nor U19567 (N_19567,N_19365,N_19326);
or U19568 (N_19568,N_19061,N_18882);
and U19569 (N_19569,N_18759,N_18937);
nor U19570 (N_19570,N_19141,N_18895);
or U19571 (N_19571,N_19346,N_19360);
and U19572 (N_19572,N_19000,N_18767);
nand U19573 (N_19573,N_19089,N_19197);
and U19574 (N_19574,N_19232,N_19369);
and U19575 (N_19575,N_18840,N_19072);
nor U19576 (N_19576,N_19134,N_19053);
nand U19577 (N_19577,N_19159,N_18770);
and U19578 (N_19578,N_19217,N_19237);
xor U19579 (N_19579,N_19316,N_18823);
nor U19580 (N_19580,N_19098,N_18963);
nand U19581 (N_19581,N_18827,N_18999);
and U19582 (N_19582,N_19015,N_18788);
xor U19583 (N_19583,N_18819,N_18775);
nand U19584 (N_19584,N_19058,N_19136);
nand U19585 (N_19585,N_19290,N_18972);
or U19586 (N_19586,N_19293,N_19363);
nand U19587 (N_19587,N_18977,N_19040);
xor U19588 (N_19588,N_18848,N_19274);
nand U19589 (N_19589,N_19048,N_18909);
xnor U19590 (N_19590,N_18752,N_19258);
or U19591 (N_19591,N_18807,N_18970);
xor U19592 (N_19592,N_19325,N_19063);
and U19593 (N_19593,N_18856,N_19179);
or U19594 (N_19594,N_18896,N_19064);
or U19595 (N_19595,N_19128,N_18846);
or U19596 (N_19596,N_18758,N_19336);
and U19597 (N_19597,N_18921,N_19372);
and U19598 (N_19598,N_18888,N_18751);
nand U19599 (N_19599,N_19059,N_19321);
nand U19600 (N_19600,N_19178,N_18905);
or U19601 (N_19601,N_19020,N_18983);
nor U19602 (N_19602,N_18876,N_19298);
nor U19603 (N_19603,N_18899,N_18911);
or U19604 (N_19604,N_19239,N_19359);
or U19605 (N_19605,N_18949,N_19093);
or U19606 (N_19606,N_19282,N_19057);
or U19607 (N_19607,N_19341,N_19264);
nand U19608 (N_19608,N_18990,N_19172);
nand U19609 (N_19609,N_18941,N_18784);
nand U19610 (N_19610,N_18757,N_18806);
or U19611 (N_19611,N_19186,N_19270);
nor U19612 (N_19612,N_19160,N_19170);
nor U19613 (N_19613,N_18878,N_19177);
or U19614 (N_19614,N_18875,N_19367);
or U19615 (N_19615,N_19348,N_19168);
xnor U19616 (N_19616,N_18867,N_18902);
nand U19617 (N_19617,N_18982,N_18886);
and U19618 (N_19618,N_19236,N_19042);
nand U19619 (N_19619,N_19323,N_19017);
and U19620 (N_19620,N_19287,N_19032);
nor U19621 (N_19621,N_18943,N_19198);
xor U19622 (N_19622,N_18940,N_19310);
nand U19623 (N_19623,N_19223,N_19068);
or U19624 (N_19624,N_19120,N_18857);
and U19625 (N_19625,N_18831,N_19173);
and U19626 (N_19626,N_19204,N_19220);
or U19627 (N_19627,N_19265,N_19203);
and U19628 (N_19628,N_19044,N_19355);
xnor U19629 (N_19629,N_18930,N_19344);
or U19630 (N_19630,N_19313,N_18816);
nor U19631 (N_19631,N_19079,N_18898);
and U19632 (N_19632,N_18808,N_19208);
nor U19633 (N_19633,N_19295,N_19167);
nor U19634 (N_19634,N_18907,N_18879);
or U19635 (N_19635,N_19299,N_19222);
and U19636 (N_19636,N_19233,N_18934);
or U19637 (N_19637,N_18887,N_19271);
and U19638 (N_19638,N_18847,N_18975);
xor U19639 (N_19639,N_19252,N_18914);
or U19640 (N_19640,N_18966,N_19109);
and U19641 (N_19641,N_19226,N_19304);
nor U19642 (N_19642,N_19088,N_19019);
or U19643 (N_19643,N_19315,N_19353);
and U19644 (N_19644,N_19322,N_19163);
or U19645 (N_19645,N_19111,N_19244);
xnor U19646 (N_19646,N_19242,N_18913);
and U19647 (N_19647,N_19006,N_18960);
nand U19648 (N_19648,N_19082,N_18969);
or U19649 (N_19649,N_19138,N_19144);
nand U19650 (N_19650,N_18763,N_19060);
nor U19651 (N_19651,N_19305,N_18923);
nor U19652 (N_19652,N_19343,N_19351);
nand U19653 (N_19653,N_18799,N_19009);
or U19654 (N_19654,N_18917,N_18892);
xor U19655 (N_19655,N_18805,N_18771);
or U19656 (N_19656,N_19147,N_19055);
nor U19657 (N_19657,N_18952,N_18947);
nand U19658 (N_19658,N_19076,N_18957);
or U19659 (N_19659,N_18801,N_19374);
or U19660 (N_19660,N_18849,N_18944);
nand U19661 (N_19661,N_19327,N_18919);
nand U19662 (N_19662,N_19190,N_18814);
nand U19663 (N_19663,N_19062,N_18916);
nand U19664 (N_19664,N_19324,N_19240);
and U19665 (N_19665,N_18841,N_18958);
or U19666 (N_19666,N_19031,N_18985);
nor U19667 (N_19667,N_18901,N_19257);
nor U19668 (N_19668,N_18865,N_18961);
nor U19669 (N_19669,N_19228,N_18880);
or U19670 (N_19670,N_18927,N_19142);
xnor U19671 (N_19671,N_19201,N_19300);
and U19672 (N_19672,N_18780,N_19035);
or U19673 (N_19673,N_19193,N_19294);
nand U19674 (N_19674,N_19269,N_18932);
or U19675 (N_19675,N_19207,N_18951);
nor U19676 (N_19676,N_18861,N_18820);
and U19677 (N_19677,N_18756,N_19192);
and U19678 (N_19678,N_18992,N_19065);
nor U19679 (N_19679,N_19036,N_18760);
and U19680 (N_19680,N_19307,N_18773);
or U19681 (N_19681,N_19249,N_19199);
nand U19682 (N_19682,N_18965,N_18854);
or U19683 (N_19683,N_19342,N_19209);
or U19684 (N_19684,N_19334,N_19297);
or U19685 (N_19685,N_19123,N_19054);
or U19686 (N_19686,N_19317,N_19037);
nand U19687 (N_19687,N_18825,N_18924);
and U19688 (N_19688,N_19326,N_19023);
nor U19689 (N_19689,N_18889,N_18918);
and U19690 (N_19690,N_19194,N_19162);
nor U19691 (N_19691,N_18919,N_19056);
xor U19692 (N_19692,N_19235,N_19369);
and U19693 (N_19693,N_18808,N_18797);
xnor U19694 (N_19694,N_19187,N_19090);
or U19695 (N_19695,N_18761,N_19180);
xor U19696 (N_19696,N_18834,N_19123);
or U19697 (N_19697,N_19138,N_19082);
nor U19698 (N_19698,N_19050,N_19206);
nand U19699 (N_19699,N_18859,N_19144);
nor U19700 (N_19700,N_18789,N_18843);
nand U19701 (N_19701,N_18799,N_19240);
nor U19702 (N_19702,N_19213,N_18941);
nor U19703 (N_19703,N_18953,N_18756);
or U19704 (N_19704,N_19157,N_18812);
xnor U19705 (N_19705,N_19359,N_19189);
nand U19706 (N_19706,N_19227,N_18923);
or U19707 (N_19707,N_18754,N_18809);
nand U19708 (N_19708,N_19001,N_19203);
xnor U19709 (N_19709,N_18750,N_18985);
or U19710 (N_19710,N_19078,N_19033);
nand U19711 (N_19711,N_18949,N_18846);
nor U19712 (N_19712,N_18903,N_18796);
and U19713 (N_19713,N_19269,N_19343);
nor U19714 (N_19714,N_19010,N_19065);
and U19715 (N_19715,N_19354,N_19251);
and U19716 (N_19716,N_19364,N_19082);
or U19717 (N_19717,N_19119,N_18987);
nor U19718 (N_19718,N_19002,N_19094);
nand U19719 (N_19719,N_19267,N_18908);
or U19720 (N_19720,N_18956,N_19016);
and U19721 (N_19721,N_19205,N_18755);
nand U19722 (N_19722,N_19200,N_19136);
or U19723 (N_19723,N_18866,N_18762);
and U19724 (N_19724,N_19181,N_18992);
nor U19725 (N_19725,N_19326,N_19035);
nor U19726 (N_19726,N_19121,N_19064);
nor U19727 (N_19727,N_19319,N_18766);
or U19728 (N_19728,N_18855,N_18838);
nand U19729 (N_19729,N_18869,N_18852);
xor U19730 (N_19730,N_19245,N_18984);
nand U19731 (N_19731,N_19096,N_18857);
and U19732 (N_19732,N_18966,N_18870);
or U19733 (N_19733,N_19143,N_19272);
or U19734 (N_19734,N_18979,N_19292);
or U19735 (N_19735,N_18983,N_18831);
nand U19736 (N_19736,N_19041,N_18789);
nand U19737 (N_19737,N_19168,N_19217);
nand U19738 (N_19738,N_19121,N_18826);
nand U19739 (N_19739,N_19211,N_19246);
and U19740 (N_19740,N_18923,N_18989);
or U19741 (N_19741,N_19226,N_18838);
nor U19742 (N_19742,N_19186,N_19156);
and U19743 (N_19743,N_18977,N_19270);
and U19744 (N_19744,N_18917,N_19161);
or U19745 (N_19745,N_18778,N_19077);
or U19746 (N_19746,N_18871,N_18913);
nand U19747 (N_19747,N_18877,N_18939);
or U19748 (N_19748,N_18934,N_18809);
and U19749 (N_19749,N_19188,N_18851);
xnor U19750 (N_19750,N_19087,N_18828);
nand U19751 (N_19751,N_19096,N_18828);
or U19752 (N_19752,N_19368,N_19028);
nor U19753 (N_19753,N_19122,N_19082);
xor U19754 (N_19754,N_18770,N_19353);
nor U19755 (N_19755,N_19235,N_19161);
nor U19756 (N_19756,N_18956,N_18855);
nor U19757 (N_19757,N_18826,N_18925);
nand U19758 (N_19758,N_19087,N_18756);
and U19759 (N_19759,N_18753,N_19091);
nand U19760 (N_19760,N_19189,N_19107);
or U19761 (N_19761,N_18887,N_18989);
nor U19762 (N_19762,N_18928,N_18889);
and U19763 (N_19763,N_18808,N_19362);
or U19764 (N_19764,N_18918,N_18753);
nor U19765 (N_19765,N_19216,N_19349);
nor U19766 (N_19766,N_19074,N_18931);
nand U19767 (N_19767,N_19252,N_19365);
xnor U19768 (N_19768,N_19001,N_18974);
xnor U19769 (N_19769,N_18753,N_18939);
nor U19770 (N_19770,N_19314,N_19172);
and U19771 (N_19771,N_18757,N_19242);
or U19772 (N_19772,N_19238,N_19215);
and U19773 (N_19773,N_18992,N_18928);
nor U19774 (N_19774,N_19224,N_19316);
and U19775 (N_19775,N_19053,N_19104);
and U19776 (N_19776,N_18874,N_19291);
or U19777 (N_19777,N_19170,N_18926);
nand U19778 (N_19778,N_19211,N_18897);
or U19779 (N_19779,N_19077,N_19192);
and U19780 (N_19780,N_19129,N_19283);
nand U19781 (N_19781,N_19235,N_18753);
or U19782 (N_19782,N_18835,N_18810);
and U19783 (N_19783,N_18889,N_19174);
and U19784 (N_19784,N_18882,N_18907);
and U19785 (N_19785,N_18879,N_18901);
nand U19786 (N_19786,N_19175,N_18800);
xor U19787 (N_19787,N_19260,N_18900);
or U19788 (N_19788,N_18951,N_19051);
nand U19789 (N_19789,N_19296,N_19298);
nand U19790 (N_19790,N_18993,N_18973);
or U19791 (N_19791,N_18853,N_18750);
xnor U19792 (N_19792,N_19155,N_18906);
nand U19793 (N_19793,N_18937,N_18917);
or U19794 (N_19794,N_19273,N_18901);
and U19795 (N_19795,N_18986,N_18796);
nand U19796 (N_19796,N_19298,N_19278);
or U19797 (N_19797,N_19298,N_19367);
xor U19798 (N_19798,N_19219,N_19191);
and U19799 (N_19799,N_19000,N_19312);
nand U19800 (N_19800,N_18814,N_19218);
and U19801 (N_19801,N_18913,N_19082);
nand U19802 (N_19802,N_19374,N_19062);
nor U19803 (N_19803,N_18796,N_19190);
xor U19804 (N_19804,N_18800,N_19358);
nor U19805 (N_19805,N_19172,N_18936);
or U19806 (N_19806,N_19148,N_18895);
nand U19807 (N_19807,N_18836,N_19131);
nand U19808 (N_19808,N_18926,N_19297);
nand U19809 (N_19809,N_19185,N_19310);
and U19810 (N_19810,N_18907,N_18812);
nand U19811 (N_19811,N_19011,N_18938);
or U19812 (N_19812,N_18978,N_19067);
or U19813 (N_19813,N_19252,N_19230);
and U19814 (N_19814,N_18775,N_19045);
or U19815 (N_19815,N_19346,N_19309);
nand U19816 (N_19816,N_19059,N_18835);
nor U19817 (N_19817,N_19290,N_18768);
nor U19818 (N_19818,N_18896,N_19308);
xnor U19819 (N_19819,N_19272,N_18970);
or U19820 (N_19820,N_18888,N_19198);
nand U19821 (N_19821,N_19157,N_18876);
nor U19822 (N_19822,N_18967,N_19340);
and U19823 (N_19823,N_18957,N_19178);
nor U19824 (N_19824,N_19227,N_19060);
nor U19825 (N_19825,N_19062,N_18811);
or U19826 (N_19826,N_19041,N_18852);
nor U19827 (N_19827,N_19164,N_18835);
xor U19828 (N_19828,N_19336,N_19012);
and U19829 (N_19829,N_18840,N_18953);
or U19830 (N_19830,N_18792,N_19247);
or U19831 (N_19831,N_19291,N_19106);
nand U19832 (N_19832,N_18770,N_19229);
and U19833 (N_19833,N_18897,N_19360);
nand U19834 (N_19834,N_19105,N_18922);
and U19835 (N_19835,N_18824,N_19256);
nor U19836 (N_19836,N_18935,N_18759);
nor U19837 (N_19837,N_19019,N_18851);
nor U19838 (N_19838,N_18900,N_19217);
and U19839 (N_19839,N_19305,N_19159);
and U19840 (N_19840,N_18923,N_19276);
nand U19841 (N_19841,N_18910,N_19272);
nor U19842 (N_19842,N_19141,N_19293);
nand U19843 (N_19843,N_19140,N_19092);
and U19844 (N_19844,N_19248,N_19358);
nand U19845 (N_19845,N_19191,N_18946);
xor U19846 (N_19846,N_18967,N_19298);
and U19847 (N_19847,N_19091,N_19360);
or U19848 (N_19848,N_19090,N_19342);
nor U19849 (N_19849,N_19111,N_18790);
nand U19850 (N_19850,N_19360,N_19046);
or U19851 (N_19851,N_18909,N_18868);
nand U19852 (N_19852,N_19254,N_18917);
nand U19853 (N_19853,N_18769,N_18946);
nor U19854 (N_19854,N_18940,N_18974);
or U19855 (N_19855,N_19053,N_19185);
nand U19856 (N_19856,N_19256,N_18959);
or U19857 (N_19857,N_18903,N_18939);
xor U19858 (N_19858,N_19090,N_19175);
nor U19859 (N_19859,N_18856,N_18839);
or U19860 (N_19860,N_18876,N_19064);
nor U19861 (N_19861,N_19186,N_19166);
or U19862 (N_19862,N_19355,N_19108);
or U19863 (N_19863,N_18815,N_18840);
nand U19864 (N_19864,N_18948,N_18993);
or U19865 (N_19865,N_19304,N_18824);
nor U19866 (N_19866,N_18944,N_19217);
nand U19867 (N_19867,N_19105,N_18815);
nor U19868 (N_19868,N_19266,N_19268);
xor U19869 (N_19869,N_19267,N_18854);
and U19870 (N_19870,N_19246,N_18836);
nand U19871 (N_19871,N_19353,N_18805);
nor U19872 (N_19872,N_18929,N_19314);
nand U19873 (N_19873,N_19264,N_18781);
xnor U19874 (N_19874,N_19037,N_19314);
nand U19875 (N_19875,N_19054,N_19200);
xnor U19876 (N_19876,N_18844,N_19251);
and U19877 (N_19877,N_18956,N_18770);
nor U19878 (N_19878,N_18823,N_18979);
nor U19879 (N_19879,N_19105,N_18915);
and U19880 (N_19880,N_18837,N_19200);
xor U19881 (N_19881,N_19205,N_19299);
nor U19882 (N_19882,N_18764,N_19264);
nor U19883 (N_19883,N_18968,N_18909);
nor U19884 (N_19884,N_19366,N_19213);
and U19885 (N_19885,N_18813,N_19298);
nand U19886 (N_19886,N_19299,N_18769);
nor U19887 (N_19887,N_18901,N_18888);
nor U19888 (N_19888,N_19372,N_19079);
nand U19889 (N_19889,N_18932,N_18761);
and U19890 (N_19890,N_19132,N_19073);
or U19891 (N_19891,N_19337,N_18902);
xor U19892 (N_19892,N_19141,N_19192);
and U19893 (N_19893,N_19151,N_19291);
xor U19894 (N_19894,N_19270,N_19355);
or U19895 (N_19895,N_18878,N_19241);
or U19896 (N_19896,N_18906,N_19100);
nand U19897 (N_19897,N_19323,N_18978);
nand U19898 (N_19898,N_19183,N_19127);
or U19899 (N_19899,N_18868,N_18758);
xor U19900 (N_19900,N_18786,N_19038);
and U19901 (N_19901,N_19180,N_19218);
and U19902 (N_19902,N_18989,N_18804);
nand U19903 (N_19903,N_19066,N_19208);
and U19904 (N_19904,N_19163,N_19181);
and U19905 (N_19905,N_18777,N_18967);
xnor U19906 (N_19906,N_18943,N_19143);
or U19907 (N_19907,N_18956,N_19227);
or U19908 (N_19908,N_19004,N_18932);
nor U19909 (N_19909,N_19041,N_19225);
and U19910 (N_19910,N_18962,N_19325);
xnor U19911 (N_19911,N_19085,N_19198);
and U19912 (N_19912,N_19011,N_19116);
and U19913 (N_19913,N_19220,N_18908);
and U19914 (N_19914,N_19004,N_18776);
and U19915 (N_19915,N_19114,N_18825);
nand U19916 (N_19916,N_19114,N_19349);
and U19917 (N_19917,N_19231,N_19110);
nor U19918 (N_19918,N_18982,N_19091);
and U19919 (N_19919,N_19277,N_18814);
or U19920 (N_19920,N_19249,N_19075);
nand U19921 (N_19921,N_19062,N_19126);
or U19922 (N_19922,N_18842,N_18871);
and U19923 (N_19923,N_19039,N_19316);
and U19924 (N_19924,N_19337,N_18895);
nor U19925 (N_19925,N_19120,N_19372);
xnor U19926 (N_19926,N_18799,N_19180);
and U19927 (N_19927,N_18833,N_18755);
or U19928 (N_19928,N_19142,N_18825);
and U19929 (N_19929,N_19170,N_19061);
nor U19930 (N_19930,N_18811,N_18919);
and U19931 (N_19931,N_18820,N_18961);
nand U19932 (N_19932,N_19180,N_18955);
or U19933 (N_19933,N_19153,N_18963);
nand U19934 (N_19934,N_18841,N_19025);
or U19935 (N_19935,N_18981,N_19194);
and U19936 (N_19936,N_19250,N_18801);
nor U19937 (N_19937,N_19368,N_18757);
nand U19938 (N_19938,N_19060,N_18916);
nand U19939 (N_19939,N_19340,N_19117);
nor U19940 (N_19940,N_18944,N_19362);
nor U19941 (N_19941,N_18842,N_19361);
nand U19942 (N_19942,N_18761,N_18850);
or U19943 (N_19943,N_19318,N_18887);
and U19944 (N_19944,N_18801,N_18788);
nor U19945 (N_19945,N_19223,N_18962);
xor U19946 (N_19946,N_18895,N_19077);
xnor U19947 (N_19947,N_19195,N_18931);
nand U19948 (N_19948,N_18954,N_18798);
or U19949 (N_19949,N_18910,N_19140);
and U19950 (N_19950,N_19309,N_19162);
or U19951 (N_19951,N_19238,N_19076);
and U19952 (N_19952,N_19304,N_19066);
and U19953 (N_19953,N_18844,N_19290);
nand U19954 (N_19954,N_19187,N_18897);
nand U19955 (N_19955,N_19224,N_19270);
or U19956 (N_19956,N_18928,N_19193);
or U19957 (N_19957,N_18833,N_19340);
xor U19958 (N_19958,N_19166,N_19153);
xor U19959 (N_19959,N_19371,N_19094);
xnor U19960 (N_19960,N_19280,N_18853);
or U19961 (N_19961,N_19085,N_18758);
nand U19962 (N_19962,N_19084,N_18767);
nand U19963 (N_19963,N_19278,N_18766);
xor U19964 (N_19964,N_19018,N_19169);
or U19965 (N_19965,N_19325,N_18774);
and U19966 (N_19966,N_19006,N_19157);
and U19967 (N_19967,N_18877,N_19250);
nor U19968 (N_19968,N_19037,N_18973);
and U19969 (N_19969,N_19257,N_18956);
nor U19970 (N_19970,N_18828,N_19339);
and U19971 (N_19971,N_19100,N_18887);
nand U19972 (N_19972,N_19150,N_19245);
nor U19973 (N_19973,N_19006,N_18842);
and U19974 (N_19974,N_19299,N_19296);
or U19975 (N_19975,N_19195,N_19270);
and U19976 (N_19976,N_19035,N_19188);
and U19977 (N_19977,N_18837,N_19048);
and U19978 (N_19978,N_18806,N_18829);
nor U19979 (N_19979,N_19266,N_19003);
nor U19980 (N_19980,N_19146,N_19278);
nand U19981 (N_19981,N_18823,N_19278);
or U19982 (N_19982,N_19152,N_19207);
or U19983 (N_19983,N_18802,N_19310);
nand U19984 (N_19984,N_18876,N_18757);
or U19985 (N_19985,N_19362,N_19311);
or U19986 (N_19986,N_19333,N_19030);
nor U19987 (N_19987,N_19347,N_19116);
nand U19988 (N_19988,N_18938,N_19200);
and U19989 (N_19989,N_19234,N_18793);
xnor U19990 (N_19990,N_19112,N_18772);
or U19991 (N_19991,N_18816,N_18857);
and U19992 (N_19992,N_18835,N_18874);
nor U19993 (N_19993,N_18782,N_19151);
or U19994 (N_19994,N_19360,N_18893);
nor U19995 (N_19995,N_18845,N_19120);
nor U19996 (N_19996,N_18867,N_18903);
or U19997 (N_19997,N_18766,N_18849);
and U19998 (N_19998,N_19328,N_19209);
nand U19999 (N_19999,N_19364,N_18807);
nor U20000 (N_20000,N_19456,N_19882);
nand U20001 (N_20001,N_19715,N_19435);
and U20002 (N_20002,N_19974,N_19551);
xor U20003 (N_20003,N_19858,N_19642);
nand U20004 (N_20004,N_19603,N_19469);
and U20005 (N_20005,N_19506,N_19756);
nor U20006 (N_20006,N_19912,N_19870);
nor U20007 (N_20007,N_19583,N_19765);
and U20008 (N_20008,N_19448,N_19830);
and U20009 (N_20009,N_19693,N_19592);
nand U20010 (N_20010,N_19658,N_19661);
nor U20011 (N_20011,N_19421,N_19723);
nor U20012 (N_20012,N_19970,N_19464);
and U20013 (N_20013,N_19695,N_19995);
nand U20014 (N_20014,N_19639,N_19800);
nand U20015 (N_20015,N_19669,N_19763);
nand U20016 (N_20016,N_19581,N_19517);
nand U20017 (N_20017,N_19805,N_19400);
nor U20018 (N_20018,N_19475,N_19522);
nand U20019 (N_20019,N_19527,N_19379);
nor U20020 (N_20020,N_19722,N_19673);
nand U20021 (N_20021,N_19503,N_19633);
nand U20022 (N_20022,N_19746,N_19494);
and U20023 (N_20023,N_19961,N_19815);
nand U20024 (N_20024,N_19457,N_19502);
nor U20025 (N_20025,N_19786,N_19836);
or U20026 (N_20026,N_19659,N_19876);
xnor U20027 (N_20027,N_19567,N_19549);
xor U20028 (N_20028,N_19634,N_19415);
nand U20029 (N_20029,N_19611,N_19663);
xor U20030 (N_20030,N_19542,N_19727);
or U20031 (N_20031,N_19788,N_19606);
and U20032 (N_20032,N_19760,N_19461);
xor U20033 (N_20033,N_19779,N_19810);
nor U20034 (N_20034,N_19431,N_19411);
and U20035 (N_20035,N_19885,N_19942);
or U20036 (N_20036,N_19685,N_19433);
or U20037 (N_20037,N_19651,N_19519);
xnor U20038 (N_20038,N_19773,N_19510);
or U20039 (N_20039,N_19934,N_19463);
nand U20040 (N_20040,N_19489,N_19476);
or U20041 (N_20041,N_19544,N_19785);
and U20042 (N_20042,N_19408,N_19670);
or U20043 (N_20043,N_19931,N_19967);
xor U20044 (N_20044,N_19832,N_19748);
or U20045 (N_20045,N_19846,N_19985);
xor U20046 (N_20046,N_19598,N_19822);
or U20047 (N_20047,N_19500,N_19621);
nand U20048 (N_20048,N_19617,N_19817);
nand U20049 (N_20049,N_19524,N_19656);
and U20050 (N_20050,N_19413,N_19787);
and U20051 (N_20051,N_19619,N_19930);
nor U20052 (N_20052,N_19466,N_19625);
and U20053 (N_20053,N_19873,N_19863);
and U20054 (N_20054,N_19736,N_19532);
xor U20055 (N_20055,N_19755,N_19399);
nand U20056 (N_20056,N_19790,N_19718);
or U20057 (N_20057,N_19759,N_19481);
nand U20058 (N_20058,N_19681,N_19537);
and U20059 (N_20059,N_19847,N_19975);
nand U20060 (N_20060,N_19450,N_19907);
and U20061 (N_20061,N_19555,N_19531);
or U20062 (N_20062,N_19593,N_19825);
nand U20063 (N_20063,N_19996,N_19483);
and U20064 (N_20064,N_19979,N_19962);
nand U20065 (N_20065,N_19726,N_19526);
xor U20066 (N_20066,N_19960,N_19808);
nor U20067 (N_20067,N_19686,N_19493);
or U20068 (N_20068,N_19430,N_19410);
nor U20069 (N_20069,N_19601,N_19791);
and U20070 (N_20070,N_19477,N_19612);
and U20071 (N_20071,N_19406,N_19711);
nand U20072 (N_20072,N_19929,N_19577);
or U20073 (N_20073,N_19576,N_19745);
nor U20074 (N_20074,N_19794,N_19487);
or U20075 (N_20075,N_19385,N_19933);
and U20076 (N_20076,N_19789,N_19798);
xnor U20077 (N_20077,N_19793,N_19602);
and U20078 (N_20078,N_19843,N_19699);
and U20079 (N_20079,N_19921,N_19888);
xor U20080 (N_20080,N_19386,N_19398);
nand U20081 (N_20081,N_19820,N_19646);
or U20082 (N_20082,N_19886,N_19495);
and U20083 (N_20083,N_19919,N_19570);
or U20084 (N_20084,N_19608,N_19378);
and U20085 (N_20085,N_19467,N_19590);
and U20086 (N_20086,N_19772,N_19432);
nor U20087 (N_20087,N_19445,N_19958);
nor U20088 (N_20088,N_19905,N_19729);
nand U20089 (N_20089,N_19868,N_19556);
or U20090 (N_20090,N_19733,N_19648);
xnor U20091 (N_20091,N_19849,N_19917);
or U20092 (N_20092,N_19471,N_19497);
nor U20093 (N_20093,N_19762,N_19998);
and U20094 (N_20094,N_19380,N_19376);
or U20095 (N_20095,N_19394,N_19383);
nand U20096 (N_20096,N_19875,N_19405);
nor U20097 (N_20097,N_19898,N_19547);
or U20098 (N_20098,N_19558,N_19935);
and U20099 (N_20099,N_19375,N_19538);
nand U20100 (N_20100,N_19384,N_19496);
and U20101 (N_20101,N_19856,N_19554);
or U20102 (N_20102,N_19480,N_19833);
and U20103 (N_20103,N_19874,N_19705);
nand U20104 (N_20104,N_19428,N_19626);
and U20105 (N_20105,N_19412,N_19507);
nand U20106 (N_20106,N_19541,N_19903);
xor U20107 (N_20107,N_19697,N_19778);
xnor U20108 (N_20108,N_19943,N_19687);
nand U20109 (N_20109,N_19986,N_19439);
xor U20110 (N_20110,N_19529,N_19473);
and U20111 (N_20111,N_19490,N_19860);
nand U20112 (N_20112,N_19546,N_19908);
and U20113 (N_20113,N_19855,N_19725);
nand U20114 (N_20114,N_19696,N_19923);
nor U20115 (N_20115,N_19769,N_19613);
nand U20116 (N_20116,N_19951,N_19774);
nor U20117 (N_20117,N_19831,N_19389);
nand U20118 (N_20118,N_19871,N_19864);
or U20119 (N_20119,N_19777,N_19989);
or U20120 (N_20120,N_19595,N_19417);
and U20121 (N_20121,N_19395,N_19586);
nor U20122 (N_20122,N_19802,N_19622);
and U20123 (N_20123,N_19580,N_19574);
or U20124 (N_20124,N_19717,N_19465);
and U20125 (N_20125,N_19927,N_19382);
nand U20126 (N_20126,N_19916,N_19978);
nand U20127 (N_20127,N_19972,N_19650);
and U20128 (N_20128,N_19819,N_19910);
or U20129 (N_20129,N_19734,N_19568);
nor U20130 (N_20130,N_19700,N_19573);
or U20131 (N_20131,N_19713,N_19928);
nand U20132 (N_20132,N_19926,N_19749);
and U20133 (N_20133,N_19614,N_19911);
and U20134 (N_20134,N_19638,N_19835);
and U20135 (N_20135,N_19904,N_19859);
nand U20136 (N_20136,N_19971,N_19414);
nor U20137 (N_20137,N_19716,N_19680);
or U20138 (N_20138,N_19643,N_19829);
nand U20139 (N_20139,N_19599,N_19754);
nand U20140 (N_20140,N_19478,N_19426);
or U20141 (N_20141,N_19637,N_19679);
and U20142 (N_20142,N_19991,N_19730);
nand U20143 (N_20143,N_19990,N_19390);
nand U20144 (N_20144,N_19533,N_19499);
nor U20145 (N_20145,N_19950,N_19557);
and U20146 (N_20146,N_19664,N_19528);
nor U20147 (N_20147,N_19803,N_19674);
or U20148 (N_20148,N_19543,N_19809);
nor U20149 (N_20149,N_19818,N_19758);
nor U20150 (N_20150,N_19429,N_19404);
or U20151 (N_20151,N_19451,N_19861);
or U20152 (N_20152,N_19980,N_19470);
and U20153 (N_20153,N_19665,N_19536);
or U20154 (N_20154,N_19492,N_19949);
and U20155 (N_20155,N_19657,N_19804);
or U20156 (N_20156,N_19811,N_19504);
xor U20157 (N_20157,N_19436,N_19963);
or U20158 (N_20158,N_19654,N_19828);
or U20159 (N_20159,N_19630,N_19566);
nor U20160 (N_20160,N_19915,N_19520);
and U20161 (N_20161,N_19629,N_19452);
or U20162 (N_20162,N_19485,N_19924);
nor U20163 (N_20163,N_19987,N_19640);
xnor U20164 (N_20164,N_19947,N_19981);
nor U20165 (N_20165,N_19735,N_19918);
or U20166 (N_20166,N_19683,N_19869);
xnor U20167 (N_20167,N_19732,N_19530);
or U20168 (N_20168,N_19563,N_19585);
or U20169 (N_20169,N_19623,N_19728);
xor U20170 (N_20170,N_19597,N_19521);
and U20171 (N_20171,N_19391,N_19427);
nand U20172 (N_20172,N_19731,N_19387);
nand U20173 (N_20173,N_19707,N_19739);
and U20174 (N_20174,N_19671,N_19899);
xnor U20175 (N_20175,N_19618,N_19653);
nor U20176 (N_20176,N_19937,N_19797);
xnor U20177 (N_20177,N_19983,N_19479);
or U20178 (N_20178,N_19887,N_19900);
and U20179 (N_20179,N_19867,N_19857);
nand U20180 (N_20180,N_19896,N_19486);
nand U20181 (N_20181,N_19396,N_19511);
or U20182 (N_20182,N_19628,N_19742);
and U20183 (N_20183,N_19824,N_19660);
nand U20184 (N_20184,N_19668,N_19969);
and U20185 (N_20185,N_19607,N_19709);
and U20186 (N_20186,N_19948,N_19616);
or U20187 (N_20187,N_19941,N_19454);
nor U20188 (N_20188,N_19743,N_19909);
nor U20189 (N_20189,N_19706,N_19582);
and U20190 (N_20190,N_19737,N_19897);
nor U20191 (N_20191,N_19977,N_19823);
nand U20192 (N_20192,N_19393,N_19594);
or U20193 (N_20193,N_19488,N_19881);
nor U20194 (N_20194,N_19635,N_19562);
nand U20195 (N_20195,N_19548,N_19596);
xnor U20196 (N_20196,N_19854,N_19509);
nand U20197 (N_20197,N_19578,N_19569);
or U20198 (N_20198,N_19973,N_19740);
or U20199 (N_20199,N_19550,N_19889);
nor U20200 (N_20200,N_19761,N_19837);
nor U20201 (N_20201,N_19534,N_19482);
nand U20202 (N_20202,N_19782,N_19631);
nor U20203 (N_20203,N_19781,N_19834);
nand U20204 (N_20204,N_19956,N_19684);
nor U20205 (N_20205,N_19560,N_19976);
nor U20206 (N_20206,N_19440,N_19826);
nand U20207 (N_20207,N_19591,N_19652);
and U20208 (N_20208,N_19453,N_19764);
nor U20209 (N_20209,N_19838,N_19766);
nor U20210 (N_20210,N_19442,N_19999);
nor U20211 (N_20211,N_19438,N_19780);
or U20212 (N_20212,N_19588,N_19879);
or U20213 (N_20213,N_19694,N_19954);
or U20214 (N_20214,N_19416,N_19702);
nand U20215 (N_20215,N_19655,N_19675);
xnor U20216 (N_20216,N_19946,N_19587);
nand U20217 (N_20217,N_19645,N_19925);
nand U20218 (N_20218,N_19559,N_19968);
nand U20219 (N_20219,N_19501,N_19610);
and U20220 (N_20220,N_19984,N_19443);
nand U20221 (N_20221,N_19561,N_19884);
nand U20222 (N_20222,N_19407,N_19845);
and U20223 (N_20223,N_19468,N_19392);
and U20224 (N_20224,N_19813,N_19690);
nor U20225 (N_20225,N_19848,N_19771);
nand U20226 (N_20226,N_19484,N_19880);
and U20227 (N_20227,N_19719,N_19724);
nor U20228 (N_20228,N_19689,N_19472);
nor U20229 (N_20229,N_19401,N_19444);
nand U20230 (N_20230,N_19553,N_19783);
or U20231 (N_20231,N_19812,N_19994);
or U20232 (N_20232,N_19377,N_19409);
nand U20233 (N_20233,N_19982,N_19784);
nor U20234 (N_20234,N_19877,N_19997);
and U20235 (N_20235,N_19814,N_19641);
nor U20236 (N_20236,N_19698,N_19701);
nor U20237 (N_20237,N_19677,N_19920);
or U20238 (N_20238,N_19418,N_19866);
and U20239 (N_20239,N_19892,N_19627);
and U20240 (N_20240,N_19840,N_19883);
or U20241 (N_20241,N_19902,N_19609);
nor U20242 (N_20242,N_19540,N_19721);
nand U20243 (N_20243,N_19842,N_19535);
nor U20244 (N_20244,N_19508,N_19523);
nor U20245 (N_20245,N_19584,N_19801);
or U20246 (N_20246,N_19872,N_19474);
and U20247 (N_20247,N_19447,N_19388);
or U20248 (N_20248,N_19959,N_19862);
nor U20249 (N_20249,N_19514,N_19545);
nand U20250 (N_20250,N_19738,N_19750);
xnor U20251 (N_20251,N_19572,N_19676);
xnor U20252 (N_20252,N_19688,N_19799);
and U20253 (N_20253,N_19712,N_19894);
nand U20254 (N_20254,N_19498,N_19604);
and U20255 (N_20255,N_19806,N_19564);
and U20256 (N_20256,N_19605,N_19796);
and U20257 (N_20257,N_19952,N_19932);
nor U20258 (N_20258,N_19767,N_19757);
nand U20259 (N_20259,N_19944,N_19397);
or U20260 (N_20260,N_19988,N_19458);
nand U20261 (N_20261,N_19692,N_19644);
and U20262 (N_20262,N_19841,N_19419);
and U20263 (N_20263,N_19459,N_19768);
nor U20264 (N_20264,N_19792,N_19922);
and U20265 (N_20265,N_19914,N_19647);
or U20266 (N_20266,N_19589,N_19853);
or U20267 (N_20267,N_19775,N_19513);
and U20268 (N_20268,N_19691,N_19525);
and U20269 (N_20269,N_19425,N_19424);
and U20270 (N_20270,N_19512,N_19662);
or U20271 (N_20271,N_19620,N_19891);
nor U20272 (N_20272,N_19491,N_19704);
nand U20273 (N_20273,N_19441,N_19955);
or U20274 (N_20274,N_19455,N_19422);
nor U20275 (N_20275,N_19518,N_19851);
or U20276 (N_20276,N_19770,N_19964);
or U20277 (N_20277,N_19741,N_19752);
nand U20278 (N_20278,N_19552,N_19462);
nor U20279 (N_20279,N_19776,N_19624);
nor U20280 (N_20280,N_19423,N_19852);
and U20281 (N_20281,N_19744,N_19460);
nor U20282 (N_20282,N_19953,N_19993);
xor U20283 (N_20283,N_19827,N_19449);
or U20284 (N_20284,N_19966,N_19901);
xnor U20285 (N_20285,N_19936,N_19649);
xor U20286 (N_20286,N_19615,N_19515);
nor U20287 (N_20287,N_19437,N_19844);
or U20288 (N_20288,N_19434,N_19539);
or U20289 (N_20289,N_19906,N_19839);
nand U20290 (N_20290,N_19667,N_19747);
or U20291 (N_20291,N_19381,N_19890);
xor U20292 (N_20292,N_19720,N_19878);
and U20293 (N_20293,N_19751,N_19420);
nand U20294 (N_20294,N_19753,N_19965);
nand U20295 (N_20295,N_19579,N_19708);
nand U20296 (N_20296,N_19632,N_19795);
and U20297 (N_20297,N_19571,N_19678);
nor U20298 (N_20298,N_19913,N_19565);
or U20299 (N_20299,N_19703,N_19666);
nor U20300 (N_20300,N_19714,N_19636);
or U20301 (N_20301,N_19600,N_19575);
nor U20302 (N_20302,N_19945,N_19807);
nor U20303 (N_20303,N_19402,N_19893);
and U20304 (N_20304,N_19865,N_19446);
nor U20305 (N_20305,N_19505,N_19403);
or U20306 (N_20306,N_19816,N_19516);
nand U20307 (N_20307,N_19938,N_19939);
nand U20308 (N_20308,N_19992,N_19940);
nor U20309 (N_20309,N_19672,N_19850);
or U20310 (N_20310,N_19895,N_19957);
xnor U20311 (N_20311,N_19710,N_19821);
nor U20312 (N_20312,N_19682,N_19881);
nor U20313 (N_20313,N_19905,N_19711);
or U20314 (N_20314,N_19666,N_19608);
or U20315 (N_20315,N_19586,N_19635);
and U20316 (N_20316,N_19796,N_19402);
and U20317 (N_20317,N_19406,N_19656);
nand U20318 (N_20318,N_19870,N_19765);
nor U20319 (N_20319,N_19434,N_19965);
nand U20320 (N_20320,N_19911,N_19796);
nor U20321 (N_20321,N_19621,N_19720);
nand U20322 (N_20322,N_19985,N_19899);
xnor U20323 (N_20323,N_19779,N_19881);
or U20324 (N_20324,N_19818,N_19571);
nand U20325 (N_20325,N_19758,N_19893);
and U20326 (N_20326,N_19705,N_19807);
xnor U20327 (N_20327,N_19784,N_19778);
xnor U20328 (N_20328,N_19972,N_19575);
nand U20329 (N_20329,N_19906,N_19812);
or U20330 (N_20330,N_19619,N_19660);
or U20331 (N_20331,N_19851,N_19527);
or U20332 (N_20332,N_19609,N_19761);
nor U20333 (N_20333,N_19478,N_19459);
nor U20334 (N_20334,N_19403,N_19921);
nand U20335 (N_20335,N_19805,N_19826);
nor U20336 (N_20336,N_19986,N_19537);
nor U20337 (N_20337,N_19674,N_19848);
nor U20338 (N_20338,N_19798,N_19618);
xor U20339 (N_20339,N_19669,N_19597);
nor U20340 (N_20340,N_19836,N_19914);
nand U20341 (N_20341,N_19692,N_19666);
and U20342 (N_20342,N_19755,N_19396);
nor U20343 (N_20343,N_19832,N_19489);
nor U20344 (N_20344,N_19420,N_19739);
nand U20345 (N_20345,N_19677,N_19989);
or U20346 (N_20346,N_19431,N_19985);
nor U20347 (N_20347,N_19788,N_19980);
xnor U20348 (N_20348,N_19677,N_19383);
nor U20349 (N_20349,N_19619,N_19896);
and U20350 (N_20350,N_19475,N_19816);
nor U20351 (N_20351,N_19986,N_19812);
nand U20352 (N_20352,N_19680,N_19808);
nand U20353 (N_20353,N_19405,N_19963);
and U20354 (N_20354,N_19812,N_19774);
nand U20355 (N_20355,N_19574,N_19535);
or U20356 (N_20356,N_19465,N_19824);
nor U20357 (N_20357,N_19827,N_19476);
nand U20358 (N_20358,N_19874,N_19918);
xnor U20359 (N_20359,N_19787,N_19562);
nand U20360 (N_20360,N_19477,N_19858);
or U20361 (N_20361,N_19870,N_19479);
and U20362 (N_20362,N_19572,N_19388);
nand U20363 (N_20363,N_19949,N_19543);
or U20364 (N_20364,N_19491,N_19546);
nor U20365 (N_20365,N_19941,N_19700);
and U20366 (N_20366,N_19724,N_19615);
and U20367 (N_20367,N_19686,N_19566);
nor U20368 (N_20368,N_19651,N_19801);
and U20369 (N_20369,N_19513,N_19823);
and U20370 (N_20370,N_19608,N_19946);
and U20371 (N_20371,N_19391,N_19839);
or U20372 (N_20372,N_19851,N_19556);
nand U20373 (N_20373,N_19976,N_19634);
xnor U20374 (N_20374,N_19785,N_19953);
nor U20375 (N_20375,N_19653,N_19408);
nor U20376 (N_20376,N_19777,N_19520);
or U20377 (N_20377,N_19610,N_19612);
nor U20378 (N_20378,N_19522,N_19806);
and U20379 (N_20379,N_19864,N_19744);
and U20380 (N_20380,N_19900,N_19557);
nor U20381 (N_20381,N_19684,N_19947);
nor U20382 (N_20382,N_19376,N_19953);
or U20383 (N_20383,N_19883,N_19942);
or U20384 (N_20384,N_19865,N_19885);
or U20385 (N_20385,N_19863,N_19673);
nand U20386 (N_20386,N_19873,N_19864);
nor U20387 (N_20387,N_19680,N_19968);
nand U20388 (N_20388,N_19433,N_19424);
and U20389 (N_20389,N_19596,N_19496);
and U20390 (N_20390,N_19986,N_19861);
nor U20391 (N_20391,N_19607,N_19741);
and U20392 (N_20392,N_19455,N_19570);
nor U20393 (N_20393,N_19776,N_19552);
or U20394 (N_20394,N_19534,N_19400);
nor U20395 (N_20395,N_19926,N_19724);
nand U20396 (N_20396,N_19589,N_19609);
and U20397 (N_20397,N_19500,N_19518);
and U20398 (N_20398,N_19706,N_19636);
nand U20399 (N_20399,N_19701,N_19973);
nand U20400 (N_20400,N_19573,N_19611);
nand U20401 (N_20401,N_19714,N_19536);
nand U20402 (N_20402,N_19945,N_19793);
and U20403 (N_20403,N_19997,N_19454);
nand U20404 (N_20404,N_19652,N_19915);
or U20405 (N_20405,N_19773,N_19579);
or U20406 (N_20406,N_19761,N_19712);
nand U20407 (N_20407,N_19552,N_19928);
xnor U20408 (N_20408,N_19576,N_19973);
nand U20409 (N_20409,N_19559,N_19944);
or U20410 (N_20410,N_19500,N_19706);
and U20411 (N_20411,N_19376,N_19780);
nand U20412 (N_20412,N_19507,N_19792);
or U20413 (N_20413,N_19932,N_19777);
nand U20414 (N_20414,N_19464,N_19744);
and U20415 (N_20415,N_19599,N_19795);
xor U20416 (N_20416,N_19617,N_19882);
xnor U20417 (N_20417,N_19572,N_19834);
or U20418 (N_20418,N_19893,N_19770);
nand U20419 (N_20419,N_19985,N_19611);
and U20420 (N_20420,N_19773,N_19689);
or U20421 (N_20421,N_19891,N_19441);
and U20422 (N_20422,N_19450,N_19522);
and U20423 (N_20423,N_19710,N_19882);
xor U20424 (N_20424,N_19552,N_19839);
nor U20425 (N_20425,N_19769,N_19933);
nand U20426 (N_20426,N_19904,N_19924);
nand U20427 (N_20427,N_19462,N_19664);
nand U20428 (N_20428,N_19986,N_19690);
or U20429 (N_20429,N_19750,N_19634);
xnor U20430 (N_20430,N_19701,N_19645);
nor U20431 (N_20431,N_19948,N_19881);
nand U20432 (N_20432,N_19422,N_19774);
nand U20433 (N_20433,N_19838,N_19555);
nor U20434 (N_20434,N_19467,N_19869);
and U20435 (N_20435,N_19461,N_19670);
or U20436 (N_20436,N_19421,N_19782);
nand U20437 (N_20437,N_19706,N_19783);
or U20438 (N_20438,N_19559,N_19408);
nor U20439 (N_20439,N_19597,N_19788);
nor U20440 (N_20440,N_19592,N_19879);
and U20441 (N_20441,N_19911,N_19389);
nor U20442 (N_20442,N_19775,N_19776);
nor U20443 (N_20443,N_19434,N_19525);
or U20444 (N_20444,N_19875,N_19619);
nor U20445 (N_20445,N_19430,N_19836);
nand U20446 (N_20446,N_19674,N_19390);
and U20447 (N_20447,N_19460,N_19747);
nor U20448 (N_20448,N_19889,N_19593);
nand U20449 (N_20449,N_19436,N_19615);
or U20450 (N_20450,N_19958,N_19800);
or U20451 (N_20451,N_19538,N_19851);
nand U20452 (N_20452,N_19728,N_19954);
or U20453 (N_20453,N_19432,N_19573);
and U20454 (N_20454,N_19946,N_19961);
and U20455 (N_20455,N_19728,N_19567);
xnor U20456 (N_20456,N_19421,N_19988);
or U20457 (N_20457,N_19836,N_19617);
and U20458 (N_20458,N_19555,N_19469);
or U20459 (N_20459,N_19680,N_19884);
or U20460 (N_20460,N_19851,N_19479);
nand U20461 (N_20461,N_19725,N_19899);
nand U20462 (N_20462,N_19988,N_19893);
nor U20463 (N_20463,N_19861,N_19756);
or U20464 (N_20464,N_19981,N_19731);
nand U20465 (N_20465,N_19760,N_19989);
and U20466 (N_20466,N_19702,N_19462);
and U20467 (N_20467,N_19966,N_19699);
nor U20468 (N_20468,N_19509,N_19485);
nand U20469 (N_20469,N_19813,N_19720);
or U20470 (N_20470,N_19939,N_19528);
nor U20471 (N_20471,N_19602,N_19659);
or U20472 (N_20472,N_19775,N_19708);
and U20473 (N_20473,N_19780,N_19930);
or U20474 (N_20474,N_19415,N_19811);
nand U20475 (N_20475,N_19510,N_19593);
or U20476 (N_20476,N_19382,N_19537);
and U20477 (N_20477,N_19613,N_19733);
and U20478 (N_20478,N_19632,N_19563);
nor U20479 (N_20479,N_19963,N_19584);
nand U20480 (N_20480,N_19584,N_19964);
nand U20481 (N_20481,N_19578,N_19826);
nor U20482 (N_20482,N_19803,N_19565);
nand U20483 (N_20483,N_19986,N_19895);
and U20484 (N_20484,N_19792,N_19769);
nand U20485 (N_20485,N_19650,N_19938);
or U20486 (N_20486,N_19978,N_19634);
nor U20487 (N_20487,N_19705,N_19812);
nand U20488 (N_20488,N_19664,N_19826);
nor U20489 (N_20489,N_19473,N_19383);
xor U20490 (N_20490,N_19932,N_19971);
nand U20491 (N_20491,N_19866,N_19857);
or U20492 (N_20492,N_19434,N_19676);
nand U20493 (N_20493,N_19477,N_19580);
nor U20494 (N_20494,N_19810,N_19807);
and U20495 (N_20495,N_19852,N_19556);
and U20496 (N_20496,N_19975,N_19733);
and U20497 (N_20497,N_19383,N_19797);
nand U20498 (N_20498,N_19753,N_19484);
and U20499 (N_20499,N_19637,N_19751);
or U20500 (N_20500,N_19577,N_19843);
xor U20501 (N_20501,N_19638,N_19831);
nand U20502 (N_20502,N_19909,N_19409);
nor U20503 (N_20503,N_19575,N_19871);
or U20504 (N_20504,N_19444,N_19870);
nand U20505 (N_20505,N_19829,N_19631);
nor U20506 (N_20506,N_19523,N_19826);
nand U20507 (N_20507,N_19481,N_19561);
and U20508 (N_20508,N_19996,N_19558);
nand U20509 (N_20509,N_19387,N_19430);
and U20510 (N_20510,N_19390,N_19878);
and U20511 (N_20511,N_19569,N_19656);
nor U20512 (N_20512,N_19776,N_19985);
xnor U20513 (N_20513,N_19598,N_19516);
nand U20514 (N_20514,N_19798,N_19835);
or U20515 (N_20515,N_19654,N_19487);
or U20516 (N_20516,N_19403,N_19902);
or U20517 (N_20517,N_19710,N_19515);
or U20518 (N_20518,N_19901,N_19533);
xor U20519 (N_20519,N_19399,N_19590);
nor U20520 (N_20520,N_19519,N_19900);
xnor U20521 (N_20521,N_19801,N_19779);
nor U20522 (N_20522,N_19656,N_19746);
nor U20523 (N_20523,N_19832,N_19442);
nand U20524 (N_20524,N_19724,N_19825);
or U20525 (N_20525,N_19382,N_19587);
or U20526 (N_20526,N_19989,N_19679);
or U20527 (N_20527,N_19379,N_19831);
nor U20528 (N_20528,N_19420,N_19871);
nand U20529 (N_20529,N_19683,N_19849);
and U20530 (N_20530,N_19668,N_19377);
xnor U20531 (N_20531,N_19885,N_19715);
and U20532 (N_20532,N_19734,N_19460);
nand U20533 (N_20533,N_19469,N_19582);
nor U20534 (N_20534,N_19893,N_19763);
or U20535 (N_20535,N_19496,N_19999);
and U20536 (N_20536,N_19630,N_19757);
nor U20537 (N_20537,N_19554,N_19617);
and U20538 (N_20538,N_19530,N_19580);
nor U20539 (N_20539,N_19878,N_19817);
and U20540 (N_20540,N_19375,N_19441);
and U20541 (N_20541,N_19549,N_19818);
nand U20542 (N_20542,N_19877,N_19423);
nor U20543 (N_20543,N_19477,N_19904);
or U20544 (N_20544,N_19383,N_19455);
xor U20545 (N_20545,N_19471,N_19445);
nor U20546 (N_20546,N_19392,N_19849);
nor U20547 (N_20547,N_19976,N_19492);
xor U20548 (N_20548,N_19511,N_19679);
or U20549 (N_20549,N_19885,N_19804);
and U20550 (N_20550,N_19760,N_19847);
or U20551 (N_20551,N_19853,N_19851);
or U20552 (N_20552,N_19856,N_19850);
and U20553 (N_20553,N_19939,N_19947);
xnor U20554 (N_20554,N_19684,N_19691);
and U20555 (N_20555,N_19948,N_19574);
nand U20556 (N_20556,N_19640,N_19899);
or U20557 (N_20557,N_19688,N_19830);
nor U20558 (N_20558,N_19393,N_19739);
nor U20559 (N_20559,N_19774,N_19695);
and U20560 (N_20560,N_19733,N_19594);
or U20561 (N_20561,N_19531,N_19703);
nand U20562 (N_20562,N_19918,N_19961);
and U20563 (N_20563,N_19740,N_19506);
or U20564 (N_20564,N_19982,N_19654);
nor U20565 (N_20565,N_19754,N_19681);
nand U20566 (N_20566,N_19878,N_19407);
or U20567 (N_20567,N_19532,N_19918);
nand U20568 (N_20568,N_19422,N_19472);
and U20569 (N_20569,N_19450,N_19409);
xnor U20570 (N_20570,N_19376,N_19443);
nor U20571 (N_20571,N_19664,N_19761);
xor U20572 (N_20572,N_19621,N_19415);
xnor U20573 (N_20573,N_19399,N_19453);
nand U20574 (N_20574,N_19683,N_19524);
or U20575 (N_20575,N_19899,N_19938);
and U20576 (N_20576,N_19709,N_19695);
nand U20577 (N_20577,N_19571,N_19872);
nand U20578 (N_20578,N_19686,N_19940);
and U20579 (N_20579,N_19995,N_19994);
nor U20580 (N_20580,N_19686,N_19396);
and U20581 (N_20581,N_19646,N_19824);
and U20582 (N_20582,N_19630,N_19913);
xnor U20583 (N_20583,N_19696,N_19709);
or U20584 (N_20584,N_19573,N_19580);
or U20585 (N_20585,N_19891,N_19687);
nor U20586 (N_20586,N_19544,N_19878);
nor U20587 (N_20587,N_19609,N_19448);
nand U20588 (N_20588,N_19727,N_19662);
or U20589 (N_20589,N_19951,N_19807);
and U20590 (N_20590,N_19521,N_19535);
nor U20591 (N_20591,N_19869,N_19722);
nand U20592 (N_20592,N_19497,N_19494);
or U20593 (N_20593,N_19920,N_19591);
or U20594 (N_20594,N_19562,N_19962);
nand U20595 (N_20595,N_19413,N_19738);
xnor U20596 (N_20596,N_19742,N_19835);
and U20597 (N_20597,N_19808,N_19745);
nor U20598 (N_20598,N_19740,N_19776);
or U20599 (N_20599,N_19617,N_19701);
nand U20600 (N_20600,N_19637,N_19688);
or U20601 (N_20601,N_19798,N_19474);
and U20602 (N_20602,N_19822,N_19527);
or U20603 (N_20603,N_19826,N_19728);
and U20604 (N_20604,N_19540,N_19658);
nor U20605 (N_20605,N_19885,N_19846);
nand U20606 (N_20606,N_19494,N_19621);
nor U20607 (N_20607,N_19974,N_19588);
and U20608 (N_20608,N_19741,N_19964);
or U20609 (N_20609,N_19884,N_19529);
nand U20610 (N_20610,N_19803,N_19980);
nor U20611 (N_20611,N_19517,N_19564);
nand U20612 (N_20612,N_19961,N_19963);
or U20613 (N_20613,N_19561,N_19974);
xnor U20614 (N_20614,N_19766,N_19854);
or U20615 (N_20615,N_19738,N_19425);
nor U20616 (N_20616,N_19984,N_19818);
nand U20617 (N_20617,N_19904,N_19615);
nand U20618 (N_20618,N_19791,N_19943);
and U20619 (N_20619,N_19926,N_19942);
nand U20620 (N_20620,N_19751,N_19651);
nand U20621 (N_20621,N_19649,N_19732);
nand U20622 (N_20622,N_19626,N_19793);
or U20623 (N_20623,N_19956,N_19895);
xor U20624 (N_20624,N_19854,N_19579);
and U20625 (N_20625,N_20526,N_20105);
nor U20626 (N_20626,N_20051,N_20549);
nand U20627 (N_20627,N_20497,N_20534);
nor U20628 (N_20628,N_20562,N_20523);
nand U20629 (N_20629,N_20250,N_20594);
and U20630 (N_20630,N_20061,N_20425);
nand U20631 (N_20631,N_20010,N_20387);
or U20632 (N_20632,N_20037,N_20403);
nand U20633 (N_20633,N_20525,N_20266);
and U20634 (N_20634,N_20230,N_20527);
xnor U20635 (N_20635,N_20193,N_20217);
and U20636 (N_20636,N_20500,N_20186);
or U20637 (N_20637,N_20420,N_20557);
or U20638 (N_20638,N_20593,N_20034);
nor U20639 (N_20639,N_20498,N_20011);
nor U20640 (N_20640,N_20394,N_20097);
nor U20641 (N_20641,N_20530,N_20453);
and U20642 (N_20642,N_20089,N_20538);
nand U20643 (N_20643,N_20617,N_20203);
or U20644 (N_20644,N_20409,N_20091);
nor U20645 (N_20645,N_20030,N_20261);
nor U20646 (N_20646,N_20080,N_20590);
nand U20647 (N_20647,N_20431,N_20302);
and U20648 (N_20648,N_20023,N_20172);
nor U20649 (N_20649,N_20459,N_20361);
nor U20650 (N_20650,N_20402,N_20352);
nor U20651 (N_20651,N_20454,N_20422);
nor U20652 (N_20652,N_20062,N_20179);
xnor U20653 (N_20653,N_20492,N_20318);
nor U20654 (N_20654,N_20413,N_20157);
or U20655 (N_20655,N_20580,N_20390);
nor U20656 (N_20656,N_20301,N_20356);
nand U20657 (N_20657,N_20605,N_20595);
or U20658 (N_20658,N_20424,N_20095);
nor U20659 (N_20659,N_20188,N_20291);
nand U20660 (N_20660,N_20353,N_20311);
and U20661 (N_20661,N_20559,N_20385);
xnor U20662 (N_20662,N_20435,N_20572);
xor U20663 (N_20663,N_20084,N_20285);
or U20664 (N_20664,N_20587,N_20345);
nor U20665 (N_20665,N_20063,N_20620);
or U20666 (N_20666,N_20462,N_20111);
nand U20667 (N_20667,N_20423,N_20539);
and U20668 (N_20668,N_20624,N_20223);
nand U20669 (N_20669,N_20263,N_20322);
and U20670 (N_20670,N_20086,N_20357);
and U20671 (N_20671,N_20524,N_20441);
xor U20672 (N_20672,N_20005,N_20582);
or U20673 (N_20673,N_20430,N_20024);
nand U20674 (N_20674,N_20589,N_20270);
or U20675 (N_20675,N_20240,N_20437);
xnor U20676 (N_20676,N_20078,N_20451);
xor U20677 (N_20677,N_20503,N_20028);
nand U20678 (N_20678,N_20610,N_20260);
and U20679 (N_20679,N_20000,N_20211);
nor U20680 (N_20680,N_20143,N_20124);
or U20681 (N_20681,N_20540,N_20395);
or U20682 (N_20682,N_20146,N_20215);
and U20683 (N_20683,N_20228,N_20517);
nor U20684 (N_20684,N_20584,N_20579);
and U20685 (N_20685,N_20221,N_20476);
and U20686 (N_20686,N_20036,N_20128);
nor U20687 (N_20687,N_20252,N_20218);
and U20688 (N_20688,N_20119,N_20065);
xnor U20689 (N_20689,N_20110,N_20327);
nand U20690 (N_20690,N_20592,N_20253);
or U20691 (N_20691,N_20207,N_20458);
or U20692 (N_20692,N_20096,N_20281);
nor U20693 (N_20693,N_20484,N_20249);
or U20694 (N_20694,N_20478,N_20090);
and U20695 (N_20695,N_20310,N_20556);
nand U20696 (N_20696,N_20305,N_20055);
and U20697 (N_20697,N_20351,N_20543);
and U20698 (N_20698,N_20536,N_20265);
and U20699 (N_20699,N_20236,N_20112);
or U20700 (N_20700,N_20012,N_20209);
nor U20701 (N_20701,N_20474,N_20100);
or U20702 (N_20702,N_20528,N_20495);
nand U20703 (N_20703,N_20013,N_20502);
and U20704 (N_20704,N_20277,N_20212);
and U20705 (N_20705,N_20558,N_20093);
nand U20706 (N_20706,N_20337,N_20407);
or U20707 (N_20707,N_20449,N_20509);
and U20708 (N_20708,N_20033,N_20074);
nand U20709 (N_20709,N_20546,N_20308);
nor U20710 (N_20710,N_20537,N_20547);
nor U20711 (N_20711,N_20071,N_20513);
or U20712 (N_20712,N_20466,N_20241);
xor U20713 (N_20713,N_20622,N_20116);
nor U20714 (N_20714,N_20300,N_20101);
and U20715 (N_20715,N_20535,N_20306);
nor U20716 (N_20716,N_20205,N_20541);
nor U20717 (N_20717,N_20246,N_20088);
xnor U20718 (N_20718,N_20072,N_20032);
nand U20719 (N_20719,N_20552,N_20098);
nand U20720 (N_20720,N_20463,N_20312);
nand U20721 (N_20721,N_20383,N_20163);
nor U20722 (N_20722,N_20048,N_20297);
nand U20723 (N_20723,N_20464,N_20563);
xor U20724 (N_20724,N_20456,N_20204);
or U20725 (N_20725,N_20560,N_20280);
nand U20726 (N_20726,N_20512,N_20618);
nor U20727 (N_20727,N_20216,N_20450);
and U20728 (N_20728,N_20576,N_20248);
or U20729 (N_20729,N_20340,N_20288);
nand U20730 (N_20730,N_20542,N_20275);
nor U20731 (N_20731,N_20371,N_20410);
nand U20732 (N_20732,N_20338,N_20184);
nor U20733 (N_20733,N_20137,N_20069);
nor U20734 (N_20734,N_20170,N_20045);
nor U20735 (N_20735,N_20479,N_20104);
or U20736 (N_20736,N_20367,N_20355);
nand U20737 (N_20737,N_20173,N_20440);
or U20738 (N_20738,N_20370,N_20508);
nand U20739 (N_20739,N_20354,N_20247);
nand U20740 (N_20740,N_20398,N_20496);
or U20741 (N_20741,N_20548,N_20416);
nor U20742 (N_20742,N_20581,N_20133);
nand U20743 (N_20743,N_20405,N_20040);
or U20744 (N_20744,N_20177,N_20342);
nand U20745 (N_20745,N_20324,N_20279);
nor U20746 (N_20746,N_20309,N_20614);
xor U20747 (N_20747,N_20469,N_20446);
or U20748 (N_20748,N_20044,N_20166);
nand U20749 (N_20749,N_20384,N_20374);
nand U20750 (N_20750,N_20145,N_20434);
nor U20751 (N_20751,N_20234,N_20235);
and U20752 (N_20752,N_20152,N_20131);
and U20753 (N_20753,N_20057,N_20176);
and U20754 (N_20754,N_20368,N_20561);
xnor U20755 (N_20755,N_20489,N_20194);
xnor U20756 (N_20756,N_20391,N_20583);
nor U20757 (N_20757,N_20518,N_20411);
nor U20758 (N_20758,N_20317,N_20202);
nor U20759 (N_20759,N_20190,N_20251);
xor U20760 (N_20760,N_20130,N_20591);
nand U20761 (N_20761,N_20161,N_20075);
nand U20762 (N_20762,N_20118,N_20514);
nor U20763 (N_20763,N_20262,N_20003);
and U20764 (N_20764,N_20087,N_20292);
or U20765 (N_20765,N_20136,N_20363);
and U20766 (N_20766,N_20042,N_20602);
nor U20767 (N_20767,N_20243,N_20393);
nand U20768 (N_20768,N_20187,N_20213);
nor U20769 (N_20769,N_20482,N_20386);
and U20770 (N_20770,N_20019,N_20094);
and U20771 (N_20771,N_20196,N_20220);
or U20772 (N_20772,N_20477,N_20388);
nand U20773 (N_20773,N_20347,N_20531);
nor U20774 (N_20774,N_20330,N_20046);
nor U20775 (N_20775,N_20507,N_20522);
nor U20776 (N_20776,N_20007,N_20242);
xnor U20777 (N_20777,N_20227,N_20615);
nand U20778 (N_20778,N_20396,N_20117);
nor U20779 (N_20779,N_20397,N_20004);
nand U20780 (N_20780,N_20264,N_20171);
nand U20781 (N_20781,N_20232,N_20102);
nor U20782 (N_20782,N_20056,N_20596);
nor U20783 (N_20783,N_20376,N_20224);
and U20784 (N_20784,N_20533,N_20006);
or U20785 (N_20785,N_20021,N_20504);
nand U20786 (N_20786,N_20417,N_20429);
nand U20787 (N_20787,N_20486,N_20083);
or U20788 (N_20788,N_20226,N_20493);
and U20789 (N_20789,N_20321,N_20269);
nand U20790 (N_20790,N_20015,N_20287);
and U20791 (N_20791,N_20554,N_20331);
xor U20792 (N_20792,N_20490,N_20014);
nand U20793 (N_20793,N_20018,N_20127);
and U20794 (N_20794,N_20336,N_20341);
or U20795 (N_20795,N_20114,N_20471);
nor U20796 (N_20796,N_20494,N_20038);
nand U20797 (N_20797,N_20043,N_20284);
nand U20798 (N_20798,N_20457,N_20076);
or U20799 (N_20799,N_20609,N_20141);
and U20800 (N_20800,N_20016,N_20029);
nand U20801 (N_20801,N_20412,N_20569);
or U20802 (N_20802,N_20421,N_20132);
and U20803 (N_20803,N_20125,N_20577);
and U20804 (N_20804,N_20597,N_20229);
nand U20805 (N_20805,N_20467,N_20320);
nand U20806 (N_20806,N_20225,N_20169);
nor U20807 (N_20807,N_20077,N_20092);
and U20808 (N_20808,N_20178,N_20189);
nand U20809 (N_20809,N_20573,N_20392);
nor U20810 (N_20810,N_20551,N_20550);
nor U20811 (N_20811,N_20574,N_20017);
nor U20812 (N_20812,N_20427,N_20366);
and U20813 (N_20813,N_20295,N_20020);
nor U20814 (N_20814,N_20135,N_20233);
nor U20815 (N_20815,N_20373,N_20109);
xor U20816 (N_20816,N_20499,N_20578);
and U20817 (N_20817,N_20360,N_20025);
and U20818 (N_20818,N_20140,N_20245);
nand U20819 (N_20819,N_20505,N_20182);
nand U20820 (N_20820,N_20365,N_20162);
and U20821 (N_20821,N_20276,N_20159);
nor U20822 (N_20822,N_20002,N_20079);
nand U20823 (N_20823,N_20286,N_20439);
or U20824 (N_20824,N_20346,N_20185);
nand U20825 (N_20825,N_20568,N_20598);
or U20826 (N_20826,N_20139,N_20473);
and U20827 (N_20827,N_20520,N_20485);
nand U20828 (N_20828,N_20444,N_20231);
nor U20829 (N_20829,N_20611,N_20335);
or U20830 (N_20830,N_20468,N_20606);
and U20831 (N_20831,N_20399,N_20448);
and U20832 (N_20832,N_20001,N_20378);
xor U20833 (N_20833,N_20601,N_20294);
nand U20834 (N_20834,N_20142,N_20419);
nand U20835 (N_20835,N_20268,N_20604);
nand U20836 (N_20836,N_20181,N_20487);
and U20837 (N_20837,N_20326,N_20244);
and U20838 (N_20838,N_20623,N_20313);
nand U20839 (N_20839,N_20586,N_20304);
nand U20840 (N_20840,N_20465,N_20274);
nand U20841 (N_20841,N_20314,N_20027);
or U20842 (N_20842,N_20362,N_20257);
nand U20843 (N_20843,N_20208,N_20436);
nand U20844 (N_20844,N_20058,N_20447);
or U20845 (N_20845,N_20156,N_20035);
nand U20846 (N_20846,N_20299,N_20290);
nand U20847 (N_20847,N_20201,N_20359);
nor U20848 (N_20848,N_20039,N_20113);
and U20849 (N_20849,N_20588,N_20147);
nor U20850 (N_20850,N_20293,N_20258);
and U20851 (N_20851,N_20339,N_20401);
or U20852 (N_20852,N_20319,N_20283);
nand U20853 (N_20853,N_20067,N_20566);
xnor U20854 (N_20854,N_20372,N_20008);
and U20855 (N_20855,N_20047,N_20452);
or U20856 (N_20856,N_20480,N_20123);
nand U20857 (N_20857,N_20380,N_20344);
nor U20858 (N_20858,N_20348,N_20174);
or U20859 (N_20859,N_20155,N_20555);
and U20860 (N_20860,N_20064,N_20418);
or U20861 (N_20861,N_20271,N_20491);
and U20862 (N_20862,N_20315,N_20022);
xnor U20863 (N_20863,N_20455,N_20134);
or U20864 (N_20864,N_20350,N_20164);
nand U20865 (N_20865,N_20150,N_20379);
or U20866 (N_20866,N_20160,N_20404);
and U20867 (N_20867,N_20389,N_20041);
nor U20868 (N_20868,N_20107,N_20129);
nor U20869 (N_20869,N_20289,N_20607);
nor U20870 (N_20870,N_20103,N_20183);
nand U20871 (N_20871,N_20564,N_20068);
xor U20872 (N_20872,N_20445,N_20323);
nor U20873 (N_20873,N_20206,N_20238);
nand U20874 (N_20874,N_20049,N_20328);
nand U20875 (N_20875,N_20358,N_20278);
nor U20876 (N_20876,N_20099,N_20428);
or U20877 (N_20877,N_20481,N_20488);
or U20878 (N_20878,N_20603,N_20443);
or U20879 (N_20879,N_20219,N_20050);
nor U20880 (N_20880,N_20138,N_20108);
nand U20881 (N_20881,N_20126,N_20151);
nor U20882 (N_20882,N_20553,N_20198);
and U20883 (N_20883,N_20199,N_20545);
nand U20884 (N_20884,N_20195,N_20165);
nand U20885 (N_20885,N_20272,N_20613);
or U20886 (N_20886,N_20377,N_20121);
xor U20887 (N_20887,N_20438,N_20009);
and U20888 (N_20888,N_20599,N_20175);
and U20889 (N_20889,N_20433,N_20532);
nor U20890 (N_20890,N_20239,N_20364);
and U20891 (N_20891,N_20307,N_20608);
nand U20892 (N_20892,N_20511,N_20059);
nor U20893 (N_20893,N_20026,N_20567);
xnor U20894 (N_20894,N_20408,N_20325);
xor U20895 (N_20895,N_20149,N_20254);
and U20896 (N_20896,N_20120,N_20483);
nand U20897 (N_20897,N_20432,N_20516);
nor U20898 (N_20898,N_20316,N_20191);
nor U20899 (N_20899,N_20515,N_20400);
or U20900 (N_20900,N_20332,N_20461);
nor U20901 (N_20901,N_20472,N_20200);
and U20902 (N_20902,N_20470,N_20053);
or U20903 (N_20903,N_20296,N_20066);
nor U20904 (N_20904,N_20054,N_20158);
or U20905 (N_20905,N_20255,N_20369);
and U20906 (N_20906,N_20060,N_20214);
nand U20907 (N_20907,N_20267,N_20475);
nor U20908 (N_20908,N_20167,N_20329);
and U20909 (N_20909,N_20154,N_20600);
or U20910 (N_20910,N_20621,N_20585);
and U20911 (N_20911,N_20381,N_20460);
xor U20912 (N_20912,N_20081,N_20616);
nand U20913 (N_20913,N_20349,N_20180);
or U20914 (N_20914,N_20073,N_20273);
or U20915 (N_20915,N_20521,N_20619);
or U20916 (N_20916,N_20501,N_20298);
nand U20917 (N_20917,N_20343,N_20506);
xnor U20918 (N_20918,N_20510,N_20575);
nand U20919 (N_20919,N_20197,N_20122);
xor U20920 (N_20920,N_20031,N_20334);
nand U20921 (N_20921,N_20222,N_20148);
nor U20922 (N_20922,N_20192,N_20070);
and U20923 (N_20923,N_20612,N_20406);
nand U20924 (N_20924,N_20259,N_20375);
nand U20925 (N_20925,N_20442,N_20571);
or U20926 (N_20926,N_20085,N_20153);
nand U20927 (N_20927,N_20082,N_20282);
nand U20928 (N_20928,N_20426,N_20237);
nor U20929 (N_20929,N_20519,N_20544);
nor U20930 (N_20930,N_20115,N_20303);
and U20931 (N_20931,N_20106,N_20529);
and U20932 (N_20932,N_20415,N_20168);
and U20933 (N_20933,N_20333,N_20565);
nor U20934 (N_20934,N_20414,N_20052);
and U20935 (N_20935,N_20210,N_20256);
nand U20936 (N_20936,N_20570,N_20144);
xor U20937 (N_20937,N_20382,N_20129);
nand U20938 (N_20938,N_20517,N_20335);
nand U20939 (N_20939,N_20339,N_20341);
nand U20940 (N_20940,N_20285,N_20185);
and U20941 (N_20941,N_20478,N_20097);
and U20942 (N_20942,N_20471,N_20078);
nor U20943 (N_20943,N_20145,N_20465);
or U20944 (N_20944,N_20174,N_20224);
or U20945 (N_20945,N_20359,N_20019);
or U20946 (N_20946,N_20061,N_20417);
nor U20947 (N_20947,N_20304,N_20130);
nand U20948 (N_20948,N_20076,N_20264);
nor U20949 (N_20949,N_20330,N_20183);
and U20950 (N_20950,N_20233,N_20144);
nor U20951 (N_20951,N_20572,N_20287);
nand U20952 (N_20952,N_20367,N_20495);
or U20953 (N_20953,N_20031,N_20320);
nand U20954 (N_20954,N_20160,N_20545);
nor U20955 (N_20955,N_20190,N_20466);
nor U20956 (N_20956,N_20002,N_20393);
and U20957 (N_20957,N_20274,N_20539);
nor U20958 (N_20958,N_20280,N_20162);
or U20959 (N_20959,N_20355,N_20253);
nor U20960 (N_20960,N_20504,N_20405);
nand U20961 (N_20961,N_20171,N_20117);
and U20962 (N_20962,N_20199,N_20250);
nor U20963 (N_20963,N_20350,N_20401);
nor U20964 (N_20964,N_20427,N_20076);
or U20965 (N_20965,N_20585,N_20060);
or U20966 (N_20966,N_20149,N_20597);
nand U20967 (N_20967,N_20466,N_20194);
nand U20968 (N_20968,N_20076,N_20081);
and U20969 (N_20969,N_20256,N_20068);
or U20970 (N_20970,N_20286,N_20575);
nor U20971 (N_20971,N_20437,N_20021);
nor U20972 (N_20972,N_20489,N_20054);
nor U20973 (N_20973,N_20043,N_20374);
xnor U20974 (N_20974,N_20598,N_20405);
nor U20975 (N_20975,N_20036,N_20262);
and U20976 (N_20976,N_20243,N_20331);
nor U20977 (N_20977,N_20428,N_20478);
and U20978 (N_20978,N_20287,N_20340);
or U20979 (N_20979,N_20513,N_20344);
nor U20980 (N_20980,N_20301,N_20220);
nand U20981 (N_20981,N_20506,N_20473);
and U20982 (N_20982,N_20484,N_20123);
nor U20983 (N_20983,N_20612,N_20036);
nand U20984 (N_20984,N_20421,N_20100);
and U20985 (N_20985,N_20412,N_20193);
nor U20986 (N_20986,N_20133,N_20142);
or U20987 (N_20987,N_20371,N_20050);
and U20988 (N_20988,N_20103,N_20250);
nor U20989 (N_20989,N_20565,N_20205);
nand U20990 (N_20990,N_20266,N_20579);
nor U20991 (N_20991,N_20125,N_20414);
and U20992 (N_20992,N_20155,N_20498);
nor U20993 (N_20993,N_20552,N_20020);
and U20994 (N_20994,N_20231,N_20251);
nor U20995 (N_20995,N_20414,N_20290);
and U20996 (N_20996,N_20226,N_20338);
nor U20997 (N_20997,N_20158,N_20055);
and U20998 (N_20998,N_20619,N_20318);
nand U20999 (N_20999,N_20503,N_20157);
nand U21000 (N_21000,N_20194,N_20373);
and U21001 (N_21001,N_20530,N_20255);
nand U21002 (N_21002,N_20385,N_20319);
xnor U21003 (N_21003,N_20361,N_20422);
and U21004 (N_21004,N_20434,N_20080);
and U21005 (N_21005,N_20367,N_20187);
nand U21006 (N_21006,N_20468,N_20356);
nor U21007 (N_21007,N_20157,N_20561);
or U21008 (N_21008,N_20582,N_20303);
and U21009 (N_21009,N_20295,N_20002);
nor U21010 (N_21010,N_20490,N_20515);
and U21011 (N_21011,N_20318,N_20254);
nor U21012 (N_21012,N_20360,N_20295);
or U21013 (N_21013,N_20272,N_20072);
and U21014 (N_21014,N_20158,N_20104);
or U21015 (N_21015,N_20242,N_20273);
nor U21016 (N_21016,N_20485,N_20127);
xnor U21017 (N_21017,N_20346,N_20165);
nor U21018 (N_21018,N_20490,N_20477);
nand U21019 (N_21019,N_20514,N_20541);
xor U21020 (N_21020,N_20282,N_20060);
or U21021 (N_21021,N_20122,N_20148);
nor U21022 (N_21022,N_20066,N_20156);
and U21023 (N_21023,N_20460,N_20468);
or U21024 (N_21024,N_20178,N_20572);
xnor U21025 (N_21025,N_20228,N_20104);
nor U21026 (N_21026,N_20309,N_20397);
nand U21027 (N_21027,N_20360,N_20205);
and U21028 (N_21028,N_20215,N_20383);
or U21029 (N_21029,N_20251,N_20252);
nand U21030 (N_21030,N_20484,N_20054);
nor U21031 (N_21031,N_20008,N_20252);
nand U21032 (N_21032,N_20457,N_20392);
and U21033 (N_21033,N_20062,N_20593);
nand U21034 (N_21034,N_20603,N_20000);
nand U21035 (N_21035,N_20204,N_20137);
nor U21036 (N_21036,N_20574,N_20443);
xnor U21037 (N_21037,N_20431,N_20048);
and U21038 (N_21038,N_20609,N_20538);
nor U21039 (N_21039,N_20158,N_20412);
nand U21040 (N_21040,N_20510,N_20475);
or U21041 (N_21041,N_20602,N_20129);
or U21042 (N_21042,N_20570,N_20246);
nor U21043 (N_21043,N_20015,N_20388);
and U21044 (N_21044,N_20104,N_20429);
nand U21045 (N_21045,N_20449,N_20412);
or U21046 (N_21046,N_20611,N_20169);
xnor U21047 (N_21047,N_20179,N_20549);
nand U21048 (N_21048,N_20454,N_20443);
and U21049 (N_21049,N_20011,N_20284);
nor U21050 (N_21050,N_20017,N_20000);
xor U21051 (N_21051,N_20281,N_20457);
and U21052 (N_21052,N_20406,N_20534);
or U21053 (N_21053,N_20115,N_20415);
nor U21054 (N_21054,N_20242,N_20378);
and U21055 (N_21055,N_20476,N_20217);
nor U21056 (N_21056,N_20037,N_20173);
nor U21057 (N_21057,N_20535,N_20295);
nor U21058 (N_21058,N_20040,N_20362);
nand U21059 (N_21059,N_20010,N_20131);
nor U21060 (N_21060,N_20524,N_20221);
nor U21061 (N_21061,N_20344,N_20174);
or U21062 (N_21062,N_20345,N_20056);
or U21063 (N_21063,N_20341,N_20277);
and U21064 (N_21064,N_20624,N_20486);
nor U21065 (N_21065,N_20156,N_20464);
and U21066 (N_21066,N_20071,N_20155);
nor U21067 (N_21067,N_20563,N_20130);
or U21068 (N_21068,N_20159,N_20401);
xor U21069 (N_21069,N_20514,N_20395);
nand U21070 (N_21070,N_20448,N_20479);
and U21071 (N_21071,N_20138,N_20348);
or U21072 (N_21072,N_20038,N_20345);
xnor U21073 (N_21073,N_20274,N_20216);
or U21074 (N_21074,N_20078,N_20061);
nor U21075 (N_21075,N_20589,N_20447);
nor U21076 (N_21076,N_20241,N_20130);
nor U21077 (N_21077,N_20556,N_20315);
and U21078 (N_21078,N_20059,N_20375);
nor U21079 (N_21079,N_20555,N_20414);
xnor U21080 (N_21080,N_20236,N_20104);
nor U21081 (N_21081,N_20435,N_20551);
and U21082 (N_21082,N_20033,N_20137);
and U21083 (N_21083,N_20243,N_20189);
nand U21084 (N_21084,N_20409,N_20396);
nand U21085 (N_21085,N_20196,N_20525);
xor U21086 (N_21086,N_20192,N_20099);
nand U21087 (N_21087,N_20448,N_20296);
or U21088 (N_21088,N_20033,N_20301);
or U21089 (N_21089,N_20176,N_20618);
or U21090 (N_21090,N_20088,N_20321);
and U21091 (N_21091,N_20524,N_20151);
nand U21092 (N_21092,N_20198,N_20583);
nor U21093 (N_21093,N_20216,N_20512);
nor U21094 (N_21094,N_20026,N_20561);
or U21095 (N_21095,N_20044,N_20214);
xnor U21096 (N_21096,N_20574,N_20090);
or U21097 (N_21097,N_20279,N_20104);
nand U21098 (N_21098,N_20477,N_20056);
or U21099 (N_21099,N_20588,N_20140);
nand U21100 (N_21100,N_20062,N_20368);
or U21101 (N_21101,N_20301,N_20556);
nor U21102 (N_21102,N_20516,N_20422);
nor U21103 (N_21103,N_20385,N_20579);
and U21104 (N_21104,N_20098,N_20022);
nand U21105 (N_21105,N_20475,N_20175);
and U21106 (N_21106,N_20187,N_20546);
nand U21107 (N_21107,N_20401,N_20082);
nand U21108 (N_21108,N_20563,N_20516);
and U21109 (N_21109,N_20332,N_20579);
and U21110 (N_21110,N_20456,N_20085);
nor U21111 (N_21111,N_20110,N_20575);
xnor U21112 (N_21112,N_20464,N_20568);
and U21113 (N_21113,N_20436,N_20538);
or U21114 (N_21114,N_20230,N_20272);
nor U21115 (N_21115,N_20608,N_20401);
and U21116 (N_21116,N_20184,N_20000);
nor U21117 (N_21117,N_20490,N_20534);
or U21118 (N_21118,N_20093,N_20529);
or U21119 (N_21119,N_20048,N_20261);
xor U21120 (N_21120,N_20168,N_20307);
nor U21121 (N_21121,N_20458,N_20612);
xnor U21122 (N_21122,N_20474,N_20406);
xnor U21123 (N_21123,N_20085,N_20602);
nand U21124 (N_21124,N_20309,N_20056);
nor U21125 (N_21125,N_20507,N_20478);
nand U21126 (N_21126,N_20399,N_20162);
nand U21127 (N_21127,N_20206,N_20177);
and U21128 (N_21128,N_20434,N_20216);
or U21129 (N_21129,N_20174,N_20145);
or U21130 (N_21130,N_20404,N_20415);
nor U21131 (N_21131,N_20241,N_20409);
nand U21132 (N_21132,N_20021,N_20458);
and U21133 (N_21133,N_20584,N_20227);
xnor U21134 (N_21134,N_20231,N_20098);
xor U21135 (N_21135,N_20556,N_20460);
or U21136 (N_21136,N_20061,N_20031);
or U21137 (N_21137,N_20435,N_20491);
and U21138 (N_21138,N_20178,N_20548);
nor U21139 (N_21139,N_20377,N_20623);
nor U21140 (N_21140,N_20243,N_20420);
nand U21141 (N_21141,N_20584,N_20142);
xnor U21142 (N_21142,N_20178,N_20017);
nand U21143 (N_21143,N_20611,N_20360);
and U21144 (N_21144,N_20384,N_20379);
or U21145 (N_21145,N_20500,N_20260);
nand U21146 (N_21146,N_20315,N_20242);
nand U21147 (N_21147,N_20616,N_20041);
or U21148 (N_21148,N_20219,N_20222);
nor U21149 (N_21149,N_20417,N_20296);
nand U21150 (N_21150,N_20614,N_20298);
and U21151 (N_21151,N_20612,N_20470);
nand U21152 (N_21152,N_20162,N_20473);
or U21153 (N_21153,N_20616,N_20410);
and U21154 (N_21154,N_20165,N_20462);
or U21155 (N_21155,N_20255,N_20344);
and U21156 (N_21156,N_20398,N_20119);
xor U21157 (N_21157,N_20507,N_20203);
and U21158 (N_21158,N_20405,N_20214);
and U21159 (N_21159,N_20033,N_20341);
nand U21160 (N_21160,N_20191,N_20574);
or U21161 (N_21161,N_20163,N_20335);
nor U21162 (N_21162,N_20324,N_20392);
and U21163 (N_21163,N_20616,N_20548);
nor U21164 (N_21164,N_20459,N_20203);
nor U21165 (N_21165,N_20361,N_20563);
nand U21166 (N_21166,N_20495,N_20118);
or U21167 (N_21167,N_20157,N_20209);
nand U21168 (N_21168,N_20331,N_20463);
nor U21169 (N_21169,N_20423,N_20519);
or U21170 (N_21170,N_20310,N_20418);
nor U21171 (N_21171,N_20375,N_20340);
or U21172 (N_21172,N_20251,N_20057);
or U21173 (N_21173,N_20034,N_20238);
or U21174 (N_21174,N_20133,N_20476);
xor U21175 (N_21175,N_20096,N_20289);
nor U21176 (N_21176,N_20317,N_20275);
nand U21177 (N_21177,N_20193,N_20521);
nand U21178 (N_21178,N_20116,N_20068);
nand U21179 (N_21179,N_20338,N_20390);
and U21180 (N_21180,N_20003,N_20059);
or U21181 (N_21181,N_20301,N_20198);
and U21182 (N_21182,N_20203,N_20473);
or U21183 (N_21183,N_20419,N_20274);
nor U21184 (N_21184,N_20275,N_20199);
nand U21185 (N_21185,N_20376,N_20024);
and U21186 (N_21186,N_20237,N_20099);
and U21187 (N_21187,N_20435,N_20596);
nand U21188 (N_21188,N_20566,N_20563);
and U21189 (N_21189,N_20356,N_20365);
and U21190 (N_21190,N_20048,N_20216);
and U21191 (N_21191,N_20569,N_20475);
nor U21192 (N_21192,N_20580,N_20199);
nor U21193 (N_21193,N_20221,N_20579);
or U21194 (N_21194,N_20150,N_20262);
xnor U21195 (N_21195,N_20339,N_20195);
nor U21196 (N_21196,N_20265,N_20556);
nor U21197 (N_21197,N_20500,N_20582);
and U21198 (N_21198,N_20202,N_20129);
nor U21199 (N_21199,N_20618,N_20029);
nand U21200 (N_21200,N_20354,N_20557);
and U21201 (N_21201,N_20304,N_20354);
nand U21202 (N_21202,N_20565,N_20219);
xor U21203 (N_21203,N_20486,N_20160);
xor U21204 (N_21204,N_20560,N_20145);
or U21205 (N_21205,N_20450,N_20055);
or U21206 (N_21206,N_20047,N_20417);
or U21207 (N_21207,N_20072,N_20339);
and U21208 (N_21208,N_20612,N_20372);
or U21209 (N_21209,N_20165,N_20588);
nor U21210 (N_21210,N_20160,N_20496);
xnor U21211 (N_21211,N_20242,N_20344);
and U21212 (N_21212,N_20450,N_20603);
or U21213 (N_21213,N_20140,N_20201);
nand U21214 (N_21214,N_20078,N_20361);
or U21215 (N_21215,N_20083,N_20195);
nor U21216 (N_21216,N_20233,N_20210);
nand U21217 (N_21217,N_20434,N_20144);
nor U21218 (N_21218,N_20328,N_20339);
xnor U21219 (N_21219,N_20507,N_20609);
or U21220 (N_21220,N_20072,N_20114);
or U21221 (N_21221,N_20299,N_20557);
nand U21222 (N_21222,N_20350,N_20580);
nand U21223 (N_21223,N_20518,N_20595);
nor U21224 (N_21224,N_20366,N_20187);
nand U21225 (N_21225,N_20462,N_20484);
nand U21226 (N_21226,N_20238,N_20240);
xor U21227 (N_21227,N_20130,N_20619);
nor U21228 (N_21228,N_20545,N_20267);
nor U21229 (N_21229,N_20445,N_20208);
nor U21230 (N_21230,N_20512,N_20533);
and U21231 (N_21231,N_20140,N_20203);
nor U21232 (N_21232,N_20033,N_20265);
nand U21233 (N_21233,N_20524,N_20428);
and U21234 (N_21234,N_20184,N_20515);
or U21235 (N_21235,N_20238,N_20073);
nor U21236 (N_21236,N_20299,N_20395);
nand U21237 (N_21237,N_20027,N_20616);
nand U21238 (N_21238,N_20365,N_20140);
nor U21239 (N_21239,N_20130,N_20546);
nor U21240 (N_21240,N_20105,N_20246);
nand U21241 (N_21241,N_20519,N_20039);
nor U21242 (N_21242,N_20569,N_20112);
and U21243 (N_21243,N_20084,N_20423);
nand U21244 (N_21244,N_20158,N_20519);
nor U21245 (N_21245,N_20314,N_20233);
nor U21246 (N_21246,N_20149,N_20286);
and U21247 (N_21247,N_20593,N_20479);
and U21248 (N_21248,N_20357,N_20087);
and U21249 (N_21249,N_20017,N_20316);
or U21250 (N_21250,N_21063,N_21172);
and U21251 (N_21251,N_20911,N_21020);
or U21252 (N_21252,N_20880,N_21129);
or U21253 (N_21253,N_20847,N_21030);
or U21254 (N_21254,N_20765,N_21083);
nor U21255 (N_21255,N_20906,N_20939);
nand U21256 (N_21256,N_21173,N_20874);
and U21257 (N_21257,N_20640,N_21061);
or U21258 (N_21258,N_21033,N_20648);
nor U21259 (N_21259,N_20698,N_20793);
or U21260 (N_21260,N_20785,N_20689);
and U21261 (N_21261,N_21140,N_20644);
and U21262 (N_21262,N_20659,N_21054);
nand U21263 (N_21263,N_20842,N_20916);
nor U21264 (N_21264,N_20780,N_21000);
and U21265 (N_21265,N_20650,N_21060);
nor U21266 (N_21266,N_21157,N_20828);
and U21267 (N_21267,N_20786,N_20773);
or U21268 (N_21268,N_21124,N_20895);
and U21269 (N_21269,N_20669,N_21099);
and U21270 (N_21270,N_20989,N_20998);
nand U21271 (N_21271,N_20812,N_20695);
and U21272 (N_21272,N_20743,N_21170);
nand U21273 (N_21273,N_20917,N_21088);
nor U21274 (N_21274,N_20902,N_20735);
and U21275 (N_21275,N_21199,N_21016);
nand U21276 (N_21276,N_21220,N_20837);
nand U21277 (N_21277,N_20870,N_20725);
or U21278 (N_21278,N_21235,N_20719);
nor U21279 (N_21279,N_21153,N_20711);
nand U21280 (N_21280,N_21209,N_21028);
and U21281 (N_21281,N_21069,N_20927);
nand U21282 (N_21282,N_21219,N_20886);
or U21283 (N_21283,N_20807,N_21085);
nor U21284 (N_21284,N_20871,N_21026);
nand U21285 (N_21285,N_20676,N_21107);
nor U21286 (N_21286,N_20996,N_21150);
nor U21287 (N_21287,N_20991,N_21188);
nand U21288 (N_21288,N_21064,N_21077);
or U21289 (N_21289,N_21213,N_21087);
xor U21290 (N_21290,N_20816,N_20701);
nand U21291 (N_21291,N_20954,N_20899);
nand U21292 (N_21292,N_20737,N_20943);
xor U21293 (N_21293,N_21056,N_20855);
nor U21294 (N_21294,N_21136,N_20882);
nor U21295 (N_21295,N_21242,N_20801);
nand U21296 (N_21296,N_21142,N_20746);
and U21297 (N_21297,N_20741,N_21146);
nor U21298 (N_21298,N_20873,N_20814);
nor U21299 (N_21299,N_20818,N_21053);
nor U21300 (N_21300,N_21217,N_20684);
nand U21301 (N_21301,N_20716,N_21108);
or U21302 (N_21302,N_20962,N_20833);
nand U21303 (N_21303,N_21223,N_20730);
nor U21304 (N_21304,N_21196,N_20686);
nand U21305 (N_21305,N_20969,N_20979);
nand U21306 (N_21306,N_20789,N_21071);
nand U21307 (N_21307,N_20849,N_21134);
and U21308 (N_21308,N_21174,N_21074);
nand U21309 (N_21309,N_20736,N_21101);
and U21310 (N_21310,N_20769,N_21021);
nand U21311 (N_21311,N_20688,N_20952);
and U21312 (N_21312,N_21078,N_21132);
and U21313 (N_21313,N_20715,N_21097);
or U21314 (N_21314,N_20885,N_20663);
nand U21315 (N_21315,N_20915,N_21232);
or U21316 (N_21316,N_21103,N_20845);
or U21317 (N_21317,N_20888,N_21156);
and U21318 (N_21318,N_20657,N_20784);
xor U21319 (N_21319,N_21158,N_20710);
nand U21320 (N_21320,N_21149,N_20980);
and U21321 (N_21321,N_20848,N_20850);
nor U21322 (N_21322,N_21043,N_20727);
nand U21323 (N_21323,N_21143,N_20664);
and U21324 (N_21324,N_20709,N_20950);
nor U21325 (N_21325,N_20700,N_21072);
nor U21326 (N_21326,N_20791,N_20973);
nor U21327 (N_21327,N_20632,N_21159);
or U21328 (N_21328,N_20796,N_20660);
nand U21329 (N_21329,N_21169,N_20827);
and U21330 (N_21330,N_20779,N_20752);
nand U21331 (N_21331,N_20909,N_21148);
nand U21332 (N_21332,N_20907,N_20914);
nor U21333 (N_21333,N_21104,N_21047);
and U21334 (N_21334,N_21122,N_21234);
and U21335 (N_21335,N_21094,N_21125);
nor U21336 (N_21336,N_20639,N_20966);
xnor U21337 (N_21337,N_20953,N_20681);
xnor U21338 (N_21338,N_20921,N_20908);
nand U21339 (N_21339,N_20815,N_21160);
xnor U21340 (N_21340,N_20750,N_21175);
or U21341 (N_21341,N_20795,N_20932);
nor U21342 (N_21342,N_21012,N_20731);
and U21343 (N_21343,N_20758,N_20840);
or U21344 (N_21344,N_21068,N_20658);
nand U21345 (N_21345,N_20949,N_20775);
nand U21346 (N_21346,N_20697,N_21184);
or U21347 (N_21347,N_21168,N_20651);
or U21348 (N_21348,N_21230,N_21163);
or U21349 (N_21349,N_21203,N_20628);
or U21350 (N_21350,N_21066,N_20728);
and U21351 (N_21351,N_20724,N_21073);
nand U21352 (N_21352,N_21067,N_20878);
nor U21353 (N_21353,N_20692,N_20889);
or U21354 (N_21354,N_20699,N_20654);
and U21355 (N_21355,N_20708,N_20768);
and U21356 (N_21356,N_20783,N_20682);
nor U21357 (N_21357,N_21001,N_21154);
xor U21358 (N_21358,N_20830,N_20971);
xor U21359 (N_21359,N_21014,N_21100);
xor U21360 (N_21360,N_20643,N_21240);
xor U21361 (N_21361,N_20981,N_21191);
nand U21362 (N_21362,N_21008,N_20819);
and U21363 (N_21363,N_20920,N_21095);
or U21364 (N_21364,N_20972,N_21005);
or U21365 (N_21365,N_21098,N_20852);
or U21366 (N_21366,N_20685,N_20987);
and U21367 (N_21367,N_20649,N_21227);
nand U21368 (N_21368,N_21057,N_20668);
or U21369 (N_21369,N_20672,N_21070);
xor U21370 (N_21370,N_20673,N_20729);
nor U21371 (N_21371,N_21086,N_20985);
and U21372 (N_21372,N_20670,N_21215);
and U21373 (N_21373,N_21007,N_21206);
and U21374 (N_21374,N_20679,N_21137);
nand U21375 (N_21375,N_20997,N_20748);
nand U21376 (N_21376,N_20900,N_21145);
or U21377 (N_21377,N_20875,N_21241);
or U21378 (N_21378,N_21109,N_20762);
and U21379 (N_21379,N_20763,N_20963);
xor U21380 (N_21380,N_20674,N_20897);
and U21381 (N_21381,N_20806,N_20732);
xor U21382 (N_21382,N_21018,N_20820);
nand U21383 (N_21383,N_20829,N_21115);
nor U21384 (N_21384,N_20778,N_20714);
and U21385 (N_21385,N_21027,N_21116);
and U21386 (N_21386,N_20945,N_20804);
and U21387 (N_21387,N_20744,N_21035);
and U21388 (N_21388,N_20792,N_20753);
nand U21389 (N_21389,N_20931,N_20671);
nand U21390 (N_21390,N_20937,N_20890);
or U21391 (N_21391,N_20879,N_20821);
nor U21392 (N_21392,N_21198,N_20754);
nor U21393 (N_21393,N_20799,N_20721);
xor U21394 (N_21394,N_20696,N_20788);
or U21395 (N_21395,N_20687,N_21092);
or U21396 (N_21396,N_20690,N_20790);
or U21397 (N_21397,N_20956,N_20771);
nand U21398 (N_21398,N_20905,N_20983);
nor U21399 (N_21399,N_21167,N_21197);
nand U21400 (N_21400,N_21046,N_20782);
and U21401 (N_21401,N_20861,N_20707);
nand U21402 (N_21402,N_20957,N_20755);
or U21403 (N_21403,N_20893,N_20946);
nand U21404 (N_21404,N_20993,N_20802);
xnor U21405 (N_21405,N_21050,N_21237);
nand U21406 (N_21406,N_21229,N_21238);
nor U21407 (N_21407,N_20960,N_20910);
and U21408 (N_21408,N_20968,N_20898);
nor U21409 (N_21409,N_20922,N_21089);
nand U21410 (N_21410,N_20913,N_21102);
or U21411 (N_21411,N_21222,N_20720);
nand U21412 (N_21412,N_21013,N_20839);
or U21413 (N_21413,N_21091,N_20817);
or U21414 (N_21414,N_20635,N_21200);
nand U21415 (N_21415,N_21009,N_20662);
nand U21416 (N_21416,N_20683,N_20749);
or U21417 (N_21417,N_21201,N_21032);
nor U21418 (N_21418,N_20666,N_20675);
and U21419 (N_21419,N_20838,N_20928);
nand U21420 (N_21420,N_21080,N_20767);
nor U21421 (N_21421,N_21117,N_20631);
or U21422 (N_21422,N_21055,N_20843);
or U21423 (N_21423,N_20941,N_21189);
or U21424 (N_21424,N_20887,N_21178);
xor U21425 (N_21425,N_20646,N_20661);
or U21426 (N_21426,N_21131,N_21042);
and U21427 (N_21427,N_21212,N_21226);
and U21428 (N_21428,N_21176,N_21161);
nor U21429 (N_21429,N_21155,N_20706);
and U21430 (N_21430,N_21133,N_20901);
and U21431 (N_21431,N_20713,N_20722);
or U21432 (N_21432,N_21211,N_21040);
nand U21433 (N_21433,N_20860,N_20726);
and U21434 (N_21434,N_21128,N_20733);
and U21435 (N_21435,N_20824,N_20854);
nand U21436 (N_21436,N_20717,N_20936);
and U21437 (N_21437,N_20857,N_21221);
and U21438 (N_21438,N_21119,N_20877);
xnor U21439 (N_21439,N_20680,N_20761);
nor U21440 (N_21440,N_21185,N_21059);
and U21441 (N_21441,N_21166,N_20864);
xor U21442 (N_21442,N_20794,N_20923);
and U21443 (N_21443,N_21048,N_20844);
and U21444 (N_21444,N_20809,N_20800);
or U21445 (N_21445,N_20652,N_20653);
and U21446 (N_21446,N_20693,N_21224);
nand U21447 (N_21447,N_21243,N_20777);
nand U21448 (N_21448,N_21110,N_20940);
nand U21449 (N_21449,N_20863,N_21180);
and U21450 (N_21450,N_21049,N_20951);
and U21451 (N_21451,N_21147,N_21138);
and U21452 (N_21452,N_20865,N_21084);
and U21453 (N_21453,N_20665,N_20647);
and U21454 (N_21454,N_21171,N_20846);
and U21455 (N_21455,N_20826,N_20787);
or U21456 (N_21456,N_20667,N_21023);
nand U21457 (N_21457,N_20772,N_21195);
and U21458 (N_21458,N_20770,N_21111);
and U21459 (N_21459,N_20919,N_20964);
xnor U21460 (N_21460,N_20625,N_20944);
xnor U21461 (N_21461,N_20740,N_21210);
xor U21462 (N_21462,N_21202,N_21123);
or U21463 (N_21463,N_20869,N_20891);
nand U21464 (N_21464,N_21231,N_21082);
nor U21465 (N_21465,N_20756,N_20984);
xnor U21466 (N_21466,N_20976,N_21062);
nand U21467 (N_21467,N_20942,N_20862);
and U21468 (N_21468,N_21118,N_20704);
nand U21469 (N_21469,N_20745,N_20645);
and U21470 (N_21470,N_20867,N_21105);
nand U21471 (N_21471,N_20641,N_21245);
and U21472 (N_21472,N_20766,N_21044);
and U21473 (N_21473,N_20866,N_20823);
and U21474 (N_21474,N_21152,N_21216);
nor U21475 (N_21475,N_21004,N_21187);
nand U21476 (N_21476,N_21041,N_21236);
nand U21477 (N_21477,N_20892,N_21003);
or U21478 (N_21478,N_21031,N_21190);
and U21479 (N_21479,N_21205,N_20859);
xnor U21480 (N_21480,N_20933,N_20884);
xnor U21481 (N_21481,N_21076,N_20831);
nand U21482 (N_21482,N_20961,N_20811);
or U21483 (N_21483,N_21052,N_21193);
nand U21484 (N_21484,N_21096,N_20982);
nand U21485 (N_21485,N_20894,N_21246);
nand U21486 (N_21486,N_20938,N_21214);
nor U21487 (N_21487,N_20856,N_20738);
nor U21488 (N_21488,N_20974,N_20896);
nor U21489 (N_21489,N_20924,N_21228);
and U21490 (N_21490,N_20970,N_21186);
or U21491 (N_21491,N_20836,N_21114);
nand U21492 (N_21492,N_21090,N_21139);
or U21493 (N_21493,N_20925,N_20760);
nand U21494 (N_21494,N_20832,N_21079);
or U21495 (N_21495,N_21051,N_20718);
and U21496 (N_21496,N_20904,N_20926);
or U21497 (N_21497,N_21151,N_20723);
xnor U21498 (N_21498,N_21075,N_20813);
nand U21499 (N_21499,N_20764,N_21218);
nor U21500 (N_21500,N_20703,N_20678);
xnor U21501 (N_21501,N_20995,N_21164);
nand U21502 (N_21502,N_21113,N_20691);
xor U21503 (N_21503,N_21022,N_20986);
and U21504 (N_21504,N_20851,N_21127);
or U21505 (N_21505,N_20903,N_20822);
nor U21506 (N_21506,N_20677,N_20978);
and U21507 (N_21507,N_20988,N_20834);
nor U21508 (N_21508,N_21239,N_21106);
nand U21509 (N_21509,N_21038,N_21162);
or U21510 (N_21510,N_20712,N_20637);
or U21511 (N_21511,N_21225,N_20739);
or U21512 (N_21512,N_20694,N_20881);
or U21513 (N_21513,N_20872,N_20705);
nand U21514 (N_21514,N_21192,N_20934);
nand U21515 (N_21515,N_21182,N_21194);
nor U21516 (N_21516,N_21029,N_20975);
or U21517 (N_21517,N_21019,N_20853);
or U21518 (N_21518,N_20990,N_21025);
nand U21519 (N_21519,N_21006,N_20965);
nor U21520 (N_21520,N_20929,N_20734);
or U21521 (N_21521,N_20994,N_20912);
nand U21522 (N_21522,N_21208,N_21002);
and U21523 (N_21523,N_21081,N_20999);
xnor U21524 (N_21524,N_21144,N_20947);
or U21525 (N_21525,N_21247,N_21165);
nand U21526 (N_21526,N_20958,N_21065);
nor U21527 (N_21527,N_20759,N_20805);
and U21528 (N_21528,N_21249,N_20918);
and U21529 (N_21529,N_20803,N_20992);
nand U21530 (N_21530,N_20747,N_20629);
nor U21531 (N_21531,N_20774,N_20967);
or U21532 (N_21532,N_20955,N_20656);
nand U21533 (N_21533,N_20876,N_21036);
or U21534 (N_21534,N_20810,N_21120);
or U21535 (N_21535,N_20808,N_21034);
nand U21536 (N_21536,N_20776,N_20627);
nand U21537 (N_21537,N_20757,N_20702);
nor U21538 (N_21538,N_21130,N_20883);
nand U21539 (N_21539,N_20634,N_21017);
or U21540 (N_21540,N_21024,N_20825);
nor U21541 (N_21541,N_21011,N_21204);
nand U21542 (N_21542,N_20626,N_20781);
and U21543 (N_21543,N_20977,N_21177);
or U21544 (N_21544,N_21112,N_21037);
and U21545 (N_21545,N_21093,N_21045);
and U21546 (N_21546,N_20633,N_20638);
or U21547 (N_21547,N_20930,N_21015);
nor U21548 (N_21548,N_21058,N_21135);
nand U21549 (N_21549,N_20959,N_20630);
or U21550 (N_21550,N_20751,N_21207);
nand U21551 (N_21551,N_20797,N_21141);
nand U21552 (N_21552,N_21010,N_21181);
or U21553 (N_21553,N_21126,N_20655);
or U21554 (N_21554,N_21244,N_20835);
and U21555 (N_21555,N_20798,N_21183);
or U21556 (N_21556,N_20858,N_21233);
or U21557 (N_21557,N_20642,N_21179);
or U21558 (N_21558,N_20742,N_21039);
nand U21559 (N_21559,N_20935,N_20841);
and U21560 (N_21560,N_21121,N_20636);
nand U21561 (N_21561,N_20948,N_21248);
or U21562 (N_21562,N_20868,N_20983);
and U21563 (N_21563,N_20958,N_21159);
nand U21564 (N_21564,N_21248,N_20777);
nor U21565 (N_21565,N_20826,N_20951);
nand U21566 (N_21566,N_21016,N_20651);
nor U21567 (N_21567,N_21117,N_20810);
nand U21568 (N_21568,N_20906,N_20736);
and U21569 (N_21569,N_21245,N_21102);
and U21570 (N_21570,N_20929,N_21180);
or U21571 (N_21571,N_21241,N_20682);
nand U21572 (N_21572,N_20789,N_20863);
nand U21573 (N_21573,N_20652,N_20955);
and U21574 (N_21574,N_21196,N_20719);
nand U21575 (N_21575,N_21148,N_20806);
or U21576 (N_21576,N_21022,N_21235);
nor U21577 (N_21577,N_20781,N_21176);
or U21578 (N_21578,N_20730,N_21151);
and U21579 (N_21579,N_21164,N_21119);
or U21580 (N_21580,N_20816,N_20705);
nor U21581 (N_21581,N_21080,N_21005);
and U21582 (N_21582,N_20763,N_21070);
xnor U21583 (N_21583,N_20790,N_21166);
or U21584 (N_21584,N_20840,N_20783);
nand U21585 (N_21585,N_21170,N_20837);
nor U21586 (N_21586,N_20662,N_21136);
or U21587 (N_21587,N_21155,N_20833);
xnor U21588 (N_21588,N_21198,N_20696);
or U21589 (N_21589,N_21121,N_20728);
and U21590 (N_21590,N_21043,N_20630);
xnor U21591 (N_21591,N_21234,N_20871);
xnor U21592 (N_21592,N_20807,N_20673);
or U21593 (N_21593,N_20860,N_20840);
or U21594 (N_21594,N_21163,N_20699);
nor U21595 (N_21595,N_21219,N_20817);
nand U21596 (N_21596,N_20908,N_20756);
nor U21597 (N_21597,N_21031,N_21088);
or U21598 (N_21598,N_20681,N_21048);
nand U21599 (N_21599,N_20650,N_20774);
xnor U21600 (N_21600,N_21010,N_20913);
and U21601 (N_21601,N_21088,N_20828);
nand U21602 (N_21602,N_20911,N_21182);
nand U21603 (N_21603,N_21023,N_20880);
and U21604 (N_21604,N_20675,N_20626);
and U21605 (N_21605,N_20686,N_21043);
nor U21606 (N_21606,N_20840,N_21108);
and U21607 (N_21607,N_21159,N_20993);
nand U21608 (N_21608,N_20886,N_20626);
nand U21609 (N_21609,N_21159,N_21224);
nand U21610 (N_21610,N_20685,N_21197);
and U21611 (N_21611,N_20627,N_20775);
or U21612 (N_21612,N_20842,N_20724);
or U21613 (N_21613,N_21030,N_21246);
and U21614 (N_21614,N_20962,N_20913);
and U21615 (N_21615,N_20946,N_21104);
nor U21616 (N_21616,N_21142,N_20871);
nor U21617 (N_21617,N_20983,N_21222);
nor U21618 (N_21618,N_21162,N_20724);
and U21619 (N_21619,N_20982,N_20792);
nand U21620 (N_21620,N_20997,N_20638);
or U21621 (N_21621,N_20842,N_21004);
nor U21622 (N_21622,N_21063,N_21114);
or U21623 (N_21623,N_20915,N_20861);
nand U21624 (N_21624,N_20738,N_21003);
nor U21625 (N_21625,N_20961,N_20684);
and U21626 (N_21626,N_21020,N_21014);
nand U21627 (N_21627,N_21157,N_21119);
or U21628 (N_21628,N_21021,N_20762);
or U21629 (N_21629,N_21039,N_20944);
nor U21630 (N_21630,N_20712,N_20767);
xor U21631 (N_21631,N_21119,N_21022);
and U21632 (N_21632,N_21204,N_20710);
and U21633 (N_21633,N_20727,N_21174);
nor U21634 (N_21634,N_20666,N_21006);
nor U21635 (N_21635,N_20654,N_20963);
and U21636 (N_21636,N_20854,N_20889);
or U21637 (N_21637,N_20935,N_21107);
nand U21638 (N_21638,N_20661,N_20766);
xor U21639 (N_21639,N_20736,N_20638);
and U21640 (N_21640,N_20742,N_21017);
and U21641 (N_21641,N_20787,N_20642);
nand U21642 (N_21642,N_21198,N_20907);
nor U21643 (N_21643,N_21226,N_21008);
or U21644 (N_21644,N_20934,N_21105);
or U21645 (N_21645,N_20853,N_20956);
and U21646 (N_21646,N_20780,N_21141);
or U21647 (N_21647,N_21129,N_21142);
xnor U21648 (N_21648,N_20906,N_21243);
or U21649 (N_21649,N_20873,N_20714);
nand U21650 (N_21650,N_20844,N_20786);
nor U21651 (N_21651,N_20863,N_20797);
nor U21652 (N_21652,N_21000,N_20750);
xor U21653 (N_21653,N_20887,N_21213);
nand U21654 (N_21654,N_20750,N_20671);
or U21655 (N_21655,N_21163,N_20924);
nand U21656 (N_21656,N_20873,N_20961);
or U21657 (N_21657,N_21003,N_20703);
or U21658 (N_21658,N_20674,N_20884);
or U21659 (N_21659,N_21231,N_20806);
nor U21660 (N_21660,N_21090,N_20951);
nor U21661 (N_21661,N_21082,N_20825);
nor U21662 (N_21662,N_21015,N_20678);
xor U21663 (N_21663,N_21103,N_21133);
or U21664 (N_21664,N_20819,N_20906);
nand U21665 (N_21665,N_20810,N_20852);
nand U21666 (N_21666,N_21129,N_20903);
nand U21667 (N_21667,N_20910,N_21015);
and U21668 (N_21668,N_21056,N_21189);
or U21669 (N_21669,N_20803,N_20761);
and U21670 (N_21670,N_21076,N_21040);
nand U21671 (N_21671,N_21021,N_20682);
or U21672 (N_21672,N_21121,N_20815);
nand U21673 (N_21673,N_20660,N_20671);
nand U21674 (N_21674,N_20845,N_20894);
or U21675 (N_21675,N_21205,N_20968);
nor U21676 (N_21676,N_20719,N_21247);
nor U21677 (N_21677,N_20945,N_21246);
nor U21678 (N_21678,N_21247,N_20954);
nand U21679 (N_21679,N_21099,N_21224);
nor U21680 (N_21680,N_21116,N_21036);
nor U21681 (N_21681,N_21236,N_20874);
and U21682 (N_21682,N_20633,N_20760);
or U21683 (N_21683,N_21212,N_21058);
or U21684 (N_21684,N_20725,N_20692);
or U21685 (N_21685,N_20886,N_20726);
or U21686 (N_21686,N_21160,N_21014);
nand U21687 (N_21687,N_20960,N_21210);
nand U21688 (N_21688,N_20737,N_20975);
xor U21689 (N_21689,N_20778,N_20986);
nand U21690 (N_21690,N_20964,N_20778);
nor U21691 (N_21691,N_20792,N_21199);
xor U21692 (N_21692,N_21066,N_20825);
xor U21693 (N_21693,N_21078,N_21128);
or U21694 (N_21694,N_21100,N_21163);
nor U21695 (N_21695,N_20790,N_21065);
nand U21696 (N_21696,N_20775,N_20833);
nand U21697 (N_21697,N_20805,N_20945);
xor U21698 (N_21698,N_20761,N_20648);
or U21699 (N_21699,N_20650,N_20929);
and U21700 (N_21700,N_20721,N_20659);
and U21701 (N_21701,N_21161,N_21077);
or U21702 (N_21702,N_21110,N_21115);
xnor U21703 (N_21703,N_20869,N_21039);
nor U21704 (N_21704,N_20946,N_21224);
nand U21705 (N_21705,N_21099,N_20959);
or U21706 (N_21706,N_20954,N_20836);
nand U21707 (N_21707,N_20859,N_21091);
nand U21708 (N_21708,N_20793,N_20707);
xor U21709 (N_21709,N_20669,N_21106);
or U21710 (N_21710,N_20661,N_21172);
and U21711 (N_21711,N_21024,N_20920);
nand U21712 (N_21712,N_20987,N_20757);
xnor U21713 (N_21713,N_20631,N_21057);
nand U21714 (N_21714,N_20632,N_21045);
and U21715 (N_21715,N_20858,N_20839);
and U21716 (N_21716,N_21168,N_21136);
xnor U21717 (N_21717,N_20794,N_21231);
nand U21718 (N_21718,N_20901,N_21238);
nor U21719 (N_21719,N_20930,N_20872);
and U21720 (N_21720,N_20780,N_20979);
nor U21721 (N_21721,N_20971,N_20834);
and U21722 (N_21722,N_21224,N_20966);
nor U21723 (N_21723,N_20784,N_20909);
nor U21724 (N_21724,N_20696,N_20898);
or U21725 (N_21725,N_21171,N_20637);
xnor U21726 (N_21726,N_21139,N_21068);
nand U21727 (N_21727,N_20928,N_20637);
or U21728 (N_21728,N_20930,N_20726);
and U21729 (N_21729,N_20856,N_20896);
or U21730 (N_21730,N_20772,N_20694);
nand U21731 (N_21731,N_20904,N_21077);
nand U21732 (N_21732,N_21215,N_20992);
nand U21733 (N_21733,N_20721,N_21171);
nor U21734 (N_21734,N_21224,N_20967);
nor U21735 (N_21735,N_20630,N_21203);
nand U21736 (N_21736,N_20696,N_20762);
and U21737 (N_21737,N_21042,N_20724);
or U21738 (N_21738,N_20950,N_20915);
nand U21739 (N_21739,N_21216,N_20866);
xnor U21740 (N_21740,N_20872,N_21135);
xnor U21741 (N_21741,N_21016,N_20760);
nand U21742 (N_21742,N_21176,N_20998);
and U21743 (N_21743,N_20733,N_21127);
nand U21744 (N_21744,N_20950,N_21161);
nor U21745 (N_21745,N_20733,N_21066);
and U21746 (N_21746,N_20765,N_21207);
nor U21747 (N_21747,N_21109,N_21142);
or U21748 (N_21748,N_21134,N_21091);
xnor U21749 (N_21749,N_20649,N_21221);
or U21750 (N_21750,N_20788,N_20821);
nor U21751 (N_21751,N_20962,N_21224);
and U21752 (N_21752,N_20813,N_20987);
nand U21753 (N_21753,N_21053,N_20875);
and U21754 (N_21754,N_20998,N_20897);
nand U21755 (N_21755,N_21052,N_21074);
nand U21756 (N_21756,N_20701,N_21065);
nand U21757 (N_21757,N_21195,N_21077);
nor U21758 (N_21758,N_20811,N_20933);
nor U21759 (N_21759,N_20959,N_21051);
nand U21760 (N_21760,N_20750,N_20667);
and U21761 (N_21761,N_21045,N_20971);
xor U21762 (N_21762,N_21071,N_21223);
or U21763 (N_21763,N_20760,N_20929);
nand U21764 (N_21764,N_20641,N_21228);
nand U21765 (N_21765,N_20968,N_20953);
or U21766 (N_21766,N_20687,N_21073);
nand U21767 (N_21767,N_20838,N_21154);
nand U21768 (N_21768,N_21195,N_20631);
nand U21769 (N_21769,N_21018,N_21197);
nand U21770 (N_21770,N_20886,N_20806);
nor U21771 (N_21771,N_20661,N_20665);
or U21772 (N_21772,N_20978,N_21212);
nand U21773 (N_21773,N_21131,N_21180);
nand U21774 (N_21774,N_21154,N_20811);
nand U21775 (N_21775,N_21242,N_20815);
xor U21776 (N_21776,N_20664,N_21074);
or U21777 (N_21777,N_20906,N_20891);
or U21778 (N_21778,N_20971,N_20785);
and U21779 (N_21779,N_21064,N_20883);
xor U21780 (N_21780,N_20750,N_20926);
and U21781 (N_21781,N_21095,N_20753);
or U21782 (N_21782,N_20678,N_21108);
or U21783 (N_21783,N_21215,N_20927);
and U21784 (N_21784,N_20934,N_21131);
nand U21785 (N_21785,N_21061,N_20906);
or U21786 (N_21786,N_20672,N_20995);
or U21787 (N_21787,N_20962,N_20767);
or U21788 (N_21788,N_20805,N_20730);
nor U21789 (N_21789,N_20991,N_21169);
nand U21790 (N_21790,N_20799,N_20759);
nand U21791 (N_21791,N_21212,N_21091);
or U21792 (N_21792,N_21020,N_20792);
and U21793 (N_21793,N_21057,N_21242);
and U21794 (N_21794,N_20663,N_20991);
nor U21795 (N_21795,N_21138,N_20807);
and U21796 (N_21796,N_21035,N_21164);
xor U21797 (N_21797,N_20731,N_20714);
or U21798 (N_21798,N_21163,N_20909);
and U21799 (N_21799,N_20654,N_21184);
or U21800 (N_21800,N_20916,N_21065);
and U21801 (N_21801,N_21091,N_21138);
or U21802 (N_21802,N_21233,N_20970);
xor U21803 (N_21803,N_21006,N_20981);
nand U21804 (N_21804,N_20796,N_20782);
or U21805 (N_21805,N_20752,N_20790);
and U21806 (N_21806,N_20764,N_20892);
nand U21807 (N_21807,N_21070,N_20647);
nand U21808 (N_21808,N_20716,N_21164);
nor U21809 (N_21809,N_20649,N_21057);
nor U21810 (N_21810,N_20648,N_20814);
nor U21811 (N_21811,N_20714,N_20687);
xnor U21812 (N_21812,N_21187,N_20940);
nor U21813 (N_21813,N_21086,N_21248);
and U21814 (N_21814,N_21019,N_21039);
and U21815 (N_21815,N_20933,N_20862);
nand U21816 (N_21816,N_21167,N_20916);
nor U21817 (N_21817,N_21035,N_21208);
nand U21818 (N_21818,N_20695,N_21231);
and U21819 (N_21819,N_20846,N_20813);
and U21820 (N_21820,N_20941,N_21025);
or U21821 (N_21821,N_21013,N_20902);
nor U21822 (N_21822,N_20986,N_20946);
nor U21823 (N_21823,N_20857,N_20780);
xnor U21824 (N_21824,N_20632,N_20947);
nand U21825 (N_21825,N_20647,N_20893);
nand U21826 (N_21826,N_20834,N_21120);
xor U21827 (N_21827,N_20735,N_20707);
or U21828 (N_21828,N_20632,N_21208);
and U21829 (N_21829,N_21000,N_20627);
nand U21830 (N_21830,N_20742,N_21048);
nand U21831 (N_21831,N_21058,N_20927);
nand U21832 (N_21832,N_20723,N_20703);
nor U21833 (N_21833,N_20753,N_21178);
or U21834 (N_21834,N_20654,N_20705);
or U21835 (N_21835,N_21193,N_21005);
nor U21836 (N_21836,N_20651,N_21156);
nor U21837 (N_21837,N_21040,N_21005);
or U21838 (N_21838,N_20807,N_20657);
nand U21839 (N_21839,N_20839,N_20894);
nand U21840 (N_21840,N_21079,N_20951);
nand U21841 (N_21841,N_21044,N_21177);
nor U21842 (N_21842,N_21022,N_20744);
or U21843 (N_21843,N_20928,N_21104);
or U21844 (N_21844,N_21082,N_21194);
or U21845 (N_21845,N_20962,N_20961);
nand U21846 (N_21846,N_20713,N_20888);
nor U21847 (N_21847,N_20653,N_21214);
and U21848 (N_21848,N_21153,N_20959);
and U21849 (N_21849,N_21242,N_20669);
nor U21850 (N_21850,N_20873,N_21189);
and U21851 (N_21851,N_21019,N_20903);
and U21852 (N_21852,N_21162,N_20739);
nand U21853 (N_21853,N_20673,N_20649);
xnor U21854 (N_21854,N_21117,N_20699);
and U21855 (N_21855,N_21022,N_20885);
and U21856 (N_21856,N_20897,N_20892);
nand U21857 (N_21857,N_20925,N_21090);
or U21858 (N_21858,N_20790,N_21107);
and U21859 (N_21859,N_20716,N_20815);
xnor U21860 (N_21860,N_20996,N_21047);
and U21861 (N_21861,N_21058,N_20818);
nor U21862 (N_21862,N_21233,N_20784);
nor U21863 (N_21863,N_21006,N_20667);
and U21864 (N_21864,N_20680,N_20750);
or U21865 (N_21865,N_21018,N_21237);
or U21866 (N_21866,N_20666,N_21152);
or U21867 (N_21867,N_21010,N_21194);
or U21868 (N_21868,N_21000,N_21172);
xnor U21869 (N_21869,N_20807,N_20839);
nand U21870 (N_21870,N_20921,N_20824);
nand U21871 (N_21871,N_21082,N_21059);
and U21872 (N_21872,N_21078,N_21024);
nor U21873 (N_21873,N_21043,N_20918);
xor U21874 (N_21874,N_20731,N_21213);
nand U21875 (N_21875,N_21724,N_21855);
or U21876 (N_21876,N_21513,N_21866);
nand U21877 (N_21877,N_21275,N_21569);
nor U21878 (N_21878,N_21350,N_21388);
nand U21879 (N_21879,N_21540,N_21771);
and U21880 (N_21880,N_21726,N_21788);
nand U21881 (N_21881,N_21523,N_21475);
xor U21882 (N_21882,N_21799,N_21666);
and U21883 (N_21883,N_21349,N_21425);
nand U21884 (N_21884,N_21426,N_21452);
and U21885 (N_21885,N_21618,N_21541);
nand U21886 (N_21886,N_21692,N_21339);
nor U21887 (N_21887,N_21585,N_21579);
xor U21888 (N_21888,N_21770,N_21826);
or U21889 (N_21889,N_21838,N_21645);
nand U21890 (N_21890,N_21470,N_21636);
and U21891 (N_21891,N_21577,N_21710);
nor U21892 (N_21892,N_21264,N_21443);
nor U21893 (N_21893,N_21345,N_21730);
nand U21894 (N_21894,N_21688,N_21564);
nand U21895 (N_21895,N_21520,N_21252);
nor U21896 (N_21896,N_21632,N_21832);
nand U21897 (N_21897,N_21760,N_21572);
nor U21898 (N_21898,N_21422,N_21630);
xor U21899 (N_21899,N_21595,N_21790);
or U21900 (N_21900,N_21481,N_21846);
nand U21901 (N_21901,N_21453,N_21720);
and U21902 (N_21902,N_21365,N_21816);
nand U21903 (N_21903,N_21483,N_21288);
nor U21904 (N_21904,N_21505,N_21712);
nor U21905 (N_21905,N_21690,N_21567);
and U21906 (N_21906,N_21717,N_21491);
nor U21907 (N_21907,N_21874,N_21589);
xor U21908 (N_21908,N_21695,N_21303);
or U21909 (N_21909,N_21551,N_21741);
and U21910 (N_21910,N_21411,N_21665);
nor U21911 (N_21911,N_21508,N_21667);
or U21912 (N_21912,N_21620,N_21829);
xnor U21913 (N_21913,N_21313,N_21344);
nor U21914 (N_21914,N_21278,N_21265);
nand U21915 (N_21915,N_21335,N_21496);
or U21916 (N_21916,N_21756,N_21650);
or U21917 (N_21917,N_21458,N_21831);
xnor U21918 (N_21918,N_21609,N_21260);
nor U21919 (N_21919,N_21372,N_21798);
or U21920 (N_21920,N_21291,N_21573);
nor U21921 (N_21921,N_21644,N_21522);
nand U21922 (N_21922,N_21765,N_21836);
and U21923 (N_21923,N_21530,N_21869);
nand U21924 (N_21924,N_21328,N_21758);
and U21925 (N_21925,N_21525,N_21557);
nand U21926 (N_21926,N_21616,N_21800);
or U21927 (N_21927,N_21423,N_21787);
or U21928 (N_21928,N_21696,N_21697);
and U21929 (N_21929,N_21818,N_21814);
nand U21930 (N_21930,N_21600,N_21333);
nand U21931 (N_21931,N_21506,N_21659);
nor U21932 (N_21932,N_21612,N_21773);
or U21933 (N_21933,N_21719,N_21369);
nor U21934 (N_21934,N_21524,N_21646);
or U21935 (N_21935,N_21619,N_21542);
and U21936 (N_21936,N_21387,N_21466);
or U21937 (N_21937,N_21509,N_21873);
xor U21938 (N_21938,N_21307,N_21680);
xnor U21939 (N_21939,N_21329,N_21316);
nor U21940 (N_21940,N_21601,N_21324);
and U21941 (N_21941,N_21497,N_21368);
nand U21942 (N_21942,N_21471,N_21849);
nor U21943 (N_21943,N_21521,N_21830);
nand U21944 (N_21944,N_21539,N_21456);
and U21945 (N_21945,N_21427,N_21574);
xor U21946 (N_21946,N_21317,N_21767);
and U21947 (N_21947,N_21312,N_21267);
nor U21948 (N_21948,N_21416,N_21362);
xor U21949 (N_21949,N_21780,N_21708);
and U21950 (N_21950,N_21559,N_21704);
or U21951 (N_21951,N_21686,N_21581);
nand U21952 (N_21952,N_21858,N_21759);
or U21953 (N_21953,N_21562,N_21584);
xnor U21954 (N_21954,N_21725,N_21284);
or U21955 (N_21955,N_21627,N_21872);
nor U21956 (N_21956,N_21446,N_21621);
or U21957 (N_21957,N_21392,N_21462);
nor U21958 (N_21958,N_21682,N_21319);
nand U21959 (N_21959,N_21555,N_21500);
xnor U21960 (N_21960,N_21401,N_21702);
nor U21961 (N_21961,N_21840,N_21430);
and U21962 (N_21962,N_21852,N_21824);
or U21963 (N_21963,N_21499,N_21810);
nand U21964 (N_21964,N_21651,N_21827);
nand U21965 (N_21965,N_21380,N_21683);
xnor U21966 (N_21966,N_21611,N_21781);
or U21967 (N_21967,N_21352,N_21763);
nand U21968 (N_21968,N_21862,N_21635);
and U21969 (N_21969,N_21302,N_21463);
nand U21970 (N_21970,N_21480,N_21703);
and U21971 (N_21971,N_21280,N_21777);
xnor U21972 (N_21972,N_21676,N_21473);
and U21973 (N_21973,N_21518,N_21399);
or U21974 (N_21974,N_21516,N_21293);
and U21975 (N_21975,N_21258,N_21642);
or U21976 (N_21976,N_21566,N_21484);
nand U21977 (N_21977,N_21454,N_21669);
nor U21978 (N_21978,N_21701,N_21511);
nand U21979 (N_21979,N_21373,N_21803);
and U21980 (N_21980,N_21277,N_21802);
nor U21981 (N_21981,N_21677,N_21591);
and U21982 (N_21982,N_21868,N_21590);
nor U21983 (N_21983,N_21825,N_21384);
nor U21984 (N_21984,N_21279,N_21778);
nand U21985 (N_21985,N_21797,N_21561);
xor U21986 (N_21986,N_21310,N_21534);
nand U21987 (N_21987,N_21447,N_21750);
and U21988 (N_21988,N_21538,N_21529);
xor U21989 (N_21989,N_21397,N_21537);
nand U21990 (N_21990,N_21658,N_21439);
nor U21991 (N_21991,N_21655,N_21582);
nand U21992 (N_21992,N_21698,N_21374);
nor U21993 (N_21993,N_21652,N_21398);
or U21994 (N_21994,N_21853,N_21863);
or U21995 (N_21995,N_21357,N_21376);
and U21996 (N_21996,N_21272,N_21570);
nand U21997 (N_21997,N_21809,N_21713);
nor U21998 (N_21998,N_21649,N_21436);
nor U21999 (N_21999,N_21297,N_21327);
and U22000 (N_22000,N_21510,N_21262);
or U22001 (N_22001,N_21848,N_21531);
and U22002 (N_22002,N_21568,N_21753);
or U22003 (N_22003,N_21338,N_21707);
nor U22004 (N_22004,N_21792,N_21586);
xnor U22005 (N_22005,N_21691,N_21294);
and U22006 (N_22006,N_21364,N_21255);
and U22007 (N_22007,N_21336,N_21761);
nor U22008 (N_22008,N_21594,N_21762);
or U22009 (N_22009,N_21304,N_21536);
nand U22010 (N_22010,N_21502,N_21261);
and U22011 (N_22011,N_21533,N_21517);
nor U22012 (N_22012,N_21501,N_21678);
or U22013 (N_22013,N_21266,N_21654);
or U22014 (N_22014,N_21837,N_21653);
nor U22015 (N_22015,N_21689,N_21526);
nor U22016 (N_22016,N_21828,N_21634);
and U22017 (N_22017,N_21340,N_21820);
or U22018 (N_22018,N_21460,N_21734);
or U22019 (N_22019,N_21854,N_21732);
and U22020 (N_22020,N_21806,N_21457);
nand U22021 (N_22021,N_21354,N_21351);
nor U22022 (N_22022,N_21550,N_21685);
and U22023 (N_22023,N_21283,N_21571);
xnor U22024 (N_22024,N_21864,N_21402);
nor U22025 (N_22025,N_21671,N_21865);
nor U22026 (N_22026,N_21598,N_21406);
and U22027 (N_22027,N_21396,N_21556);
nor U22028 (N_22028,N_21735,N_21450);
nor U22029 (N_22029,N_21709,N_21812);
and U22030 (N_22030,N_21487,N_21378);
nor U22031 (N_22031,N_21727,N_21821);
xor U22032 (N_22032,N_21699,N_21552);
and U22033 (N_22033,N_21469,N_21285);
xor U22034 (N_22034,N_21856,N_21546);
or U22035 (N_22035,N_21554,N_21747);
nand U22036 (N_22036,N_21668,N_21723);
xnor U22037 (N_22037,N_21461,N_21485);
and U22038 (N_22038,N_21415,N_21322);
and U22039 (N_22039,N_21610,N_21438);
nor U22040 (N_22040,N_21599,N_21254);
nor U22041 (N_22041,N_21251,N_21718);
or U22042 (N_22042,N_21558,N_21754);
and U22043 (N_22043,N_21867,N_21628);
or U22044 (N_22044,N_21451,N_21395);
nand U22045 (N_22045,N_21811,N_21318);
nor U22046 (N_22046,N_21661,N_21519);
xnor U22047 (N_22047,N_21860,N_21640);
nand U22048 (N_22048,N_21563,N_21468);
nor U22049 (N_22049,N_21488,N_21622);
nor U22050 (N_22050,N_21679,N_21490);
and U22051 (N_22051,N_21626,N_21363);
or U22052 (N_22052,N_21409,N_21602);
nand U22053 (N_22053,N_21663,N_21250);
nand U22054 (N_22054,N_21694,N_21419);
and U22055 (N_22055,N_21670,N_21711);
nand U22056 (N_22056,N_21791,N_21737);
nand U22057 (N_22057,N_21326,N_21472);
nand U22058 (N_22058,N_21445,N_21638);
or U22059 (N_22059,N_21389,N_21549);
and U22060 (N_22060,N_21859,N_21745);
nand U22061 (N_22061,N_21257,N_21629);
nor U22062 (N_22062,N_21393,N_21833);
nand U22063 (N_22063,N_21334,N_21861);
and U22064 (N_22064,N_21432,N_21332);
or U22065 (N_22065,N_21377,N_21404);
or U22066 (N_22066,N_21715,N_21641);
nand U22067 (N_22067,N_21623,N_21444);
and U22068 (N_22068,N_21330,N_21347);
nand U22069 (N_22069,N_21437,N_21259);
xnor U22070 (N_22070,N_21504,N_21687);
nand U22071 (N_22071,N_21295,N_21413);
and U22072 (N_22072,N_21822,N_21731);
nand U22073 (N_22073,N_21361,N_21606);
or U22074 (N_22074,N_21410,N_21576);
nor U22075 (N_22075,N_21603,N_21742);
xnor U22076 (N_22076,N_21286,N_21604);
or U22077 (N_22077,N_21841,N_21281);
and U22078 (N_22078,N_21370,N_21657);
nand U22079 (N_22079,N_21845,N_21588);
nor U22080 (N_22080,N_21309,N_21779);
or U22081 (N_22081,N_21424,N_21331);
and U22082 (N_22082,N_21320,N_21360);
nand U22083 (N_22083,N_21477,N_21273);
or U22084 (N_22084,N_21749,N_21507);
nand U22085 (N_22085,N_21740,N_21674);
or U22086 (N_22086,N_21407,N_21714);
and U22087 (N_22087,N_21728,N_21722);
and U22088 (N_22088,N_21514,N_21476);
and U22089 (N_22089,N_21418,N_21819);
nor U22090 (N_22090,N_21575,N_21721);
nor U22091 (N_22091,N_21434,N_21315);
and U22092 (N_22092,N_21493,N_21786);
or U22093 (N_22093,N_21381,N_21528);
and U22094 (N_22094,N_21449,N_21417);
and U22095 (N_22095,N_21435,N_21560);
or U22096 (N_22096,N_21341,N_21512);
nor U22097 (N_22097,N_21346,N_21637);
nand U22098 (N_22098,N_21597,N_21394);
nor U22099 (N_22099,N_21489,N_21433);
or U22100 (N_22100,N_21639,N_21768);
or U22101 (N_22101,N_21795,N_21835);
nand U22102 (N_22102,N_21343,N_21276);
xor U22103 (N_22103,N_21353,N_21431);
nor U22104 (N_22104,N_21390,N_21801);
nor U22105 (N_22105,N_21751,N_21371);
nor U22106 (N_22106,N_21543,N_21583);
nor U22107 (N_22107,N_21796,N_21308);
nor U22108 (N_22108,N_21624,N_21478);
xor U22109 (N_22109,N_21614,N_21282);
nand U22110 (N_22110,N_21305,N_21383);
nand U22111 (N_22111,N_21736,N_21672);
and U22112 (N_22112,N_21405,N_21817);
or U22113 (N_22113,N_21775,N_21843);
or U22114 (N_22114,N_21693,N_21467);
or U22115 (N_22115,N_21733,N_21776);
xnor U22116 (N_22116,N_21857,N_21785);
nand U22117 (N_22117,N_21643,N_21580);
and U22118 (N_22118,N_21300,N_21355);
and U22119 (N_22119,N_21738,N_21474);
nand U22120 (N_22120,N_21366,N_21660);
or U22121 (N_22121,N_21544,N_21772);
xor U22122 (N_22122,N_21356,N_21794);
or U22123 (N_22123,N_21684,N_21593);
xor U22124 (N_22124,N_21782,N_21631);
nand U22125 (N_22125,N_21408,N_21705);
nand U22126 (N_22126,N_21565,N_21268);
nand U22127 (N_22127,N_21805,N_21442);
nand U22128 (N_22128,N_21448,N_21535);
nand U22129 (N_22129,N_21391,N_21850);
xor U22130 (N_22130,N_21306,N_21783);
nor U22131 (N_22131,N_21301,N_21764);
and U22132 (N_22132,N_21479,N_21414);
or U22133 (N_22133,N_21789,N_21337);
xnor U22134 (N_22134,N_21292,N_21842);
nor U22135 (N_22135,N_21321,N_21385);
nor U22136 (N_22136,N_21441,N_21287);
or U22137 (N_22137,N_21808,N_21547);
or U22138 (N_22138,N_21253,N_21605);
xnor U22139 (N_22139,N_21495,N_21608);
or U22140 (N_22140,N_21342,N_21348);
and U22141 (N_22141,N_21617,N_21420);
or U22142 (N_22142,N_21527,N_21289);
and U22143 (N_22143,N_21375,N_21774);
or U22144 (N_22144,N_21807,N_21766);
or U22145 (N_22145,N_21311,N_21325);
nor U22146 (N_22146,N_21748,N_21625);
and U22147 (N_22147,N_21615,N_21664);
nand U22148 (N_22148,N_21769,N_21486);
nand U22149 (N_22149,N_21656,N_21847);
nand U22150 (N_22150,N_21823,N_21358);
nor U22151 (N_22151,N_21412,N_21844);
or U22152 (N_22152,N_21743,N_21314);
and U22153 (N_22153,N_21700,N_21256);
nand U22154 (N_22154,N_21834,N_21729);
nand U22155 (N_22155,N_21403,N_21613);
nor U22156 (N_22156,N_21744,N_21648);
nor U22157 (N_22157,N_21553,N_21271);
nand U22158 (N_22158,N_21675,N_21382);
nand U22159 (N_22159,N_21784,N_21739);
or U22160 (N_22160,N_21465,N_21270);
nand U22161 (N_22161,N_21813,N_21662);
nor U22162 (N_22162,N_21804,N_21400);
nand U22163 (N_22163,N_21673,N_21274);
and U22164 (N_22164,N_21793,N_21428);
nor U22165 (N_22165,N_21532,N_21503);
or U22166 (N_22166,N_21871,N_21746);
nor U22167 (N_22167,N_21716,N_21548);
nand U22168 (N_22168,N_21299,N_21607);
nor U22169 (N_22169,N_21757,N_21296);
nor U22170 (N_22170,N_21269,N_21494);
nor U22171 (N_22171,N_21429,N_21578);
nor U22172 (N_22172,N_21596,N_21359);
nor U22173 (N_22173,N_21681,N_21367);
nor U22174 (N_22174,N_21587,N_21482);
nor U22175 (N_22175,N_21647,N_21870);
and U22176 (N_22176,N_21323,N_21755);
nor U22177 (N_22177,N_21290,N_21752);
or U22178 (N_22178,N_21815,N_21851);
xnor U22179 (N_22179,N_21421,N_21379);
nand U22180 (N_22180,N_21298,N_21455);
and U22181 (N_22181,N_21633,N_21839);
and U22182 (N_22182,N_21498,N_21515);
or U22183 (N_22183,N_21459,N_21592);
or U22184 (N_22184,N_21464,N_21263);
xor U22185 (N_22185,N_21545,N_21706);
nor U22186 (N_22186,N_21386,N_21492);
or U22187 (N_22187,N_21440,N_21821);
nor U22188 (N_22188,N_21672,N_21598);
nor U22189 (N_22189,N_21871,N_21302);
nand U22190 (N_22190,N_21331,N_21372);
or U22191 (N_22191,N_21358,N_21774);
nand U22192 (N_22192,N_21411,N_21293);
or U22193 (N_22193,N_21455,N_21502);
and U22194 (N_22194,N_21318,N_21681);
nor U22195 (N_22195,N_21393,N_21267);
or U22196 (N_22196,N_21769,N_21270);
nor U22197 (N_22197,N_21468,N_21803);
nand U22198 (N_22198,N_21553,N_21545);
or U22199 (N_22199,N_21314,N_21569);
nand U22200 (N_22200,N_21379,N_21381);
and U22201 (N_22201,N_21456,N_21726);
nand U22202 (N_22202,N_21783,N_21361);
nand U22203 (N_22203,N_21346,N_21592);
or U22204 (N_22204,N_21389,N_21763);
nor U22205 (N_22205,N_21474,N_21687);
nand U22206 (N_22206,N_21701,N_21780);
or U22207 (N_22207,N_21390,N_21773);
nor U22208 (N_22208,N_21622,N_21601);
or U22209 (N_22209,N_21731,N_21539);
or U22210 (N_22210,N_21612,N_21706);
nand U22211 (N_22211,N_21573,N_21360);
nor U22212 (N_22212,N_21351,N_21512);
nand U22213 (N_22213,N_21579,N_21385);
nand U22214 (N_22214,N_21550,N_21347);
or U22215 (N_22215,N_21323,N_21612);
and U22216 (N_22216,N_21282,N_21724);
or U22217 (N_22217,N_21497,N_21321);
xnor U22218 (N_22218,N_21661,N_21803);
xnor U22219 (N_22219,N_21411,N_21354);
nand U22220 (N_22220,N_21294,N_21473);
and U22221 (N_22221,N_21405,N_21685);
or U22222 (N_22222,N_21744,N_21260);
or U22223 (N_22223,N_21724,N_21370);
xor U22224 (N_22224,N_21775,N_21688);
nor U22225 (N_22225,N_21446,N_21772);
or U22226 (N_22226,N_21510,N_21331);
or U22227 (N_22227,N_21661,N_21521);
nor U22228 (N_22228,N_21860,N_21826);
nor U22229 (N_22229,N_21702,N_21256);
or U22230 (N_22230,N_21416,N_21582);
nand U22231 (N_22231,N_21444,N_21626);
or U22232 (N_22232,N_21639,N_21369);
nand U22233 (N_22233,N_21653,N_21331);
or U22234 (N_22234,N_21451,N_21798);
or U22235 (N_22235,N_21708,N_21282);
and U22236 (N_22236,N_21380,N_21337);
or U22237 (N_22237,N_21813,N_21704);
or U22238 (N_22238,N_21649,N_21722);
and U22239 (N_22239,N_21287,N_21337);
nor U22240 (N_22240,N_21777,N_21855);
or U22241 (N_22241,N_21682,N_21592);
or U22242 (N_22242,N_21868,N_21694);
or U22243 (N_22243,N_21299,N_21760);
and U22244 (N_22244,N_21290,N_21351);
and U22245 (N_22245,N_21549,N_21295);
and U22246 (N_22246,N_21353,N_21350);
xnor U22247 (N_22247,N_21515,N_21526);
and U22248 (N_22248,N_21600,N_21683);
and U22249 (N_22249,N_21638,N_21593);
nor U22250 (N_22250,N_21638,N_21740);
and U22251 (N_22251,N_21826,N_21367);
nand U22252 (N_22252,N_21602,N_21826);
or U22253 (N_22253,N_21858,N_21866);
or U22254 (N_22254,N_21657,N_21866);
nand U22255 (N_22255,N_21453,N_21630);
xnor U22256 (N_22256,N_21830,N_21562);
xnor U22257 (N_22257,N_21625,N_21375);
or U22258 (N_22258,N_21421,N_21714);
nor U22259 (N_22259,N_21829,N_21871);
nand U22260 (N_22260,N_21372,N_21567);
or U22261 (N_22261,N_21258,N_21708);
or U22262 (N_22262,N_21365,N_21510);
nor U22263 (N_22263,N_21762,N_21698);
or U22264 (N_22264,N_21718,N_21707);
or U22265 (N_22265,N_21720,N_21323);
or U22266 (N_22266,N_21801,N_21523);
or U22267 (N_22267,N_21608,N_21705);
nor U22268 (N_22268,N_21472,N_21831);
or U22269 (N_22269,N_21531,N_21661);
and U22270 (N_22270,N_21699,N_21335);
nor U22271 (N_22271,N_21326,N_21782);
nand U22272 (N_22272,N_21290,N_21624);
and U22273 (N_22273,N_21414,N_21867);
xnor U22274 (N_22274,N_21473,N_21418);
nand U22275 (N_22275,N_21832,N_21838);
or U22276 (N_22276,N_21604,N_21792);
nand U22277 (N_22277,N_21791,N_21838);
and U22278 (N_22278,N_21598,N_21572);
or U22279 (N_22279,N_21556,N_21376);
nor U22280 (N_22280,N_21757,N_21324);
nand U22281 (N_22281,N_21653,N_21696);
nor U22282 (N_22282,N_21669,N_21336);
or U22283 (N_22283,N_21867,N_21644);
nor U22284 (N_22284,N_21834,N_21680);
nor U22285 (N_22285,N_21748,N_21461);
xnor U22286 (N_22286,N_21569,N_21605);
xnor U22287 (N_22287,N_21562,N_21255);
and U22288 (N_22288,N_21444,N_21515);
or U22289 (N_22289,N_21560,N_21273);
nor U22290 (N_22290,N_21753,N_21396);
and U22291 (N_22291,N_21750,N_21848);
nand U22292 (N_22292,N_21391,N_21468);
and U22293 (N_22293,N_21720,N_21500);
or U22294 (N_22294,N_21740,N_21258);
nand U22295 (N_22295,N_21680,N_21554);
nand U22296 (N_22296,N_21359,N_21712);
and U22297 (N_22297,N_21569,N_21692);
and U22298 (N_22298,N_21718,N_21649);
xor U22299 (N_22299,N_21504,N_21695);
nor U22300 (N_22300,N_21505,N_21853);
and U22301 (N_22301,N_21421,N_21375);
or U22302 (N_22302,N_21726,N_21347);
nand U22303 (N_22303,N_21594,N_21389);
nand U22304 (N_22304,N_21723,N_21793);
xor U22305 (N_22305,N_21360,N_21542);
or U22306 (N_22306,N_21609,N_21688);
xor U22307 (N_22307,N_21389,N_21305);
or U22308 (N_22308,N_21572,N_21725);
nand U22309 (N_22309,N_21273,N_21386);
nor U22310 (N_22310,N_21278,N_21508);
nand U22311 (N_22311,N_21592,N_21675);
nand U22312 (N_22312,N_21700,N_21781);
and U22313 (N_22313,N_21563,N_21270);
xor U22314 (N_22314,N_21700,N_21346);
xnor U22315 (N_22315,N_21319,N_21553);
or U22316 (N_22316,N_21848,N_21810);
nand U22317 (N_22317,N_21455,N_21702);
xnor U22318 (N_22318,N_21310,N_21386);
and U22319 (N_22319,N_21556,N_21387);
xor U22320 (N_22320,N_21323,N_21753);
or U22321 (N_22321,N_21768,N_21600);
nor U22322 (N_22322,N_21520,N_21528);
and U22323 (N_22323,N_21342,N_21471);
and U22324 (N_22324,N_21837,N_21706);
nand U22325 (N_22325,N_21480,N_21592);
xor U22326 (N_22326,N_21321,N_21778);
nor U22327 (N_22327,N_21612,N_21698);
nor U22328 (N_22328,N_21816,N_21843);
and U22329 (N_22329,N_21735,N_21262);
nor U22330 (N_22330,N_21865,N_21832);
nand U22331 (N_22331,N_21555,N_21473);
or U22332 (N_22332,N_21585,N_21694);
xnor U22333 (N_22333,N_21826,N_21765);
or U22334 (N_22334,N_21420,N_21320);
or U22335 (N_22335,N_21465,N_21322);
or U22336 (N_22336,N_21498,N_21377);
nor U22337 (N_22337,N_21828,N_21651);
nand U22338 (N_22338,N_21785,N_21789);
and U22339 (N_22339,N_21536,N_21454);
xor U22340 (N_22340,N_21807,N_21838);
or U22341 (N_22341,N_21502,N_21256);
and U22342 (N_22342,N_21633,N_21796);
nor U22343 (N_22343,N_21277,N_21554);
and U22344 (N_22344,N_21406,N_21350);
and U22345 (N_22345,N_21773,N_21274);
nor U22346 (N_22346,N_21395,N_21525);
nor U22347 (N_22347,N_21575,N_21463);
nor U22348 (N_22348,N_21542,N_21644);
nor U22349 (N_22349,N_21537,N_21605);
nor U22350 (N_22350,N_21530,N_21671);
nand U22351 (N_22351,N_21486,N_21319);
and U22352 (N_22352,N_21704,N_21310);
or U22353 (N_22353,N_21408,N_21356);
nor U22354 (N_22354,N_21756,N_21579);
nor U22355 (N_22355,N_21255,N_21684);
xor U22356 (N_22356,N_21809,N_21276);
nand U22357 (N_22357,N_21323,N_21696);
nand U22358 (N_22358,N_21790,N_21384);
and U22359 (N_22359,N_21433,N_21627);
and U22360 (N_22360,N_21602,N_21771);
nand U22361 (N_22361,N_21303,N_21324);
nand U22362 (N_22362,N_21283,N_21533);
and U22363 (N_22363,N_21706,N_21862);
xnor U22364 (N_22364,N_21848,N_21596);
nor U22365 (N_22365,N_21713,N_21382);
and U22366 (N_22366,N_21672,N_21544);
nor U22367 (N_22367,N_21401,N_21804);
nand U22368 (N_22368,N_21298,N_21369);
xor U22369 (N_22369,N_21544,N_21400);
nand U22370 (N_22370,N_21361,N_21767);
nor U22371 (N_22371,N_21277,N_21489);
nand U22372 (N_22372,N_21691,N_21335);
xor U22373 (N_22373,N_21271,N_21618);
nand U22374 (N_22374,N_21330,N_21305);
nor U22375 (N_22375,N_21450,N_21623);
or U22376 (N_22376,N_21507,N_21512);
nor U22377 (N_22377,N_21553,N_21694);
or U22378 (N_22378,N_21423,N_21538);
nand U22379 (N_22379,N_21384,N_21639);
xnor U22380 (N_22380,N_21311,N_21763);
xor U22381 (N_22381,N_21689,N_21278);
nand U22382 (N_22382,N_21724,N_21733);
and U22383 (N_22383,N_21564,N_21585);
or U22384 (N_22384,N_21480,N_21607);
and U22385 (N_22385,N_21720,N_21679);
nor U22386 (N_22386,N_21797,N_21474);
nor U22387 (N_22387,N_21805,N_21405);
or U22388 (N_22388,N_21616,N_21361);
nand U22389 (N_22389,N_21815,N_21487);
nor U22390 (N_22390,N_21478,N_21399);
xnor U22391 (N_22391,N_21536,N_21668);
xnor U22392 (N_22392,N_21671,N_21641);
nand U22393 (N_22393,N_21457,N_21322);
xor U22394 (N_22394,N_21424,N_21583);
and U22395 (N_22395,N_21358,N_21437);
or U22396 (N_22396,N_21585,N_21512);
xnor U22397 (N_22397,N_21833,N_21790);
and U22398 (N_22398,N_21340,N_21512);
xnor U22399 (N_22399,N_21454,N_21727);
and U22400 (N_22400,N_21754,N_21797);
or U22401 (N_22401,N_21648,N_21308);
nor U22402 (N_22402,N_21793,N_21337);
or U22403 (N_22403,N_21845,N_21710);
nor U22404 (N_22404,N_21588,N_21764);
xnor U22405 (N_22405,N_21792,N_21270);
nor U22406 (N_22406,N_21787,N_21584);
and U22407 (N_22407,N_21707,N_21658);
nor U22408 (N_22408,N_21495,N_21622);
nor U22409 (N_22409,N_21689,N_21575);
or U22410 (N_22410,N_21501,N_21418);
xor U22411 (N_22411,N_21327,N_21448);
or U22412 (N_22412,N_21837,N_21791);
and U22413 (N_22413,N_21543,N_21766);
or U22414 (N_22414,N_21644,N_21494);
nand U22415 (N_22415,N_21698,N_21370);
nor U22416 (N_22416,N_21637,N_21796);
and U22417 (N_22417,N_21624,N_21796);
nand U22418 (N_22418,N_21524,N_21761);
nand U22419 (N_22419,N_21829,N_21780);
nor U22420 (N_22420,N_21742,N_21442);
nor U22421 (N_22421,N_21538,N_21560);
and U22422 (N_22422,N_21750,N_21499);
and U22423 (N_22423,N_21857,N_21310);
and U22424 (N_22424,N_21465,N_21519);
or U22425 (N_22425,N_21749,N_21340);
or U22426 (N_22426,N_21848,N_21587);
nand U22427 (N_22427,N_21800,N_21664);
or U22428 (N_22428,N_21296,N_21859);
and U22429 (N_22429,N_21698,N_21833);
nor U22430 (N_22430,N_21668,N_21394);
or U22431 (N_22431,N_21627,N_21453);
nor U22432 (N_22432,N_21414,N_21571);
or U22433 (N_22433,N_21778,N_21413);
and U22434 (N_22434,N_21797,N_21277);
and U22435 (N_22435,N_21264,N_21395);
nand U22436 (N_22436,N_21569,N_21646);
or U22437 (N_22437,N_21527,N_21543);
or U22438 (N_22438,N_21739,N_21419);
nand U22439 (N_22439,N_21284,N_21859);
and U22440 (N_22440,N_21265,N_21789);
nor U22441 (N_22441,N_21827,N_21579);
or U22442 (N_22442,N_21284,N_21863);
nand U22443 (N_22443,N_21541,N_21379);
or U22444 (N_22444,N_21715,N_21304);
nor U22445 (N_22445,N_21603,N_21638);
and U22446 (N_22446,N_21706,N_21762);
and U22447 (N_22447,N_21534,N_21417);
and U22448 (N_22448,N_21844,N_21398);
nand U22449 (N_22449,N_21787,N_21260);
or U22450 (N_22450,N_21643,N_21575);
nor U22451 (N_22451,N_21850,N_21852);
nand U22452 (N_22452,N_21740,N_21499);
nor U22453 (N_22453,N_21759,N_21775);
and U22454 (N_22454,N_21401,N_21478);
nor U22455 (N_22455,N_21482,N_21565);
nand U22456 (N_22456,N_21390,N_21558);
nor U22457 (N_22457,N_21815,N_21826);
and U22458 (N_22458,N_21592,N_21406);
nor U22459 (N_22459,N_21746,N_21657);
nor U22460 (N_22460,N_21710,N_21515);
or U22461 (N_22461,N_21370,N_21525);
or U22462 (N_22462,N_21671,N_21604);
and U22463 (N_22463,N_21812,N_21579);
nor U22464 (N_22464,N_21310,N_21741);
nand U22465 (N_22465,N_21660,N_21414);
nor U22466 (N_22466,N_21711,N_21722);
or U22467 (N_22467,N_21491,N_21257);
nand U22468 (N_22468,N_21511,N_21420);
and U22469 (N_22469,N_21691,N_21581);
or U22470 (N_22470,N_21318,N_21532);
nand U22471 (N_22471,N_21645,N_21840);
and U22472 (N_22472,N_21260,N_21722);
nor U22473 (N_22473,N_21747,N_21264);
nor U22474 (N_22474,N_21284,N_21374);
and U22475 (N_22475,N_21797,N_21314);
and U22476 (N_22476,N_21757,N_21817);
nand U22477 (N_22477,N_21394,N_21686);
and U22478 (N_22478,N_21702,N_21264);
nor U22479 (N_22479,N_21649,N_21276);
or U22480 (N_22480,N_21780,N_21743);
and U22481 (N_22481,N_21631,N_21380);
nor U22482 (N_22482,N_21612,N_21581);
nand U22483 (N_22483,N_21564,N_21621);
nand U22484 (N_22484,N_21427,N_21807);
or U22485 (N_22485,N_21432,N_21631);
and U22486 (N_22486,N_21351,N_21253);
xnor U22487 (N_22487,N_21428,N_21264);
or U22488 (N_22488,N_21872,N_21383);
nand U22489 (N_22489,N_21784,N_21534);
and U22490 (N_22490,N_21544,N_21623);
nand U22491 (N_22491,N_21484,N_21652);
nand U22492 (N_22492,N_21836,N_21484);
nand U22493 (N_22493,N_21438,N_21708);
and U22494 (N_22494,N_21750,N_21599);
nand U22495 (N_22495,N_21329,N_21708);
or U22496 (N_22496,N_21330,N_21781);
nand U22497 (N_22497,N_21675,N_21713);
nor U22498 (N_22498,N_21605,N_21651);
nand U22499 (N_22499,N_21310,N_21512);
nor U22500 (N_22500,N_22071,N_21974);
and U22501 (N_22501,N_22161,N_21899);
or U22502 (N_22502,N_22331,N_22407);
xor U22503 (N_22503,N_21971,N_21889);
nand U22504 (N_22504,N_22116,N_22356);
or U22505 (N_22505,N_21962,N_22387);
nor U22506 (N_22506,N_21888,N_22283);
nor U22507 (N_22507,N_22250,N_22058);
nand U22508 (N_22508,N_22307,N_22281);
and U22509 (N_22509,N_22496,N_21891);
and U22510 (N_22510,N_21900,N_22017);
and U22511 (N_22511,N_21917,N_22171);
or U22512 (N_22512,N_22188,N_22470);
nor U22513 (N_22513,N_22094,N_22135);
and U22514 (N_22514,N_22463,N_21928);
nand U22515 (N_22515,N_21943,N_22298);
nand U22516 (N_22516,N_22284,N_22297);
or U22517 (N_22517,N_21919,N_22055);
xnor U22518 (N_22518,N_22193,N_22028);
nor U22519 (N_22519,N_22372,N_22380);
and U22520 (N_22520,N_22385,N_22275);
nand U22521 (N_22521,N_22333,N_22304);
xor U22522 (N_22522,N_22424,N_22123);
nor U22523 (N_22523,N_22020,N_22126);
xor U22524 (N_22524,N_22257,N_22241);
or U22525 (N_22525,N_22411,N_22070);
and U22526 (N_22526,N_22162,N_21975);
nand U22527 (N_22527,N_21969,N_22471);
or U22528 (N_22528,N_21979,N_22122);
or U22529 (N_22529,N_22446,N_22037);
nor U22530 (N_22530,N_22209,N_22415);
and U22531 (N_22531,N_21881,N_22190);
xor U22532 (N_22532,N_22497,N_21988);
nor U22533 (N_22533,N_21993,N_21960);
and U22534 (N_22534,N_21876,N_22339);
or U22535 (N_22535,N_22472,N_22486);
nand U22536 (N_22536,N_22233,N_22400);
and U22537 (N_22537,N_22069,N_22234);
nor U22538 (N_22538,N_22273,N_22264);
or U22539 (N_22539,N_22416,N_22431);
nand U22540 (N_22540,N_22433,N_22279);
nand U22541 (N_22541,N_22350,N_22453);
or U22542 (N_22542,N_22317,N_21910);
nand U22543 (N_22543,N_22063,N_22391);
nand U22544 (N_22544,N_22054,N_22398);
xnor U22545 (N_22545,N_22202,N_21905);
or U22546 (N_22546,N_22258,N_22127);
or U22547 (N_22547,N_22410,N_22167);
and U22548 (N_22548,N_22376,N_22456);
nor U22549 (N_22549,N_21977,N_21995);
and U22550 (N_22550,N_22201,N_22206);
nand U22551 (N_22551,N_22011,N_22319);
nand U22552 (N_22552,N_22445,N_21992);
nand U22553 (N_22553,N_22146,N_22378);
nand U22554 (N_22554,N_22321,N_22053);
and U22555 (N_22555,N_21902,N_21875);
and U22556 (N_22556,N_22080,N_22314);
nor U22557 (N_22557,N_21950,N_22352);
nor U22558 (N_22558,N_22389,N_22148);
nand U22559 (N_22559,N_22216,N_22493);
and U22560 (N_22560,N_22084,N_22213);
nor U22561 (N_22561,N_21967,N_21944);
or U22562 (N_22562,N_22406,N_22021);
nor U22563 (N_22563,N_22425,N_22499);
xor U22564 (N_22564,N_22031,N_22318);
nand U22565 (N_22565,N_22034,N_22403);
nand U22566 (N_22566,N_21980,N_21983);
or U22567 (N_22567,N_22417,N_21914);
and U22568 (N_22568,N_22220,N_22191);
or U22569 (N_22569,N_22165,N_22289);
or U22570 (N_22570,N_21999,N_22211);
nor U22571 (N_22571,N_21965,N_22105);
nor U22572 (N_22572,N_22237,N_22335);
nand U22573 (N_22573,N_21940,N_22256);
or U22574 (N_22574,N_22061,N_21963);
or U22575 (N_22575,N_22093,N_22262);
nor U22576 (N_22576,N_22434,N_21895);
xnor U22577 (N_22577,N_22461,N_22251);
nor U22578 (N_22578,N_22014,N_22296);
nand U22579 (N_22579,N_22033,N_22484);
nand U22580 (N_22580,N_21985,N_22179);
or U22581 (N_22581,N_22108,N_22128);
nor U22582 (N_22582,N_21938,N_22156);
or U22583 (N_22583,N_22255,N_22479);
or U22584 (N_22584,N_22157,N_22150);
xnor U22585 (N_22585,N_22344,N_21883);
nor U22586 (N_22586,N_22130,N_22343);
nand U22587 (N_22587,N_21916,N_22012);
or U22588 (N_22588,N_22426,N_21949);
and U22589 (N_22589,N_21987,N_22361);
and U22590 (N_22590,N_22199,N_22002);
or U22591 (N_22591,N_22207,N_21922);
and U22592 (N_22592,N_22480,N_21972);
nand U22593 (N_22593,N_22138,N_22267);
nor U22594 (N_22594,N_22409,N_22325);
or U22595 (N_22595,N_22090,N_22113);
nor U22596 (N_22596,N_22030,N_22334);
xnor U22597 (N_22597,N_22439,N_22098);
xnor U22598 (N_22598,N_22462,N_22384);
and U22599 (N_22599,N_22373,N_22215);
nand U22600 (N_22600,N_22290,N_22327);
nand U22601 (N_22601,N_22124,N_22354);
or U22602 (N_22602,N_22222,N_22112);
and U22603 (N_22603,N_22375,N_22442);
and U22604 (N_22604,N_22026,N_22200);
nand U22605 (N_22605,N_22007,N_22395);
or U22606 (N_22606,N_21935,N_21920);
and U22607 (N_22607,N_21904,N_22009);
nor U22608 (N_22608,N_22302,N_22239);
nand U22609 (N_22609,N_22035,N_21903);
nor U22610 (N_22610,N_22322,N_21966);
and U22611 (N_22611,N_22455,N_22265);
nor U22612 (N_22612,N_22274,N_21898);
nor U22613 (N_22613,N_22042,N_21939);
xnor U22614 (N_22614,N_22203,N_21887);
nand U22615 (N_22615,N_22485,N_22192);
nor U22616 (N_22616,N_22172,N_22248);
or U22617 (N_22617,N_22025,N_22107);
nor U22618 (N_22618,N_22114,N_22360);
or U22619 (N_22619,N_22176,N_21970);
or U22620 (N_22620,N_22086,N_22096);
nor U22621 (N_22621,N_22082,N_22346);
and U22622 (N_22622,N_22219,N_22492);
nor U22623 (N_22623,N_22303,N_22300);
or U22624 (N_22624,N_22121,N_22115);
or U22625 (N_22625,N_22271,N_22057);
nand U22626 (N_22626,N_22197,N_22357);
and U22627 (N_22627,N_22364,N_22097);
nand U22628 (N_22628,N_22422,N_22323);
nor U22629 (N_22629,N_22109,N_22168);
nand U22630 (N_22630,N_21986,N_22224);
xor U22631 (N_22631,N_22247,N_22029);
or U22632 (N_22632,N_22338,N_21880);
and U22633 (N_22633,N_22137,N_22189);
nand U22634 (N_22634,N_22280,N_22382);
and U22635 (N_22635,N_22078,N_22062);
nand U22636 (N_22636,N_22003,N_21981);
and U22637 (N_22637,N_22181,N_21933);
nand U22638 (N_22638,N_22088,N_21953);
and U22639 (N_22639,N_22367,N_21877);
nor U22640 (N_22640,N_22074,N_21958);
nor U22641 (N_22641,N_22301,N_22469);
or U22642 (N_22642,N_22381,N_21982);
or U22643 (N_22643,N_22246,N_21911);
xnor U22644 (N_22644,N_22464,N_21990);
nor U22645 (N_22645,N_22091,N_21954);
nand U22646 (N_22646,N_22066,N_22312);
nor U22647 (N_22647,N_22473,N_21913);
xor U22648 (N_22648,N_22475,N_22056);
or U22649 (N_22649,N_22141,N_22177);
xnor U22650 (N_22650,N_22299,N_22068);
and U22651 (N_22651,N_22491,N_22019);
nor U22652 (N_22652,N_22404,N_22428);
or U22653 (N_22653,N_21946,N_22359);
xor U22654 (N_22654,N_22419,N_22489);
xnor U22655 (N_22655,N_22379,N_22187);
and U22656 (N_22656,N_21937,N_22240);
and U22657 (N_22657,N_22328,N_22119);
nand U22658 (N_22658,N_21994,N_22261);
xnor U22659 (N_22659,N_22362,N_22111);
and U22660 (N_22660,N_22402,N_21955);
and U22661 (N_22661,N_22164,N_22392);
nand U22662 (N_22662,N_22468,N_22345);
nand U22663 (N_22663,N_21976,N_22390);
or U22664 (N_22664,N_22447,N_21908);
nand U22665 (N_22665,N_21930,N_22120);
nand U22666 (N_22666,N_22236,N_22494);
or U22667 (N_22667,N_22399,N_22221);
and U22668 (N_22668,N_22254,N_22488);
nand U22669 (N_22669,N_22170,N_22351);
or U22670 (N_22670,N_22089,N_22110);
or U22671 (N_22671,N_21984,N_22401);
or U22672 (N_22672,N_22151,N_21893);
nor U22673 (N_22673,N_21956,N_21957);
or U22674 (N_22674,N_21978,N_22073);
and U22675 (N_22675,N_22450,N_22481);
or U22676 (N_22676,N_22045,N_22336);
nand U22677 (N_22677,N_21924,N_22460);
and U22678 (N_22678,N_22394,N_22173);
and U22679 (N_22679,N_22160,N_21948);
and U22680 (N_22680,N_22133,N_22324);
xnor U22681 (N_22681,N_22064,N_22243);
nor U22682 (N_22682,N_22018,N_22340);
and U22683 (N_22683,N_22075,N_22405);
and U22684 (N_22684,N_22022,N_22212);
and U22685 (N_22685,N_22449,N_21932);
nand U22686 (N_22686,N_22429,N_22016);
nand U22687 (N_22687,N_22326,N_22388);
nor U22688 (N_22688,N_22269,N_22152);
or U22689 (N_22689,N_22142,N_22059);
nor U22690 (N_22690,N_22316,N_22228);
nor U22691 (N_22691,N_22015,N_22467);
nand U22692 (N_22692,N_22125,N_21952);
nor U22693 (N_22693,N_22498,N_22013);
and U22694 (N_22694,N_22085,N_22214);
nor U22695 (N_22695,N_22039,N_22046);
or U22696 (N_22696,N_21942,N_22052);
nor U22697 (N_22697,N_22077,N_22330);
nand U22698 (N_22698,N_22286,N_22474);
nand U22699 (N_22699,N_21897,N_22076);
or U22700 (N_22700,N_22348,N_22329);
nor U22701 (N_22701,N_22000,N_22358);
nand U22702 (N_22702,N_22332,N_22414);
or U22703 (N_22703,N_22159,N_22366);
or U22704 (N_22704,N_22368,N_22272);
or U22705 (N_22705,N_22288,N_22095);
and U22706 (N_22706,N_21931,N_22166);
nor U22707 (N_22707,N_22249,N_22418);
or U22708 (N_22708,N_22079,N_21885);
and U22709 (N_22709,N_22072,N_21892);
or U22710 (N_22710,N_22435,N_22309);
xor U22711 (N_22711,N_22306,N_22099);
or U22712 (N_22712,N_22010,N_22310);
nor U22713 (N_22713,N_22315,N_22490);
nor U22714 (N_22714,N_22397,N_22038);
nand U22715 (N_22715,N_22454,N_22184);
nor U22716 (N_22716,N_22140,N_21927);
and U22717 (N_22717,N_22001,N_22432);
or U22718 (N_22718,N_22466,N_22421);
and U22719 (N_22719,N_22266,N_22452);
and U22720 (N_22720,N_22194,N_22185);
or U22721 (N_22721,N_22436,N_22223);
and U22722 (N_22722,N_21936,N_22291);
and U22723 (N_22723,N_21959,N_22006);
or U22724 (N_22724,N_21934,N_21890);
nand U22725 (N_22725,N_21918,N_21964);
and U22726 (N_22726,N_21921,N_22129);
or U22727 (N_22727,N_22065,N_22292);
or U22728 (N_22728,N_22036,N_22374);
nand U22729 (N_22729,N_22476,N_22451);
nand U22730 (N_22730,N_22103,N_21973);
nor U22731 (N_22731,N_22448,N_22051);
nor U22732 (N_22732,N_22440,N_22347);
nand U22733 (N_22733,N_22365,N_22174);
xor U22734 (N_22734,N_22369,N_22465);
nand U22735 (N_22735,N_21884,N_22023);
nand U22736 (N_22736,N_22139,N_21989);
nand U22737 (N_22737,N_22218,N_22259);
xnor U22738 (N_22738,N_22060,N_22204);
or U22739 (N_22739,N_22270,N_22242);
and U22740 (N_22740,N_22305,N_22155);
nand U22741 (N_22741,N_22229,N_22134);
nor U22742 (N_22742,N_22295,N_21907);
nor U22743 (N_22743,N_21878,N_22044);
nor U22744 (N_22744,N_22081,N_22438);
and U22745 (N_22745,N_22226,N_22196);
nand U22746 (N_22746,N_21991,N_22118);
nor U22747 (N_22747,N_22198,N_22131);
xor U22748 (N_22748,N_22370,N_22377);
or U22749 (N_22749,N_22050,N_22144);
nor U22750 (N_22750,N_22032,N_21901);
nor U22751 (N_22751,N_22430,N_21906);
and U22752 (N_22752,N_22393,N_22363);
and U22753 (N_22753,N_22482,N_22231);
nand U22754 (N_22754,N_22477,N_22483);
nand U22755 (N_22755,N_22282,N_22276);
and U22756 (N_22756,N_22353,N_21923);
xor U22757 (N_22757,N_22100,N_22024);
and U22758 (N_22758,N_22412,N_22106);
nand U22759 (N_22759,N_22238,N_22041);
nand U22760 (N_22760,N_22427,N_22175);
xnor U22761 (N_22761,N_22320,N_22153);
and U22762 (N_22762,N_22067,N_22230);
and U22763 (N_22763,N_21925,N_21879);
and U22764 (N_22764,N_22263,N_22355);
nand U22765 (N_22765,N_22313,N_22423);
nand U22766 (N_22766,N_22386,N_22208);
and U22767 (N_22767,N_22217,N_22040);
nor U22768 (N_22768,N_22420,N_21961);
nor U22769 (N_22769,N_22158,N_22154);
xor U22770 (N_22770,N_22186,N_22285);
nand U22771 (N_22771,N_22102,N_22205);
nor U22772 (N_22772,N_21886,N_22235);
xor U22773 (N_22773,N_22260,N_22311);
nand U22774 (N_22774,N_22101,N_22008);
nor U22775 (N_22775,N_22252,N_22443);
xnor U22776 (N_22776,N_21909,N_22225);
nor U22777 (N_22777,N_21912,N_21926);
or U22778 (N_22778,N_21998,N_21947);
xor U22779 (N_22779,N_21929,N_22293);
and U22780 (N_22780,N_22047,N_22143);
or U22781 (N_22781,N_21997,N_22244);
nor U22782 (N_22782,N_22227,N_22396);
nand U22783 (N_22783,N_22278,N_22049);
nor U22784 (N_22784,N_21882,N_22341);
nand U22785 (N_22785,N_22444,N_22337);
nand U22786 (N_22786,N_22210,N_22232);
and U22787 (N_22787,N_22005,N_21996);
nand U22788 (N_22788,N_22027,N_22132);
or U22789 (N_22789,N_21894,N_22043);
nor U22790 (N_22790,N_21951,N_22163);
nand U22791 (N_22791,N_22268,N_22253);
nand U22792 (N_22792,N_22083,N_21945);
nand U22793 (N_22793,N_22048,N_22408);
and U22794 (N_22794,N_22183,N_22087);
nor U22795 (N_22795,N_22308,N_22169);
and U22796 (N_22796,N_22487,N_22277);
nand U22797 (N_22797,N_22457,N_22478);
or U22798 (N_22798,N_22136,N_22178);
nand U22799 (N_22799,N_22349,N_21915);
xnor U22800 (N_22800,N_22180,N_22458);
nor U22801 (N_22801,N_22245,N_22413);
nand U22802 (N_22802,N_22004,N_22495);
xnor U22803 (N_22803,N_22147,N_22383);
or U22804 (N_22804,N_21968,N_22117);
and U22805 (N_22805,N_22371,N_21941);
nor U22806 (N_22806,N_22459,N_22182);
nand U22807 (N_22807,N_22342,N_22441);
or U22808 (N_22808,N_22287,N_21896);
nor U22809 (N_22809,N_22195,N_22104);
or U22810 (N_22810,N_22092,N_22437);
nand U22811 (N_22811,N_22149,N_22294);
and U22812 (N_22812,N_22145,N_22226);
nand U22813 (N_22813,N_22477,N_22031);
xnor U22814 (N_22814,N_22315,N_22399);
and U22815 (N_22815,N_22167,N_22030);
nor U22816 (N_22816,N_22015,N_22165);
nor U22817 (N_22817,N_22383,N_21985);
or U22818 (N_22818,N_22258,N_22232);
nor U22819 (N_22819,N_21946,N_22351);
and U22820 (N_22820,N_22404,N_22499);
nand U22821 (N_22821,N_22180,N_22296);
nor U22822 (N_22822,N_22069,N_22276);
and U22823 (N_22823,N_22481,N_22215);
nor U22824 (N_22824,N_22227,N_21997);
or U22825 (N_22825,N_22278,N_22144);
xor U22826 (N_22826,N_22421,N_21900);
and U22827 (N_22827,N_22192,N_22408);
and U22828 (N_22828,N_22337,N_22197);
or U22829 (N_22829,N_21997,N_22124);
xnor U22830 (N_22830,N_21875,N_22017);
or U22831 (N_22831,N_22117,N_22419);
and U22832 (N_22832,N_21923,N_21918);
or U22833 (N_22833,N_22043,N_22498);
nand U22834 (N_22834,N_22298,N_22480);
nand U22835 (N_22835,N_22365,N_22380);
and U22836 (N_22836,N_22137,N_22492);
and U22837 (N_22837,N_22033,N_21902);
xor U22838 (N_22838,N_22148,N_22275);
or U22839 (N_22839,N_22209,N_21915);
and U22840 (N_22840,N_22344,N_22247);
nor U22841 (N_22841,N_22375,N_21975);
nand U22842 (N_22842,N_22383,N_22394);
or U22843 (N_22843,N_22396,N_22289);
or U22844 (N_22844,N_22492,N_22406);
nand U22845 (N_22845,N_22298,N_22471);
and U22846 (N_22846,N_22254,N_22142);
or U22847 (N_22847,N_22479,N_21946);
nand U22848 (N_22848,N_21961,N_22023);
and U22849 (N_22849,N_21891,N_21969);
and U22850 (N_22850,N_22114,N_22202);
and U22851 (N_22851,N_22418,N_22239);
and U22852 (N_22852,N_22102,N_21927);
nor U22853 (N_22853,N_22351,N_22044);
nor U22854 (N_22854,N_22427,N_22042);
nor U22855 (N_22855,N_21992,N_22181);
nand U22856 (N_22856,N_22261,N_22437);
and U22857 (N_22857,N_22459,N_22170);
or U22858 (N_22858,N_21924,N_22369);
and U22859 (N_22859,N_22418,N_22166);
nand U22860 (N_22860,N_22324,N_22033);
or U22861 (N_22861,N_21930,N_21947);
or U22862 (N_22862,N_22418,N_21948);
and U22863 (N_22863,N_22348,N_22133);
nand U22864 (N_22864,N_22090,N_22455);
or U22865 (N_22865,N_22267,N_22486);
nand U22866 (N_22866,N_21924,N_22251);
and U22867 (N_22867,N_22486,N_22390);
and U22868 (N_22868,N_22213,N_21979);
nand U22869 (N_22869,N_22065,N_22151);
or U22870 (N_22870,N_22291,N_22324);
or U22871 (N_22871,N_22230,N_22471);
nor U22872 (N_22872,N_22440,N_22096);
or U22873 (N_22873,N_22318,N_21993);
nand U22874 (N_22874,N_22445,N_22357);
nand U22875 (N_22875,N_22380,N_22150);
nor U22876 (N_22876,N_22120,N_22377);
nand U22877 (N_22877,N_21963,N_21923);
or U22878 (N_22878,N_22446,N_22334);
nand U22879 (N_22879,N_21969,N_22195);
xnor U22880 (N_22880,N_22191,N_22200);
nand U22881 (N_22881,N_21884,N_22084);
and U22882 (N_22882,N_22002,N_22470);
and U22883 (N_22883,N_22224,N_21950);
or U22884 (N_22884,N_22457,N_22274);
or U22885 (N_22885,N_21980,N_22375);
nor U22886 (N_22886,N_21894,N_22437);
nor U22887 (N_22887,N_22206,N_22280);
or U22888 (N_22888,N_22304,N_22158);
nor U22889 (N_22889,N_22204,N_21899);
and U22890 (N_22890,N_22127,N_22038);
or U22891 (N_22891,N_22388,N_22378);
xor U22892 (N_22892,N_22380,N_22387);
nor U22893 (N_22893,N_22017,N_21985);
and U22894 (N_22894,N_22358,N_22108);
or U22895 (N_22895,N_22364,N_22379);
nand U22896 (N_22896,N_22480,N_22347);
nand U22897 (N_22897,N_22450,N_22056);
nand U22898 (N_22898,N_22366,N_22022);
xnor U22899 (N_22899,N_22062,N_22167);
or U22900 (N_22900,N_22477,N_22030);
nand U22901 (N_22901,N_22259,N_22072);
nor U22902 (N_22902,N_22202,N_21889);
and U22903 (N_22903,N_21931,N_22282);
and U22904 (N_22904,N_21923,N_22233);
or U22905 (N_22905,N_22002,N_21920);
nor U22906 (N_22906,N_21941,N_22321);
nor U22907 (N_22907,N_22262,N_22492);
and U22908 (N_22908,N_21960,N_22240);
or U22909 (N_22909,N_22108,N_22028);
nor U22910 (N_22910,N_22461,N_21889);
and U22911 (N_22911,N_21954,N_22177);
or U22912 (N_22912,N_21898,N_22276);
or U22913 (N_22913,N_22271,N_21994);
nor U22914 (N_22914,N_22100,N_21886);
nor U22915 (N_22915,N_22235,N_21899);
nor U22916 (N_22916,N_22020,N_21980);
nor U22917 (N_22917,N_22305,N_22040);
nor U22918 (N_22918,N_22261,N_21901);
xnor U22919 (N_22919,N_22109,N_21932);
nor U22920 (N_22920,N_21976,N_22031);
nor U22921 (N_22921,N_22059,N_21940);
xor U22922 (N_22922,N_22477,N_22434);
nand U22923 (N_22923,N_22443,N_22195);
and U22924 (N_22924,N_22112,N_22239);
and U22925 (N_22925,N_22428,N_22431);
and U22926 (N_22926,N_22161,N_22358);
and U22927 (N_22927,N_22021,N_22171);
and U22928 (N_22928,N_22317,N_21885);
nor U22929 (N_22929,N_22438,N_22341);
nor U22930 (N_22930,N_22468,N_22363);
or U22931 (N_22931,N_22117,N_22231);
xnor U22932 (N_22932,N_22357,N_22461);
nor U22933 (N_22933,N_22411,N_21889);
nand U22934 (N_22934,N_22018,N_22386);
or U22935 (N_22935,N_22169,N_22126);
and U22936 (N_22936,N_22148,N_22471);
or U22937 (N_22937,N_22447,N_21918);
nand U22938 (N_22938,N_22253,N_22363);
nor U22939 (N_22939,N_22327,N_22361);
and U22940 (N_22940,N_22323,N_22281);
or U22941 (N_22941,N_22198,N_21904);
xnor U22942 (N_22942,N_22376,N_22323);
nand U22943 (N_22943,N_22488,N_21943);
nor U22944 (N_22944,N_21950,N_22312);
nand U22945 (N_22945,N_22010,N_22489);
and U22946 (N_22946,N_22328,N_21970);
nor U22947 (N_22947,N_22041,N_22018);
and U22948 (N_22948,N_21976,N_22353);
and U22949 (N_22949,N_21972,N_22417);
and U22950 (N_22950,N_22372,N_22195);
nor U22951 (N_22951,N_22078,N_22364);
and U22952 (N_22952,N_22425,N_22412);
nor U22953 (N_22953,N_21895,N_22281);
and U22954 (N_22954,N_22460,N_22477);
or U22955 (N_22955,N_21932,N_22246);
nor U22956 (N_22956,N_22122,N_21896);
nand U22957 (N_22957,N_22436,N_22407);
nand U22958 (N_22958,N_22130,N_21882);
nand U22959 (N_22959,N_22097,N_22162);
and U22960 (N_22960,N_22159,N_22199);
or U22961 (N_22961,N_22161,N_22313);
nor U22962 (N_22962,N_22356,N_22494);
nor U22963 (N_22963,N_21951,N_21879);
or U22964 (N_22964,N_22203,N_22369);
and U22965 (N_22965,N_22133,N_22156);
or U22966 (N_22966,N_22260,N_22347);
nand U22967 (N_22967,N_22146,N_22118);
and U22968 (N_22968,N_22049,N_21977);
and U22969 (N_22969,N_22375,N_22395);
nor U22970 (N_22970,N_22027,N_22407);
nand U22971 (N_22971,N_22055,N_22347);
and U22972 (N_22972,N_21980,N_22085);
nand U22973 (N_22973,N_22432,N_22039);
and U22974 (N_22974,N_22171,N_22229);
nand U22975 (N_22975,N_21980,N_22078);
or U22976 (N_22976,N_22391,N_22291);
nand U22977 (N_22977,N_22420,N_22253);
nor U22978 (N_22978,N_22428,N_22154);
and U22979 (N_22979,N_22221,N_22178);
xnor U22980 (N_22980,N_22204,N_21959);
nand U22981 (N_22981,N_22441,N_22462);
or U22982 (N_22982,N_21916,N_21996);
or U22983 (N_22983,N_22434,N_22341);
or U22984 (N_22984,N_21915,N_22415);
or U22985 (N_22985,N_21909,N_22365);
and U22986 (N_22986,N_22393,N_22486);
nand U22987 (N_22987,N_22183,N_22069);
or U22988 (N_22988,N_22089,N_22215);
nor U22989 (N_22989,N_22083,N_21878);
nor U22990 (N_22990,N_22277,N_21998);
and U22991 (N_22991,N_22499,N_22232);
nor U22992 (N_22992,N_21940,N_22110);
nor U22993 (N_22993,N_21920,N_21911);
or U22994 (N_22994,N_22012,N_21978);
or U22995 (N_22995,N_21999,N_22428);
or U22996 (N_22996,N_22472,N_21883);
or U22997 (N_22997,N_22182,N_22037);
nand U22998 (N_22998,N_22212,N_22075);
nand U22999 (N_22999,N_22175,N_22461);
or U23000 (N_23000,N_22137,N_21969);
and U23001 (N_23001,N_21898,N_22066);
nand U23002 (N_23002,N_22101,N_22231);
nor U23003 (N_23003,N_21978,N_22479);
nand U23004 (N_23004,N_21887,N_22225);
nand U23005 (N_23005,N_21893,N_21970);
nor U23006 (N_23006,N_21934,N_21991);
or U23007 (N_23007,N_22320,N_22303);
and U23008 (N_23008,N_22375,N_22061);
and U23009 (N_23009,N_21975,N_22457);
xor U23010 (N_23010,N_22377,N_22100);
nor U23011 (N_23011,N_22306,N_21928);
and U23012 (N_23012,N_22087,N_22313);
nand U23013 (N_23013,N_21983,N_22076);
nor U23014 (N_23014,N_22495,N_22222);
or U23015 (N_23015,N_21993,N_22415);
nor U23016 (N_23016,N_22491,N_22280);
nand U23017 (N_23017,N_21893,N_21922);
or U23018 (N_23018,N_22455,N_22247);
nor U23019 (N_23019,N_22090,N_21956);
nor U23020 (N_23020,N_21918,N_22499);
and U23021 (N_23021,N_22170,N_22492);
nor U23022 (N_23022,N_22416,N_22352);
or U23023 (N_23023,N_22279,N_22262);
or U23024 (N_23024,N_22160,N_22318);
xnor U23025 (N_23025,N_22448,N_22254);
or U23026 (N_23026,N_22025,N_22319);
nor U23027 (N_23027,N_21875,N_22298);
xnor U23028 (N_23028,N_22062,N_22137);
nand U23029 (N_23029,N_22079,N_22376);
nand U23030 (N_23030,N_22356,N_21910);
nand U23031 (N_23031,N_22123,N_21920);
and U23032 (N_23032,N_22007,N_21930);
nor U23033 (N_23033,N_22479,N_22043);
or U23034 (N_23034,N_21883,N_21941);
nand U23035 (N_23035,N_22033,N_22354);
nor U23036 (N_23036,N_22050,N_22070);
nand U23037 (N_23037,N_21912,N_22447);
and U23038 (N_23038,N_22398,N_22396);
nand U23039 (N_23039,N_22141,N_22442);
or U23040 (N_23040,N_22292,N_21902);
and U23041 (N_23041,N_21915,N_22275);
nor U23042 (N_23042,N_22345,N_22288);
or U23043 (N_23043,N_22131,N_22070);
nand U23044 (N_23044,N_22276,N_22075);
nand U23045 (N_23045,N_22148,N_21896);
and U23046 (N_23046,N_22343,N_22009);
nand U23047 (N_23047,N_22089,N_22475);
nor U23048 (N_23048,N_21939,N_22214);
or U23049 (N_23049,N_22484,N_22377);
nand U23050 (N_23050,N_22052,N_22152);
nand U23051 (N_23051,N_22066,N_22159);
and U23052 (N_23052,N_22380,N_21940);
xnor U23053 (N_23053,N_22150,N_21939);
nand U23054 (N_23054,N_22233,N_22162);
nor U23055 (N_23055,N_22449,N_22216);
nand U23056 (N_23056,N_22383,N_22378);
nor U23057 (N_23057,N_22420,N_22122);
nor U23058 (N_23058,N_22429,N_22195);
xnor U23059 (N_23059,N_22222,N_21916);
or U23060 (N_23060,N_21994,N_22299);
or U23061 (N_23061,N_22226,N_21989);
and U23062 (N_23062,N_22009,N_22099);
nand U23063 (N_23063,N_22046,N_22286);
nand U23064 (N_23064,N_22146,N_22298);
nand U23065 (N_23065,N_22168,N_22294);
and U23066 (N_23066,N_22307,N_22366);
nor U23067 (N_23067,N_22225,N_22230);
or U23068 (N_23068,N_22413,N_22058);
nor U23069 (N_23069,N_22213,N_22090);
and U23070 (N_23070,N_22048,N_21891);
or U23071 (N_23071,N_22463,N_22151);
and U23072 (N_23072,N_22039,N_21915);
nor U23073 (N_23073,N_22300,N_22290);
nand U23074 (N_23074,N_22197,N_21890);
xnor U23075 (N_23075,N_22399,N_22349);
nand U23076 (N_23076,N_22455,N_22336);
nand U23077 (N_23077,N_21978,N_22407);
nand U23078 (N_23078,N_22485,N_22034);
xor U23079 (N_23079,N_22477,N_22256);
nor U23080 (N_23080,N_22263,N_22334);
and U23081 (N_23081,N_21948,N_22026);
or U23082 (N_23082,N_22387,N_22323);
xnor U23083 (N_23083,N_22439,N_21939);
or U23084 (N_23084,N_22472,N_22102);
xnor U23085 (N_23085,N_22195,N_21977);
xnor U23086 (N_23086,N_22268,N_22066);
nand U23087 (N_23087,N_22372,N_22279);
nand U23088 (N_23088,N_22158,N_22404);
xnor U23089 (N_23089,N_22015,N_21990);
or U23090 (N_23090,N_22090,N_22182);
and U23091 (N_23091,N_21989,N_22444);
nand U23092 (N_23092,N_22003,N_22399);
nor U23093 (N_23093,N_22272,N_21991);
or U23094 (N_23094,N_22167,N_22141);
and U23095 (N_23095,N_22019,N_21991);
and U23096 (N_23096,N_22383,N_22421);
nand U23097 (N_23097,N_21924,N_22141);
nand U23098 (N_23098,N_22457,N_21898);
nand U23099 (N_23099,N_22346,N_22046);
nand U23100 (N_23100,N_22001,N_22163);
nor U23101 (N_23101,N_22221,N_22189);
nor U23102 (N_23102,N_22073,N_22259);
nand U23103 (N_23103,N_22272,N_21888);
nor U23104 (N_23104,N_21963,N_22033);
nand U23105 (N_23105,N_22295,N_21950);
or U23106 (N_23106,N_21996,N_22299);
or U23107 (N_23107,N_22058,N_22161);
nor U23108 (N_23108,N_21936,N_22094);
nor U23109 (N_23109,N_22046,N_22309);
xor U23110 (N_23110,N_22311,N_22297);
nor U23111 (N_23111,N_22385,N_22320);
and U23112 (N_23112,N_22446,N_22437);
nand U23113 (N_23113,N_22490,N_22263);
nor U23114 (N_23114,N_22324,N_22000);
nand U23115 (N_23115,N_22497,N_22178);
and U23116 (N_23116,N_22163,N_21918);
nand U23117 (N_23117,N_22355,N_21918);
or U23118 (N_23118,N_22355,N_22155);
or U23119 (N_23119,N_22324,N_22319);
and U23120 (N_23120,N_22133,N_21922);
and U23121 (N_23121,N_22480,N_22030);
nand U23122 (N_23122,N_22354,N_22318);
or U23123 (N_23123,N_22236,N_21942);
or U23124 (N_23124,N_22078,N_21987);
nor U23125 (N_23125,N_22999,N_23053);
and U23126 (N_23126,N_22534,N_23027);
nand U23127 (N_23127,N_22882,N_22877);
xnor U23128 (N_23128,N_22626,N_22685);
nor U23129 (N_23129,N_23059,N_22529);
xnor U23130 (N_23130,N_22824,N_22989);
nand U23131 (N_23131,N_22931,N_23012);
xnor U23132 (N_23132,N_22893,N_22725);
or U23133 (N_23133,N_22610,N_23111);
and U23134 (N_23134,N_22602,N_22535);
or U23135 (N_23135,N_22703,N_22672);
nand U23136 (N_23136,N_22954,N_22810);
or U23137 (N_23137,N_22904,N_22953);
and U23138 (N_23138,N_22781,N_22899);
nor U23139 (N_23139,N_22597,N_22874);
nor U23140 (N_23140,N_22812,N_22895);
xor U23141 (N_23141,N_23023,N_22774);
nor U23142 (N_23142,N_22546,N_22927);
nand U23143 (N_23143,N_22928,N_22753);
and U23144 (N_23144,N_23078,N_23104);
and U23145 (N_23145,N_22545,N_23112);
or U23146 (N_23146,N_22518,N_23101);
xnor U23147 (N_23147,N_23081,N_23113);
and U23148 (N_23148,N_22601,N_22512);
nand U23149 (N_23149,N_22817,N_22581);
and U23150 (N_23150,N_23123,N_23061);
or U23151 (N_23151,N_22773,N_22830);
and U23152 (N_23152,N_22802,N_22868);
and U23153 (N_23153,N_23007,N_22573);
nor U23154 (N_23154,N_22662,N_22629);
and U23155 (N_23155,N_23000,N_22917);
and U23156 (N_23156,N_22972,N_22798);
nor U23157 (N_23157,N_22743,N_22655);
nor U23158 (N_23158,N_22656,N_22825);
or U23159 (N_23159,N_23041,N_22912);
nor U23160 (N_23160,N_22619,N_22814);
and U23161 (N_23161,N_22716,N_23122);
xnor U23162 (N_23162,N_22659,N_22704);
and U23163 (N_23163,N_23074,N_22555);
or U23164 (N_23164,N_22959,N_22682);
and U23165 (N_23165,N_23062,N_22724);
nand U23166 (N_23166,N_22971,N_22762);
and U23167 (N_23167,N_22625,N_22617);
nor U23168 (N_23168,N_22640,N_22652);
nand U23169 (N_23169,N_22985,N_22551);
or U23170 (N_23170,N_22562,N_23048);
nor U23171 (N_23171,N_22938,N_22970);
and U23172 (N_23172,N_22805,N_23108);
and U23173 (N_23173,N_22708,N_22542);
xnor U23174 (N_23174,N_23109,N_22891);
nand U23175 (N_23175,N_22641,N_22896);
or U23176 (N_23176,N_23090,N_22850);
or U23177 (N_23177,N_22963,N_22821);
or U23178 (N_23178,N_22568,N_22583);
xnor U23179 (N_23179,N_22744,N_22711);
nor U23180 (N_23180,N_22500,N_22785);
and U23181 (N_23181,N_22582,N_22738);
or U23182 (N_23182,N_22979,N_22691);
nand U23183 (N_23183,N_22782,N_22967);
nor U23184 (N_23184,N_22906,N_22661);
nand U23185 (N_23185,N_22504,N_22571);
or U23186 (N_23186,N_22794,N_22514);
nor U23187 (N_23187,N_22903,N_22865);
nor U23188 (N_23188,N_22921,N_22540);
nor U23189 (N_23189,N_22943,N_22949);
nor U23190 (N_23190,N_22537,N_22630);
xor U23191 (N_23191,N_22517,N_22520);
and U23192 (N_23192,N_22627,N_22740);
and U23193 (N_23193,N_23076,N_22969);
nor U23194 (N_23194,N_22635,N_22855);
nand U23195 (N_23195,N_22705,N_22956);
and U23196 (N_23196,N_23045,N_22647);
and U23197 (N_23197,N_22516,N_22763);
nor U23198 (N_23198,N_22838,N_22673);
nor U23199 (N_23199,N_22797,N_23051);
and U23200 (N_23200,N_22840,N_22766);
and U23201 (N_23201,N_22747,N_23057);
and U23202 (N_23202,N_22547,N_22778);
or U23203 (N_23203,N_22684,N_22987);
and U23204 (N_23204,N_23064,N_22722);
and U23205 (N_23205,N_23063,N_22780);
and U23206 (N_23206,N_22845,N_22689);
and U23207 (N_23207,N_23005,N_22631);
or U23208 (N_23208,N_22788,N_23086);
nor U23209 (N_23209,N_22580,N_22613);
or U23210 (N_23210,N_22622,N_22595);
nand U23211 (N_23211,N_22885,N_23088);
and U23212 (N_23212,N_22732,N_22660);
or U23213 (N_23213,N_23031,N_22968);
xnor U23214 (N_23214,N_22694,N_22526);
nand U23215 (N_23215,N_23029,N_22707);
nor U23216 (N_23216,N_22519,N_23004);
nand U23217 (N_23217,N_22842,N_22950);
xor U23218 (N_23218,N_22604,N_22721);
and U23219 (N_23219,N_22822,N_22952);
or U23220 (N_23220,N_22643,N_22752);
nor U23221 (N_23221,N_22974,N_22991);
or U23222 (N_23222,N_22570,N_22853);
nor U23223 (N_23223,N_22650,N_22786);
or U23224 (N_23224,N_23014,N_22897);
nor U23225 (N_23225,N_22592,N_22523);
nor U23226 (N_23226,N_23065,N_22541);
and U23227 (N_23227,N_22533,N_22936);
xnor U23228 (N_23228,N_22951,N_22873);
nand U23229 (N_23229,N_22569,N_22737);
nor U23230 (N_23230,N_23049,N_23073);
and U23231 (N_23231,N_22962,N_23105);
nor U23232 (N_23232,N_22879,N_22657);
nor U23233 (N_23233,N_22579,N_22875);
nand U23234 (N_23234,N_22699,N_22795);
nor U23235 (N_23235,N_22964,N_22848);
nand U23236 (N_23236,N_22771,N_22857);
nand U23237 (N_23237,N_22709,N_22819);
xor U23238 (N_23238,N_22847,N_23124);
and U23239 (N_23239,N_23037,N_22813);
and U23240 (N_23240,N_23042,N_22767);
and U23241 (N_23241,N_23050,N_23075);
and U23242 (N_23242,N_22671,N_22557);
and U23243 (N_23243,N_22596,N_22664);
nor U23244 (N_23244,N_22787,N_22586);
or U23245 (N_23245,N_22980,N_23019);
nor U23246 (N_23246,N_22900,N_22828);
and U23247 (N_23247,N_22544,N_22560);
and U23248 (N_23248,N_22772,N_22730);
nand U23249 (N_23249,N_22901,N_23055);
and U23250 (N_23250,N_22930,N_22733);
and U23251 (N_23251,N_22715,N_22841);
xnor U23252 (N_23252,N_22666,N_22701);
nand U23253 (N_23253,N_22536,N_22552);
nand U23254 (N_23254,N_22688,N_22881);
and U23255 (N_23255,N_23046,N_22779);
or U23256 (N_23256,N_23082,N_22898);
xnor U23257 (N_23257,N_22940,N_22909);
nand U23258 (N_23258,N_23093,N_22808);
and U23259 (N_23259,N_22521,N_22843);
or U23260 (N_23260,N_22578,N_22777);
nand U23261 (N_23261,N_22994,N_22508);
and U23262 (N_23262,N_22978,N_22863);
nand U23263 (N_23263,N_22804,N_22892);
nor U23264 (N_23264,N_23119,N_22746);
nand U23265 (N_23265,N_22776,N_23038);
and U23266 (N_23266,N_22572,N_22644);
nand U23267 (N_23267,N_23094,N_22558);
or U23268 (N_23268,N_22648,N_23039);
nor U23269 (N_23269,N_23121,N_23043);
nor U23270 (N_23270,N_23110,N_22503);
or U23271 (N_23271,N_22690,N_22736);
nor U23272 (N_23272,N_22658,N_22966);
and U23273 (N_23273,N_23016,N_23098);
nor U23274 (N_23274,N_22836,N_22770);
or U23275 (N_23275,N_23102,N_22567);
nand U23276 (N_23276,N_23072,N_22758);
nor U23277 (N_23277,N_22574,N_22769);
xnor U23278 (N_23278,N_23116,N_22826);
nand U23279 (N_23279,N_22871,N_23085);
nand U23280 (N_23280,N_22591,N_22982);
nor U23281 (N_23281,N_22618,N_22696);
nand U23282 (N_23282,N_22575,N_22686);
nor U23283 (N_23283,N_22607,N_22501);
xnor U23284 (N_23284,N_23036,N_22761);
or U23285 (N_23285,N_22549,N_22913);
nor U23286 (N_23286,N_22669,N_22965);
and U23287 (N_23287,N_23106,N_22554);
nand U23288 (N_23288,N_22911,N_22883);
nor U23289 (N_23289,N_22624,N_22829);
nor U23290 (N_23290,N_22515,N_22734);
and U23291 (N_23291,N_22933,N_22889);
and U23292 (N_23292,N_22634,N_22870);
nor U23293 (N_23293,N_23080,N_22697);
or U23294 (N_23294,N_22564,N_22990);
nand U23295 (N_23295,N_22937,N_22509);
and U23296 (N_23296,N_22852,N_22706);
and U23297 (N_23297,N_22944,N_22839);
nand U23298 (N_23298,N_22750,N_22615);
nand U23299 (N_23299,N_23009,N_23115);
and U23300 (N_23300,N_23071,N_23002);
and U23301 (N_23301,N_22947,N_23054);
or U23302 (N_23302,N_22620,N_22609);
nor U23303 (N_23303,N_22886,N_22693);
nand U23304 (N_23304,N_22816,N_22680);
xnor U23305 (N_23305,N_22731,N_22832);
and U23306 (N_23306,N_22675,N_22550);
and U23307 (N_23307,N_22757,N_22603);
and U23308 (N_23308,N_22806,N_22612);
nor U23309 (N_23309,N_23015,N_23096);
and U23310 (N_23310,N_22745,N_22638);
and U23311 (N_23311,N_22649,N_22981);
or U23312 (N_23312,N_22506,N_23099);
nand U23313 (N_23313,N_22760,N_22559);
nor U23314 (N_23314,N_23103,N_22945);
nand U23315 (N_23315,N_22908,N_22632);
nor U23316 (N_23316,N_22667,N_22677);
nor U23317 (N_23317,N_22880,N_22932);
or U23318 (N_23318,N_22513,N_22992);
or U23319 (N_23319,N_22924,N_22553);
and U23320 (N_23320,N_22869,N_22790);
or U23321 (N_23321,N_23044,N_22543);
nor U23322 (N_23322,N_22888,N_22565);
nor U23323 (N_23323,N_23060,N_22961);
xor U23324 (N_23324,N_23058,N_23040);
nor U23325 (N_23325,N_22742,N_22914);
or U23326 (N_23326,N_23067,N_22934);
and U23327 (N_23327,N_22942,N_23003);
or U23328 (N_23328,N_22867,N_22524);
nor U23329 (N_23329,N_22726,N_23089);
nand U23330 (N_23330,N_22872,N_22803);
and U23331 (N_23331,N_22692,N_23091);
and U23332 (N_23332,N_22585,N_22801);
and U23333 (N_23333,N_22700,N_22876);
or U23334 (N_23334,N_22628,N_22918);
nor U23335 (N_23335,N_22957,N_22751);
xor U23336 (N_23336,N_22846,N_22837);
nand U23337 (N_23337,N_22941,N_22718);
nor U23338 (N_23338,N_23069,N_23100);
nand U23339 (N_23339,N_22854,N_23013);
nor U23340 (N_23340,N_22584,N_22977);
nand U23341 (N_23341,N_23026,N_23087);
and U23342 (N_23342,N_23083,N_22939);
nor U23343 (N_23343,N_22670,N_23084);
or U23344 (N_23344,N_23120,N_22823);
nor U23345 (N_23345,N_23032,N_22831);
nor U23346 (N_23346,N_23024,N_23092);
and U23347 (N_23347,N_22948,N_23008);
xor U23348 (N_23348,N_22633,N_23021);
or U23349 (N_23349,N_22919,N_22783);
nor U23350 (N_23350,N_22946,N_22807);
or U23351 (N_23351,N_22820,N_22717);
nand U23352 (N_23352,N_22663,N_22858);
nand U23353 (N_23353,N_22594,N_22866);
and U23354 (N_23354,N_22756,N_22502);
nor U23355 (N_23355,N_22527,N_22525);
nand U23356 (N_23356,N_22986,N_22678);
xor U23357 (N_23357,N_22835,N_22566);
xor U23358 (N_23358,N_23047,N_22683);
and U23359 (N_23359,N_22507,N_22920);
and U23360 (N_23360,N_22606,N_22983);
or U23361 (N_23361,N_22621,N_22702);
xor U23362 (N_23362,N_22811,N_22935);
nor U23363 (N_23363,N_23070,N_22614);
xor U23364 (N_23364,N_22735,N_22522);
and U23365 (N_23365,N_22639,N_22590);
nand U23366 (N_23366,N_23025,N_22642);
nor U23367 (N_23367,N_22844,N_22860);
or U23368 (N_23368,N_22729,N_22834);
or U23369 (N_23369,N_23056,N_22587);
nand U23370 (N_23370,N_22796,N_22793);
and U23371 (N_23371,N_22764,N_23001);
xor U23372 (N_23372,N_22576,N_22556);
or U23373 (N_23373,N_23118,N_22799);
and U23374 (N_23374,N_22789,N_22728);
nand U23375 (N_23375,N_23097,N_22884);
nor U23376 (N_23376,N_22925,N_22637);
xnor U23377 (N_23377,N_22636,N_22748);
or U23378 (N_23378,N_22818,N_23107);
nand U23379 (N_23379,N_22720,N_22645);
nand U23380 (N_23380,N_22741,N_22993);
nand U23381 (N_23381,N_22600,N_22973);
or U23382 (N_23382,N_22599,N_22651);
nand U23383 (N_23383,N_23028,N_22510);
nor U23384 (N_23384,N_22988,N_22710);
nor U23385 (N_23385,N_22538,N_22563);
nor U23386 (N_23386,N_23117,N_22907);
nand U23387 (N_23387,N_22713,N_22681);
nor U23388 (N_23388,N_23010,N_22851);
xor U23389 (N_23389,N_22887,N_22668);
nor U23390 (N_23390,N_22695,N_22791);
or U23391 (N_23391,N_22984,N_22712);
nand U23392 (N_23392,N_22997,N_22598);
nor U23393 (N_23393,N_22775,N_23114);
nor U23394 (N_23394,N_23017,N_22915);
xnor U23395 (N_23395,N_22676,N_22577);
xnor U23396 (N_23396,N_22916,N_22539);
or U23397 (N_23397,N_23018,N_23077);
nor U23398 (N_23398,N_22995,N_22910);
nand U23399 (N_23399,N_22698,N_23095);
nor U23400 (N_23400,N_23022,N_22976);
nand U23401 (N_23401,N_22723,N_22862);
nor U23402 (N_23402,N_22765,N_22589);
and U23403 (N_23403,N_22905,N_22792);
nor U23404 (N_23404,N_22674,N_22809);
and U23405 (N_23405,N_22714,N_22859);
nor U23406 (N_23406,N_22593,N_23033);
or U23407 (N_23407,N_22727,N_22530);
or U23408 (N_23408,N_22960,N_22608);
or U23409 (N_23409,N_22611,N_22922);
or U23410 (N_23410,N_22849,N_23066);
nand U23411 (N_23411,N_22996,N_23035);
and U23412 (N_23412,N_22890,N_22864);
nor U23413 (N_23413,N_22861,N_22505);
nor U23414 (N_23414,N_22561,N_22929);
xnor U23415 (N_23415,N_22827,N_22588);
and U23416 (N_23416,N_23030,N_22755);
nand U23417 (N_23417,N_22955,N_22654);
and U23418 (N_23418,N_22616,N_22902);
nor U23419 (N_23419,N_22719,N_22878);
nor U23420 (N_23420,N_23020,N_22531);
nor U23421 (N_23421,N_22665,N_22926);
nand U23422 (N_23422,N_22894,N_23011);
nor U23423 (N_23423,N_22605,N_22923);
nand U23424 (N_23424,N_22856,N_22759);
and U23425 (N_23425,N_23006,N_23052);
nand U23426 (N_23426,N_23034,N_22739);
or U23427 (N_23427,N_22687,N_22784);
and U23428 (N_23428,N_22768,N_22548);
or U23429 (N_23429,N_22623,N_23068);
nand U23430 (N_23430,N_22653,N_22975);
and U23431 (N_23431,N_22800,N_22958);
or U23432 (N_23432,N_22749,N_23079);
nor U23433 (N_23433,N_22646,N_22528);
nor U23434 (N_23434,N_22754,N_22998);
xor U23435 (N_23435,N_22679,N_22532);
nor U23436 (N_23436,N_22833,N_22815);
and U23437 (N_23437,N_22511,N_22768);
nand U23438 (N_23438,N_22878,N_22614);
and U23439 (N_23439,N_22822,N_22842);
xor U23440 (N_23440,N_22769,N_22819);
nor U23441 (N_23441,N_23073,N_23078);
and U23442 (N_23442,N_22840,N_22663);
nor U23443 (N_23443,N_22987,N_22673);
nand U23444 (N_23444,N_22970,N_22618);
nand U23445 (N_23445,N_22740,N_23046);
or U23446 (N_23446,N_22827,N_22553);
or U23447 (N_23447,N_23091,N_22988);
xnor U23448 (N_23448,N_22897,N_22604);
or U23449 (N_23449,N_22746,N_22683);
and U23450 (N_23450,N_22666,N_22564);
and U23451 (N_23451,N_22798,N_23102);
nand U23452 (N_23452,N_23005,N_22600);
xnor U23453 (N_23453,N_22625,N_22896);
nor U23454 (N_23454,N_22627,N_22519);
and U23455 (N_23455,N_23119,N_22979);
nor U23456 (N_23456,N_22678,N_22828);
nor U23457 (N_23457,N_22675,N_22965);
and U23458 (N_23458,N_22999,N_23076);
nor U23459 (N_23459,N_22536,N_22964);
and U23460 (N_23460,N_22563,N_23122);
and U23461 (N_23461,N_23073,N_22730);
nor U23462 (N_23462,N_22707,N_23025);
nand U23463 (N_23463,N_22896,N_22779);
and U23464 (N_23464,N_22676,N_22548);
or U23465 (N_23465,N_23026,N_22621);
nor U23466 (N_23466,N_23005,N_22546);
nand U23467 (N_23467,N_23050,N_22878);
nor U23468 (N_23468,N_22877,N_22753);
and U23469 (N_23469,N_22950,N_23078);
nor U23470 (N_23470,N_22874,N_22647);
nor U23471 (N_23471,N_22538,N_22855);
nand U23472 (N_23472,N_22918,N_22840);
or U23473 (N_23473,N_22806,N_22811);
nor U23474 (N_23474,N_22512,N_22855);
nor U23475 (N_23475,N_22584,N_22582);
and U23476 (N_23476,N_22796,N_23045);
and U23477 (N_23477,N_22539,N_22500);
nor U23478 (N_23478,N_22755,N_23034);
nand U23479 (N_23479,N_23102,N_22867);
nor U23480 (N_23480,N_22709,N_22560);
nand U23481 (N_23481,N_22997,N_22637);
or U23482 (N_23482,N_22779,N_22951);
nor U23483 (N_23483,N_22555,N_23089);
or U23484 (N_23484,N_22815,N_23000);
nor U23485 (N_23485,N_22663,N_22576);
or U23486 (N_23486,N_22923,N_22627);
nor U23487 (N_23487,N_22992,N_22923);
and U23488 (N_23488,N_22998,N_22601);
nor U23489 (N_23489,N_22927,N_22588);
and U23490 (N_23490,N_22630,N_22675);
and U23491 (N_23491,N_23056,N_22756);
xor U23492 (N_23492,N_22993,N_22586);
and U23493 (N_23493,N_22893,N_23022);
or U23494 (N_23494,N_22514,N_22727);
or U23495 (N_23495,N_22926,N_23067);
or U23496 (N_23496,N_22768,N_22681);
nand U23497 (N_23497,N_23122,N_22520);
and U23498 (N_23498,N_23013,N_22689);
or U23499 (N_23499,N_22937,N_22814);
and U23500 (N_23500,N_22659,N_22558);
nor U23501 (N_23501,N_22626,N_22909);
and U23502 (N_23502,N_22918,N_22560);
nor U23503 (N_23503,N_23122,N_22562);
or U23504 (N_23504,N_22668,N_23033);
nor U23505 (N_23505,N_22863,N_23041);
and U23506 (N_23506,N_22912,N_22909);
or U23507 (N_23507,N_22938,N_22992);
xnor U23508 (N_23508,N_22597,N_22904);
xnor U23509 (N_23509,N_22702,N_22644);
or U23510 (N_23510,N_22963,N_22738);
nand U23511 (N_23511,N_22829,N_22988);
or U23512 (N_23512,N_23082,N_22877);
nor U23513 (N_23513,N_23025,N_22597);
or U23514 (N_23514,N_22722,N_22760);
nand U23515 (N_23515,N_22887,N_22766);
and U23516 (N_23516,N_22936,N_22689);
nor U23517 (N_23517,N_22620,N_22700);
nor U23518 (N_23518,N_22963,N_22762);
nand U23519 (N_23519,N_22686,N_22997);
nor U23520 (N_23520,N_22647,N_22860);
and U23521 (N_23521,N_22988,N_23038);
or U23522 (N_23522,N_22972,N_22832);
and U23523 (N_23523,N_22731,N_22684);
xnor U23524 (N_23524,N_22500,N_22868);
nor U23525 (N_23525,N_22893,N_22727);
nor U23526 (N_23526,N_22775,N_22828);
nor U23527 (N_23527,N_22718,N_22553);
xnor U23528 (N_23528,N_22757,N_23002);
nor U23529 (N_23529,N_22764,N_22568);
xnor U23530 (N_23530,N_22684,N_22599);
nor U23531 (N_23531,N_22812,N_22609);
and U23532 (N_23532,N_22597,N_23123);
and U23533 (N_23533,N_23037,N_22582);
nand U23534 (N_23534,N_22670,N_22511);
or U23535 (N_23535,N_22641,N_22893);
and U23536 (N_23536,N_22816,N_22826);
or U23537 (N_23537,N_22527,N_22934);
nand U23538 (N_23538,N_22520,N_22956);
or U23539 (N_23539,N_22510,N_22588);
nand U23540 (N_23540,N_22599,N_22739);
nand U23541 (N_23541,N_22909,N_22502);
or U23542 (N_23542,N_22979,N_22899);
and U23543 (N_23543,N_22980,N_22582);
nand U23544 (N_23544,N_22654,N_22882);
or U23545 (N_23545,N_23054,N_22771);
or U23546 (N_23546,N_22607,N_22650);
nor U23547 (N_23547,N_22672,N_22797);
xor U23548 (N_23548,N_22654,N_22873);
nand U23549 (N_23549,N_23094,N_22842);
and U23550 (N_23550,N_22674,N_22730);
nand U23551 (N_23551,N_23004,N_22548);
or U23552 (N_23552,N_23087,N_22583);
nand U23553 (N_23553,N_22771,N_23111);
nor U23554 (N_23554,N_23035,N_22654);
nand U23555 (N_23555,N_22689,N_22628);
or U23556 (N_23556,N_22803,N_22549);
and U23557 (N_23557,N_22904,N_22782);
and U23558 (N_23558,N_22537,N_22584);
nand U23559 (N_23559,N_22974,N_22697);
nor U23560 (N_23560,N_22978,N_22834);
nand U23561 (N_23561,N_22538,N_22585);
nor U23562 (N_23562,N_23123,N_22917);
xnor U23563 (N_23563,N_22562,N_22937);
nor U23564 (N_23564,N_22504,N_22731);
and U23565 (N_23565,N_22563,N_22951);
and U23566 (N_23566,N_22737,N_23033);
nor U23567 (N_23567,N_22838,N_22522);
and U23568 (N_23568,N_22509,N_23004);
or U23569 (N_23569,N_22836,N_22842);
nor U23570 (N_23570,N_22606,N_23057);
or U23571 (N_23571,N_23111,N_23010);
and U23572 (N_23572,N_22757,N_23081);
nor U23573 (N_23573,N_22607,N_22917);
nor U23574 (N_23574,N_23045,N_22539);
xor U23575 (N_23575,N_23047,N_22699);
and U23576 (N_23576,N_22881,N_22763);
nor U23577 (N_23577,N_22534,N_22514);
nand U23578 (N_23578,N_22838,N_22718);
or U23579 (N_23579,N_22884,N_22785);
nand U23580 (N_23580,N_23081,N_22793);
nor U23581 (N_23581,N_22737,N_22931);
nor U23582 (N_23582,N_22732,N_23069);
xnor U23583 (N_23583,N_22922,N_22612);
nand U23584 (N_23584,N_22949,N_22791);
nor U23585 (N_23585,N_22943,N_23085);
xor U23586 (N_23586,N_22728,N_22937);
or U23587 (N_23587,N_22507,N_22513);
or U23588 (N_23588,N_22983,N_22970);
and U23589 (N_23589,N_23008,N_22892);
nand U23590 (N_23590,N_22954,N_23092);
nand U23591 (N_23591,N_22963,N_22888);
nor U23592 (N_23592,N_23001,N_22605);
nor U23593 (N_23593,N_23043,N_22727);
nor U23594 (N_23594,N_22554,N_22550);
or U23595 (N_23595,N_23053,N_23005);
or U23596 (N_23596,N_22988,N_22612);
and U23597 (N_23597,N_23046,N_23110);
nand U23598 (N_23598,N_22802,N_22593);
and U23599 (N_23599,N_22780,N_23098);
and U23600 (N_23600,N_22528,N_22647);
and U23601 (N_23601,N_22932,N_22709);
or U23602 (N_23602,N_22838,N_22967);
or U23603 (N_23603,N_22932,N_22961);
and U23604 (N_23604,N_22856,N_23113);
nor U23605 (N_23605,N_22606,N_22852);
xor U23606 (N_23606,N_22552,N_22700);
or U23607 (N_23607,N_22612,N_23036);
nor U23608 (N_23608,N_23113,N_22773);
or U23609 (N_23609,N_22623,N_22567);
nand U23610 (N_23610,N_23115,N_23054);
nor U23611 (N_23611,N_23120,N_22633);
nand U23612 (N_23612,N_22654,N_22990);
nor U23613 (N_23613,N_23054,N_22847);
or U23614 (N_23614,N_22626,N_22818);
and U23615 (N_23615,N_22646,N_22966);
and U23616 (N_23616,N_22895,N_22789);
and U23617 (N_23617,N_22991,N_22533);
nand U23618 (N_23618,N_22913,N_22918);
or U23619 (N_23619,N_22868,N_22709);
nand U23620 (N_23620,N_22746,N_22698);
and U23621 (N_23621,N_22688,N_23105);
nand U23622 (N_23622,N_22917,N_23122);
and U23623 (N_23623,N_22669,N_22874);
nand U23624 (N_23624,N_22867,N_23058);
nand U23625 (N_23625,N_22672,N_22743);
nand U23626 (N_23626,N_22971,N_22613);
nand U23627 (N_23627,N_22849,N_22595);
or U23628 (N_23628,N_22681,N_22562);
nor U23629 (N_23629,N_22731,N_23108);
nand U23630 (N_23630,N_22783,N_23054);
and U23631 (N_23631,N_22862,N_22549);
and U23632 (N_23632,N_22862,N_22886);
nor U23633 (N_23633,N_23008,N_23110);
nor U23634 (N_23634,N_22503,N_22688);
nor U23635 (N_23635,N_22947,N_22700);
nand U23636 (N_23636,N_22909,N_22775);
xnor U23637 (N_23637,N_22801,N_23105);
nor U23638 (N_23638,N_22819,N_22679);
or U23639 (N_23639,N_22643,N_22968);
xor U23640 (N_23640,N_22898,N_23049);
and U23641 (N_23641,N_22982,N_22569);
nor U23642 (N_23642,N_22920,N_23111);
xor U23643 (N_23643,N_23062,N_22578);
nand U23644 (N_23644,N_22590,N_23005);
nand U23645 (N_23645,N_23025,N_22860);
or U23646 (N_23646,N_22775,N_22760);
nor U23647 (N_23647,N_22791,N_22650);
nand U23648 (N_23648,N_22775,N_22652);
and U23649 (N_23649,N_22600,N_22902);
or U23650 (N_23650,N_22853,N_22995);
and U23651 (N_23651,N_22879,N_22941);
nor U23652 (N_23652,N_22536,N_22791);
nand U23653 (N_23653,N_23070,N_22785);
nor U23654 (N_23654,N_22659,N_23062);
nor U23655 (N_23655,N_22895,N_22827);
and U23656 (N_23656,N_22514,N_22746);
or U23657 (N_23657,N_22750,N_22819);
or U23658 (N_23658,N_22524,N_22671);
or U23659 (N_23659,N_22916,N_22853);
and U23660 (N_23660,N_23049,N_23050);
and U23661 (N_23661,N_22509,N_22830);
xor U23662 (N_23662,N_23014,N_23034);
nand U23663 (N_23663,N_22734,N_22656);
and U23664 (N_23664,N_22626,N_22729);
or U23665 (N_23665,N_23087,N_22960);
or U23666 (N_23666,N_23009,N_22558);
nand U23667 (N_23667,N_22841,N_22633);
xnor U23668 (N_23668,N_23085,N_22617);
xnor U23669 (N_23669,N_22754,N_23107);
or U23670 (N_23670,N_22638,N_23119);
and U23671 (N_23671,N_22688,N_22615);
xor U23672 (N_23672,N_22761,N_22629);
nand U23673 (N_23673,N_22873,N_22739);
nor U23674 (N_23674,N_22700,N_22820);
or U23675 (N_23675,N_22586,N_22776);
nor U23676 (N_23676,N_22849,N_22810);
or U23677 (N_23677,N_23109,N_22934);
nor U23678 (N_23678,N_22893,N_22913);
nand U23679 (N_23679,N_22709,N_22684);
or U23680 (N_23680,N_22543,N_22723);
nand U23681 (N_23681,N_23047,N_22739);
xor U23682 (N_23682,N_22803,N_22988);
xor U23683 (N_23683,N_22612,N_22881);
xnor U23684 (N_23684,N_23078,N_22820);
and U23685 (N_23685,N_22742,N_22937);
and U23686 (N_23686,N_22893,N_22606);
nor U23687 (N_23687,N_22774,N_22869);
nor U23688 (N_23688,N_22595,N_22901);
or U23689 (N_23689,N_23064,N_22813);
nor U23690 (N_23690,N_22677,N_23121);
or U23691 (N_23691,N_22663,N_22681);
nor U23692 (N_23692,N_23074,N_22664);
nand U23693 (N_23693,N_22602,N_22527);
and U23694 (N_23694,N_22717,N_23119);
and U23695 (N_23695,N_23118,N_23005);
and U23696 (N_23696,N_22845,N_22520);
nand U23697 (N_23697,N_23110,N_23033);
nand U23698 (N_23698,N_22979,N_22887);
nor U23699 (N_23699,N_22882,N_22700);
nor U23700 (N_23700,N_23012,N_22826);
or U23701 (N_23701,N_22596,N_22829);
or U23702 (N_23702,N_23006,N_22909);
xor U23703 (N_23703,N_22608,N_23016);
or U23704 (N_23704,N_23026,N_22894);
nand U23705 (N_23705,N_22774,N_22618);
and U23706 (N_23706,N_22879,N_22564);
nor U23707 (N_23707,N_22905,N_22737);
nor U23708 (N_23708,N_23030,N_22718);
or U23709 (N_23709,N_22878,N_22673);
nor U23710 (N_23710,N_22968,N_22772);
or U23711 (N_23711,N_22535,N_22960);
or U23712 (N_23712,N_22702,N_22611);
or U23713 (N_23713,N_23070,N_22735);
nor U23714 (N_23714,N_22617,N_22879);
and U23715 (N_23715,N_22979,N_22811);
and U23716 (N_23716,N_22921,N_22977);
nor U23717 (N_23717,N_22759,N_23102);
or U23718 (N_23718,N_23096,N_22803);
nand U23719 (N_23719,N_22721,N_22623);
xor U23720 (N_23720,N_22600,N_22669);
nand U23721 (N_23721,N_22968,N_22610);
nand U23722 (N_23722,N_22891,N_22859);
nand U23723 (N_23723,N_22840,N_22821);
and U23724 (N_23724,N_22898,N_23015);
nand U23725 (N_23725,N_22640,N_23010);
nand U23726 (N_23726,N_23111,N_22883);
or U23727 (N_23727,N_22525,N_22984);
or U23728 (N_23728,N_22584,N_22764);
nand U23729 (N_23729,N_22548,N_23079);
or U23730 (N_23730,N_22504,N_22826);
nor U23731 (N_23731,N_22665,N_22649);
and U23732 (N_23732,N_22926,N_23000);
nor U23733 (N_23733,N_22959,N_22802);
and U23734 (N_23734,N_22884,N_23022);
and U23735 (N_23735,N_22535,N_22619);
nor U23736 (N_23736,N_22601,N_22608);
and U23737 (N_23737,N_23004,N_22863);
nor U23738 (N_23738,N_22873,N_22663);
nand U23739 (N_23739,N_22743,N_22573);
nor U23740 (N_23740,N_23076,N_23067);
nand U23741 (N_23741,N_22943,N_22784);
nor U23742 (N_23742,N_23087,N_22846);
nor U23743 (N_23743,N_22539,N_22553);
xor U23744 (N_23744,N_22647,N_22852);
nand U23745 (N_23745,N_23000,N_22658);
nor U23746 (N_23746,N_22531,N_22733);
nand U23747 (N_23747,N_22856,N_22502);
or U23748 (N_23748,N_22719,N_22685);
nor U23749 (N_23749,N_22588,N_22963);
or U23750 (N_23750,N_23474,N_23710);
or U23751 (N_23751,N_23545,N_23567);
nand U23752 (N_23752,N_23221,N_23126);
and U23753 (N_23753,N_23262,N_23329);
and U23754 (N_23754,N_23463,N_23723);
or U23755 (N_23755,N_23226,N_23747);
and U23756 (N_23756,N_23610,N_23658);
nand U23757 (N_23757,N_23568,N_23408);
or U23758 (N_23758,N_23456,N_23331);
or U23759 (N_23759,N_23500,N_23523);
and U23760 (N_23760,N_23376,N_23427);
nand U23761 (N_23761,N_23302,N_23194);
and U23762 (N_23762,N_23664,N_23692);
nand U23763 (N_23763,N_23406,N_23395);
nand U23764 (N_23764,N_23219,N_23193);
xor U23765 (N_23765,N_23371,N_23158);
nor U23766 (N_23766,N_23538,N_23187);
nor U23767 (N_23767,N_23480,N_23272);
and U23768 (N_23768,N_23301,N_23624);
nor U23769 (N_23769,N_23482,N_23281);
nand U23770 (N_23770,N_23127,N_23398);
and U23771 (N_23771,N_23288,N_23514);
nor U23772 (N_23772,N_23240,N_23731);
nor U23773 (N_23773,N_23481,N_23612);
nor U23774 (N_23774,N_23393,N_23615);
nand U23775 (N_23775,N_23591,N_23254);
and U23776 (N_23776,N_23597,N_23143);
xor U23777 (N_23777,N_23222,N_23726);
nand U23778 (N_23778,N_23330,N_23423);
nor U23779 (N_23779,N_23713,N_23182);
xnor U23780 (N_23780,N_23571,N_23552);
nor U23781 (N_23781,N_23244,N_23327);
nand U23782 (N_23782,N_23241,N_23672);
xnor U23783 (N_23783,N_23377,N_23201);
or U23784 (N_23784,N_23231,N_23239);
nand U23785 (N_23785,N_23172,N_23163);
nand U23786 (N_23786,N_23146,N_23652);
nor U23787 (N_23787,N_23602,N_23333);
nor U23788 (N_23788,N_23196,N_23447);
xnor U23789 (N_23789,N_23295,N_23347);
or U23790 (N_23790,N_23375,N_23342);
or U23791 (N_23791,N_23677,N_23698);
and U23792 (N_23792,N_23186,N_23515);
or U23793 (N_23793,N_23412,N_23562);
nand U23794 (N_23794,N_23598,N_23687);
nand U23795 (N_23795,N_23669,N_23537);
or U23796 (N_23796,N_23583,N_23703);
nor U23797 (N_23797,N_23697,N_23223);
and U23798 (N_23798,N_23259,N_23180);
nand U23799 (N_23799,N_23540,N_23305);
nand U23800 (N_23800,N_23472,N_23142);
nor U23801 (N_23801,N_23264,N_23550);
or U23802 (N_23802,N_23149,N_23506);
and U23803 (N_23803,N_23434,N_23576);
and U23804 (N_23804,N_23654,N_23720);
or U23805 (N_23805,N_23675,N_23736);
nand U23806 (N_23806,N_23138,N_23251);
and U23807 (N_23807,N_23352,N_23715);
nand U23808 (N_23808,N_23509,N_23185);
xor U23809 (N_23809,N_23269,N_23220);
and U23810 (N_23810,N_23348,N_23203);
nor U23811 (N_23811,N_23508,N_23202);
and U23812 (N_23812,N_23199,N_23385);
nand U23813 (N_23813,N_23601,N_23666);
nand U23814 (N_23814,N_23643,N_23246);
nand U23815 (N_23815,N_23167,N_23326);
and U23816 (N_23816,N_23581,N_23455);
xor U23817 (N_23817,N_23526,N_23634);
nor U23818 (N_23818,N_23743,N_23569);
nand U23819 (N_23819,N_23245,N_23700);
nand U23820 (N_23820,N_23641,N_23466);
nor U23821 (N_23821,N_23378,N_23467);
or U23822 (N_23822,N_23527,N_23594);
or U23823 (N_23823,N_23656,N_23243);
xor U23824 (N_23824,N_23546,N_23418);
or U23825 (N_23825,N_23315,N_23283);
and U23826 (N_23826,N_23425,N_23516);
nand U23827 (N_23827,N_23582,N_23608);
and U23828 (N_23828,N_23183,N_23670);
nor U23829 (N_23829,N_23536,N_23213);
nor U23830 (N_23830,N_23618,N_23438);
nor U23831 (N_23831,N_23486,N_23528);
or U23832 (N_23832,N_23225,N_23464);
or U23833 (N_23833,N_23135,N_23188);
or U23834 (N_23834,N_23603,N_23533);
nor U23835 (N_23835,N_23717,N_23144);
nor U23836 (N_23836,N_23334,N_23555);
nor U23837 (N_23837,N_23367,N_23255);
and U23838 (N_23838,N_23414,N_23492);
nand U23839 (N_23839,N_23745,N_23746);
nor U23840 (N_23840,N_23340,N_23577);
or U23841 (N_23841,N_23310,N_23517);
and U23842 (N_23842,N_23534,N_23630);
and U23843 (N_23843,N_23542,N_23729);
nand U23844 (N_23844,N_23169,N_23626);
nand U23845 (N_23845,N_23140,N_23179);
xor U23846 (N_23846,N_23308,N_23679);
nor U23847 (N_23847,N_23356,N_23446);
and U23848 (N_23848,N_23477,N_23312);
nor U23849 (N_23849,N_23361,N_23566);
and U23850 (N_23850,N_23659,N_23646);
xnor U23851 (N_23851,N_23572,N_23724);
nor U23852 (N_23852,N_23397,N_23354);
nand U23853 (N_23853,N_23580,N_23696);
or U23854 (N_23854,N_23217,N_23357);
or U23855 (N_23855,N_23307,N_23740);
and U23856 (N_23856,N_23504,N_23741);
nand U23857 (N_23857,N_23197,N_23475);
or U23858 (N_23858,N_23265,N_23511);
and U23859 (N_23859,N_23407,N_23599);
or U23860 (N_23860,N_23323,N_23707);
xnor U23861 (N_23861,N_23725,N_23131);
or U23862 (N_23862,N_23564,N_23152);
or U23863 (N_23863,N_23284,N_23619);
nand U23864 (N_23864,N_23400,N_23346);
and U23865 (N_23865,N_23620,N_23294);
or U23866 (N_23866,N_23297,N_23543);
xnor U23867 (N_23867,N_23595,N_23683);
and U23868 (N_23868,N_23271,N_23399);
and U23869 (N_23869,N_23175,N_23607);
and U23870 (N_23870,N_23128,N_23212);
and U23871 (N_23871,N_23671,N_23476);
nand U23872 (N_23872,N_23667,N_23507);
or U23873 (N_23873,N_23473,N_23621);
and U23874 (N_23874,N_23350,N_23579);
nor U23875 (N_23875,N_23553,N_23332);
or U23876 (N_23876,N_23177,N_23639);
nand U23877 (N_23877,N_23233,N_23458);
and U23878 (N_23878,N_23200,N_23693);
xor U23879 (N_23879,N_23338,N_23403);
and U23880 (N_23880,N_23642,N_23211);
nand U23881 (N_23881,N_23487,N_23653);
and U23882 (N_23882,N_23409,N_23208);
nor U23883 (N_23883,N_23335,N_23428);
nand U23884 (N_23884,N_23228,N_23465);
xor U23885 (N_23885,N_23268,N_23229);
nand U23886 (N_23886,N_23558,N_23578);
or U23887 (N_23887,N_23242,N_23633);
or U23888 (N_23888,N_23270,N_23366);
or U23889 (N_23889,N_23640,N_23535);
or U23890 (N_23890,N_23164,N_23277);
xor U23891 (N_23891,N_23629,N_23593);
xor U23892 (N_23892,N_23496,N_23422);
or U23893 (N_23893,N_23449,N_23660);
nand U23894 (N_23894,N_23604,N_23650);
nand U23895 (N_23895,N_23573,N_23320);
or U23896 (N_23896,N_23191,N_23337);
or U23897 (N_23897,N_23325,N_23370);
nor U23898 (N_23898,N_23549,N_23575);
nor U23899 (N_23899,N_23735,N_23737);
nand U23900 (N_23900,N_23360,N_23234);
or U23901 (N_23901,N_23631,N_23627);
or U23902 (N_23902,N_23719,N_23645);
or U23903 (N_23903,N_23168,N_23133);
and U23904 (N_23904,N_23444,N_23362);
or U23905 (N_23905,N_23749,N_23391);
or U23906 (N_23906,N_23450,N_23192);
nand U23907 (N_23907,N_23129,N_23730);
or U23908 (N_23908,N_23299,N_23290);
or U23909 (N_23909,N_23153,N_23184);
and U23910 (N_23910,N_23285,N_23695);
and U23911 (N_23911,N_23166,N_23318);
or U23912 (N_23912,N_23556,N_23278);
and U23913 (N_23913,N_23457,N_23432);
or U23914 (N_23914,N_23637,N_23702);
and U23915 (N_23915,N_23328,N_23235);
nand U23916 (N_23916,N_23260,N_23287);
nand U23917 (N_23917,N_23663,N_23258);
nor U23918 (N_23918,N_23137,N_23648);
nor U23919 (N_23919,N_23539,N_23379);
or U23920 (N_23920,N_23586,N_23681);
nor U23921 (N_23921,N_23214,N_23635);
xnor U23922 (N_23922,N_23505,N_23661);
and U23923 (N_23923,N_23439,N_23417);
nor U23924 (N_23924,N_23532,N_23321);
nor U23925 (N_23925,N_23657,N_23388);
nand U23926 (N_23926,N_23596,N_23261);
nand U23927 (N_23927,N_23709,N_23491);
nor U23928 (N_23928,N_23130,N_23319);
or U23929 (N_23929,N_23704,N_23522);
and U23930 (N_23930,N_23588,N_23712);
nor U23931 (N_23931,N_23413,N_23565);
xor U23932 (N_23932,N_23364,N_23410);
and U23933 (N_23933,N_23353,N_23714);
xor U23934 (N_23934,N_23324,N_23380);
nand U23935 (N_23935,N_23402,N_23690);
and U23936 (N_23936,N_23382,N_23561);
nand U23937 (N_23937,N_23685,N_23253);
and U23938 (N_23938,N_23150,N_23744);
and U23939 (N_23939,N_23623,N_23125);
nand U23940 (N_23940,N_23512,N_23676);
nand U23941 (N_23941,N_23300,N_23174);
nor U23942 (N_23942,N_23273,N_23574);
and U23943 (N_23943,N_23738,N_23311);
nor U23944 (N_23944,N_23363,N_23647);
xnor U23945 (N_23945,N_23727,N_23453);
and U23946 (N_23946,N_23605,N_23651);
or U23947 (N_23947,N_23237,N_23665);
or U23948 (N_23948,N_23563,N_23430);
or U23949 (N_23949,N_23435,N_23470);
or U23950 (N_23950,N_23718,N_23613);
or U23951 (N_23951,N_23368,N_23419);
nor U23952 (N_23952,N_23339,N_23655);
nor U23953 (N_23953,N_23173,N_23673);
nand U23954 (N_23954,N_23494,N_23441);
or U23955 (N_23955,N_23165,N_23383);
and U23956 (N_23956,N_23279,N_23424);
or U23957 (N_23957,N_23694,N_23493);
or U23958 (N_23958,N_23345,N_23230);
nand U23959 (N_23959,N_23498,N_23195);
nand U23960 (N_23960,N_23742,N_23147);
xnor U23961 (N_23961,N_23734,N_23384);
and U23962 (N_23962,N_23181,N_23286);
or U23963 (N_23963,N_23547,N_23436);
nor U23964 (N_23964,N_23374,N_23448);
or U23965 (N_23965,N_23190,N_23132);
and U23966 (N_23966,N_23708,N_23349);
xor U23967 (N_23967,N_23411,N_23392);
and U23968 (N_23968,N_23682,N_23298);
and U23969 (N_23969,N_23401,N_23248);
or U23970 (N_23970,N_23587,N_23691);
and U23971 (N_23971,N_23267,N_23557);
nor U23972 (N_23972,N_23250,N_23289);
nand U23973 (N_23973,N_23592,N_23559);
and U23974 (N_23974,N_23151,N_23322);
and U23975 (N_23975,N_23554,N_23748);
and U23976 (N_23976,N_23451,N_23524);
nor U23977 (N_23977,N_23684,N_23495);
nor U23978 (N_23978,N_23644,N_23282);
and U23979 (N_23979,N_23236,N_23148);
and U23980 (N_23980,N_23513,N_23351);
nand U23981 (N_23981,N_23699,N_23689);
xor U23982 (N_23982,N_23204,N_23688);
nand U23983 (N_23983,N_23716,N_23161);
or U23984 (N_23984,N_23280,N_23154);
or U23985 (N_23985,N_23421,N_23291);
nor U23986 (N_23986,N_23454,N_23485);
nand U23987 (N_23987,N_23420,N_23306);
nand U23988 (N_23988,N_23227,N_23632);
nand U23989 (N_23989,N_23462,N_23484);
or U23990 (N_23990,N_23317,N_23590);
and U23991 (N_23991,N_23461,N_23359);
and U23992 (N_23992,N_23157,N_23215);
xnor U23993 (N_23993,N_23343,N_23452);
and U23994 (N_23994,N_23459,N_23155);
or U23995 (N_23995,N_23218,N_23560);
nor U23996 (N_23996,N_23649,N_23209);
nand U23997 (N_23997,N_23488,N_23156);
and U23998 (N_23998,N_23293,N_23674);
and U23999 (N_23999,N_23404,N_23551);
nand U24000 (N_24000,N_23739,N_23711);
or U24001 (N_24001,N_23178,N_23232);
and U24002 (N_24002,N_23609,N_23489);
nand U24003 (N_24003,N_23636,N_23381);
nor U24004 (N_24004,N_23510,N_23387);
xnor U24005 (N_24005,N_23274,N_23701);
nor U24006 (N_24006,N_23159,N_23266);
nor U24007 (N_24007,N_23443,N_23134);
nand U24008 (N_24008,N_23316,N_23314);
or U24009 (N_24009,N_23499,N_23389);
nand U24010 (N_24010,N_23405,N_23396);
or U24011 (N_24011,N_23622,N_23584);
or U24012 (N_24012,N_23503,N_23722);
and U24013 (N_24013,N_23136,N_23386);
and U24014 (N_24014,N_23252,N_23431);
nand U24015 (N_24015,N_23373,N_23468);
nand U24016 (N_24016,N_23176,N_23479);
and U24017 (N_24017,N_23390,N_23589);
and U24018 (N_24018,N_23478,N_23531);
or U24019 (N_24019,N_23616,N_23313);
nor U24020 (N_24020,N_23292,N_23336);
nand U24021 (N_24021,N_23600,N_23548);
nor U24022 (N_24022,N_23483,N_23570);
nand U24023 (N_24023,N_23525,N_23705);
nor U24024 (N_24024,N_23426,N_23490);
or U24025 (N_24025,N_23706,N_23606);
or U24026 (N_24026,N_23445,N_23249);
nand U24027 (N_24027,N_23309,N_23247);
and U24028 (N_24028,N_23519,N_23257);
nor U24029 (N_24029,N_23617,N_23372);
or U24030 (N_24030,N_23585,N_23721);
or U24031 (N_24031,N_23530,N_23275);
and U24032 (N_24032,N_23521,N_23415);
xnor U24033 (N_24033,N_23303,N_23141);
and U24034 (N_24034,N_23341,N_23469);
and U24035 (N_24035,N_23638,N_23440);
and U24036 (N_24036,N_23520,N_23502);
and U24037 (N_24037,N_23369,N_23437);
nor U24038 (N_24038,N_23442,N_23518);
and U24039 (N_24039,N_23296,N_23139);
nand U24040 (N_24040,N_23614,N_23205);
nand U24041 (N_24041,N_23678,N_23662);
and U24042 (N_24042,N_23344,N_23732);
and U24043 (N_24043,N_23628,N_23501);
or U24044 (N_24044,N_23433,N_23668);
nand U24045 (N_24045,N_23224,N_23210);
and U24046 (N_24046,N_23170,N_23206);
nand U24047 (N_24047,N_23611,N_23529);
nand U24048 (N_24048,N_23686,N_23733);
nand U24049 (N_24049,N_23416,N_23544);
nand U24050 (N_24050,N_23171,N_23460);
or U24051 (N_24051,N_23160,N_23276);
or U24052 (N_24052,N_23198,N_23304);
nand U24053 (N_24053,N_23471,N_23189);
nor U24054 (N_24054,N_23394,N_23162);
xnor U24055 (N_24055,N_23355,N_23365);
and U24056 (N_24056,N_23625,N_23256);
and U24057 (N_24057,N_23541,N_23207);
and U24058 (N_24058,N_23238,N_23358);
nand U24059 (N_24059,N_23145,N_23728);
nand U24060 (N_24060,N_23429,N_23263);
and U24061 (N_24061,N_23497,N_23680);
nor U24062 (N_24062,N_23216,N_23382);
or U24063 (N_24063,N_23378,N_23431);
or U24064 (N_24064,N_23717,N_23525);
nand U24065 (N_24065,N_23399,N_23393);
or U24066 (N_24066,N_23603,N_23260);
xor U24067 (N_24067,N_23373,N_23403);
nand U24068 (N_24068,N_23505,N_23623);
nor U24069 (N_24069,N_23450,N_23558);
and U24070 (N_24070,N_23496,N_23655);
and U24071 (N_24071,N_23736,N_23275);
or U24072 (N_24072,N_23666,N_23589);
nor U24073 (N_24073,N_23637,N_23585);
and U24074 (N_24074,N_23231,N_23749);
and U24075 (N_24075,N_23351,N_23217);
and U24076 (N_24076,N_23226,N_23352);
nand U24077 (N_24077,N_23327,N_23264);
nor U24078 (N_24078,N_23233,N_23387);
nor U24079 (N_24079,N_23630,N_23327);
nand U24080 (N_24080,N_23602,N_23254);
or U24081 (N_24081,N_23734,N_23534);
nand U24082 (N_24082,N_23626,N_23689);
and U24083 (N_24083,N_23538,N_23658);
and U24084 (N_24084,N_23736,N_23185);
nor U24085 (N_24085,N_23285,N_23198);
or U24086 (N_24086,N_23166,N_23459);
nor U24087 (N_24087,N_23355,N_23126);
nor U24088 (N_24088,N_23698,N_23354);
nor U24089 (N_24089,N_23748,N_23258);
nand U24090 (N_24090,N_23443,N_23562);
or U24091 (N_24091,N_23287,N_23632);
nor U24092 (N_24092,N_23270,N_23513);
or U24093 (N_24093,N_23178,N_23651);
or U24094 (N_24094,N_23373,N_23270);
or U24095 (N_24095,N_23706,N_23601);
nand U24096 (N_24096,N_23492,N_23160);
nand U24097 (N_24097,N_23546,N_23186);
nand U24098 (N_24098,N_23517,N_23732);
and U24099 (N_24099,N_23665,N_23277);
xor U24100 (N_24100,N_23437,N_23469);
nand U24101 (N_24101,N_23341,N_23747);
nand U24102 (N_24102,N_23547,N_23308);
nor U24103 (N_24103,N_23236,N_23417);
nor U24104 (N_24104,N_23411,N_23540);
nor U24105 (N_24105,N_23211,N_23705);
xnor U24106 (N_24106,N_23657,N_23299);
nor U24107 (N_24107,N_23551,N_23614);
and U24108 (N_24108,N_23632,N_23733);
and U24109 (N_24109,N_23184,N_23612);
and U24110 (N_24110,N_23243,N_23601);
nand U24111 (N_24111,N_23242,N_23596);
nor U24112 (N_24112,N_23182,N_23595);
nand U24113 (N_24113,N_23679,N_23739);
or U24114 (N_24114,N_23335,N_23130);
and U24115 (N_24115,N_23315,N_23338);
and U24116 (N_24116,N_23526,N_23213);
or U24117 (N_24117,N_23634,N_23624);
or U24118 (N_24118,N_23477,N_23137);
or U24119 (N_24119,N_23732,N_23583);
nor U24120 (N_24120,N_23174,N_23144);
xnor U24121 (N_24121,N_23604,N_23173);
xor U24122 (N_24122,N_23307,N_23496);
nor U24123 (N_24123,N_23197,N_23383);
nor U24124 (N_24124,N_23381,N_23327);
xnor U24125 (N_24125,N_23609,N_23346);
nand U24126 (N_24126,N_23345,N_23716);
and U24127 (N_24127,N_23467,N_23638);
or U24128 (N_24128,N_23420,N_23156);
nand U24129 (N_24129,N_23479,N_23295);
and U24130 (N_24130,N_23666,N_23623);
nor U24131 (N_24131,N_23231,N_23310);
nand U24132 (N_24132,N_23604,N_23722);
and U24133 (N_24133,N_23328,N_23133);
nor U24134 (N_24134,N_23136,N_23264);
nor U24135 (N_24135,N_23500,N_23724);
and U24136 (N_24136,N_23726,N_23205);
nand U24137 (N_24137,N_23544,N_23199);
or U24138 (N_24138,N_23518,N_23486);
nor U24139 (N_24139,N_23393,N_23162);
nor U24140 (N_24140,N_23461,N_23274);
nor U24141 (N_24141,N_23457,N_23532);
nor U24142 (N_24142,N_23714,N_23646);
xnor U24143 (N_24143,N_23685,N_23245);
nor U24144 (N_24144,N_23401,N_23450);
and U24145 (N_24145,N_23708,N_23164);
or U24146 (N_24146,N_23353,N_23559);
and U24147 (N_24147,N_23292,N_23441);
nor U24148 (N_24148,N_23630,N_23610);
nor U24149 (N_24149,N_23720,N_23680);
nand U24150 (N_24150,N_23412,N_23172);
or U24151 (N_24151,N_23213,N_23429);
or U24152 (N_24152,N_23685,N_23363);
and U24153 (N_24153,N_23135,N_23507);
or U24154 (N_24154,N_23324,N_23495);
xnor U24155 (N_24155,N_23568,N_23405);
xor U24156 (N_24156,N_23661,N_23383);
nor U24157 (N_24157,N_23541,N_23712);
or U24158 (N_24158,N_23412,N_23707);
nor U24159 (N_24159,N_23619,N_23724);
and U24160 (N_24160,N_23589,N_23582);
xor U24161 (N_24161,N_23143,N_23271);
and U24162 (N_24162,N_23580,N_23284);
or U24163 (N_24163,N_23560,N_23188);
nor U24164 (N_24164,N_23237,N_23196);
or U24165 (N_24165,N_23145,N_23216);
nand U24166 (N_24166,N_23365,N_23532);
or U24167 (N_24167,N_23669,N_23379);
nor U24168 (N_24168,N_23390,N_23543);
nor U24169 (N_24169,N_23154,N_23466);
xor U24170 (N_24170,N_23220,N_23213);
nand U24171 (N_24171,N_23162,N_23358);
xor U24172 (N_24172,N_23544,N_23135);
or U24173 (N_24173,N_23229,N_23285);
xnor U24174 (N_24174,N_23303,N_23145);
nand U24175 (N_24175,N_23298,N_23313);
or U24176 (N_24176,N_23620,N_23659);
nor U24177 (N_24177,N_23276,N_23242);
nand U24178 (N_24178,N_23162,N_23578);
and U24179 (N_24179,N_23491,N_23229);
nand U24180 (N_24180,N_23172,N_23265);
nand U24181 (N_24181,N_23137,N_23218);
and U24182 (N_24182,N_23281,N_23286);
and U24183 (N_24183,N_23193,N_23531);
xor U24184 (N_24184,N_23679,N_23295);
xnor U24185 (N_24185,N_23296,N_23651);
and U24186 (N_24186,N_23217,N_23683);
nor U24187 (N_24187,N_23533,N_23662);
nand U24188 (N_24188,N_23136,N_23413);
nor U24189 (N_24189,N_23710,N_23146);
nand U24190 (N_24190,N_23190,N_23209);
and U24191 (N_24191,N_23588,N_23276);
nor U24192 (N_24192,N_23729,N_23163);
and U24193 (N_24193,N_23441,N_23479);
nand U24194 (N_24194,N_23643,N_23199);
nand U24195 (N_24195,N_23446,N_23211);
nand U24196 (N_24196,N_23701,N_23480);
or U24197 (N_24197,N_23270,N_23336);
nor U24198 (N_24198,N_23582,N_23623);
nor U24199 (N_24199,N_23368,N_23466);
or U24200 (N_24200,N_23194,N_23211);
or U24201 (N_24201,N_23307,N_23144);
nor U24202 (N_24202,N_23468,N_23301);
nand U24203 (N_24203,N_23154,N_23583);
nor U24204 (N_24204,N_23212,N_23740);
nor U24205 (N_24205,N_23489,N_23601);
nor U24206 (N_24206,N_23670,N_23423);
nor U24207 (N_24207,N_23470,N_23549);
nor U24208 (N_24208,N_23645,N_23434);
nand U24209 (N_24209,N_23548,N_23166);
nor U24210 (N_24210,N_23369,N_23169);
or U24211 (N_24211,N_23671,N_23276);
nand U24212 (N_24212,N_23169,N_23358);
or U24213 (N_24213,N_23719,N_23299);
or U24214 (N_24214,N_23327,N_23366);
or U24215 (N_24215,N_23352,N_23659);
and U24216 (N_24216,N_23607,N_23416);
nor U24217 (N_24217,N_23346,N_23348);
and U24218 (N_24218,N_23353,N_23329);
nor U24219 (N_24219,N_23670,N_23208);
and U24220 (N_24220,N_23552,N_23578);
nor U24221 (N_24221,N_23359,N_23182);
xor U24222 (N_24222,N_23465,N_23405);
nand U24223 (N_24223,N_23187,N_23499);
nor U24224 (N_24224,N_23549,N_23151);
or U24225 (N_24225,N_23201,N_23164);
and U24226 (N_24226,N_23468,N_23306);
or U24227 (N_24227,N_23630,N_23523);
nand U24228 (N_24228,N_23125,N_23631);
and U24229 (N_24229,N_23517,N_23136);
and U24230 (N_24230,N_23636,N_23380);
nand U24231 (N_24231,N_23373,N_23157);
xnor U24232 (N_24232,N_23721,N_23345);
nand U24233 (N_24233,N_23659,N_23361);
nor U24234 (N_24234,N_23561,N_23644);
and U24235 (N_24235,N_23617,N_23163);
or U24236 (N_24236,N_23533,N_23453);
nor U24237 (N_24237,N_23271,N_23393);
and U24238 (N_24238,N_23127,N_23427);
nand U24239 (N_24239,N_23519,N_23732);
nand U24240 (N_24240,N_23479,N_23579);
and U24241 (N_24241,N_23661,N_23655);
nand U24242 (N_24242,N_23382,N_23208);
and U24243 (N_24243,N_23300,N_23531);
and U24244 (N_24244,N_23454,N_23219);
and U24245 (N_24245,N_23459,N_23549);
nand U24246 (N_24246,N_23342,N_23712);
and U24247 (N_24247,N_23530,N_23619);
nand U24248 (N_24248,N_23390,N_23635);
and U24249 (N_24249,N_23139,N_23179);
and U24250 (N_24250,N_23580,N_23151);
nor U24251 (N_24251,N_23126,N_23602);
and U24252 (N_24252,N_23152,N_23281);
nand U24253 (N_24253,N_23536,N_23587);
or U24254 (N_24254,N_23334,N_23496);
or U24255 (N_24255,N_23677,N_23380);
nor U24256 (N_24256,N_23627,N_23521);
nor U24257 (N_24257,N_23254,N_23235);
nand U24258 (N_24258,N_23329,N_23161);
or U24259 (N_24259,N_23452,N_23611);
nand U24260 (N_24260,N_23384,N_23433);
nor U24261 (N_24261,N_23326,N_23295);
nand U24262 (N_24262,N_23653,N_23435);
nand U24263 (N_24263,N_23618,N_23336);
or U24264 (N_24264,N_23734,N_23287);
or U24265 (N_24265,N_23268,N_23736);
and U24266 (N_24266,N_23225,N_23581);
nand U24267 (N_24267,N_23715,N_23573);
or U24268 (N_24268,N_23711,N_23141);
or U24269 (N_24269,N_23264,N_23402);
nor U24270 (N_24270,N_23330,N_23530);
and U24271 (N_24271,N_23350,N_23180);
nand U24272 (N_24272,N_23462,N_23666);
nor U24273 (N_24273,N_23137,N_23334);
nor U24274 (N_24274,N_23448,N_23486);
or U24275 (N_24275,N_23245,N_23144);
nor U24276 (N_24276,N_23270,N_23633);
nor U24277 (N_24277,N_23709,N_23241);
nor U24278 (N_24278,N_23268,N_23545);
or U24279 (N_24279,N_23476,N_23555);
and U24280 (N_24280,N_23589,N_23145);
and U24281 (N_24281,N_23258,N_23266);
or U24282 (N_24282,N_23341,N_23322);
and U24283 (N_24283,N_23703,N_23150);
nor U24284 (N_24284,N_23157,N_23479);
xnor U24285 (N_24285,N_23154,N_23215);
and U24286 (N_24286,N_23152,N_23713);
nand U24287 (N_24287,N_23163,N_23321);
nor U24288 (N_24288,N_23158,N_23333);
and U24289 (N_24289,N_23132,N_23724);
nor U24290 (N_24290,N_23563,N_23648);
nor U24291 (N_24291,N_23453,N_23438);
nor U24292 (N_24292,N_23571,N_23727);
or U24293 (N_24293,N_23270,N_23718);
xor U24294 (N_24294,N_23417,N_23391);
nor U24295 (N_24295,N_23542,N_23338);
nor U24296 (N_24296,N_23695,N_23190);
and U24297 (N_24297,N_23430,N_23137);
or U24298 (N_24298,N_23129,N_23246);
and U24299 (N_24299,N_23511,N_23603);
nor U24300 (N_24300,N_23145,N_23299);
or U24301 (N_24301,N_23421,N_23344);
xnor U24302 (N_24302,N_23602,N_23354);
nand U24303 (N_24303,N_23224,N_23140);
or U24304 (N_24304,N_23485,N_23433);
or U24305 (N_24305,N_23160,N_23525);
nand U24306 (N_24306,N_23706,N_23699);
nand U24307 (N_24307,N_23541,N_23206);
and U24308 (N_24308,N_23659,N_23359);
and U24309 (N_24309,N_23594,N_23184);
or U24310 (N_24310,N_23125,N_23707);
and U24311 (N_24311,N_23140,N_23476);
nor U24312 (N_24312,N_23506,N_23308);
nor U24313 (N_24313,N_23361,N_23609);
nor U24314 (N_24314,N_23465,N_23311);
nor U24315 (N_24315,N_23484,N_23517);
and U24316 (N_24316,N_23749,N_23615);
nand U24317 (N_24317,N_23528,N_23641);
and U24318 (N_24318,N_23415,N_23361);
or U24319 (N_24319,N_23533,N_23288);
and U24320 (N_24320,N_23215,N_23143);
and U24321 (N_24321,N_23615,N_23715);
and U24322 (N_24322,N_23405,N_23349);
and U24323 (N_24323,N_23563,N_23384);
nand U24324 (N_24324,N_23381,N_23333);
and U24325 (N_24325,N_23235,N_23156);
or U24326 (N_24326,N_23293,N_23333);
and U24327 (N_24327,N_23138,N_23387);
and U24328 (N_24328,N_23412,N_23324);
nand U24329 (N_24329,N_23273,N_23420);
nand U24330 (N_24330,N_23712,N_23698);
or U24331 (N_24331,N_23419,N_23645);
or U24332 (N_24332,N_23698,N_23587);
nor U24333 (N_24333,N_23588,N_23422);
nand U24334 (N_24334,N_23374,N_23282);
nor U24335 (N_24335,N_23529,N_23254);
nand U24336 (N_24336,N_23135,N_23384);
nand U24337 (N_24337,N_23549,N_23734);
nor U24338 (N_24338,N_23638,N_23385);
nand U24339 (N_24339,N_23730,N_23269);
nand U24340 (N_24340,N_23310,N_23505);
nor U24341 (N_24341,N_23619,N_23277);
nor U24342 (N_24342,N_23616,N_23299);
nor U24343 (N_24343,N_23302,N_23184);
and U24344 (N_24344,N_23603,N_23195);
xnor U24345 (N_24345,N_23335,N_23569);
xor U24346 (N_24346,N_23741,N_23252);
nor U24347 (N_24347,N_23445,N_23349);
nor U24348 (N_24348,N_23710,N_23438);
nor U24349 (N_24349,N_23231,N_23479);
and U24350 (N_24350,N_23608,N_23493);
nand U24351 (N_24351,N_23671,N_23727);
and U24352 (N_24352,N_23624,N_23725);
and U24353 (N_24353,N_23316,N_23265);
and U24354 (N_24354,N_23434,N_23547);
nand U24355 (N_24355,N_23432,N_23735);
nor U24356 (N_24356,N_23673,N_23691);
or U24357 (N_24357,N_23482,N_23315);
nand U24358 (N_24358,N_23685,N_23456);
nand U24359 (N_24359,N_23316,N_23502);
xor U24360 (N_24360,N_23419,N_23344);
nor U24361 (N_24361,N_23634,N_23348);
nor U24362 (N_24362,N_23541,N_23703);
and U24363 (N_24363,N_23531,N_23729);
and U24364 (N_24364,N_23622,N_23509);
nand U24365 (N_24365,N_23301,N_23184);
nor U24366 (N_24366,N_23439,N_23225);
nand U24367 (N_24367,N_23304,N_23681);
or U24368 (N_24368,N_23598,N_23566);
and U24369 (N_24369,N_23740,N_23520);
and U24370 (N_24370,N_23183,N_23330);
and U24371 (N_24371,N_23735,N_23144);
or U24372 (N_24372,N_23640,N_23151);
or U24373 (N_24373,N_23230,N_23653);
nor U24374 (N_24374,N_23196,N_23696);
nor U24375 (N_24375,N_24038,N_23980);
or U24376 (N_24376,N_24051,N_24317);
nor U24377 (N_24377,N_24031,N_24015);
nor U24378 (N_24378,N_24194,N_24359);
or U24379 (N_24379,N_24082,N_24237);
and U24380 (N_24380,N_24132,N_24252);
xnor U24381 (N_24381,N_23913,N_24049);
nand U24382 (N_24382,N_23796,N_23857);
nor U24383 (N_24383,N_23903,N_23832);
nand U24384 (N_24384,N_23861,N_24297);
nor U24385 (N_24385,N_23917,N_24060);
nand U24386 (N_24386,N_23815,N_24287);
xnor U24387 (N_24387,N_24222,N_24165);
or U24388 (N_24388,N_24105,N_24032);
and U24389 (N_24389,N_24339,N_24346);
nor U24390 (N_24390,N_23873,N_24184);
or U24391 (N_24391,N_24009,N_24335);
nand U24392 (N_24392,N_24199,N_23764);
and U24393 (N_24393,N_23817,N_24083);
nand U24394 (N_24394,N_24182,N_24154);
or U24395 (N_24395,N_23860,N_24330);
nor U24396 (N_24396,N_23943,N_24073);
nand U24397 (N_24397,N_24269,N_23887);
or U24398 (N_24398,N_23897,N_24300);
and U24399 (N_24399,N_23834,N_24155);
and U24400 (N_24400,N_23852,N_23811);
nand U24401 (N_24401,N_23894,N_23848);
and U24402 (N_24402,N_24058,N_24217);
and U24403 (N_24403,N_23807,N_24246);
and U24404 (N_24404,N_24340,N_24245);
nor U24405 (N_24405,N_23843,N_23778);
nand U24406 (N_24406,N_23877,N_23761);
and U24407 (N_24407,N_24003,N_24100);
or U24408 (N_24408,N_23758,N_23909);
and U24409 (N_24409,N_24183,N_24069);
or U24410 (N_24410,N_24364,N_23823);
and U24411 (N_24411,N_24004,N_24224);
and U24412 (N_24412,N_24355,N_24232);
and U24413 (N_24413,N_24257,N_23846);
or U24414 (N_24414,N_23774,N_23939);
and U24415 (N_24415,N_23979,N_23889);
nor U24416 (N_24416,N_24170,N_24005);
nor U24417 (N_24417,N_24316,N_24039);
nor U24418 (N_24418,N_24333,N_24261);
nand U24419 (N_24419,N_24278,N_23930);
and U24420 (N_24420,N_24077,N_24197);
xnor U24421 (N_24421,N_24080,N_24162);
or U24422 (N_24422,N_23773,N_24268);
xnor U24423 (N_24423,N_24271,N_24090);
or U24424 (N_24424,N_23858,N_24305);
nand U24425 (N_24425,N_24334,N_24052);
or U24426 (N_24426,N_24117,N_23756);
nand U24427 (N_24427,N_23967,N_24088);
nand U24428 (N_24428,N_23993,N_23997);
nor U24429 (N_24429,N_24275,N_23986);
nor U24430 (N_24430,N_24153,N_23779);
and U24431 (N_24431,N_23760,N_23931);
nor U24432 (N_24432,N_24327,N_24023);
xnor U24433 (N_24433,N_24281,N_24322);
nand U24434 (N_24434,N_23914,N_23870);
and U24435 (N_24435,N_24181,N_23900);
and U24436 (N_24436,N_24091,N_23780);
xor U24437 (N_24437,N_24021,N_23942);
nor U24438 (N_24438,N_24228,N_23782);
xnor U24439 (N_24439,N_23927,N_23835);
nand U24440 (N_24440,N_23820,N_24213);
xnor U24441 (N_24441,N_24185,N_24172);
nand U24442 (N_24442,N_23824,N_23847);
nand U24443 (N_24443,N_24121,N_23786);
xnor U24444 (N_24444,N_23803,N_23766);
nand U24445 (N_24445,N_23819,N_24012);
nand U24446 (N_24446,N_23798,N_24027);
xnor U24447 (N_24447,N_24212,N_24141);
and U24448 (N_24448,N_24247,N_24156);
xor U24449 (N_24449,N_24095,N_24353);
or U24450 (N_24450,N_24298,N_24304);
nand U24451 (N_24451,N_24243,N_24289);
nand U24452 (N_24452,N_24351,N_24253);
or U24453 (N_24453,N_24215,N_23789);
nor U24454 (N_24454,N_24010,N_23921);
and U24455 (N_24455,N_24089,N_24230);
nor U24456 (N_24456,N_23985,N_24254);
and U24457 (N_24457,N_23959,N_24323);
nand U24458 (N_24458,N_24071,N_23783);
or U24459 (N_24459,N_24102,N_24244);
nand U24460 (N_24460,N_24349,N_24180);
nor U24461 (N_24461,N_24099,N_24129);
xnor U24462 (N_24462,N_24219,N_24079);
or U24463 (N_24463,N_24277,N_23935);
and U24464 (N_24464,N_23953,N_24249);
and U24465 (N_24465,N_24081,N_24190);
or U24466 (N_24466,N_23987,N_24104);
nand U24467 (N_24467,N_23941,N_23904);
nor U24468 (N_24468,N_23973,N_24065);
and U24469 (N_24469,N_24362,N_23944);
or U24470 (N_24470,N_24200,N_23795);
nor U24471 (N_24471,N_24036,N_24033);
and U24472 (N_24472,N_24087,N_24236);
xor U24473 (N_24473,N_23864,N_23755);
or U24474 (N_24474,N_24177,N_24028);
nand U24475 (N_24475,N_24035,N_24341);
and U24476 (N_24476,N_23933,N_24358);
and U24477 (N_24477,N_23814,N_23912);
or U24478 (N_24478,N_24143,N_24186);
or U24479 (N_24479,N_23837,N_24319);
nor U24480 (N_24480,N_24315,N_23785);
xor U24481 (N_24481,N_23853,N_24365);
xnor U24482 (N_24482,N_24054,N_23911);
or U24483 (N_24483,N_23775,N_23996);
nor U24484 (N_24484,N_24285,N_23830);
and U24485 (N_24485,N_24343,N_24210);
or U24486 (N_24486,N_24361,N_24125);
and U24487 (N_24487,N_23949,N_23876);
and U24488 (N_24488,N_24013,N_24274);
or U24489 (N_24489,N_24115,N_24167);
and U24490 (N_24490,N_24324,N_23884);
and U24491 (N_24491,N_23809,N_24356);
or U24492 (N_24492,N_24188,N_23866);
or U24493 (N_24493,N_23763,N_24290);
or U24494 (N_24494,N_23910,N_24112);
and U24495 (N_24495,N_24189,N_24096);
or U24496 (N_24496,N_24286,N_23802);
or U24497 (N_24497,N_24279,N_24270);
nand U24498 (N_24498,N_24347,N_24329);
nor U24499 (N_24499,N_24331,N_23862);
or U24500 (N_24500,N_24136,N_23799);
or U24501 (N_24501,N_24223,N_23883);
nand U24502 (N_24502,N_24256,N_24007);
and U24503 (N_24503,N_24248,N_23998);
and U24504 (N_24504,N_23836,N_23947);
or U24505 (N_24505,N_24152,N_24016);
and U24506 (N_24506,N_24166,N_24160);
nand U24507 (N_24507,N_24229,N_24370);
and U24508 (N_24508,N_23788,N_23869);
nor U24509 (N_24509,N_23838,N_24344);
or U24510 (N_24510,N_23984,N_23962);
nor U24511 (N_24511,N_24137,N_23922);
or U24512 (N_24512,N_23964,N_23898);
or U24513 (N_24513,N_23994,N_23988);
nor U24514 (N_24514,N_24225,N_23963);
nand U24515 (N_24515,N_23951,N_23833);
nand U24516 (N_24516,N_24325,N_24231);
or U24517 (N_24517,N_24306,N_23906);
or U24518 (N_24518,N_24118,N_24050);
xor U24519 (N_24519,N_23825,N_24303);
or U24520 (N_24520,N_24158,N_24207);
and U24521 (N_24521,N_24284,N_24126);
nor U24522 (N_24522,N_23874,N_23981);
or U24523 (N_24523,N_24000,N_24368);
or U24524 (N_24524,N_24187,N_23810);
and U24525 (N_24525,N_24057,N_23916);
and U24526 (N_24526,N_24174,N_23793);
and U24527 (N_24527,N_23970,N_24101);
and U24528 (N_24528,N_24134,N_24116);
nor U24529 (N_24529,N_24250,N_24046);
or U24530 (N_24530,N_23851,N_23950);
and U24531 (N_24531,N_23940,N_24374);
xnor U24532 (N_24532,N_23938,N_23752);
or U24533 (N_24533,N_23865,N_24075);
or U24534 (N_24534,N_23875,N_23850);
or U24535 (N_24535,N_24241,N_24056);
nor U24536 (N_24536,N_24321,N_23845);
nor U24537 (N_24537,N_24192,N_23977);
and U24538 (N_24538,N_23965,N_23954);
or U24539 (N_24539,N_23829,N_24045);
or U24540 (N_24540,N_23777,N_24150);
nand U24541 (N_24541,N_23902,N_23975);
nand U24542 (N_24542,N_23881,N_24017);
nand U24543 (N_24543,N_23856,N_23831);
nand U24544 (N_24544,N_24266,N_23983);
and U24545 (N_24545,N_24074,N_24064);
or U24546 (N_24546,N_23957,N_24363);
nand U24547 (N_24547,N_23772,N_24264);
xor U24548 (N_24548,N_24119,N_24086);
nand U24549 (N_24549,N_24204,N_24318);
or U24550 (N_24550,N_24366,N_24265);
nor U24551 (N_24551,N_24313,N_24020);
or U24552 (N_24552,N_24288,N_23936);
nand U24553 (N_24553,N_24085,N_24221);
or U24554 (N_24554,N_24048,N_24320);
nor U24555 (N_24555,N_23885,N_23867);
nand U24556 (N_24556,N_23968,N_24336);
nand U24557 (N_24557,N_24067,N_23892);
and U24558 (N_24558,N_23769,N_24131);
nand U24559 (N_24559,N_23839,N_24171);
nand U24560 (N_24560,N_23888,N_24201);
nand U24561 (N_24561,N_23976,N_23896);
nand U24562 (N_24562,N_23751,N_24063);
nor U24563 (N_24563,N_24114,N_24342);
nor U24564 (N_24564,N_24214,N_24337);
or U24565 (N_24565,N_23908,N_24242);
and U24566 (N_24566,N_24372,N_24299);
nand U24567 (N_24567,N_24123,N_24014);
nor U24568 (N_24568,N_23934,N_24161);
and U24569 (N_24569,N_24110,N_24084);
nor U24570 (N_24570,N_24019,N_24024);
nand U24571 (N_24571,N_24220,N_24196);
and U24572 (N_24572,N_23762,N_24163);
or U24573 (N_24573,N_24072,N_24111);
xor U24574 (N_24574,N_23805,N_24149);
and U24575 (N_24575,N_23989,N_24168);
and U24576 (N_24576,N_24272,N_23932);
or U24577 (N_24577,N_24280,N_24146);
nand U24578 (N_24578,N_24109,N_23750);
nor U24579 (N_24579,N_23859,N_23781);
nor U24580 (N_24580,N_24276,N_24178);
and U24581 (N_24581,N_24053,N_23841);
nor U24582 (N_24582,N_24002,N_23840);
xor U24583 (N_24583,N_23791,N_23828);
nand U24584 (N_24584,N_24025,N_24294);
xnor U24585 (N_24585,N_23999,N_23971);
and U24586 (N_24586,N_23816,N_24240);
nor U24587 (N_24587,N_24292,N_24120);
xnor U24588 (N_24588,N_23784,N_24176);
xor U24589 (N_24589,N_23891,N_24309);
and U24590 (N_24590,N_24147,N_24234);
nand U24591 (N_24591,N_23905,N_23868);
or U24592 (N_24592,N_23915,N_24040);
or U24593 (N_24593,N_23926,N_23826);
nor U24594 (N_24594,N_23958,N_24042);
nand U24595 (N_24595,N_24338,N_23920);
nor U24596 (N_24596,N_24206,N_23923);
nor U24597 (N_24597,N_24282,N_23879);
or U24598 (N_24598,N_24267,N_23899);
nor U24599 (N_24599,N_24259,N_24041);
or U24600 (N_24600,N_24238,N_24108);
nor U24601 (N_24601,N_23928,N_24173);
and U24602 (N_24602,N_23863,N_24037);
nor U24603 (N_24603,N_23880,N_24133);
and U24604 (N_24604,N_24357,N_24293);
nor U24605 (N_24605,N_24059,N_23907);
nor U24606 (N_24606,N_23992,N_23991);
nor U24607 (N_24607,N_24026,N_23893);
or U24608 (N_24608,N_23844,N_24062);
and U24609 (N_24609,N_24151,N_24179);
nor U24610 (N_24610,N_23800,N_24130);
xnor U24611 (N_24611,N_24233,N_23995);
nor U24612 (N_24612,N_24211,N_24097);
or U24613 (N_24613,N_23806,N_23849);
nor U24614 (N_24614,N_24312,N_23872);
or U24615 (N_24615,N_24260,N_24218);
and U24616 (N_24616,N_24070,N_24198);
or U24617 (N_24617,N_24140,N_23842);
nor U24618 (N_24618,N_23978,N_23776);
nor U24619 (N_24619,N_24227,N_23765);
nand U24620 (N_24620,N_24001,N_24209);
nor U24621 (N_24621,N_24202,N_23969);
and U24622 (N_24622,N_24191,N_23925);
xnor U24623 (N_24623,N_23787,N_24078);
nor U24624 (N_24624,N_23878,N_24008);
and U24625 (N_24625,N_24044,N_23797);
xnor U24626 (N_24626,N_24103,N_24367);
or U24627 (N_24627,N_24148,N_23767);
and U24628 (N_24628,N_24030,N_24255);
or U24629 (N_24629,N_24029,N_23945);
nor U24630 (N_24630,N_24142,N_24226);
nor U24631 (N_24631,N_23818,N_24128);
nand U24632 (N_24632,N_24308,N_24135);
or U24633 (N_24633,N_24157,N_24076);
nor U24634 (N_24634,N_23768,N_24068);
nor U24635 (N_24635,N_24360,N_23801);
xor U24636 (N_24636,N_23753,N_24113);
nor U24637 (N_24637,N_23946,N_23961);
and U24638 (N_24638,N_24159,N_23808);
xor U24639 (N_24639,N_24175,N_24273);
and U24640 (N_24640,N_23890,N_23794);
and U24641 (N_24641,N_24043,N_23822);
nor U24642 (N_24642,N_24066,N_23972);
and U24643 (N_24643,N_23919,N_24018);
nor U24644 (N_24644,N_23960,N_24034);
and U24645 (N_24645,N_24369,N_23770);
nor U24646 (N_24646,N_23918,N_23882);
and U24647 (N_24647,N_24195,N_24055);
and U24648 (N_24648,N_24314,N_24203);
nor U24649 (N_24649,N_23955,N_23937);
or U24650 (N_24650,N_24345,N_24022);
or U24651 (N_24651,N_24006,N_23854);
nor U24652 (N_24652,N_24124,N_24350);
nand U24653 (N_24653,N_24326,N_24296);
nor U24654 (N_24654,N_24169,N_23792);
or U24655 (N_24655,N_23974,N_24307);
nor U24656 (N_24656,N_23827,N_23929);
and U24657 (N_24657,N_24235,N_24371);
nor U24658 (N_24658,N_23790,N_24144);
or U24659 (N_24659,N_24258,N_24092);
and U24660 (N_24660,N_23771,N_24216);
xor U24661 (N_24661,N_24283,N_23757);
nand U24662 (N_24662,N_23813,N_24193);
xnor U24663 (N_24663,N_24047,N_23821);
nor U24664 (N_24664,N_24352,N_24164);
and U24665 (N_24665,N_23871,N_24208);
or U24666 (N_24666,N_23895,N_24106);
nor U24667 (N_24667,N_24310,N_24094);
and U24668 (N_24668,N_24011,N_23855);
or U24669 (N_24669,N_23754,N_23924);
or U24670 (N_24670,N_24122,N_24373);
nor U24671 (N_24671,N_23759,N_24311);
nor U24672 (N_24672,N_24262,N_23966);
or U24673 (N_24673,N_23952,N_23982);
and U24674 (N_24674,N_24328,N_24145);
or U24675 (N_24675,N_24138,N_23990);
or U24676 (N_24676,N_23812,N_24107);
or U24677 (N_24677,N_24301,N_24098);
nor U24678 (N_24678,N_24251,N_24302);
and U24679 (N_24679,N_24139,N_24348);
or U24680 (N_24680,N_24239,N_24295);
nand U24681 (N_24681,N_24127,N_24291);
xor U24682 (N_24682,N_23948,N_24263);
and U24683 (N_24683,N_23956,N_24061);
nand U24684 (N_24684,N_24205,N_23886);
xor U24685 (N_24685,N_23804,N_24332);
nand U24686 (N_24686,N_24093,N_24354);
nor U24687 (N_24687,N_23901,N_24326);
or U24688 (N_24688,N_23892,N_24200);
and U24689 (N_24689,N_23980,N_23918);
nor U24690 (N_24690,N_24367,N_24160);
xor U24691 (N_24691,N_24186,N_23855);
nand U24692 (N_24692,N_24132,N_24035);
or U24693 (N_24693,N_23789,N_24045);
or U24694 (N_24694,N_24141,N_24299);
and U24695 (N_24695,N_24173,N_24327);
nor U24696 (N_24696,N_23933,N_23900);
or U24697 (N_24697,N_24259,N_24004);
and U24698 (N_24698,N_23902,N_24366);
nor U24699 (N_24699,N_23921,N_24350);
or U24700 (N_24700,N_23919,N_24355);
or U24701 (N_24701,N_23751,N_23930);
nand U24702 (N_24702,N_23956,N_24330);
nand U24703 (N_24703,N_23991,N_24213);
nand U24704 (N_24704,N_24256,N_23854);
xnor U24705 (N_24705,N_23868,N_24151);
nand U24706 (N_24706,N_24187,N_24083);
nand U24707 (N_24707,N_24269,N_23781);
xor U24708 (N_24708,N_24034,N_24271);
nor U24709 (N_24709,N_23941,N_24164);
nand U24710 (N_24710,N_23931,N_24304);
or U24711 (N_24711,N_24016,N_23932);
nand U24712 (N_24712,N_24170,N_24211);
nor U24713 (N_24713,N_24175,N_24002);
or U24714 (N_24714,N_24238,N_24150);
nor U24715 (N_24715,N_23837,N_23820);
and U24716 (N_24716,N_24337,N_23874);
and U24717 (N_24717,N_23803,N_24240);
or U24718 (N_24718,N_24137,N_24190);
xor U24719 (N_24719,N_23936,N_24107);
xor U24720 (N_24720,N_23887,N_24046);
nand U24721 (N_24721,N_23987,N_24189);
and U24722 (N_24722,N_24134,N_24104);
or U24723 (N_24723,N_24169,N_24277);
or U24724 (N_24724,N_24177,N_23863);
nand U24725 (N_24725,N_24298,N_23856);
nor U24726 (N_24726,N_23767,N_24120);
and U24727 (N_24727,N_24152,N_24162);
and U24728 (N_24728,N_24271,N_24316);
nor U24729 (N_24729,N_23822,N_24065);
or U24730 (N_24730,N_23763,N_23961);
nand U24731 (N_24731,N_24192,N_24221);
or U24732 (N_24732,N_23880,N_24156);
and U24733 (N_24733,N_24001,N_24003);
or U24734 (N_24734,N_24138,N_23971);
nand U24735 (N_24735,N_23883,N_24211);
nor U24736 (N_24736,N_24295,N_24315);
nand U24737 (N_24737,N_24367,N_23879);
nand U24738 (N_24738,N_24100,N_24029);
and U24739 (N_24739,N_23908,N_24287);
nand U24740 (N_24740,N_24235,N_23921);
and U24741 (N_24741,N_24307,N_24160);
nand U24742 (N_24742,N_23844,N_24287);
xor U24743 (N_24743,N_23900,N_24258);
and U24744 (N_24744,N_23752,N_24248);
or U24745 (N_24745,N_24012,N_23768);
nor U24746 (N_24746,N_23797,N_24232);
or U24747 (N_24747,N_24301,N_23945);
nand U24748 (N_24748,N_23904,N_23936);
or U24749 (N_24749,N_24110,N_23834);
nand U24750 (N_24750,N_24243,N_24275);
xor U24751 (N_24751,N_24242,N_24298);
or U24752 (N_24752,N_23751,N_23912);
nor U24753 (N_24753,N_24335,N_24197);
nand U24754 (N_24754,N_24114,N_24065);
nor U24755 (N_24755,N_24140,N_24076);
xnor U24756 (N_24756,N_24172,N_23930);
and U24757 (N_24757,N_23955,N_24372);
and U24758 (N_24758,N_23757,N_23909);
nor U24759 (N_24759,N_23916,N_23946);
or U24760 (N_24760,N_24221,N_24158);
nand U24761 (N_24761,N_24216,N_23928);
and U24762 (N_24762,N_24322,N_23992);
nand U24763 (N_24763,N_23774,N_24373);
and U24764 (N_24764,N_24236,N_24021);
xor U24765 (N_24765,N_23847,N_23851);
nand U24766 (N_24766,N_24095,N_23996);
nand U24767 (N_24767,N_24187,N_24367);
and U24768 (N_24768,N_23926,N_24340);
nand U24769 (N_24769,N_24290,N_24024);
nor U24770 (N_24770,N_23944,N_24269);
and U24771 (N_24771,N_24359,N_23781);
and U24772 (N_24772,N_24164,N_24191);
or U24773 (N_24773,N_24286,N_24045);
and U24774 (N_24774,N_24278,N_23819);
nor U24775 (N_24775,N_23993,N_23985);
nand U24776 (N_24776,N_24347,N_24281);
nor U24777 (N_24777,N_24263,N_24328);
nand U24778 (N_24778,N_24373,N_23929);
nor U24779 (N_24779,N_23857,N_24326);
or U24780 (N_24780,N_23788,N_24308);
and U24781 (N_24781,N_23761,N_24171);
or U24782 (N_24782,N_24153,N_23803);
and U24783 (N_24783,N_23935,N_23857);
and U24784 (N_24784,N_24003,N_24301);
nor U24785 (N_24785,N_24283,N_23765);
nor U24786 (N_24786,N_23953,N_23969);
nand U24787 (N_24787,N_23973,N_24072);
and U24788 (N_24788,N_23885,N_23760);
nand U24789 (N_24789,N_24015,N_24270);
nor U24790 (N_24790,N_23918,N_23894);
xor U24791 (N_24791,N_24286,N_24330);
nor U24792 (N_24792,N_23825,N_24046);
and U24793 (N_24793,N_24018,N_24059);
or U24794 (N_24794,N_24345,N_23992);
nor U24795 (N_24795,N_23925,N_24027);
nand U24796 (N_24796,N_24283,N_24188);
or U24797 (N_24797,N_24365,N_23999);
xnor U24798 (N_24798,N_23791,N_23849);
nand U24799 (N_24799,N_23856,N_24367);
nand U24800 (N_24800,N_23903,N_23870);
nand U24801 (N_24801,N_23830,N_23865);
and U24802 (N_24802,N_24319,N_23787);
or U24803 (N_24803,N_24372,N_23813);
nor U24804 (N_24804,N_23894,N_23866);
or U24805 (N_24805,N_24074,N_24263);
or U24806 (N_24806,N_23858,N_24017);
and U24807 (N_24807,N_24056,N_23762);
and U24808 (N_24808,N_23999,N_24336);
xor U24809 (N_24809,N_24186,N_24013);
nand U24810 (N_24810,N_24238,N_24070);
xor U24811 (N_24811,N_24040,N_24334);
and U24812 (N_24812,N_24092,N_24362);
nor U24813 (N_24813,N_23942,N_23785);
nor U24814 (N_24814,N_24001,N_24091);
nand U24815 (N_24815,N_24275,N_24064);
and U24816 (N_24816,N_23918,N_23784);
and U24817 (N_24817,N_23961,N_23785);
nor U24818 (N_24818,N_23760,N_24294);
xnor U24819 (N_24819,N_24284,N_23919);
or U24820 (N_24820,N_23860,N_23902);
and U24821 (N_24821,N_24042,N_24077);
nand U24822 (N_24822,N_23832,N_24302);
nor U24823 (N_24823,N_24158,N_23866);
and U24824 (N_24824,N_24109,N_23777);
or U24825 (N_24825,N_24294,N_23755);
and U24826 (N_24826,N_24254,N_23882);
nand U24827 (N_24827,N_24174,N_24295);
or U24828 (N_24828,N_23970,N_24262);
or U24829 (N_24829,N_24373,N_23869);
and U24830 (N_24830,N_24342,N_24256);
nor U24831 (N_24831,N_24120,N_24116);
nand U24832 (N_24832,N_23869,N_23813);
nand U24833 (N_24833,N_24165,N_23918);
nand U24834 (N_24834,N_24088,N_24059);
or U24835 (N_24835,N_24307,N_24242);
nand U24836 (N_24836,N_24170,N_24146);
and U24837 (N_24837,N_24228,N_23888);
and U24838 (N_24838,N_23994,N_24329);
and U24839 (N_24839,N_24225,N_23880);
or U24840 (N_24840,N_24068,N_23937);
nor U24841 (N_24841,N_24154,N_23801);
or U24842 (N_24842,N_23806,N_23870);
and U24843 (N_24843,N_24051,N_24234);
or U24844 (N_24844,N_24022,N_24083);
and U24845 (N_24845,N_24111,N_24328);
and U24846 (N_24846,N_23855,N_24037);
nor U24847 (N_24847,N_24010,N_24036);
nand U24848 (N_24848,N_24021,N_23947);
nand U24849 (N_24849,N_24108,N_24153);
and U24850 (N_24850,N_24374,N_24325);
and U24851 (N_24851,N_24163,N_24138);
nand U24852 (N_24852,N_23754,N_24217);
xnor U24853 (N_24853,N_23989,N_24236);
or U24854 (N_24854,N_23891,N_24358);
nand U24855 (N_24855,N_24174,N_23963);
nand U24856 (N_24856,N_23817,N_23982);
or U24857 (N_24857,N_24037,N_24200);
and U24858 (N_24858,N_24091,N_24112);
and U24859 (N_24859,N_24331,N_24170);
and U24860 (N_24860,N_24289,N_24188);
and U24861 (N_24861,N_24310,N_24350);
nor U24862 (N_24862,N_24352,N_23953);
nand U24863 (N_24863,N_23861,N_23999);
nand U24864 (N_24864,N_23841,N_23785);
nand U24865 (N_24865,N_23975,N_24028);
nand U24866 (N_24866,N_24187,N_24012);
and U24867 (N_24867,N_23871,N_23990);
nand U24868 (N_24868,N_24039,N_24088);
or U24869 (N_24869,N_24273,N_23977);
or U24870 (N_24870,N_24142,N_23924);
and U24871 (N_24871,N_24029,N_23893);
or U24872 (N_24872,N_23919,N_24295);
or U24873 (N_24873,N_23779,N_23937);
xor U24874 (N_24874,N_23934,N_24170);
xnor U24875 (N_24875,N_23993,N_23820);
nand U24876 (N_24876,N_24219,N_24103);
nor U24877 (N_24877,N_24185,N_24120);
nor U24878 (N_24878,N_24310,N_24165);
and U24879 (N_24879,N_23825,N_23841);
nand U24880 (N_24880,N_24304,N_24036);
nor U24881 (N_24881,N_23901,N_24286);
nor U24882 (N_24882,N_23887,N_24143);
and U24883 (N_24883,N_24192,N_24185);
nand U24884 (N_24884,N_23914,N_24155);
or U24885 (N_24885,N_24374,N_24086);
or U24886 (N_24886,N_23898,N_24212);
and U24887 (N_24887,N_23792,N_24065);
nor U24888 (N_24888,N_24339,N_23943);
xor U24889 (N_24889,N_23867,N_24047);
nand U24890 (N_24890,N_23886,N_24141);
or U24891 (N_24891,N_24251,N_24230);
or U24892 (N_24892,N_24368,N_24063);
and U24893 (N_24893,N_23837,N_24004);
nand U24894 (N_24894,N_23849,N_24075);
or U24895 (N_24895,N_23986,N_23863);
or U24896 (N_24896,N_24137,N_23820);
nand U24897 (N_24897,N_24258,N_24341);
nand U24898 (N_24898,N_24068,N_24031);
and U24899 (N_24899,N_24124,N_24198);
or U24900 (N_24900,N_24297,N_23943);
nor U24901 (N_24901,N_23962,N_24102);
nand U24902 (N_24902,N_24253,N_24042);
nand U24903 (N_24903,N_24279,N_23830);
and U24904 (N_24904,N_24057,N_24142);
nor U24905 (N_24905,N_23774,N_24229);
nand U24906 (N_24906,N_24014,N_23878);
or U24907 (N_24907,N_23816,N_24119);
xor U24908 (N_24908,N_24165,N_24364);
nand U24909 (N_24909,N_24091,N_24016);
nor U24910 (N_24910,N_24222,N_23753);
xor U24911 (N_24911,N_24348,N_23803);
and U24912 (N_24912,N_24086,N_24361);
and U24913 (N_24913,N_24189,N_23946);
and U24914 (N_24914,N_23926,N_24185);
xnor U24915 (N_24915,N_23773,N_24255);
and U24916 (N_24916,N_24281,N_24033);
nor U24917 (N_24917,N_23857,N_23838);
nand U24918 (N_24918,N_24144,N_23991);
nor U24919 (N_24919,N_24293,N_24180);
or U24920 (N_24920,N_24184,N_24082);
or U24921 (N_24921,N_23754,N_24270);
and U24922 (N_24922,N_23893,N_23873);
nor U24923 (N_24923,N_24261,N_24101);
nand U24924 (N_24924,N_24279,N_24091);
nand U24925 (N_24925,N_23974,N_24127);
nand U24926 (N_24926,N_23940,N_24136);
nor U24927 (N_24927,N_24298,N_24337);
nor U24928 (N_24928,N_24130,N_23855);
or U24929 (N_24929,N_23901,N_24275);
and U24930 (N_24930,N_24064,N_24356);
nor U24931 (N_24931,N_24026,N_24276);
xor U24932 (N_24932,N_24033,N_23834);
and U24933 (N_24933,N_24193,N_24206);
or U24934 (N_24934,N_24135,N_24235);
or U24935 (N_24935,N_24151,N_24201);
nand U24936 (N_24936,N_24110,N_23956);
and U24937 (N_24937,N_23795,N_24095);
and U24938 (N_24938,N_23942,N_24022);
nand U24939 (N_24939,N_24000,N_24317);
nor U24940 (N_24940,N_23887,N_24369);
xor U24941 (N_24941,N_24256,N_23813);
xor U24942 (N_24942,N_23991,N_24004);
or U24943 (N_24943,N_23835,N_23814);
nand U24944 (N_24944,N_24239,N_23754);
or U24945 (N_24945,N_23762,N_23808);
nor U24946 (N_24946,N_23767,N_23754);
or U24947 (N_24947,N_24122,N_24071);
nand U24948 (N_24948,N_24200,N_24204);
and U24949 (N_24949,N_24069,N_24144);
and U24950 (N_24950,N_24210,N_24140);
nor U24951 (N_24951,N_24146,N_24258);
nand U24952 (N_24952,N_24225,N_24367);
nand U24953 (N_24953,N_23821,N_24290);
or U24954 (N_24954,N_24354,N_23878);
xnor U24955 (N_24955,N_23774,N_24284);
or U24956 (N_24956,N_23999,N_24235);
or U24957 (N_24957,N_24031,N_24368);
or U24958 (N_24958,N_24233,N_23864);
or U24959 (N_24959,N_24297,N_24017);
nor U24960 (N_24960,N_24003,N_24125);
nand U24961 (N_24961,N_24070,N_23955);
and U24962 (N_24962,N_23771,N_23880);
nand U24963 (N_24963,N_24074,N_24061);
nand U24964 (N_24964,N_24288,N_23912);
and U24965 (N_24965,N_24128,N_23903);
nand U24966 (N_24966,N_23966,N_24141);
nor U24967 (N_24967,N_24223,N_23903);
nand U24968 (N_24968,N_23762,N_24032);
nor U24969 (N_24969,N_24018,N_23861);
or U24970 (N_24970,N_24364,N_23891);
nor U24971 (N_24971,N_24298,N_24002);
nor U24972 (N_24972,N_24111,N_24269);
nor U24973 (N_24973,N_23855,N_24318);
or U24974 (N_24974,N_24222,N_24321);
or U24975 (N_24975,N_23994,N_24004);
and U24976 (N_24976,N_24091,N_24023);
nor U24977 (N_24977,N_24164,N_23893);
or U24978 (N_24978,N_24197,N_24319);
and U24979 (N_24979,N_23957,N_24198);
nand U24980 (N_24980,N_24093,N_24078);
xnor U24981 (N_24981,N_24222,N_24247);
xnor U24982 (N_24982,N_24234,N_23889);
nand U24983 (N_24983,N_23959,N_24110);
xnor U24984 (N_24984,N_23926,N_24248);
nor U24985 (N_24985,N_24137,N_24142);
and U24986 (N_24986,N_24171,N_23852);
xor U24987 (N_24987,N_23913,N_24262);
nor U24988 (N_24988,N_24345,N_24202);
or U24989 (N_24989,N_24157,N_23775);
or U24990 (N_24990,N_24242,N_24174);
xnor U24991 (N_24991,N_24224,N_23979);
and U24992 (N_24992,N_24056,N_23980);
xnor U24993 (N_24993,N_24115,N_23930);
xnor U24994 (N_24994,N_23825,N_24084);
nand U24995 (N_24995,N_23834,N_24043);
nor U24996 (N_24996,N_24033,N_24172);
nor U24997 (N_24997,N_24057,N_23958);
and U24998 (N_24998,N_24186,N_23789);
nor U24999 (N_24999,N_24186,N_23850);
nand UO_0 (O_0,N_24674,N_24758);
nand UO_1 (O_1,N_24418,N_24620);
nand UO_2 (O_2,N_24527,N_24425);
nand UO_3 (O_3,N_24486,N_24537);
nand UO_4 (O_4,N_24877,N_24495);
or UO_5 (O_5,N_24848,N_24704);
or UO_6 (O_6,N_24725,N_24503);
xnor UO_7 (O_7,N_24582,N_24429);
or UO_8 (O_8,N_24903,N_24439);
nand UO_9 (O_9,N_24679,N_24424);
xor UO_10 (O_10,N_24880,N_24638);
nor UO_11 (O_11,N_24755,N_24635);
nand UO_12 (O_12,N_24502,N_24749);
nor UO_13 (O_13,N_24783,N_24383);
nand UO_14 (O_14,N_24487,N_24696);
nand UO_15 (O_15,N_24776,N_24798);
and UO_16 (O_16,N_24551,N_24957);
and UO_17 (O_17,N_24835,N_24869);
and UO_18 (O_18,N_24651,N_24691);
xor UO_19 (O_19,N_24575,N_24587);
and UO_20 (O_20,N_24452,N_24540);
and UO_21 (O_21,N_24985,N_24398);
nand UO_22 (O_22,N_24834,N_24456);
or UO_23 (O_23,N_24618,N_24397);
or UO_24 (O_24,N_24546,N_24663);
nor UO_25 (O_25,N_24440,N_24443);
nor UO_26 (O_26,N_24931,N_24402);
or UO_27 (O_27,N_24606,N_24570);
nor UO_28 (O_28,N_24925,N_24380);
and UO_29 (O_29,N_24799,N_24581);
and UO_30 (O_30,N_24464,N_24761);
nand UO_31 (O_31,N_24808,N_24775);
nand UO_32 (O_32,N_24700,N_24394);
or UO_33 (O_33,N_24555,N_24870);
and UO_34 (O_34,N_24917,N_24906);
nor UO_35 (O_35,N_24868,N_24396);
nor UO_36 (O_36,N_24384,N_24516);
nor UO_37 (O_37,N_24935,N_24554);
nand UO_38 (O_38,N_24839,N_24722);
nand UO_39 (O_39,N_24428,N_24523);
nor UO_40 (O_40,N_24403,N_24496);
or UO_41 (O_41,N_24492,N_24619);
nor UO_42 (O_42,N_24945,N_24994);
nand UO_43 (O_43,N_24934,N_24597);
nand UO_44 (O_44,N_24455,N_24735);
nand UO_45 (O_45,N_24874,N_24557);
and UO_46 (O_46,N_24784,N_24797);
nand UO_47 (O_47,N_24665,N_24416);
or UO_48 (O_48,N_24721,N_24594);
or UO_49 (O_49,N_24560,N_24435);
nor UO_50 (O_50,N_24386,N_24680);
or UO_51 (O_51,N_24658,N_24387);
or UO_52 (O_52,N_24927,N_24982);
xnor UO_53 (O_53,N_24686,N_24672);
nor UO_54 (O_54,N_24675,N_24987);
and UO_55 (O_55,N_24731,N_24623);
or UO_56 (O_56,N_24565,N_24669);
and UO_57 (O_57,N_24460,N_24611);
nor UO_58 (O_58,N_24461,N_24790);
and UO_59 (O_59,N_24437,N_24795);
xnor UO_60 (O_60,N_24643,N_24718);
and UO_61 (O_61,N_24729,N_24533);
or UO_62 (O_62,N_24964,N_24791);
nand UO_63 (O_63,N_24626,N_24726);
and UO_64 (O_64,N_24891,N_24730);
nand UO_65 (O_65,N_24932,N_24534);
nand UO_66 (O_66,N_24766,N_24639);
nor UO_67 (O_67,N_24656,N_24996);
nor UO_68 (O_68,N_24600,N_24878);
xor UO_69 (O_69,N_24796,N_24992);
and UO_70 (O_70,N_24779,N_24750);
nand UO_71 (O_71,N_24979,N_24655);
and UO_72 (O_72,N_24813,N_24482);
nor UO_73 (O_73,N_24804,N_24548);
nand UO_74 (O_74,N_24821,N_24715);
nor UO_75 (O_75,N_24599,N_24532);
or UO_76 (O_76,N_24884,N_24958);
nand UO_77 (O_77,N_24559,N_24765);
nand UO_78 (O_78,N_24449,N_24688);
nand UO_79 (O_79,N_24382,N_24636);
nand UO_80 (O_80,N_24612,N_24511);
and UO_81 (O_81,N_24415,N_24450);
and UO_82 (O_82,N_24944,N_24955);
nand UO_83 (O_83,N_24828,N_24531);
and UO_84 (O_84,N_24810,N_24385);
or UO_85 (O_85,N_24393,N_24769);
nor UO_86 (O_86,N_24774,N_24602);
or UO_87 (O_87,N_24522,N_24981);
nor UO_88 (O_88,N_24608,N_24832);
or UO_89 (O_89,N_24660,N_24629);
xor UO_90 (O_90,N_24589,N_24598);
and UO_91 (O_91,N_24409,N_24719);
or UO_92 (O_92,N_24407,N_24567);
nand UO_93 (O_93,N_24843,N_24610);
nor UO_94 (O_94,N_24717,N_24458);
or UO_95 (O_95,N_24543,N_24481);
nand UO_96 (O_96,N_24904,N_24800);
nand UO_97 (O_97,N_24512,N_24921);
nor UO_98 (O_98,N_24485,N_24603);
or UO_99 (O_99,N_24916,N_24661);
or UO_100 (O_100,N_24975,N_24470);
nand UO_101 (O_101,N_24818,N_24707);
nand UO_102 (O_102,N_24965,N_24484);
nor UO_103 (O_103,N_24571,N_24708);
nor UO_104 (O_104,N_24744,N_24712);
xnor UO_105 (O_105,N_24561,N_24617);
nand UO_106 (O_106,N_24986,N_24837);
and UO_107 (O_107,N_24941,N_24701);
or UO_108 (O_108,N_24506,N_24914);
nor UO_109 (O_109,N_24666,N_24950);
nand UO_110 (O_110,N_24499,N_24919);
and UO_111 (O_111,N_24634,N_24866);
nand UO_112 (O_112,N_24911,N_24882);
or UO_113 (O_113,N_24959,N_24938);
and UO_114 (O_114,N_24631,N_24539);
and UO_115 (O_115,N_24451,N_24789);
xnor UO_116 (O_116,N_24759,N_24844);
nor UO_117 (O_117,N_24434,N_24671);
or UO_118 (O_118,N_24438,N_24969);
nand UO_119 (O_119,N_24857,N_24886);
nor UO_120 (O_120,N_24713,N_24662);
and UO_121 (O_121,N_24420,N_24659);
and UO_122 (O_122,N_24505,N_24836);
nand UO_123 (O_123,N_24419,N_24859);
and UO_124 (O_124,N_24967,N_24745);
or UO_125 (O_125,N_24920,N_24573);
nor UO_126 (O_126,N_24991,N_24995);
nor UO_127 (O_127,N_24652,N_24683);
nor UO_128 (O_128,N_24754,N_24817);
nor UO_129 (O_129,N_24621,N_24595);
or UO_130 (O_130,N_24794,N_24901);
nand UO_131 (O_131,N_24445,N_24478);
or UO_132 (O_132,N_24980,N_24871);
and UO_133 (O_133,N_24777,N_24740);
and UO_134 (O_134,N_24410,N_24695);
and UO_135 (O_135,N_24929,N_24973);
nor UO_136 (O_136,N_24466,N_24593);
or UO_137 (O_137,N_24687,N_24862);
xnor UO_138 (O_138,N_24806,N_24840);
nand UO_139 (O_139,N_24809,N_24743);
nand UO_140 (O_140,N_24865,N_24389);
nand UO_141 (O_141,N_24628,N_24942);
or UO_142 (O_142,N_24490,N_24569);
or UO_143 (O_143,N_24703,N_24741);
nor UO_144 (O_144,N_24430,N_24391);
or UO_145 (O_145,N_24918,N_24885);
or UO_146 (O_146,N_24702,N_24549);
or UO_147 (O_147,N_24412,N_24530);
and UO_148 (O_148,N_24851,N_24524);
or UO_149 (O_149,N_24781,N_24641);
or UO_150 (O_150,N_24547,N_24579);
or UO_151 (O_151,N_24845,N_24898);
and UO_152 (O_152,N_24446,N_24902);
xnor UO_153 (O_153,N_24477,N_24494);
nand UO_154 (O_154,N_24545,N_24580);
xor UO_155 (O_155,N_24948,N_24786);
and UO_156 (O_156,N_24802,N_24578);
nor UO_157 (O_157,N_24946,N_24910);
nor UO_158 (O_158,N_24408,N_24879);
or UO_159 (O_159,N_24792,N_24767);
nor UO_160 (O_160,N_24762,N_24780);
or UO_161 (O_161,N_24960,N_24616);
nor UO_162 (O_162,N_24913,N_24785);
nor UO_163 (O_163,N_24480,N_24649);
nand UO_164 (O_164,N_24814,N_24983);
or UO_165 (O_165,N_24771,N_24811);
xor UO_166 (O_166,N_24515,N_24710);
and UO_167 (O_167,N_24928,N_24388);
nand UO_168 (O_168,N_24820,N_24924);
and UO_169 (O_169,N_24552,N_24847);
or UO_170 (O_170,N_24693,N_24807);
or UO_171 (O_171,N_24956,N_24550);
or UO_172 (O_172,N_24400,N_24907);
or UO_173 (O_173,N_24463,N_24732);
and UO_174 (O_174,N_24970,N_24473);
nand UO_175 (O_175,N_24801,N_24645);
nor UO_176 (O_176,N_24444,N_24873);
or UO_177 (O_177,N_24887,N_24816);
or UO_178 (O_178,N_24605,N_24827);
and UO_179 (O_179,N_24926,N_24949);
nand UO_180 (O_180,N_24971,N_24815);
or UO_181 (O_181,N_24888,N_24413);
or UO_182 (O_182,N_24897,N_24431);
nand UO_183 (O_183,N_24772,N_24627);
xnor UO_184 (O_184,N_24376,N_24930);
nand UO_185 (O_185,N_24805,N_24854);
nand UO_186 (O_186,N_24940,N_24459);
nand UO_187 (O_187,N_24465,N_24842);
nand UO_188 (O_188,N_24538,N_24890);
or UO_189 (O_189,N_24905,N_24736);
or UO_190 (O_190,N_24768,N_24936);
nand UO_191 (O_191,N_24838,N_24584);
xnor UO_192 (O_192,N_24984,N_24937);
nor UO_193 (O_193,N_24472,N_24414);
nand UO_194 (O_194,N_24609,N_24734);
nand UO_195 (O_195,N_24760,N_24667);
nor UO_196 (O_196,N_24588,N_24867);
nand UO_197 (O_197,N_24471,N_24863);
or UO_198 (O_198,N_24698,N_24640);
nor UO_199 (O_199,N_24999,N_24633);
nand UO_200 (O_200,N_24853,N_24697);
nand UO_201 (O_201,N_24556,N_24513);
nand UO_202 (O_202,N_24764,N_24507);
or UO_203 (O_203,N_24733,N_24432);
nor UO_204 (O_204,N_24423,N_24558);
nor UO_205 (O_205,N_24630,N_24390);
nand UO_206 (O_206,N_24690,N_24751);
nand UO_207 (O_207,N_24900,N_24966);
xnor UO_208 (O_208,N_24642,N_24467);
or UO_209 (O_209,N_24462,N_24893);
nor UO_210 (O_210,N_24824,N_24685);
xnor UO_211 (O_211,N_24379,N_24586);
xor UO_212 (O_212,N_24668,N_24829);
nand UO_213 (O_213,N_24520,N_24562);
and UO_214 (O_214,N_24535,N_24782);
nand UO_215 (O_215,N_24968,N_24553);
nor UO_216 (O_216,N_24525,N_24474);
or UO_217 (O_217,N_24541,N_24846);
nor UO_218 (O_218,N_24988,N_24997);
nor UO_219 (O_219,N_24684,N_24493);
xor UO_220 (O_220,N_24881,N_24442);
nand UO_221 (O_221,N_24699,N_24664);
or UO_222 (O_222,N_24411,N_24508);
nand UO_223 (O_223,N_24457,N_24706);
nor UO_224 (O_224,N_24453,N_24395);
nor UO_225 (O_225,N_24488,N_24963);
and UO_226 (O_226,N_24822,N_24738);
nand UO_227 (O_227,N_24475,N_24756);
nor UO_228 (O_228,N_24433,N_24489);
nand UO_229 (O_229,N_24521,N_24625);
or UO_230 (O_230,N_24681,N_24517);
and UO_231 (O_231,N_24504,N_24404);
or UO_232 (O_232,N_24747,N_24943);
or UO_233 (O_233,N_24908,N_24447);
or UO_234 (O_234,N_24978,N_24825);
and UO_235 (O_235,N_24613,N_24875);
and UO_236 (O_236,N_24739,N_24401);
or UO_237 (O_237,N_24876,N_24912);
xor UO_238 (O_238,N_24590,N_24381);
and UO_239 (O_239,N_24972,N_24954);
nand UO_240 (O_240,N_24757,N_24711);
or UO_241 (O_241,N_24427,N_24654);
or UO_242 (O_242,N_24849,N_24894);
or UO_243 (O_243,N_24607,N_24637);
nand UO_244 (O_244,N_24787,N_24468);
or UO_245 (O_245,N_24514,N_24566);
xnor UO_246 (O_246,N_24860,N_24933);
nand UO_247 (O_247,N_24501,N_24644);
nor UO_248 (O_248,N_24421,N_24422);
or UO_249 (O_249,N_24563,N_24510);
or UO_250 (O_250,N_24773,N_24826);
and UO_251 (O_251,N_24491,N_24778);
nand UO_252 (O_252,N_24479,N_24497);
and UO_253 (O_253,N_24748,N_24694);
or UO_254 (O_254,N_24648,N_24377);
and UO_255 (O_255,N_24378,N_24406);
and UO_256 (O_256,N_24714,N_24572);
or UO_257 (O_257,N_24939,N_24819);
or UO_258 (O_258,N_24709,N_24909);
xnor UO_259 (O_259,N_24646,N_24728);
and UO_260 (O_260,N_24989,N_24962);
nor UO_261 (O_261,N_24417,N_24544);
nand UO_262 (O_262,N_24632,N_24746);
nand UO_263 (O_263,N_24705,N_24682);
xnor UO_264 (O_264,N_24724,N_24568);
nor UO_265 (O_265,N_24528,N_24993);
or UO_266 (O_266,N_24673,N_24896);
or UO_267 (O_267,N_24864,N_24476);
or UO_268 (O_268,N_24624,N_24720);
and UO_269 (O_269,N_24850,N_24615);
nand UO_270 (O_270,N_24823,N_24585);
and UO_271 (O_271,N_24852,N_24405);
or UO_272 (O_272,N_24596,N_24752);
and UO_273 (O_273,N_24500,N_24895);
and UO_274 (O_274,N_24998,N_24526);
and UO_275 (O_275,N_24375,N_24892);
nor UO_276 (O_276,N_24650,N_24855);
xnor UO_277 (O_277,N_24812,N_24856);
nor UO_278 (O_278,N_24426,N_24604);
xor UO_279 (O_279,N_24872,N_24436);
xor UO_280 (O_280,N_24399,N_24737);
and UO_281 (O_281,N_24601,N_24454);
and UO_282 (O_282,N_24542,N_24653);
and UO_283 (O_283,N_24951,N_24469);
nand UO_284 (O_284,N_24961,N_24577);
nand UO_285 (O_285,N_24536,N_24923);
and UO_286 (O_286,N_24670,N_24899);
nor UO_287 (O_287,N_24622,N_24716);
and UO_288 (O_288,N_24592,N_24915);
xnor UO_289 (O_289,N_24753,N_24831);
xor UO_290 (O_290,N_24990,N_24830);
nor UO_291 (O_291,N_24788,N_24976);
xor UO_292 (O_292,N_24483,N_24922);
or UO_293 (O_293,N_24519,N_24678);
nand UO_294 (O_294,N_24529,N_24498);
nand UO_295 (O_295,N_24564,N_24614);
and UO_296 (O_296,N_24952,N_24742);
or UO_297 (O_297,N_24858,N_24509);
and UO_298 (O_298,N_24689,N_24974);
or UO_299 (O_299,N_24574,N_24953);
nor UO_300 (O_300,N_24676,N_24833);
nand UO_301 (O_301,N_24647,N_24576);
nand UO_302 (O_302,N_24591,N_24763);
and UO_303 (O_303,N_24518,N_24677);
and UO_304 (O_304,N_24770,N_24723);
nand UO_305 (O_305,N_24692,N_24583);
nor UO_306 (O_306,N_24977,N_24657);
nor UO_307 (O_307,N_24889,N_24727);
or UO_308 (O_308,N_24947,N_24861);
or UO_309 (O_309,N_24841,N_24883);
nand UO_310 (O_310,N_24793,N_24448);
nor UO_311 (O_311,N_24441,N_24803);
or UO_312 (O_312,N_24392,N_24518);
or UO_313 (O_313,N_24384,N_24573);
nand UO_314 (O_314,N_24768,N_24804);
xor UO_315 (O_315,N_24772,N_24786);
and UO_316 (O_316,N_24707,N_24907);
nor UO_317 (O_317,N_24952,N_24388);
nor UO_318 (O_318,N_24722,N_24947);
nor UO_319 (O_319,N_24937,N_24593);
or UO_320 (O_320,N_24767,N_24403);
or UO_321 (O_321,N_24932,N_24607);
or UO_322 (O_322,N_24558,N_24569);
and UO_323 (O_323,N_24741,N_24686);
and UO_324 (O_324,N_24717,N_24412);
nor UO_325 (O_325,N_24565,N_24412);
or UO_326 (O_326,N_24918,N_24955);
nand UO_327 (O_327,N_24919,N_24484);
and UO_328 (O_328,N_24717,N_24550);
nand UO_329 (O_329,N_24863,N_24788);
nand UO_330 (O_330,N_24961,N_24900);
and UO_331 (O_331,N_24388,N_24691);
xnor UO_332 (O_332,N_24612,N_24746);
nand UO_333 (O_333,N_24424,N_24587);
and UO_334 (O_334,N_24388,N_24929);
nor UO_335 (O_335,N_24424,N_24495);
nand UO_336 (O_336,N_24954,N_24991);
or UO_337 (O_337,N_24910,N_24945);
nor UO_338 (O_338,N_24713,N_24899);
or UO_339 (O_339,N_24788,N_24793);
xnor UO_340 (O_340,N_24939,N_24775);
nand UO_341 (O_341,N_24770,N_24677);
nor UO_342 (O_342,N_24743,N_24534);
nand UO_343 (O_343,N_24416,N_24886);
or UO_344 (O_344,N_24558,N_24665);
nor UO_345 (O_345,N_24679,N_24386);
nor UO_346 (O_346,N_24641,N_24797);
and UO_347 (O_347,N_24556,N_24602);
xor UO_348 (O_348,N_24825,N_24529);
nand UO_349 (O_349,N_24961,N_24615);
nand UO_350 (O_350,N_24388,N_24920);
or UO_351 (O_351,N_24619,N_24876);
nor UO_352 (O_352,N_24736,N_24443);
or UO_353 (O_353,N_24955,N_24679);
xor UO_354 (O_354,N_24534,N_24712);
xor UO_355 (O_355,N_24463,N_24809);
nand UO_356 (O_356,N_24391,N_24424);
xor UO_357 (O_357,N_24477,N_24929);
nand UO_358 (O_358,N_24683,N_24735);
nand UO_359 (O_359,N_24663,N_24481);
nor UO_360 (O_360,N_24956,N_24968);
nand UO_361 (O_361,N_24473,N_24563);
nor UO_362 (O_362,N_24909,N_24438);
nor UO_363 (O_363,N_24445,N_24767);
nand UO_364 (O_364,N_24855,N_24985);
and UO_365 (O_365,N_24479,N_24424);
xor UO_366 (O_366,N_24992,N_24970);
nor UO_367 (O_367,N_24477,N_24386);
nand UO_368 (O_368,N_24451,N_24919);
nor UO_369 (O_369,N_24751,N_24786);
or UO_370 (O_370,N_24776,N_24454);
and UO_371 (O_371,N_24648,N_24689);
nand UO_372 (O_372,N_24940,N_24447);
nor UO_373 (O_373,N_24959,N_24931);
and UO_374 (O_374,N_24970,N_24905);
nor UO_375 (O_375,N_24513,N_24913);
nand UO_376 (O_376,N_24639,N_24992);
nor UO_377 (O_377,N_24852,N_24831);
or UO_378 (O_378,N_24836,N_24819);
nand UO_379 (O_379,N_24690,N_24866);
and UO_380 (O_380,N_24939,N_24763);
or UO_381 (O_381,N_24777,N_24812);
or UO_382 (O_382,N_24974,N_24481);
nand UO_383 (O_383,N_24686,N_24748);
nor UO_384 (O_384,N_24506,N_24629);
nor UO_385 (O_385,N_24820,N_24946);
nor UO_386 (O_386,N_24654,N_24603);
or UO_387 (O_387,N_24862,N_24625);
and UO_388 (O_388,N_24879,N_24420);
or UO_389 (O_389,N_24787,N_24570);
nor UO_390 (O_390,N_24875,N_24654);
nor UO_391 (O_391,N_24603,N_24694);
nor UO_392 (O_392,N_24384,N_24559);
nor UO_393 (O_393,N_24750,N_24736);
or UO_394 (O_394,N_24561,N_24786);
nand UO_395 (O_395,N_24575,N_24798);
or UO_396 (O_396,N_24854,N_24961);
or UO_397 (O_397,N_24648,N_24678);
nor UO_398 (O_398,N_24384,N_24836);
or UO_399 (O_399,N_24788,N_24626);
or UO_400 (O_400,N_24520,N_24971);
nor UO_401 (O_401,N_24798,N_24416);
nand UO_402 (O_402,N_24871,N_24578);
or UO_403 (O_403,N_24761,N_24883);
nor UO_404 (O_404,N_24533,N_24906);
nand UO_405 (O_405,N_24394,N_24950);
or UO_406 (O_406,N_24834,N_24576);
nor UO_407 (O_407,N_24573,N_24710);
and UO_408 (O_408,N_24557,N_24845);
and UO_409 (O_409,N_24831,N_24870);
or UO_410 (O_410,N_24831,N_24704);
nand UO_411 (O_411,N_24449,N_24438);
or UO_412 (O_412,N_24913,N_24682);
nor UO_413 (O_413,N_24819,N_24974);
and UO_414 (O_414,N_24583,N_24744);
and UO_415 (O_415,N_24460,N_24989);
or UO_416 (O_416,N_24439,N_24456);
and UO_417 (O_417,N_24599,N_24785);
and UO_418 (O_418,N_24963,N_24625);
and UO_419 (O_419,N_24928,N_24972);
or UO_420 (O_420,N_24615,N_24433);
and UO_421 (O_421,N_24943,N_24822);
and UO_422 (O_422,N_24757,N_24776);
nor UO_423 (O_423,N_24794,N_24524);
nand UO_424 (O_424,N_24409,N_24957);
and UO_425 (O_425,N_24492,N_24412);
or UO_426 (O_426,N_24475,N_24851);
nor UO_427 (O_427,N_24696,N_24511);
nand UO_428 (O_428,N_24522,N_24513);
or UO_429 (O_429,N_24711,N_24592);
nand UO_430 (O_430,N_24740,N_24398);
xnor UO_431 (O_431,N_24891,N_24913);
nor UO_432 (O_432,N_24924,N_24432);
nand UO_433 (O_433,N_24394,N_24593);
and UO_434 (O_434,N_24509,N_24408);
and UO_435 (O_435,N_24782,N_24573);
or UO_436 (O_436,N_24940,N_24728);
and UO_437 (O_437,N_24614,N_24811);
xnor UO_438 (O_438,N_24485,N_24474);
xor UO_439 (O_439,N_24948,N_24721);
nand UO_440 (O_440,N_24455,N_24489);
or UO_441 (O_441,N_24606,N_24491);
nand UO_442 (O_442,N_24746,N_24691);
or UO_443 (O_443,N_24425,N_24489);
nor UO_444 (O_444,N_24619,N_24825);
nor UO_445 (O_445,N_24507,N_24844);
nor UO_446 (O_446,N_24993,N_24390);
nor UO_447 (O_447,N_24631,N_24923);
and UO_448 (O_448,N_24661,N_24404);
or UO_449 (O_449,N_24558,N_24962);
or UO_450 (O_450,N_24518,N_24785);
nand UO_451 (O_451,N_24489,N_24387);
nand UO_452 (O_452,N_24409,N_24435);
nor UO_453 (O_453,N_24708,N_24472);
nor UO_454 (O_454,N_24810,N_24907);
or UO_455 (O_455,N_24593,N_24532);
and UO_456 (O_456,N_24829,N_24418);
xnor UO_457 (O_457,N_24515,N_24717);
nand UO_458 (O_458,N_24700,N_24856);
or UO_459 (O_459,N_24671,N_24899);
nor UO_460 (O_460,N_24621,N_24758);
or UO_461 (O_461,N_24823,N_24977);
nor UO_462 (O_462,N_24433,N_24824);
xnor UO_463 (O_463,N_24783,N_24409);
xor UO_464 (O_464,N_24936,N_24531);
nand UO_465 (O_465,N_24749,N_24694);
or UO_466 (O_466,N_24735,N_24602);
nor UO_467 (O_467,N_24946,N_24760);
xor UO_468 (O_468,N_24581,N_24627);
and UO_469 (O_469,N_24794,N_24912);
and UO_470 (O_470,N_24516,N_24940);
and UO_471 (O_471,N_24704,N_24891);
and UO_472 (O_472,N_24736,N_24899);
and UO_473 (O_473,N_24640,N_24879);
nor UO_474 (O_474,N_24515,N_24782);
nor UO_475 (O_475,N_24958,N_24950);
and UO_476 (O_476,N_24527,N_24669);
nor UO_477 (O_477,N_24695,N_24799);
or UO_478 (O_478,N_24810,N_24432);
and UO_479 (O_479,N_24469,N_24598);
and UO_480 (O_480,N_24615,N_24936);
nand UO_481 (O_481,N_24408,N_24711);
and UO_482 (O_482,N_24703,N_24801);
nand UO_483 (O_483,N_24842,N_24688);
nand UO_484 (O_484,N_24787,N_24732);
nor UO_485 (O_485,N_24397,N_24741);
or UO_486 (O_486,N_24470,N_24766);
or UO_487 (O_487,N_24494,N_24906);
nand UO_488 (O_488,N_24848,N_24865);
and UO_489 (O_489,N_24664,N_24557);
or UO_490 (O_490,N_24662,N_24944);
and UO_491 (O_491,N_24467,N_24646);
and UO_492 (O_492,N_24764,N_24670);
nor UO_493 (O_493,N_24521,N_24542);
or UO_494 (O_494,N_24386,N_24879);
and UO_495 (O_495,N_24991,N_24403);
and UO_496 (O_496,N_24951,N_24561);
or UO_497 (O_497,N_24497,N_24804);
nor UO_498 (O_498,N_24461,N_24486);
and UO_499 (O_499,N_24895,N_24661);
nand UO_500 (O_500,N_24424,N_24455);
xnor UO_501 (O_501,N_24895,N_24523);
nand UO_502 (O_502,N_24756,N_24650);
xor UO_503 (O_503,N_24988,N_24753);
and UO_504 (O_504,N_24593,N_24833);
nand UO_505 (O_505,N_24827,N_24393);
and UO_506 (O_506,N_24812,N_24509);
nand UO_507 (O_507,N_24764,N_24403);
nand UO_508 (O_508,N_24893,N_24841);
nand UO_509 (O_509,N_24774,N_24891);
nand UO_510 (O_510,N_24799,N_24537);
or UO_511 (O_511,N_24429,N_24848);
and UO_512 (O_512,N_24387,N_24921);
and UO_513 (O_513,N_24975,N_24456);
and UO_514 (O_514,N_24408,N_24650);
or UO_515 (O_515,N_24602,N_24672);
nor UO_516 (O_516,N_24479,N_24687);
or UO_517 (O_517,N_24874,N_24720);
nor UO_518 (O_518,N_24635,N_24844);
nor UO_519 (O_519,N_24379,N_24782);
or UO_520 (O_520,N_24902,N_24600);
and UO_521 (O_521,N_24583,N_24924);
nand UO_522 (O_522,N_24627,N_24886);
nor UO_523 (O_523,N_24688,N_24573);
xnor UO_524 (O_524,N_24510,N_24727);
nand UO_525 (O_525,N_24951,N_24625);
and UO_526 (O_526,N_24399,N_24678);
nor UO_527 (O_527,N_24434,N_24411);
or UO_528 (O_528,N_24384,N_24960);
or UO_529 (O_529,N_24931,N_24811);
or UO_530 (O_530,N_24609,N_24668);
and UO_531 (O_531,N_24935,N_24708);
and UO_532 (O_532,N_24699,N_24794);
nor UO_533 (O_533,N_24829,N_24712);
or UO_534 (O_534,N_24502,N_24966);
and UO_535 (O_535,N_24492,N_24791);
nor UO_536 (O_536,N_24508,N_24566);
xnor UO_537 (O_537,N_24964,N_24829);
and UO_538 (O_538,N_24660,N_24477);
nand UO_539 (O_539,N_24948,N_24997);
xor UO_540 (O_540,N_24696,N_24439);
nand UO_541 (O_541,N_24713,N_24803);
and UO_542 (O_542,N_24694,N_24800);
nor UO_543 (O_543,N_24714,N_24395);
or UO_544 (O_544,N_24680,N_24743);
nand UO_545 (O_545,N_24945,N_24724);
nand UO_546 (O_546,N_24736,N_24789);
and UO_547 (O_547,N_24668,N_24564);
or UO_548 (O_548,N_24438,N_24486);
and UO_549 (O_549,N_24895,N_24676);
nand UO_550 (O_550,N_24390,N_24577);
nor UO_551 (O_551,N_24982,N_24589);
xor UO_552 (O_552,N_24967,N_24697);
xor UO_553 (O_553,N_24654,N_24771);
nand UO_554 (O_554,N_24726,N_24988);
nor UO_555 (O_555,N_24974,N_24873);
or UO_556 (O_556,N_24817,N_24680);
or UO_557 (O_557,N_24698,N_24685);
or UO_558 (O_558,N_24916,N_24963);
or UO_559 (O_559,N_24516,N_24549);
or UO_560 (O_560,N_24514,N_24855);
or UO_561 (O_561,N_24910,N_24776);
or UO_562 (O_562,N_24617,N_24398);
or UO_563 (O_563,N_24971,N_24756);
and UO_564 (O_564,N_24709,N_24672);
or UO_565 (O_565,N_24506,N_24874);
or UO_566 (O_566,N_24842,N_24552);
nor UO_567 (O_567,N_24532,N_24747);
and UO_568 (O_568,N_24657,N_24877);
or UO_569 (O_569,N_24884,N_24487);
and UO_570 (O_570,N_24446,N_24494);
or UO_571 (O_571,N_24876,N_24919);
nor UO_572 (O_572,N_24605,N_24488);
nor UO_573 (O_573,N_24875,N_24447);
and UO_574 (O_574,N_24868,N_24454);
and UO_575 (O_575,N_24917,N_24776);
nand UO_576 (O_576,N_24966,N_24875);
and UO_577 (O_577,N_24924,N_24571);
and UO_578 (O_578,N_24959,N_24540);
and UO_579 (O_579,N_24406,N_24534);
xnor UO_580 (O_580,N_24764,N_24972);
nand UO_581 (O_581,N_24647,N_24766);
nand UO_582 (O_582,N_24400,N_24721);
and UO_583 (O_583,N_24569,N_24662);
and UO_584 (O_584,N_24770,N_24810);
and UO_585 (O_585,N_24553,N_24900);
and UO_586 (O_586,N_24612,N_24930);
or UO_587 (O_587,N_24527,N_24672);
or UO_588 (O_588,N_24574,N_24520);
nor UO_589 (O_589,N_24949,N_24495);
and UO_590 (O_590,N_24857,N_24447);
nand UO_591 (O_591,N_24983,N_24876);
nor UO_592 (O_592,N_24427,N_24466);
and UO_593 (O_593,N_24586,N_24853);
or UO_594 (O_594,N_24593,N_24602);
and UO_595 (O_595,N_24970,N_24688);
xnor UO_596 (O_596,N_24530,N_24989);
or UO_597 (O_597,N_24516,N_24874);
or UO_598 (O_598,N_24462,N_24428);
nor UO_599 (O_599,N_24597,N_24731);
nand UO_600 (O_600,N_24689,N_24383);
and UO_601 (O_601,N_24521,N_24752);
nand UO_602 (O_602,N_24481,N_24857);
nor UO_603 (O_603,N_24574,N_24776);
and UO_604 (O_604,N_24735,N_24436);
nor UO_605 (O_605,N_24586,N_24558);
or UO_606 (O_606,N_24978,N_24758);
nand UO_607 (O_607,N_24463,N_24712);
or UO_608 (O_608,N_24820,N_24377);
nor UO_609 (O_609,N_24841,N_24671);
nor UO_610 (O_610,N_24807,N_24682);
nor UO_611 (O_611,N_24571,N_24724);
nand UO_612 (O_612,N_24448,N_24575);
nand UO_613 (O_613,N_24894,N_24584);
or UO_614 (O_614,N_24974,N_24614);
or UO_615 (O_615,N_24542,N_24548);
or UO_616 (O_616,N_24776,N_24985);
nor UO_617 (O_617,N_24791,N_24924);
nand UO_618 (O_618,N_24464,N_24872);
nor UO_619 (O_619,N_24816,N_24635);
nand UO_620 (O_620,N_24939,N_24635);
or UO_621 (O_621,N_24842,N_24627);
nand UO_622 (O_622,N_24503,N_24387);
and UO_623 (O_623,N_24474,N_24427);
and UO_624 (O_624,N_24989,N_24959);
nand UO_625 (O_625,N_24689,N_24551);
nor UO_626 (O_626,N_24739,N_24847);
nand UO_627 (O_627,N_24421,N_24941);
and UO_628 (O_628,N_24384,N_24561);
xnor UO_629 (O_629,N_24436,N_24579);
xnor UO_630 (O_630,N_24502,N_24523);
and UO_631 (O_631,N_24587,N_24860);
nor UO_632 (O_632,N_24543,N_24538);
nand UO_633 (O_633,N_24777,N_24469);
nand UO_634 (O_634,N_24734,N_24831);
or UO_635 (O_635,N_24729,N_24453);
nor UO_636 (O_636,N_24581,N_24584);
and UO_637 (O_637,N_24964,N_24517);
xnor UO_638 (O_638,N_24479,N_24419);
nand UO_639 (O_639,N_24403,N_24789);
or UO_640 (O_640,N_24543,N_24881);
nand UO_641 (O_641,N_24558,N_24787);
nand UO_642 (O_642,N_24623,N_24522);
and UO_643 (O_643,N_24662,N_24444);
nand UO_644 (O_644,N_24416,N_24923);
nor UO_645 (O_645,N_24936,N_24409);
xnor UO_646 (O_646,N_24458,N_24805);
nor UO_647 (O_647,N_24447,N_24729);
or UO_648 (O_648,N_24774,N_24999);
nor UO_649 (O_649,N_24894,N_24743);
or UO_650 (O_650,N_24559,N_24644);
nand UO_651 (O_651,N_24913,N_24739);
nand UO_652 (O_652,N_24669,N_24971);
nor UO_653 (O_653,N_24512,N_24784);
nand UO_654 (O_654,N_24974,N_24461);
or UO_655 (O_655,N_24613,N_24433);
nor UO_656 (O_656,N_24477,N_24787);
or UO_657 (O_657,N_24773,N_24712);
nand UO_658 (O_658,N_24545,N_24558);
nand UO_659 (O_659,N_24920,N_24792);
nor UO_660 (O_660,N_24406,N_24857);
and UO_661 (O_661,N_24389,N_24630);
and UO_662 (O_662,N_24667,N_24422);
nor UO_663 (O_663,N_24738,N_24706);
and UO_664 (O_664,N_24896,N_24439);
or UO_665 (O_665,N_24772,N_24683);
nand UO_666 (O_666,N_24771,N_24571);
nand UO_667 (O_667,N_24551,N_24644);
or UO_668 (O_668,N_24596,N_24978);
nand UO_669 (O_669,N_24541,N_24837);
xnor UO_670 (O_670,N_24583,N_24580);
nand UO_671 (O_671,N_24415,N_24538);
nand UO_672 (O_672,N_24634,N_24854);
and UO_673 (O_673,N_24794,N_24764);
and UO_674 (O_674,N_24775,N_24936);
or UO_675 (O_675,N_24619,N_24429);
nor UO_676 (O_676,N_24716,N_24448);
or UO_677 (O_677,N_24423,N_24858);
and UO_678 (O_678,N_24688,N_24620);
nand UO_679 (O_679,N_24701,N_24546);
nand UO_680 (O_680,N_24930,N_24685);
or UO_681 (O_681,N_24741,N_24725);
or UO_682 (O_682,N_24414,N_24701);
or UO_683 (O_683,N_24434,N_24605);
or UO_684 (O_684,N_24709,N_24566);
nor UO_685 (O_685,N_24483,N_24931);
nor UO_686 (O_686,N_24783,N_24496);
and UO_687 (O_687,N_24783,N_24802);
xnor UO_688 (O_688,N_24607,N_24938);
and UO_689 (O_689,N_24929,N_24386);
nand UO_690 (O_690,N_24577,N_24546);
and UO_691 (O_691,N_24519,N_24637);
xor UO_692 (O_692,N_24972,N_24456);
nand UO_693 (O_693,N_24629,N_24805);
or UO_694 (O_694,N_24825,N_24949);
nor UO_695 (O_695,N_24709,N_24754);
or UO_696 (O_696,N_24538,N_24715);
nand UO_697 (O_697,N_24737,N_24739);
or UO_698 (O_698,N_24919,N_24818);
and UO_699 (O_699,N_24585,N_24939);
nand UO_700 (O_700,N_24690,N_24693);
xor UO_701 (O_701,N_24884,N_24435);
nand UO_702 (O_702,N_24847,N_24977);
or UO_703 (O_703,N_24816,N_24486);
nor UO_704 (O_704,N_24536,N_24874);
nand UO_705 (O_705,N_24751,N_24445);
nand UO_706 (O_706,N_24806,N_24876);
nor UO_707 (O_707,N_24923,N_24945);
nor UO_708 (O_708,N_24434,N_24618);
nand UO_709 (O_709,N_24597,N_24928);
nand UO_710 (O_710,N_24926,N_24517);
nor UO_711 (O_711,N_24964,N_24983);
nor UO_712 (O_712,N_24705,N_24535);
xor UO_713 (O_713,N_24812,N_24377);
nor UO_714 (O_714,N_24897,N_24574);
or UO_715 (O_715,N_24867,N_24440);
nand UO_716 (O_716,N_24810,N_24956);
and UO_717 (O_717,N_24779,N_24762);
nand UO_718 (O_718,N_24434,N_24888);
nor UO_719 (O_719,N_24831,N_24494);
or UO_720 (O_720,N_24536,N_24602);
nand UO_721 (O_721,N_24406,N_24941);
nand UO_722 (O_722,N_24678,N_24925);
nor UO_723 (O_723,N_24556,N_24820);
or UO_724 (O_724,N_24559,N_24771);
nand UO_725 (O_725,N_24946,N_24643);
xnor UO_726 (O_726,N_24947,N_24457);
nand UO_727 (O_727,N_24824,N_24579);
xor UO_728 (O_728,N_24754,N_24639);
xor UO_729 (O_729,N_24962,N_24973);
nand UO_730 (O_730,N_24756,N_24995);
or UO_731 (O_731,N_24853,N_24595);
or UO_732 (O_732,N_24705,N_24937);
nand UO_733 (O_733,N_24710,N_24411);
or UO_734 (O_734,N_24902,N_24580);
xnor UO_735 (O_735,N_24723,N_24931);
nor UO_736 (O_736,N_24489,N_24976);
nand UO_737 (O_737,N_24529,N_24455);
or UO_738 (O_738,N_24517,N_24618);
nor UO_739 (O_739,N_24769,N_24794);
nand UO_740 (O_740,N_24630,N_24937);
or UO_741 (O_741,N_24520,N_24598);
nand UO_742 (O_742,N_24903,N_24953);
or UO_743 (O_743,N_24843,N_24638);
nor UO_744 (O_744,N_24487,N_24452);
nand UO_745 (O_745,N_24923,N_24857);
nor UO_746 (O_746,N_24936,N_24524);
nand UO_747 (O_747,N_24922,N_24606);
and UO_748 (O_748,N_24775,N_24900);
and UO_749 (O_749,N_24525,N_24548);
and UO_750 (O_750,N_24759,N_24968);
nor UO_751 (O_751,N_24982,N_24972);
or UO_752 (O_752,N_24394,N_24829);
nand UO_753 (O_753,N_24678,N_24414);
nor UO_754 (O_754,N_24505,N_24933);
xor UO_755 (O_755,N_24735,N_24765);
nor UO_756 (O_756,N_24652,N_24740);
and UO_757 (O_757,N_24617,N_24828);
and UO_758 (O_758,N_24842,N_24956);
nor UO_759 (O_759,N_24971,N_24844);
nand UO_760 (O_760,N_24511,N_24744);
nand UO_761 (O_761,N_24543,N_24569);
xor UO_762 (O_762,N_24423,N_24735);
xor UO_763 (O_763,N_24954,N_24417);
and UO_764 (O_764,N_24887,N_24634);
and UO_765 (O_765,N_24581,N_24426);
nand UO_766 (O_766,N_24840,N_24454);
nand UO_767 (O_767,N_24636,N_24511);
nand UO_768 (O_768,N_24476,N_24588);
nand UO_769 (O_769,N_24422,N_24617);
nand UO_770 (O_770,N_24773,N_24900);
and UO_771 (O_771,N_24938,N_24736);
and UO_772 (O_772,N_24823,N_24687);
and UO_773 (O_773,N_24655,N_24910);
or UO_774 (O_774,N_24735,N_24411);
and UO_775 (O_775,N_24845,N_24491);
xor UO_776 (O_776,N_24891,N_24388);
and UO_777 (O_777,N_24827,N_24502);
nor UO_778 (O_778,N_24616,N_24941);
nand UO_779 (O_779,N_24691,N_24979);
xor UO_780 (O_780,N_24421,N_24908);
and UO_781 (O_781,N_24495,N_24973);
or UO_782 (O_782,N_24964,N_24947);
nor UO_783 (O_783,N_24477,N_24771);
nor UO_784 (O_784,N_24864,N_24647);
or UO_785 (O_785,N_24827,N_24831);
or UO_786 (O_786,N_24696,N_24630);
and UO_787 (O_787,N_24667,N_24721);
xor UO_788 (O_788,N_24539,N_24732);
and UO_789 (O_789,N_24571,N_24668);
nor UO_790 (O_790,N_24714,N_24736);
or UO_791 (O_791,N_24946,N_24929);
and UO_792 (O_792,N_24916,N_24726);
or UO_793 (O_793,N_24967,N_24577);
nand UO_794 (O_794,N_24428,N_24863);
or UO_795 (O_795,N_24843,N_24642);
or UO_796 (O_796,N_24948,N_24459);
nand UO_797 (O_797,N_24645,N_24598);
nand UO_798 (O_798,N_24700,N_24637);
nor UO_799 (O_799,N_24432,N_24539);
xor UO_800 (O_800,N_24713,N_24931);
xnor UO_801 (O_801,N_24688,N_24949);
nand UO_802 (O_802,N_24821,N_24950);
and UO_803 (O_803,N_24906,N_24564);
xor UO_804 (O_804,N_24748,N_24552);
and UO_805 (O_805,N_24897,N_24654);
nand UO_806 (O_806,N_24846,N_24506);
and UO_807 (O_807,N_24437,N_24770);
nand UO_808 (O_808,N_24738,N_24917);
nor UO_809 (O_809,N_24808,N_24625);
nand UO_810 (O_810,N_24433,N_24814);
nand UO_811 (O_811,N_24858,N_24664);
or UO_812 (O_812,N_24525,N_24792);
and UO_813 (O_813,N_24992,N_24749);
nand UO_814 (O_814,N_24700,N_24633);
and UO_815 (O_815,N_24902,N_24382);
and UO_816 (O_816,N_24782,N_24925);
and UO_817 (O_817,N_24761,N_24957);
nor UO_818 (O_818,N_24976,N_24854);
or UO_819 (O_819,N_24666,N_24599);
or UO_820 (O_820,N_24571,N_24572);
xor UO_821 (O_821,N_24991,N_24634);
or UO_822 (O_822,N_24708,N_24532);
nand UO_823 (O_823,N_24762,N_24745);
nand UO_824 (O_824,N_24860,N_24741);
or UO_825 (O_825,N_24393,N_24891);
nand UO_826 (O_826,N_24795,N_24523);
and UO_827 (O_827,N_24825,N_24571);
and UO_828 (O_828,N_24401,N_24409);
nand UO_829 (O_829,N_24615,N_24570);
or UO_830 (O_830,N_24473,N_24492);
and UO_831 (O_831,N_24466,N_24412);
nor UO_832 (O_832,N_24620,N_24402);
nand UO_833 (O_833,N_24483,N_24638);
and UO_834 (O_834,N_24629,N_24999);
nand UO_835 (O_835,N_24826,N_24640);
nand UO_836 (O_836,N_24936,N_24647);
and UO_837 (O_837,N_24457,N_24925);
nand UO_838 (O_838,N_24846,N_24558);
or UO_839 (O_839,N_24708,N_24840);
xnor UO_840 (O_840,N_24418,N_24775);
nor UO_841 (O_841,N_24968,N_24625);
nor UO_842 (O_842,N_24988,N_24655);
or UO_843 (O_843,N_24506,N_24782);
xor UO_844 (O_844,N_24736,N_24571);
or UO_845 (O_845,N_24950,N_24962);
nor UO_846 (O_846,N_24913,N_24796);
and UO_847 (O_847,N_24831,N_24500);
and UO_848 (O_848,N_24564,N_24608);
xor UO_849 (O_849,N_24553,N_24624);
nand UO_850 (O_850,N_24499,N_24694);
nor UO_851 (O_851,N_24458,N_24623);
or UO_852 (O_852,N_24574,N_24494);
nor UO_853 (O_853,N_24585,N_24868);
nand UO_854 (O_854,N_24884,N_24802);
nor UO_855 (O_855,N_24915,N_24997);
nand UO_856 (O_856,N_24737,N_24865);
or UO_857 (O_857,N_24932,N_24961);
nand UO_858 (O_858,N_24848,N_24646);
nor UO_859 (O_859,N_24606,N_24659);
and UO_860 (O_860,N_24768,N_24923);
or UO_861 (O_861,N_24404,N_24470);
nand UO_862 (O_862,N_24947,N_24419);
xnor UO_863 (O_863,N_24467,N_24423);
nand UO_864 (O_864,N_24589,N_24400);
and UO_865 (O_865,N_24706,N_24761);
nand UO_866 (O_866,N_24396,N_24823);
nor UO_867 (O_867,N_24430,N_24980);
and UO_868 (O_868,N_24990,N_24645);
and UO_869 (O_869,N_24467,N_24906);
or UO_870 (O_870,N_24758,N_24885);
nand UO_871 (O_871,N_24401,N_24931);
xor UO_872 (O_872,N_24610,N_24768);
nand UO_873 (O_873,N_24532,N_24709);
and UO_874 (O_874,N_24517,N_24586);
and UO_875 (O_875,N_24828,N_24405);
or UO_876 (O_876,N_24922,N_24808);
xnor UO_877 (O_877,N_24828,N_24557);
nand UO_878 (O_878,N_24656,N_24629);
or UO_879 (O_879,N_24427,N_24877);
nor UO_880 (O_880,N_24673,N_24847);
nand UO_881 (O_881,N_24656,N_24671);
or UO_882 (O_882,N_24472,N_24430);
xnor UO_883 (O_883,N_24931,N_24818);
nand UO_884 (O_884,N_24566,N_24526);
nand UO_885 (O_885,N_24485,N_24561);
and UO_886 (O_886,N_24467,N_24904);
nand UO_887 (O_887,N_24473,N_24659);
and UO_888 (O_888,N_24411,N_24804);
nor UO_889 (O_889,N_24684,N_24743);
and UO_890 (O_890,N_24458,N_24948);
or UO_891 (O_891,N_24488,N_24427);
nor UO_892 (O_892,N_24668,N_24407);
or UO_893 (O_893,N_24384,N_24938);
nand UO_894 (O_894,N_24932,N_24832);
nor UO_895 (O_895,N_24909,N_24799);
nor UO_896 (O_896,N_24597,N_24868);
and UO_897 (O_897,N_24971,N_24984);
or UO_898 (O_898,N_24895,N_24936);
nor UO_899 (O_899,N_24776,N_24442);
nand UO_900 (O_900,N_24533,N_24919);
and UO_901 (O_901,N_24569,N_24561);
or UO_902 (O_902,N_24602,N_24758);
or UO_903 (O_903,N_24524,N_24612);
nand UO_904 (O_904,N_24868,N_24611);
xnor UO_905 (O_905,N_24897,N_24644);
or UO_906 (O_906,N_24777,N_24511);
nor UO_907 (O_907,N_24953,N_24441);
or UO_908 (O_908,N_24745,N_24748);
or UO_909 (O_909,N_24662,N_24639);
or UO_910 (O_910,N_24973,N_24990);
or UO_911 (O_911,N_24955,N_24623);
and UO_912 (O_912,N_24828,N_24621);
nand UO_913 (O_913,N_24978,N_24723);
and UO_914 (O_914,N_24991,N_24488);
or UO_915 (O_915,N_24597,N_24823);
nor UO_916 (O_916,N_24781,N_24954);
or UO_917 (O_917,N_24530,N_24855);
and UO_918 (O_918,N_24677,N_24979);
and UO_919 (O_919,N_24621,N_24737);
nand UO_920 (O_920,N_24770,N_24788);
and UO_921 (O_921,N_24929,N_24683);
nor UO_922 (O_922,N_24613,N_24883);
nor UO_923 (O_923,N_24958,N_24993);
and UO_924 (O_924,N_24571,N_24782);
nor UO_925 (O_925,N_24533,N_24463);
nor UO_926 (O_926,N_24868,N_24563);
nor UO_927 (O_927,N_24929,N_24987);
or UO_928 (O_928,N_24488,N_24776);
xnor UO_929 (O_929,N_24390,N_24964);
nor UO_930 (O_930,N_24883,N_24860);
or UO_931 (O_931,N_24581,N_24504);
and UO_932 (O_932,N_24806,N_24560);
or UO_933 (O_933,N_24935,N_24604);
xnor UO_934 (O_934,N_24993,N_24877);
and UO_935 (O_935,N_24909,N_24755);
and UO_936 (O_936,N_24497,N_24389);
and UO_937 (O_937,N_24736,N_24460);
nor UO_938 (O_938,N_24412,N_24596);
nor UO_939 (O_939,N_24822,N_24613);
nand UO_940 (O_940,N_24852,N_24816);
and UO_941 (O_941,N_24431,N_24946);
and UO_942 (O_942,N_24544,N_24524);
nand UO_943 (O_943,N_24890,N_24611);
nor UO_944 (O_944,N_24436,N_24413);
nor UO_945 (O_945,N_24725,N_24557);
or UO_946 (O_946,N_24502,N_24498);
nand UO_947 (O_947,N_24769,N_24924);
or UO_948 (O_948,N_24809,N_24818);
and UO_949 (O_949,N_24700,N_24432);
or UO_950 (O_950,N_24670,N_24389);
and UO_951 (O_951,N_24627,N_24966);
nand UO_952 (O_952,N_24641,N_24492);
nand UO_953 (O_953,N_24973,N_24452);
or UO_954 (O_954,N_24926,N_24869);
or UO_955 (O_955,N_24815,N_24527);
or UO_956 (O_956,N_24402,N_24989);
nor UO_957 (O_957,N_24495,N_24918);
nand UO_958 (O_958,N_24849,N_24810);
and UO_959 (O_959,N_24799,N_24663);
and UO_960 (O_960,N_24516,N_24480);
xor UO_961 (O_961,N_24896,N_24999);
and UO_962 (O_962,N_24435,N_24812);
or UO_963 (O_963,N_24588,N_24704);
nand UO_964 (O_964,N_24725,N_24510);
nand UO_965 (O_965,N_24637,N_24797);
or UO_966 (O_966,N_24418,N_24587);
or UO_967 (O_967,N_24645,N_24718);
nand UO_968 (O_968,N_24775,N_24730);
or UO_969 (O_969,N_24555,N_24402);
nor UO_970 (O_970,N_24571,N_24517);
and UO_971 (O_971,N_24523,N_24565);
nand UO_972 (O_972,N_24785,N_24539);
nor UO_973 (O_973,N_24403,N_24810);
nand UO_974 (O_974,N_24850,N_24456);
nand UO_975 (O_975,N_24596,N_24729);
or UO_976 (O_976,N_24775,N_24871);
or UO_977 (O_977,N_24858,N_24636);
nor UO_978 (O_978,N_24630,N_24385);
nor UO_979 (O_979,N_24725,N_24846);
nor UO_980 (O_980,N_24728,N_24632);
nand UO_981 (O_981,N_24924,N_24934);
xor UO_982 (O_982,N_24464,N_24437);
or UO_983 (O_983,N_24874,N_24812);
and UO_984 (O_984,N_24983,N_24656);
or UO_985 (O_985,N_24598,N_24969);
and UO_986 (O_986,N_24851,N_24921);
or UO_987 (O_987,N_24587,N_24915);
nand UO_988 (O_988,N_24974,N_24514);
and UO_989 (O_989,N_24704,N_24640);
nor UO_990 (O_990,N_24919,N_24979);
nand UO_991 (O_991,N_24543,N_24749);
nor UO_992 (O_992,N_24942,N_24393);
and UO_993 (O_993,N_24435,N_24794);
or UO_994 (O_994,N_24600,N_24891);
nand UO_995 (O_995,N_24442,N_24954);
nand UO_996 (O_996,N_24788,N_24921);
xor UO_997 (O_997,N_24442,N_24612);
xnor UO_998 (O_998,N_24428,N_24797);
or UO_999 (O_999,N_24929,N_24541);
and UO_1000 (O_1000,N_24851,N_24958);
xnor UO_1001 (O_1001,N_24559,N_24419);
and UO_1002 (O_1002,N_24397,N_24404);
xnor UO_1003 (O_1003,N_24929,N_24594);
xnor UO_1004 (O_1004,N_24777,N_24632);
nand UO_1005 (O_1005,N_24479,N_24631);
nand UO_1006 (O_1006,N_24940,N_24507);
and UO_1007 (O_1007,N_24820,N_24453);
and UO_1008 (O_1008,N_24975,N_24710);
nor UO_1009 (O_1009,N_24809,N_24624);
nand UO_1010 (O_1010,N_24692,N_24867);
and UO_1011 (O_1011,N_24944,N_24538);
nor UO_1012 (O_1012,N_24933,N_24980);
and UO_1013 (O_1013,N_24657,N_24586);
xnor UO_1014 (O_1014,N_24764,N_24428);
nor UO_1015 (O_1015,N_24805,N_24711);
or UO_1016 (O_1016,N_24511,N_24601);
or UO_1017 (O_1017,N_24781,N_24405);
nand UO_1018 (O_1018,N_24812,N_24986);
nand UO_1019 (O_1019,N_24988,N_24862);
and UO_1020 (O_1020,N_24861,N_24650);
and UO_1021 (O_1021,N_24505,N_24865);
nor UO_1022 (O_1022,N_24558,N_24620);
nor UO_1023 (O_1023,N_24415,N_24623);
xor UO_1024 (O_1024,N_24985,N_24984);
nand UO_1025 (O_1025,N_24435,N_24856);
nor UO_1026 (O_1026,N_24420,N_24517);
nor UO_1027 (O_1027,N_24546,N_24705);
nand UO_1028 (O_1028,N_24817,N_24684);
or UO_1029 (O_1029,N_24390,N_24995);
nand UO_1030 (O_1030,N_24747,N_24744);
xnor UO_1031 (O_1031,N_24443,N_24641);
nand UO_1032 (O_1032,N_24416,N_24574);
nand UO_1033 (O_1033,N_24486,N_24910);
and UO_1034 (O_1034,N_24909,N_24974);
nor UO_1035 (O_1035,N_24518,N_24859);
nor UO_1036 (O_1036,N_24598,N_24505);
nor UO_1037 (O_1037,N_24855,N_24786);
or UO_1038 (O_1038,N_24690,N_24908);
nand UO_1039 (O_1039,N_24380,N_24717);
nor UO_1040 (O_1040,N_24430,N_24561);
xnor UO_1041 (O_1041,N_24960,N_24553);
or UO_1042 (O_1042,N_24442,N_24833);
xor UO_1043 (O_1043,N_24557,N_24385);
nand UO_1044 (O_1044,N_24478,N_24586);
nand UO_1045 (O_1045,N_24924,N_24764);
and UO_1046 (O_1046,N_24523,N_24509);
nor UO_1047 (O_1047,N_24644,N_24631);
xnor UO_1048 (O_1048,N_24801,N_24397);
nand UO_1049 (O_1049,N_24754,N_24758);
or UO_1050 (O_1050,N_24975,N_24977);
or UO_1051 (O_1051,N_24535,N_24974);
nand UO_1052 (O_1052,N_24680,N_24753);
nor UO_1053 (O_1053,N_24714,N_24917);
nor UO_1054 (O_1054,N_24393,N_24816);
xor UO_1055 (O_1055,N_24505,N_24393);
nand UO_1056 (O_1056,N_24939,N_24550);
or UO_1057 (O_1057,N_24891,N_24560);
or UO_1058 (O_1058,N_24679,N_24620);
or UO_1059 (O_1059,N_24377,N_24759);
nand UO_1060 (O_1060,N_24955,N_24748);
nor UO_1061 (O_1061,N_24909,N_24562);
or UO_1062 (O_1062,N_24560,N_24430);
nand UO_1063 (O_1063,N_24518,N_24435);
nand UO_1064 (O_1064,N_24645,N_24936);
nand UO_1065 (O_1065,N_24714,N_24442);
and UO_1066 (O_1066,N_24825,N_24883);
xor UO_1067 (O_1067,N_24574,N_24591);
and UO_1068 (O_1068,N_24400,N_24475);
or UO_1069 (O_1069,N_24782,N_24757);
or UO_1070 (O_1070,N_24560,N_24745);
nand UO_1071 (O_1071,N_24681,N_24866);
xor UO_1072 (O_1072,N_24866,N_24540);
and UO_1073 (O_1073,N_24483,N_24976);
nor UO_1074 (O_1074,N_24426,N_24763);
nor UO_1075 (O_1075,N_24842,N_24701);
and UO_1076 (O_1076,N_24502,N_24436);
and UO_1077 (O_1077,N_24909,N_24384);
nand UO_1078 (O_1078,N_24427,N_24828);
xnor UO_1079 (O_1079,N_24425,N_24431);
nor UO_1080 (O_1080,N_24389,N_24681);
or UO_1081 (O_1081,N_24835,N_24760);
and UO_1082 (O_1082,N_24614,N_24568);
or UO_1083 (O_1083,N_24473,N_24945);
or UO_1084 (O_1084,N_24880,N_24410);
xor UO_1085 (O_1085,N_24672,N_24937);
xor UO_1086 (O_1086,N_24906,N_24891);
or UO_1087 (O_1087,N_24850,N_24626);
nor UO_1088 (O_1088,N_24962,N_24643);
nand UO_1089 (O_1089,N_24953,N_24723);
xnor UO_1090 (O_1090,N_24786,N_24806);
nand UO_1091 (O_1091,N_24726,N_24675);
xor UO_1092 (O_1092,N_24433,N_24543);
or UO_1093 (O_1093,N_24924,N_24424);
nor UO_1094 (O_1094,N_24917,N_24655);
and UO_1095 (O_1095,N_24945,N_24795);
nand UO_1096 (O_1096,N_24375,N_24696);
or UO_1097 (O_1097,N_24400,N_24438);
nand UO_1098 (O_1098,N_24457,N_24595);
and UO_1099 (O_1099,N_24914,N_24696);
nand UO_1100 (O_1100,N_24502,N_24381);
nand UO_1101 (O_1101,N_24780,N_24632);
or UO_1102 (O_1102,N_24612,N_24849);
nor UO_1103 (O_1103,N_24777,N_24891);
nor UO_1104 (O_1104,N_24826,N_24883);
nand UO_1105 (O_1105,N_24904,N_24955);
nand UO_1106 (O_1106,N_24948,N_24558);
nor UO_1107 (O_1107,N_24798,N_24550);
nor UO_1108 (O_1108,N_24485,N_24768);
nand UO_1109 (O_1109,N_24726,N_24858);
or UO_1110 (O_1110,N_24924,N_24827);
xnor UO_1111 (O_1111,N_24679,N_24626);
xnor UO_1112 (O_1112,N_24541,N_24583);
nand UO_1113 (O_1113,N_24777,N_24778);
and UO_1114 (O_1114,N_24484,N_24573);
or UO_1115 (O_1115,N_24965,N_24682);
nor UO_1116 (O_1116,N_24388,N_24959);
and UO_1117 (O_1117,N_24777,N_24766);
nand UO_1118 (O_1118,N_24972,N_24794);
xnor UO_1119 (O_1119,N_24893,N_24375);
nand UO_1120 (O_1120,N_24970,N_24754);
nand UO_1121 (O_1121,N_24617,N_24415);
or UO_1122 (O_1122,N_24882,N_24852);
nand UO_1123 (O_1123,N_24586,N_24616);
and UO_1124 (O_1124,N_24649,N_24934);
xnor UO_1125 (O_1125,N_24506,N_24799);
or UO_1126 (O_1126,N_24701,N_24916);
xor UO_1127 (O_1127,N_24631,N_24906);
xor UO_1128 (O_1128,N_24425,N_24890);
xnor UO_1129 (O_1129,N_24969,N_24544);
nand UO_1130 (O_1130,N_24958,N_24809);
and UO_1131 (O_1131,N_24492,N_24650);
or UO_1132 (O_1132,N_24490,N_24576);
xnor UO_1133 (O_1133,N_24515,N_24388);
or UO_1134 (O_1134,N_24569,N_24575);
nand UO_1135 (O_1135,N_24783,N_24931);
nand UO_1136 (O_1136,N_24834,N_24394);
nand UO_1137 (O_1137,N_24656,N_24499);
or UO_1138 (O_1138,N_24746,N_24490);
or UO_1139 (O_1139,N_24720,N_24680);
xor UO_1140 (O_1140,N_24779,N_24456);
nor UO_1141 (O_1141,N_24786,N_24981);
and UO_1142 (O_1142,N_24473,N_24977);
nand UO_1143 (O_1143,N_24411,N_24527);
nand UO_1144 (O_1144,N_24541,N_24860);
nand UO_1145 (O_1145,N_24575,N_24620);
nand UO_1146 (O_1146,N_24479,N_24901);
xnor UO_1147 (O_1147,N_24467,N_24869);
and UO_1148 (O_1148,N_24474,N_24697);
nor UO_1149 (O_1149,N_24595,N_24638);
or UO_1150 (O_1150,N_24445,N_24410);
xor UO_1151 (O_1151,N_24743,N_24884);
nand UO_1152 (O_1152,N_24553,N_24966);
nand UO_1153 (O_1153,N_24731,N_24796);
nand UO_1154 (O_1154,N_24661,N_24851);
or UO_1155 (O_1155,N_24983,N_24674);
nor UO_1156 (O_1156,N_24751,N_24420);
and UO_1157 (O_1157,N_24854,N_24849);
nand UO_1158 (O_1158,N_24782,N_24467);
nand UO_1159 (O_1159,N_24933,N_24519);
and UO_1160 (O_1160,N_24653,N_24586);
nor UO_1161 (O_1161,N_24498,N_24589);
and UO_1162 (O_1162,N_24404,N_24629);
nor UO_1163 (O_1163,N_24988,N_24418);
xnor UO_1164 (O_1164,N_24919,N_24989);
nor UO_1165 (O_1165,N_24867,N_24514);
nand UO_1166 (O_1166,N_24660,N_24444);
and UO_1167 (O_1167,N_24824,N_24488);
nor UO_1168 (O_1168,N_24528,N_24704);
and UO_1169 (O_1169,N_24573,N_24799);
and UO_1170 (O_1170,N_24490,N_24561);
nand UO_1171 (O_1171,N_24826,N_24814);
and UO_1172 (O_1172,N_24986,N_24437);
and UO_1173 (O_1173,N_24589,N_24879);
or UO_1174 (O_1174,N_24919,N_24917);
nor UO_1175 (O_1175,N_24707,N_24654);
or UO_1176 (O_1176,N_24695,N_24813);
nand UO_1177 (O_1177,N_24410,N_24572);
nand UO_1178 (O_1178,N_24763,N_24600);
nor UO_1179 (O_1179,N_24971,N_24871);
or UO_1180 (O_1180,N_24679,N_24514);
nand UO_1181 (O_1181,N_24746,N_24694);
and UO_1182 (O_1182,N_24891,N_24685);
nor UO_1183 (O_1183,N_24576,N_24612);
and UO_1184 (O_1184,N_24403,N_24600);
nand UO_1185 (O_1185,N_24749,N_24884);
and UO_1186 (O_1186,N_24593,N_24776);
or UO_1187 (O_1187,N_24892,N_24471);
nand UO_1188 (O_1188,N_24822,N_24435);
nor UO_1189 (O_1189,N_24702,N_24564);
and UO_1190 (O_1190,N_24916,N_24448);
nor UO_1191 (O_1191,N_24578,N_24979);
or UO_1192 (O_1192,N_24630,N_24599);
nor UO_1193 (O_1193,N_24704,N_24536);
nor UO_1194 (O_1194,N_24922,N_24795);
xnor UO_1195 (O_1195,N_24757,N_24687);
nand UO_1196 (O_1196,N_24575,N_24622);
or UO_1197 (O_1197,N_24590,N_24887);
or UO_1198 (O_1198,N_24416,N_24378);
nand UO_1199 (O_1199,N_24987,N_24537);
or UO_1200 (O_1200,N_24644,N_24862);
xnor UO_1201 (O_1201,N_24488,N_24692);
and UO_1202 (O_1202,N_24891,N_24838);
and UO_1203 (O_1203,N_24824,N_24847);
or UO_1204 (O_1204,N_24591,N_24839);
or UO_1205 (O_1205,N_24794,N_24933);
nand UO_1206 (O_1206,N_24567,N_24814);
xor UO_1207 (O_1207,N_24415,N_24466);
or UO_1208 (O_1208,N_24672,N_24830);
or UO_1209 (O_1209,N_24391,N_24723);
and UO_1210 (O_1210,N_24506,N_24438);
and UO_1211 (O_1211,N_24650,N_24666);
or UO_1212 (O_1212,N_24879,N_24797);
or UO_1213 (O_1213,N_24857,N_24814);
nand UO_1214 (O_1214,N_24902,N_24744);
or UO_1215 (O_1215,N_24454,N_24410);
nor UO_1216 (O_1216,N_24648,N_24851);
nand UO_1217 (O_1217,N_24908,N_24463);
nor UO_1218 (O_1218,N_24464,N_24951);
nand UO_1219 (O_1219,N_24470,N_24860);
and UO_1220 (O_1220,N_24526,N_24673);
and UO_1221 (O_1221,N_24751,N_24970);
nand UO_1222 (O_1222,N_24481,N_24826);
nand UO_1223 (O_1223,N_24687,N_24554);
nand UO_1224 (O_1224,N_24508,N_24964);
nand UO_1225 (O_1225,N_24666,N_24592);
and UO_1226 (O_1226,N_24826,N_24764);
nand UO_1227 (O_1227,N_24855,N_24543);
or UO_1228 (O_1228,N_24404,N_24576);
and UO_1229 (O_1229,N_24780,N_24681);
nand UO_1230 (O_1230,N_24778,N_24794);
nand UO_1231 (O_1231,N_24611,N_24493);
nand UO_1232 (O_1232,N_24706,N_24737);
nor UO_1233 (O_1233,N_24755,N_24971);
or UO_1234 (O_1234,N_24469,N_24966);
xnor UO_1235 (O_1235,N_24953,N_24606);
and UO_1236 (O_1236,N_24395,N_24660);
nand UO_1237 (O_1237,N_24394,N_24613);
or UO_1238 (O_1238,N_24839,N_24951);
nand UO_1239 (O_1239,N_24996,N_24801);
nor UO_1240 (O_1240,N_24860,N_24736);
and UO_1241 (O_1241,N_24447,N_24511);
xnor UO_1242 (O_1242,N_24814,N_24757);
xnor UO_1243 (O_1243,N_24900,N_24866);
nand UO_1244 (O_1244,N_24375,N_24934);
xnor UO_1245 (O_1245,N_24976,N_24830);
nand UO_1246 (O_1246,N_24856,N_24807);
or UO_1247 (O_1247,N_24860,N_24895);
or UO_1248 (O_1248,N_24813,N_24617);
or UO_1249 (O_1249,N_24971,N_24816);
nor UO_1250 (O_1250,N_24694,N_24471);
nand UO_1251 (O_1251,N_24894,N_24395);
nor UO_1252 (O_1252,N_24733,N_24799);
nand UO_1253 (O_1253,N_24712,N_24938);
nor UO_1254 (O_1254,N_24773,N_24612);
and UO_1255 (O_1255,N_24885,N_24588);
nor UO_1256 (O_1256,N_24971,N_24678);
or UO_1257 (O_1257,N_24422,N_24590);
nand UO_1258 (O_1258,N_24493,N_24593);
nor UO_1259 (O_1259,N_24444,N_24789);
nor UO_1260 (O_1260,N_24996,N_24463);
nand UO_1261 (O_1261,N_24623,N_24636);
or UO_1262 (O_1262,N_24898,N_24475);
or UO_1263 (O_1263,N_24573,N_24742);
nor UO_1264 (O_1264,N_24613,N_24468);
and UO_1265 (O_1265,N_24863,N_24927);
or UO_1266 (O_1266,N_24668,N_24847);
nand UO_1267 (O_1267,N_24594,N_24486);
nor UO_1268 (O_1268,N_24670,N_24850);
nor UO_1269 (O_1269,N_24376,N_24993);
nand UO_1270 (O_1270,N_24631,N_24578);
or UO_1271 (O_1271,N_24655,N_24703);
nor UO_1272 (O_1272,N_24634,N_24605);
nand UO_1273 (O_1273,N_24376,N_24871);
or UO_1274 (O_1274,N_24540,N_24603);
nor UO_1275 (O_1275,N_24526,N_24770);
nand UO_1276 (O_1276,N_24917,N_24563);
nand UO_1277 (O_1277,N_24378,N_24805);
or UO_1278 (O_1278,N_24586,N_24757);
or UO_1279 (O_1279,N_24756,N_24957);
nand UO_1280 (O_1280,N_24586,N_24416);
or UO_1281 (O_1281,N_24802,N_24692);
nor UO_1282 (O_1282,N_24467,N_24881);
nand UO_1283 (O_1283,N_24604,N_24889);
nand UO_1284 (O_1284,N_24468,N_24685);
nand UO_1285 (O_1285,N_24588,N_24406);
or UO_1286 (O_1286,N_24633,N_24406);
and UO_1287 (O_1287,N_24720,N_24969);
nor UO_1288 (O_1288,N_24820,N_24664);
nand UO_1289 (O_1289,N_24772,N_24459);
nor UO_1290 (O_1290,N_24672,N_24829);
nand UO_1291 (O_1291,N_24822,N_24419);
xor UO_1292 (O_1292,N_24492,N_24796);
and UO_1293 (O_1293,N_24480,N_24742);
and UO_1294 (O_1294,N_24475,N_24992);
xnor UO_1295 (O_1295,N_24412,N_24407);
and UO_1296 (O_1296,N_24762,N_24533);
xnor UO_1297 (O_1297,N_24891,N_24723);
nand UO_1298 (O_1298,N_24560,N_24515);
nor UO_1299 (O_1299,N_24765,N_24618);
and UO_1300 (O_1300,N_24687,N_24766);
and UO_1301 (O_1301,N_24666,N_24904);
or UO_1302 (O_1302,N_24410,N_24847);
nor UO_1303 (O_1303,N_24410,N_24820);
and UO_1304 (O_1304,N_24519,N_24838);
and UO_1305 (O_1305,N_24995,N_24736);
or UO_1306 (O_1306,N_24999,N_24469);
and UO_1307 (O_1307,N_24497,N_24793);
nor UO_1308 (O_1308,N_24611,N_24536);
xor UO_1309 (O_1309,N_24886,N_24985);
nor UO_1310 (O_1310,N_24896,N_24410);
nor UO_1311 (O_1311,N_24723,N_24454);
and UO_1312 (O_1312,N_24554,N_24900);
nand UO_1313 (O_1313,N_24424,N_24742);
nand UO_1314 (O_1314,N_24729,N_24467);
or UO_1315 (O_1315,N_24413,N_24483);
nand UO_1316 (O_1316,N_24725,N_24533);
nand UO_1317 (O_1317,N_24511,N_24476);
or UO_1318 (O_1318,N_24752,N_24637);
nand UO_1319 (O_1319,N_24947,N_24539);
nand UO_1320 (O_1320,N_24524,N_24735);
nand UO_1321 (O_1321,N_24581,N_24501);
nor UO_1322 (O_1322,N_24423,N_24664);
and UO_1323 (O_1323,N_24980,N_24821);
and UO_1324 (O_1324,N_24712,N_24651);
and UO_1325 (O_1325,N_24819,N_24401);
or UO_1326 (O_1326,N_24942,N_24420);
or UO_1327 (O_1327,N_24817,N_24888);
xnor UO_1328 (O_1328,N_24603,N_24831);
or UO_1329 (O_1329,N_24939,N_24382);
and UO_1330 (O_1330,N_24853,N_24421);
or UO_1331 (O_1331,N_24573,N_24387);
and UO_1332 (O_1332,N_24501,N_24830);
and UO_1333 (O_1333,N_24433,N_24576);
nor UO_1334 (O_1334,N_24574,N_24842);
and UO_1335 (O_1335,N_24726,N_24551);
nor UO_1336 (O_1336,N_24651,N_24711);
nor UO_1337 (O_1337,N_24489,N_24415);
nor UO_1338 (O_1338,N_24563,N_24431);
and UO_1339 (O_1339,N_24636,N_24421);
nand UO_1340 (O_1340,N_24818,N_24861);
nor UO_1341 (O_1341,N_24771,N_24649);
and UO_1342 (O_1342,N_24784,N_24856);
and UO_1343 (O_1343,N_24587,N_24453);
nor UO_1344 (O_1344,N_24981,N_24756);
or UO_1345 (O_1345,N_24398,N_24669);
nor UO_1346 (O_1346,N_24930,N_24433);
nand UO_1347 (O_1347,N_24815,N_24379);
or UO_1348 (O_1348,N_24889,N_24637);
or UO_1349 (O_1349,N_24414,N_24588);
or UO_1350 (O_1350,N_24859,N_24607);
nor UO_1351 (O_1351,N_24445,N_24525);
or UO_1352 (O_1352,N_24411,N_24438);
nand UO_1353 (O_1353,N_24424,N_24648);
xnor UO_1354 (O_1354,N_24973,N_24457);
nor UO_1355 (O_1355,N_24550,N_24783);
or UO_1356 (O_1356,N_24863,N_24618);
nand UO_1357 (O_1357,N_24398,N_24756);
nor UO_1358 (O_1358,N_24650,N_24710);
nand UO_1359 (O_1359,N_24763,N_24735);
nor UO_1360 (O_1360,N_24940,N_24930);
or UO_1361 (O_1361,N_24611,N_24396);
nand UO_1362 (O_1362,N_24783,N_24828);
nand UO_1363 (O_1363,N_24679,N_24821);
and UO_1364 (O_1364,N_24844,N_24666);
or UO_1365 (O_1365,N_24380,N_24866);
and UO_1366 (O_1366,N_24665,N_24431);
or UO_1367 (O_1367,N_24478,N_24466);
xnor UO_1368 (O_1368,N_24743,N_24643);
and UO_1369 (O_1369,N_24826,N_24774);
nor UO_1370 (O_1370,N_24661,N_24646);
nor UO_1371 (O_1371,N_24921,N_24445);
or UO_1372 (O_1372,N_24662,N_24390);
nor UO_1373 (O_1373,N_24578,N_24390);
or UO_1374 (O_1374,N_24624,N_24604);
nand UO_1375 (O_1375,N_24945,N_24774);
nor UO_1376 (O_1376,N_24961,N_24933);
nand UO_1377 (O_1377,N_24657,N_24899);
or UO_1378 (O_1378,N_24740,N_24396);
or UO_1379 (O_1379,N_24578,N_24416);
and UO_1380 (O_1380,N_24495,N_24833);
xnor UO_1381 (O_1381,N_24707,N_24586);
or UO_1382 (O_1382,N_24499,N_24769);
or UO_1383 (O_1383,N_24739,N_24609);
or UO_1384 (O_1384,N_24655,N_24791);
and UO_1385 (O_1385,N_24998,N_24534);
or UO_1386 (O_1386,N_24584,N_24998);
or UO_1387 (O_1387,N_24513,N_24960);
nand UO_1388 (O_1388,N_24495,N_24528);
nor UO_1389 (O_1389,N_24957,N_24764);
nand UO_1390 (O_1390,N_24910,N_24540);
xor UO_1391 (O_1391,N_24870,N_24792);
nor UO_1392 (O_1392,N_24725,N_24988);
nor UO_1393 (O_1393,N_24993,N_24637);
nand UO_1394 (O_1394,N_24882,N_24868);
or UO_1395 (O_1395,N_24742,N_24763);
nand UO_1396 (O_1396,N_24559,N_24409);
and UO_1397 (O_1397,N_24893,N_24810);
nand UO_1398 (O_1398,N_24695,N_24522);
and UO_1399 (O_1399,N_24968,N_24398);
and UO_1400 (O_1400,N_24478,N_24896);
xor UO_1401 (O_1401,N_24891,N_24573);
or UO_1402 (O_1402,N_24840,N_24817);
nor UO_1403 (O_1403,N_24456,N_24686);
nand UO_1404 (O_1404,N_24441,N_24429);
nor UO_1405 (O_1405,N_24627,N_24717);
nand UO_1406 (O_1406,N_24494,N_24914);
xnor UO_1407 (O_1407,N_24537,N_24908);
nor UO_1408 (O_1408,N_24615,N_24643);
nor UO_1409 (O_1409,N_24771,N_24609);
nor UO_1410 (O_1410,N_24702,N_24496);
nor UO_1411 (O_1411,N_24740,N_24938);
and UO_1412 (O_1412,N_24596,N_24501);
nor UO_1413 (O_1413,N_24420,N_24723);
nand UO_1414 (O_1414,N_24509,N_24875);
and UO_1415 (O_1415,N_24971,N_24798);
xor UO_1416 (O_1416,N_24905,N_24517);
nor UO_1417 (O_1417,N_24523,N_24498);
or UO_1418 (O_1418,N_24416,N_24951);
or UO_1419 (O_1419,N_24509,N_24539);
and UO_1420 (O_1420,N_24946,N_24838);
nor UO_1421 (O_1421,N_24554,N_24988);
nor UO_1422 (O_1422,N_24486,N_24859);
and UO_1423 (O_1423,N_24684,N_24404);
or UO_1424 (O_1424,N_24774,N_24939);
xnor UO_1425 (O_1425,N_24733,N_24666);
nor UO_1426 (O_1426,N_24383,N_24609);
nand UO_1427 (O_1427,N_24573,N_24637);
and UO_1428 (O_1428,N_24985,N_24902);
or UO_1429 (O_1429,N_24380,N_24965);
or UO_1430 (O_1430,N_24946,N_24673);
or UO_1431 (O_1431,N_24503,N_24995);
xnor UO_1432 (O_1432,N_24447,N_24892);
xor UO_1433 (O_1433,N_24831,N_24713);
and UO_1434 (O_1434,N_24751,N_24562);
nor UO_1435 (O_1435,N_24515,N_24571);
nand UO_1436 (O_1436,N_24559,N_24774);
or UO_1437 (O_1437,N_24681,N_24889);
and UO_1438 (O_1438,N_24737,N_24506);
nand UO_1439 (O_1439,N_24405,N_24989);
and UO_1440 (O_1440,N_24936,N_24383);
or UO_1441 (O_1441,N_24940,N_24949);
and UO_1442 (O_1442,N_24628,N_24850);
and UO_1443 (O_1443,N_24955,N_24563);
nor UO_1444 (O_1444,N_24825,N_24431);
nand UO_1445 (O_1445,N_24916,N_24435);
and UO_1446 (O_1446,N_24931,N_24930);
or UO_1447 (O_1447,N_24858,N_24380);
nand UO_1448 (O_1448,N_24846,N_24918);
or UO_1449 (O_1449,N_24631,N_24747);
and UO_1450 (O_1450,N_24400,N_24507);
nor UO_1451 (O_1451,N_24971,N_24610);
and UO_1452 (O_1452,N_24625,N_24699);
and UO_1453 (O_1453,N_24691,N_24548);
or UO_1454 (O_1454,N_24585,N_24668);
or UO_1455 (O_1455,N_24681,N_24979);
and UO_1456 (O_1456,N_24534,N_24897);
and UO_1457 (O_1457,N_24578,N_24854);
xnor UO_1458 (O_1458,N_24749,N_24844);
and UO_1459 (O_1459,N_24658,N_24452);
nand UO_1460 (O_1460,N_24841,N_24600);
nor UO_1461 (O_1461,N_24594,N_24997);
or UO_1462 (O_1462,N_24548,N_24661);
and UO_1463 (O_1463,N_24940,N_24635);
nand UO_1464 (O_1464,N_24849,N_24914);
nor UO_1465 (O_1465,N_24948,N_24995);
xnor UO_1466 (O_1466,N_24688,N_24926);
or UO_1467 (O_1467,N_24676,N_24407);
or UO_1468 (O_1468,N_24759,N_24552);
nand UO_1469 (O_1469,N_24439,N_24402);
xnor UO_1470 (O_1470,N_24749,N_24906);
nand UO_1471 (O_1471,N_24799,N_24875);
and UO_1472 (O_1472,N_24649,N_24863);
nor UO_1473 (O_1473,N_24690,N_24454);
nand UO_1474 (O_1474,N_24572,N_24954);
and UO_1475 (O_1475,N_24802,N_24737);
nor UO_1476 (O_1476,N_24395,N_24768);
or UO_1477 (O_1477,N_24538,N_24994);
nand UO_1478 (O_1478,N_24676,N_24636);
or UO_1479 (O_1479,N_24821,N_24417);
nand UO_1480 (O_1480,N_24461,N_24777);
or UO_1481 (O_1481,N_24451,N_24864);
and UO_1482 (O_1482,N_24959,N_24822);
and UO_1483 (O_1483,N_24531,N_24934);
nor UO_1484 (O_1484,N_24394,N_24697);
nand UO_1485 (O_1485,N_24809,N_24857);
nor UO_1486 (O_1486,N_24999,N_24400);
xor UO_1487 (O_1487,N_24645,N_24907);
nor UO_1488 (O_1488,N_24637,N_24902);
and UO_1489 (O_1489,N_24425,N_24477);
or UO_1490 (O_1490,N_24683,N_24727);
or UO_1491 (O_1491,N_24902,N_24386);
and UO_1492 (O_1492,N_24378,N_24551);
or UO_1493 (O_1493,N_24935,N_24949);
nand UO_1494 (O_1494,N_24566,N_24376);
nor UO_1495 (O_1495,N_24904,N_24650);
or UO_1496 (O_1496,N_24774,N_24725);
nand UO_1497 (O_1497,N_24392,N_24506);
nor UO_1498 (O_1498,N_24608,N_24515);
nand UO_1499 (O_1499,N_24513,N_24645);
nor UO_1500 (O_1500,N_24620,N_24978);
and UO_1501 (O_1501,N_24803,N_24862);
nor UO_1502 (O_1502,N_24922,N_24718);
and UO_1503 (O_1503,N_24681,N_24833);
or UO_1504 (O_1504,N_24938,N_24923);
and UO_1505 (O_1505,N_24473,N_24850);
xor UO_1506 (O_1506,N_24811,N_24663);
or UO_1507 (O_1507,N_24934,N_24955);
and UO_1508 (O_1508,N_24467,N_24599);
nor UO_1509 (O_1509,N_24780,N_24501);
or UO_1510 (O_1510,N_24817,N_24693);
and UO_1511 (O_1511,N_24535,N_24662);
nand UO_1512 (O_1512,N_24956,N_24504);
and UO_1513 (O_1513,N_24683,N_24472);
nand UO_1514 (O_1514,N_24838,N_24748);
and UO_1515 (O_1515,N_24972,N_24493);
and UO_1516 (O_1516,N_24785,N_24774);
nor UO_1517 (O_1517,N_24821,N_24447);
and UO_1518 (O_1518,N_24893,N_24618);
or UO_1519 (O_1519,N_24687,N_24967);
and UO_1520 (O_1520,N_24943,N_24734);
or UO_1521 (O_1521,N_24788,N_24404);
nor UO_1522 (O_1522,N_24521,N_24986);
nor UO_1523 (O_1523,N_24616,N_24901);
and UO_1524 (O_1524,N_24642,N_24561);
nor UO_1525 (O_1525,N_24699,N_24878);
nand UO_1526 (O_1526,N_24559,N_24776);
nand UO_1527 (O_1527,N_24377,N_24478);
or UO_1528 (O_1528,N_24593,N_24668);
or UO_1529 (O_1529,N_24670,N_24663);
and UO_1530 (O_1530,N_24599,N_24560);
nand UO_1531 (O_1531,N_24643,N_24815);
nor UO_1532 (O_1532,N_24827,N_24491);
and UO_1533 (O_1533,N_24720,N_24589);
and UO_1534 (O_1534,N_24545,N_24967);
and UO_1535 (O_1535,N_24886,N_24839);
nor UO_1536 (O_1536,N_24419,N_24633);
or UO_1537 (O_1537,N_24489,N_24881);
nand UO_1538 (O_1538,N_24809,N_24391);
and UO_1539 (O_1539,N_24669,N_24482);
nand UO_1540 (O_1540,N_24569,N_24727);
nor UO_1541 (O_1541,N_24530,N_24835);
nand UO_1542 (O_1542,N_24920,N_24719);
and UO_1543 (O_1543,N_24414,N_24948);
nor UO_1544 (O_1544,N_24800,N_24726);
nand UO_1545 (O_1545,N_24860,N_24832);
or UO_1546 (O_1546,N_24800,N_24938);
nor UO_1547 (O_1547,N_24777,N_24761);
or UO_1548 (O_1548,N_24425,N_24869);
or UO_1549 (O_1549,N_24402,N_24895);
nor UO_1550 (O_1550,N_24816,N_24905);
nand UO_1551 (O_1551,N_24775,N_24729);
xor UO_1552 (O_1552,N_24441,N_24666);
and UO_1553 (O_1553,N_24702,N_24405);
and UO_1554 (O_1554,N_24858,N_24803);
and UO_1555 (O_1555,N_24560,N_24494);
or UO_1556 (O_1556,N_24727,N_24604);
nand UO_1557 (O_1557,N_24519,N_24435);
xor UO_1558 (O_1558,N_24415,N_24924);
or UO_1559 (O_1559,N_24635,N_24778);
and UO_1560 (O_1560,N_24845,N_24765);
or UO_1561 (O_1561,N_24383,N_24867);
or UO_1562 (O_1562,N_24510,N_24518);
nor UO_1563 (O_1563,N_24785,N_24447);
or UO_1564 (O_1564,N_24412,N_24974);
or UO_1565 (O_1565,N_24610,N_24481);
nor UO_1566 (O_1566,N_24904,N_24391);
nand UO_1567 (O_1567,N_24542,N_24953);
or UO_1568 (O_1568,N_24664,N_24430);
nand UO_1569 (O_1569,N_24525,N_24522);
nor UO_1570 (O_1570,N_24633,N_24590);
nand UO_1571 (O_1571,N_24869,N_24439);
nand UO_1572 (O_1572,N_24797,N_24510);
nor UO_1573 (O_1573,N_24742,N_24797);
or UO_1574 (O_1574,N_24589,N_24931);
and UO_1575 (O_1575,N_24411,N_24801);
or UO_1576 (O_1576,N_24575,N_24872);
or UO_1577 (O_1577,N_24405,N_24909);
xor UO_1578 (O_1578,N_24687,N_24838);
and UO_1579 (O_1579,N_24438,N_24868);
and UO_1580 (O_1580,N_24881,N_24920);
or UO_1581 (O_1581,N_24488,N_24849);
nor UO_1582 (O_1582,N_24730,N_24541);
nand UO_1583 (O_1583,N_24933,N_24969);
and UO_1584 (O_1584,N_24880,N_24845);
and UO_1585 (O_1585,N_24978,N_24599);
nor UO_1586 (O_1586,N_24383,N_24865);
nor UO_1587 (O_1587,N_24858,N_24454);
nor UO_1588 (O_1588,N_24983,N_24755);
nor UO_1589 (O_1589,N_24522,N_24978);
or UO_1590 (O_1590,N_24800,N_24654);
or UO_1591 (O_1591,N_24844,N_24643);
nor UO_1592 (O_1592,N_24951,N_24976);
and UO_1593 (O_1593,N_24608,N_24787);
and UO_1594 (O_1594,N_24478,N_24597);
nand UO_1595 (O_1595,N_24508,N_24592);
or UO_1596 (O_1596,N_24888,N_24381);
and UO_1597 (O_1597,N_24585,N_24822);
or UO_1598 (O_1598,N_24393,N_24713);
xnor UO_1599 (O_1599,N_24717,N_24795);
and UO_1600 (O_1600,N_24517,N_24748);
nand UO_1601 (O_1601,N_24460,N_24449);
nand UO_1602 (O_1602,N_24500,N_24570);
and UO_1603 (O_1603,N_24966,N_24640);
nor UO_1604 (O_1604,N_24836,N_24466);
xnor UO_1605 (O_1605,N_24724,N_24630);
nor UO_1606 (O_1606,N_24901,N_24693);
nand UO_1607 (O_1607,N_24639,N_24642);
or UO_1608 (O_1608,N_24402,N_24944);
and UO_1609 (O_1609,N_24618,N_24642);
nor UO_1610 (O_1610,N_24565,N_24806);
nor UO_1611 (O_1611,N_24875,N_24489);
nand UO_1612 (O_1612,N_24385,N_24939);
nor UO_1613 (O_1613,N_24712,N_24529);
or UO_1614 (O_1614,N_24978,N_24608);
or UO_1615 (O_1615,N_24665,N_24563);
nand UO_1616 (O_1616,N_24409,N_24677);
nor UO_1617 (O_1617,N_24954,N_24600);
nor UO_1618 (O_1618,N_24530,N_24632);
or UO_1619 (O_1619,N_24579,N_24811);
and UO_1620 (O_1620,N_24887,N_24607);
or UO_1621 (O_1621,N_24462,N_24840);
or UO_1622 (O_1622,N_24956,N_24894);
and UO_1623 (O_1623,N_24932,N_24636);
or UO_1624 (O_1624,N_24915,N_24511);
and UO_1625 (O_1625,N_24489,N_24385);
nor UO_1626 (O_1626,N_24584,N_24473);
nand UO_1627 (O_1627,N_24842,N_24967);
nand UO_1628 (O_1628,N_24557,N_24931);
or UO_1629 (O_1629,N_24693,N_24685);
nor UO_1630 (O_1630,N_24462,N_24834);
nor UO_1631 (O_1631,N_24966,N_24386);
nand UO_1632 (O_1632,N_24772,N_24842);
and UO_1633 (O_1633,N_24564,N_24922);
or UO_1634 (O_1634,N_24989,N_24825);
nand UO_1635 (O_1635,N_24935,N_24904);
nand UO_1636 (O_1636,N_24837,N_24479);
or UO_1637 (O_1637,N_24865,N_24798);
nor UO_1638 (O_1638,N_24482,N_24598);
nand UO_1639 (O_1639,N_24541,N_24627);
or UO_1640 (O_1640,N_24431,N_24463);
nand UO_1641 (O_1641,N_24820,N_24632);
and UO_1642 (O_1642,N_24902,N_24863);
or UO_1643 (O_1643,N_24388,N_24736);
or UO_1644 (O_1644,N_24377,N_24861);
and UO_1645 (O_1645,N_24971,N_24508);
nor UO_1646 (O_1646,N_24726,N_24986);
nor UO_1647 (O_1647,N_24950,N_24988);
xnor UO_1648 (O_1648,N_24771,N_24557);
nor UO_1649 (O_1649,N_24793,N_24462);
nand UO_1650 (O_1650,N_24756,N_24940);
nor UO_1651 (O_1651,N_24456,N_24941);
nor UO_1652 (O_1652,N_24891,N_24553);
and UO_1653 (O_1653,N_24689,N_24841);
or UO_1654 (O_1654,N_24880,N_24945);
xor UO_1655 (O_1655,N_24626,N_24814);
or UO_1656 (O_1656,N_24899,N_24804);
nand UO_1657 (O_1657,N_24771,N_24865);
nand UO_1658 (O_1658,N_24547,N_24737);
nand UO_1659 (O_1659,N_24847,N_24767);
or UO_1660 (O_1660,N_24573,N_24733);
nand UO_1661 (O_1661,N_24634,N_24697);
xnor UO_1662 (O_1662,N_24914,N_24643);
nor UO_1663 (O_1663,N_24461,N_24637);
and UO_1664 (O_1664,N_24839,N_24751);
nand UO_1665 (O_1665,N_24586,N_24827);
or UO_1666 (O_1666,N_24733,N_24911);
or UO_1667 (O_1667,N_24467,N_24549);
nand UO_1668 (O_1668,N_24536,N_24944);
nand UO_1669 (O_1669,N_24800,N_24651);
and UO_1670 (O_1670,N_24538,N_24517);
xnor UO_1671 (O_1671,N_24543,N_24813);
xor UO_1672 (O_1672,N_24956,N_24397);
nor UO_1673 (O_1673,N_24531,N_24701);
nor UO_1674 (O_1674,N_24581,N_24594);
or UO_1675 (O_1675,N_24458,N_24481);
nand UO_1676 (O_1676,N_24461,N_24505);
or UO_1677 (O_1677,N_24589,N_24831);
and UO_1678 (O_1678,N_24399,N_24383);
and UO_1679 (O_1679,N_24433,N_24511);
nand UO_1680 (O_1680,N_24482,N_24402);
nor UO_1681 (O_1681,N_24591,N_24495);
or UO_1682 (O_1682,N_24760,N_24916);
and UO_1683 (O_1683,N_24462,N_24838);
or UO_1684 (O_1684,N_24572,N_24563);
nor UO_1685 (O_1685,N_24477,N_24675);
nor UO_1686 (O_1686,N_24800,N_24577);
nor UO_1687 (O_1687,N_24986,N_24737);
and UO_1688 (O_1688,N_24858,N_24961);
nand UO_1689 (O_1689,N_24554,N_24404);
and UO_1690 (O_1690,N_24574,N_24414);
nor UO_1691 (O_1691,N_24751,N_24430);
nand UO_1692 (O_1692,N_24541,N_24933);
nor UO_1693 (O_1693,N_24470,N_24857);
nand UO_1694 (O_1694,N_24573,N_24706);
and UO_1695 (O_1695,N_24595,N_24866);
or UO_1696 (O_1696,N_24789,N_24438);
and UO_1697 (O_1697,N_24613,N_24859);
and UO_1698 (O_1698,N_24625,N_24462);
nor UO_1699 (O_1699,N_24581,N_24522);
and UO_1700 (O_1700,N_24764,N_24733);
nor UO_1701 (O_1701,N_24536,N_24470);
and UO_1702 (O_1702,N_24848,N_24765);
and UO_1703 (O_1703,N_24877,N_24836);
xor UO_1704 (O_1704,N_24793,N_24695);
nor UO_1705 (O_1705,N_24615,N_24766);
and UO_1706 (O_1706,N_24936,N_24514);
and UO_1707 (O_1707,N_24734,N_24473);
or UO_1708 (O_1708,N_24813,N_24726);
and UO_1709 (O_1709,N_24755,N_24399);
or UO_1710 (O_1710,N_24582,N_24848);
nor UO_1711 (O_1711,N_24528,N_24721);
xnor UO_1712 (O_1712,N_24618,N_24565);
and UO_1713 (O_1713,N_24507,N_24392);
or UO_1714 (O_1714,N_24434,N_24931);
or UO_1715 (O_1715,N_24882,N_24560);
and UO_1716 (O_1716,N_24946,N_24396);
nor UO_1717 (O_1717,N_24444,N_24622);
nand UO_1718 (O_1718,N_24745,N_24539);
nor UO_1719 (O_1719,N_24797,N_24505);
nor UO_1720 (O_1720,N_24535,N_24533);
nand UO_1721 (O_1721,N_24856,N_24608);
and UO_1722 (O_1722,N_24832,N_24603);
xnor UO_1723 (O_1723,N_24417,N_24690);
nor UO_1724 (O_1724,N_24889,N_24495);
nor UO_1725 (O_1725,N_24488,N_24647);
or UO_1726 (O_1726,N_24533,N_24393);
or UO_1727 (O_1727,N_24840,N_24559);
nand UO_1728 (O_1728,N_24831,N_24993);
nor UO_1729 (O_1729,N_24741,N_24600);
or UO_1730 (O_1730,N_24862,N_24943);
and UO_1731 (O_1731,N_24771,N_24621);
and UO_1732 (O_1732,N_24468,N_24375);
and UO_1733 (O_1733,N_24785,N_24755);
nor UO_1734 (O_1734,N_24868,N_24414);
nand UO_1735 (O_1735,N_24386,N_24595);
nand UO_1736 (O_1736,N_24604,N_24753);
nand UO_1737 (O_1737,N_24528,N_24401);
nor UO_1738 (O_1738,N_24393,N_24520);
nor UO_1739 (O_1739,N_24577,N_24998);
and UO_1740 (O_1740,N_24743,N_24545);
and UO_1741 (O_1741,N_24516,N_24897);
nor UO_1742 (O_1742,N_24540,N_24899);
or UO_1743 (O_1743,N_24958,N_24714);
and UO_1744 (O_1744,N_24403,N_24740);
and UO_1745 (O_1745,N_24533,N_24794);
or UO_1746 (O_1746,N_24980,N_24907);
xor UO_1747 (O_1747,N_24632,N_24935);
nor UO_1748 (O_1748,N_24978,N_24973);
and UO_1749 (O_1749,N_24875,N_24721);
and UO_1750 (O_1750,N_24379,N_24378);
nor UO_1751 (O_1751,N_24857,N_24981);
and UO_1752 (O_1752,N_24887,N_24930);
and UO_1753 (O_1753,N_24957,N_24729);
nor UO_1754 (O_1754,N_24428,N_24859);
or UO_1755 (O_1755,N_24480,N_24942);
nor UO_1756 (O_1756,N_24927,N_24620);
nand UO_1757 (O_1757,N_24516,N_24784);
or UO_1758 (O_1758,N_24507,N_24669);
nor UO_1759 (O_1759,N_24834,N_24699);
nor UO_1760 (O_1760,N_24922,N_24524);
nor UO_1761 (O_1761,N_24876,N_24855);
and UO_1762 (O_1762,N_24386,N_24841);
or UO_1763 (O_1763,N_24684,N_24978);
or UO_1764 (O_1764,N_24461,N_24946);
and UO_1765 (O_1765,N_24521,N_24530);
or UO_1766 (O_1766,N_24819,N_24901);
nand UO_1767 (O_1767,N_24495,N_24661);
nor UO_1768 (O_1768,N_24914,N_24838);
or UO_1769 (O_1769,N_24950,N_24405);
nand UO_1770 (O_1770,N_24722,N_24493);
nand UO_1771 (O_1771,N_24688,N_24964);
nor UO_1772 (O_1772,N_24726,N_24932);
nor UO_1773 (O_1773,N_24614,N_24853);
nor UO_1774 (O_1774,N_24480,N_24913);
nand UO_1775 (O_1775,N_24817,N_24418);
nand UO_1776 (O_1776,N_24899,N_24759);
and UO_1777 (O_1777,N_24505,N_24502);
nor UO_1778 (O_1778,N_24612,N_24726);
or UO_1779 (O_1779,N_24802,N_24558);
nand UO_1780 (O_1780,N_24764,N_24635);
nor UO_1781 (O_1781,N_24871,N_24812);
nor UO_1782 (O_1782,N_24434,N_24872);
and UO_1783 (O_1783,N_24907,N_24918);
xor UO_1784 (O_1784,N_24623,N_24843);
nand UO_1785 (O_1785,N_24391,N_24561);
and UO_1786 (O_1786,N_24421,N_24844);
xnor UO_1787 (O_1787,N_24730,N_24881);
xnor UO_1788 (O_1788,N_24943,N_24643);
nand UO_1789 (O_1789,N_24615,N_24624);
nand UO_1790 (O_1790,N_24589,N_24535);
and UO_1791 (O_1791,N_24909,N_24864);
or UO_1792 (O_1792,N_24412,N_24585);
and UO_1793 (O_1793,N_24985,N_24635);
nand UO_1794 (O_1794,N_24831,N_24391);
xor UO_1795 (O_1795,N_24720,N_24950);
or UO_1796 (O_1796,N_24518,N_24713);
xnor UO_1797 (O_1797,N_24766,N_24653);
xor UO_1798 (O_1798,N_24678,N_24687);
and UO_1799 (O_1799,N_24397,N_24968);
and UO_1800 (O_1800,N_24435,N_24888);
or UO_1801 (O_1801,N_24679,N_24480);
or UO_1802 (O_1802,N_24933,N_24453);
nand UO_1803 (O_1803,N_24786,N_24671);
nor UO_1804 (O_1804,N_24555,N_24687);
or UO_1805 (O_1805,N_24569,N_24472);
nand UO_1806 (O_1806,N_24955,N_24697);
xnor UO_1807 (O_1807,N_24679,N_24649);
or UO_1808 (O_1808,N_24816,N_24703);
or UO_1809 (O_1809,N_24648,N_24815);
or UO_1810 (O_1810,N_24995,N_24610);
and UO_1811 (O_1811,N_24977,N_24555);
nor UO_1812 (O_1812,N_24867,N_24880);
nand UO_1813 (O_1813,N_24814,N_24841);
nand UO_1814 (O_1814,N_24724,N_24801);
and UO_1815 (O_1815,N_24773,N_24590);
nor UO_1816 (O_1816,N_24790,N_24994);
nand UO_1817 (O_1817,N_24376,N_24701);
nor UO_1818 (O_1818,N_24835,N_24636);
and UO_1819 (O_1819,N_24929,N_24671);
nor UO_1820 (O_1820,N_24508,N_24937);
or UO_1821 (O_1821,N_24738,N_24474);
nand UO_1822 (O_1822,N_24530,N_24639);
xnor UO_1823 (O_1823,N_24812,N_24783);
nand UO_1824 (O_1824,N_24710,N_24983);
and UO_1825 (O_1825,N_24773,N_24823);
nor UO_1826 (O_1826,N_24580,N_24637);
nor UO_1827 (O_1827,N_24817,N_24492);
nand UO_1828 (O_1828,N_24536,N_24499);
and UO_1829 (O_1829,N_24667,N_24476);
and UO_1830 (O_1830,N_24905,N_24548);
xor UO_1831 (O_1831,N_24470,N_24418);
nand UO_1832 (O_1832,N_24427,N_24836);
nor UO_1833 (O_1833,N_24778,N_24463);
nor UO_1834 (O_1834,N_24815,N_24415);
xnor UO_1835 (O_1835,N_24708,N_24598);
and UO_1836 (O_1836,N_24781,N_24490);
nor UO_1837 (O_1837,N_24408,N_24802);
or UO_1838 (O_1838,N_24376,N_24975);
nor UO_1839 (O_1839,N_24597,N_24807);
nor UO_1840 (O_1840,N_24453,N_24747);
or UO_1841 (O_1841,N_24925,N_24442);
nor UO_1842 (O_1842,N_24536,N_24619);
xor UO_1843 (O_1843,N_24855,N_24848);
or UO_1844 (O_1844,N_24434,N_24525);
and UO_1845 (O_1845,N_24517,N_24501);
xor UO_1846 (O_1846,N_24837,N_24880);
or UO_1847 (O_1847,N_24522,N_24985);
and UO_1848 (O_1848,N_24532,N_24844);
or UO_1849 (O_1849,N_24759,N_24729);
and UO_1850 (O_1850,N_24652,N_24406);
nand UO_1851 (O_1851,N_24446,N_24504);
and UO_1852 (O_1852,N_24661,N_24805);
and UO_1853 (O_1853,N_24903,N_24522);
nand UO_1854 (O_1854,N_24435,N_24883);
nand UO_1855 (O_1855,N_24587,N_24635);
nand UO_1856 (O_1856,N_24552,N_24670);
or UO_1857 (O_1857,N_24820,N_24644);
nor UO_1858 (O_1858,N_24938,N_24696);
nor UO_1859 (O_1859,N_24473,N_24629);
or UO_1860 (O_1860,N_24510,N_24796);
xor UO_1861 (O_1861,N_24823,N_24994);
nand UO_1862 (O_1862,N_24846,N_24441);
nor UO_1863 (O_1863,N_24901,N_24787);
and UO_1864 (O_1864,N_24477,N_24738);
and UO_1865 (O_1865,N_24733,N_24559);
and UO_1866 (O_1866,N_24645,N_24882);
or UO_1867 (O_1867,N_24747,N_24558);
nor UO_1868 (O_1868,N_24473,N_24730);
nor UO_1869 (O_1869,N_24383,N_24842);
nand UO_1870 (O_1870,N_24486,N_24705);
or UO_1871 (O_1871,N_24604,N_24792);
nand UO_1872 (O_1872,N_24730,N_24410);
xor UO_1873 (O_1873,N_24990,N_24394);
nor UO_1874 (O_1874,N_24806,N_24440);
nor UO_1875 (O_1875,N_24404,N_24527);
and UO_1876 (O_1876,N_24930,N_24557);
nand UO_1877 (O_1877,N_24606,N_24444);
or UO_1878 (O_1878,N_24956,N_24784);
nand UO_1879 (O_1879,N_24772,N_24723);
or UO_1880 (O_1880,N_24860,N_24649);
or UO_1881 (O_1881,N_24794,N_24902);
nor UO_1882 (O_1882,N_24515,N_24903);
and UO_1883 (O_1883,N_24450,N_24629);
nand UO_1884 (O_1884,N_24403,N_24454);
nand UO_1885 (O_1885,N_24993,N_24964);
or UO_1886 (O_1886,N_24395,N_24763);
and UO_1887 (O_1887,N_24664,N_24726);
nor UO_1888 (O_1888,N_24380,N_24649);
and UO_1889 (O_1889,N_24669,N_24943);
nor UO_1890 (O_1890,N_24831,N_24544);
or UO_1891 (O_1891,N_24999,N_24617);
or UO_1892 (O_1892,N_24726,N_24860);
nand UO_1893 (O_1893,N_24623,N_24819);
or UO_1894 (O_1894,N_24610,N_24486);
and UO_1895 (O_1895,N_24763,N_24672);
nor UO_1896 (O_1896,N_24871,N_24735);
or UO_1897 (O_1897,N_24483,N_24649);
xor UO_1898 (O_1898,N_24589,N_24674);
nor UO_1899 (O_1899,N_24473,N_24926);
and UO_1900 (O_1900,N_24967,N_24958);
nand UO_1901 (O_1901,N_24966,N_24416);
or UO_1902 (O_1902,N_24722,N_24897);
nand UO_1903 (O_1903,N_24671,N_24775);
and UO_1904 (O_1904,N_24582,N_24821);
nand UO_1905 (O_1905,N_24681,N_24666);
nor UO_1906 (O_1906,N_24791,N_24598);
nor UO_1907 (O_1907,N_24795,N_24989);
nor UO_1908 (O_1908,N_24468,N_24662);
nand UO_1909 (O_1909,N_24750,N_24885);
nor UO_1910 (O_1910,N_24427,N_24553);
nand UO_1911 (O_1911,N_24376,N_24729);
nor UO_1912 (O_1912,N_24666,N_24988);
nand UO_1913 (O_1913,N_24525,N_24797);
and UO_1914 (O_1914,N_24825,N_24899);
or UO_1915 (O_1915,N_24381,N_24767);
nor UO_1916 (O_1916,N_24601,N_24733);
nor UO_1917 (O_1917,N_24762,N_24973);
nand UO_1918 (O_1918,N_24814,N_24451);
nand UO_1919 (O_1919,N_24446,N_24432);
nor UO_1920 (O_1920,N_24818,N_24391);
nand UO_1921 (O_1921,N_24450,N_24696);
nor UO_1922 (O_1922,N_24604,N_24714);
and UO_1923 (O_1923,N_24815,N_24929);
nand UO_1924 (O_1924,N_24996,N_24710);
and UO_1925 (O_1925,N_24948,N_24584);
and UO_1926 (O_1926,N_24494,N_24414);
nand UO_1927 (O_1927,N_24583,N_24730);
or UO_1928 (O_1928,N_24569,N_24801);
and UO_1929 (O_1929,N_24697,N_24871);
and UO_1930 (O_1930,N_24713,N_24743);
nor UO_1931 (O_1931,N_24859,N_24710);
and UO_1932 (O_1932,N_24646,N_24735);
and UO_1933 (O_1933,N_24976,N_24382);
nand UO_1934 (O_1934,N_24622,N_24789);
nand UO_1935 (O_1935,N_24611,N_24943);
nand UO_1936 (O_1936,N_24897,N_24443);
nor UO_1937 (O_1937,N_24931,N_24903);
nor UO_1938 (O_1938,N_24823,N_24677);
xor UO_1939 (O_1939,N_24861,N_24488);
or UO_1940 (O_1940,N_24952,N_24461);
or UO_1941 (O_1941,N_24766,N_24791);
nor UO_1942 (O_1942,N_24882,N_24379);
nand UO_1943 (O_1943,N_24622,N_24691);
and UO_1944 (O_1944,N_24489,N_24453);
nand UO_1945 (O_1945,N_24756,N_24969);
nor UO_1946 (O_1946,N_24930,N_24742);
or UO_1947 (O_1947,N_24404,N_24870);
nand UO_1948 (O_1948,N_24879,N_24666);
nor UO_1949 (O_1949,N_24412,N_24716);
xor UO_1950 (O_1950,N_24581,N_24755);
or UO_1951 (O_1951,N_24769,N_24514);
xnor UO_1952 (O_1952,N_24528,N_24729);
xor UO_1953 (O_1953,N_24490,N_24660);
nor UO_1954 (O_1954,N_24746,N_24613);
and UO_1955 (O_1955,N_24811,N_24551);
and UO_1956 (O_1956,N_24874,N_24927);
and UO_1957 (O_1957,N_24511,N_24574);
nand UO_1958 (O_1958,N_24809,N_24387);
or UO_1959 (O_1959,N_24554,N_24955);
or UO_1960 (O_1960,N_24502,N_24974);
xnor UO_1961 (O_1961,N_24691,N_24592);
or UO_1962 (O_1962,N_24869,N_24487);
or UO_1963 (O_1963,N_24701,N_24869);
nor UO_1964 (O_1964,N_24790,N_24472);
nor UO_1965 (O_1965,N_24472,N_24545);
or UO_1966 (O_1966,N_24740,N_24817);
nor UO_1967 (O_1967,N_24784,N_24521);
nand UO_1968 (O_1968,N_24640,N_24714);
xnor UO_1969 (O_1969,N_24536,N_24618);
and UO_1970 (O_1970,N_24828,N_24500);
nor UO_1971 (O_1971,N_24443,N_24396);
nor UO_1972 (O_1972,N_24383,N_24644);
nor UO_1973 (O_1973,N_24405,N_24477);
nand UO_1974 (O_1974,N_24400,N_24925);
nand UO_1975 (O_1975,N_24570,N_24553);
nand UO_1976 (O_1976,N_24618,N_24572);
or UO_1977 (O_1977,N_24823,N_24921);
nor UO_1978 (O_1978,N_24690,N_24885);
nand UO_1979 (O_1979,N_24987,N_24856);
nor UO_1980 (O_1980,N_24555,N_24618);
nor UO_1981 (O_1981,N_24752,N_24452);
nor UO_1982 (O_1982,N_24614,N_24916);
nand UO_1983 (O_1983,N_24787,N_24464);
nor UO_1984 (O_1984,N_24786,N_24563);
or UO_1985 (O_1985,N_24941,N_24425);
or UO_1986 (O_1986,N_24645,N_24424);
xnor UO_1987 (O_1987,N_24402,N_24745);
and UO_1988 (O_1988,N_24705,N_24460);
and UO_1989 (O_1989,N_24606,N_24879);
nand UO_1990 (O_1990,N_24622,N_24776);
nor UO_1991 (O_1991,N_24822,N_24611);
or UO_1992 (O_1992,N_24640,N_24516);
nand UO_1993 (O_1993,N_24740,N_24642);
and UO_1994 (O_1994,N_24916,N_24952);
or UO_1995 (O_1995,N_24854,N_24789);
or UO_1996 (O_1996,N_24813,N_24376);
xor UO_1997 (O_1997,N_24756,N_24652);
and UO_1998 (O_1998,N_24999,N_24502);
and UO_1999 (O_1999,N_24909,N_24956);
nand UO_2000 (O_2000,N_24819,N_24920);
nor UO_2001 (O_2001,N_24492,N_24785);
or UO_2002 (O_2002,N_24585,N_24672);
or UO_2003 (O_2003,N_24713,N_24721);
or UO_2004 (O_2004,N_24818,N_24664);
nor UO_2005 (O_2005,N_24789,N_24765);
nand UO_2006 (O_2006,N_24673,N_24793);
nand UO_2007 (O_2007,N_24860,N_24948);
nand UO_2008 (O_2008,N_24902,N_24542);
nand UO_2009 (O_2009,N_24802,N_24602);
nand UO_2010 (O_2010,N_24384,N_24995);
or UO_2011 (O_2011,N_24615,N_24781);
xnor UO_2012 (O_2012,N_24627,N_24526);
nor UO_2013 (O_2013,N_24425,N_24981);
nor UO_2014 (O_2014,N_24930,N_24520);
nor UO_2015 (O_2015,N_24964,N_24607);
xor UO_2016 (O_2016,N_24433,N_24496);
or UO_2017 (O_2017,N_24512,N_24644);
nor UO_2018 (O_2018,N_24570,N_24978);
and UO_2019 (O_2019,N_24682,N_24648);
and UO_2020 (O_2020,N_24978,N_24831);
nor UO_2021 (O_2021,N_24485,N_24753);
and UO_2022 (O_2022,N_24529,N_24659);
nor UO_2023 (O_2023,N_24637,N_24406);
xor UO_2024 (O_2024,N_24549,N_24749);
or UO_2025 (O_2025,N_24991,N_24927);
nor UO_2026 (O_2026,N_24408,N_24508);
and UO_2027 (O_2027,N_24636,N_24522);
xnor UO_2028 (O_2028,N_24477,N_24911);
nand UO_2029 (O_2029,N_24954,N_24806);
nor UO_2030 (O_2030,N_24642,N_24525);
and UO_2031 (O_2031,N_24465,N_24859);
and UO_2032 (O_2032,N_24423,N_24468);
and UO_2033 (O_2033,N_24911,N_24951);
or UO_2034 (O_2034,N_24587,N_24447);
nor UO_2035 (O_2035,N_24804,N_24935);
and UO_2036 (O_2036,N_24654,N_24434);
xor UO_2037 (O_2037,N_24666,N_24530);
nand UO_2038 (O_2038,N_24724,N_24704);
or UO_2039 (O_2039,N_24808,N_24722);
xnor UO_2040 (O_2040,N_24790,N_24629);
and UO_2041 (O_2041,N_24375,N_24697);
and UO_2042 (O_2042,N_24447,N_24457);
nor UO_2043 (O_2043,N_24642,N_24482);
nand UO_2044 (O_2044,N_24587,N_24948);
nor UO_2045 (O_2045,N_24803,N_24569);
or UO_2046 (O_2046,N_24562,N_24705);
nor UO_2047 (O_2047,N_24589,N_24438);
nand UO_2048 (O_2048,N_24461,N_24599);
nand UO_2049 (O_2049,N_24386,N_24624);
nor UO_2050 (O_2050,N_24993,N_24927);
nand UO_2051 (O_2051,N_24848,N_24927);
and UO_2052 (O_2052,N_24459,N_24988);
or UO_2053 (O_2053,N_24560,N_24444);
and UO_2054 (O_2054,N_24780,N_24835);
and UO_2055 (O_2055,N_24632,N_24959);
nor UO_2056 (O_2056,N_24895,N_24971);
and UO_2057 (O_2057,N_24872,N_24878);
and UO_2058 (O_2058,N_24881,N_24569);
or UO_2059 (O_2059,N_24761,N_24416);
nor UO_2060 (O_2060,N_24874,N_24742);
or UO_2061 (O_2061,N_24511,N_24672);
xnor UO_2062 (O_2062,N_24919,N_24538);
nand UO_2063 (O_2063,N_24720,N_24862);
nand UO_2064 (O_2064,N_24558,N_24968);
or UO_2065 (O_2065,N_24963,N_24427);
nor UO_2066 (O_2066,N_24589,N_24414);
nor UO_2067 (O_2067,N_24763,N_24750);
and UO_2068 (O_2068,N_24846,N_24944);
nand UO_2069 (O_2069,N_24890,N_24977);
and UO_2070 (O_2070,N_24382,N_24889);
and UO_2071 (O_2071,N_24852,N_24992);
nand UO_2072 (O_2072,N_24596,N_24979);
nor UO_2073 (O_2073,N_24849,N_24756);
nand UO_2074 (O_2074,N_24710,N_24664);
or UO_2075 (O_2075,N_24444,N_24781);
or UO_2076 (O_2076,N_24940,N_24883);
and UO_2077 (O_2077,N_24472,N_24859);
xnor UO_2078 (O_2078,N_24417,N_24454);
nand UO_2079 (O_2079,N_24541,N_24482);
and UO_2080 (O_2080,N_24508,N_24527);
or UO_2081 (O_2081,N_24392,N_24983);
and UO_2082 (O_2082,N_24437,N_24825);
or UO_2083 (O_2083,N_24825,N_24509);
nor UO_2084 (O_2084,N_24545,N_24913);
and UO_2085 (O_2085,N_24545,N_24725);
and UO_2086 (O_2086,N_24885,N_24749);
nand UO_2087 (O_2087,N_24603,N_24643);
or UO_2088 (O_2088,N_24815,N_24652);
nand UO_2089 (O_2089,N_24612,N_24407);
and UO_2090 (O_2090,N_24936,N_24955);
nand UO_2091 (O_2091,N_24824,N_24682);
or UO_2092 (O_2092,N_24752,N_24916);
nand UO_2093 (O_2093,N_24505,N_24795);
nor UO_2094 (O_2094,N_24505,N_24552);
nand UO_2095 (O_2095,N_24725,N_24945);
and UO_2096 (O_2096,N_24733,N_24751);
nor UO_2097 (O_2097,N_24924,N_24896);
nand UO_2098 (O_2098,N_24913,N_24946);
nand UO_2099 (O_2099,N_24911,N_24781);
or UO_2100 (O_2100,N_24529,N_24530);
nor UO_2101 (O_2101,N_24820,N_24547);
nor UO_2102 (O_2102,N_24990,N_24880);
or UO_2103 (O_2103,N_24950,N_24989);
nor UO_2104 (O_2104,N_24513,N_24519);
and UO_2105 (O_2105,N_24996,N_24496);
or UO_2106 (O_2106,N_24888,N_24615);
and UO_2107 (O_2107,N_24563,N_24932);
nor UO_2108 (O_2108,N_24549,N_24975);
or UO_2109 (O_2109,N_24735,N_24751);
or UO_2110 (O_2110,N_24686,N_24866);
or UO_2111 (O_2111,N_24957,N_24632);
or UO_2112 (O_2112,N_24976,N_24544);
xor UO_2113 (O_2113,N_24587,N_24606);
and UO_2114 (O_2114,N_24631,N_24449);
nor UO_2115 (O_2115,N_24922,N_24540);
xnor UO_2116 (O_2116,N_24452,N_24668);
nand UO_2117 (O_2117,N_24749,N_24725);
or UO_2118 (O_2118,N_24436,N_24768);
nand UO_2119 (O_2119,N_24860,N_24445);
xnor UO_2120 (O_2120,N_24777,N_24779);
nor UO_2121 (O_2121,N_24523,N_24644);
and UO_2122 (O_2122,N_24632,N_24571);
or UO_2123 (O_2123,N_24586,N_24392);
and UO_2124 (O_2124,N_24989,N_24771);
or UO_2125 (O_2125,N_24418,N_24452);
or UO_2126 (O_2126,N_24838,N_24912);
or UO_2127 (O_2127,N_24441,N_24847);
and UO_2128 (O_2128,N_24880,N_24402);
and UO_2129 (O_2129,N_24451,N_24450);
or UO_2130 (O_2130,N_24851,N_24387);
or UO_2131 (O_2131,N_24422,N_24401);
and UO_2132 (O_2132,N_24546,N_24537);
nand UO_2133 (O_2133,N_24865,N_24614);
nor UO_2134 (O_2134,N_24672,N_24395);
and UO_2135 (O_2135,N_24872,N_24586);
nand UO_2136 (O_2136,N_24987,N_24430);
nand UO_2137 (O_2137,N_24910,N_24937);
nor UO_2138 (O_2138,N_24837,N_24611);
and UO_2139 (O_2139,N_24445,N_24982);
and UO_2140 (O_2140,N_24706,N_24912);
nand UO_2141 (O_2141,N_24619,N_24455);
nor UO_2142 (O_2142,N_24769,N_24737);
nand UO_2143 (O_2143,N_24936,N_24725);
and UO_2144 (O_2144,N_24994,N_24484);
xnor UO_2145 (O_2145,N_24475,N_24956);
and UO_2146 (O_2146,N_24964,N_24406);
nor UO_2147 (O_2147,N_24748,N_24536);
or UO_2148 (O_2148,N_24951,N_24747);
nor UO_2149 (O_2149,N_24986,N_24395);
or UO_2150 (O_2150,N_24387,N_24865);
and UO_2151 (O_2151,N_24584,N_24976);
and UO_2152 (O_2152,N_24722,N_24771);
and UO_2153 (O_2153,N_24876,N_24417);
and UO_2154 (O_2154,N_24733,N_24807);
or UO_2155 (O_2155,N_24573,N_24625);
or UO_2156 (O_2156,N_24767,N_24567);
or UO_2157 (O_2157,N_24609,N_24725);
or UO_2158 (O_2158,N_24590,N_24465);
and UO_2159 (O_2159,N_24529,N_24502);
nor UO_2160 (O_2160,N_24426,N_24444);
or UO_2161 (O_2161,N_24840,N_24777);
nand UO_2162 (O_2162,N_24798,N_24479);
nand UO_2163 (O_2163,N_24862,N_24936);
nor UO_2164 (O_2164,N_24924,N_24709);
and UO_2165 (O_2165,N_24621,N_24704);
or UO_2166 (O_2166,N_24848,N_24579);
nand UO_2167 (O_2167,N_24690,N_24558);
or UO_2168 (O_2168,N_24660,N_24948);
nor UO_2169 (O_2169,N_24870,N_24815);
and UO_2170 (O_2170,N_24700,N_24712);
and UO_2171 (O_2171,N_24974,N_24688);
or UO_2172 (O_2172,N_24994,N_24890);
and UO_2173 (O_2173,N_24909,N_24644);
or UO_2174 (O_2174,N_24417,N_24552);
or UO_2175 (O_2175,N_24901,N_24595);
and UO_2176 (O_2176,N_24717,N_24468);
nand UO_2177 (O_2177,N_24854,N_24503);
or UO_2178 (O_2178,N_24753,N_24484);
or UO_2179 (O_2179,N_24398,N_24947);
or UO_2180 (O_2180,N_24916,N_24665);
or UO_2181 (O_2181,N_24788,N_24517);
and UO_2182 (O_2182,N_24380,N_24395);
nand UO_2183 (O_2183,N_24628,N_24920);
nand UO_2184 (O_2184,N_24449,N_24396);
and UO_2185 (O_2185,N_24876,N_24393);
and UO_2186 (O_2186,N_24698,N_24426);
or UO_2187 (O_2187,N_24769,N_24607);
nor UO_2188 (O_2188,N_24963,N_24701);
and UO_2189 (O_2189,N_24737,N_24544);
xnor UO_2190 (O_2190,N_24442,N_24444);
or UO_2191 (O_2191,N_24622,N_24800);
nand UO_2192 (O_2192,N_24798,N_24752);
and UO_2193 (O_2193,N_24397,N_24700);
or UO_2194 (O_2194,N_24424,N_24826);
and UO_2195 (O_2195,N_24659,N_24464);
and UO_2196 (O_2196,N_24901,N_24784);
nand UO_2197 (O_2197,N_24998,N_24484);
nand UO_2198 (O_2198,N_24384,N_24884);
nand UO_2199 (O_2199,N_24953,N_24925);
or UO_2200 (O_2200,N_24618,N_24996);
nand UO_2201 (O_2201,N_24468,N_24969);
nand UO_2202 (O_2202,N_24888,N_24853);
xor UO_2203 (O_2203,N_24729,N_24480);
nor UO_2204 (O_2204,N_24545,N_24583);
or UO_2205 (O_2205,N_24696,N_24816);
nand UO_2206 (O_2206,N_24565,N_24630);
or UO_2207 (O_2207,N_24971,N_24732);
or UO_2208 (O_2208,N_24618,N_24601);
nand UO_2209 (O_2209,N_24892,N_24633);
and UO_2210 (O_2210,N_24486,N_24649);
nor UO_2211 (O_2211,N_24445,N_24651);
and UO_2212 (O_2212,N_24749,N_24763);
xor UO_2213 (O_2213,N_24528,N_24825);
and UO_2214 (O_2214,N_24761,N_24614);
and UO_2215 (O_2215,N_24865,N_24927);
nor UO_2216 (O_2216,N_24965,N_24466);
nor UO_2217 (O_2217,N_24820,N_24746);
or UO_2218 (O_2218,N_24557,N_24376);
nand UO_2219 (O_2219,N_24526,N_24736);
and UO_2220 (O_2220,N_24478,N_24980);
and UO_2221 (O_2221,N_24815,N_24664);
nand UO_2222 (O_2222,N_24814,N_24538);
nor UO_2223 (O_2223,N_24461,N_24963);
or UO_2224 (O_2224,N_24904,N_24950);
nor UO_2225 (O_2225,N_24890,N_24561);
or UO_2226 (O_2226,N_24975,N_24768);
nor UO_2227 (O_2227,N_24626,N_24704);
and UO_2228 (O_2228,N_24643,N_24632);
xnor UO_2229 (O_2229,N_24615,N_24863);
and UO_2230 (O_2230,N_24594,N_24931);
or UO_2231 (O_2231,N_24498,N_24987);
nor UO_2232 (O_2232,N_24973,N_24941);
nor UO_2233 (O_2233,N_24599,N_24514);
xor UO_2234 (O_2234,N_24982,N_24459);
nor UO_2235 (O_2235,N_24869,N_24504);
nand UO_2236 (O_2236,N_24963,N_24678);
nand UO_2237 (O_2237,N_24616,N_24427);
and UO_2238 (O_2238,N_24619,N_24633);
xnor UO_2239 (O_2239,N_24751,N_24704);
or UO_2240 (O_2240,N_24945,N_24809);
or UO_2241 (O_2241,N_24933,N_24662);
nor UO_2242 (O_2242,N_24996,N_24667);
or UO_2243 (O_2243,N_24381,N_24721);
and UO_2244 (O_2244,N_24975,N_24943);
xnor UO_2245 (O_2245,N_24915,N_24978);
or UO_2246 (O_2246,N_24790,N_24808);
nand UO_2247 (O_2247,N_24441,N_24519);
or UO_2248 (O_2248,N_24471,N_24385);
and UO_2249 (O_2249,N_24665,N_24937);
or UO_2250 (O_2250,N_24914,N_24876);
and UO_2251 (O_2251,N_24401,N_24786);
xor UO_2252 (O_2252,N_24926,N_24758);
or UO_2253 (O_2253,N_24498,N_24670);
nand UO_2254 (O_2254,N_24793,N_24490);
and UO_2255 (O_2255,N_24519,N_24920);
nand UO_2256 (O_2256,N_24570,N_24757);
or UO_2257 (O_2257,N_24473,N_24435);
nand UO_2258 (O_2258,N_24579,N_24495);
nand UO_2259 (O_2259,N_24509,N_24791);
or UO_2260 (O_2260,N_24797,N_24467);
xnor UO_2261 (O_2261,N_24621,N_24799);
and UO_2262 (O_2262,N_24461,N_24693);
and UO_2263 (O_2263,N_24868,N_24634);
or UO_2264 (O_2264,N_24706,N_24748);
and UO_2265 (O_2265,N_24835,N_24576);
nor UO_2266 (O_2266,N_24620,N_24914);
nor UO_2267 (O_2267,N_24973,N_24902);
and UO_2268 (O_2268,N_24948,N_24960);
and UO_2269 (O_2269,N_24515,N_24693);
and UO_2270 (O_2270,N_24688,N_24934);
xor UO_2271 (O_2271,N_24995,N_24780);
nand UO_2272 (O_2272,N_24428,N_24679);
xor UO_2273 (O_2273,N_24396,N_24639);
nor UO_2274 (O_2274,N_24717,N_24614);
and UO_2275 (O_2275,N_24857,N_24465);
and UO_2276 (O_2276,N_24745,N_24698);
and UO_2277 (O_2277,N_24480,N_24428);
xnor UO_2278 (O_2278,N_24827,N_24993);
nand UO_2279 (O_2279,N_24523,N_24598);
and UO_2280 (O_2280,N_24975,N_24572);
nand UO_2281 (O_2281,N_24448,N_24927);
nor UO_2282 (O_2282,N_24423,N_24854);
and UO_2283 (O_2283,N_24894,N_24481);
nand UO_2284 (O_2284,N_24713,N_24483);
nand UO_2285 (O_2285,N_24395,N_24976);
nand UO_2286 (O_2286,N_24823,N_24628);
nor UO_2287 (O_2287,N_24444,N_24580);
nand UO_2288 (O_2288,N_24453,N_24651);
nor UO_2289 (O_2289,N_24871,N_24471);
nand UO_2290 (O_2290,N_24577,N_24561);
and UO_2291 (O_2291,N_24443,N_24769);
nand UO_2292 (O_2292,N_24483,N_24798);
nand UO_2293 (O_2293,N_24895,N_24743);
or UO_2294 (O_2294,N_24888,N_24961);
and UO_2295 (O_2295,N_24505,N_24570);
nand UO_2296 (O_2296,N_24848,N_24602);
and UO_2297 (O_2297,N_24931,N_24456);
nand UO_2298 (O_2298,N_24862,N_24985);
and UO_2299 (O_2299,N_24915,N_24972);
and UO_2300 (O_2300,N_24590,N_24375);
or UO_2301 (O_2301,N_24961,N_24467);
or UO_2302 (O_2302,N_24869,N_24653);
or UO_2303 (O_2303,N_24638,N_24993);
and UO_2304 (O_2304,N_24734,N_24688);
or UO_2305 (O_2305,N_24890,N_24831);
xor UO_2306 (O_2306,N_24624,N_24455);
nor UO_2307 (O_2307,N_24693,N_24521);
nor UO_2308 (O_2308,N_24760,N_24566);
and UO_2309 (O_2309,N_24896,N_24473);
nor UO_2310 (O_2310,N_24712,N_24788);
nor UO_2311 (O_2311,N_24596,N_24570);
nand UO_2312 (O_2312,N_24562,N_24734);
and UO_2313 (O_2313,N_24915,N_24544);
nor UO_2314 (O_2314,N_24866,N_24580);
or UO_2315 (O_2315,N_24801,N_24697);
or UO_2316 (O_2316,N_24930,N_24440);
nand UO_2317 (O_2317,N_24556,N_24703);
and UO_2318 (O_2318,N_24417,N_24864);
nand UO_2319 (O_2319,N_24839,N_24942);
nand UO_2320 (O_2320,N_24418,N_24692);
nor UO_2321 (O_2321,N_24379,N_24598);
nand UO_2322 (O_2322,N_24402,N_24775);
nand UO_2323 (O_2323,N_24840,N_24846);
and UO_2324 (O_2324,N_24678,N_24794);
xnor UO_2325 (O_2325,N_24418,N_24917);
nor UO_2326 (O_2326,N_24511,N_24425);
nand UO_2327 (O_2327,N_24763,N_24848);
nand UO_2328 (O_2328,N_24503,N_24975);
or UO_2329 (O_2329,N_24378,N_24577);
and UO_2330 (O_2330,N_24720,N_24875);
nand UO_2331 (O_2331,N_24558,N_24543);
or UO_2332 (O_2332,N_24724,N_24454);
nor UO_2333 (O_2333,N_24534,N_24841);
and UO_2334 (O_2334,N_24541,N_24849);
and UO_2335 (O_2335,N_24854,N_24485);
and UO_2336 (O_2336,N_24721,N_24417);
nor UO_2337 (O_2337,N_24617,N_24539);
nor UO_2338 (O_2338,N_24682,N_24820);
and UO_2339 (O_2339,N_24940,N_24736);
nand UO_2340 (O_2340,N_24684,N_24822);
xor UO_2341 (O_2341,N_24827,N_24932);
nor UO_2342 (O_2342,N_24930,N_24487);
or UO_2343 (O_2343,N_24517,N_24841);
xnor UO_2344 (O_2344,N_24748,N_24503);
and UO_2345 (O_2345,N_24849,N_24895);
or UO_2346 (O_2346,N_24926,N_24652);
nand UO_2347 (O_2347,N_24544,N_24575);
nand UO_2348 (O_2348,N_24434,N_24802);
and UO_2349 (O_2349,N_24830,N_24520);
nor UO_2350 (O_2350,N_24614,N_24386);
nand UO_2351 (O_2351,N_24811,N_24406);
nor UO_2352 (O_2352,N_24549,N_24973);
and UO_2353 (O_2353,N_24448,N_24557);
and UO_2354 (O_2354,N_24634,N_24787);
and UO_2355 (O_2355,N_24814,N_24443);
and UO_2356 (O_2356,N_24559,N_24712);
or UO_2357 (O_2357,N_24758,N_24762);
xnor UO_2358 (O_2358,N_24497,N_24951);
nor UO_2359 (O_2359,N_24584,N_24482);
or UO_2360 (O_2360,N_24787,N_24826);
or UO_2361 (O_2361,N_24765,N_24602);
or UO_2362 (O_2362,N_24459,N_24526);
nand UO_2363 (O_2363,N_24985,N_24832);
nor UO_2364 (O_2364,N_24555,N_24397);
xor UO_2365 (O_2365,N_24955,N_24389);
and UO_2366 (O_2366,N_24934,N_24871);
or UO_2367 (O_2367,N_24899,N_24895);
or UO_2368 (O_2368,N_24850,N_24723);
and UO_2369 (O_2369,N_24792,N_24892);
or UO_2370 (O_2370,N_24531,N_24417);
nand UO_2371 (O_2371,N_24883,N_24815);
or UO_2372 (O_2372,N_24875,N_24979);
nor UO_2373 (O_2373,N_24550,N_24790);
nand UO_2374 (O_2374,N_24709,N_24624);
xor UO_2375 (O_2375,N_24919,N_24781);
nor UO_2376 (O_2376,N_24924,N_24406);
or UO_2377 (O_2377,N_24375,N_24939);
nor UO_2378 (O_2378,N_24918,N_24882);
or UO_2379 (O_2379,N_24382,N_24826);
nand UO_2380 (O_2380,N_24660,N_24812);
nand UO_2381 (O_2381,N_24902,N_24554);
or UO_2382 (O_2382,N_24915,N_24578);
nand UO_2383 (O_2383,N_24816,N_24836);
and UO_2384 (O_2384,N_24684,N_24500);
or UO_2385 (O_2385,N_24985,N_24730);
and UO_2386 (O_2386,N_24836,N_24528);
and UO_2387 (O_2387,N_24887,N_24965);
nand UO_2388 (O_2388,N_24580,N_24407);
nand UO_2389 (O_2389,N_24709,N_24398);
and UO_2390 (O_2390,N_24759,N_24557);
nor UO_2391 (O_2391,N_24843,N_24625);
and UO_2392 (O_2392,N_24951,N_24485);
nand UO_2393 (O_2393,N_24890,N_24743);
xnor UO_2394 (O_2394,N_24499,N_24687);
or UO_2395 (O_2395,N_24744,N_24669);
nor UO_2396 (O_2396,N_24839,N_24849);
or UO_2397 (O_2397,N_24394,N_24384);
or UO_2398 (O_2398,N_24993,N_24985);
or UO_2399 (O_2399,N_24463,N_24928);
nand UO_2400 (O_2400,N_24486,N_24835);
and UO_2401 (O_2401,N_24878,N_24539);
or UO_2402 (O_2402,N_24542,N_24564);
nor UO_2403 (O_2403,N_24558,N_24593);
xor UO_2404 (O_2404,N_24967,N_24917);
or UO_2405 (O_2405,N_24749,N_24705);
and UO_2406 (O_2406,N_24508,N_24812);
and UO_2407 (O_2407,N_24389,N_24520);
nand UO_2408 (O_2408,N_24715,N_24546);
nor UO_2409 (O_2409,N_24866,N_24949);
or UO_2410 (O_2410,N_24437,N_24751);
and UO_2411 (O_2411,N_24830,N_24726);
nand UO_2412 (O_2412,N_24463,N_24960);
nand UO_2413 (O_2413,N_24906,N_24473);
nand UO_2414 (O_2414,N_24949,N_24811);
and UO_2415 (O_2415,N_24944,N_24683);
nand UO_2416 (O_2416,N_24580,N_24442);
nand UO_2417 (O_2417,N_24814,N_24563);
nand UO_2418 (O_2418,N_24443,N_24494);
or UO_2419 (O_2419,N_24735,N_24461);
xnor UO_2420 (O_2420,N_24522,N_24827);
nor UO_2421 (O_2421,N_24459,N_24894);
nand UO_2422 (O_2422,N_24786,N_24763);
xnor UO_2423 (O_2423,N_24632,N_24778);
and UO_2424 (O_2424,N_24541,N_24380);
or UO_2425 (O_2425,N_24773,N_24859);
nor UO_2426 (O_2426,N_24720,N_24745);
nor UO_2427 (O_2427,N_24864,N_24916);
or UO_2428 (O_2428,N_24650,N_24624);
and UO_2429 (O_2429,N_24738,N_24405);
and UO_2430 (O_2430,N_24838,N_24749);
and UO_2431 (O_2431,N_24468,N_24840);
or UO_2432 (O_2432,N_24479,N_24820);
or UO_2433 (O_2433,N_24468,N_24573);
nor UO_2434 (O_2434,N_24434,N_24564);
nor UO_2435 (O_2435,N_24896,N_24778);
nor UO_2436 (O_2436,N_24604,N_24476);
nand UO_2437 (O_2437,N_24856,N_24844);
nand UO_2438 (O_2438,N_24828,N_24377);
and UO_2439 (O_2439,N_24686,N_24858);
and UO_2440 (O_2440,N_24944,N_24587);
nand UO_2441 (O_2441,N_24794,N_24718);
nand UO_2442 (O_2442,N_24591,N_24947);
nor UO_2443 (O_2443,N_24701,N_24572);
xor UO_2444 (O_2444,N_24906,N_24881);
or UO_2445 (O_2445,N_24848,N_24608);
or UO_2446 (O_2446,N_24741,N_24934);
and UO_2447 (O_2447,N_24793,N_24888);
and UO_2448 (O_2448,N_24638,N_24639);
or UO_2449 (O_2449,N_24607,N_24928);
or UO_2450 (O_2450,N_24391,N_24419);
nor UO_2451 (O_2451,N_24521,N_24808);
nor UO_2452 (O_2452,N_24469,N_24470);
or UO_2453 (O_2453,N_24997,N_24735);
and UO_2454 (O_2454,N_24748,N_24631);
xnor UO_2455 (O_2455,N_24907,N_24624);
or UO_2456 (O_2456,N_24462,N_24835);
nor UO_2457 (O_2457,N_24682,N_24724);
xor UO_2458 (O_2458,N_24938,N_24921);
nand UO_2459 (O_2459,N_24608,N_24849);
nand UO_2460 (O_2460,N_24451,N_24963);
nor UO_2461 (O_2461,N_24491,N_24898);
nand UO_2462 (O_2462,N_24489,N_24398);
and UO_2463 (O_2463,N_24608,N_24689);
or UO_2464 (O_2464,N_24966,N_24508);
nor UO_2465 (O_2465,N_24592,N_24448);
and UO_2466 (O_2466,N_24431,N_24924);
and UO_2467 (O_2467,N_24634,N_24955);
and UO_2468 (O_2468,N_24829,N_24484);
or UO_2469 (O_2469,N_24687,N_24683);
nand UO_2470 (O_2470,N_24396,N_24768);
nand UO_2471 (O_2471,N_24991,N_24431);
nand UO_2472 (O_2472,N_24975,N_24389);
nand UO_2473 (O_2473,N_24990,N_24602);
and UO_2474 (O_2474,N_24885,N_24575);
nor UO_2475 (O_2475,N_24816,N_24678);
nor UO_2476 (O_2476,N_24621,N_24470);
nor UO_2477 (O_2477,N_24817,N_24952);
nor UO_2478 (O_2478,N_24712,N_24588);
and UO_2479 (O_2479,N_24380,N_24735);
nor UO_2480 (O_2480,N_24445,N_24387);
and UO_2481 (O_2481,N_24419,N_24871);
or UO_2482 (O_2482,N_24990,N_24996);
nand UO_2483 (O_2483,N_24805,N_24719);
or UO_2484 (O_2484,N_24417,N_24604);
xnor UO_2485 (O_2485,N_24469,N_24781);
and UO_2486 (O_2486,N_24788,N_24555);
and UO_2487 (O_2487,N_24908,N_24572);
nor UO_2488 (O_2488,N_24646,N_24641);
nand UO_2489 (O_2489,N_24710,N_24947);
or UO_2490 (O_2490,N_24843,N_24798);
xnor UO_2491 (O_2491,N_24942,N_24471);
nor UO_2492 (O_2492,N_24952,N_24733);
nor UO_2493 (O_2493,N_24438,N_24586);
nor UO_2494 (O_2494,N_24883,N_24487);
nor UO_2495 (O_2495,N_24920,N_24655);
or UO_2496 (O_2496,N_24799,N_24510);
nand UO_2497 (O_2497,N_24644,N_24832);
and UO_2498 (O_2498,N_24801,N_24926);
or UO_2499 (O_2499,N_24939,N_24861);
or UO_2500 (O_2500,N_24625,N_24733);
and UO_2501 (O_2501,N_24608,N_24547);
or UO_2502 (O_2502,N_24936,N_24934);
xor UO_2503 (O_2503,N_24403,N_24869);
xnor UO_2504 (O_2504,N_24767,N_24851);
or UO_2505 (O_2505,N_24587,N_24778);
and UO_2506 (O_2506,N_24710,N_24621);
and UO_2507 (O_2507,N_24455,N_24486);
and UO_2508 (O_2508,N_24513,N_24765);
nand UO_2509 (O_2509,N_24599,N_24414);
or UO_2510 (O_2510,N_24531,N_24877);
or UO_2511 (O_2511,N_24853,N_24531);
nand UO_2512 (O_2512,N_24584,N_24758);
nand UO_2513 (O_2513,N_24987,N_24977);
and UO_2514 (O_2514,N_24823,N_24930);
nor UO_2515 (O_2515,N_24608,N_24378);
nor UO_2516 (O_2516,N_24895,N_24699);
nand UO_2517 (O_2517,N_24756,N_24390);
and UO_2518 (O_2518,N_24980,N_24828);
and UO_2519 (O_2519,N_24630,N_24881);
nor UO_2520 (O_2520,N_24906,N_24652);
or UO_2521 (O_2521,N_24928,N_24494);
and UO_2522 (O_2522,N_24521,N_24502);
or UO_2523 (O_2523,N_24822,N_24732);
nor UO_2524 (O_2524,N_24938,N_24996);
nor UO_2525 (O_2525,N_24519,N_24922);
and UO_2526 (O_2526,N_24723,N_24524);
nand UO_2527 (O_2527,N_24700,N_24834);
nor UO_2528 (O_2528,N_24913,N_24404);
xor UO_2529 (O_2529,N_24563,N_24697);
nor UO_2530 (O_2530,N_24958,N_24840);
nor UO_2531 (O_2531,N_24594,N_24778);
nand UO_2532 (O_2532,N_24689,N_24505);
or UO_2533 (O_2533,N_24718,N_24938);
nor UO_2534 (O_2534,N_24576,N_24915);
nor UO_2535 (O_2535,N_24704,N_24475);
or UO_2536 (O_2536,N_24590,N_24893);
nand UO_2537 (O_2537,N_24690,N_24811);
nor UO_2538 (O_2538,N_24607,N_24540);
or UO_2539 (O_2539,N_24664,N_24501);
xor UO_2540 (O_2540,N_24700,N_24533);
nand UO_2541 (O_2541,N_24787,N_24616);
nor UO_2542 (O_2542,N_24650,N_24945);
xor UO_2543 (O_2543,N_24726,N_24575);
xnor UO_2544 (O_2544,N_24981,N_24673);
or UO_2545 (O_2545,N_24751,N_24457);
or UO_2546 (O_2546,N_24543,N_24505);
nand UO_2547 (O_2547,N_24637,N_24831);
nor UO_2548 (O_2548,N_24543,N_24682);
xor UO_2549 (O_2549,N_24387,N_24926);
nor UO_2550 (O_2550,N_24435,N_24829);
and UO_2551 (O_2551,N_24946,N_24529);
and UO_2552 (O_2552,N_24918,N_24834);
and UO_2553 (O_2553,N_24620,N_24811);
or UO_2554 (O_2554,N_24471,N_24532);
nor UO_2555 (O_2555,N_24625,N_24897);
xor UO_2556 (O_2556,N_24506,N_24526);
nand UO_2557 (O_2557,N_24639,N_24744);
xnor UO_2558 (O_2558,N_24894,N_24844);
xnor UO_2559 (O_2559,N_24824,N_24969);
xnor UO_2560 (O_2560,N_24583,N_24870);
or UO_2561 (O_2561,N_24572,N_24858);
nor UO_2562 (O_2562,N_24991,N_24525);
nand UO_2563 (O_2563,N_24648,N_24969);
nand UO_2564 (O_2564,N_24528,N_24972);
or UO_2565 (O_2565,N_24992,N_24451);
and UO_2566 (O_2566,N_24499,N_24901);
or UO_2567 (O_2567,N_24882,N_24644);
nor UO_2568 (O_2568,N_24998,N_24437);
and UO_2569 (O_2569,N_24572,N_24413);
nor UO_2570 (O_2570,N_24537,N_24566);
and UO_2571 (O_2571,N_24463,N_24492);
or UO_2572 (O_2572,N_24988,N_24903);
nand UO_2573 (O_2573,N_24553,N_24749);
nand UO_2574 (O_2574,N_24552,N_24467);
and UO_2575 (O_2575,N_24677,N_24753);
nand UO_2576 (O_2576,N_24626,N_24932);
nor UO_2577 (O_2577,N_24467,N_24747);
or UO_2578 (O_2578,N_24642,N_24699);
nand UO_2579 (O_2579,N_24897,N_24573);
nand UO_2580 (O_2580,N_24787,N_24795);
nand UO_2581 (O_2581,N_24810,N_24787);
nand UO_2582 (O_2582,N_24548,N_24657);
nand UO_2583 (O_2583,N_24497,N_24923);
and UO_2584 (O_2584,N_24406,N_24390);
or UO_2585 (O_2585,N_24990,N_24453);
or UO_2586 (O_2586,N_24788,N_24537);
or UO_2587 (O_2587,N_24444,N_24540);
nor UO_2588 (O_2588,N_24589,N_24918);
and UO_2589 (O_2589,N_24536,N_24953);
nor UO_2590 (O_2590,N_24453,N_24600);
or UO_2591 (O_2591,N_24708,N_24773);
nand UO_2592 (O_2592,N_24885,N_24516);
xnor UO_2593 (O_2593,N_24765,N_24383);
nand UO_2594 (O_2594,N_24888,N_24648);
xor UO_2595 (O_2595,N_24500,N_24834);
nor UO_2596 (O_2596,N_24526,N_24612);
nor UO_2597 (O_2597,N_24613,N_24763);
nor UO_2598 (O_2598,N_24626,N_24710);
or UO_2599 (O_2599,N_24967,N_24538);
xor UO_2600 (O_2600,N_24790,N_24910);
nand UO_2601 (O_2601,N_24849,N_24877);
xor UO_2602 (O_2602,N_24914,N_24492);
nor UO_2603 (O_2603,N_24723,N_24858);
nor UO_2604 (O_2604,N_24505,N_24474);
nand UO_2605 (O_2605,N_24942,N_24487);
and UO_2606 (O_2606,N_24530,N_24600);
nor UO_2607 (O_2607,N_24616,N_24806);
and UO_2608 (O_2608,N_24678,N_24631);
nand UO_2609 (O_2609,N_24408,N_24759);
nor UO_2610 (O_2610,N_24833,N_24634);
nand UO_2611 (O_2611,N_24517,N_24450);
or UO_2612 (O_2612,N_24720,N_24376);
xnor UO_2613 (O_2613,N_24433,N_24747);
or UO_2614 (O_2614,N_24418,N_24398);
nor UO_2615 (O_2615,N_24550,N_24660);
nor UO_2616 (O_2616,N_24784,N_24559);
nor UO_2617 (O_2617,N_24987,N_24652);
nor UO_2618 (O_2618,N_24623,N_24913);
xor UO_2619 (O_2619,N_24860,N_24388);
nand UO_2620 (O_2620,N_24915,N_24976);
and UO_2621 (O_2621,N_24678,N_24386);
or UO_2622 (O_2622,N_24680,N_24939);
nand UO_2623 (O_2623,N_24981,N_24830);
or UO_2624 (O_2624,N_24580,N_24915);
and UO_2625 (O_2625,N_24692,N_24683);
and UO_2626 (O_2626,N_24600,N_24375);
or UO_2627 (O_2627,N_24494,N_24873);
xor UO_2628 (O_2628,N_24533,N_24415);
and UO_2629 (O_2629,N_24735,N_24575);
or UO_2630 (O_2630,N_24495,N_24778);
nand UO_2631 (O_2631,N_24488,N_24567);
and UO_2632 (O_2632,N_24966,N_24567);
and UO_2633 (O_2633,N_24654,N_24809);
nand UO_2634 (O_2634,N_24762,N_24781);
xor UO_2635 (O_2635,N_24642,N_24947);
xnor UO_2636 (O_2636,N_24569,N_24827);
or UO_2637 (O_2637,N_24841,N_24458);
nor UO_2638 (O_2638,N_24847,N_24879);
or UO_2639 (O_2639,N_24695,N_24869);
nor UO_2640 (O_2640,N_24462,N_24419);
nand UO_2641 (O_2641,N_24555,N_24928);
and UO_2642 (O_2642,N_24805,N_24798);
nor UO_2643 (O_2643,N_24624,N_24573);
and UO_2644 (O_2644,N_24399,N_24417);
and UO_2645 (O_2645,N_24782,N_24624);
and UO_2646 (O_2646,N_24943,N_24737);
and UO_2647 (O_2647,N_24379,N_24535);
nor UO_2648 (O_2648,N_24976,N_24646);
or UO_2649 (O_2649,N_24975,N_24966);
nor UO_2650 (O_2650,N_24614,N_24499);
and UO_2651 (O_2651,N_24523,N_24496);
nand UO_2652 (O_2652,N_24667,N_24817);
nand UO_2653 (O_2653,N_24610,N_24463);
nor UO_2654 (O_2654,N_24982,N_24609);
nand UO_2655 (O_2655,N_24402,N_24981);
nor UO_2656 (O_2656,N_24383,N_24411);
xor UO_2657 (O_2657,N_24759,N_24655);
or UO_2658 (O_2658,N_24902,N_24664);
nand UO_2659 (O_2659,N_24889,N_24934);
or UO_2660 (O_2660,N_24884,N_24523);
nand UO_2661 (O_2661,N_24419,N_24620);
and UO_2662 (O_2662,N_24946,N_24874);
nand UO_2663 (O_2663,N_24686,N_24914);
or UO_2664 (O_2664,N_24658,N_24755);
and UO_2665 (O_2665,N_24949,N_24477);
and UO_2666 (O_2666,N_24566,N_24888);
and UO_2667 (O_2667,N_24683,N_24455);
xor UO_2668 (O_2668,N_24824,N_24749);
nand UO_2669 (O_2669,N_24608,N_24866);
and UO_2670 (O_2670,N_24603,N_24751);
nand UO_2671 (O_2671,N_24457,N_24928);
nor UO_2672 (O_2672,N_24479,N_24511);
nor UO_2673 (O_2673,N_24896,N_24551);
or UO_2674 (O_2674,N_24530,N_24786);
and UO_2675 (O_2675,N_24446,N_24417);
xor UO_2676 (O_2676,N_24608,N_24936);
or UO_2677 (O_2677,N_24916,N_24666);
nor UO_2678 (O_2678,N_24620,N_24609);
nand UO_2679 (O_2679,N_24957,N_24719);
nor UO_2680 (O_2680,N_24702,N_24640);
and UO_2681 (O_2681,N_24928,N_24398);
and UO_2682 (O_2682,N_24913,N_24445);
nor UO_2683 (O_2683,N_24506,N_24870);
and UO_2684 (O_2684,N_24755,N_24874);
or UO_2685 (O_2685,N_24581,N_24520);
and UO_2686 (O_2686,N_24420,N_24791);
or UO_2687 (O_2687,N_24556,N_24674);
and UO_2688 (O_2688,N_24784,N_24489);
nor UO_2689 (O_2689,N_24565,N_24701);
nor UO_2690 (O_2690,N_24375,N_24489);
nand UO_2691 (O_2691,N_24695,N_24510);
nor UO_2692 (O_2692,N_24947,N_24986);
nand UO_2693 (O_2693,N_24463,N_24894);
and UO_2694 (O_2694,N_24771,N_24611);
or UO_2695 (O_2695,N_24939,N_24795);
nor UO_2696 (O_2696,N_24680,N_24776);
or UO_2697 (O_2697,N_24740,N_24910);
nor UO_2698 (O_2698,N_24765,N_24974);
xnor UO_2699 (O_2699,N_24906,N_24797);
nor UO_2700 (O_2700,N_24541,N_24875);
nand UO_2701 (O_2701,N_24484,N_24904);
nor UO_2702 (O_2702,N_24674,N_24916);
or UO_2703 (O_2703,N_24983,N_24857);
nor UO_2704 (O_2704,N_24956,N_24671);
nor UO_2705 (O_2705,N_24585,N_24721);
nor UO_2706 (O_2706,N_24937,N_24482);
and UO_2707 (O_2707,N_24430,N_24654);
and UO_2708 (O_2708,N_24583,N_24546);
nand UO_2709 (O_2709,N_24868,N_24785);
nor UO_2710 (O_2710,N_24772,N_24444);
nor UO_2711 (O_2711,N_24759,N_24592);
nand UO_2712 (O_2712,N_24523,N_24793);
xor UO_2713 (O_2713,N_24923,N_24808);
or UO_2714 (O_2714,N_24949,N_24834);
xnor UO_2715 (O_2715,N_24927,N_24870);
or UO_2716 (O_2716,N_24805,N_24706);
and UO_2717 (O_2717,N_24441,N_24724);
and UO_2718 (O_2718,N_24923,N_24517);
nand UO_2719 (O_2719,N_24625,N_24507);
or UO_2720 (O_2720,N_24666,N_24670);
and UO_2721 (O_2721,N_24519,N_24432);
or UO_2722 (O_2722,N_24983,N_24875);
nand UO_2723 (O_2723,N_24394,N_24403);
nor UO_2724 (O_2724,N_24386,N_24998);
and UO_2725 (O_2725,N_24840,N_24568);
or UO_2726 (O_2726,N_24732,N_24591);
or UO_2727 (O_2727,N_24718,N_24666);
and UO_2728 (O_2728,N_24543,N_24965);
xor UO_2729 (O_2729,N_24641,N_24425);
and UO_2730 (O_2730,N_24382,N_24606);
nor UO_2731 (O_2731,N_24588,N_24510);
nor UO_2732 (O_2732,N_24652,N_24589);
and UO_2733 (O_2733,N_24787,N_24497);
nor UO_2734 (O_2734,N_24924,N_24691);
nand UO_2735 (O_2735,N_24386,N_24399);
or UO_2736 (O_2736,N_24421,N_24768);
nor UO_2737 (O_2737,N_24633,N_24911);
nand UO_2738 (O_2738,N_24694,N_24667);
nor UO_2739 (O_2739,N_24631,N_24540);
and UO_2740 (O_2740,N_24767,N_24545);
and UO_2741 (O_2741,N_24757,N_24461);
xor UO_2742 (O_2742,N_24564,N_24465);
nor UO_2743 (O_2743,N_24421,N_24823);
nor UO_2744 (O_2744,N_24839,N_24578);
nor UO_2745 (O_2745,N_24381,N_24422);
and UO_2746 (O_2746,N_24612,N_24715);
nand UO_2747 (O_2747,N_24713,N_24827);
nand UO_2748 (O_2748,N_24998,N_24749);
and UO_2749 (O_2749,N_24702,N_24617);
and UO_2750 (O_2750,N_24899,N_24714);
nand UO_2751 (O_2751,N_24852,N_24702);
nor UO_2752 (O_2752,N_24532,N_24950);
nand UO_2753 (O_2753,N_24904,N_24497);
nor UO_2754 (O_2754,N_24432,N_24805);
and UO_2755 (O_2755,N_24863,N_24555);
and UO_2756 (O_2756,N_24443,N_24661);
nand UO_2757 (O_2757,N_24539,N_24529);
nand UO_2758 (O_2758,N_24974,N_24548);
or UO_2759 (O_2759,N_24726,N_24930);
or UO_2760 (O_2760,N_24623,N_24531);
nor UO_2761 (O_2761,N_24521,N_24546);
or UO_2762 (O_2762,N_24840,N_24621);
nor UO_2763 (O_2763,N_24798,N_24935);
or UO_2764 (O_2764,N_24844,N_24980);
nor UO_2765 (O_2765,N_24415,N_24483);
nand UO_2766 (O_2766,N_24995,N_24860);
and UO_2767 (O_2767,N_24379,N_24607);
nor UO_2768 (O_2768,N_24665,N_24733);
or UO_2769 (O_2769,N_24980,N_24638);
or UO_2770 (O_2770,N_24586,N_24951);
nand UO_2771 (O_2771,N_24418,N_24766);
nand UO_2772 (O_2772,N_24701,N_24856);
xor UO_2773 (O_2773,N_24784,N_24461);
or UO_2774 (O_2774,N_24764,N_24766);
xnor UO_2775 (O_2775,N_24844,N_24415);
nand UO_2776 (O_2776,N_24447,N_24389);
nor UO_2777 (O_2777,N_24383,N_24863);
or UO_2778 (O_2778,N_24454,N_24828);
or UO_2779 (O_2779,N_24900,N_24598);
or UO_2780 (O_2780,N_24839,N_24698);
and UO_2781 (O_2781,N_24804,N_24689);
nand UO_2782 (O_2782,N_24459,N_24873);
nor UO_2783 (O_2783,N_24546,N_24837);
xnor UO_2784 (O_2784,N_24902,N_24893);
nand UO_2785 (O_2785,N_24710,N_24546);
nor UO_2786 (O_2786,N_24976,N_24478);
nand UO_2787 (O_2787,N_24662,N_24830);
and UO_2788 (O_2788,N_24820,N_24534);
nor UO_2789 (O_2789,N_24516,N_24835);
nand UO_2790 (O_2790,N_24478,N_24512);
nor UO_2791 (O_2791,N_24597,N_24427);
and UO_2792 (O_2792,N_24729,N_24650);
and UO_2793 (O_2793,N_24634,N_24673);
xnor UO_2794 (O_2794,N_24513,N_24627);
nand UO_2795 (O_2795,N_24564,N_24476);
nand UO_2796 (O_2796,N_24725,N_24887);
nand UO_2797 (O_2797,N_24972,N_24810);
nand UO_2798 (O_2798,N_24951,N_24613);
nand UO_2799 (O_2799,N_24817,N_24475);
nand UO_2800 (O_2800,N_24721,N_24903);
nand UO_2801 (O_2801,N_24414,N_24927);
or UO_2802 (O_2802,N_24538,N_24418);
nor UO_2803 (O_2803,N_24421,N_24738);
nand UO_2804 (O_2804,N_24406,N_24454);
nor UO_2805 (O_2805,N_24957,N_24992);
nor UO_2806 (O_2806,N_24384,N_24599);
or UO_2807 (O_2807,N_24464,N_24419);
and UO_2808 (O_2808,N_24813,N_24460);
xor UO_2809 (O_2809,N_24528,N_24862);
nand UO_2810 (O_2810,N_24464,N_24417);
nand UO_2811 (O_2811,N_24619,N_24605);
nor UO_2812 (O_2812,N_24820,N_24618);
nand UO_2813 (O_2813,N_24562,N_24988);
nand UO_2814 (O_2814,N_24977,N_24617);
nor UO_2815 (O_2815,N_24710,N_24796);
and UO_2816 (O_2816,N_24553,N_24412);
and UO_2817 (O_2817,N_24994,N_24935);
and UO_2818 (O_2818,N_24682,N_24507);
or UO_2819 (O_2819,N_24750,N_24457);
nor UO_2820 (O_2820,N_24676,N_24437);
nor UO_2821 (O_2821,N_24764,N_24478);
nor UO_2822 (O_2822,N_24660,N_24379);
xor UO_2823 (O_2823,N_24418,N_24609);
and UO_2824 (O_2824,N_24787,N_24557);
nand UO_2825 (O_2825,N_24535,N_24671);
nand UO_2826 (O_2826,N_24436,N_24834);
and UO_2827 (O_2827,N_24969,N_24526);
and UO_2828 (O_2828,N_24445,N_24838);
nor UO_2829 (O_2829,N_24556,N_24480);
and UO_2830 (O_2830,N_24485,N_24703);
or UO_2831 (O_2831,N_24583,N_24912);
and UO_2832 (O_2832,N_24982,N_24977);
xnor UO_2833 (O_2833,N_24574,N_24611);
nand UO_2834 (O_2834,N_24533,N_24904);
and UO_2835 (O_2835,N_24855,N_24470);
nand UO_2836 (O_2836,N_24776,N_24446);
or UO_2837 (O_2837,N_24444,N_24476);
nor UO_2838 (O_2838,N_24564,N_24941);
nand UO_2839 (O_2839,N_24538,N_24843);
xor UO_2840 (O_2840,N_24397,N_24945);
or UO_2841 (O_2841,N_24760,N_24492);
nand UO_2842 (O_2842,N_24959,N_24669);
or UO_2843 (O_2843,N_24457,N_24856);
or UO_2844 (O_2844,N_24857,N_24907);
nand UO_2845 (O_2845,N_24733,N_24945);
or UO_2846 (O_2846,N_24942,N_24474);
nor UO_2847 (O_2847,N_24813,N_24890);
nand UO_2848 (O_2848,N_24875,N_24463);
and UO_2849 (O_2849,N_24718,N_24612);
or UO_2850 (O_2850,N_24978,N_24781);
and UO_2851 (O_2851,N_24406,N_24914);
nand UO_2852 (O_2852,N_24809,N_24877);
nand UO_2853 (O_2853,N_24760,N_24622);
nand UO_2854 (O_2854,N_24447,N_24796);
or UO_2855 (O_2855,N_24421,N_24664);
or UO_2856 (O_2856,N_24817,N_24942);
or UO_2857 (O_2857,N_24854,N_24773);
and UO_2858 (O_2858,N_24867,N_24966);
and UO_2859 (O_2859,N_24779,N_24459);
or UO_2860 (O_2860,N_24874,N_24436);
nor UO_2861 (O_2861,N_24475,N_24553);
and UO_2862 (O_2862,N_24790,N_24991);
xnor UO_2863 (O_2863,N_24442,N_24880);
or UO_2864 (O_2864,N_24798,N_24641);
nand UO_2865 (O_2865,N_24651,N_24874);
nor UO_2866 (O_2866,N_24466,N_24750);
nor UO_2867 (O_2867,N_24400,N_24510);
nor UO_2868 (O_2868,N_24948,N_24710);
nor UO_2869 (O_2869,N_24430,N_24826);
nor UO_2870 (O_2870,N_24546,N_24561);
nand UO_2871 (O_2871,N_24688,N_24529);
nand UO_2872 (O_2872,N_24760,N_24409);
or UO_2873 (O_2873,N_24737,N_24412);
and UO_2874 (O_2874,N_24793,N_24384);
nor UO_2875 (O_2875,N_24804,N_24982);
or UO_2876 (O_2876,N_24915,N_24827);
and UO_2877 (O_2877,N_24533,N_24697);
and UO_2878 (O_2878,N_24566,N_24555);
or UO_2879 (O_2879,N_24952,N_24500);
and UO_2880 (O_2880,N_24516,N_24954);
or UO_2881 (O_2881,N_24868,N_24458);
nor UO_2882 (O_2882,N_24634,N_24770);
and UO_2883 (O_2883,N_24705,N_24502);
nand UO_2884 (O_2884,N_24780,N_24572);
or UO_2885 (O_2885,N_24451,N_24924);
and UO_2886 (O_2886,N_24943,N_24718);
and UO_2887 (O_2887,N_24554,N_24414);
nor UO_2888 (O_2888,N_24558,N_24748);
and UO_2889 (O_2889,N_24655,N_24934);
and UO_2890 (O_2890,N_24445,N_24715);
and UO_2891 (O_2891,N_24609,N_24621);
and UO_2892 (O_2892,N_24610,N_24545);
xor UO_2893 (O_2893,N_24598,N_24508);
or UO_2894 (O_2894,N_24791,N_24843);
or UO_2895 (O_2895,N_24559,N_24405);
xnor UO_2896 (O_2896,N_24598,N_24832);
or UO_2897 (O_2897,N_24794,N_24793);
or UO_2898 (O_2898,N_24754,N_24775);
xnor UO_2899 (O_2899,N_24997,N_24897);
nor UO_2900 (O_2900,N_24394,N_24775);
nand UO_2901 (O_2901,N_24579,N_24619);
nor UO_2902 (O_2902,N_24469,N_24479);
nand UO_2903 (O_2903,N_24490,N_24497);
or UO_2904 (O_2904,N_24691,N_24419);
nand UO_2905 (O_2905,N_24631,N_24941);
nor UO_2906 (O_2906,N_24987,N_24871);
nor UO_2907 (O_2907,N_24879,N_24751);
or UO_2908 (O_2908,N_24488,N_24707);
nand UO_2909 (O_2909,N_24869,N_24417);
or UO_2910 (O_2910,N_24935,N_24731);
nor UO_2911 (O_2911,N_24999,N_24484);
nor UO_2912 (O_2912,N_24694,N_24850);
or UO_2913 (O_2913,N_24484,N_24905);
nand UO_2914 (O_2914,N_24509,N_24892);
nand UO_2915 (O_2915,N_24599,N_24506);
nor UO_2916 (O_2916,N_24846,N_24509);
nor UO_2917 (O_2917,N_24481,N_24687);
nand UO_2918 (O_2918,N_24580,N_24451);
nand UO_2919 (O_2919,N_24575,N_24631);
and UO_2920 (O_2920,N_24452,N_24644);
xor UO_2921 (O_2921,N_24495,N_24413);
and UO_2922 (O_2922,N_24560,N_24482);
and UO_2923 (O_2923,N_24771,N_24913);
nor UO_2924 (O_2924,N_24791,N_24953);
and UO_2925 (O_2925,N_24721,N_24602);
or UO_2926 (O_2926,N_24875,N_24988);
and UO_2927 (O_2927,N_24537,N_24586);
xnor UO_2928 (O_2928,N_24657,N_24823);
and UO_2929 (O_2929,N_24381,N_24441);
nor UO_2930 (O_2930,N_24409,N_24844);
xor UO_2931 (O_2931,N_24437,N_24477);
nand UO_2932 (O_2932,N_24967,N_24989);
nor UO_2933 (O_2933,N_24570,N_24628);
nor UO_2934 (O_2934,N_24803,N_24876);
and UO_2935 (O_2935,N_24888,N_24665);
xor UO_2936 (O_2936,N_24887,N_24453);
or UO_2937 (O_2937,N_24537,N_24535);
or UO_2938 (O_2938,N_24397,N_24898);
nor UO_2939 (O_2939,N_24761,N_24375);
and UO_2940 (O_2940,N_24898,N_24512);
and UO_2941 (O_2941,N_24535,N_24479);
or UO_2942 (O_2942,N_24871,N_24979);
and UO_2943 (O_2943,N_24872,N_24930);
nor UO_2944 (O_2944,N_24558,N_24715);
or UO_2945 (O_2945,N_24629,N_24380);
nor UO_2946 (O_2946,N_24546,N_24698);
nand UO_2947 (O_2947,N_24637,N_24694);
nand UO_2948 (O_2948,N_24409,N_24725);
and UO_2949 (O_2949,N_24787,N_24690);
or UO_2950 (O_2950,N_24562,N_24776);
nor UO_2951 (O_2951,N_24626,N_24884);
nor UO_2952 (O_2952,N_24444,N_24741);
or UO_2953 (O_2953,N_24766,N_24717);
or UO_2954 (O_2954,N_24450,N_24726);
nor UO_2955 (O_2955,N_24885,N_24727);
nand UO_2956 (O_2956,N_24934,N_24388);
xnor UO_2957 (O_2957,N_24675,N_24643);
or UO_2958 (O_2958,N_24929,N_24618);
and UO_2959 (O_2959,N_24969,N_24385);
or UO_2960 (O_2960,N_24960,N_24664);
nand UO_2961 (O_2961,N_24580,N_24475);
nor UO_2962 (O_2962,N_24691,N_24460);
nand UO_2963 (O_2963,N_24958,N_24448);
or UO_2964 (O_2964,N_24741,N_24661);
and UO_2965 (O_2965,N_24629,N_24832);
nand UO_2966 (O_2966,N_24702,N_24883);
nor UO_2967 (O_2967,N_24584,N_24483);
xor UO_2968 (O_2968,N_24688,N_24437);
or UO_2969 (O_2969,N_24971,N_24463);
and UO_2970 (O_2970,N_24535,N_24559);
nor UO_2971 (O_2971,N_24452,N_24945);
xor UO_2972 (O_2972,N_24917,N_24437);
nor UO_2973 (O_2973,N_24839,N_24732);
xnor UO_2974 (O_2974,N_24846,N_24566);
nand UO_2975 (O_2975,N_24715,N_24801);
or UO_2976 (O_2976,N_24760,N_24533);
nand UO_2977 (O_2977,N_24686,N_24380);
and UO_2978 (O_2978,N_24912,N_24402);
xnor UO_2979 (O_2979,N_24921,N_24514);
or UO_2980 (O_2980,N_24689,N_24500);
nand UO_2981 (O_2981,N_24502,N_24440);
and UO_2982 (O_2982,N_24979,N_24429);
or UO_2983 (O_2983,N_24468,N_24543);
or UO_2984 (O_2984,N_24794,N_24654);
or UO_2985 (O_2985,N_24810,N_24596);
or UO_2986 (O_2986,N_24606,N_24699);
nor UO_2987 (O_2987,N_24388,N_24380);
nand UO_2988 (O_2988,N_24819,N_24659);
xnor UO_2989 (O_2989,N_24650,N_24657);
or UO_2990 (O_2990,N_24391,N_24690);
and UO_2991 (O_2991,N_24687,N_24409);
or UO_2992 (O_2992,N_24669,N_24768);
or UO_2993 (O_2993,N_24821,N_24783);
or UO_2994 (O_2994,N_24572,N_24777);
and UO_2995 (O_2995,N_24783,N_24979);
nand UO_2996 (O_2996,N_24573,N_24825);
nand UO_2997 (O_2997,N_24693,N_24529);
nor UO_2998 (O_2998,N_24947,N_24980);
nor UO_2999 (O_2999,N_24449,N_24819);
endmodule