module basic_750_5000_1000_10_levels_2xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_535,In_390);
or U1 (N_1,In_698,In_514);
and U2 (N_2,In_428,In_440);
or U3 (N_3,In_749,In_153);
nand U4 (N_4,In_742,In_500);
nor U5 (N_5,In_11,In_323);
or U6 (N_6,In_561,In_690);
nand U7 (N_7,In_348,In_733);
xnor U8 (N_8,In_493,In_705);
or U9 (N_9,In_687,In_701);
nand U10 (N_10,In_100,In_329);
or U11 (N_11,In_360,In_22);
and U12 (N_12,In_251,In_73);
xnor U13 (N_13,In_16,In_572);
and U14 (N_14,In_651,In_363);
and U15 (N_15,In_290,In_60);
and U16 (N_16,In_693,In_124);
nand U17 (N_17,In_478,In_497);
nand U18 (N_18,In_120,In_51);
nand U19 (N_19,In_242,In_315);
nor U20 (N_20,In_117,In_410);
and U21 (N_21,In_660,In_585);
or U22 (N_22,In_353,In_339);
nor U23 (N_23,In_154,In_181);
nand U24 (N_24,In_89,In_375);
nor U25 (N_25,In_383,In_683);
and U26 (N_26,In_14,In_308);
and U27 (N_27,In_175,In_487);
nand U28 (N_28,In_80,In_593);
nor U29 (N_29,In_692,In_189);
and U30 (N_30,In_295,In_451);
nand U31 (N_31,In_657,In_634);
nand U32 (N_32,In_261,In_185);
nand U33 (N_33,In_1,In_522);
nand U34 (N_34,In_187,In_145);
and U35 (N_35,In_574,In_267);
nand U36 (N_36,In_531,In_157);
nor U37 (N_37,In_695,In_337);
and U38 (N_38,In_538,In_639);
and U39 (N_39,In_352,In_626);
nand U40 (N_40,In_438,In_503);
nor U41 (N_41,In_196,In_677);
and U42 (N_42,In_617,In_653);
nand U43 (N_43,In_411,In_463);
nor U44 (N_44,In_130,In_443);
or U45 (N_45,In_466,In_311);
nor U46 (N_46,In_654,In_663);
and U47 (N_47,In_128,In_256);
nor U48 (N_48,In_179,In_480);
nor U49 (N_49,In_725,In_288);
nand U50 (N_50,In_621,In_243);
or U51 (N_51,In_36,In_3);
nor U52 (N_52,In_482,In_301);
or U53 (N_53,In_43,In_155);
and U54 (N_54,In_598,In_414);
nor U55 (N_55,In_183,In_165);
nand U56 (N_56,In_380,In_214);
or U57 (N_57,In_647,In_268);
and U58 (N_58,In_282,In_401);
and U59 (N_59,In_442,In_605);
nor U60 (N_60,In_52,In_686);
or U61 (N_61,In_333,In_250);
nand U62 (N_62,In_211,In_118);
and U63 (N_63,In_545,In_426);
nor U64 (N_64,In_32,In_404);
and U65 (N_65,In_659,In_412);
nor U66 (N_66,In_330,In_37);
nor U67 (N_67,In_48,In_46);
or U68 (N_68,In_257,In_361);
nand U69 (N_69,In_416,In_544);
or U70 (N_70,In_523,In_540);
and U71 (N_71,In_205,In_381);
nand U72 (N_72,In_174,In_345);
nor U73 (N_73,In_619,In_533);
nand U74 (N_74,In_467,In_58);
and U75 (N_75,In_423,In_57);
nor U76 (N_76,In_370,In_335);
nand U77 (N_77,In_312,In_527);
or U78 (N_78,In_332,In_20);
nor U79 (N_79,In_114,In_304);
and U80 (N_80,In_539,In_13);
nand U81 (N_81,In_0,In_296);
and U82 (N_82,In_642,In_292);
and U83 (N_83,In_618,In_373);
or U84 (N_84,In_392,In_699);
and U85 (N_85,In_650,In_581);
nand U86 (N_86,In_286,In_240);
nand U87 (N_87,In_158,In_355);
and U88 (N_88,In_177,In_310);
nor U89 (N_89,In_230,In_673);
and U90 (N_90,In_204,In_351);
and U91 (N_91,In_190,In_324);
or U92 (N_92,In_244,In_568);
nand U93 (N_93,In_403,In_417);
nor U94 (N_94,In_629,In_364);
or U95 (N_95,In_488,In_726);
or U96 (N_96,In_8,In_309);
nor U97 (N_97,In_41,In_342);
or U98 (N_98,In_649,In_162);
and U99 (N_99,In_79,In_265);
nor U100 (N_100,In_389,In_449);
or U101 (N_101,In_139,In_570);
nor U102 (N_102,In_253,In_528);
and U103 (N_103,In_624,In_447);
and U104 (N_104,In_529,In_547);
nand U105 (N_105,In_602,In_94);
and U106 (N_106,In_241,In_317);
nand U107 (N_107,In_446,In_633);
or U108 (N_108,In_26,In_648);
nand U109 (N_109,In_402,In_325);
and U110 (N_110,In_313,In_49);
and U111 (N_111,In_521,In_15);
nor U112 (N_112,In_548,In_149);
xor U113 (N_113,In_623,In_543);
nand U114 (N_114,In_279,In_209);
xnor U115 (N_115,In_280,In_7);
nand U116 (N_116,In_559,In_391);
nand U117 (N_117,In_587,In_688);
nor U118 (N_118,In_70,In_56);
nand U119 (N_119,In_628,In_249);
nor U120 (N_120,In_69,In_591);
and U121 (N_121,In_576,In_397);
nor U122 (N_122,In_512,In_638);
nand U123 (N_123,In_456,In_563);
nand U124 (N_124,In_81,In_431);
nand U125 (N_125,In_458,In_129);
nand U126 (N_126,In_374,In_588);
and U127 (N_127,In_247,In_93);
nor U128 (N_128,In_142,In_746);
and U129 (N_129,In_72,In_65);
and U130 (N_130,In_468,In_106);
xor U131 (N_131,In_112,In_387);
or U132 (N_132,In_107,In_67);
nand U133 (N_133,In_105,In_55);
nand U134 (N_134,In_481,In_422);
and U135 (N_135,In_223,In_10);
or U136 (N_136,In_729,In_151);
nor U137 (N_137,In_327,In_741);
or U138 (N_138,In_747,In_109);
nor U139 (N_139,In_691,In_731);
and U140 (N_140,In_645,In_314);
nand U141 (N_141,In_224,In_719);
and U142 (N_142,In_409,In_732);
nor U143 (N_143,In_516,In_226);
and U144 (N_144,In_276,In_511);
and U145 (N_145,In_385,In_513);
and U146 (N_146,In_668,In_465);
and U147 (N_147,In_349,In_703);
or U148 (N_148,In_245,In_667);
nand U149 (N_149,In_297,In_672);
nor U150 (N_150,In_195,In_554);
and U151 (N_151,In_640,In_86);
nand U152 (N_152,In_376,In_104);
and U153 (N_153,In_289,In_121);
nand U154 (N_154,In_437,In_435);
or U155 (N_155,In_358,In_33);
nand U156 (N_156,In_494,In_225);
or U157 (N_157,In_708,In_291);
and U158 (N_158,In_182,In_168);
and U159 (N_159,In_62,In_546);
nor U160 (N_160,In_486,In_103);
nor U161 (N_161,In_408,In_90);
or U162 (N_162,In_459,In_346);
nand U163 (N_163,In_713,In_116);
nor U164 (N_164,In_405,In_125);
or U165 (N_165,In_508,In_50);
nand U166 (N_166,In_433,In_192);
or U167 (N_167,In_160,In_365);
and U168 (N_168,In_441,In_206);
and U169 (N_169,In_338,In_322);
xnor U170 (N_170,In_550,In_284);
nand U171 (N_171,In_236,In_212);
nor U172 (N_172,In_340,In_658);
or U173 (N_173,In_501,In_630);
nor U174 (N_174,In_450,In_717);
nand U175 (N_175,In_586,In_287);
nor U176 (N_176,In_606,In_252);
or U177 (N_177,In_607,In_172);
or U178 (N_178,In_328,In_6);
or U179 (N_179,In_115,In_439);
or U180 (N_180,In_716,In_263);
or U181 (N_181,In_88,In_98);
or U182 (N_182,In_24,In_156);
nand U183 (N_183,In_394,In_643);
nor U184 (N_184,In_294,In_565);
and U185 (N_185,In_743,In_674);
nand U186 (N_186,In_278,In_470);
nand U187 (N_187,In_184,In_59);
nand U188 (N_188,In_293,In_302);
and U189 (N_189,In_61,In_525);
or U190 (N_190,In_455,In_191);
or U191 (N_191,In_661,In_347);
and U192 (N_192,In_343,In_331);
xor U193 (N_193,In_709,In_534);
nand U194 (N_194,In_722,In_97);
nor U195 (N_195,In_715,In_359);
and U196 (N_196,In_551,In_697);
nor U197 (N_197,In_113,In_696);
nor U198 (N_198,In_300,In_202);
nand U199 (N_199,In_530,In_307);
or U200 (N_200,In_232,In_738);
xnor U201 (N_201,In_398,In_178);
and U202 (N_202,In_453,In_47);
or U203 (N_203,In_150,In_135);
nor U204 (N_204,In_163,In_372);
nor U205 (N_205,In_499,In_532);
nor U206 (N_206,In_234,In_622);
nand U207 (N_207,In_694,In_171);
and U208 (N_208,In_173,In_371);
nor U209 (N_209,In_415,In_474);
or U210 (N_210,In_608,In_542);
nor U211 (N_211,In_12,In_111);
nor U212 (N_212,In_445,In_737);
xnor U213 (N_213,In_655,In_711);
nor U214 (N_214,In_569,In_469);
nor U215 (N_215,In_199,In_53);
nor U216 (N_216,In_38,In_498);
or U217 (N_217,In_666,In_727);
nand U218 (N_218,In_258,In_320);
nand U219 (N_219,In_613,In_203);
and U220 (N_220,In_396,In_644);
nor U221 (N_221,In_386,In_40);
or U222 (N_222,In_44,In_420);
nand U223 (N_223,In_4,In_636);
or U224 (N_224,In_573,In_367);
and U225 (N_225,In_369,In_176);
nand U226 (N_226,In_427,In_123);
nand U227 (N_227,In_495,In_518);
or U228 (N_228,In_736,In_600);
nand U229 (N_229,In_334,In_259);
nand U230 (N_230,In_595,In_509);
and U231 (N_231,In_75,In_616);
and U232 (N_232,In_641,In_96);
and U233 (N_233,In_266,In_164);
or U234 (N_234,In_601,In_552);
or U235 (N_235,In_589,In_670);
or U236 (N_236,In_744,In_366);
nand U237 (N_237,In_676,In_134);
and U238 (N_238,In_68,In_611);
nand U239 (N_239,In_418,In_235);
nand U240 (N_240,In_193,In_39);
xor U241 (N_241,In_248,In_144);
xor U242 (N_242,In_87,In_632);
and U243 (N_243,In_198,In_133);
nor U244 (N_244,In_555,In_524);
nand U245 (N_245,In_305,In_146);
nor U246 (N_246,In_707,In_567);
or U247 (N_247,In_461,In_669);
nor U248 (N_248,In_505,In_34);
nand U249 (N_249,In_406,In_471);
nand U250 (N_250,In_664,In_710);
nand U251 (N_251,In_84,In_132);
nor U252 (N_252,In_491,In_614);
and U253 (N_253,In_444,In_99);
or U254 (N_254,In_473,In_679);
or U255 (N_255,In_739,In_485);
or U256 (N_256,In_228,In_42);
or U257 (N_257,In_354,In_101);
and U258 (N_258,In_64,In_421);
nor U259 (N_259,In_510,In_652);
nand U260 (N_260,In_239,In_635);
nor U261 (N_261,In_395,In_77);
or U262 (N_262,In_273,In_603);
nand U263 (N_263,In_76,In_148);
xor U264 (N_264,In_682,In_400);
nor U265 (N_265,In_194,In_745);
xor U266 (N_266,In_303,In_233);
nor U267 (N_267,In_92,In_489);
nor U268 (N_268,In_558,In_384);
and U269 (N_269,In_169,In_63);
nor U270 (N_270,In_718,In_271);
xnor U271 (N_271,In_662,In_319);
and U272 (N_272,In_637,In_583);
nor U273 (N_273,In_45,In_393);
xnor U274 (N_274,In_377,In_143);
or U275 (N_275,In_584,In_141);
and U276 (N_276,In_326,In_460);
or U277 (N_277,In_425,In_216);
nand U278 (N_278,In_186,In_432);
or U279 (N_279,In_298,In_188);
and U280 (N_280,In_5,In_272);
and U281 (N_281,In_388,In_28);
and U282 (N_282,In_122,In_483);
nand U283 (N_283,In_571,In_200);
or U284 (N_284,In_656,In_452);
and U285 (N_285,In_379,In_27);
nand U286 (N_286,In_597,In_54);
or U287 (N_287,In_556,In_25);
and U288 (N_288,In_476,In_430);
or U289 (N_289,In_706,In_227);
nor U290 (N_290,In_23,In_612);
and U291 (N_291,In_578,In_734);
nand U292 (N_292,In_368,In_2);
nor U293 (N_293,In_102,In_429);
nor U294 (N_294,In_299,In_237);
nor U295 (N_295,In_213,In_167);
nand U296 (N_296,In_475,In_285);
and U297 (N_297,In_318,In_520);
or U298 (N_298,In_350,In_566);
or U299 (N_299,In_604,In_714);
nand U300 (N_300,In_9,In_424);
and U301 (N_301,In_399,In_207);
and U302 (N_302,In_484,In_219);
and U303 (N_303,In_526,In_577);
or U304 (N_304,In_564,In_17);
and U305 (N_305,In_229,In_197);
nand U306 (N_306,In_557,In_31);
or U307 (N_307,In_274,In_454);
nor U308 (N_308,In_126,In_541);
nor U309 (N_309,In_721,In_675);
nand U310 (N_310,In_689,In_594);
or U311 (N_311,In_221,In_702);
nor U312 (N_312,In_479,In_210);
nand U313 (N_313,In_728,In_477);
and U314 (N_314,In_136,In_19);
or U315 (N_315,In_208,In_246);
nand U316 (N_316,In_723,In_110);
or U317 (N_317,In_95,In_161);
xnor U318 (N_318,In_434,In_536);
nand U319 (N_319,In_217,In_553);
nor U320 (N_320,In_599,In_665);
or U321 (N_321,In_562,In_131);
xor U322 (N_322,In_82,In_74);
nand U323 (N_323,In_724,In_492);
and U324 (N_324,In_506,In_21);
nand U325 (N_325,In_378,In_306);
and U326 (N_326,In_462,In_419);
and U327 (N_327,In_646,In_704);
and U328 (N_328,In_740,In_218);
nor U329 (N_329,In_283,In_344);
nand U330 (N_330,In_596,In_472);
or U331 (N_331,In_671,In_407);
nand U332 (N_332,In_254,In_270);
nand U333 (N_333,In_700,In_575);
xor U334 (N_334,In_490,In_83);
nor U335 (N_335,In_277,In_140);
or U336 (N_336,In_159,In_255);
or U337 (N_337,In_582,In_91);
nand U338 (N_338,In_262,In_362);
and U339 (N_339,In_627,In_504);
or U340 (N_340,In_264,In_537);
nand U341 (N_341,In_684,In_138);
nand U342 (N_342,In_29,In_464);
or U343 (N_343,In_201,In_517);
and U344 (N_344,In_382,In_260);
nor U345 (N_345,In_590,In_137);
or U346 (N_346,In_620,In_85);
and U347 (N_347,In_357,In_712);
or U348 (N_348,In_316,In_119);
and U349 (N_349,In_108,In_560);
xnor U350 (N_350,In_610,In_615);
or U351 (N_351,In_180,In_631);
or U352 (N_352,In_502,In_275);
or U353 (N_353,In_222,In_127);
and U354 (N_354,In_147,In_18);
nor U355 (N_355,In_457,In_231);
and U356 (N_356,In_321,In_609);
and U357 (N_357,In_549,In_681);
nor U358 (N_358,In_281,In_215);
nor U359 (N_359,In_238,In_66);
or U360 (N_360,In_152,In_30);
and U361 (N_361,In_436,In_625);
nand U362 (N_362,In_748,In_35);
or U363 (N_363,In_515,In_519);
xnor U364 (N_364,In_448,In_735);
nand U365 (N_365,In_71,In_580);
nand U366 (N_366,In_220,In_78);
or U367 (N_367,In_680,In_685);
or U368 (N_368,In_336,In_507);
or U369 (N_369,In_720,In_341);
nand U370 (N_370,In_592,In_678);
nand U371 (N_371,In_269,In_356);
or U372 (N_372,In_496,In_413);
and U373 (N_373,In_730,In_166);
nor U374 (N_374,In_579,In_170);
nor U375 (N_375,In_251,In_374);
or U376 (N_376,In_63,In_157);
and U377 (N_377,In_662,In_77);
nor U378 (N_378,In_728,In_414);
and U379 (N_379,In_704,In_71);
nor U380 (N_380,In_162,In_340);
nand U381 (N_381,In_620,In_299);
nor U382 (N_382,In_621,In_225);
xor U383 (N_383,In_12,In_683);
or U384 (N_384,In_15,In_166);
and U385 (N_385,In_459,In_221);
nor U386 (N_386,In_328,In_173);
nand U387 (N_387,In_379,In_306);
and U388 (N_388,In_382,In_550);
or U389 (N_389,In_448,In_517);
or U390 (N_390,In_107,In_473);
or U391 (N_391,In_430,In_365);
nand U392 (N_392,In_547,In_96);
nor U393 (N_393,In_174,In_163);
or U394 (N_394,In_400,In_228);
or U395 (N_395,In_676,In_62);
nand U396 (N_396,In_78,In_671);
and U397 (N_397,In_382,In_309);
nor U398 (N_398,In_239,In_339);
nand U399 (N_399,In_267,In_310);
nor U400 (N_400,In_378,In_225);
and U401 (N_401,In_445,In_472);
or U402 (N_402,In_105,In_140);
nor U403 (N_403,In_110,In_504);
nor U404 (N_404,In_666,In_395);
nand U405 (N_405,In_217,In_670);
and U406 (N_406,In_393,In_243);
and U407 (N_407,In_678,In_180);
nor U408 (N_408,In_720,In_464);
nor U409 (N_409,In_629,In_615);
nand U410 (N_410,In_561,In_241);
and U411 (N_411,In_193,In_70);
nor U412 (N_412,In_351,In_580);
or U413 (N_413,In_646,In_304);
and U414 (N_414,In_22,In_674);
or U415 (N_415,In_298,In_15);
and U416 (N_416,In_223,In_526);
and U417 (N_417,In_288,In_523);
or U418 (N_418,In_273,In_412);
and U419 (N_419,In_743,In_724);
or U420 (N_420,In_434,In_712);
nand U421 (N_421,In_685,In_621);
nor U422 (N_422,In_64,In_31);
nand U423 (N_423,In_107,In_470);
or U424 (N_424,In_649,In_231);
or U425 (N_425,In_635,In_682);
and U426 (N_426,In_216,In_738);
and U427 (N_427,In_683,In_339);
nor U428 (N_428,In_343,In_734);
nand U429 (N_429,In_48,In_275);
and U430 (N_430,In_415,In_3);
or U431 (N_431,In_235,In_705);
or U432 (N_432,In_26,In_315);
and U433 (N_433,In_628,In_544);
or U434 (N_434,In_98,In_312);
xnor U435 (N_435,In_236,In_183);
or U436 (N_436,In_268,In_150);
nor U437 (N_437,In_310,In_78);
or U438 (N_438,In_166,In_91);
nand U439 (N_439,In_387,In_708);
and U440 (N_440,In_375,In_590);
and U441 (N_441,In_424,In_498);
nor U442 (N_442,In_468,In_168);
nor U443 (N_443,In_709,In_133);
nand U444 (N_444,In_539,In_289);
or U445 (N_445,In_223,In_250);
and U446 (N_446,In_429,In_655);
or U447 (N_447,In_469,In_694);
or U448 (N_448,In_140,In_598);
nor U449 (N_449,In_298,In_155);
or U450 (N_450,In_414,In_489);
nor U451 (N_451,In_383,In_242);
and U452 (N_452,In_204,In_561);
and U453 (N_453,In_586,In_379);
or U454 (N_454,In_183,In_670);
nor U455 (N_455,In_135,In_498);
nand U456 (N_456,In_196,In_657);
and U457 (N_457,In_702,In_71);
nand U458 (N_458,In_737,In_277);
or U459 (N_459,In_332,In_623);
and U460 (N_460,In_266,In_15);
and U461 (N_461,In_154,In_106);
and U462 (N_462,In_491,In_0);
nor U463 (N_463,In_578,In_468);
or U464 (N_464,In_366,In_225);
nor U465 (N_465,In_205,In_519);
or U466 (N_466,In_360,In_349);
nor U467 (N_467,In_613,In_242);
nor U468 (N_468,In_182,In_284);
nor U469 (N_469,In_591,In_594);
nor U470 (N_470,In_642,In_724);
nor U471 (N_471,In_208,In_199);
and U472 (N_472,In_371,In_315);
nand U473 (N_473,In_503,In_151);
nand U474 (N_474,In_426,In_333);
and U475 (N_475,In_667,In_3);
nor U476 (N_476,In_210,In_577);
nand U477 (N_477,In_207,In_176);
nand U478 (N_478,In_94,In_26);
or U479 (N_479,In_6,In_321);
nor U480 (N_480,In_613,In_541);
or U481 (N_481,In_24,In_164);
nand U482 (N_482,In_388,In_632);
or U483 (N_483,In_8,In_453);
nor U484 (N_484,In_519,In_619);
nand U485 (N_485,In_682,In_144);
nand U486 (N_486,In_364,In_425);
or U487 (N_487,In_112,In_608);
xor U488 (N_488,In_726,In_470);
nor U489 (N_489,In_229,In_603);
nor U490 (N_490,In_728,In_464);
nand U491 (N_491,In_498,In_471);
or U492 (N_492,In_97,In_688);
or U493 (N_493,In_205,In_717);
and U494 (N_494,In_663,In_435);
or U495 (N_495,In_279,In_28);
nor U496 (N_496,In_459,In_403);
or U497 (N_497,In_302,In_515);
or U498 (N_498,In_608,In_152);
or U499 (N_499,In_372,In_682);
or U500 (N_500,N_66,N_401);
nor U501 (N_501,N_187,N_125);
nand U502 (N_502,N_152,N_90);
xnor U503 (N_503,N_218,N_161);
or U504 (N_504,N_157,N_143);
and U505 (N_505,N_131,N_438);
and U506 (N_506,N_198,N_23);
nand U507 (N_507,N_113,N_81);
nand U508 (N_508,N_459,N_291);
and U509 (N_509,N_282,N_83);
nand U510 (N_510,N_457,N_173);
nor U511 (N_511,N_384,N_179);
nand U512 (N_512,N_15,N_123);
nand U513 (N_513,N_344,N_59);
or U514 (N_514,N_16,N_400);
and U515 (N_515,N_73,N_463);
or U516 (N_516,N_475,N_424);
nand U517 (N_517,N_281,N_102);
or U518 (N_518,N_294,N_144);
nand U519 (N_519,N_120,N_452);
nor U520 (N_520,N_350,N_174);
nor U521 (N_521,N_255,N_379);
or U522 (N_522,N_377,N_347);
or U523 (N_523,N_56,N_65);
and U524 (N_524,N_52,N_7);
and U525 (N_525,N_54,N_462);
and U526 (N_526,N_469,N_220);
and U527 (N_527,N_481,N_437);
nand U528 (N_528,N_349,N_235);
or U529 (N_529,N_177,N_62);
or U530 (N_530,N_12,N_250);
nand U531 (N_531,N_151,N_121);
xor U532 (N_532,N_86,N_35);
nor U533 (N_533,N_9,N_283);
or U534 (N_534,N_210,N_140);
nor U535 (N_535,N_323,N_136);
or U536 (N_536,N_486,N_166);
or U537 (N_537,N_146,N_28);
or U538 (N_538,N_404,N_48);
nand U539 (N_539,N_130,N_163);
nor U540 (N_540,N_359,N_270);
nand U541 (N_541,N_362,N_178);
nand U542 (N_542,N_190,N_422);
and U543 (N_543,N_464,N_292);
nand U544 (N_544,N_162,N_388);
nor U545 (N_545,N_318,N_216);
and U546 (N_546,N_207,N_293);
nand U547 (N_547,N_105,N_399);
nor U548 (N_548,N_180,N_407);
or U549 (N_549,N_484,N_149);
and U550 (N_550,N_492,N_249);
nor U551 (N_551,N_355,N_443);
and U552 (N_552,N_31,N_203);
nand U553 (N_553,N_34,N_251);
nand U554 (N_554,N_369,N_159);
or U555 (N_555,N_8,N_253);
and U556 (N_556,N_106,N_184);
nor U557 (N_557,N_188,N_317);
or U558 (N_558,N_273,N_238);
and U559 (N_559,N_169,N_389);
and U560 (N_560,N_122,N_1);
or U561 (N_561,N_425,N_470);
nor U562 (N_562,N_234,N_468);
or U563 (N_563,N_473,N_372);
nand U564 (N_564,N_435,N_27);
and U565 (N_565,N_440,N_418);
and U566 (N_566,N_115,N_441);
nand U567 (N_567,N_415,N_303);
and U568 (N_568,N_431,N_398);
or U569 (N_569,N_236,N_211);
nand U570 (N_570,N_320,N_154);
or U571 (N_571,N_454,N_204);
and U572 (N_572,N_447,N_380);
and U573 (N_573,N_314,N_432);
xnor U574 (N_574,N_20,N_206);
and U575 (N_575,N_313,N_370);
nor U576 (N_576,N_227,N_279);
nor U577 (N_577,N_107,N_57);
nand U578 (N_578,N_499,N_6);
nand U579 (N_579,N_256,N_332);
or U580 (N_580,N_44,N_358);
nor U581 (N_581,N_479,N_112);
nor U582 (N_582,N_199,N_406);
and U583 (N_583,N_191,N_386);
nor U584 (N_584,N_427,N_259);
nor U585 (N_585,N_11,N_382);
and U586 (N_586,N_480,N_476);
nand U587 (N_587,N_272,N_421);
xnor U588 (N_588,N_465,N_45);
or U589 (N_589,N_153,N_391);
or U590 (N_590,N_101,N_30);
nor U591 (N_591,N_74,N_63);
nor U592 (N_592,N_429,N_430);
and U593 (N_593,N_69,N_47);
nor U594 (N_594,N_232,N_129);
and U595 (N_595,N_110,N_396);
and U596 (N_596,N_26,N_436);
or U597 (N_597,N_82,N_330);
or U598 (N_598,N_319,N_497);
or U599 (N_599,N_245,N_375);
nand U600 (N_600,N_61,N_127);
xnor U601 (N_601,N_395,N_37);
nor U602 (N_602,N_21,N_394);
nand U603 (N_603,N_420,N_116);
nand U604 (N_604,N_247,N_142);
nand U605 (N_605,N_13,N_495);
and U606 (N_606,N_494,N_439);
or U607 (N_607,N_94,N_242);
nor U608 (N_608,N_402,N_84);
or U609 (N_609,N_450,N_434);
or U610 (N_610,N_442,N_186);
and U611 (N_611,N_53,N_241);
and U612 (N_612,N_147,N_298);
xnor U613 (N_613,N_328,N_285);
and U614 (N_614,N_222,N_171);
nand U615 (N_615,N_364,N_240);
and U616 (N_616,N_351,N_77);
nor U617 (N_617,N_296,N_280);
and U618 (N_618,N_458,N_416);
or U619 (N_619,N_490,N_10);
or U620 (N_620,N_327,N_145);
or U621 (N_621,N_378,N_5);
nor U622 (N_622,N_194,N_267);
or U623 (N_623,N_217,N_2);
nor U624 (N_624,N_325,N_55);
nand U625 (N_625,N_239,N_111);
or U626 (N_626,N_271,N_445);
xor U627 (N_627,N_338,N_329);
nor U628 (N_628,N_284,N_76);
or U629 (N_629,N_301,N_138);
nand U630 (N_630,N_353,N_118);
nor U631 (N_631,N_97,N_170);
or U632 (N_632,N_451,N_262);
and U633 (N_633,N_100,N_354);
nand U634 (N_634,N_117,N_444);
nand U635 (N_635,N_258,N_172);
and U636 (N_636,N_288,N_383);
nand U637 (N_637,N_29,N_41);
and U638 (N_638,N_201,N_365);
and U639 (N_639,N_336,N_104);
nand U640 (N_640,N_189,N_374);
nand U641 (N_641,N_43,N_150);
and U642 (N_642,N_40,N_334);
nand U643 (N_643,N_483,N_363);
or U644 (N_644,N_64,N_265);
nand U645 (N_645,N_167,N_79);
or U646 (N_646,N_185,N_75);
or U647 (N_647,N_335,N_196);
nand U648 (N_648,N_89,N_299);
or U649 (N_649,N_51,N_132);
and U650 (N_650,N_304,N_148);
or U651 (N_651,N_164,N_496);
and U652 (N_652,N_460,N_228);
nor U653 (N_653,N_230,N_96);
and U654 (N_654,N_19,N_278);
and U655 (N_655,N_307,N_139);
or U656 (N_656,N_60,N_70);
or U657 (N_657,N_345,N_205);
or U658 (N_658,N_192,N_485);
or U659 (N_659,N_175,N_126);
nor U660 (N_660,N_300,N_393);
nand U661 (N_661,N_254,N_333);
nand U662 (N_662,N_478,N_493);
or U663 (N_663,N_103,N_133);
nor U664 (N_664,N_233,N_331);
nand U665 (N_665,N_448,N_474);
or U666 (N_666,N_3,N_455);
and U667 (N_667,N_346,N_263);
and U668 (N_668,N_489,N_165);
or U669 (N_669,N_356,N_456);
or U670 (N_670,N_276,N_176);
or U671 (N_671,N_33,N_309);
nor U672 (N_672,N_22,N_397);
and U673 (N_673,N_321,N_326);
nor U674 (N_674,N_17,N_38);
nand U675 (N_675,N_260,N_36);
or U676 (N_676,N_295,N_310);
nand U677 (N_677,N_18,N_141);
nor U678 (N_678,N_417,N_32);
nand U679 (N_679,N_261,N_498);
and U680 (N_680,N_467,N_376);
and U681 (N_681,N_305,N_412);
or U682 (N_682,N_58,N_99);
or U683 (N_683,N_49,N_72);
nand U684 (N_684,N_315,N_67);
nand U685 (N_685,N_231,N_366);
or U686 (N_686,N_252,N_472);
and U687 (N_687,N_368,N_24);
nor U688 (N_688,N_109,N_392);
nand U689 (N_689,N_491,N_428);
and U690 (N_690,N_373,N_208);
nor U691 (N_691,N_182,N_277);
and U692 (N_692,N_266,N_357);
nor U693 (N_693,N_168,N_246);
nand U694 (N_694,N_243,N_135);
nand U695 (N_695,N_248,N_257);
or U696 (N_696,N_223,N_411);
or U697 (N_697,N_488,N_487);
and U698 (N_698,N_155,N_446);
and U699 (N_699,N_200,N_87);
nand U700 (N_700,N_324,N_92);
and U701 (N_701,N_25,N_156);
nor U702 (N_702,N_337,N_95);
nand U703 (N_703,N_371,N_46);
and U704 (N_704,N_449,N_409);
and U705 (N_705,N_426,N_181);
nand U706 (N_706,N_114,N_237);
and U707 (N_707,N_405,N_80);
and U708 (N_708,N_134,N_229);
or U709 (N_709,N_306,N_224);
nor U710 (N_710,N_202,N_322);
or U711 (N_711,N_119,N_341);
nand U712 (N_712,N_312,N_286);
nand U713 (N_713,N_453,N_225);
nand U714 (N_714,N_423,N_352);
nor U715 (N_715,N_197,N_264);
nand U716 (N_716,N_71,N_195);
and U717 (N_717,N_42,N_466);
and U718 (N_718,N_93,N_269);
nor U719 (N_719,N_124,N_311);
and U720 (N_720,N_244,N_0);
nor U721 (N_721,N_482,N_4);
or U722 (N_722,N_137,N_128);
nand U723 (N_723,N_477,N_78);
or U724 (N_724,N_343,N_214);
or U725 (N_725,N_433,N_226);
nand U726 (N_726,N_360,N_160);
and U727 (N_727,N_410,N_39);
and U728 (N_728,N_297,N_471);
and U729 (N_729,N_339,N_14);
or U730 (N_730,N_91,N_414);
nor U731 (N_731,N_88,N_390);
nor U732 (N_732,N_268,N_183);
nor U733 (N_733,N_387,N_221);
nor U734 (N_734,N_275,N_408);
and U735 (N_735,N_308,N_289);
and U736 (N_736,N_403,N_348);
nor U737 (N_737,N_287,N_219);
or U738 (N_738,N_419,N_193);
nand U739 (N_739,N_108,N_213);
and U740 (N_740,N_158,N_367);
and U741 (N_741,N_209,N_98);
or U742 (N_742,N_381,N_302);
and U743 (N_743,N_50,N_342);
or U744 (N_744,N_274,N_361);
xor U745 (N_745,N_212,N_290);
nand U746 (N_746,N_215,N_340);
nor U747 (N_747,N_385,N_68);
nand U748 (N_748,N_85,N_461);
nor U749 (N_749,N_413,N_316);
nor U750 (N_750,N_291,N_311);
nor U751 (N_751,N_437,N_32);
or U752 (N_752,N_277,N_160);
nand U753 (N_753,N_189,N_290);
nor U754 (N_754,N_369,N_238);
or U755 (N_755,N_300,N_443);
nor U756 (N_756,N_366,N_462);
or U757 (N_757,N_428,N_66);
nor U758 (N_758,N_300,N_372);
xor U759 (N_759,N_48,N_471);
nand U760 (N_760,N_122,N_191);
nand U761 (N_761,N_272,N_266);
nand U762 (N_762,N_48,N_129);
or U763 (N_763,N_491,N_1);
nor U764 (N_764,N_334,N_165);
nor U765 (N_765,N_75,N_21);
and U766 (N_766,N_298,N_78);
nor U767 (N_767,N_20,N_40);
nor U768 (N_768,N_312,N_212);
nand U769 (N_769,N_270,N_276);
nor U770 (N_770,N_209,N_367);
nand U771 (N_771,N_135,N_171);
or U772 (N_772,N_248,N_94);
or U773 (N_773,N_321,N_262);
xor U774 (N_774,N_355,N_133);
nor U775 (N_775,N_296,N_90);
nand U776 (N_776,N_253,N_312);
or U777 (N_777,N_84,N_332);
nand U778 (N_778,N_316,N_362);
xor U779 (N_779,N_429,N_352);
nand U780 (N_780,N_219,N_446);
or U781 (N_781,N_296,N_113);
or U782 (N_782,N_264,N_133);
and U783 (N_783,N_133,N_456);
and U784 (N_784,N_174,N_39);
nor U785 (N_785,N_472,N_486);
and U786 (N_786,N_203,N_299);
nor U787 (N_787,N_239,N_181);
or U788 (N_788,N_479,N_484);
xnor U789 (N_789,N_130,N_59);
and U790 (N_790,N_355,N_110);
nand U791 (N_791,N_222,N_422);
nand U792 (N_792,N_333,N_451);
and U793 (N_793,N_278,N_110);
nor U794 (N_794,N_232,N_140);
or U795 (N_795,N_194,N_50);
xor U796 (N_796,N_395,N_314);
or U797 (N_797,N_152,N_128);
or U798 (N_798,N_488,N_352);
nand U799 (N_799,N_136,N_193);
nand U800 (N_800,N_475,N_260);
nand U801 (N_801,N_350,N_204);
and U802 (N_802,N_6,N_80);
nand U803 (N_803,N_187,N_441);
xnor U804 (N_804,N_416,N_241);
or U805 (N_805,N_470,N_245);
or U806 (N_806,N_196,N_109);
nand U807 (N_807,N_31,N_17);
or U808 (N_808,N_404,N_364);
nor U809 (N_809,N_63,N_80);
or U810 (N_810,N_210,N_334);
nand U811 (N_811,N_447,N_303);
or U812 (N_812,N_201,N_455);
nor U813 (N_813,N_131,N_468);
nand U814 (N_814,N_81,N_161);
or U815 (N_815,N_453,N_234);
or U816 (N_816,N_235,N_238);
nor U817 (N_817,N_178,N_439);
or U818 (N_818,N_496,N_19);
and U819 (N_819,N_79,N_352);
nand U820 (N_820,N_305,N_149);
and U821 (N_821,N_207,N_338);
nor U822 (N_822,N_12,N_71);
or U823 (N_823,N_114,N_497);
nor U824 (N_824,N_435,N_122);
nand U825 (N_825,N_135,N_463);
or U826 (N_826,N_334,N_46);
nand U827 (N_827,N_364,N_147);
nand U828 (N_828,N_224,N_276);
and U829 (N_829,N_403,N_440);
or U830 (N_830,N_80,N_49);
nor U831 (N_831,N_194,N_302);
or U832 (N_832,N_21,N_342);
nand U833 (N_833,N_254,N_127);
nor U834 (N_834,N_288,N_265);
nand U835 (N_835,N_151,N_293);
or U836 (N_836,N_342,N_48);
nand U837 (N_837,N_231,N_246);
or U838 (N_838,N_198,N_201);
and U839 (N_839,N_151,N_105);
nor U840 (N_840,N_249,N_129);
nor U841 (N_841,N_178,N_237);
nand U842 (N_842,N_462,N_384);
and U843 (N_843,N_248,N_333);
nand U844 (N_844,N_80,N_243);
nor U845 (N_845,N_287,N_451);
or U846 (N_846,N_367,N_66);
nand U847 (N_847,N_44,N_112);
nor U848 (N_848,N_159,N_318);
or U849 (N_849,N_305,N_119);
and U850 (N_850,N_94,N_53);
nand U851 (N_851,N_17,N_7);
nor U852 (N_852,N_270,N_338);
nor U853 (N_853,N_471,N_230);
nand U854 (N_854,N_465,N_229);
nand U855 (N_855,N_7,N_177);
xor U856 (N_856,N_320,N_221);
or U857 (N_857,N_491,N_67);
nand U858 (N_858,N_403,N_164);
nand U859 (N_859,N_60,N_134);
nand U860 (N_860,N_56,N_269);
or U861 (N_861,N_344,N_458);
nor U862 (N_862,N_145,N_345);
nand U863 (N_863,N_280,N_250);
nand U864 (N_864,N_367,N_419);
and U865 (N_865,N_252,N_259);
nand U866 (N_866,N_96,N_194);
or U867 (N_867,N_366,N_330);
and U868 (N_868,N_114,N_192);
or U869 (N_869,N_181,N_153);
nor U870 (N_870,N_412,N_158);
or U871 (N_871,N_385,N_297);
nor U872 (N_872,N_222,N_365);
and U873 (N_873,N_123,N_156);
or U874 (N_874,N_276,N_490);
and U875 (N_875,N_125,N_299);
or U876 (N_876,N_248,N_448);
nand U877 (N_877,N_463,N_415);
nor U878 (N_878,N_95,N_58);
or U879 (N_879,N_146,N_137);
or U880 (N_880,N_257,N_251);
or U881 (N_881,N_300,N_294);
nor U882 (N_882,N_134,N_84);
and U883 (N_883,N_292,N_236);
nor U884 (N_884,N_116,N_414);
nand U885 (N_885,N_12,N_473);
nand U886 (N_886,N_310,N_280);
nand U887 (N_887,N_187,N_129);
and U888 (N_888,N_460,N_100);
nand U889 (N_889,N_465,N_160);
and U890 (N_890,N_257,N_218);
and U891 (N_891,N_287,N_128);
and U892 (N_892,N_149,N_389);
or U893 (N_893,N_323,N_398);
nor U894 (N_894,N_449,N_301);
and U895 (N_895,N_313,N_159);
nor U896 (N_896,N_426,N_240);
nand U897 (N_897,N_426,N_43);
or U898 (N_898,N_221,N_346);
or U899 (N_899,N_429,N_424);
nor U900 (N_900,N_133,N_6);
and U901 (N_901,N_478,N_383);
nand U902 (N_902,N_374,N_262);
and U903 (N_903,N_370,N_465);
nor U904 (N_904,N_339,N_180);
nand U905 (N_905,N_287,N_480);
and U906 (N_906,N_158,N_197);
nand U907 (N_907,N_292,N_162);
nand U908 (N_908,N_166,N_330);
and U909 (N_909,N_10,N_51);
nand U910 (N_910,N_181,N_24);
nand U911 (N_911,N_308,N_101);
or U912 (N_912,N_45,N_25);
or U913 (N_913,N_88,N_444);
nand U914 (N_914,N_474,N_472);
nand U915 (N_915,N_60,N_69);
and U916 (N_916,N_425,N_364);
nor U917 (N_917,N_259,N_34);
and U918 (N_918,N_181,N_220);
nand U919 (N_919,N_252,N_192);
and U920 (N_920,N_310,N_127);
and U921 (N_921,N_263,N_378);
nor U922 (N_922,N_212,N_306);
or U923 (N_923,N_190,N_421);
or U924 (N_924,N_298,N_462);
and U925 (N_925,N_82,N_114);
and U926 (N_926,N_89,N_402);
and U927 (N_927,N_244,N_217);
nor U928 (N_928,N_177,N_216);
or U929 (N_929,N_305,N_273);
or U930 (N_930,N_157,N_316);
or U931 (N_931,N_247,N_310);
nand U932 (N_932,N_404,N_417);
nor U933 (N_933,N_123,N_260);
xnor U934 (N_934,N_185,N_129);
nand U935 (N_935,N_426,N_215);
nor U936 (N_936,N_422,N_106);
nor U937 (N_937,N_78,N_317);
nor U938 (N_938,N_6,N_205);
and U939 (N_939,N_26,N_254);
and U940 (N_940,N_338,N_389);
nand U941 (N_941,N_142,N_280);
or U942 (N_942,N_128,N_256);
nand U943 (N_943,N_71,N_269);
nand U944 (N_944,N_424,N_167);
or U945 (N_945,N_396,N_381);
and U946 (N_946,N_269,N_48);
and U947 (N_947,N_169,N_494);
or U948 (N_948,N_437,N_238);
and U949 (N_949,N_322,N_194);
or U950 (N_950,N_9,N_49);
and U951 (N_951,N_364,N_133);
and U952 (N_952,N_245,N_216);
and U953 (N_953,N_181,N_165);
nor U954 (N_954,N_398,N_21);
nand U955 (N_955,N_287,N_286);
nand U956 (N_956,N_345,N_317);
nor U957 (N_957,N_180,N_194);
nor U958 (N_958,N_178,N_331);
nand U959 (N_959,N_144,N_175);
or U960 (N_960,N_160,N_221);
and U961 (N_961,N_491,N_217);
nor U962 (N_962,N_76,N_211);
nand U963 (N_963,N_439,N_491);
nor U964 (N_964,N_8,N_63);
or U965 (N_965,N_298,N_287);
nand U966 (N_966,N_278,N_153);
or U967 (N_967,N_428,N_338);
nand U968 (N_968,N_233,N_99);
and U969 (N_969,N_88,N_348);
nand U970 (N_970,N_374,N_485);
or U971 (N_971,N_242,N_23);
nand U972 (N_972,N_126,N_461);
nand U973 (N_973,N_23,N_175);
and U974 (N_974,N_168,N_236);
or U975 (N_975,N_150,N_225);
or U976 (N_976,N_411,N_302);
nor U977 (N_977,N_487,N_483);
nor U978 (N_978,N_363,N_262);
or U979 (N_979,N_105,N_381);
nand U980 (N_980,N_236,N_213);
nand U981 (N_981,N_439,N_45);
nor U982 (N_982,N_209,N_362);
or U983 (N_983,N_221,N_347);
or U984 (N_984,N_393,N_23);
nor U985 (N_985,N_467,N_45);
or U986 (N_986,N_122,N_256);
nor U987 (N_987,N_399,N_363);
and U988 (N_988,N_265,N_163);
or U989 (N_989,N_34,N_272);
or U990 (N_990,N_159,N_138);
nor U991 (N_991,N_52,N_33);
nand U992 (N_992,N_499,N_106);
nor U993 (N_993,N_1,N_407);
nand U994 (N_994,N_6,N_105);
or U995 (N_995,N_322,N_125);
and U996 (N_996,N_19,N_323);
or U997 (N_997,N_279,N_197);
or U998 (N_998,N_268,N_207);
nor U999 (N_999,N_161,N_86);
and U1000 (N_1000,N_773,N_828);
and U1001 (N_1001,N_730,N_623);
nand U1002 (N_1002,N_936,N_832);
nor U1003 (N_1003,N_666,N_823);
nor U1004 (N_1004,N_541,N_703);
or U1005 (N_1005,N_903,N_533);
or U1006 (N_1006,N_977,N_993);
or U1007 (N_1007,N_561,N_725);
nor U1008 (N_1008,N_749,N_577);
nor U1009 (N_1009,N_945,N_804);
nand U1010 (N_1010,N_879,N_991);
nor U1011 (N_1011,N_846,N_701);
nor U1012 (N_1012,N_967,N_508);
or U1013 (N_1013,N_691,N_658);
nor U1014 (N_1014,N_865,N_517);
nand U1015 (N_1015,N_621,N_891);
nor U1016 (N_1016,N_969,N_628);
and U1017 (N_1017,N_767,N_734);
nand U1018 (N_1018,N_932,N_751);
nor U1019 (N_1019,N_952,N_852);
or U1020 (N_1020,N_567,N_896);
or U1021 (N_1021,N_801,N_984);
nor U1022 (N_1022,N_604,N_797);
and U1023 (N_1023,N_563,N_880);
or U1024 (N_1024,N_715,N_868);
nand U1025 (N_1025,N_862,N_968);
nor U1026 (N_1026,N_694,N_783);
nand U1027 (N_1027,N_627,N_927);
and U1028 (N_1028,N_809,N_673);
nor U1029 (N_1029,N_720,N_521);
or U1030 (N_1030,N_559,N_842);
and U1031 (N_1031,N_959,N_500);
or U1032 (N_1032,N_939,N_989);
or U1033 (N_1033,N_682,N_651);
nand U1034 (N_1034,N_883,N_978);
and U1035 (N_1035,N_565,N_585);
or U1036 (N_1036,N_740,N_607);
and U1037 (N_1037,N_768,N_550);
nor U1038 (N_1038,N_830,N_934);
nand U1039 (N_1039,N_716,N_683);
nand U1040 (N_1040,N_547,N_839);
and U1041 (N_1041,N_856,N_753);
nand U1042 (N_1042,N_670,N_906);
or U1043 (N_1043,N_609,N_810);
and U1044 (N_1044,N_871,N_546);
or U1045 (N_1045,N_723,N_955);
nand U1046 (N_1046,N_974,N_829);
nor U1047 (N_1047,N_631,N_921);
and U1048 (N_1048,N_728,N_573);
nor U1049 (N_1049,N_746,N_739);
xnor U1050 (N_1050,N_877,N_685);
nor U1051 (N_1051,N_820,N_827);
nor U1052 (N_1052,N_910,N_617);
and U1053 (N_1053,N_745,N_613);
and U1054 (N_1054,N_888,N_931);
nor U1055 (N_1055,N_900,N_679);
and U1056 (N_1056,N_553,N_853);
nor U1057 (N_1057,N_712,N_596);
nand U1058 (N_1058,N_755,N_776);
and U1059 (N_1059,N_634,N_743);
or U1060 (N_1060,N_710,N_992);
xnor U1061 (N_1061,N_807,N_702);
and U1062 (N_1062,N_618,N_624);
or U1063 (N_1063,N_652,N_733);
or U1064 (N_1064,N_552,N_873);
and U1065 (N_1065,N_953,N_878);
and U1066 (N_1066,N_537,N_648);
and U1067 (N_1067,N_835,N_539);
nor U1068 (N_1068,N_695,N_737);
and U1069 (N_1069,N_824,N_686);
and U1070 (N_1070,N_971,N_844);
or U1071 (N_1071,N_731,N_678);
nand U1072 (N_1072,N_518,N_980);
nor U1073 (N_1073,N_528,N_660);
and U1074 (N_1074,N_812,N_764);
nor U1075 (N_1075,N_503,N_549);
or U1076 (N_1076,N_647,N_640);
and U1077 (N_1077,N_704,N_510);
and U1078 (N_1078,N_570,N_988);
nor U1079 (N_1079,N_770,N_905);
and U1080 (N_1080,N_895,N_719);
and U1081 (N_1081,N_632,N_775);
nor U1082 (N_1082,N_555,N_505);
and U1083 (N_1083,N_635,N_795);
and U1084 (N_1084,N_736,N_982);
and U1085 (N_1085,N_506,N_501);
or U1086 (N_1086,N_522,N_851);
nand U1087 (N_1087,N_688,N_709);
and U1088 (N_1088,N_697,N_571);
or U1089 (N_1089,N_645,N_881);
and U1090 (N_1090,N_575,N_706);
nor U1091 (N_1091,N_630,N_664);
nor U1092 (N_1092,N_983,N_930);
nor U1093 (N_1093,N_512,N_513);
nor U1094 (N_1094,N_687,N_885);
or U1095 (N_1095,N_909,N_857);
nor U1096 (N_1096,N_556,N_754);
nor U1097 (N_1097,N_920,N_580);
or U1098 (N_1098,N_833,N_538);
or U1099 (N_1099,N_592,N_629);
or U1100 (N_1100,N_961,N_574);
nor U1101 (N_1101,N_562,N_707);
nor U1102 (N_1102,N_884,N_711);
nor U1103 (N_1103,N_886,N_898);
or U1104 (N_1104,N_855,N_717);
or U1105 (N_1105,N_787,N_525);
nor U1106 (N_1106,N_665,N_843);
or U1107 (N_1107,N_826,N_515);
and U1108 (N_1108,N_625,N_560);
or U1109 (N_1109,N_591,N_511);
or U1110 (N_1110,N_803,N_774);
and U1111 (N_1111,N_662,N_516);
or U1112 (N_1112,N_684,N_698);
nor U1113 (N_1113,N_756,N_780);
nand U1114 (N_1114,N_994,N_784);
and U1115 (N_1115,N_760,N_849);
and U1116 (N_1116,N_966,N_817);
nand U1117 (N_1117,N_970,N_502);
nand U1118 (N_1118,N_946,N_638);
nand U1119 (N_1119,N_578,N_779);
or U1120 (N_1120,N_519,N_527);
and U1121 (N_1121,N_860,N_566);
or U1122 (N_1122,N_981,N_656);
or U1123 (N_1123,N_786,N_785);
nor U1124 (N_1124,N_700,N_811);
nand U1125 (N_1125,N_752,N_689);
nor U1126 (N_1126,N_606,N_761);
or U1127 (N_1127,N_897,N_996);
or U1128 (N_1128,N_864,N_813);
nor U1129 (N_1129,N_986,N_821);
nand U1130 (N_1130,N_997,N_777);
nand U1131 (N_1131,N_536,N_680);
or U1132 (N_1132,N_637,N_799);
nor U1133 (N_1133,N_985,N_861);
nor U1134 (N_1134,N_845,N_890);
nand U1135 (N_1135,N_766,N_584);
nor U1136 (N_1136,N_876,N_741);
nand U1137 (N_1137,N_998,N_520);
nand U1138 (N_1138,N_605,N_659);
and U1139 (N_1139,N_887,N_894);
nor U1140 (N_1140,N_612,N_672);
nor U1141 (N_1141,N_935,N_912);
nor U1142 (N_1142,N_579,N_973);
or U1143 (N_1143,N_972,N_681);
nor U1144 (N_1144,N_708,N_557);
or U1145 (N_1145,N_558,N_526);
nand U1146 (N_1146,N_742,N_507);
and U1147 (N_1147,N_763,N_610);
nand U1148 (N_1148,N_951,N_913);
and U1149 (N_1149,N_722,N_590);
and U1150 (N_1150,N_616,N_564);
nand U1151 (N_1151,N_714,N_958);
or U1152 (N_1152,N_948,N_671);
nand U1153 (N_1153,N_915,N_765);
or U1154 (N_1154,N_940,N_987);
and U1155 (N_1155,N_944,N_954);
or U1156 (N_1156,N_854,N_990);
nand U1157 (N_1157,N_595,N_837);
and U1158 (N_1158,N_923,N_601);
and U1159 (N_1159,N_841,N_794);
and U1160 (N_1160,N_790,N_614);
nand U1161 (N_1161,N_622,N_646);
and U1162 (N_1162,N_676,N_863);
nor U1163 (N_1163,N_836,N_545);
nor U1164 (N_1164,N_576,N_781);
nor U1165 (N_1165,N_892,N_732);
or U1166 (N_1166,N_534,N_875);
and U1167 (N_1167,N_729,N_509);
or U1168 (N_1168,N_544,N_995);
and U1169 (N_1169,N_802,N_872);
or U1170 (N_1170,N_619,N_769);
nand U1171 (N_1171,N_963,N_568);
nor U1172 (N_1172,N_911,N_735);
and U1173 (N_1173,N_999,N_788);
or U1174 (N_1174,N_942,N_960);
or U1175 (N_1175,N_599,N_800);
or U1176 (N_1176,N_908,N_747);
and U1177 (N_1177,N_918,N_589);
and U1178 (N_1178,N_615,N_705);
or U1179 (N_1179,N_639,N_620);
or U1180 (N_1180,N_548,N_805);
xor U1181 (N_1181,N_975,N_713);
nand U1182 (N_1182,N_693,N_882);
or U1183 (N_1183,N_937,N_667);
nor U1184 (N_1184,N_523,N_602);
nand U1185 (N_1185,N_793,N_586);
and U1186 (N_1186,N_772,N_956);
or U1187 (N_1187,N_831,N_692);
nand U1188 (N_1188,N_641,N_529);
nand U1189 (N_1189,N_941,N_587);
nand U1190 (N_1190,N_924,N_626);
nor U1191 (N_1191,N_581,N_850);
or U1192 (N_1192,N_504,N_950);
nand U1193 (N_1193,N_674,N_771);
or U1194 (N_1194,N_919,N_928);
and U1195 (N_1195,N_916,N_738);
nand U1196 (N_1196,N_866,N_904);
nor U1197 (N_1197,N_531,N_814);
and U1198 (N_1198,N_762,N_668);
or U1199 (N_1199,N_840,N_902);
xor U1200 (N_1200,N_653,N_778);
nor U1201 (N_1201,N_543,N_669);
nand U1202 (N_1202,N_791,N_644);
nand U1203 (N_1203,N_650,N_907);
nor U1204 (N_1204,N_816,N_929);
or U1205 (N_1205,N_655,N_677);
nand U1206 (N_1206,N_654,N_914);
nand U1207 (N_1207,N_847,N_750);
or U1208 (N_1208,N_572,N_597);
nand U1209 (N_1209,N_661,N_893);
xnor U1210 (N_1210,N_796,N_726);
nor U1211 (N_1211,N_757,N_696);
nor U1212 (N_1212,N_808,N_569);
nor U1213 (N_1213,N_643,N_699);
and U1214 (N_1214,N_593,N_925);
nor U1215 (N_1215,N_798,N_542);
and U1216 (N_1216,N_514,N_869);
nor U1217 (N_1217,N_551,N_806);
nand U1218 (N_1218,N_964,N_949);
and U1219 (N_1219,N_976,N_834);
nor U1220 (N_1220,N_594,N_957);
nor U1221 (N_1221,N_926,N_782);
or U1222 (N_1222,N_727,N_965);
nand U1223 (N_1223,N_663,N_748);
nor U1224 (N_1224,N_943,N_867);
or U1225 (N_1225,N_858,N_822);
and U1226 (N_1226,N_608,N_582);
and U1227 (N_1227,N_583,N_917);
and U1228 (N_1228,N_721,N_838);
or U1229 (N_1229,N_524,N_899);
nand U1230 (N_1230,N_870,N_611);
nor U1231 (N_1231,N_598,N_554);
nor U1232 (N_1232,N_815,N_759);
or U1233 (N_1233,N_744,N_718);
nor U1234 (N_1234,N_535,N_633);
nor U1235 (N_1235,N_922,N_532);
nand U1236 (N_1236,N_649,N_825);
or U1237 (N_1237,N_603,N_933);
and U1238 (N_1238,N_979,N_938);
nor U1239 (N_1239,N_962,N_848);
or U1240 (N_1240,N_724,N_758);
nand U1241 (N_1241,N_540,N_642);
or U1242 (N_1242,N_636,N_818);
nand U1243 (N_1243,N_675,N_588);
and U1244 (N_1244,N_874,N_901);
or U1245 (N_1245,N_947,N_792);
nor U1246 (N_1246,N_859,N_690);
nor U1247 (N_1247,N_600,N_889);
nand U1248 (N_1248,N_819,N_530);
nand U1249 (N_1249,N_789,N_657);
nor U1250 (N_1250,N_970,N_582);
and U1251 (N_1251,N_842,N_730);
or U1252 (N_1252,N_825,N_918);
nand U1253 (N_1253,N_961,N_648);
nand U1254 (N_1254,N_562,N_871);
nor U1255 (N_1255,N_842,N_719);
nand U1256 (N_1256,N_745,N_602);
or U1257 (N_1257,N_927,N_594);
nand U1258 (N_1258,N_596,N_594);
or U1259 (N_1259,N_841,N_943);
nand U1260 (N_1260,N_531,N_672);
nor U1261 (N_1261,N_603,N_851);
nor U1262 (N_1262,N_807,N_923);
nor U1263 (N_1263,N_796,N_868);
nor U1264 (N_1264,N_883,N_844);
and U1265 (N_1265,N_774,N_607);
nand U1266 (N_1266,N_926,N_731);
nor U1267 (N_1267,N_658,N_768);
and U1268 (N_1268,N_773,N_956);
nand U1269 (N_1269,N_803,N_970);
nor U1270 (N_1270,N_972,N_803);
and U1271 (N_1271,N_587,N_727);
nand U1272 (N_1272,N_958,N_572);
and U1273 (N_1273,N_776,N_579);
nand U1274 (N_1274,N_861,N_766);
nand U1275 (N_1275,N_804,N_556);
and U1276 (N_1276,N_914,N_655);
nand U1277 (N_1277,N_721,N_588);
nor U1278 (N_1278,N_842,N_517);
and U1279 (N_1279,N_557,N_871);
or U1280 (N_1280,N_891,N_748);
and U1281 (N_1281,N_947,N_993);
nor U1282 (N_1282,N_869,N_602);
xnor U1283 (N_1283,N_987,N_515);
or U1284 (N_1284,N_731,N_542);
and U1285 (N_1285,N_897,N_637);
nor U1286 (N_1286,N_696,N_753);
nand U1287 (N_1287,N_784,N_563);
nor U1288 (N_1288,N_791,N_722);
nor U1289 (N_1289,N_971,N_634);
nand U1290 (N_1290,N_520,N_646);
and U1291 (N_1291,N_743,N_785);
nor U1292 (N_1292,N_749,N_623);
or U1293 (N_1293,N_556,N_634);
xor U1294 (N_1294,N_804,N_577);
nand U1295 (N_1295,N_777,N_763);
nor U1296 (N_1296,N_740,N_774);
and U1297 (N_1297,N_744,N_774);
nand U1298 (N_1298,N_986,N_595);
and U1299 (N_1299,N_709,N_952);
and U1300 (N_1300,N_978,N_530);
and U1301 (N_1301,N_580,N_996);
nor U1302 (N_1302,N_537,N_659);
nand U1303 (N_1303,N_661,N_678);
or U1304 (N_1304,N_939,N_636);
and U1305 (N_1305,N_898,N_512);
and U1306 (N_1306,N_775,N_657);
or U1307 (N_1307,N_555,N_669);
nor U1308 (N_1308,N_608,N_676);
and U1309 (N_1309,N_636,N_811);
nor U1310 (N_1310,N_960,N_870);
nand U1311 (N_1311,N_705,N_908);
and U1312 (N_1312,N_548,N_616);
xnor U1313 (N_1313,N_909,N_842);
nor U1314 (N_1314,N_776,N_721);
nor U1315 (N_1315,N_662,N_576);
nor U1316 (N_1316,N_974,N_890);
nor U1317 (N_1317,N_623,N_755);
nor U1318 (N_1318,N_537,N_775);
nand U1319 (N_1319,N_652,N_638);
and U1320 (N_1320,N_581,N_647);
xnor U1321 (N_1321,N_631,N_743);
nor U1322 (N_1322,N_613,N_937);
nor U1323 (N_1323,N_648,N_984);
and U1324 (N_1324,N_927,N_574);
or U1325 (N_1325,N_666,N_929);
or U1326 (N_1326,N_933,N_883);
and U1327 (N_1327,N_745,N_821);
xnor U1328 (N_1328,N_856,N_516);
or U1329 (N_1329,N_567,N_963);
nand U1330 (N_1330,N_667,N_506);
nand U1331 (N_1331,N_769,N_795);
or U1332 (N_1332,N_560,N_553);
nand U1333 (N_1333,N_565,N_632);
nand U1334 (N_1334,N_540,N_897);
nor U1335 (N_1335,N_841,N_705);
and U1336 (N_1336,N_793,N_511);
nand U1337 (N_1337,N_947,N_583);
nand U1338 (N_1338,N_854,N_570);
nand U1339 (N_1339,N_971,N_763);
or U1340 (N_1340,N_787,N_672);
nand U1341 (N_1341,N_845,N_833);
nor U1342 (N_1342,N_899,N_576);
nor U1343 (N_1343,N_928,N_960);
nand U1344 (N_1344,N_583,N_966);
and U1345 (N_1345,N_709,N_956);
or U1346 (N_1346,N_711,N_731);
nor U1347 (N_1347,N_533,N_591);
and U1348 (N_1348,N_934,N_870);
nor U1349 (N_1349,N_606,N_553);
nor U1350 (N_1350,N_710,N_788);
nand U1351 (N_1351,N_720,N_648);
nor U1352 (N_1352,N_512,N_674);
nor U1353 (N_1353,N_704,N_596);
nor U1354 (N_1354,N_861,N_922);
or U1355 (N_1355,N_509,N_511);
or U1356 (N_1356,N_681,N_658);
or U1357 (N_1357,N_555,N_914);
nor U1358 (N_1358,N_574,N_520);
nand U1359 (N_1359,N_620,N_741);
and U1360 (N_1360,N_535,N_581);
nor U1361 (N_1361,N_837,N_900);
nor U1362 (N_1362,N_551,N_552);
nor U1363 (N_1363,N_726,N_941);
nand U1364 (N_1364,N_965,N_532);
nor U1365 (N_1365,N_757,N_602);
nand U1366 (N_1366,N_975,N_935);
and U1367 (N_1367,N_656,N_549);
nand U1368 (N_1368,N_653,N_590);
nor U1369 (N_1369,N_873,N_553);
nand U1370 (N_1370,N_817,N_814);
or U1371 (N_1371,N_815,N_975);
or U1372 (N_1372,N_816,N_815);
nor U1373 (N_1373,N_968,N_597);
and U1374 (N_1374,N_619,N_834);
xnor U1375 (N_1375,N_783,N_985);
or U1376 (N_1376,N_978,N_677);
or U1377 (N_1377,N_938,N_678);
and U1378 (N_1378,N_761,N_852);
nor U1379 (N_1379,N_713,N_719);
or U1380 (N_1380,N_700,N_573);
nor U1381 (N_1381,N_542,N_605);
xnor U1382 (N_1382,N_870,N_982);
nor U1383 (N_1383,N_948,N_905);
or U1384 (N_1384,N_675,N_647);
and U1385 (N_1385,N_522,N_612);
and U1386 (N_1386,N_533,N_578);
nor U1387 (N_1387,N_894,N_626);
and U1388 (N_1388,N_914,N_523);
and U1389 (N_1389,N_865,N_520);
and U1390 (N_1390,N_731,N_746);
nor U1391 (N_1391,N_632,N_605);
and U1392 (N_1392,N_502,N_798);
nor U1393 (N_1393,N_515,N_848);
nand U1394 (N_1394,N_824,N_705);
nand U1395 (N_1395,N_870,N_811);
nand U1396 (N_1396,N_841,N_925);
and U1397 (N_1397,N_929,N_886);
nor U1398 (N_1398,N_505,N_566);
nand U1399 (N_1399,N_612,N_682);
and U1400 (N_1400,N_696,N_706);
or U1401 (N_1401,N_774,N_844);
nor U1402 (N_1402,N_603,N_559);
nand U1403 (N_1403,N_870,N_635);
or U1404 (N_1404,N_754,N_833);
nor U1405 (N_1405,N_785,N_798);
nand U1406 (N_1406,N_800,N_633);
xor U1407 (N_1407,N_509,N_695);
nor U1408 (N_1408,N_867,N_915);
xnor U1409 (N_1409,N_669,N_736);
nor U1410 (N_1410,N_742,N_574);
and U1411 (N_1411,N_870,N_890);
nor U1412 (N_1412,N_518,N_680);
or U1413 (N_1413,N_930,N_985);
or U1414 (N_1414,N_999,N_703);
nand U1415 (N_1415,N_809,N_981);
nor U1416 (N_1416,N_500,N_706);
and U1417 (N_1417,N_783,N_697);
nand U1418 (N_1418,N_912,N_968);
or U1419 (N_1419,N_977,N_969);
nor U1420 (N_1420,N_939,N_907);
nand U1421 (N_1421,N_659,N_615);
or U1422 (N_1422,N_672,N_743);
nor U1423 (N_1423,N_570,N_648);
nor U1424 (N_1424,N_897,N_676);
or U1425 (N_1425,N_920,N_765);
nor U1426 (N_1426,N_808,N_880);
or U1427 (N_1427,N_997,N_699);
and U1428 (N_1428,N_920,N_557);
or U1429 (N_1429,N_777,N_805);
nand U1430 (N_1430,N_759,N_880);
nand U1431 (N_1431,N_543,N_546);
nand U1432 (N_1432,N_530,N_735);
nand U1433 (N_1433,N_704,N_609);
nor U1434 (N_1434,N_557,N_878);
and U1435 (N_1435,N_922,N_907);
nand U1436 (N_1436,N_642,N_660);
nor U1437 (N_1437,N_820,N_999);
xnor U1438 (N_1438,N_580,N_556);
or U1439 (N_1439,N_878,N_933);
and U1440 (N_1440,N_865,N_991);
and U1441 (N_1441,N_600,N_986);
nor U1442 (N_1442,N_891,N_602);
and U1443 (N_1443,N_712,N_585);
nand U1444 (N_1444,N_779,N_715);
and U1445 (N_1445,N_640,N_637);
or U1446 (N_1446,N_760,N_792);
or U1447 (N_1447,N_919,N_531);
nand U1448 (N_1448,N_744,N_902);
nand U1449 (N_1449,N_971,N_935);
and U1450 (N_1450,N_540,N_818);
nor U1451 (N_1451,N_615,N_606);
and U1452 (N_1452,N_953,N_800);
nand U1453 (N_1453,N_839,N_836);
or U1454 (N_1454,N_761,N_939);
nand U1455 (N_1455,N_982,N_672);
or U1456 (N_1456,N_983,N_670);
nand U1457 (N_1457,N_577,N_844);
nand U1458 (N_1458,N_870,N_797);
nor U1459 (N_1459,N_665,N_910);
and U1460 (N_1460,N_595,N_614);
or U1461 (N_1461,N_878,N_823);
or U1462 (N_1462,N_833,N_589);
or U1463 (N_1463,N_939,N_536);
nand U1464 (N_1464,N_882,N_602);
and U1465 (N_1465,N_658,N_831);
and U1466 (N_1466,N_603,N_707);
nand U1467 (N_1467,N_966,N_730);
or U1468 (N_1468,N_845,N_770);
nor U1469 (N_1469,N_874,N_843);
nor U1470 (N_1470,N_674,N_763);
nand U1471 (N_1471,N_858,N_998);
nor U1472 (N_1472,N_873,N_930);
nand U1473 (N_1473,N_911,N_742);
and U1474 (N_1474,N_901,N_896);
nand U1475 (N_1475,N_667,N_886);
nor U1476 (N_1476,N_877,N_638);
and U1477 (N_1477,N_999,N_581);
or U1478 (N_1478,N_985,N_758);
xnor U1479 (N_1479,N_735,N_896);
nand U1480 (N_1480,N_502,N_615);
and U1481 (N_1481,N_739,N_960);
and U1482 (N_1482,N_969,N_908);
xnor U1483 (N_1483,N_818,N_983);
and U1484 (N_1484,N_503,N_852);
and U1485 (N_1485,N_740,N_901);
nand U1486 (N_1486,N_556,N_864);
nand U1487 (N_1487,N_970,N_595);
and U1488 (N_1488,N_753,N_736);
nand U1489 (N_1489,N_614,N_733);
or U1490 (N_1490,N_824,N_802);
and U1491 (N_1491,N_819,N_667);
or U1492 (N_1492,N_701,N_616);
nand U1493 (N_1493,N_943,N_935);
nor U1494 (N_1494,N_718,N_687);
and U1495 (N_1495,N_894,N_959);
or U1496 (N_1496,N_609,N_832);
nand U1497 (N_1497,N_902,N_934);
nor U1498 (N_1498,N_766,N_768);
or U1499 (N_1499,N_762,N_670);
xor U1500 (N_1500,N_1105,N_1322);
nor U1501 (N_1501,N_1005,N_1064);
and U1502 (N_1502,N_1439,N_1112);
nor U1503 (N_1503,N_1458,N_1072);
nor U1504 (N_1504,N_1130,N_1109);
or U1505 (N_1505,N_1317,N_1283);
or U1506 (N_1506,N_1304,N_1110);
xor U1507 (N_1507,N_1205,N_1416);
nand U1508 (N_1508,N_1312,N_1356);
or U1509 (N_1509,N_1122,N_1261);
xnor U1510 (N_1510,N_1101,N_1329);
and U1511 (N_1511,N_1021,N_1031);
and U1512 (N_1512,N_1196,N_1246);
nand U1513 (N_1513,N_1438,N_1314);
and U1514 (N_1514,N_1455,N_1431);
nor U1515 (N_1515,N_1429,N_1425);
or U1516 (N_1516,N_1282,N_1121);
and U1517 (N_1517,N_1010,N_1019);
nand U1518 (N_1518,N_1147,N_1288);
nand U1519 (N_1519,N_1287,N_1223);
nor U1520 (N_1520,N_1332,N_1368);
nor U1521 (N_1521,N_1488,N_1046);
and U1522 (N_1522,N_1178,N_1417);
nand U1523 (N_1523,N_1289,N_1389);
nand U1524 (N_1524,N_1373,N_1259);
and U1525 (N_1525,N_1040,N_1348);
nand U1526 (N_1526,N_1263,N_1254);
and U1527 (N_1527,N_1024,N_1371);
xor U1528 (N_1528,N_1074,N_1483);
nor U1529 (N_1529,N_1187,N_1100);
nor U1530 (N_1530,N_1142,N_1041);
or U1531 (N_1531,N_1065,N_1071);
or U1532 (N_1532,N_1229,N_1159);
nor U1533 (N_1533,N_1061,N_1042);
nor U1534 (N_1534,N_1292,N_1001);
nand U1535 (N_1535,N_1244,N_1009);
nor U1536 (N_1536,N_1491,N_1272);
nor U1537 (N_1537,N_1043,N_1111);
and U1538 (N_1538,N_1301,N_1191);
nor U1539 (N_1539,N_1423,N_1481);
and U1540 (N_1540,N_1123,N_1233);
and U1541 (N_1541,N_1498,N_1459);
nand U1542 (N_1542,N_1426,N_1214);
or U1543 (N_1543,N_1236,N_1091);
and U1544 (N_1544,N_1250,N_1392);
or U1545 (N_1545,N_1231,N_1474);
nand U1546 (N_1546,N_1321,N_1369);
xor U1547 (N_1547,N_1313,N_1144);
or U1548 (N_1548,N_1410,N_1281);
nand U1549 (N_1549,N_1385,N_1028);
nand U1550 (N_1550,N_1052,N_1357);
nand U1551 (N_1551,N_1038,N_1255);
and U1552 (N_1552,N_1405,N_1493);
and U1553 (N_1553,N_1413,N_1396);
nand U1554 (N_1554,N_1190,N_1402);
nor U1555 (N_1555,N_1175,N_1445);
or U1556 (N_1556,N_1352,N_1027);
nand U1557 (N_1557,N_1343,N_1427);
and U1558 (N_1558,N_1486,N_1390);
nor U1559 (N_1559,N_1117,N_1443);
and U1560 (N_1560,N_1238,N_1218);
xnor U1561 (N_1561,N_1471,N_1157);
and U1562 (N_1562,N_1472,N_1068);
nor U1563 (N_1563,N_1376,N_1387);
or U1564 (N_1564,N_1129,N_1036);
or U1565 (N_1565,N_1222,N_1085);
nor U1566 (N_1566,N_1268,N_1184);
nand U1567 (N_1567,N_1464,N_1497);
and U1568 (N_1568,N_1059,N_1465);
nand U1569 (N_1569,N_1119,N_1367);
nor U1570 (N_1570,N_1437,N_1219);
nor U1571 (N_1571,N_1393,N_1362);
or U1572 (N_1572,N_1020,N_1099);
nor U1573 (N_1573,N_1490,N_1168);
or U1574 (N_1574,N_1243,N_1118);
or U1575 (N_1575,N_1169,N_1489);
nand U1576 (N_1576,N_1424,N_1325);
nor U1577 (N_1577,N_1299,N_1284);
nor U1578 (N_1578,N_1311,N_1355);
or U1579 (N_1579,N_1492,N_1276);
nand U1580 (N_1580,N_1225,N_1409);
nor U1581 (N_1581,N_1240,N_1432);
or U1582 (N_1582,N_1015,N_1192);
and U1583 (N_1583,N_1251,N_1440);
or U1584 (N_1584,N_1349,N_1460);
and U1585 (N_1585,N_1278,N_1346);
xor U1586 (N_1586,N_1477,N_1073);
nand U1587 (N_1587,N_1331,N_1418);
and U1588 (N_1588,N_1476,N_1485);
nor U1589 (N_1589,N_1442,N_1145);
or U1590 (N_1590,N_1307,N_1083);
nand U1591 (N_1591,N_1297,N_1163);
nand U1592 (N_1592,N_1473,N_1138);
and U1593 (N_1593,N_1401,N_1300);
nand U1594 (N_1594,N_1048,N_1279);
and U1595 (N_1595,N_1080,N_1003);
nor U1596 (N_1596,N_1245,N_1228);
nor U1597 (N_1597,N_1412,N_1058);
nor U1598 (N_1598,N_1347,N_1204);
and U1599 (N_1599,N_1155,N_1088);
and U1600 (N_1600,N_1221,N_1333);
and U1601 (N_1601,N_1057,N_1198);
or U1602 (N_1602,N_1395,N_1170);
xor U1603 (N_1603,N_1203,N_1388);
and U1604 (N_1604,N_1306,N_1496);
nor U1605 (N_1605,N_1081,N_1149);
nand U1606 (N_1606,N_1360,N_1450);
nand U1607 (N_1607,N_1340,N_1107);
and U1608 (N_1608,N_1146,N_1158);
or U1609 (N_1609,N_1454,N_1139);
nor U1610 (N_1610,N_1098,N_1078);
nand U1611 (N_1611,N_1293,N_1125);
nand U1612 (N_1612,N_1495,N_1186);
and U1613 (N_1613,N_1089,N_1013);
or U1614 (N_1614,N_1411,N_1093);
nor U1615 (N_1615,N_1366,N_1232);
nand U1616 (N_1616,N_1258,N_1039);
or U1617 (N_1617,N_1239,N_1398);
or U1618 (N_1618,N_1188,N_1051);
or U1619 (N_1619,N_1358,N_1176);
and U1620 (N_1620,N_1422,N_1103);
or U1621 (N_1621,N_1270,N_1049);
and U1622 (N_1622,N_1004,N_1453);
or U1623 (N_1623,N_1044,N_1115);
nand U1624 (N_1624,N_1160,N_1179);
nor U1625 (N_1625,N_1319,N_1202);
nand U1626 (N_1626,N_1226,N_1235);
nand U1627 (N_1627,N_1032,N_1494);
and U1628 (N_1628,N_1183,N_1165);
and U1629 (N_1629,N_1137,N_1253);
and U1630 (N_1630,N_1060,N_1308);
nand U1631 (N_1631,N_1391,N_1189);
and U1632 (N_1632,N_1377,N_1249);
nor U1633 (N_1633,N_1014,N_1095);
or U1634 (N_1634,N_1403,N_1127);
and U1635 (N_1635,N_1126,N_1256);
nand U1636 (N_1636,N_1215,N_1033);
and U1637 (N_1637,N_1242,N_1153);
nand U1638 (N_1638,N_1108,N_1007);
nand U1639 (N_1639,N_1327,N_1234);
and U1640 (N_1640,N_1478,N_1482);
and U1641 (N_1641,N_1378,N_1008);
nor U1642 (N_1642,N_1267,N_1208);
nor U1643 (N_1643,N_1150,N_1034);
and U1644 (N_1644,N_1269,N_1151);
xnor U1645 (N_1645,N_1381,N_1141);
and U1646 (N_1646,N_1404,N_1456);
nand U1647 (N_1647,N_1419,N_1448);
xor U1648 (N_1648,N_1323,N_1156);
xor U1649 (N_1649,N_1320,N_1280);
or U1650 (N_1650,N_1140,N_1173);
nor U1651 (N_1651,N_1045,N_1029);
and U1652 (N_1652,N_1247,N_1285);
nor U1653 (N_1653,N_1361,N_1104);
nor U1654 (N_1654,N_1075,N_1069);
xnor U1655 (N_1655,N_1182,N_1224);
nor U1656 (N_1656,N_1309,N_1067);
and U1657 (N_1657,N_1161,N_1000);
and U1658 (N_1658,N_1096,N_1180);
nand U1659 (N_1659,N_1116,N_1386);
nor U1660 (N_1660,N_1076,N_1216);
nand U1661 (N_1661,N_1408,N_1206);
and U1662 (N_1662,N_1446,N_1047);
or U1663 (N_1663,N_1197,N_1016);
and U1664 (N_1664,N_1185,N_1466);
and U1665 (N_1665,N_1181,N_1394);
or U1666 (N_1666,N_1382,N_1266);
and U1667 (N_1667,N_1209,N_1022);
nand U1668 (N_1668,N_1164,N_1484);
nor U1669 (N_1669,N_1342,N_1444);
or U1670 (N_1670,N_1227,N_1274);
or U1671 (N_1671,N_1248,N_1436);
nor U1672 (N_1672,N_1400,N_1054);
or U1673 (N_1673,N_1406,N_1372);
nand U1674 (N_1674,N_1262,N_1207);
and U1675 (N_1675,N_1026,N_1449);
nor U1676 (N_1676,N_1066,N_1201);
and U1677 (N_1677,N_1050,N_1345);
nand U1678 (N_1678,N_1296,N_1193);
nor U1679 (N_1679,N_1002,N_1037);
or U1680 (N_1680,N_1452,N_1177);
or U1681 (N_1681,N_1467,N_1303);
or U1682 (N_1682,N_1433,N_1035);
nand U1683 (N_1683,N_1328,N_1434);
nand U1684 (N_1684,N_1351,N_1220);
and U1685 (N_1685,N_1023,N_1017);
nand U1686 (N_1686,N_1171,N_1124);
and U1687 (N_1687,N_1344,N_1135);
nor U1688 (N_1688,N_1338,N_1375);
nand U1689 (N_1689,N_1154,N_1336);
nand U1690 (N_1690,N_1326,N_1475);
and U1691 (N_1691,N_1379,N_1430);
or U1692 (N_1692,N_1363,N_1011);
or U1693 (N_1693,N_1148,N_1428);
nand U1694 (N_1694,N_1469,N_1102);
or U1695 (N_1695,N_1370,N_1077);
nand U1696 (N_1696,N_1480,N_1133);
and U1697 (N_1697,N_1241,N_1166);
or U1698 (N_1698,N_1252,N_1260);
and U1699 (N_1699,N_1337,N_1479);
nor U1700 (N_1700,N_1062,N_1174);
or U1701 (N_1701,N_1053,N_1120);
and U1702 (N_1702,N_1499,N_1167);
nand U1703 (N_1703,N_1082,N_1414);
nor U1704 (N_1704,N_1315,N_1063);
or U1705 (N_1705,N_1086,N_1025);
nand U1706 (N_1706,N_1273,N_1237);
xnor U1707 (N_1707,N_1441,N_1397);
nand U1708 (N_1708,N_1462,N_1407);
or U1709 (N_1709,N_1055,N_1463);
nand U1710 (N_1710,N_1350,N_1341);
and U1711 (N_1711,N_1200,N_1114);
or U1712 (N_1712,N_1470,N_1374);
xnor U1713 (N_1713,N_1018,N_1457);
or U1714 (N_1714,N_1195,N_1291);
or U1715 (N_1715,N_1217,N_1305);
nand U1716 (N_1716,N_1415,N_1084);
nor U1717 (N_1717,N_1451,N_1132);
nand U1718 (N_1718,N_1334,N_1364);
and U1719 (N_1719,N_1230,N_1079);
or U1720 (N_1720,N_1090,N_1210);
nand U1721 (N_1721,N_1318,N_1257);
nand U1722 (N_1722,N_1468,N_1435);
nor U1723 (N_1723,N_1113,N_1136);
nand U1724 (N_1724,N_1295,N_1383);
nor U1725 (N_1725,N_1030,N_1290);
and U1726 (N_1726,N_1172,N_1012);
nand U1727 (N_1727,N_1087,N_1365);
and U1728 (N_1728,N_1212,N_1152);
nor U1729 (N_1729,N_1399,N_1265);
nand U1730 (N_1730,N_1194,N_1006);
nand U1731 (N_1731,N_1353,N_1339);
nand U1732 (N_1732,N_1277,N_1094);
nand U1733 (N_1733,N_1092,N_1447);
nand U1734 (N_1734,N_1134,N_1264);
nor U1735 (N_1735,N_1384,N_1302);
or U1736 (N_1736,N_1421,N_1106);
nor U1737 (N_1737,N_1097,N_1310);
nor U1738 (N_1738,N_1275,N_1271);
nor U1739 (N_1739,N_1354,N_1286);
nand U1740 (N_1740,N_1461,N_1298);
nand U1741 (N_1741,N_1131,N_1316);
nor U1742 (N_1742,N_1330,N_1324);
nand U1743 (N_1743,N_1143,N_1213);
nor U1744 (N_1744,N_1294,N_1199);
or U1745 (N_1745,N_1211,N_1487);
and U1746 (N_1746,N_1380,N_1070);
nor U1747 (N_1747,N_1056,N_1162);
and U1748 (N_1748,N_1420,N_1335);
or U1749 (N_1749,N_1128,N_1359);
nand U1750 (N_1750,N_1386,N_1166);
nor U1751 (N_1751,N_1189,N_1135);
nor U1752 (N_1752,N_1151,N_1465);
or U1753 (N_1753,N_1230,N_1479);
and U1754 (N_1754,N_1327,N_1095);
nand U1755 (N_1755,N_1332,N_1187);
nand U1756 (N_1756,N_1215,N_1031);
and U1757 (N_1757,N_1401,N_1222);
and U1758 (N_1758,N_1373,N_1334);
or U1759 (N_1759,N_1103,N_1409);
and U1760 (N_1760,N_1458,N_1078);
or U1761 (N_1761,N_1334,N_1031);
or U1762 (N_1762,N_1316,N_1475);
or U1763 (N_1763,N_1071,N_1055);
nor U1764 (N_1764,N_1421,N_1408);
nor U1765 (N_1765,N_1036,N_1390);
or U1766 (N_1766,N_1071,N_1388);
nand U1767 (N_1767,N_1471,N_1242);
nor U1768 (N_1768,N_1415,N_1035);
nand U1769 (N_1769,N_1371,N_1288);
and U1770 (N_1770,N_1399,N_1382);
xnor U1771 (N_1771,N_1204,N_1097);
and U1772 (N_1772,N_1412,N_1086);
nand U1773 (N_1773,N_1145,N_1315);
or U1774 (N_1774,N_1251,N_1050);
nor U1775 (N_1775,N_1409,N_1052);
nor U1776 (N_1776,N_1489,N_1325);
nor U1777 (N_1777,N_1108,N_1015);
and U1778 (N_1778,N_1303,N_1211);
nand U1779 (N_1779,N_1438,N_1059);
nand U1780 (N_1780,N_1429,N_1317);
nor U1781 (N_1781,N_1266,N_1195);
and U1782 (N_1782,N_1120,N_1405);
nor U1783 (N_1783,N_1161,N_1450);
and U1784 (N_1784,N_1082,N_1295);
or U1785 (N_1785,N_1105,N_1320);
or U1786 (N_1786,N_1330,N_1137);
nor U1787 (N_1787,N_1015,N_1163);
and U1788 (N_1788,N_1397,N_1255);
or U1789 (N_1789,N_1192,N_1016);
and U1790 (N_1790,N_1438,N_1136);
and U1791 (N_1791,N_1030,N_1024);
nor U1792 (N_1792,N_1404,N_1061);
or U1793 (N_1793,N_1482,N_1260);
or U1794 (N_1794,N_1473,N_1380);
or U1795 (N_1795,N_1356,N_1184);
nand U1796 (N_1796,N_1171,N_1399);
or U1797 (N_1797,N_1321,N_1462);
nand U1798 (N_1798,N_1257,N_1142);
or U1799 (N_1799,N_1163,N_1056);
nor U1800 (N_1800,N_1275,N_1320);
or U1801 (N_1801,N_1462,N_1143);
nand U1802 (N_1802,N_1317,N_1350);
nor U1803 (N_1803,N_1415,N_1349);
and U1804 (N_1804,N_1062,N_1465);
or U1805 (N_1805,N_1005,N_1398);
or U1806 (N_1806,N_1433,N_1251);
nand U1807 (N_1807,N_1370,N_1204);
nor U1808 (N_1808,N_1289,N_1121);
nor U1809 (N_1809,N_1454,N_1153);
and U1810 (N_1810,N_1265,N_1424);
and U1811 (N_1811,N_1437,N_1063);
xnor U1812 (N_1812,N_1423,N_1004);
or U1813 (N_1813,N_1399,N_1434);
nand U1814 (N_1814,N_1034,N_1430);
and U1815 (N_1815,N_1206,N_1100);
nor U1816 (N_1816,N_1038,N_1235);
nand U1817 (N_1817,N_1106,N_1157);
nor U1818 (N_1818,N_1013,N_1051);
nand U1819 (N_1819,N_1121,N_1342);
nor U1820 (N_1820,N_1411,N_1011);
nand U1821 (N_1821,N_1243,N_1117);
nor U1822 (N_1822,N_1387,N_1378);
or U1823 (N_1823,N_1495,N_1358);
xnor U1824 (N_1824,N_1078,N_1393);
nor U1825 (N_1825,N_1481,N_1098);
or U1826 (N_1826,N_1357,N_1365);
xor U1827 (N_1827,N_1337,N_1197);
and U1828 (N_1828,N_1157,N_1456);
nand U1829 (N_1829,N_1344,N_1427);
nand U1830 (N_1830,N_1401,N_1034);
or U1831 (N_1831,N_1295,N_1412);
nand U1832 (N_1832,N_1182,N_1418);
and U1833 (N_1833,N_1478,N_1423);
or U1834 (N_1834,N_1166,N_1419);
nand U1835 (N_1835,N_1181,N_1436);
nor U1836 (N_1836,N_1076,N_1209);
or U1837 (N_1837,N_1376,N_1054);
nor U1838 (N_1838,N_1371,N_1139);
nand U1839 (N_1839,N_1323,N_1146);
nand U1840 (N_1840,N_1059,N_1436);
nand U1841 (N_1841,N_1438,N_1371);
and U1842 (N_1842,N_1484,N_1231);
nand U1843 (N_1843,N_1199,N_1214);
nor U1844 (N_1844,N_1083,N_1458);
or U1845 (N_1845,N_1209,N_1152);
and U1846 (N_1846,N_1081,N_1436);
nor U1847 (N_1847,N_1000,N_1274);
nor U1848 (N_1848,N_1121,N_1062);
nor U1849 (N_1849,N_1160,N_1093);
and U1850 (N_1850,N_1014,N_1417);
nand U1851 (N_1851,N_1331,N_1373);
xnor U1852 (N_1852,N_1287,N_1389);
nand U1853 (N_1853,N_1462,N_1302);
xor U1854 (N_1854,N_1198,N_1035);
nand U1855 (N_1855,N_1190,N_1492);
nor U1856 (N_1856,N_1233,N_1105);
and U1857 (N_1857,N_1204,N_1402);
nand U1858 (N_1858,N_1234,N_1433);
and U1859 (N_1859,N_1190,N_1439);
nor U1860 (N_1860,N_1296,N_1073);
nand U1861 (N_1861,N_1227,N_1327);
nor U1862 (N_1862,N_1236,N_1127);
nor U1863 (N_1863,N_1021,N_1033);
and U1864 (N_1864,N_1228,N_1042);
or U1865 (N_1865,N_1216,N_1045);
or U1866 (N_1866,N_1432,N_1462);
nand U1867 (N_1867,N_1072,N_1480);
and U1868 (N_1868,N_1044,N_1224);
and U1869 (N_1869,N_1470,N_1069);
nand U1870 (N_1870,N_1288,N_1481);
or U1871 (N_1871,N_1354,N_1275);
and U1872 (N_1872,N_1443,N_1046);
nor U1873 (N_1873,N_1398,N_1012);
or U1874 (N_1874,N_1358,N_1344);
nor U1875 (N_1875,N_1483,N_1055);
and U1876 (N_1876,N_1094,N_1187);
xnor U1877 (N_1877,N_1495,N_1315);
nor U1878 (N_1878,N_1425,N_1325);
nand U1879 (N_1879,N_1167,N_1133);
and U1880 (N_1880,N_1355,N_1493);
or U1881 (N_1881,N_1165,N_1001);
and U1882 (N_1882,N_1184,N_1171);
or U1883 (N_1883,N_1109,N_1281);
and U1884 (N_1884,N_1113,N_1448);
nand U1885 (N_1885,N_1098,N_1321);
nor U1886 (N_1886,N_1133,N_1062);
nand U1887 (N_1887,N_1212,N_1258);
nor U1888 (N_1888,N_1038,N_1179);
nor U1889 (N_1889,N_1159,N_1174);
and U1890 (N_1890,N_1471,N_1255);
and U1891 (N_1891,N_1270,N_1017);
nor U1892 (N_1892,N_1167,N_1321);
nand U1893 (N_1893,N_1324,N_1412);
xnor U1894 (N_1894,N_1153,N_1037);
nand U1895 (N_1895,N_1300,N_1239);
or U1896 (N_1896,N_1291,N_1496);
nand U1897 (N_1897,N_1311,N_1380);
or U1898 (N_1898,N_1299,N_1033);
and U1899 (N_1899,N_1146,N_1047);
nor U1900 (N_1900,N_1135,N_1470);
xnor U1901 (N_1901,N_1075,N_1483);
or U1902 (N_1902,N_1255,N_1291);
or U1903 (N_1903,N_1235,N_1451);
nor U1904 (N_1904,N_1265,N_1296);
or U1905 (N_1905,N_1056,N_1083);
and U1906 (N_1906,N_1258,N_1256);
nand U1907 (N_1907,N_1061,N_1262);
or U1908 (N_1908,N_1093,N_1255);
or U1909 (N_1909,N_1239,N_1169);
nand U1910 (N_1910,N_1411,N_1499);
nor U1911 (N_1911,N_1410,N_1284);
or U1912 (N_1912,N_1447,N_1091);
nor U1913 (N_1913,N_1287,N_1447);
and U1914 (N_1914,N_1120,N_1372);
nor U1915 (N_1915,N_1232,N_1310);
and U1916 (N_1916,N_1457,N_1117);
nor U1917 (N_1917,N_1473,N_1123);
and U1918 (N_1918,N_1053,N_1415);
or U1919 (N_1919,N_1244,N_1356);
nor U1920 (N_1920,N_1113,N_1056);
nand U1921 (N_1921,N_1272,N_1411);
and U1922 (N_1922,N_1192,N_1499);
nor U1923 (N_1923,N_1024,N_1008);
and U1924 (N_1924,N_1211,N_1271);
nand U1925 (N_1925,N_1483,N_1239);
and U1926 (N_1926,N_1242,N_1199);
and U1927 (N_1927,N_1022,N_1173);
or U1928 (N_1928,N_1339,N_1458);
nand U1929 (N_1929,N_1104,N_1054);
and U1930 (N_1930,N_1207,N_1213);
or U1931 (N_1931,N_1358,N_1250);
nor U1932 (N_1932,N_1091,N_1469);
or U1933 (N_1933,N_1350,N_1213);
and U1934 (N_1934,N_1346,N_1283);
nor U1935 (N_1935,N_1275,N_1223);
or U1936 (N_1936,N_1343,N_1384);
nand U1937 (N_1937,N_1279,N_1114);
nand U1938 (N_1938,N_1036,N_1464);
nand U1939 (N_1939,N_1259,N_1186);
and U1940 (N_1940,N_1403,N_1044);
nor U1941 (N_1941,N_1164,N_1255);
or U1942 (N_1942,N_1346,N_1153);
nor U1943 (N_1943,N_1312,N_1405);
nor U1944 (N_1944,N_1393,N_1295);
and U1945 (N_1945,N_1360,N_1228);
nand U1946 (N_1946,N_1022,N_1189);
or U1947 (N_1947,N_1041,N_1382);
or U1948 (N_1948,N_1172,N_1031);
nor U1949 (N_1949,N_1078,N_1485);
and U1950 (N_1950,N_1160,N_1327);
and U1951 (N_1951,N_1296,N_1330);
and U1952 (N_1952,N_1226,N_1110);
nand U1953 (N_1953,N_1159,N_1233);
nand U1954 (N_1954,N_1135,N_1207);
and U1955 (N_1955,N_1307,N_1124);
nor U1956 (N_1956,N_1376,N_1488);
or U1957 (N_1957,N_1390,N_1161);
and U1958 (N_1958,N_1356,N_1268);
nand U1959 (N_1959,N_1317,N_1144);
nand U1960 (N_1960,N_1366,N_1022);
and U1961 (N_1961,N_1196,N_1375);
nand U1962 (N_1962,N_1023,N_1315);
nand U1963 (N_1963,N_1375,N_1496);
nor U1964 (N_1964,N_1096,N_1421);
nor U1965 (N_1965,N_1019,N_1383);
and U1966 (N_1966,N_1387,N_1496);
and U1967 (N_1967,N_1481,N_1278);
nor U1968 (N_1968,N_1093,N_1343);
or U1969 (N_1969,N_1086,N_1315);
nand U1970 (N_1970,N_1172,N_1315);
or U1971 (N_1971,N_1315,N_1472);
nor U1972 (N_1972,N_1272,N_1075);
nor U1973 (N_1973,N_1196,N_1305);
or U1974 (N_1974,N_1219,N_1184);
or U1975 (N_1975,N_1340,N_1344);
or U1976 (N_1976,N_1081,N_1048);
or U1977 (N_1977,N_1458,N_1423);
and U1978 (N_1978,N_1257,N_1475);
xor U1979 (N_1979,N_1183,N_1231);
and U1980 (N_1980,N_1229,N_1189);
or U1981 (N_1981,N_1410,N_1419);
or U1982 (N_1982,N_1362,N_1306);
or U1983 (N_1983,N_1246,N_1295);
or U1984 (N_1984,N_1480,N_1046);
nor U1985 (N_1985,N_1184,N_1406);
nand U1986 (N_1986,N_1450,N_1149);
nor U1987 (N_1987,N_1075,N_1277);
nand U1988 (N_1988,N_1411,N_1169);
nor U1989 (N_1989,N_1372,N_1416);
nand U1990 (N_1990,N_1064,N_1307);
or U1991 (N_1991,N_1464,N_1139);
nor U1992 (N_1992,N_1060,N_1113);
nor U1993 (N_1993,N_1197,N_1376);
nand U1994 (N_1994,N_1106,N_1215);
nand U1995 (N_1995,N_1260,N_1429);
nand U1996 (N_1996,N_1257,N_1457);
or U1997 (N_1997,N_1389,N_1034);
and U1998 (N_1998,N_1039,N_1450);
and U1999 (N_1999,N_1354,N_1366);
xnor U2000 (N_2000,N_1827,N_1610);
nor U2001 (N_2001,N_1686,N_1917);
and U2002 (N_2002,N_1582,N_1990);
and U2003 (N_2003,N_1746,N_1898);
or U2004 (N_2004,N_1574,N_1517);
nand U2005 (N_2005,N_1885,N_1659);
and U2006 (N_2006,N_1835,N_1942);
or U2007 (N_2007,N_1542,N_1941);
nor U2008 (N_2008,N_1645,N_1638);
nor U2009 (N_2009,N_1628,N_1794);
nor U2010 (N_2010,N_1979,N_1796);
nor U2011 (N_2011,N_1823,N_1683);
and U2012 (N_2012,N_1616,N_1673);
nor U2013 (N_2013,N_1602,N_1579);
or U2014 (N_2014,N_1671,N_1844);
and U2015 (N_2015,N_1732,N_1553);
nand U2016 (N_2016,N_1782,N_1750);
and U2017 (N_2017,N_1825,N_1536);
or U2018 (N_2018,N_1731,N_1666);
or U2019 (N_2019,N_1648,N_1967);
nand U2020 (N_2020,N_1787,N_1716);
or U2021 (N_2021,N_1888,N_1846);
or U2022 (N_2022,N_1678,N_1832);
nor U2023 (N_2023,N_1996,N_1593);
nand U2024 (N_2024,N_1961,N_1710);
or U2025 (N_2025,N_1854,N_1758);
nand U2026 (N_2026,N_1535,N_1781);
nor U2027 (N_2027,N_1540,N_1926);
and U2028 (N_2028,N_1580,N_1989);
and U2029 (N_2029,N_1864,N_1798);
nand U2030 (N_2030,N_1664,N_1637);
nand U2031 (N_2031,N_1919,N_1913);
xnor U2032 (N_2032,N_1760,N_1887);
and U2033 (N_2033,N_1713,N_1661);
and U2034 (N_2034,N_1721,N_1784);
nand U2035 (N_2035,N_1631,N_1501);
xor U2036 (N_2036,N_1998,N_1868);
and U2037 (N_2037,N_1959,N_1972);
nand U2038 (N_2038,N_1896,N_1875);
and U2039 (N_2039,N_1783,N_1807);
nor U2040 (N_2040,N_1764,N_1903);
nor U2041 (N_2041,N_1838,N_1573);
nand U2042 (N_2042,N_1692,N_1563);
nor U2043 (N_2043,N_1995,N_1656);
xnor U2044 (N_2044,N_1867,N_1655);
or U2045 (N_2045,N_1589,N_1911);
nand U2046 (N_2046,N_1761,N_1733);
nor U2047 (N_2047,N_1667,N_1634);
xnor U2048 (N_2048,N_1943,N_1650);
nand U2049 (N_2049,N_1584,N_1891);
nor U2050 (N_2050,N_1675,N_1663);
nand U2051 (N_2051,N_1946,N_1636);
or U2052 (N_2052,N_1630,N_1785);
xnor U2053 (N_2053,N_1882,N_1518);
or U2054 (N_2054,N_1546,N_1551);
and U2055 (N_2055,N_1811,N_1618);
nor U2056 (N_2056,N_1775,N_1510);
and U2057 (N_2057,N_1830,N_1519);
nand U2058 (N_2058,N_1842,N_1806);
and U2059 (N_2059,N_1873,N_1822);
nor U2060 (N_2060,N_1951,N_1590);
nand U2061 (N_2061,N_1607,N_1994);
nor U2062 (N_2062,N_1984,N_1562);
and U2063 (N_2063,N_1642,N_1841);
xnor U2064 (N_2064,N_1687,N_1568);
or U2065 (N_2065,N_1978,N_1670);
nand U2066 (N_2066,N_1737,N_1526);
nor U2067 (N_2067,N_1970,N_1725);
and U2068 (N_2068,N_1500,N_1576);
or U2069 (N_2069,N_1833,N_1528);
nand U2070 (N_2070,N_1522,N_1914);
nand U2071 (N_2071,N_1587,N_1985);
nor U2072 (N_2072,N_1677,N_1708);
xor U2073 (N_2073,N_1759,N_1803);
and U2074 (N_2074,N_1726,N_1707);
nand U2075 (N_2075,N_1814,N_1554);
nor U2076 (N_2076,N_1639,N_1925);
or U2077 (N_2077,N_1955,N_1578);
and U2078 (N_2078,N_1701,N_1815);
nand U2079 (N_2079,N_1818,N_1819);
and U2080 (N_2080,N_1795,N_1641);
or U2081 (N_2081,N_1693,N_1715);
and U2082 (N_2082,N_1852,N_1559);
or U2083 (N_2083,N_1921,N_1586);
nand U2084 (N_2084,N_1859,N_1709);
nor U2085 (N_2085,N_1702,N_1679);
and U2086 (N_2086,N_1876,N_1899);
nand U2087 (N_2087,N_1747,N_1699);
nand U2088 (N_2088,N_1769,N_1626);
nand U2089 (N_2089,N_1717,N_1912);
and U2090 (N_2090,N_1541,N_1694);
nand U2091 (N_2091,N_1991,N_1968);
nor U2092 (N_2092,N_1558,N_1892);
nor U2093 (N_2093,N_1848,N_1965);
and U2094 (N_2094,N_1521,N_1604);
nor U2095 (N_2095,N_1722,N_1539);
or U2096 (N_2096,N_1765,N_1964);
and U2097 (N_2097,N_1625,N_1640);
or U2098 (N_2098,N_1997,N_1860);
and U2099 (N_2099,N_1880,N_1533);
nand U2100 (N_2100,N_1662,N_1776);
nand U2101 (N_2101,N_1564,N_1691);
and U2102 (N_2102,N_1895,N_1986);
or U2103 (N_2103,N_1740,N_1719);
or U2104 (N_2104,N_1947,N_1894);
or U2105 (N_2105,N_1729,N_1936);
nand U2106 (N_2106,N_1767,N_1527);
or U2107 (N_2107,N_1883,N_1665);
nor U2108 (N_2108,N_1723,N_1752);
nand U2109 (N_2109,N_1930,N_1613);
nand U2110 (N_2110,N_1742,N_1870);
and U2111 (N_2111,N_1847,N_1504);
and U2112 (N_2112,N_1976,N_1952);
and U2113 (N_2113,N_1572,N_1538);
nand U2114 (N_2114,N_1697,N_1547);
nor U2115 (N_2115,N_1931,N_1674);
or U2116 (N_2116,N_1916,N_1700);
nand U2117 (N_2117,N_1906,N_1884);
nand U2118 (N_2118,N_1856,N_1608);
nor U2119 (N_2119,N_1975,N_1766);
nor U2120 (N_2120,N_1513,N_1754);
nor U2121 (N_2121,N_1817,N_1609);
nand U2122 (N_2122,N_1770,N_1657);
and U2123 (N_2123,N_1757,N_1736);
nand U2124 (N_2124,N_1591,N_1577);
and U2125 (N_2125,N_1804,N_1744);
nor U2126 (N_2126,N_1548,N_1935);
nor U2127 (N_2127,N_1704,N_1845);
and U2128 (N_2128,N_1508,N_1531);
and U2129 (N_2129,N_1646,N_1890);
and U2130 (N_2130,N_1515,N_1592);
or U2131 (N_2131,N_1843,N_1774);
and U2132 (N_2132,N_1872,N_1617);
nand U2133 (N_2133,N_1809,N_1960);
nand U2134 (N_2134,N_1571,N_1810);
nand U2135 (N_2135,N_1599,N_1566);
xnor U2136 (N_2136,N_1824,N_1669);
and U2137 (N_2137,N_1944,N_1505);
nor U2138 (N_2138,N_1971,N_1922);
nand U2139 (N_2139,N_1581,N_1793);
nor U2140 (N_2140,N_1749,N_1762);
nor U2141 (N_2141,N_1556,N_1711);
nand U2142 (N_2142,N_1881,N_1605);
or U2143 (N_2143,N_1988,N_1603);
nor U2144 (N_2144,N_1956,N_1768);
nor U2145 (N_2145,N_1569,N_1612);
nand U2146 (N_2146,N_1857,N_1954);
nand U2147 (N_2147,N_1871,N_1739);
or U2148 (N_2148,N_1950,N_1743);
nand U2149 (N_2149,N_1816,N_1753);
nor U2150 (N_2150,N_1866,N_1712);
nor U2151 (N_2151,N_1703,N_1649);
nand U2152 (N_2152,N_1973,N_1685);
nor U2153 (N_2153,N_1619,N_1530);
and U2154 (N_2154,N_1738,N_1920);
nor U2155 (N_2155,N_1836,N_1902);
nand U2156 (N_2156,N_1779,N_1643);
xor U2157 (N_2157,N_1982,N_1858);
xor U2158 (N_2158,N_1909,N_1654);
or U2159 (N_2159,N_1908,N_1727);
nand U2160 (N_2160,N_1869,N_1735);
and U2161 (N_2161,N_1834,N_1681);
xor U2162 (N_2162,N_1658,N_1745);
nor U2163 (N_2163,N_1840,N_1940);
nor U2164 (N_2164,N_1969,N_1651);
and U2165 (N_2165,N_1755,N_1910);
or U2166 (N_2166,N_1821,N_1791);
or U2167 (N_2167,N_1934,N_1588);
nand U2168 (N_2168,N_1855,N_1839);
nand U2169 (N_2169,N_1644,N_1748);
or U2170 (N_2170,N_1583,N_1615);
nand U2171 (N_2171,N_1682,N_1861);
or U2172 (N_2172,N_1544,N_1698);
or U2173 (N_2173,N_1904,N_1596);
or U2174 (N_2174,N_1585,N_1621);
nor U2175 (N_2175,N_1983,N_1620);
and U2176 (N_2176,N_1557,N_1632);
xor U2177 (N_2177,N_1614,N_1751);
and U2178 (N_2178,N_1532,N_1647);
nor U2179 (N_2179,N_1777,N_1907);
nand U2180 (N_2180,N_1805,N_1741);
nand U2181 (N_2181,N_1652,N_1966);
and U2182 (N_2182,N_1993,N_1690);
nor U2183 (N_2183,N_1594,N_1831);
nand U2184 (N_2184,N_1812,N_1676);
xnor U2185 (N_2185,N_1850,N_1958);
nand U2186 (N_2186,N_1992,N_1889);
nor U2187 (N_2187,N_1980,N_1520);
nor U2188 (N_2188,N_1606,N_1549);
and U2189 (N_2189,N_1624,N_1865);
and U2190 (N_2190,N_1598,N_1780);
and U2191 (N_2191,N_1627,N_1689);
nor U2192 (N_2192,N_1863,N_1826);
nor U2193 (N_2193,N_1957,N_1706);
and U2194 (N_2194,N_1837,N_1684);
and U2195 (N_2195,N_1789,N_1511);
or U2196 (N_2196,N_1977,N_1820);
and U2197 (N_2197,N_1509,N_1962);
and U2198 (N_2198,N_1561,N_1567);
nand U2199 (N_2199,N_1808,N_1945);
or U2200 (N_2200,N_1849,N_1877);
or U2201 (N_2201,N_1611,N_1705);
and U2202 (N_2202,N_1575,N_1622);
or U2203 (N_2203,N_1905,N_1529);
or U2204 (N_2204,N_1555,N_1653);
nor U2205 (N_2205,N_1786,N_1773);
xnor U2206 (N_2206,N_1688,N_1525);
and U2207 (N_2207,N_1801,N_1829);
nand U2208 (N_2208,N_1623,N_1695);
xor U2209 (N_2209,N_1629,N_1503);
nor U2210 (N_2210,N_1734,N_1999);
nor U2211 (N_2211,N_1918,N_1728);
nor U2212 (N_2212,N_1799,N_1927);
and U2213 (N_2213,N_1595,N_1720);
nor U2214 (N_2214,N_1928,N_1696);
nand U2215 (N_2215,N_1502,N_1797);
or U2216 (N_2216,N_1552,N_1974);
and U2217 (N_2217,N_1948,N_1937);
nand U2218 (N_2218,N_1813,N_1828);
or U2219 (N_2219,N_1963,N_1788);
and U2220 (N_2220,N_1771,N_1512);
nor U2221 (N_2221,N_1893,N_1724);
nand U2222 (N_2222,N_1874,N_1900);
or U2223 (N_2223,N_1514,N_1802);
nand U2224 (N_2224,N_1672,N_1901);
nand U2225 (N_2225,N_1534,N_1790);
nor U2226 (N_2226,N_1800,N_1600);
nand U2227 (N_2227,N_1792,N_1853);
or U2228 (N_2228,N_1680,N_1516);
and U2229 (N_2229,N_1714,N_1862);
xor U2230 (N_2230,N_1886,N_1543);
or U2231 (N_2231,N_1523,N_1550);
nor U2232 (N_2232,N_1597,N_1851);
nor U2233 (N_2233,N_1537,N_1633);
nand U2234 (N_2234,N_1915,N_1524);
nor U2235 (N_2235,N_1763,N_1635);
or U2236 (N_2236,N_1506,N_1560);
or U2237 (N_2237,N_1929,N_1601);
or U2238 (N_2238,N_1730,N_1938);
nor U2239 (N_2239,N_1756,N_1897);
and U2240 (N_2240,N_1924,N_1570);
nor U2241 (N_2241,N_1981,N_1933);
nand U2242 (N_2242,N_1772,N_1668);
nor U2243 (N_2243,N_1718,N_1987);
nor U2244 (N_2244,N_1923,N_1660);
and U2245 (N_2245,N_1545,N_1932);
nor U2246 (N_2246,N_1879,N_1953);
or U2247 (N_2247,N_1565,N_1878);
or U2248 (N_2248,N_1939,N_1507);
or U2249 (N_2249,N_1949,N_1778);
nor U2250 (N_2250,N_1628,N_1687);
or U2251 (N_2251,N_1884,N_1868);
nand U2252 (N_2252,N_1994,N_1888);
nor U2253 (N_2253,N_1668,N_1832);
and U2254 (N_2254,N_1620,N_1994);
and U2255 (N_2255,N_1557,N_1838);
nand U2256 (N_2256,N_1597,N_1617);
and U2257 (N_2257,N_1576,N_1931);
xnor U2258 (N_2258,N_1596,N_1921);
or U2259 (N_2259,N_1753,N_1959);
or U2260 (N_2260,N_1833,N_1639);
or U2261 (N_2261,N_1682,N_1928);
nor U2262 (N_2262,N_1913,N_1544);
and U2263 (N_2263,N_1965,N_1782);
nand U2264 (N_2264,N_1502,N_1801);
nand U2265 (N_2265,N_1866,N_1872);
nand U2266 (N_2266,N_1682,N_1997);
nand U2267 (N_2267,N_1710,N_1934);
nand U2268 (N_2268,N_1667,N_1763);
or U2269 (N_2269,N_1769,N_1515);
nand U2270 (N_2270,N_1668,N_1606);
nor U2271 (N_2271,N_1723,N_1946);
nor U2272 (N_2272,N_1800,N_1607);
nand U2273 (N_2273,N_1722,N_1678);
nor U2274 (N_2274,N_1729,N_1863);
nor U2275 (N_2275,N_1939,N_1658);
and U2276 (N_2276,N_1532,N_1994);
nand U2277 (N_2277,N_1591,N_1909);
and U2278 (N_2278,N_1530,N_1820);
nor U2279 (N_2279,N_1637,N_1778);
nor U2280 (N_2280,N_1914,N_1989);
and U2281 (N_2281,N_1612,N_1554);
and U2282 (N_2282,N_1777,N_1945);
and U2283 (N_2283,N_1559,N_1888);
and U2284 (N_2284,N_1872,N_1602);
or U2285 (N_2285,N_1512,N_1838);
or U2286 (N_2286,N_1619,N_1734);
nor U2287 (N_2287,N_1852,N_1504);
xor U2288 (N_2288,N_1585,N_1830);
or U2289 (N_2289,N_1566,N_1812);
nor U2290 (N_2290,N_1985,N_1504);
and U2291 (N_2291,N_1857,N_1830);
nand U2292 (N_2292,N_1865,N_1906);
or U2293 (N_2293,N_1588,N_1543);
nand U2294 (N_2294,N_1503,N_1979);
or U2295 (N_2295,N_1665,N_1661);
or U2296 (N_2296,N_1589,N_1525);
nor U2297 (N_2297,N_1634,N_1576);
nand U2298 (N_2298,N_1743,N_1772);
or U2299 (N_2299,N_1694,N_1964);
nor U2300 (N_2300,N_1539,N_1720);
nand U2301 (N_2301,N_1787,N_1686);
or U2302 (N_2302,N_1556,N_1509);
and U2303 (N_2303,N_1977,N_1863);
nor U2304 (N_2304,N_1569,N_1766);
nor U2305 (N_2305,N_1871,N_1623);
and U2306 (N_2306,N_1553,N_1876);
or U2307 (N_2307,N_1745,N_1637);
and U2308 (N_2308,N_1553,N_1520);
nand U2309 (N_2309,N_1852,N_1985);
nor U2310 (N_2310,N_1903,N_1804);
or U2311 (N_2311,N_1702,N_1937);
and U2312 (N_2312,N_1609,N_1845);
nand U2313 (N_2313,N_1892,N_1691);
or U2314 (N_2314,N_1588,N_1798);
nand U2315 (N_2315,N_1782,N_1920);
and U2316 (N_2316,N_1823,N_1725);
and U2317 (N_2317,N_1527,N_1646);
or U2318 (N_2318,N_1730,N_1744);
and U2319 (N_2319,N_1633,N_1538);
nand U2320 (N_2320,N_1844,N_1862);
and U2321 (N_2321,N_1727,N_1802);
and U2322 (N_2322,N_1992,N_1854);
nor U2323 (N_2323,N_1805,N_1814);
or U2324 (N_2324,N_1550,N_1657);
nand U2325 (N_2325,N_1950,N_1988);
or U2326 (N_2326,N_1888,N_1663);
or U2327 (N_2327,N_1747,N_1512);
or U2328 (N_2328,N_1536,N_1601);
and U2329 (N_2329,N_1914,N_1715);
nor U2330 (N_2330,N_1995,N_1677);
and U2331 (N_2331,N_1869,N_1922);
and U2332 (N_2332,N_1928,N_1827);
nor U2333 (N_2333,N_1905,N_1721);
and U2334 (N_2334,N_1820,N_1660);
and U2335 (N_2335,N_1741,N_1597);
and U2336 (N_2336,N_1602,N_1994);
nor U2337 (N_2337,N_1958,N_1809);
or U2338 (N_2338,N_1959,N_1983);
nand U2339 (N_2339,N_1914,N_1661);
nor U2340 (N_2340,N_1982,N_1632);
and U2341 (N_2341,N_1724,N_1512);
xnor U2342 (N_2342,N_1966,N_1779);
and U2343 (N_2343,N_1814,N_1859);
nand U2344 (N_2344,N_1522,N_1695);
and U2345 (N_2345,N_1768,N_1647);
and U2346 (N_2346,N_1562,N_1771);
nor U2347 (N_2347,N_1757,N_1737);
or U2348 (N_2348,N_1890,N_1815);
xnor U2349 (N_2349,N_1923,N_1826);
nand U2350 (N_2350,N_1651,N_1959);
xor U2351 (N_2351,N_1598,N_1663);
and U2352 (N_2352,N_1863,N_1883);
xnor U2353 (N_2353,N_1644,N_1917);
nor U2354 (N_2354,N_1972,N_1799);
or U2355 (N_2355,N_1902,N_1803);
and U2356 (N_2356,N_1676,N_1523);
or U2357 (N_2357,N_1933,N_1923);
or U2358 (N_2358,N_1850,N_1503);
nor U2359 (N_2359,N_1641,N_1605);
nand U2360 (N_2360,N_1993,N_1767);
and U2361 (N_2361,N_1524,N_1589);
and U2362 (N_2362,N_1723,N_1603);
and U2363 (N_2363,N_1554,N_1611);
or U2364 (N_2364,N_1959,N_1535);
xor U2365 (N_2365,N_1553,N_1919);
nor U2366 (N_2366,N_1614,N_1814);
nand U2367 (N_2367,N_1890,N_1569);
and U2368 (N_2368,N_1826,N_1594);
and U2369 (N_2369,N_1685,N_1787);
nor U2370 (N_2370,N_1883,N_1951);
or U2371 (N_2371,N_1745,N_1654);
or U2372 (N_2372,N_1723,N_1806);
nor U2373 (N_2373,N_1904,N_1949);
nor U2374 (N_2374,N_1555,N_1854);
nor U2375 (N_2375,N_1716,N_1696);
nor U2376 (N_2376,N_1648,N_1819);
or U2377 (N_2377,N_1908,N_1538);
or U2378 (N_2378,N_1751,N_1683);
nand U2379 (N_2379,N_1664,N_1567);
nor U2380 (N_2380,N_1792,N_1885);
or U2381 (N_2381,N_1775,N_1590);
nand U2382 (N_2382,N_1935,N_1639);
and U2383 (N_2383,N_1770,N_1794);
nand U2384 (N_2384,N_1684,N_1672);
or U2385 (N_2385,N_1818,N_1766);
and U2386 (N_2386,N_1890,N_1797);
nor U2387 (N_2387,N_1505,N_1856);
nor U2388 (N_2388,N_1561,N_1972);
nand U2389 (N_2389,N_1846,N_1617);
or U2390 (N_2390,N_1775,N_1914);
nand U2391 (N_2391,N_1796,N_1923);
and U2392 (N_2392,N_1512,N_1998);
or U2393 (N_2393,N_1624,N_1787);
and U2394 (N_2394,N_1838,N_1931);
nand U2395 (N_2395,N_1934,N_1754);
nor U2396 (N_2396,N_1722,N_1985);
or U2397 (N_2397,N_1850,N_1518);
nor U2398 (N_2398,N_1994,N_1549);
and U2399 (N_2399,N_1878,N_1843);
or U2400 (N_2400,N_1789,N_1843);
or U2401 (N_2401,N_1671,N_1579);
nand U2402 (N_2402,N_1802,N_1531);
or U2403 (N_2403,N_1679,N_1878);
or U2404 (N_2404,N_1917,N_1624);
or U2405 (N_2405,N_1597,N_1747);
nand U2406 (N_2406,N_1578,N_1825);
nor U2407 (N_2407,N_1505,N_1681);
nor U2408 (N_2408,N_1686,N_1557);
nor U2409 (N_2409,N_1705,N_1736);
nor U2410 (N_2410,N_1760,N_1720);
nand U2411 (N_2411,N_1810,N_1695);
and U2412 (N_2412,N_1587,N_1794);
nor U2413 (N_2413,N_1638,N_1776);
or U2414 (N_2414,N_1888,N_1734);
or U2415 (N_2415,N_1517,N_1973);
or U2416 (N_2416,N_1818,N_1823);
nor U2417 (N_2417,N_1843,N_1665);
nand U2418 (N_2418,N_1962,N_1627);
and U2419 (N_2419,N_1862,N_1650);
and U2420 (N_2420,N_1538,N_1776);
nand U2421 (N_2421,N_1888,N_1664);
or U2422 (N_2422,N_1954,N_1965);
and U2423 (N_2423,N_1955,N_1808);
or U2424 (N_2424,N_1652,N_1585);
or U2425 (N_2425,N_1996,N_1901);
or U2426 (N_2426,N_1524,N_1611);
xnor U2427 (N_2427,N_1804,N_1912);
nor U2428 (N_2428,N_1550,N_1933);
or U2429 (N_2429,N_1800,N_1655);
xnor U2430 (N_2430,N_1911,N_1728);
nor U2431 (N_2431,N_1660,N_1727);
or U2432 (N_2432,N_1711,N_1843);
nand U2433 (N_2433,N_1534,N_1825);
or U2434 (N_2434,N_1905,N_1758);
nor U2435 (N_2435,N_1980,N_1726);
nor U2436 (N_2436,N_1864,N_1707);
nor U2437 (N_2437,N_1809,N_1989);
and U2438 (N_2438,N_1885,N_1993);
nor U2439 (N_2439,N_1835,N_1707);
nor U2440 (N_2440,N_1801,N_1748);
and U2441 (N_2441,N_1946,N_1533);
nor U2442 (N_2442,N_1601,N_1856);
nor U2443 (N_2443,N_1574,N_1748);
or U2444 (N_2444,N_1507,N_1544);
nor U2445 (N_2445,N_1546,N_1544);
nand U2446 (N_2446,N_1634,N_1784);
nor U2447 (N_2447,N_1921,N_1655);
or U2448 (N_2448,N_1767,N_1637);
and U2449 (N_2449,N_1530,N_1566);
or U2450 (N_2450,N_1576,N_1821);
and U2451 (N_2451,N_1538,N_1506);
or U2452 (N_2452,N_1930,N_1707);
nor U2453 (N_2453,N_1919,N_1691);
and U2454 (N_2454,N_1724,N_1706);
nand U2455 (N_2455,N_1849,N_1622);
and U2456 (N_2456,N_1906,N_1752);
and U2457 (N_2457,N_1633,N_1923);
or U2458 (N_2458,N_1865,N_1680);
and U2459 (N_2459,N_1593,N_1622);
and U2460 (N_2460,N_1577,N_1568);
nor U2461 (N_2461,N_1890,N_1945);
xnor U2462 (N_2462,N_1866,N_1543);
nand U2463 (N_2463,N_1524,N_1810);
or U2464 (N_2464,N_1993,N_1521);
nand U2465 (N_2465,N_1513,N_1745);
nand U2466 (N_2466,N_1536,N_1986);
or U2467 (N_2467,N_1857,N_1925);
nand U2468 (N_2468,N_1622,N_1650);
nand U2469 (N_2469,N_1715,N_1849);
xor U2470 (N_2470,N_1647,N_1751);
or U2471 (N_2471,N_1600,N_1531);
and U2472 (N_2472,N_1872,N_1962);
nand U2473 (N_2473,N_1629,N_1807);
or U2474 (N_2474,N_1690,N_1525);
and U2475 (N_2475,N_1937,N_1979);
and U2476 (N_2476,N_1785,N_1933);
and U2477 (N_2477,N_1692,N_1695);
nand U2478 (N_2478,N_1920,N_1686);
or U2479 (N_2479,N_1552,N_1619);
or U2480 (N_2480,N_1568,N_1725);
or U2481 (N_2481,N_1607,N_1575);
nand U2482 (N_2482,N_1741,N_1664);
or U2483 (N_2483,N_1591,N_1977);
nor U2484 (N_2484,N_1506,N_1642);
and U2485 (N_2485,N_1784,N_1951);
or U2486 (N_2486,N_1675,N_1961);
or U2487 (N_2487,N_1672,N_1728);
nor U2488 (N_2488,N_1693,N_1961);
or U2489 (N_2489,N_1551,N_1504);
or U2490 (N_2490,N_1904,N_1953);
nand U2491 (N_2491,N_1915,N_1549);
and U2492 (N_2492,N_1929,N_1666);
and U2493 (N_2493,N_1930,N_1777);
and U2494 (N_2494,N_1842,N_1544);
or U2495 (N_2495,N_1851,N_1739);
nor U2496 (N_2496,N_1876,N_1817);
and U2497 (N_2497,N_1539,N_1956);
nor U2498 (N_2498,N_1667,N_1508);
or U2499 (N_2499,N_1844,N_1841);
nand U2500 (N_2500,N_2418,N_2212);
nand U2501 (N_2501,N_2216,N_2182);
nor U2502 (N_2502,N_2225,N_2483);
nand U2503 (N_2503,N_2438,N_2346);
nand U2504 (N_2504,N_2058,N_2349);
nor U2505 (N_2505,N_2037,N_2307);
nor U2506 (N_2506,N_2296,N_2211);
nor U2507 (N_2507,N_2300,N_2371);
or U2508 (N_2508,N_2080,N_2039);
nand U2509 (N_2509,N_2098,N_2056);
and U2510 (N_2510,N_2199,N_2284);
nor U2511 (N_2511,N_2028,N_2352);
nor U2512 (N_2512,N_2153,N_2087);
nor U2513 (N_2513,N_2413,N_2150);
nand U2514 (N_2514,N_2137,N_2391);
and U2515 (N_2515,N_2126,N_2492);
nand U2516 (N_2516,N_2267,N_2079);
nor U2517 (N_2517,N_2077,N_2240);
nand U2518 (N_2518,N_2421,N_2074);
xnor U2519 (N_2519,N_2390,N_2471);
nor U2520 (N_2520,N_2232,N_2345);
nor U2521 (N_2521,N_2067,N_2168);
xor U2522 (N_2522,N_2209,N_2289);
or U2523 (N_2523,N_2254,N_2044);
or U2524 (N_2524,N_2218,N_2249);
nor U2525 (N_2525,N_2172,N_2157);
nand U2526 (N_2526,N_2226,N_2432);
and U2527 (N_2527,N_2151,N_2487);
or U2528 (N_2528,N_2395,N_2445);
nor U2529 (N_2529,N_2140,N_2177);
or U2530 (N_2530,N_2207,N_2295);
nand U2531 (N_2531,N_2021,N_2447);
or U2532 (N_2532,N_2308,N_2405);
nor U2533 (N_2533,N_2241,N_2129);
or U2534 (N_2534,N_2132,N_2486);
nor U2535 (N_2535,N_2115,N_2061);
nand U2536 (N_2536,N_2223,N_2313);
nand U2537 (N_2537,N_2312,N_2416);
nand U2538 (N_2538,N_2449,N_2222);
and U2539 (N_2539,N_2347,N_2382);
nor U2540 (N_2540,N_2431,N_2377);
nand U2541 (N_2541,N_2474,N_2165);
nand U2542 (N_2542,N_2263,N_2496);
and U2543 (N_2543,N_2442,N_2237);
or U2544 (N_2544,N_2453,N_2446);
nand U2545 (N_2545,N_2135,N_2023);
and U2546 (N_2546,N_2299,N_2310);
nor U2547 (N_2547,N_2428,N_2429);
nor U2548 (N_2548,N_2214,N_2489);
and U2549 (N_2549,N_2354,N_2494);
nand U2550 (N_2550,N_2201,N_2411);
or U2551 (N_2551,N_2005,N_2319);
nand U2552 (N_2552,N_2478,N_2049);
nand U2553 (N_2553,N_2130,N_2235);
nor U2554 (N_2554,N_2440,N_2205);
or U2555 (N_2555,N_2069,N_2465);
xor U2556 (N_2556,N_2099,N_2188);
or U2557 (N_2557,N_2381,N_2460);
nand U2558 (N_2558,N_2253,N_2053);
nand U2559 (N_2559,N_2359,N_2191);
nor U2560 (N_2560,N_2084,N_2327);
nor U2561 (N_2561,N_2458,N_2063);
nand U2562 (N_2562,N_2055,N_2376);
nand U2563 (N_2563,N_2092,N_2259);
and U2564 (N_2564,N_2178,N_2015);
nand U2565 (N_2565,N_2244,N_2324);
nand U2566 (N_2566,N_2000,N_2043);
nand U2567 (N_2567,N_2139,N_2422);
nor U2568 (N_2568,N_2481,N_2258);
or U2569 (N_2569,N_2409,N_2325);
or U2570 (N_2570,N_2384,N_2329);
and U2571 (N_2571,N_2113,N_2336);
nor U2572 (N_2572,N_2142,N_2022);
and U2573 (N_2573,N_2260,N_2499);
and U2574 (N_2574,N_2148,N_2497);
nor U2575 (N_2575,N_2001,N_2356);
nand U2576 (N_2576,N_2170,N_2275);
nand U2577 (N_2577,N_2255,N_2357);
and U2578 (N_2578,N_2062,N_2366);
nor U2579 (N_2579,N_2025,N_2332);
nand U2580 (N_2580,N_2206,N_2468);
or U2581 (N_2581,N_2368,N_2270);
and U2582 (N_2582,N_2152,N_2108);
and U2583 (N_2583,N_2027,N_2333);
nand U2584 (N_2584,N_2339,N_2475);
nor U2585 (N_2585,N_2125,N_2195);
and U2586 (N_2586,N_2387,N_2197);
xnor U2587 (N_2587,N_2190,N_2102);
and U2588 (N_2588,N_2277,N_2109);
nand U2589 (N_2589,N_2407,N_2479);
and U2590 (N_2590,N_2457,N_2330);
and U2591 (N_2591,N_2451,N_2236);
nand U2592 (N_2592,N_2276,N_2250);
and U2593 (N_2593,N_2193,N_2246);
nor U2594 (N_2594,N_2101,N_2004);
nand U2595 (N_2595,N_2105,N_2184);
or U2596 (N_2596,N_2408,N_2385);
and U2597 (N_2597,N_2302,N_2012);
or U2598 (N_2598,N_2454,N_2426);
and U2599 (N_2599,N_2133,N_2213);
nor U2600 (N_2600,N_2287,N_2118);
nand U2601 (N_2601,N_2396,N_2059);
and U2602 (N_2602,N_2323,N_2116);
and U2603 (N_2603,N_2233,N_2161);
or U2604 (N_2604,N_2141,N_2427);
nand U2605 (N_2605,N_2181,N_2176);
nand U2606 (N_2606,N_2169,N_2401);
and U2607 (N_2607,N_2495,N_2078);
nand U2608 (N_2608,N_2219,N_2341);
and U2609 (N_2609,N_2159,N_2180);
xnor U2610 (N_2610,N_2171,N_2488);
xor U2611 (N_2611,N_2154,N_2064);
or U2612 (N_2612,N_2072,N_2472);
or U2613 (N_2613,N_2412,N_2298);
nand U2614 (N_2614,N_2361,N_2315);
nand U2615 (N_2615,N_2014,N_2322);
nand U2616 (N_2616,N_2038,N_2490);
and U2617 (N_2617,N_2045,N_2110);
or U2618 (N_2618,N_2173,N_2117);
and U2619 (N_2619,N_2456,N_2441);
nor U2620 (N_2620,N_2245,N_2477);
xor U2621 (N_2621,N_2283,N_2402);
nor U2622 (N_2622,N_2434,N_2484);
nor U2623 (N_2623,N_2268,N_2466);
xor U2624 (N_2624,N_2394,N_2318);
or U2625 (N_2625,N_2397,N_2210);
or U2626 (N_2626,N_2485,N_2155);
nor U2627 (N_2627,N_2128,N_2208);
nand U2628 (N_2628,N_2452,N_2301);
or U2629 (N_2629,N_2389,N_2363);
nand U2630 (N_2630,N_2399,N_2158);
nor U2631 (N_2631,N_2034,N_2417);
or U2632 (N_2632,N_2439,N_2370);
and U2633 (N_2633,N_2493,N_2247);
nand U2634 (N_2634,N_2229,N_2328);
nand U2635 (N_2635,N_2362,N_2279);
or U2636 (N_2636,N_2112,N_2095);
and U2637 (N_2637,N_2261,N_2054);
nor U2638 (N_2638,N_2175,N_2424);
nand U2639 (N_2639,N_2187,N_2273);
and U2640 (N_2640,N_2076,N_2234);
nand U2641 (N_2641,N_2430,N_2437);
or U2642 (N_2642,N_2463,N_2192);
and U2643 (N_2643,N_2119,N_2075);
nor U2644 (N_2644,N_2353,N_2406);
nor U2645 (N_2645,N_2285,N_2278);
nor U2646 (N_2646,N_2435,N_2462);
or U2647 (N_2647,N_2337,N_2280);
nor U2648 (N_2648,N_2017,N_2138);
or U2649 (N_2649,N_2290,N_2364);
nor U2650 (N_2650,N_2414,N_2344);
and U2651 (N_2651,N_2160,N_2060);
and U2652 (N_2652,N_2145,N_2403);
or U2653 (N_2653,N_2008,N_2068);
or U2654 (N_2654,N_2262,N_2048);
and U2655 (N_2655,N_2269,N_2470);
or U2656 (N_2656,N_2179,N_2392);
nand U2657 (N_2657,N_2450,N_2291);
and U2658 (N_2658,N_2018,N_2448);
or U2659 (N_2659,N_2030,N_2114);
nand U2660 (N_2660,N_2163,N_2200);
nor U2661 (N_2661,N_2097,N_2010);
or U2662 (N_2662,N_2026,N_2265);
nor U2663 (N_2663,N_2239,N_2041);
nor U2664 (N_2664,N_2007,N_2002);
xnor U2665 (N_2665,N_2257,N_2057);
or U2666 (N_2666,N_2309,N_2013);
nand U2667 (N_2667,N_2100,N_2256);
nand U2668 (N_2668,N_2033,N_2029);
and U2669 (N_2669,N_2081,N_2185);
or U2670 (N_2670,N_2380,N_2016);
nor U2671 (N_2671,N_2374,N_2147);
or U2672 (N_2672,N_2198,N_2303);
nor U2673 (N_2673,N_2335,N_2167);
nor U2674 (N_2674,N_2360,N_2351);
xor U2675 (N_2675,N_2051,N_2252);
nand U2676 (N_2676,N_2024,N_2317);
and U2677 (N_2677,N_2086,N_2204);
and U2678 (N_2678,N_2415,N_2123);
nand U2679 (N_2679,N_2433,N_2386);
and U2680 (N_2680,N_2294,N_2202);
nor U2681 (N_2681,N_2293,N_2047);
or U2682 (N_2682,N_2003,N_2009);
nor U2683 (N_2683,N_2383,N_2476);
nor U2684 (N_2684,N_2071,N_2243);
nor U2685 (N_2685,N_2443,N_2127);
and U2686 (N_2686,N_2404,N_2073);
or U2687 (N_2687,N_2050,N_2297);
and U2688 (N_2688,N_2350,N_2019);
nor U2689 (N_2689,N_2122,N_2321);
and U2690 (N_2690,N_2091,N_2085);
or U2691 (N_2691,N_2316,N_2420);
nand U2692 (N_2692,N_2436,N_2036);
and U2693 (N_2693,N_2032,N_2183);
and U2694 (N_2694,N_2035,N_2134);
nand U2695 (N_2695,N_2146,N_2372);
and U2696 (N_2696,N_2094,N_2046);
nor U2697 (N_2697,N_2228,N_2189);
nand U2698 (N_2698,N_2286,N_2461);
and U2699 (N_2699,N_2238,N_2083);
or U2700 (N_2700,N_2455,N_2375);
nor U2701 (N_2701,N_2281,N_2338);
or U2702 (N_2702,N_2220,N_2480);
nand U2703 (N_2703,N_2367,N_2162);
nor U2704 (N_2704,N_2111,N_2006);
and U2705 (N_2705,N_2031,N_2136);
nand U2706 (N_2706,N_2215,N_2304);
and U2707 (N_2707,N_2469,N_2444);
nor U2708 (N_2708,N_2231,N_2340);
nor U2709 (N_2709,N_2288,N_2311);
nor U2710 (N_2710,N_2410,N_2348);
and U2711 (N_2711,N_2326,N_2282);
or U2712 (N_2712,N_2082,N_2143);
nor U2713 (N_2713,N_2274,N_2089);
and U2714 (N_2714,N_2272,N_2149);
and U2715 (N_2715,N_2164,N_2106);
nor U2716 (N_2716,N_2242,N_2388);
nor U2717 (N_2717,N_2482,N_2196);
nand U2718 (N_2718,N_2186,N_2203);
nand U2719 (N_2719,N_2369,N_2096);
and U2720 (N_2720,N_2491,N_2042);
and U2721 (N_2721,N_2464,N_2227);
or U2722 (N_2722,N_2090,N_2121);
or U2723 (N_2723,N_2378,N_2107);
and U2724 (N_2724,N_2156,N_2305);
nor U2725 (N_2725,N_2314,N_2251);
or U2726 (N_2726,N_2358,N_2343);
xor U2727 (N_2727,N_2070,N_2419);
and U2728 (N_2728,N_2365,N_2355);
and U2729 (N_2729,N_2271,N_2459);
nor U2730 (N_2730,N_2103,N_2124);
nand U2731 (N_2731,N_2373,N_2342);
or U2732 (N_2732,N_2264,N_2292);
nand U2733 (N_2733,N_2066,N_2248);
or U2734 (N_2734,N_2467,N_2425);
and U2735 (N_2735,N_2104,N_2320);
or U2736 (N_2736,N_2306,N_2334);
and U2737 (N_2737,N_2088,N_2144);
xnor U2738 (N_2738,N_2040,N_2052);
nor U2739 (N_2739,N_2498,N_2120);
nor U2740 (N_2740,N_2065,N_2221);
xor U2741 (N_2741,N_2174,N_2224);
nor U2742 (N_2742,N_2266,N_2423);
and U2743 (N_2743,N_2131,N_2020);
nand U2744 (N_2744,N_2166,N_2400);
and U2745 (N_2745,N_2217,N_2011);
nand U2746 (N_2746,N_2473,N_2398);
and U2747 (N_2747,N_2230,N_2093);
or U2748 (N_2748,N_2331,N_2393);
or U2749 (N_2749,N_2194,N_2379);
or U2750 (N_2750,N_2168,N_2428);
or U2751 (N_2751,N_2051,N_2032);
nor U2752 (N_2752,N_2026,N_2145);
xor U2753 (N_2753,N_2319,N_2245);
or U2754 (N_2754,N_2298,N_2034);
and U2755 (N_2755,N_2369,N_2053);
and U2756 (N_2756,N_2265,N_2073);
and U2757 (N_2757,N_2248,N_2401);
nand U2758 (N_2758,N_2484,N_2177);
or U2759 (N_2759,N_2074,N_2087);
nor U2760 (N_2760,N_2089,N_2382);
and U2761 (N_2761,N_2478,N_2380);
and U2762 (N_2762,N_2300,N_2474);
and U2763 (N_2763,N_2266,N_2058);
or U2764 (N_2764,N_2493,N_2173);
or U2765 (N_2765,N_2299,N_2099);
nor U2766 (N_2766,N_2494,N_2067);
or U2767 (N_2767,N_2238,N_2420);
nand U2768 (N_2768,N_2145,N_2378);
nand U2769 (N_2769,N_2209,N_2207);
nor U2770 (N_2770,N_2114,N_2474);
and U2771 (N_2771,N_2087,N_2261);
or U2772 (N_2772,N_2021,N_2068);
nor U2773 (N_2773,N_2189,N_2119);
and U2774 (N_2774,N_2407,N_2341);
nand U2775 (N_2775,N_2499,N_2157);
nand U2776 (N_2776,N_2406,N_2313);
and U2777 (N_2777,N_2120,N_2086);
nor U2778 (N_2778,N_2127,N_2291);
nand U2779 (N_2779,N_2309,N_2063);
and U2780 (N_2780,N_2360,N_2057);
nand U2781 (N_2781,N_2169,N_2114);
and U2782 (N_2782,N_2305,N_2434);
and U2783 (N_2783,N_2269,N_2432);
nand U2784 (N_2784,N_2032,N_2030);
or U2785 (N_2785,N_2490,N_2034);
and U2786 (N_2786,N_2155,N_2120);
or U2787 (N_2787,N_2272,N_2358);
or U2788 (N_2788,N_2008,N_2211);
and U2789 (N_2789,N_2274,N_2415);
and U2790 (N_2790,N_2041,N_2047);
nand U2791 (N_2791,N_2136,N_2367);
or U2792 (N_2792,N_2171,N_2458);
or U2793 (N_2793,N_2345,N_2420);
and U2794 (N_2794,N_2042,N_2020);
nand U2795 (N_2795,N_2305,N_2218);
and U2796 (N_2796,N_2259,N_2167);
or U2797 (N_2797,N_2188,N_2317);
nand U2798 (N_2798,N_2342,N_2168);
nor U2799 (N_2799,N_2240,N_2061);
nor U2800 (N_2800,N_2287,N_2456);
and U2801 (N_2801,N_2243,N_2434);
nand U2802 (N_2802,N_2260,N_2421);
and U2803 (N_2803,N_2026,N_2004);
nand U2804 (N_2804,N_2051,N_2321);
nor U2805 (N_2805,N_2195,N_2313);
and U2806 (N_2806,N_2317,N_2483);
and U2807 (N_2807,N_2277,N_2045);
and U2808 (N_2808,N_2361,N_2004);
and U2809 (N_2809,N_2114,N_2266);
nand U2810 (N_2810,N_2129,N_2353);
nor U2811 (N_2811,N_2325,N_2104);
nand U2812 (N_2812,N_2329,N_2404);
nor U2813 (N_2813,N_2304,N_2085);
nand U2814 (N_2814,N_2456,N_2033);
nor U2815 (N_2815,N_2416,N_2472);
or U2816 (N_2816,N_2093,N_2076);
nor U2817 (N_2817,N_2493,N_2164);
and U2818 (N_2818,N_2205,N_2116);
or U2819 (N_2819,N_2436,N_2223);
nor U2820 (N_2820,N_2261,N_2069);
nand U2821 (N_2821,N_2211,N_2275);
nor U2822 (N_2822,N_2383,N_2296);
and U2823 (N_2823,N_2287,N_2176);
and U2824 (N_2824,N_2470,N_2029);
nor U2825 (N_2825,N_2256,N_2452);
nand U2826 (N_2826,N_2458,N_2013);
nor U2827 (N_2827,N_2157,N_2216);
or U2828 (N_2828,N_2042,N_2087);
and U2829 (N_2829,N_2105,N_2189);
nor U2830 (N_2830,N_2408,N_2094);
nor U2831 (N_2831,N_2003,N_2476);
nor U2832 (N_2832,N_2290,N_2492);
or U2833 (N_2833,N_2024,N_2058);
or U2834 (N_2834,N_2379,N_2238);
or U2835 (N_2835,N_2064,N_2423);
nor U2836 (N_2836,N_2073,N_2475);
xnor U2837 (N_2837,N_2321,N_2140);
nand U2838 (N_2838,N_2183,N_2482);
or U2839 (N_2839,N_2181,N_2234);
or U2840 (N_2840,N_2388,N_2369);
nor U2841 (N_2841,N_2046,N_2323);
and U2842 (N_2842,N_2373,N_2107);
and U2843 (N_2843,N_2243,N_2231);
or U2844 (N_2844,N_2149,N_2014);
nand U2845 (N_2845,N_2462,N_2039);
nor U2846 (N_2846,N_2214,N_2455);
or U2847 (N_2847,N_2462,N_2333);
and U2848 (N_2848,N_2255,N_2441);
nor U2849 (N_2849,N_2438,N_2046);
nand U2850 (N_2850,N_2444,N_2488);
nand U2851 (N_2851,N_2188,N_2362);
or U2852 (N_2852,N_2453,N_2135);
nand U2853 (N_2853,N_2265,N_2055);
nor U2854 (N_2854,N_2276,N_2059);
and U2855 (N_2855,N_2010,N_2403);
and U2856 (N_2856,N_2126,N_2185);
or U2857 (N_2857,N_2003,N_2211);
and U2858 (N_2858,N_2091,N_2280);
nor U2859 (N_2859,N_2229,N_2120);
and U2860 (N_2860,N_2017,N_2375);
nor U2861 (N_2861,N_2484,N_2096);
nor U2862 (N_2862,N_2406,N_2089);
nor U2863 (N_2863,N_2263,N_2377);
nand U2864 (N_2864,N_2395,N_2210);
nand U2865 (N_2865,N_2492,N_2062);
nor U2866 (N_2866,N_2030,N_2082);
xor U2867 (N_2867,N_2245,N_2316);
nand U2868 (N_2868,N_2040,N_2402);
nor U2869 (N_2869,N_2256,N_2483);
nor U2870 (N_2870,N_2316,N_2085);
nand U2871 (N_2871,N_2112,N_2119);
nor U2872 (N_2872,N_2325,N_2075);
nor U2873 (N_2873,N_2005,N_2028);
nor U2874 (N_2874,N_2267,N_2378);
nand U2875 (N_2875,N_2088,N_2184);
and U2876 (N_2876,N_2221,N_2227);
and U2877 (N_2877,N_2294,N_2094);
and U2878 (N_2878,N_2409,N_2186);
nand U2879 (N_2879,N_2104,N_2451);
and U2880 (N_2880,N_2411,N_2036);
nor U2881 (N_2881,N_2233,N_2130);
nand U2882 (N_2882,N_2123,N_2393);
and U2883 (N_2883,N_2287,N_2416);
nor U2884 (N_2884,N_2294,N_2024);
or U2885 (N_2885,N_2298,N_2455);
nor U2886 (N_2886,N_2091,N_2303);
or U2887 (N_2887,N_2005,N_2369);
or U2888 (N_2888,N_2044,N_2451);
or U2889 (N_2889,N_2492,N_2186);
nand U2890 (N_2890,N_2204,N_2274);
and U2891 (N_2891,N_2017,N_2285);
nor U2892 (N_2892,N_2115,N_2085);
and U2893 (N_2893,N_2486,N_2444);
and U2894 (N_2894,N_2271,N_2338);
xnor U2895 (N_2895,N_2023,N_2441);
nand U2896 (N_2896,N_2030,N_2300);
and U2897 (N_2897,N_2111,N_2080);
nor U2898 (N_2898,N_2455,N_2094);
nor U2899 (N_2899,N_2065,N_2346);
or U2900 (N_2900,N_2496,N_2127);
or U2901 (N_2901,N_2221,N_2102);
nand U2902 (N_2902,N_2454,N_2334);
nand U2903 (N_2903,N_2229,N_2263);
nand U2904 (N_2904,N_2471,N_2165);
or U2905 (N_2905,N_2253,N_2077);
xor U2906 (N_2906,N_2380,N_2131);
nand U2907 (N_2907,N_2245,N_2323);
and U2908 (N_2908,N_2135,N_2165);
and U2909 (N_2909,N_2009,N_2125);
nor U2910 (N_2910,N_2269,N_2281);
or U2911 (N_2911,N_2263,N_2178);
nor U2912 (N_2912,N_2145,N_2288);
and U2913 (N_2913,N_2001,N_2253);
nor U2914 (N_2914,N_2432,N_2464);
and U2915 (N_2915,N_2385,N_2290);
or U2916 (N_2916,N_2430,N_2498);
nor U2917 (N_2917,N_2215,N_2011);
or U2918 (N_2918,N_2401,N_2119);
and U2919 (N_2919,N_2052,N_2200);
nor U2920 (N_2920,N_2131,N_2017);
and U2921 (N_2921,N_2149,N_2090);
nand U2922 (N_2922,N_2177,N_2267);
nor U2923 (N_2923,N_2298,N_2014);
nand U2924 (N_2924,N_2017,N_2305);
and U2925 (N_2925,N_2273,N_2177);
nor U2926 (N_2926,N_2181,N_2459);
or U2927 (N_2927,N_2070,N_2069);
or U2928 (N_2928,N_2275,N_2005);
and U2929 (N_2929,N_2054,N_2124);
and U2930 (N_2930,N_2044,N_2358);
or U2931 (N_2931,N_2296,N_2287);
nand U2932 (N_2932,N_2426,N_2441);
and U2933 (N_2933,N_2216,N_2387);
or U2934 (N_2934,N_2346,N_2437);
nand U2935 (N_2935,N_2436,N_2161);
and U2936 (N_2936,N_2379,N_2340);
and U2937 (N_2937,N_2481,N_2034);
nor U2938 (N_2938,N_2015,N_2268);
or U2939 (N_2939,N_2484,N_2072);
nand U2940 (N_2940,N_2378,N_2417);
or U2941 (N_2941,N_2193,N_2468);
or U2942 (N_2942,N_2077,N_2015);
nand U2943 (N_2943,N_2331,N_2276);
nor U2944 (N_2944,N_2017,N_2127);
nor U2945 (N_2945,N_2186,N_2150);
nor U2946 (N_2946,N_2022,N_2487);
nand U2947 (N_2947,N_2395,N_2472);
nand U2948 (N_2948,N_2440,N_2025);
and U2949 (N_2949,N_2385,N_2458);
and U2950 (N_2950,N_2343,N_2132);
and U2951 (N_2951,N_2466,N_2049);
or U2952 (N_2952,N_2153,N_2205);
nand U2953 (N_2953,N_2111,N_2202);
or U2954 (N_2954,N_2212,N_2308);
or U2955 (N_2955,N_2426,N_2123);
or U2956 (N_2956,N_2015,N_2285);
nand U2957 (N_2957,N_2049,N_2034);
nor U2958 (N_2958,N_2468,N_2479);
and U2959 (N_2959,N_2298,N_2144);
nor U2960 (N_2960,N_2120,N_2009);
nor U2961 (N_2961,N_2420,N_2104);
and U2962 (N_2962,N_2357,N_2294);
or U2963 (N_2963,N_2169,N_2321);
nor U2964 (N_2964,N_2440,N_2277);
nand U2965 (N_2965,N_2062,N_2278);
nand U2966 (N_2966,N_2145,N_2241);
nor U2967 (N_2967,N_2328,N_2028);
and U2968 (N_2968,N_2117,N_2494);
nor U2969 (N_2969,N_2104,N_2365);
nor U2970 (N_2970,N_2008,N_2219);
nor U2971 (N_2971,N_2293,N_2160);
and U2972 (N_2972,N_2214,N_2255);
or U2973 (N_2973,N_2087,N_2301);
and U2974 (N_2974,N_2437,N_2065);
and U2975 (N_2975,N_2416,N_2358);
nand U2976 (N_2976,N_2127,N_2390);
and U2977 (N_2977,N_2300,N_2352);
nor U2978 (N_2978,N_2307,N_2293);
nand U2979 (N_2979,N_2356,N_2042);
or U2980 (N_2980,N_2037,N_2215);
and U2981 (N_2981,N_2151,N_2394);
nand U2982 (N_2982,N_2335,N_2366);
nand U2983 (N_2983,N_2138,N_2122);
nand U2984 (N_2984,N_2155,N_2072);
and U2985 (N_2985,N_2218,N_2256);
and U2986 (N_2986,N_2351,N_2207);
nor U2987 (N_2987,N_2485,N_2413);
or U2988 (N_2988,N_2297,N_2330);
and U2989 (N_2989,N_2343,N_2481);
and U2990 (N_2990,N_2132,N_2269);
nor U2991 (N_2991,N_2168,N_2092);
nor U2992 (N_2992,N_2053,N_2475);
and U2993 (N_2993,N_2100,N_2209);
or U2994 (N_2994,N_2186,N_2486);
or U2995 (N_2995,N_2327,N_2003);
or U2996 (N_2996,N_2030,N_2308);
nand U2997 (N_2997,N_2116,N_2109);
nand U2998 (N_2998,N_2111,N_2259);
or U2999 (N_2999,N_2393,N_2081);
and U3000 (N_3000,N_2645,N_2997);
xor U3001 (N_3001,N_2905,N_2708);
or U3002 (N_3002,N_2747,N_2989);
nand U3003 (N_3003,N_2845,N_2912);
and U3004 (N_3004,N_2643,N_2504);
nor U3005 (N_3005,N_2739,N_2808);
nor U3006 (N_3006,N_2733,N_2562);
or U3007 (N_3007,N_2571,N_2896);
and U3008 (N_3008,N_2518,N_2732);
or U3009 (N_3009,N_2952,N_2671);
xor U3010 (N_3010,N_2786,N_2678);
and U3011 (N_3011,N_2741,N_2855);
or U3012 (N_3012,N_2771,N_2692);
xor U3013 (N_3013,N_2667,N_2535);
and U3014 (N_3014,N_2584,N_2615);
or U3015 (N_3015,N_2529,N_2889);
nor U3016 (N_3016,N_2996,N_2956);
and U3017 (N_3017,N_2661,N_2795);
or U3018 (N_3018,N_2742,N_2632);
nand U3019 (N_3019,N_2903,N_2718);
nand U3020 (N_3020,N_2960,N_2804);
nand U3021 (N_3021,N_2843,N_2800);
and U3022 (N_3022,N_2983,N_2590);
nand U3023 (N_3023,N_2720,N_2908);
nand U3024 (N_3024,N_2766,N_2592);
nand U3025 (N_3025,N_2920,N_2677);
nor U3026 (N_3026,N_2775,N_2927);
nand U3027 (N_3027,N_2639,N_2698);
xnor U3028 (N_3028,N_2807,N_2982);
and U3029 (N_3029,N_2713,N_2743);
nor U3030 (N_3030,N_2744,N_2527);
and U3031 (N_3031,N_2803,N_2506);
or U3032 (N_3032,N_2642,N_2847);
xnor U3033 (N_3033,N_2971,N_2925);
nand U3034 (N_3034,N_2919,N_2611);
or U3035 (N_3035,N_2710,N_2703);
or U3036 (N_3036,N_2900,N_2687);
and U3037 (N_3037,N_2605,N_2964);
and U3038 (N_3038,N_2649,N_2929);
or U3039 (N_3039,N_2559,N_2898);
and U3040 (N_3040,N_2676,N_2561);
or U3041 (N_3041,N_2748,N_2773);
and U3042 (N_3042,N_2746,N_2838);
nand U3043 (N_3043,N_2503,N_2769);
and U3044 (N_3044,N_2831,N_2709);
nor U3045 (N_3045,N_2542,N_2862);
or U3046 (N_3046,N_2635,N_2958);
nand U3047 (N_3047,N_2754,N_2995);
nor U3048 (N_3048,N_2655,N_2824);
nand U3049 (N_3049,N_2953,N_2814);
nand U3050 (N_3050,N_2609,N_2602);
nor U3051 (N_3051,N_2863,N_2729);
or U3052 (N_3052,N_2500,N_2523);
nor U3053 (N_3053,N_2767,N_2586);
nor U3054 (N_3054,N_2944,N_2646);
and U3055 (N_3055,N_2805,N_2897);
xor U3056 (N_3056,N_2670,N_2869);
or U3057 (N_3057,N_2999,N_2726);
and U3058 (N_3058,N_2672,N_2848);
or U3059 (N_3059,N_2641,N_2839);
nor U3060 (N_3060,N_2505,N_2806);
nor U3061 (N_3061,N_2730,N_2521);
or U3062 (N_3062,N_2719,N_2531);
or U3063 (N_3063,N_2928,N_2954);
or U3064 (N_3064,N_2614,N_2731);
or U3065 (N_3065,N_2755,N_2516);
nand U3066 (N_3066,N_2626,N_2660);
and U3067 (N_3067,N_2631,N_2616);
nand U3068 (N_3068,N_2696,N_2986);
and U3069 (N_3069,N_2890,N_2858);
or U3070 (N_3070,N_2913,N_2572);
and U3071 (N_3071,N_2946,N_2520);
or U3072 (N_3072,N_2910,N_2809);
or U3073 (N_3073,N_2644,N_2966);
or U3074 (N_3074,N_2884,N_2875);
nor U3075 (N_3075,N_2549,N_2797);
or U3076 (N_3076,N_2622,N_2935);
nor U3077 (N_3077,N_2981,N_2510);
and U3078 (N_3078,N_2885,N_2714);
nor U3079 (N_3079,N_2711,N_2528);
nor U3080 (N_3080,N_2994,N_2853);
nor U3081 (N_3081,N_2914,N_2817);
xor U3082 (N_3082,N_2553,N_2856);
or U3083 (N_3083,N_2756,N_2801);
nand U3084 (N_3084,N_2544,N_2790);
nand U3085 (N_3085,N_2704,N_2979);
and U3086 (N_3086,N_2737,N_2793);
nor U3087 (N_3087,N_2923,N_2618);
nor U3088 (N_3088,N_2728,N_2826);
nor U3089 (N_3089,N_2859,N_2892);
or U3090 (N_3090,N_2513,N_2991);
nor U3091 (N_3091,N_2695,N_2955);
nand U3092 (N_3092,N_2582,N_2587);
nor U3093 (N_3093,N_2552,N_2844);
or U3094 (N_3094,N_2624,N_2723);
or U3095 (N_3095,N_2872,N_2595);
nand U3096 (N_3096,N_2781,N_2974);
xnor U3097 (N_3097,N_2691,N_2822);
nor U3098 (N_3098,N_2870,N_2757);
nand U3099 (N_3099,N_2721,N_2734);
nand U3100 (N_3100,N_2789,N_2599);
or U3101 (N_3101,N_2752,N_2705);
nand U3102 (N_3102,N_2621,N_2796);
or U3103 (N_3103,N_2819,N_2736);
or U3104 (N_3104,N_2835,N_2947);
nand U3105 (N_3105,N_2768,N_2603);
and U3106 (N_3106,N_2998,N_2735);
and U3107 (N_3107,N_2891,N_2868);
or U3108 (N_3108,N_2681,N_2950);
nand U3109 (N_3109,N_2895,N_2802);
nand U3110 (N_3110,N_2545,N_2640);
and U3111 (N_3111,N_2576,N_2990);
and U3112 (N_3112,N_2598,N_2828);
nor U3113 (N_3113,N_2680,N_2988);
xor U3114 (N_3114,N_2770,N_2765);
and U3115 (N_3115,N_2820,N_2985);
nand U3116 (N_3116,N_2568,N_2575);
nor U3117 (N_3117,N_2763,N_2970);
and U3118 (N_3118,N_2604,N_2532);
and U3119 (N_3119,N_2668,N_2537);
and U3120 (N_3120,N_2810,N_2688);
nand U3121 (N_3121,N_2893,N_2579);
or U3122 (N_3122,N_2593,N_2788);
xnor U3123 (N_3123,N_2894,N_2569);
nor U3124 (N_3124,N_2550,N_2627);
and U3125 (N_3125,N_2785,N_2509);
nand U3126 (N_3126,N_2556,N_2507);
or U3127 (N_3127,N_2682,N_2846);
nand U3128 (N_3128,N_2663,N_2623);
nand U3129 (N_3129,N_2749,N_2578);
and U3130 (N_3130,N_2530,N_2865);
and U3131 (N_3131,N_2969,N_2648);
nor U3132 (N_3132,N_2638,N_2906);
nand U3133 (N_3133,N_2980,N_2717);
nor U3134 (N_3134,N_2606,N_2782);
nand U3135 (N_3135,N_2750,N_2887);
and U3136 (N_3136,N_2787,N_2617);
nand U3137 (N_3137,N_2918,N_2697);
nand U3138 (N_3138,N_2931,N_2904);
nand U3139 (N_3139,N_2907,N_2613);
nor U3140 (N_3140,N_2777,N_2674);
nor U3141 (N_3141,N_2634,N_2973);
nand U3142 (N_3142,N_2876,N_2664);
nand U3143 (N_3143,N_2857,N_2759);
nor U3144 (N_3144,N_2938,N_2546);
xor U3145 (N_3145,N_2673,N_2564);
or U3146 (N_3146,N_2701,N_2880);
and U3147 (N_3147,N_2502,N_2783);
and U3148 (N_3148,N_2707,N_2877);
xor U3149 (N_3149,N_2833,N_2962);
nor U3150 (N_3150,N_2526,N_2840);
nand U3151 (N_3151,N_2849,N_2882);
xor U3152 (N_3152,N_2524,N_2596);
or U3153 (N_3153,N_2751,N_2647);
and U3154 (N_3154,N_2725,N_2818);
or U3155 (N_3155,N_2570,N_2861);
nand U3156 (N_3156,N_2968,N_2597);
and U3157 (N_3157,N_2939,N_2560);
nor U3158 (N_3158,N_2916,N_2554);
xor U3159 (N_3159,N_2656,N_2658);
nor U3160 (N_3160,N_2540,N_2784);
xor U3161 (N_3161,N_2629,N_2934);
and U3162 (N_3162,N_2949,N_2827);
and U3163 (N_3163,N_2825,N_2883);
nand U3164 (N_3164,N_2965,N_2779);
nor U3165 (N_3165,N_2901,N_2702);
or U3166 (N_3166,N_2851,N_2565);
or U3167 (N_3167,N_2555,N_2573);
nand U3168 (N_3168,N_2685,N_2984);
or U3169 (N_3169,N_2588,N_2992);
and U3170 (N_3170,N_2791,N_2583);
nor U3171 (N_3171,N_2548,N_2881);
and U3172 (N_3172,N_2963,N_2812);
and U3173 (N_3173,N_2610,N_2879);
nor U3174 (N_3174,N_2515,N_2601);
nand U3175 (N_3175,N_2620,N_2874);
nand U3176 (N_3176,N_2888,N_2651);
nand U3177 (N_3177,N_2712,N_2836);
nor U3178 (N_3178,N_2987,N_2666);
nor U3179 (N_3179,N_2608,N_2563);
nor U3180 (N_3180,N_2866,N_2976);
nand U3181 (N_3181,N_2580,N_2937);
nor U3182 (N_3182,N_2940,N_2689);
nor U3183 (N_3183,N_2821,N_2959);
nor U3184 (N_3184,N_2977,N_2878);
and U3185 (N_3185,N_2508,N_2792);
and U3186 (N_3186,N_2860,N_2841);
and U3187 (N_3187,N_2941,N_2753);
nor U3188 (N_3188,N_2899,N_2993);
nor U3189 (N_3189,N_2514,N_2972);
and U3190 (N_3190,N_2652,N_2830);
nor U3191 (N_3191,N_2745,N_2811);
and U3192 (N_3192,N_2815,N_2600);
or U3193 (N_3193,N_2536,N_2886);
nor U3194 (N_3194,N_2716,N_2538);
nor U3195 (N_3195,N_2758,N_2636);
and U3196 (N_3196,N_2942,N_2630);
and U3197 (N_3197,N_2921,N_2567);
and U3198 (N_3198,N_2961,N_2778);
and U3199 (N_3199,N_2837,N_2715);
nand U3200 (N_3200,N_2724,N_2936);
nor U3201 (N_3201,N_2924,N_2543);
nand U3202 (N_3202,N_2512,N_2541);
or U3203 (N_3203,N_2589,N_2700);
nand U3204 (N_3204,N_2915,N_2653);
or U3205 (N_3205,N_2585,N_2637);
or U3206 (N_3206,N_2776,N_2650);
xnor U3207 (N_3207,N_2581,N_2619);
and U3208 (N_3208,N_2799,N_2519);
or U3209 (N_3209,N_2774,N_2511);
or U3210 (N_3210,N_2762,N_2612);
or U3211 (N_3211,N_2657,N_2917);
or U3212 (N_3212,N_2686,N_2539);
or U3213 (N_3213,N_2690,N_2957);
or U3214 (N_3214,N_2558,N_2761);
nor U3215 (N_3215,N_2798,N_2557);
or U3216 (N_3216,N_2832,N_2930);
or U3217 (N_3217,N_2699,N_2607);
nand U3218 (N_3218,N_2722,N_2864);
or U3219 (N_3219,N_2625,N_2829);
nand U3220 (N_3220,N_2501,N_2943);
nand U3221 (N_3221,N_2654,N_2764);
or U3222 (N_3222,N_2675,N_2873);
or U3223 (N_3223,N_2547,N_2684);
nand U3224 (N_3224,N_2706,N_2911);
nand U3225 (N_3225,N_2594,N_2693);
and U3226 (N_3226,N_2926,N_2517);
and U3227 (N_3227,N_2850,N_2694);
or U3228 (N_3228,N_2948,N_2727);
or U3229 (N_3229,N_2933,N_2922);
nor U3230 (N_3230,N_2772,N_2871);
nor U3231 (N_3231,N_2816,N_2577);
or U3232 (N_3232,N_2967,N_2854);
nand U3233 (N_3233,N_2780,N_2738);
nor U3234 (N_3234,N_2522,N_2975);
and U3235 (N_3235,N_2633,N_2813);
nor U3236 (N_3236,N_2683,N_2909);
and U3237 (N_3237,N_2525,N_2945);
or U3238 (N_3238,N_2842,N_2534);
or U3239 (N_3239,N_2852,N_2794);
and U3240 (N_3240,N_2978,N_2628);
or U3241 (N_3241,N_2740,N_2662);
and U3242 (N_3242,N_2669,N_2823);
nand U3243 (N_3243,N_2533,N_2566);
or U3244 (N_3244,N_2902,N_2551);
and U3245 (N_3245,N_2951,N_2760);
and U3246 (N_3246,N_2932,N_2834);
nor U3247 (N_3247,N_2659,N_2591);
and U3248 (N_3248,N_2665,N_2679);
and U3249 (N_3249,N_2574,N_2867);
nand U3250 (N_3250,N_2796,N_2919);
or U3251 (N_3251,N_2986,N_2540);
or U3252 (N_3252,N_2856,N_2542);
or U3253 (N_3253,N_2501,N_2538);
xor U3254 (N_3254,N_2547,N_2658);
or U3255 (N_3255,N_2862,N_2835);
or U3256 (N_3256,N_2525,N_2522);
or U3257 (N_3257,N_2706,N_2869);
xor U3258 (N_3258,N_2661,N_2722);
and U3259 (N_3259,N_2709,N_2919);
or U3260 (N_3260,N_2664,N_2837);
nor U3261 (N_3261,N_2610,N_2795);
and U3262 (N_3262,N_2656,N_2509);
nor U3263 (N_3263,N_2940,N_2757);
and U3264 (N_3264,N_2702,N_2677);
nand U3265 (N_3265,N_2980,N_2894);
and U3266 (N_3266,N_2652,N_2683);
nand U3267 (N_3267,N_2837,N_2595);
nor U3268 (N_3268,N_2667,N_2677);
or U3269 (N_3269,N_2557,N_2582);
nand U3270 (N_3270,N_2762,N_2922);
nor U3271 (N_3271,N_2757,N_2982);
nand U3272 (N_3272,N_2787,N_2824);
and U3273 (N_3273,N_2504,N_2889);
and U3274 (N_3274,N_2981,N_2501);
or U3275 (N_3275,N_2740,N_2586);
nand U3276 (N_3276,N_2923,N_2738);
or U3277 (N_3277,N_2794,N_2966);
nand U3278 (N_3278,N_2987,N_2953);
or U3279 (N_3279,N_2675,N_2678);
nor U3280 (N_3280,N_2556,N_2950);
nor U3281 (N_3281,N_2629,N_2968);
nor U3282 (N_3282,N_2791,N_2605);
nor U3283 (N_3283,N_2510,N_2874);
and U3284 (N_3284,N_2763,N_2524);
nand U3285 (N_3285,N_2851,N_2502);
nand U3286 (N_3286,N_2960,N_2928);
nor U3287 (N_3287,N_2679,N_2688);
nand U3288 (N_3288,N_2858,N_2703);
and U3289 (N_3289,N_2526,N_2850);
and U3290 (N_3290,N_2567,N_2688);
and U3291 (N_3291,N_2743,N_2716);
nor U3292 (N_3292,N_2854,N_2788);
nand U3293 (N_3293,N_2788,N_2933);
xor U3294 (N_3294,N_2998,N_2861);
nor U3295 (N_3295,N_2769,N_2852);
and U3296 (N_3296,N_2812,N_2952);
nand U3297 (N_3297,N_2756,N_2606);
and U3298 (N_3298,N_2627,N_2504);
and U3299 (N_3299,N_2766,N_2829);
nor U3300 (N_3300,N_2903,N_2789);
nand U3301 (N_3301,N_2915,N_2942);
nor U3302 (N_3302,N_2966,N_2837);
nor U3303 (N_3303,N_2726,N_2978);
nor U3304 (N_3304,N_2700,N_2829);
or U3305 (N_3305,N_2669,N_2695);
or U3306 (N_3306,N_2823,N_2836);
and U3307 (N_3307,N_2903,N_2684);
nor U3308 (N_3308,N_2928,N_2583);
and U3309 (N_3309,N_2608,N_2856);
or U3310 (N_3310,N_2886,N_2608);
nand U3311 (N_3311,N_2695,N_2621);
or U3312 (N_3312,N_2576,N_2953);
and U3313 (N_3313,N_2704,N_2559);
nor U3314 (N_3314,N_2857,N_2664);
nor U3315 (N_3315,N_2686,N_2946);
or U3316 (N_3316,N_2945,N_2534);
or U3317 (N_3317,N_2859,N_2803);
and U3318 (N_3318,N_2657,N_2618);
nor U3319 (N_3319,N_2885,N_2596);
or U3320 (N_3320,N_2996,N_2600);
or U3321 (N_3321,N_2697,N_2570);
or U3322 (N_3322,N_2551,N_2771);
nand U3323 (N_3323,N_2769,N_2649);
xnor U3324 (N_3324,N_2831,N_2874);
and U3325 (N_3325,N_2777,N_2942);
nand U3326 (N_3326,N_2710,N_2732);
nand U3327 (N_3327,N_2908,N_2709);
or U3328 (N_3328,N_2724,N_2922);
nor U3329 (N_3329,N_2848,N_2880);
and U3330 (N_3330,N_2520,N_2954);
and U3331 (N_3331,N_2689,N_2976);
nand U3332 (N_3332,N_2974,N_2982);
nor U3333 (N_3333,N_2529,N_2807);
nand U3334 (N_3334,N_2968,N_2786);
and U3335 (N_3335,N_2838,N_2813);
nand U3336 (N_3336,N_2629,N_2661);
and U3337 (N_3337,N_2700,N_2815);
or U3338 (N_3338,N_2740,N_2954);
nand U3339 (N_3339,N_2938,N_2570);
nor U3340 (N_3340,N_2724,N_2683);
or U3341 (N_3341,N_2695,N_2767);
nor U3342 (N_3342,N_2798,N_2809);
or U3343 (N_3343,N_2877,N_2517);
and U3344 (N_3344,N_2927,N_2807);
or U3345 (N_3345,N_2701,N_2531);
nand U3346 (N_3346,N_2556,N_2635);
or U3347 (N_3347,N_2684,N_2591);
nand U3348 (N_3348,N_2898,N_2609);
and U3349 (N_3349,N_2670,N_2687);
nor U3350 (N_3350,N_2564,N_2759);
or U3351 (N_3351,N_2730,N_2870);
and U3352 (N_3352,N_2533,N_2727);
and U3353 (N_3353,N_2771,N_2891);
or U3354 (N_3354,N_2977,N_2570);
or U3355 (N_3355,N_2678,N_2956);
nor U3356 (N_3356,N_2607,N_2585);
nand U3357 (N_3357,N_2583,N_2764);
and U3358 (N_3358,N_2846,N_2739);
nand U3359 (N_3359,N_2507,N_2600);
or U3360 (N_3360,N_2660,N_2932);
nor U3361 (N_3361,N_2607,N_2719);
nor U3362 (N_3362,N_2973,N_2870);
and U3363 (N_3363,N_2818,N_2557);
xor U3364 (N_3364,N_2832,N_2824);
nor U3365 (N_3365,N_2819,N_2582);
and U3366 (N_3366,N_2605,N_2706);
nand U3367 (N_3367,N_2886,N_2575);
and U3368 (N_3368,N_2558,N_2878);
and U3369 (N_3369,N_2933,N_2531);
or U3370 (N_3370,N_2854,N_2963);
or U3371 (N_3371,N_2907,N_2762);
nand U3372 (N_3372,N_2588,N_2647);
and U3373 (N_3373,N_2736,N_2978);
nor U3374 (N_3374,N_2868,N_2779);
nor U3375 (N_3375,N_2676,N_2600);
nand U3376 (N_3376,N_2987,N_2664);
or U3377 (N_3377,N_2706,N_2682);
and U3378 (N_3378,N_2715,N_2976);
or U3379 (N_3379,N_2516,N_2571);
or U3380 (N_3380,N_2713,N_2563);
or U3381 (N_3381,N_2556,N_2768);
and U3382 (N_3382,N_2578,N_2758);
or U3383 (N_3383,N_2759,N_2925);
nor U3384 (N_3384,N_2560,N_2683);
xnor U3385 (N_3385,N_2780,N_2550);
or U3386 (N_3386,N_2675,N_2727);
and U3387 (N_3387,N_2661,N_2997);
or U3388 (N_3388,N_2544,N_2625);
nor U3389 (N_3389,N_2612,N_2832);
and U3390 (N_3390,N_2904,N_2757);
nor U3391 (N_3391,N_2998,N_2652);
or U3392 (N_3392,N_2929,N_2950);
xor U3393 (N_3393,N_2604,N_2824);
nor U3394 (N_3394,N_2749,N_2634);
nor U3395 (N_3395,N_2969,N_2956);
or U3396 (N_3396,N_2995,N_2556);
nand U3397 (N_3397,N_2876,N_2581);
or U3398 (N_3398,N_2882,N_2624);
or U3399 (N_3399,N_2924,N_2768);
nor U3400 (N_3400,N_2808,N_2623);
nor U3401 (N_3401,N_2962,N_2999);
nand U3402 (N_3402,N_2507,N_2877);
nand U3403 (N_3403,N_2959,N_2671);
nand U3404 (N_3404,N_2561,N_2533);
nand U3405 (N_3405,N_2655,N_2978);
nor U3406 (N_3406,N_2903,N_2768);
nor U3407 (N_3407,N_2831,N_2731);
or U3408 (N_3408,N_2994,N_2903);
or U3409 (N_3409,N_2791,N_2966);
nor U3410 (N_3410,N_2945,N_2879);
nand U3411 (N_3411,N_2809,N_2550);
or U3412 (N_3412,N_2674,N_2717);
nand U3413 (N_3413,N_2507,N_2832);
nand U3414 (N_3414,N_2740,N_2513);
nor U3415 (N_3415,N_2990,N_2967);
and U3416 (N_3416,N_2512,N_2879);
or U3417 (N_3417,N_2532,N_2818);
nor U3418 (N_3418,N_2771,N_2682);
nand U3419 (N_3419,N_2970,N_2611);
or U3420 (N_3420,N_2794,N_2532);
nor U3421 (N_3421,N_2723,N_2814);
or U3422 (N_3422,N_2523,N_2626);
and U3423 (N_3423,N_2671,N_2843);
or U3424 (N_3424,N_2615,N_2837);
and U3425 (N_3425,N_2626,N_2983);
or U3426 (N_3426,N_2592,N_2992);
nor U3427 (N_3427,N_2817,N_2839);
or U3428 (N_3428,N_2704,N_2703);
nor U3429 (N_3429,N_2766,N_2512);
nand U3430 (N_3430,N_2632,N_2964);
and U3431 (N_3431,N_2750,N_2703);
or U3432 (N_3432,N_2619,N_2778);
and U3433 (N_3433,N_2920,N_2999);
nor U3434 (N_3434,N_2937,N_2929);
and U3435 (N_3435,N_2946,N_2901);
nand U3436 (N_3436,N_2738,N_2849);
or U3437 (N_3437,N_2878,N_2918);
nor U3438 (N_3438,N_2647,N_2650);
or U3439 (N_3439,N_2541,N_2830);
nand U3440 (N_3440,N_2921,N_2746);
or U3441 (N_3441,N_2857,N_2566);
nor U3442 (N_3442,N_2720,N_2541);
nor U3443 (N_3443,N_2590,N_2740);
and U3444 (N_3444,N_2593,N_2543);
nand U3445 (N_3445,N_2808,N_2641);
and U3446 (N_3446,N_2926,N_2845);
nand U3447 (N_3447,N_2909,N_2655);
nand U3448 (N_3448,N_2791,N_2836);
nand U3449 (N_3449,N_2541,N_2632);
nor U3450 (N_3450,N_2581,N_2802);
and U3451 (N_3451,N_2829,N_2980);
nand U3452 (N_3452,N_2894,N_2757);
or U3453 (N_3453,N_2509,N_2592);
nor U3454 (N_3454,N_2711,N_2701);
and U3455 (N_3455,N_2660,N_2596);
xor U3456 (N_3456,N_2706,N_2688);
nor U3457 (N_3457,N_2980,N_2781);
nor U3458 (N_3458,N_2700,N_2527);
and U3459 (N_3459,N_2520,N_2916);
or U3460 (N_3460,N_2946,N_2841);
or U3461 (N_3461,N_2634,N_2534);
nand U3462 (N_3462,N_2894,N_2794);
or U3463 (N_3463,N_2941,N_2655);
nor U3464 (N_3464,N_2763,N_2807);
nor U3465 (N_3465,N_2661,N_2943);
nor U3466 (N_3466,N_2546,N_2644);
or U3467 (N_3467,N_2657,N_2635);
nor U3468 (N_3468,N_2743,N_2773);
or U3469 (N_3469,N_2803,N_2874);
nor U3470 (N_3470,N_2964,N_2631);
xor U3471 (N_3471,N_2867,N_2520);
nand U3472 (N_3472,N_2744,N_2878);
and U3473 (N_3473,N_2962,N_2888);
or U3474 (N_3474,N_2500,N_2646);
nor U3475 (N_3475,N_2796,N_2582);
or U3476 (N_3476,N_2564,N_2669);
nand U3477 (N_3477,N_2599,N_2935);
and U3478 (N_3478,N_2663,N_2604);
and U3479 (N_3479,N_2829,N_2599);
nand U3480 (N_3480,N_2549,N_2732);
or U3481 (N_3481,N_2649,N_2503);
and U3482 (N_3482,N_2743,N_2620);
nor U3483 (N_3483,N_2824,N_2742);
or U3484 (N_3484,N_2881,N_2555);
or U3485 (N_3485,N_2901,N_2766);
and U3486 (N_3486,N_2959,N_2757);
or U3487 (N_3487,N_2664,N_2924);
or U3488 (N_3488,N_2793,N_2650);
nand U3489 (N_3489,N_2728,N_2904);
or U3490 (N_3490,N_2671,N_2505);
or U3491 (N_3491,N_2782,N_2981);
and U3492 (N_3492,N_2963,N_2570);
or U3493 (N_3493,N_2722,N_2608);
nor U3494 (N_3494,N_2712,N_2642);
nor U3495 (N_3495,N_2938,N_2735);
or U3496 (N_3496,N_2643,N_2515);
or U3497 (N_3497,N_2780,N_2626);
nand U3498 (N_3498,N_2925,N_2811);
nor U3499 (N_3499,N_2912,N_2928);
and U3500 (N_3500,N_3208,N_3290);
or U3501 (N_3501,N_3334,N_3162);
nor U3502 (N_3502,N_3373,N_3492);
nand U3503 (N_3503,N_3420,N_3143);
or U3504 (N_3504,N_3391,N_3140);
nor U3505 (N_3505,N_3103,N_3308);
nand U3506 (N_3506,N_3266,N_3360);
or U3507 (N_3507,N_3458,N_3242);
nand U3508 (N_3508,N_3216,N_3304);
or U3509 (N_3509,N_3476,N_3269);
or U3510 (N_3510,N_3010,N_3037);
nor U3511 (N_3511,N_3370,N_3261);
nor U3512 (N_3512,N_3418,N_3267);
nor U3513 (N_3513,N_3053,N_3486);
nor U3514 (N_3514,N_3227,N_3243);
nand U3515 (N_3515,N_3152,N_3041);
and U3516 (N_3516,N_3314,N_3043);
nand U3517 (N_3517,N_3089,N_3045);
or U3518 (N_3518,N_3113,N_3099);
nor U3519 (N_3519,N_3477,N_3275);
and U3520 (N_3520,N_3487,N_3461);
nor U3521 (N_3521,N_3249,N_3198);
or U3522 (N_3522,N_3051,N_3022);
and U3523 (N_3523,N_3212,N_3398);
nor U3524 (N_3524,N_3450,N_3497);
xnor U3525 (N_3525,N_3276,N_3006);
nand U3526 (N_3526,N_3186,N_3352);
and U3527 (N_3527,N_3258,N_3170);
nand U3528 (N_3528,N_3288,N_3335);
nor U3529 (N_3529,N_3072,N_3439);
or U3530 (N_3530,N_3076,N_3021);
xor U3531 (N_3531,N_3218,N_3361);
nand U3532 (N_3532,N_3473,N_3091);
and U3533 (N_3533,N_3374,N_3322);
nand U3534 (N_3534,N_3027,N_3074);
or U3535 (N_3535,N_3038,N_3171);
and U3536 (N_3536,N_3465,N_3491);
nor U3537 (N_3537,N_3025,N_3395);
or U3538 (N_3538,N_3470,N_3084);
or U3539 (N_3539,N_3070,N_3100);
or U3540 (N_3540,N_3150,N_3196);
or U3541 (N_3541,N_3182,N_3286);
nand U3542 (N_3542,N_3189,N_3158);
nand U3543 (N_3543,N_3007,N_3188);
and U3544 (N_3544,N_3325,N_3036);
or U3545 (N_3545,N_3475,N_3108);
or U3546 (N_3546,N_3207,N_3134);
or U3547 (N_3547,N_3396,N_3382);
nand U3548 (N_3548,N_3190,N_3318);
nand U3549 (N_3549,N_3077,N_3431);
and U3550 (N_3550,N_3468,N_3333);
or U3551 (N_3551,N_3236,N_3016);
xnor U3552 (N_3552,N_3411,N_3058);
nand U3553 (N_3553,N_3394,N_3067);
nand U3554 (N_3554,N_3295,N_3346);
and U3555 (N_3555,N_3359,N_3093);
nand U3556 (N_3556,N_3422,N_3105);
nor U3557 (N_3557,N_3264,N_3408);
or U3558 (N_3558,N_3173,N_3272);
nand U3559 (N_3559,N_3324,N_3141);
nor U3560 (N_3560,N_3149,N_3485);
nand U3561 (N_3561,N_3353,N_3079);
nand U3562 (N_3562,N_3030,N_3148);
nor U3563 (N_3563,N_3047,N_3087);
nor U3564 (N_3564,N_3187,N_3104);
or U3565 (N_3565,N_3313,N_3315);
or U3566 (N_3566,N_3032,N_3445);
nand U3567 (N_3567,N_3112,N_3349);
xnor U3568 (N_3568,N_3493,N_3042);
nand U3569 (N_3569,N_3035,N_3452);
or U3570 (N_3570,N_3000,N_3110);
and U3571 (N_3571,N_3316,N_3034);
or U3572 (N_3572,N_3066,N_3031);
or U3573 (N_3573,N_3217,N_3252);
nor U3574 (N_3574,N_3244,N_3142);
or U3575 (N_3575,N_3240,N_3092);
or U3576 (N_3576,N_3434,N_3209);
nand U3577 (N_3577,N_3024,N_3192);
nand U3578 (N_3578,N_3341,N_3495);
nand U3579 (N_3579,N_3081,N_3116);
nor U3580 (N_3580,N_3416,N_3063);
nand U3581 (N_3581,N_3097,N_3046);
and U3582 (N_3582,N_3481,N_3156);
nor U3583 (N_3583,N_3375,N_3415);
or U3584 (N_3584,N_3277,N_3008);
nand U3585 (N_3585,N_3191,N_3090);
nand U3586 (N_3586,N_3062,N_3471);
nand U3587 (N_3587,N_3137,N_3178);
nor U3588 (N_3588,N_3466,N_3366);
nand U3589 (N_3589,N_3123,N_3238);
nand U3590 (N_3590,N_3273,N_3203);
and U3591 (N_3591,N_3457,N_3289);
nand U3592 (N_3592,N_3443,N_3132);
nor U3593 (N_3593,N_3383,N_3417);
xnor U3594 (N_3594,N_3159,N_3448);
and U3595 (N_3595,N_3280,N_3454);
nand U3596 (N_3596,N_3131,N_3489);
or U3597 (N_3597,N_3300,N_3384);
nor U3598 (N_3598,N_3393,N_3262);
or U3599 (N_3599,N_3407,N_3474);
nand U3600 (N_3600,N_3480,N_3145);
nor U3601 (N_3601,N_3163,N_3128);
or U3602 (N_3602,N_3364,N_3444);
xor U3603 (N_3603,N_3193,N_3181);
nor U3604 (N_3604,N_3301,N_3488);
nor U3605 (N_3605,N_3009,N_3328);
and U3606 (N_3606,N_3307,N_3257);
xnor U3607 (N_3607,N_3026,N_3119);
or U3608 (N_3608,N_3365,N_3094);
and U3609 (N_3609,N_3342,N_3437);
nand U3610 (N_3610,N_3409,N_3124);
nor U3611 (N_3611,N_3390,N_3378);
or U3612 (N_3612,N_3101,N_3185);
and U3613 (N_3613,N_3327,N_3166);
or U3614 (N_3614,N_3494,N_3020);
nand U3615 (N_3615,N_3179,N_3268);
and U3616 (N_3616,N_3326,N_3138);
nor U3617 (N_3617,N_3061,N_3048);
or U3618 (N_3618,N_3376,N_3496);
and U3619 (N_3619,N_3338,N_3019);
and U3620 (N_3620,N_3028,N_3371);
nor U3621 (N_3621,N_3282,N_3451);
nand U3622 (N_3622,N_3049,N_3293);
or U3623 (N_3623,N_3175,N_3424);
and U3624 (N_3624,N_3117,N_3115);
nand U3625 (N_3625,N_3214,N_3436);
nand U3626 (N_3626,N_3018,N_3292);
nor U3627 (N_3627,N_3385,N_3146);
nor U3628 (N_3628,N_3168,N_3005);
nand U3629 (N_3629,N_3050,N_3336);
nor U3630 (N_3630,N_3464,N_3291);
and U3631 (N_3631,N_3402,N_3004);
and U3632 (N_3632,N_3372,N_3201);
nor U3633 (N_3633,N_3498,N_3265);
nand U3634 (N_3634,N_3220,N_3380);
nand U3635 (N_3635,N_3073,N_3446);
nand U3636 (N_3636,N_3161,N_3144);
nor U3637 (N_3637,N_3102,N_3154);
nor U3638 (N_3638,N_3320,N_3427);
and U3639 (N_3639,N_3235,N_3263);
and U3640 (N_3640,N_3428,N_3096);
nand U3641 (N_3641,N_3248,N_3177);
nor U3642 (N_3642,N_3403,N_3270);
or U3643 (N_3643,N_3453,N_3147);
nand U3644 (N_3644,N_3195,N_3284);
nand U3645 (N_3645,N_3086,N_3151);
and U3646 (N_3646,N_3127,N_3069);
xnor U3647 (N_3647,N_3440,N_3245);
nand U3648 (N_3648,N_3347,N_3044);
nor U3649 (N_3649,N_3205,N_3377);
and U3650 (N_3650,N_3438,N_3223);
xnor U3651 (N_3651,N_3065,N_3399);
nand U3652 (N_3652,N_3331,N_3351);
or U3653 (N_3653,N_3157,N_3056);
or U3654 (N_3654,N_3472,N_3088);
or U3655 (N_3655,N_3467,N_3126);
nand U3656 (N_3656,N_3194,N_3226);
nand U3657 (N_3657,N_3368,N_3029);
nor U3658 (N_3658,N_3358,N_3160);
or U3659 (N_3659,N_3283,N_3312);
and U3660 (N_3660,N_3469,N_3456);
nand U3661 (N_3661,N_3350,N_3345);
or U3662 (N_3662,N_3299,N_3463);
or U3663 (N_3663,N_3183,N_3059);
nor U3664 (N_3664,N_3302,N_3397);
nor U3665 (N_3665,N_3211,N_3329);
and U3666 (N_3666,N_3122,N_3017);
nand U3667 (N_3667,N_3224,N_3165);
nand U3668 (N_3668,N_3432,N_3459);
and U3669 (N_3669,N_3139,N_3230);
and U3670 (N_3670,N_3323,N_3033);
nor U3671 (N_3671,N_3023,N_3111);
nand U3672 (N_3672,N_3169,N_3387);
nand U3673 (N_3673,N_3479,N_3256);
or U3674 (N_3674,N_3319,N_3241);
nand U3675 (N_3675,N_3490,N_3106);
or U3676 (N_3676,N_3085,N_3362);
xor U3677 (N_3677,N_3071,N_3015);
and U3678 (N_3678,N_3484,N_3098);
nand U3679 (N_3679,N_3250,N_3389);
nand U3680 (N_3680,N_3260,N_3210);
and U3681 (N_3681,N_3057,N_3414);
nand U3682 (N_3682,N_3309,N_3136);
nor U3683 (N_3683,N_3392,N_3413);
nor U3684 (N_3684,N_3388,N_3234);
or U3685 (N_3685,N_3426,N_3013);
and U3686 (N_3686,N_3172,N_3012);
or U3687 (N_3687,N_3499,N_3204);
and U3688 (N_3688,N_3251,N_3221);
or U3689 (N_3689,N_3297,N_3274);
nor U3690 (N_3690,N_3294,N_3213);
nor U3691 (N_3691,N_3180,N_3460);
or U3692 (N_3692,N_3311,N_3206);
or U3693 (N_3693,N_3441,N_3412);
nor U3694 (N_3694,N_3425,N_3231);
and U3695 (N_3695,N_3014,N_3400);
or U3696 (N_3696,N_3433,N_3011);
nand U3697 (N_3697,N_3068,N_3135);
or U3698 (N_3698,N_3303,N_3287);
nand U3699 (N_3699,N_3040,N_3176);
or U3700 (N_3700,N_3125,N_3174);
nand U3701 (N_3701,N_3430,N_3133);
nand U3702 (N_3702,N_3121,N_3321);
and U3703 (N_3703,N_3404,N_3306);
and U3704 (N_3704,N_3386,N_3167);
and U3705 (N_3705,N_3330,N_3202);
and U3706 (N_3706,N_3344,N_3109);
or U3707 (N_3707,N_3199,N_3219);
or U3708 (N_3708,N_3222,N_3055);
nand U3709 (N_3709,N_3423,N_3083);
nor U3710 (N_3710,N_3225,N_3060);
nor U3711 (N_3711,N_3357,N_3164);
nor U3712 (N_3712,N_3184,N_3410);
and U3713 (N_3713,N_3002,N_3340);
or U3714 (N_3714,N_3356,N_3075);
nor U3715 (N_3715,N_3405,N_3332);
nor U3716 (N_3716,N_3455,N_3379);
and U3717 (N_3717,N_3442,N_3429);
nand U3718 (N_3718,N_3401,N_3310);
and U3719 (N_3719,N_3285,N_3197);
or U3720 (N_3720,N_3130,N_3153);
and U3721 (N_3721,N_3054,N_3449);
nand U3722 (N_3722,N_3253,N_3228);
and U3723 (N_3723,N_3255,N_3200);
and U3724 (N_3724,N_3237,N_3118);
and U3725 (N_3725,N_3246,N_3229);
nor U3726 (N_3726,N_3039,N_3483);
nor U3727 (N_3727,N_3363,N_3337);
nor U3728 (N_3728,N_3120,N_3155);
nand U3729 (N_3729,N_3129,N_3259);
nand U3730 (N_3730,N_3233,N_3271);
nand U3731 (N_3731,N_3064,N_3281);
and U3732 (N_3732,N_3052,N_3419);
and U3733 (N_3733,N_3298,N_3279);
nand U3734 (N_3734,N_3232,N_3114);
nand U3735 (N_3735,N_3317,N_3478);
and U3736 (N_3736,N_3355,N_3482);
xor U3737 (N_3737,N_3080,N_3339);
nand U3738 (N_3738,N_3095,N_3215);
or U3739 (N_3739,N_3406,N_3435);
nand U3740 (N_3740,N_3107,N_3247);
nand U3741 (N_3741,N_3369,N_3367);
and U3742 (N_3742,N_3296,N_3254);
or U3743 (N_3743,N_3305,N_3082);
nand U3744 (N_3744,N_3239,N_3354);
or U3745 (N_3745,N_3381,N_3447);
and U3746 (N_3746,N_3278,N_3348);
nor U3747 (N_3747,N_3078,N_3421);
or U3748 (N_3748,N_3343,N_3001);
nor U3749 (N_3749,N_3462,N_3003);
nand U3750 (N_3750,N_3066,N_3117);
or U3751 (N_3751,N_3246,N_3161);
or U3752 (N_3752,N_3406,N_3150);
nor U3753 (N_3753,N_3123,N_3206);
nor U3754 (N_3754,N_3052,N_3071);
or U3755 (N_3755,N_3481,N_3329);
and U3756 (N_3756,N_3357,N_3407);
or U3757 (N_3757,N_3233,N_3141);
nor U3758 (N_3758,N_3361,N_3382);
and U3759 (N_3759,N_3491,N_3041);
or U3760 (N_3760,N_3030,N_3388);
or U3761 (N_3761,N_3312,N_3111);
or U3762 (N_3762,N_3433,N_3009);
and U3763 (N_3763,N_3029,N_3291);
and U3764 (N_3764,N_3053,N_3028);
and U3765 (N_3765,N_3295,N_3242);
nand U3766 (N_3766,N_3429,N_3303);
or U3767 (N_3767,N_3215,N_3469);
or U3768 (N_3768,N_3017,N_3030);
or U3769 (N_3769,N_3010,N_3299);
or U3770 (N_3770,N_3343,N_3287);
nor U3771 (N_3771,N_3182,N_3190);
nand U3772 (N_3772,N_3479,N_3371);
nand U3773 (N_3773,N_3408,N_3370);
nor U3774 (N_3774,N_3090,N_3343);
nand U3775 (N_3775,N_3272,N_3136);
nand U3776 (N_3776,N_3357,N_3415);
and U3777 (N_3777,N_3270,N_3465);
nor U3778 (N_3778,N_3174,N_3010);
xnor U3779 (N_3779,N_3279,N_3171);
and U3780 (N_3780,N_3451,N_3106);
and U3781 (N_3781,N_3065,N_3152);
and U3782 (N_3782,N_3147,N_3011);
nor U3783 (N_3783,N_3212,N_3327);
or U3784 (N_3784,N_3393,N_3305);
and U3785 (N_3785,N_3278,N_3362);
nor U3786 (N_3786,N_3232,N_3167);
nor U3787 (N_3787,N_3285,N_3123);
or U3788 (N_3788,N_3265,N_3085);
or U3789 (N_3789,N_3227,N_3072);
nand U3790 (N_3790,N_3214,N_3156);
and U3791 (N_3791,N_3357,N_3487);
and U3792 (N_3792,N_3116,N_3210);
and U3793 (N_3793,N_3478,N_3149);
nor U3794 (N_3794,N_3343,N_3364);
nand U3795 (N_3795,N_3209,N_3126);
nor U3796 (N_3796,N_3386,N_3136);
nor U3797 (N_3797,N_3494,N_3181);
and U3798 (N_3798,N_3079,N_3369);
nand U3799 (N_3799,N_3233,N_3478);
and U3800 (N_3800,N_3461,N_3309);
nand U3801 (N_3801,N_3459,N_3052);
nor U3802 (N_3802,N_3160,N_3201);
or U3803 (N_3803,N_3168,N_3380);
nand U3804 (N_3804,N_3331,N_3281);
or U3805 (N_3805,N_3264,N_3072);
nor U3806 (N_3806,N_3171,N_3378);
and U3807 (N_3807,N_3128,N_3412);
nor U3808 (N_3808,N_3012,N_3090);
nor U3809 (N_3809,N_3408,N_3214);
nor U3810 (N_3810,N_3050,N_3220);
nand U3811 (N_3811,N_3343,N_3054);
nor U3812 (N_3812,N_3445,N_3197);
or U3813 (N_3813,N_3379,N_3398);
nor U3814 (N_3814,N_3193,N_3307);
nor U3815 (N_3815,N_3148,N_3266);
and U3816 (N_3816,N_3107,N_3211);
nor U3817 (N_3817,N_3106,N_3134);
and U3818 (N_3818,N_3357,N_3066);
or U3819 (N_3819,N_3032,N_3093);
or U3820 (N_3820,N_3387,N_3383);
nand U3821 (N_3821,N_3399,N_3129);
nor U3822 (N_3822,N_3120,N_3274);
nor U3823 (N_3823,N_3202,N_3430);
nand U3824 (N_3824,N_3296,N_3251);
nor U3825 (N_3825,N_3255,N_3145);
nand U3826 (N_3826,N_3270,N_3244);
and U3827 (N_3827,N_3221,N_3372);
and U3828 (N_3828,N_3331,N_3144);
xor U3829 (N_3829,N_3465,N_3468);
nand U3830 (N_3830,N_3472,N_3349);
nand U3831 (N_3831,N_3354,N_3265);
nor U3832 (N_3832,N_3222,N_3336);
and U3833 (N_3833,N_3108,N_3450);
or U3834 (N_3834,N_3231,N_3464);
and U3835 (N_3835,N_3410,N_3235);
or U3836 (N_3836,N_3413,N_3363);
nor U3837 (N_3837,N_3334,N_3064);
and U3838 (N_3838,N_3230,N_3186);
nor U3839 (N_3839,N_3421,N_3094);
or U3840 (N_3840,N_3067,N_3202);
nand U3841 (N_3841,N_3037,N_3394);
nor U3842 (N_3842,N_3291,N_3395);
and U3843 (N_3843,N_3416,N_3136);
or U3844 (N_3844,N_3497,N_3473);
nand U3845 (N_3845,N_3107,N_3281);
and U3846 (N_3846,N_3039,N_3304);
nand U3847 (N_3847,N_3251,N_3081);
or U3848 (N_3848,N_3353,N_3205);
or U3849 (N_3849,N_3183,N_3423);
or U3850 (N_3850,N_3331,N_3261);
nand U3851 (N_3851,N_3275,N_3076);
nand U3852 (N_3852,N_3230,N_3132);
nand U3853 (N_3853,N_3225,N_3240);
nand U3854 (N_3854,N_3424,N_3161);
nand U3855 (N_3855,N_3263,N_3365);
or U3856 (N_3856,N_3259,N_3340);
nand U3857 (N_3857,N_3391,N_3138);
nor U3858 (N_3858,N_3151,N_3354);
nor U3859 (N_3859,N_3240,N_3270);
nor U3860 (N_3860,N_3141,N_3068);
or U3861 (N_3861,N_3438,N_3193);
nand U3862 (N_3862,N_3230,N_3398);
and U3863 (N_3863,N_3098,N_3306);
nor U3864 (N_3864,N_3223,N_3277);
and U3865 (N_3865,N_3485,N_3174);
and U3866 (N_3866,N_3063,N_3041);
and U3867 (N_3867,N_3097,N_3147);
and U3868 (N_3868,N_3024,N_3494);
nand U3869 (N_3869,N_3045,N_3234);
nand U3870 (N_3870,N_3466,N_3126);
xor U3871 (N_3871,N_3031,N_3120);
and U3872 (N_3872,N_3094,N_3295);
or U3873 (N_3873,N_3060,N_3449);
or U3874 (N_3874,N_3205,N_3486);
and U3875 (N_3875,N_3001,N_3309);
and U3876 (N_3876,N_3125,N_3456);
xnor U3877 (N_3877,N_3103,N_3043);
nor U3878 (N_3878,N_3424,N_3152);
nor U3879 (N_3879,N_3358,N_3254);
and U3880 (N_3880,N_3166,N_3095);
and U3881 (N_3881,N_3288,N_3416);
or U3882 (N_3882,N_3491,N_3125);
nand U3883 (N_3883,N_3296,N_3063);
and U3884 (N_3884,N_3222,N_3057);
nand U3885 (N_3885,N_3245,N_3032);
and U3886 (N_3886,N_3399,N_3219);
nand U3887 (N_3887,N_3159,N_3153);
nor U3888 (N_3888,N_3299,N_3295);
nand U3889 (N_3889,N_3495,N_3055);
nand U3890 (N_3890,N_3079,N_3472);
nor U3891 (N_3891,N_3180,N_3489);
or U3892 (N_3892,N_3308,N_3299);
nand U3893 (N_3893,N_3320,N_3323);
and U3894 (N_3894,N_3005,N_3309);
and U3895 (N_3895,N_3181,N_3386);
nor U3896 (N_3896,N_3406,N_3025);
xor U3897 (N_3897,N_3081,N_3267);
and U3898 (N_3898,N_3171,N_3198);
nor U3899 (N_3899,N_3167,N_3360);
or U3900 (N_3900,N_3011,N_3209);
or U3901 (N_3901,N_3203,N_3431);
or U3902 (N_3902,N_3082,N_3315);
and U3903 (N_3903,N_3053,N_3315);
nor U3904 (N_3904,N_3461,N_3164);
or U3905 (N_3905,N_3061,N_3450);
and U3906 (N_3906,N_3129,N_3470);
nor U3907 (N_3907,N_3467,N_3095);
nor U3908 (N_3908,N_3067,N_3048);
nor U3909 (N_3909,N_3239,N_3190);
nand U3910 (N_3910,N_3190,N_3345);
nand U3911 (N_3911,N_3471,N_3076);
xnor U3912 (N_3912,N_3326,N_3387);
and U3913 (N_3913,N_3471,N_3485);
nand U3914 (N_3914,N_3034,N_3270);
nor U3915 (N_3915,N_3346,N_3083);
nand U3916 (N_3916,N_3398,N_3346);
or U3917 (N_3917,N_3098,N_3418);
nand U3918 (N_3918,N_3104,N_3010);
nand U3919 (N_3919,N_3145,N_3406);
or U3920 (N_3920,N_3086,N_3007);
and U3921 (N_3921,N_3131,N_3286);
and U3922 (N_3922,N_3337,N_3147);
nor U3923 (N_3923,N_3360,N_3285);
nand U3924 (N_3924,N_3354,N_3355);
nor U3925 (N_3925,N_3265,N_3396);
and U3926 (N_3926,N_3087,N_3394);
nor U3927 (N_3927,N_3134,N_3080);
nand U3928 (N_3928,N_3474,N_3241);
nand U3929 (N_3929,N_3461,N_3495);
nor U3930 (N_3930,N_3467,N_3227);
and U3931 (N_3931,N_3240,N_3132);
nor U3932 (N_3932,N_3320,N_3062);
nand U3933 (N_3933,N_3373,N_3125);
or U3934 (N_3934,N_3452,N_3126);
nor U3935 (N_3935,N_3350,N_3405);
nand U3936 (N_3936,N_3130,N_3391);
xnor U3937 (N_3937,N_3468,N_3210);
or U3938 (N_3938,N_3100,N_3435);
and U3939 (N_3939,N_3334,N_3354);
nor U3940 (N_3940,N_3026,N_3493);
nand U3941 (N_3941,N_3009,N_3486);
or U3942 (N_3942,N_3048,N_3131);
nor U3943 (N_3943,N_3026,N_3365);
nor U3944 (N_3944,N_3495,N_3408);
nor U3945 (N_3945,N_3098,N_3298);
and U3946 (N_3946,N_3314,N_3131);
nor U3947 (N_3947,N_3321,N_3305);
nor U3948 (N_3948,N_3417,N_3298);
nand U3949 (N_3949,N_3345,N_3014);
or U3950 (N_3950,N_3295,N_3312);
or U3951 (N_3951,N_3099,N_3186);
and U3952 (N_3952,N_3247,N_3063);
nand U3953 (N_3953,N_3266,N_3251);
nor U3954 (N_3954,N_3485,N_3026);
or U3955 (N_3955,N_3223,N_3230);
nor U3956 (N_3956,N_3187,N_3250);
nor U3957 (N_3957,N_3091,N_3128);
or U3958 (N_3958,N_3185,N_3175);
or U3959 (N_3959,N_3141,N_3221);
nand U3960 (N_3960,N_3105,N_3397);
and U3961 (N_3961,N_3222,N_3388);
or U3962 (N_3962,N_3140,N_3430);
nor U3963 (N_3963,N_3027,N_3081);
and U3964 (N_3964,N_3208,N_3299);
or U3965 (N_3965,N_3180,N_3322);
or U3966 (N_3966,N_3242,N_3192);
nand U3967 (N_3967,N_3455,N_3300);
nor U3968 (N_3968,N_3032,N_3000);
or U3969 (N_3969,N_3002,N_3012);
or U3970 (N_3970,N_3242,N_3369);
and U3971 (N_3971,N_3006,N_3411);
nand U3972 (N_3972,N_3472,N_3300);
nor U3973 (N_3973,N_3095,N_3272);
nand U3974 (N_3974,N_3388,N_3426);
nor U3975 (N_3975,N_3044,N_3003);
nand U3976 (N_3976,N_3174,N_3032);
or U3977 (N_3977,N_3452,N_3281);
or U3978 (N_3978,N_3337,N_3297);
or U3979 (N_3979,N_3367,N_3386);
nand U3980 (N_3980,N_3162,N_3360);
or U3981 (N_3981,N_3351,N_3059);
and U3982 (N_3982,N_3270,N_3097);
and U3983 (N_3983,N_3127,N_3369);
and U3984 (N_3984,N_3178,N_3068);
nor U3985 (N_3985,N_3422,N_3255);
and U3986 (N_3986,N_3108,N_3452);
and U3987 (N_3987,N_3379,N_3381);
or U3988 (N_3988,N_3473,N_3376);
or U3989 (N_3989,N_3247,N_3485);
nand U3990 (N_3990,N_3447,N_3320);
nor U3991 (N_3991,N_3379,N_3123);
or U3992 (N_3992,N_3097,N_3168);
and U3993 (N_3993,N_3064,N_3349);
and U3994 (N_3994,N_3302,N_3069);
and U3995 (N_3995,N_3482,N_3431);
and U3996 (N_3996,N_3316,N_3487);
nor U3997 (N_3997,N_3347,N_3411);
nor U3998 (N_3998,N_3404,N_3158);
nor U3999 (N_3999,N_3160,N_3349);
nor U4000 (N_4000,N_3878,N_3919);
xnor U4001 (N_4001,N_3613,N_3676);
or U4002 (N_4002,N_3629,N_3913);
or U4003 (N_4003,N_3831,N_3936);
nand U4004 (N_4004,N_3882,N_3589);
xor U4005 (N_4005,N_3517,N_3925);
nand U4006 (N_4006,N_3844,N_3937);
nand U4007 (N_4007,N_3569,N_3969);
or U4008 (N_4008,N_3781,N_3588);
nor U4009 (N_4009,N_3624,N_3680);
nor U4010 (N_4010,N_3957,N_3533);
or U4011 (N_4011,N_3574,N_3714);
nor U4012 (N_4012,N_3631,N_3880);
nand U4013 (N_4013,N_3861,N_3618);
or U4014 (N_4014,N_3557,N_3756);
nand U4015 (N_4015,N_3621,N_3702);
and U4016 (N_4016,N_3724,N_3535);
or U4017 (N_4017,N_3839,N_3924);
nor U4018 (N_4018,N_3748,N_3635);
nor U4019 (N_4019,N_3863,N_3633);
nor U4020 (N_4020,N_3955,N_3565);
and U4021 (N_4021,N_3835,N_3587);
nor U4022 (N_4022,N_3653,N_3775);
or U4023 (N_4023,N_3703,N_3753);
nor U4024 (N_4024,N_3763,N_3547);
nand U4025 (N_4025,N_3738,N_3644);
nor U4026 (N_4026,N_3899,N_3729);
and U4027 (N_4027,N_3776,N_3512);
or U4028 (N_4028,N_3843,N_3812);
and U4029 (N_4029,N_3968,N_3834);
and U4030 (N_4030,N_3874,N_3506);
or U4031 (N_4031,N_3890,N_3966);
nand U4032 (N_4032,N_3599,N_3509);
or U4033 (N_4033,N_3755,N_3879);
and U4034 (N_4034,N_3668,N_3672);
or U4035 (N_4035,N_3981,N_3671);
or U4036 (N_4036,N_3986,N_3773);
xnor U4037 (N_4037,N_3989,N_3933);
xnor U4038 (N_4038,N_3605,N_3850);
or U4039 (N_4039,N_3941,N_3751);
nand U4040 (N_4040,N_3750,N_3660);
nand U4041 (N_4041,N_3600,N_3868);
or U4042 (N_4042,N_3571,N_3687);
nor U4043 (N_4043,N_3708,N_3523);
nand U4044 (N_4044,N_3577,N_3749);
or U4045 (N_4045,N_3760,N_3594);
or U4046 (N_4046,N_3764,N_3570);
nand U4047 (N_4047,N_3884,N_3910);
and U4048 (N_4048,N_3527,N_3978);
nand U4049 (N_4049,N_3946,N_3746);
or U4050 (N_4050,N_3581,N_3980);
nor U4051 (N_4051,N_3711,N_3656);
xnor U4052 (N_4052,N_3740,N_3950);
nand U4053 (N_4053,N_3922,N_3897);
nand U4054 (N_4054,N_3757,N_3584);
and U4055 (N_4055,N_3848,N_3603);
or U4056 (N_4056,N_3615,N_3716);
nand U4057 (N_4057,N_3513,N_3530);
nor U4058 (N_4058,N_3625,N_3885);
or U4059 (N_4059,N_3858,N_3709);
nand U4060 (N_4060,N_3705,N_3999);
nand U4061 (N_4061,N_3555,N_3860);
and U4062 (N_4062,N_3893,N_3731);
nand U4063 (N_4063,N_3862,N_3632);
or U4064 (N_4064,N_3501,N_3568);
and U4065 (N_4065,N_3659,N_3872);
nand U4066 (N_4066,N_3820,N_3744);
and U4067 (N_4067,N_3601,N_3567);
or U4068 (N_4068,N_3840,N_3892);
nor U4069 (N_4069,N_3602,N_3847);
nor U4070 (N_4070,N_3528,N_3507);
nand U4071 (N_4071,N_3944,N_3909);
nand U4072 (N_4072,N_3675,N_3636);
nand U4073 (N_4073,N_3611,N_3802);
nor U4074 (N_4074,N_3550,N_3593);
or U4075 (N_4075,N_3901,N_3795);
and U4076 (N_4076,N_3699,N_3595);
nor U4077 (N_4077,N_3647,N_3855);
and U4078 (N_4078,N_3526,N_3640);
or U4079 (N_4079,N_3622,N_3681);
and U4080 (N_4080,N_3902,N_3511);
nand U4081 (N_4081,N_3789,N_3832);
or U4082 (N_4082,N_3679,N_3674);
nand U4083 (N_4083,N_3984,N_3650);
and U4084 (N_4084,N_3772,N_3995);
and U4085 (N_4085,N_3572,N_3634);
nand U4086 (N_4086,N_3792,N_3742);
and U4087 (N_4087,N_3685,N_3726);
nand U4088 (N_4088,N_3975,N_3964);
nor U4089 (N_4089,N_3816,N_3918);
or U4090 (N_4090,N_3962,N_3700);
nand U4091 (N_4091,N_3585,N_3707);
xnor U4092 (N_4092,N_3906,N_3551);
xor U4093 (N_4093,N_3616,N_3544);
nor U4094 (N_4094,N_3898,N_3651);
and U4095 (N_4095,N_3943,N_3727);
and U4096 (N_4096,N_3940,N_3607);
or U4097 (N_4097,N_3721,N_3733);
nor U4098 (N_4098,N_3983,N_3626);
nor U4099 (N_4099,N_3719,N_3911);
nand U4100 (N_4100,N_3683,N_3871);
or U4101 (N_4101,N_3710,N_3852);
and U4102 (N_4102,N_3520,N_3536);
nand U4103 (N_4103,N_3876,N_3896);
and U4104 (N_4104,N_3737,N_3851);
or U4105 (N_4105,N_3643,N_3967);
and U4106 (N_4106,N_3809,N_3697);
or U4107 (N_4107,N_3998,N_3974);
and U4108 (N_4108,N_3556,N_3889);
and U4109 (N_4109,N_3838,N_3688);
and U4110 (N_4110,N_3873,N_3785);
xnor U4111 (N_4111,N_3928,N_3591);
nand U4112 (N_4112,N_3560,N_3662);
and U4113 (N_4113,N_3658,N_3916);
nor U4114 (N_4114,N_3519,N_3692);
nand U4115 (N_4115,N_3657,N_3768);
or U4116 (N_4116,N_3783,N_3821);
and U4117 (N_4117,N_3508,N_3583);
nor U4118 (N_4118,N_3796,N_3881);
nand U4119 (N_4119,N_3597,N_3867);
or U4120 (N_4120,N_3539,N_3542);
or U4121 (N_4121,N_3942,N_3664);
nor U4122 (N_4122,N_3985,N_3759);
and U4123 (N_4123,N_3690,N_3915);
and U4124 (N_4124,N_3661,N_3713);
and U4125 (N_4125,N_3804,N_3805);
nand U4126 (N_4126,N_3514,N_3817);
or U4127 (N_4127,N_3865,N_3648);
nor U4128 (N_4128,N_3537,N_3563);
nand U4129 (N_4129,N_3515,N_3504);
or U4130 (N_4130,N_3818,N_3842);
nor U4131 (N_4131,N_3931,N_3770);
and U4132 (N_4132,N_3689,N_3694);
or U4133 (N_4133,N_3698,N_3610);
or U4134 (N_4134,N_3997,N_3900);
nor U4135 (N_4135,N_3609,N_3988);
or U4136 (N_4136,N_3604,N_3956);
nor U4137 (N_4137,N_3786,N_3866);
or U4138 (N_4138,N_3534,N_3573);
or U4139 (N_4139,N_3546,N_3830);
or U4140 (N_4140,N_3628,N_3532);
nor U4141 (N_4141,N_3845,N_3903);
and U4142 (N_4142,N_3833,N_3972);
and U4143 (N_4143,N_3883,N_3641);
or U4144 (N_4144,N_3828,N_3991);
or U4145 (N_4145,N_3951,N_3723);
nor U4146 (N_4146,N_3525,N_3758);
or U4147 (N_4147,N_3778,N_3645);
nand U4148 (N_4148,N_3678,N_3728);
nor U4149 (N_4149,N_3920,N_3917);
nand U4150 (N_4150,N_3979,N_3766);
nand U4151 (N_4151,N_3500,N_3971);
nand U4152 (N_4152,N_3576,N_3806);
or U4153 (N_4153,N_3620,N_3666);
or U4154 (N_4154,N_3538,N_3811);
nor U4155 (N_4155,N_3958,N_3667);
nand U4156 (N_4156,N_3965,N_3543);
or U4157 (N_4157,N_3977,N_3586);
nand U4158 (N_4158,N_3747,N_3935);
and U4159 (N_4159,N_3794,N_3887);
nor U4160 (N_4160,N_3797,N_3566);
nand U4161 (N_4161,N_3859,N_3695);
nor U4162 (N_4162,N_3822,N_3559);
nor U4163 (N_4163,N_3947,N_3790);
xor U4164 (N_4164,N_3548,N_3655);
and U4165 (N_4165,N_3800,N_3743);
nor U4166 (N_4166,N_3929,N_3803);
nor U4167 (N_4167,N_3754,N_3725);
nor U4168 (N_4168,N_3562,N_3665);
or U4169 (N_4169,N_3788,N_3907);
nand U4170 (N_4170,N_3619,N_3718);
nand U4171 (N_4171,N_3934,N_3735);
nand U4172 (N_4172,N_3580,N_3992);
nand U4173 (N_4173,N_3837,N_3720);
nand U4174 (N_4174,N_3734,N_3627);
nor U4175 (N_4175,N_3684,N_3518);
nand U4176 (N_4176,N_3953,N_3875);
nand U4177 (N_4177,N_3706,N_3612);
and U4178 (N_4178,N_3891,N_3701);
nand U4179 (N_4179,N_3669,N_3696);
nor U4180 (N_4180,N_3853,N_3846);
and U4181 (N_4181,N_3505,N_3782);
or U4182 (N_4182,N_3704,N_3787);
and U4183 (N_4183,N_3793,N_3693);
and U4184 (N_4184,N_3960,N_3904);
or U4185 (N_4185,N_3654,N_3730);
or U4186 (N_4186,N_3745,N_3545);
nand U4187 (N_4187,N_3712,N_3982);
nand U4188 (N_4188,N_3663,N_3912);
nor U4189 (N_4189,N_3774,N_3529);
nand U4190 (N_4190,N_3938,N_3976);
nor U4191 (N_4191,N_3606,N_3762);
and U4192 (N_4192,N_3948,N_3810);
nor U4193 (N_4193,N_3639,N_3895);
nor U4194 (N_4194,N_3854,N_3791);
and U4195 (N_4195,N_3814,N_3558);
or U4196 (N_4196,N_3932,N_3784);
and U4197 (N_4197,N_3561,N_3638);
nand U4198 (N_4198,N_3522,N_3823);
and U4199 (N_4199,N_3717,N_3973);
and U4200 (N_4200,N_3825,N_3767);
or U4201 (N_4201,N_3914,N_3670);
and U4202 (N_4202,N_3908,N_3614);
nor U4203 (N_4203,N_3864,N_3780);
and U4204 (N_4204,N_3815,N_3637);
and U4205 (N_4205,N_3799,N_3813);
nor U4206 (N_4206,N_3798,N_3722);
and U4207 (N_4207,N_3769,N_3970);
nor U4208 (N_4208,N_3779,N_3959);
nand U4209 (N_4209,N_3579,N_3877);
and U4210 (N_4210,N_3888,N_3596);
nor U4211 (N_4211,N_3869,N_3554);
nor U4212 (N_4212,N_3549,N_3553);
xor U4213 (N_4213,N_3930,N_3777);
or U4214 (N_4214,N_3961,N_3949);
or U4215 (N_4215,N_3598,N_3715);
or U4216 (N_4216,N_3510,N_3945);
nor U4217 (N_4217,N_3590,N_3836);
nor U4218 (N_4218,N_3617,N_3927);
nand U4219 (N_4219,N_3524,N_3923);
nand U4220 (N_4220,N_3856,N_3739);
and U4221 (N_4221,N_3686,N_3926);
nor U4222 (N_4222,N_3954,N_3582);
or U4223 (N_4223,N_3531,N_3552);
or U4224 (N_4224,N_3808,N_3649);
nand U4225 (N_4225,N_3578,N_3765);
and U4226 (N_4226,N_3963,N_3673);
or U4227 (N_4227,N_3608,N_3503);
nand U4228 (N_4228,N_3819,N_3801);
nor U4229 (N_4229,N_3752,N_3732);
nor U4230 (N_4230,N_3592,N_3642);
and U4231 (N_4231,N_3996,N_3807);
and U4232 (N_4232,N_3646,N_3886);
or U4233 (N_4233,N_3829,N_3826);
nand U4234 (N_4234,N_3736,N_3741);
or U4235 (N_4235,N_3841,N_3952);
nand U4236 (N_4236,N_3682,N_3771);
or U4237 (N_4237,N_3521,N_3827);
or U4238 (N_4238,N_3516,N_3623);
or U4239 (N_4239,N_3824,N_3630);
xor U4240 (N_4240,N_3870,N_3990);
or U4241 (N_4241,N_3652,N_3691);
nor U4242 (N_4242,N_3921,N_3849);
or U4243 (N_4243,N_3905,N_3575);
and U4244 (N_4244,N_3761,N_3993);
and U4245 (N_4245,N_3994,N_3857);
and U4246 (N_4246,N_3677,N_3540);
nor U4247 (N_4247,N_3502,N_3987);
and U4248 (N_4248,N_3894,N_3564);
nand U4249 (N_4249,N_3541,N_3939);
nor U4250 (N_4250,N_3932,N_3813);
nor U4251 (N_4251,N_3758,N_3914);
nor U4252 (N_4252,N_3747,N_3527);
nor U4253 (N_4253,N_3687,N_3760);
xnor U4254 (N_4254,N_3808,N_3522);
nor U4255 (N_4255,N_3654,N_3801);
nor U4256 (N_4256,N_3598,N_3931);
and U4257 (N_4257,N_3775,N_3924);
and U4258 (N_4258,N_3696,N_3821);
or U4259 (N_4259,N_3652,N_3916);
or U4260 (N_4260,N_3756,N_3881);
xnor U4261 (N_4261,N_3906,N_3724);
nor U4262 (N_4262,N_3966,N_3604);
nand U4263 (N_4263,N_3987,N_3848);
or U4264 (N_4264,N_3685,N_3681);
and U4265 (N_4265,N_3628,N_3854);
or U4266 (N_4266,N_3559,N_3984);
nand U4267 (N_4267,N_3881,N_3566);
nor U4268 (N_4268,N_3965,N_3537);
nand U4269 (N_4269,N_3922,N_3643);
nor U4270 (N_4270,N_3916,N_3946);
and U4271 (N_4271,N_3794,N_3633);
nor U4272 (N_4272,N_3630,N_3803);
and U4273 (N_4273,N_3964,N_3872);
or U4274 (N_4274,N_3960,N_3825);
or U4275 (N_4275,N_3981,N_3623);
and U4276 (N_4276,N_3520,N_3684);
or U4277 (N_4277,N_3551,N_3958);
nor U4278 (N_4278,N_3525,N_3778);
nand U4279 (N_4279,N_3777,N_3523);
or U4280 (N_4280,N_3826,N_3897);
or U4281 (N_4281,N_3899,N_3747);
or U4282 (N_4282,N_3968,N_3700);
nor U4283 (N_4283,N_3690,N_3574);
nor U4284 (N_4284,N_3616,N_3743);
nor U4285 (N_4285,N_3520,N_3808);
nand U4286 (N_4286,N_3519,N_3568);
nor U4287 (N_4287,N_3720,N_3786);
nor U4288 (N_4288,N_3753,N_3859);
nand U4289 (N_4289,N_3646,N_3971);
nor U4290 (N_4290,N_3665,N_3907);
nand U4291 (N_4291,N_3671,N_3534);
or U4292 (N_4292,N_3839,N_3506);
nor U4293 (N_4293,N_3976,N_3726);
nand U4294 (N_4294,N_3733,N_3826);
nor U4295 (N_4295,N_3616,N_3916);
or U4296 (N_4296,N_3750,N_3747);
and U4297 (N_4297,N_3925,N_3931);
and U4298 (N_4298,N_3656,N_3842);
nor U4299 (N_4299,N_3927,N_3603);
or U4300 (N_4300,N_3912,N_3671);
or U4301 (N_4301,N_3997,N_3550);
nor U4302 (N_4302,N_3829,N_3627);
and U4303 (N_4303,N_3573,N_3769);
nand U4304 (N_4304,N_3777,N_3812);
nor U4305 (N_4305,N_3910,N_3955);
or U4306 (N_4306,N_3913,N_3930);
and U4307 (N_4307,N_3828,N_3913);
and U4308 (N_4308,N_3529,N_3948);
nor U4309 (N_4309,N_3551,N_3525);
nand U4310 (N_4310,N_3585,N_3519);
nor U4311 (N_4311,N_3710,N_3703);
nor U4312 (N_4312,N_3751,N_3657);
nand U4313 (N_4313,N_3745,N_3638);
and U4314 (N_4314,N_3593,N_3970);
and U4315 (N_4315,N_3650,N_3610);
or U4316 (N_4316,N_3503,N_3759);
and U4317 (N_4317,N_3944,N_3813);
and U4318 (N_4318,N_3899,N_3720);
nor U4319 (N_4319,N_3528,N_3573);
nor U4320 (N_4320,N_3840,N_3882);
nand U4321 (N_4321,N_3931,N_3675);
and U4322 (N_4322,N_3912,N_3686);
nand U4323 (N_4323,N_3957,N_3766);
or U4324 (N_4324,N_3663,N_3536);
nand U4325 (N_4325,N_3986,N_3880);
nand U4326 (N_4326,N_3870,N_3501);
or U4327 (N_4327,N_3861,N_3573);
nor U4328 (N_4328,N_3847,N_3991);
or U4329 (N_4329,N_3852,N_3825);
nor U4330 (N_4330,N_3619,N_3939);
nand U4331 (N_4331,N_3918,N_3618);
nand U4332 (N_4332,N_3653,N_3986);
or U4333 (N_4333,N_3956,N_3551);
and U4334 (N_4334,N_3907,N_3557);
nor U4335 (N_4335,N_3897,N_3784);
nor U4336 (N_4336,N_3535,N_3898);
nor U4337 (N_4337,N_3888,N_3504);
nor U4338 (N_4338,N_3603,N_3563);
nor U4339 (N_4339,N_3993,N_3700);
nand U4340 (N_4340,N_3811,N_3661);
and U4341 (N_4341,N_3689,N_3561);
nand U4342 (N_4342,N_3564,N_3548);
and U4343 (N_4343,N_3834,N_3660);
or U4344 (N_4344,N_3549,N_3956);
nand U4345 (N_4345,N_3974,N_3565);
and U4346 (N_4346,N_3961,N_3946);
or U4347 (N_4347,N_3872,N_3781);
nor U4348 (N_4348,N_3677,N_3511);
nor U4349 (N_4349,N_3836,N_3937);
or U4350 (N_4350,N_3635,N_3682);
or U4351 (N_4351,N_3977,N_3873);
and U4352 (N_4352,N_3715,N_3825);
nand U4353 (N_4353,N_3792,N_3519);
nor U4354 (N_4354,N_3785,N_3733);
or U4355 (N_4355,N_3658,N_3971);
nand U4356 (N_4356,N_3615,N_3996);
nand U4357 (N_4357,N_3678,N_3677);
and U4358 (N_4358,N_3757,N_3547);
nand U4359 (N_4359,N_3872,N_3641);
or U4360 (N_4360,N_3979,N_3780);
nand U4361 (N_4361,N_3808,N_3961);
and U4362 (N_4362,N_3971,N_3788);
nand U4363 (N_4363,N_3629,N_3736);
or U4364 (N_4364,N_3977,N_3678);
nand U4365 (N_4365,N_3599,N_3813);
nor U4366 (N_4366,N_3573,N_3832);
or U4367 (N_4367,N_3857,N_3738);
or U4368 (N_4368,N_3864,N_3537);
nand U4369 (N_4369,N_3733,N_3635);
nor U4370 (N_4370,N_3846,N_3520);
nand U4371 (N_4371,N_3521,N_3558);
and U4372 (N_4372,N_3888,N_3560);
and U4373 (N_4373,N_3865,N_3517);
and U4374 (N_4374,N_3763,N_3799);
xor U4375 (N_4375,N_3524,N_3946);
nand U4376 (N_4376,N_3767,N_3871);
and U4377 (N_4377,N_3569,N_3652);
and U4378 (N_4378,N_3800,N_3902);
nor U4379 (N_4379,N_3868,N_3848);
nand U4380 (N_4380,N_3750,N_3823);
and U4381 (N_4381,N_3972,N_3879);
nor U4382 (N_4382,N_3937,N_3577);
nor U4383 (N_4383,N_3629,N_3993);
and U4384 (N_4384,N_3695,N_3946);
or U4385 (N_4385,N_3656,N_3719);
nand U4386 (N_4386,N_3779,N_3817);
or U4387 (N_4387,N_3607,N_3943);
nor U4388 (N_4388,N_3945,N_3855);
nor U4389 (N_4389,N_3639,N_3869);
nand U4390 (N_4390,N_3801,N_3524);
nor U4391 (N_4391,N_3737,N_3822);
nor U4392 (N_4392,N_3735,N_3873);
nor U4393 (N_4393,N_3666,N_3657);
and U4394 (N_4394,N_3739,N_3922);
nand U4395 (N_4395,N_3887,N_3896);
nor U4396 (N_4396,N_3788,N_3976);
and U4397 (N_4397,N_3503,N_3629);
or U4398 (N_4398,N_3873,N_3737);
and U4399 (N_4399,N_3516,N_3540);
nand U4400 (N_4400,N_3917,N_3989);
and U4401 (N_4401,N_3873,N_3948);
nand U4402 (N_4402,N_3884,N_3914);
nand U4403 (N_4403,N_3620,N_3767);
nand U4404 (N_4404,N_3968,N_3915);
nand U4405 (N_4405,N_3555,N_3779);
and U4406 (N_4406,N_3953,N_3617);
or U4407 (N_4407,N_3564,N_3672);
nor U4408 (N_4408,N_3682,N_3738);
or U4409 (N_4409,N_3680,N_3756);
nor U4410 (N_4410,N_3575,N_3784);
or U4411 (N_4411,N_3849,N_3963);
nand U4412 (N_4412,N_3998,N_3806);
nand U4413 (N_4413,N_3671,N_3845);
xnor U4414 (N_4414,N_3715,N_3721);
nor U4415 (N_4415,N_3527,N_3901);
nand U4416 (N_4416,N_3919,N_3710);
or U4417 (N_4417,N_3796,N_3512);
and U4418 (N_4418,N_3993,N_3784);
nand U4419 (N_4419,N_3567,N_3960);
nand U4420 (N_4420,N_3870,N_3855);
or U4421 (N_4421,N_3518,N_3597);
nand U4422 (N_4422,N_3843,N_3948);
or U4423 (N_4423,N_3740,N_3648);
or U4424 (N_4424,N_3551,N_3901);
nor U4425 (N_4425,N_3502,N_3769);
nor U4426 (N_4426,N_3865,N_3919);
and U4427 (N_4427,N_3762,N_3593);
and U4428 (N_4428,N_3789,N_3973);
xor U4429 (N_4429,N_3532,N_3812);
or U4430 (N_4430,N_3750,N_3504);
nand U4431 (N_4431,N_3787,N_3880);
nor U4432 (N_4432,N_3835,N_3664);
and U4433 (N_4433,N_3826,N_3623);
or U4434 (N_4434,N_3954,N_3828);
or U4435 (N_4435,N_3967,N_3818);
and U4436 (N_4436,N_3610,N_3904);
xor U4437 (N_4437,N_3783,N_3548);
nor U4438 (N_4438,N_3770,N_3808);
nand U4439 (N_4439,N_3734,N_3895);
nor U4440 (N_4440,N_3681,N_3997);
xnor U4441 (N_4441,N_3983,N_3743);
and U4442 (N_4442,N_3980,N_3987);
nor U4443 (N_4443,N_3888,N_3723);
nor U4444 (N_4444,N_3849,N_3854);
and U4445 (N_4445,N_3964,N_3682);
or U4446 (N_4446,N_3676,N_3776);
nand U4447 (N_4447,N_3811,N_3563);
or U4448 (N_4448,N_3758,N_3916);
and U4449 (N_4449,N_3765,N_3610);
nand U4450 (N_4450,N_3701,N_3963);
nor U4451 (N_4451,N_3547,N_3561);
nand U4452 (N_4452,N_3503,N_3585);
nor U4453 (N_4453,N_3624,N_3972);
or U4454 (N_4454,N_3758,N_3692);
and U4455 (N_4455,N_3729,N_3630);
or U4456 (N_4456,N_3629,N_3517);
or U4457 (N_4457,N_3977,N_3711);
or U4458 (N_4458,N_3792,N_3562);
nand U4459 (N_4459,N_3984,N_3666);
nand U4460 (N_4460,N_3844,N_3919);
nand U4461 (N_4461,N_3968,N_3702);
nand U4462 (N_4462,N_3715,N_3714);
nor U4463 (N_4463,N_3651,N_3531);
nand U4464 (N_4464,N_3732,N_3812);
nand U4465 (N_4465,N_3500,N_3514);
nand U4466 (N_4466,N_3705,N_3799);
or U4467 (N_4467,N_3964,N_3620);
nor U4468 (N_4468,N_3855,N_3847);
nand U4469 (N_4469,N_3803,N_3807);
nor U4470 (N_4470,N_3864,N_3913);
and U4471 (N_4471,N_3943,N_3893);
nand U4472 (N_4472,N_3898,N_3928);
nor U4473 (N_4473,N_3828,N_3509);
or U4474 (N_4474,N_3658,N_3554);
and U4475 (N_4475,N_3937,N_3767);
nor U4476 (N_4476,N_3566,N_3755);
nor U4477 (N_4477,N_3942,N_3708);
nor U4478 (N_4478,N_3790,N_3678);
or U4479 (N_4479,N_3511,N_3684);
or U4480 (N_4480,N_3742,N_3905);
or U4481 (N_4481,N_3511,N_3549);
and U4482 (N_4482,N_3949,N_3552);
nor U4483 (N_4483,N_3735,N_3790);
nand U4484 (N_4484,N_3647,N_3736);
and U4485 (N_4485,N_3823,N_3642);
xnor U4486 (N_4486,N_3972,N_3724);
and U4487 (N_4487,N_3849,N_3807);
or U4488 (N_4488,N_3563,N_3630);
nor U4489 (N_4489,N_3698,N_3634);
and U4490 (N_4490,N_3908,N_3528);
and U4491 (N_4491,N_3993,N_3687);
xnor U4492 (N_4492,N_3548,N_3927);
or U4493 (N_4493,N_3802,N_3525);
nor U4494 (N_4494,N_3644,N_3552);
or U4495 (N_4495,N_3962,N_3975);
and U4496 (N_4496,N_3504,N_3547);
nand U4497 (N_4497,N_3620,N_3786);
nand U4498 (N_4498,N_3529,N_3658);
and U4499 (N_4499,N_3643,N_3909);
and U4500 (N_4500,N_4443,N_4007);
nor U4501 (N_4501,N_4215,N_4413);
nand U4502 (N_4502,N_4161,N_4323);
and U4503 (N_4503,N_4091,N_4481);
nand U4504 (N_4504,N_4005,N_4027);
or U4505 (N_4505,N_4442,N_4146);
nor U4506 (N_4506,N_4054,N_4402);
nor U4507 (N_4507,N_4259,N_4378);
nor U4508 (N_4508,N_4181,N_4238);
nor U4509 (N_4509,N_4368,N_4468);
or U4510 (N_4510,N_4486,N_4334);
and U4511 (N_4511,N_4319,N_4218);
or U4512 (N_4512,N_4429,N_4423);
and U4513 (N_4513,N_4278,N_4120);
and U4514 (N_4514,N_4310,N_4361);
or U4515 (N_4515,N_4052,N_4014);
or U4516 (N_4516,N_4456,N_4381);
or U4517 (N_4517,N_4089,N_4153);
or U4518 (N_4518,N_4158,N_4465);
nor U4519 (N_4519,N_4197,N_4366);
nand U4520 (N_4520,N_4239,N_4017);
nand U4521 (N_4521,N_4093,N_4096);
nand U4522 (N_4522,N_4241,N_4204);
nand U4523 (N_4523,N_4471,N_4225);
xor U4524 (N_4524,N_4491,N_4011);
nor U4525 (N_4525,N_4316,N_4437);
and U4526 (N_4526,N_4286,N_4212);
or U4527 (N_4527,N_4490,N_4026);
and U4528 (N_4528,N_4336,N_4352);
and U4529 (N_4529,N_4305,N_4317);
nor U4530 (N_4530,N_4045,N_4388);
or U4531 (N_4531,N_4010,N_4337);
or U4532 (N_4532,N_4015,N_4495);
nor U4533 (N_4533,N_4119,N_4099);
or U4534 (N_4534,N_4331,N_4249);
nor U4535 (N_4535,N_4482,N_4136);
and U4536 (N_4536,N_4232,N_4357);
and U4537 (N_4537,N_4433,N_4302);
nor U4538 (N_4538,N_4447,N_4365);
nand U4539 (N_4539,N_4375,N_4090);
nand U4540 (N_4540,N_4285,N_4419);
and U4541 (N_4541,N_4198,N_4424);
nand U4542 (N_4542,N_4410,N_4455);
nor U4543 (N_4543,N_4369,N_4343);
nor U4544 (N_4544,N_4408,N_4039);
or U4545 (N_4545,N_4248,N_4370);
nand U4546 (N_4546,N_4494,N_4498);
or U4547 (N_4547,N_4290,N_4418);
or U4548 (N_4548,N_4002,N_4301);
nor U4549 (N_4549,N_4036,N_4349);
nor U4550 (N_4550,N_4012,N_4013);
nor U4551 (N_4551,N_4439,N_4115);
xor U4552 (N_4552,N_4327,N_4462);
nand U4553 (N_4553,N_4004,N_4463);
or U4554 (N_4554,N_4214,N_4438);
nand U4555 (N_4555,N_4194,N_4195);
nor U4556 (N_4556,N_4492,N_4441);
nor U4557 (N_4557,N_4143,N_4114);
nor U4558 (N_4558,N_4269,N_4001);
nand U4559 (N_4559,N_4294,N_4245);
and U4560 (N_4560,N_4071,N_4341);
nor U4561 (N_4561,N_4458,N_4333);
and U4562 (N_4562,N_4080,N_4309);
or U4563 (N_4563,N_4038,N_4450);
nor U4564 (N_4564,N_4461,N_4340);
nand U4565 (N_4565,N_4281,N_4129);
nand U4566 (N_4566,N_4395,N_4379);
and U4567 (N_4567,N_4076,N_4100);
and U4568 (N_4568,N_4047,N_4466);
nor U4569 (N_4569,N_4344,N_4237);
nand U4570 (N_4570,N_4354,N_4289);
nand U4571 (N_4571,N_4219,N_4131);
or U4572 (N_4572,N_4191,N_4164);
nor U4573 (N_4573,N_4411,N_4396);
xnor U4574 (N_4574,N_4072,N_4168);
nand U4575 (N_4575,N_4306,N_4148);
and U4576 (N_4576,N_4020,N_4185);
and U4577 (N_4577,N_4223,N_4454);
or U4578 (N_4578,N_4162,N_4489);
nand U4579 (N_4579,N_4431,N_4170);
and U4580 (N_4580,N_4347,N_4070);
and U4581 (N_4581,N_4151,N_4280);
nand U4582 (N_4582,N_4044,N_4417);
nor U4583 (N_4583,N_4311,N_4243);
or U4584 (N_4584,N_4404,N_4128);
nand U4585 (N_4585,N_4159,N_4430);
nor U4586 (N_4586,N_4085,N_4130);
nor U4587 (N_4587,N_4200,N_4444);
or U4588 (N_4588,N_4043,N_4042);
and U4589 (N_4589,N_4307,N_4029);
nor U4590 (N_4590,N_4160,N_4426);
nand U4591 (N_4591,N_4380,N_4371);
nor U4592 (N_4592,N_4264,N_4436);
or U4593 (N_4593,N_4165,N_4066);
and U4594 (N_4594,N_4457,N_4116);
nand U4595 (N_4595,N_4152,N_4324);
and U4596 (N_4596,N_4171,N_4113);
or U4597 (N_4597,N_4183,N_4332);
nand U4598 (N_4598,N_4288,N_4094);
nor U4599 (N_4599,N_4067,N_4390);
nor U4600 (N_4600,N_4263,N_4240);
nand U4601 (N_4601,N_4435,N_4321);
nor U4602 (N_4602,N_4300,N_4303);
nor U4603 (N_4603,N_4377,N_4355);
nand U4604 (N_4604,N_4033,N_4261);
and U4605 (N_4605,N_4330,N_4393);
and U4606 (N_4606,N_4421,N_4068);
nor U4607 (N_4607,N_4470,N_4220);
or U4608 (N_4608,N_4206,N_4253);
nor U4609 (N_4609,N_4174,N_4273);
or U4610 (N_4610,N_4107,N_4325);
nor U4611 (N_4611,N_4422,N_4267);
or U4612 (N_4612,N_4078,N_4359);
and U4613 (N_4613,N_4226,N_4022);
or U4614 (N_4614,N_4362,N_4252);
and U4615 (N_4615,N_4360,N_4057);
and U4616 (N_4616,N_4414,N_4477);
nand U4617 (N_4617,N_4497,N_4084);
and U4618 (N_4618,N_4265,N_4081);
nand U4619 (N_4619,N_4405,N_4231);
nor U4620 (N_4620,N_4192,N_4193);
nand U4621 (N_4621,N_4060,N_4478);
nand U4622 (N_4622,N_4222,N_4299);
xnor U4623 (N_4623,N_4182,N_4098);
and U4624 (N_4624,N_4363,N_4262);
nand U4625 (N_4625,N_4139,N_4127);
nand U4626 (N_4626,N_4480,N_4034);
or U4627 (N_4627,N_4254,N_4079);
and U4628 (N_4628,N_4035,N_4075);
and U4629 (N_4629,N_4172,N_4040);
nor U4630 (N_4630,N_4025,N_4287);
nand U4631 (N_4631,N_4399,N_4415);
and U4632 (N_4632,N_4266,N_4485);
nand U4633 (N_4633,N_4353,N_4228);
and U4634 (N_4634,N_4432,N_4157);
and U4635 (N_4635,N_4207,N_4112);
xnor U4636 (N_4636,N_4208,N_4135);
and U4637 (N_4637,N_4268,N_4169);
and U4638 (N_4638,N_4202,N_4367);
nand U4639 (N_4639,N_4235,N_4297);
nor U4640 (N_4640,N_4484,N_4211);
and U4641 (N_4641,N_4190,N_4255);
and U4642 (N_4642,N_4087,N_4213);
or U4643 (N_4643,N_4082,N_4279);
nor U4644 (N_4644,N_4346,N_4106);
or U4645 (N_4645,N_4217,N_4083);
and U4646 (N_4646,N_4257,N_4406);
or U4647 (N_4647,N_4053,N_4453);
or U4648 (N_4648,N_4448,N_4137);
or U4649 (N_4649,N_4400,N_4451);
and U4650 (N_4650,N_4144,N_4282);
and U4651 (N_4651,N_4440,N_4474);
and U4652 (N_4652,N_4251,N_4108);
and U4653 (N_4653,N_4296,N_4175);
xor U4654 (N_4654,N_4409,N_4372);
or U4655 (N_4655,N_4356,N_4102);
nor U4656 (N_4656,N_4224,N_4187);
nor U4657 (N_4657,N_4304,N_4059);
and U4658 (N_4658,N_4358,N_4063);
or U4659 (N_4659,N_4348,N_4184);
or U4660 (N_4660,N_4003,N_4322);
nand U4661 (N_4661,N_4061,N_4313);
and U4662 (N_4662,N_4389,N_4350);
nor U4663 (N_4663,N_4140,N_4064);
nor U4664 (N_4664,N_4205,N_4420);
nand U4665 (N_4665,N_4101,N_4464);
nand U4666 (N_4666,N_4074,N_4176);
or U4667 (N_4667,N_4167,N_4121);
nand U4668 (N_4668,N_4046,N_4021);
or U4669 (N_4669,N_4401,N_4385);
nor U4670 (N_4670,N_4156,N_4318);
and U4671 (N_4671,N_4446,N_4242);
nor U4672 (N_4672,N_4229,N_4284);
nor U4673 (N_4673,N_4086,N_4326);
nand U4674 (N_4674,N_4339,N_4308);
nor U4675 (N_4675,N_4221,N_4179);
nand U4676 (N_4676,N_4077,N_4111);
or U4677 (N_4677,N_4145,N_4428);
or U4678 (N_4678,N_4293,N_4479);
or U4679 (N_4679,N_4103,N_4459);
nand U4680 (N_4680,N_4382,N_4342);
nor U4681 (N_4681,N_4178,N_4016);
or U4682 (N_4682,N_4298,N_4030);
or U4683 (N_4683,N_4291,N_4397);
and U4684 (N_4684,N_4493,N_4351);
or U4685 (N_4685,N_4199,N_4449);
or U4686 (N_4686,N_4201,N_4391);
nor U4687 (N_4687,N_4260,N_4155);
nand U4688 (N_4688,N_4234,N_4233);
nand U4689 (N_4689,N_4122,N_4270);
or U4690 (N_4690,N_4006,N_4376);
or U4691 (N_4691,N_4150,N_4024);
and U4692 (N_4692,N_4055,N_4472);
nand U4693 (N_4693,N_4188,N_4277);
or U4694 (N_4694,N_4018,N_4345);
nor U4695 (N_4695,N_4227,N_4275);
or U4696 (N_4696,N_4475,N_4216);
or U4697 (N_4697,N_4123,N_4283);
nor U4698 (N_4698,N_4032,N_4488);
nand U4699 (N_4699,N_4460,N_4434);
xor U4700 (N_4700,N_4445,N_4019);
nor U4701 (N_4701,N_4403,N_4088);
nand U4702 (N_4702,N_4487,N_4117);
or U4703 (N_4703,N_4023,N_4364);
or U4704 (N_4704,N_4320,N_4166);
nand U4705 (N_4705,N_4095,N_4118);
nor U4706 (N_4706,N_4271,N_4250);
nor U4707 (N_4707,N_4452,N_4392);
and U4708 (N_4708,N_4209,N_4110);
or U4709 (N_4709,N_4163,N_4050);
nor U4710 (N_4710,N_4272,N_4028);
nor U4711 (N_4711,N_4138,N_4000);
nor U4712 (N_4712,N_4469,N_4314);
nand U4713 (N_4713,N_4180,N_4008);
nand U4714 (N_4714,N_4186,N_4274);
xor U4715 (N_4715,N_4189,N_4483);
nand U4716 (N_4716,N_4105,N_4384);
nor U4717 (N_4717,N_4246,N_4173);
nand U4718 (N_4718,N_4387,N_4467);
and U4719 (N_4719,N_4276,N_4125);
and U4720 (N_4720,N_4412,N_4329);
nor U4721 (N_4721,N_4132,N_4048);
or U4722 (N_4722,N_4009,N_4258);
or U4723 (N_4723,N_4065,N_4092);
and U4724 (N_4724,N_4154,N_4338);
and U4725 (N_4725,N_4407,N_4499);
or U4726 (N_4726,N_4058,N_4425);
and U4727 (N_4727,N_4124,N_4315);
and U4728 (N_4728,N_4037,N_4386);
or U4729 (N_4729,N_4373,N_4398);
or U4730 (N_4730,N_4051,N_4416);
or U4731 (N_4731,N_4177,N_4335);
or U4732 (N_4732,N_4210,N_4049);
and U4733 (N_4733,N_4247,N_4383);
nor U4734 (N_4734,N_4141,N_4196);
nor U4735 (N_4735,N_4133,N_4097);
or U4736 (N_4736,N_4109,N_4236);
nand U4737 (N_4737,N_4295,N_4041);
nor U4738 (N_4738,N_4031,N_4147);
nor U4739 (N_4739,N_4073,N_4056);
nor U4740 (N_4740,N_4230,N_4069);
and U4741 (N_4741,N_4473,N_4134);
nor U4742 (N_4742,N_4374,N_4244);
nand U4743 (N_4743,N_4427,N_4256);
and U4744 (N_4744,N_4142,N_4476);
nand U4745 (N_4745,N_4394,N_4104);
nor U4746 (N_4746,N_4328,N_4312);
nand U4747 (N_4747,N_4496,N_4203);
and U4748 (N_4748,N_4292,N_4062);
nand U4749 (N_4749,N_4126,N_4149);
and U4750 (N_4750,N_4185,N_4076);
or U4751 (N_4751,N_4222,N_4115);
or U4752 (N_4752,N_4350,N_4280);
nand U4753 (N_4753,N_4334,N_4181);
or U4754 (N_4754,N_4337,N_4174);
nor U4755 (N_4755,N_4200,N_4265);
nand U4756 (N_4756,N_4402,N_4130);
and U4757 (N_4757,N_4085,N_4093);
nor U4758 (N_4758,N_4348,N_4325);
or U4759 (N_4759,N_4434,N_4055);
and U4760 (N_4760,N_4071,N_4284);
nor U4761 (N_4761,N_4267,N_4044);
nand U4762 (N_4762,N_4166,N_4343);
or U4763 (N_4763,N_4382,N_4200);
nand U4764 (N_4764,N_4006,N_4009);
nand U4765 (N_4765,N_4459,N_4380);
or U4766 (N_4766,N_4423,N_4133);
xor U4767 (N_4767,N_4062,N_4246);
nand U4768 (N_4768,N_4072,N_4036);
nand U4769 (N_4769,N_4332,N_4077);
and U4770 (N_4770,N_4339,N_4215);
xor U4771 (N_4771,N_4158,N_4369);
and U4772 (N_4772,N_4050,N_4086);
or U4773 (N_4773,N_4441,N_4216);
or U4774 (N_4774,N_4460,N_4375);
nor U4775 (N_4775,N_4049,N_4175);
and U4776 (N_4776,N_4302,N_4329);
or U4777 (N_4777,N_4266,N_4176);
and U4778 (N_4778,N_4406,N_4255);
nor U4779 (N_4779,N_4456,N_4429);
nand U4780 (N_4780,N_4256,N_4060);
and U4781 (N_4781,N_4307,N_4453);
or U4782 (N_4782,N_4157,N_4470);
nand U4783 (N_4783,N_4189,N_4304);
nand U4784 (N_4784,N_4453,N_4352);
nand U4785 (N_4785,N_4396,N_4273);
nor U4786 (N_4786,N_4214,N_4446);
nor U4787 (N_4787,N_4423,N_4255);
and U4788 (N_4788,N_4333,N_4496);
nor U4789 (N_4789,N_4395,N_4064);
nor U4790 (N_4790,N_4291,N_4119);
nor U4791 (N_4791,N_4493,N_4482);
and U4792 (N_4792,N_4474,N_4205);
nor U4793 (N_4793,N_4360,N_4306);
and U4794 (N_4794,N_4329,N_4130);
or U4795 (N_4795,N_4315,N_4298);
and U4796 (N_4796,N_4095,N_4322);
nand U4797 (N_4797,N_4201,N_4222);
xor U4798 (N_4798,N_4132,N_4180);
nand U4799 (N_4799,N_4253,N_4458);
nor U4800 (N_4800,N_4484,N_4075);
or U4801 (N_4801,N_4462,N_4084);
nor U4802 (N_4802,N_4464,N_4229);
nor U4803 (N_4803,N_4255,N_4198);
nor U4804 (N_4804,N_4294,N_4306);
and U4805 (N_4805,N_4395,N_4080);
nor U4806 (N_4806,N_4419,N_4261);
nor U4807 (N_4807,N_4383,N_4424);
nand U4808 (N_4808,N_4291,N_4123);
nand U4809 (N_4809,N_4068,N_4459);
or U4810 (N_4810,N_4072,N_4181);
and U4811 (N_4811,N_4235,N_4090);
and U4812 (N_4812,N_4272,N_4030);
or U4813 (N_4813,N_4367,N_4155);
nand U4814 (N_4814,N_4482,N_4146);
or U4815 (N_4815,N_4102,N_4340);
nand U4816 (N_4816,N_4096,N_4421);
nand U4817 (N_4817,N_4361,N_4379);
nand U4818 (N_4818,N_4158,N_4146);
nand U4819 (N_4819,N_4491,N_4388);
nand U4820 (N_4820,N_4212,N_4025);
and U4821 (N_4821,N_4051,N_4012);
nand U4822 (N_4822,N_4471,N_4196);
or U4823 (N_4823,N_4194,N_4066);
nor U4824 (N_4824,N_4380,N_4048);
nand U4825 (N_4825,N_4239,N_4140);
or U4826 (N_4826,N_4109,N_4077);
nor U4827 (N_4827,N_4024,N_4175);
nand U4828 (N_4828,N_4194,N_4485);
nor U4829 (N_4829,N_4117,N_4114);
nor U4830 (N_4830,N_4106,N_4188);
nor U4831 (N_4831,N_4184,N_4361);
or U4832 (N_4832,N_4128,N_4449);
nor U4833 (N_4833,N_4440,N_4281);
xnor U4834 (N_4834,N_4200,N_4297);
or U4835 (N_4835,N_4415,N_4067);
and U4836 (N_4836,N_4306,N_4273);
and U4837 (N_4837,N_4131,N_4416);
nand U4838 (N_4838,N_4392,N_4358);
nand U4839 (N_4839,N_4052,N_4149);
and U4840 (N_4840,N_4156,N_4419);
nor U4841 (N_4841,N_4326,N_4291);
nand U4842 (N_4842,N_4139,N_4447);
xor U4843 (N_4843,N_4055,N_4368);
nor U4844 (N_4844,N_4133,N_4477);
nand U4845 (N_4845,N_4141,N_4025);
and U4846 (N_4846,N_4148,N_4192);
and U4847 (N_4847,N_4082,N_4050);
or U4848 (N_4848,N_4166,N_4353);
and U4849 (N_4849,N_4482,N_4117);
or U4850 (N_4850,N_4279,N_4046);
nor U4851 (N_4851,N_4277,N_4316);
or U4852 (N_4852,N_4254,N_4048);
nand U4853 (N_4853,N_4244,N_4354);
nor U4854 (N_4854,N_4029,N_4296);
nand U4855 (N_4855,N_4449,N_4197);
nor U4856 (N_4856,N_4367,N_4377);
nand U4857 (N_4857,N_4163,N_4228);
nand U4858 (N_4858,N_4157,N_4134);
or U4859 (N_4859,N_4382,N_4384);
nand U4860 (N_4860,N_4419,N_4153);
or U4861 (N_4861,N_4388,N_4449);
nand U4862 (N_4862,N_4258,N_4065);
nor U4863 (N_4863,N_4251,N_4481);
or U4864 (N_4864,N_4030,N_4125);
nand U4865 (N_4865,N_4024,N_4087);
and U4866 (N_4866,N_4312,N_4024);
and U4867 (N_4867,N_4158,N_4301);
and U4868 (N_4868,N_4110,N_4313);
nand U4869 (N_4869,N_4031,N_4397);
nor U4870 (N_4870,N_4143,N_4445);
nand U4871 (N_4871,N_4222,N_4282);
nand U4872 (N_4872,N_4019,N_4217);
or U4873 (N_4873,N_4275,N_4265);
or U4874 (N_4874,N_4025,N_4356);
and U4875 (N_4875,N_4332,N_4373);
nand U4876 (N_4876,N_4362,N_4083);
and U4877 (N_4877,N_4218,N_4159);
or U4878 (N_4878,N_4332,N_4010);
and U4879 (N_4879,N_4091,N_4338);
nor U4880 (N_4880,N_4168,N_4050);
or U4881 (N_4881,N_4312,N_4323);
nand U4882 (N_4882,N_4423,N_4158);
or U4883 (N_4883,N_4410,N_4385);
nand U4884 (N_4884,N_4485,N_4222);
and U4885 (N_4885,N_4498,N_4163);
nor U4886 (N_4886,N_4339,N_4319);
nand U4887 (N_4887,N_4185,N_4434);
and U4888 (N_4888,N_4193,N_4167);
and U4889 (N_4889,N_4263,N_4246);
nor U4890 (N_4890,N_4391,N_4347);
nand U4891 (N_4891,N_4117,N_4288);
nand U4892 (N_4892,N_4486,N_4386);
and U4893 (N_4893,N_4257,N_4006);
nor U4894 (N_4894,N_4394,N_4177);
nor U4895 (N_4895,N_4456,N_4461);
nor U4896 (N_4896,N_4248,N_4153);
xnor U4897 (N_4897,N_4453,N_4173);
and U4898 (N_4898,N_4356,N_4208);
or U4899 (N_4899,N_4376,N_4412);
or U4900 (N_4900,N_4196,N_4383);
and U4901 (N_4901,N_4398,N_4428);
nand U4902 (N_4902,N_4343,N_4314);
and U4903 (N_4903,N_4306,N_4302);
xor U4904 (N_4904,N_4064,N_4050);
and U4905 (N_4905,N_4173,N_4118);
nor U4906 (N_4906,N_4166,N_4107);
or U4907 (N_4907,N_4492,N_4283);
and U4908 (N_4908,N_4167,N_4217);
and U4909 (N_4909,N_4229,N_4067);
nor U4910 (N_4910,N_4464,N_4343);
or U4911 (N_4911,N_4329,N_4177);
and U4912 (N_4912,N_4048,N_4467);
nand U4913 (N_4913,N_4235,N_4134);
or U4914 (N_4914,N_4405,N_4226);
nand U4915 (N_4915,N_4153,N_4377);
or U4916 (N_4916,N_4325,N_4152);
nor U4917 (N_4917,N_4194,N_4218);
and U4918 (N_4918,N_4261,N_4327);
xnor U4919 (N_4919,N_4116,N_4232);
nand U4920 (N_4920,N_4313,N_4184);
and U4921 (N_4921,N_4326,N_4188);
nor U4922 (N_4922,N_4322,N_4383);
nor U4923 (N_4923,N_4146,N_4249);
nand U4924 (N_4924,N_4274,N_4479);
and U4925 (N_4925,N_4169,N_4316);
and U4926 (N_4926,N_4134,N_4472);
nor U4927 (N_4927,N_4402,N_4034);
nand U4928 (N_4928,N_4481,N_4488);
nand U4929 (N_4929,N_4016,N_4127);
nor U4930 (N_4930,N_4243,N_4472);
nor U4931 (N_4931,N_4433,N_4446);
nand U4932 (N_4932,N_4440,N_4167);
nor U4933 (N_4933,N_4337,N_4481);
nor U4934 (N_4934,N_4027,N_4242);
nand U4935 (N_4935,N_4205,N_4344);
and U4936 (N_4936,N_4289,N_4255);
or U4937 (N_4937,N_4436,N_4340);
and U4938 (N_4938,N_4311,N_4269);
nand U4939 (N_4939,N_4051,N_4350);
or U4940 (N_4940,N_4199,N_4050);
nand U4941 (N_4941,N_4007,N_4102);
and U4942 (N_4942,N_4071,N_4427);
nor U4943 (N_4943,N_4348,N_4317);
and U4944 (N_4944,N_4434,N_4294);
or U4945 (N_4945,N_4219,N_4416);
nand U4946 (N_4946,N_4283,N_4479);
or U4947 (N_4947,N_4061,N_4004);
nor U4948 (N_4948,N_4294,N_4264);
nand U4949 (N_4949,N_4006,N_4390);
and U4950 (N_4950,N_4395,N_4493);
nor U4951 (N_4951,N_4102,N_4234);
and U4952 (N_4952,N_4000,N_4226);
nand U4953 (N_4953,N_4135,N_4214);
and U4954 (N_4954,N_4194,N_4263);
and U4955 (N_4955,N_4377,N_4045);
nor U4956 (N_4956,N_4230,N_4006);
or U4957 (N_4957,N_4481,N_4472);
or U4958 (N_4958,N_4381,N_4026);
or U4959 (N_4959,N_4206,N_4314);
and U4960 (N_4960,N_4366,N_4331);
nand U4961 (N_4961,N_4191,N_4202);
or U4962 (N_4962,N_4293,N_4167);
nand U4963 (N_4963,N_4143,N_4193);
or U4964 (N_4964,N_4499,N_4205);
xor U4965 (N_4965,N_4285,N_4353);
nor U4966 (N_4966,N_4326,N_4126);
and U4967 (N_4967,N_4472,N_4207);
nand U4968 (N_4968,N_4320,N_4200);
xor U4969 (N_4969,N_4177,N_4398);
and U4970 (N_4970,N_4274,N_4280);
and U4971 (N_4971,N_4295,N_4398);
and U4972 (N_4972,N_4079,N_4080);
xor U4973 (N_4973,N_4142,N_4314);
and U4974 (N_4974,N_4120,N_4039);
or U4975 (N_4975,N_4392,N_4136);
and U4976 (N_4976,N_4234,N_4124);
or U4977 (N_4977,N_4139,N_4343);
nand U4978 (N_4978,N_4164,N_4157);
nand U4979 (N_4979,N_4458,N_4126);
or U4980 (N_4980,N_4163,N_4457);
and U4981 (N_4981,N_4235,N_4382);
nand U4982 (N_4982,N_4158,N_4175);
or U4983 (N_4983,N_4473,N_4276);
or U4984 (N_4984,N_4430,N_4047);
nand U4985 (N_4985,N_4413,N_4203);
nand U4986 (N_4986,N_4405,N_4196);
or U4987 (N_4987,N_4477,N_4209);
nor U4988 (N_4988,N_4027,N_4049);
or U4989 (N_4989,N_4081,N_4217);
nand U4990 (N_4990,N_4374,N_4441);
or U4991 (N_4991,N_4045,N_4199);
nor U4992 (N_4992,N_4251,N_4087);
and U4993 (N_4993,N_4152,N_4239);
and U4994 (N_4994,N_4332,N_4293);
nand U4995 (N_4995,N_4494,N_4112);
and U4996 (N_4996,N_4433,N_4314);
and U4997 (N_4997,N_4406,N_4178);
nor U4998 (N_4998,N_4326,N_4299);
or U4999 (N_4999,N_4451,N_4260);
nand UO_0 (O_0,N_4719,N_4822);
or UO_1 (O_1,N_4895,N_4912);
nand UO_2 (O_2,N_4825,N_4990);
or UO_3 (O_3,N_4622,N_4562);
or UO_4 (O_4,N_4801,N_4734);
or UO_5 (O_5,N_4699,N_4884);
and UO_6 (O_6,N_4978,N_4854);
or UO_7 (O_7,N_4867,N_4810);
or UO_8 (O_8,N_4824,N_4977);
and UO_9 (O_9,N_4539,N_4563);
nand UO_10 (O_10,N_4740,N_4842);
or UO_11 (O_11,N_4905,N_4812);
nor UO_12 (O_12,N_4580,N_4898);
nand UO_13 (O_13,N_4526,N_4722);
or UO_14 (O_14,N_4676,N_4733);
nand UO_15 (O_15,N_4889,N_4806);
or UO_16 (O_16,N_4992,N_4883);
and UO_17 (O_17,N_4590,N_4642);
or UO_18 (O_18,N_4843,N_4512);
nor UO_19 (O_19,N_4848,N_4829);
nor UO_20 (O_20,N_4773,N_4947);
and UO_21 (O_21,N_4763,N_4881);
xor UO_22 (O_22,N_4805,N_4823);
or UO_23 (O_23,N_4581,N_4543);
or UO_24 (O_24,N_4891,N_4717);
and UO_25 (O_25,N_4983,N_4863);
and UO_26 (O_26,N_4568,N_4885);
nor UO_27 (O_27,N_4862,N_4737);
nor UO_28 (O_28,N_4944,N_4841);
nor UO_29 (O_29,N_4925,N_4815);
nor UO_30 (O_30,N_4633,N_4922);
and UO_31 (O_31,N_4711,N_4975);
xor UO_32 (O_32,N_4914,N_4900);
xor UO_33 (O_33,N_4954,N_4890);
nand UO_34 (O_34,N_4816,N_4538);
nor UO_35 (O_35,N_4830,N_4675);
or UO_36 (O_36,N_4566,N_4820);
nor UO_37 (O_37,N_4686,N_4533);
or UO_38 (O_38,N_4764,N_4521);
nand UO_39 (O_39,N_4915,N_4778);
or UO_40 (O_40,N_4859,N_4638);
nor UO_41 (O_41,N_4772,N_4594);
nand UO_42 (O_42,N_4652,N_4794);
and UO_43 (O_43,N_4808,N_4786);
nand UO_44 (O_44,N_4523,N_4920);
or UO_45 (O_45,N_4952,N_4597);
nand UO_46 (O_46,N_4760,N_4758);
and UO_47 (O_47,N_4720,N_4860);
or UO_48 (O_48,N_4683,N_4766);
nand UO_49 (O_49,N_4588,N_4958);
or UO_50 (O_50,N_4714,N_4565);
nand UO_51 (O_51,N_4853,N_4871);
nand UO_52 (O_52,N_4716,N_4630);
nand UO_53 (O_53,N_4564,N_4991);
nor UO_54 (O_54,N_4660,N_4602);
nand UO_55 (O_55,N_4583,N_4902);
nand UO_56 (O_56,N_4743,N_4636);
or UO_57 (O_57,N_4657,N_4706);
nor UO_58 (O_58,N_4738,N_4730);
nand UO_59 (O_59,N_4577,N_4600);
nor UO_60 (O_60,N_4641,N_4570);
nand UO_61 (O_61,N_4963,N_4554);
or UO_62 (O_62,N_4851,N_4504);
or UO_63 (O_63,N_4974,N_4864);
or UO_64 (O_64,N_4695,N_4627);
nor UO_65 (O_65,N_4544,N_4793);
nand UO_66 (O_66,N_4712,N_4585);
xor UO_67 (O_67,N_4846,N_4610);
or UO_68 (O_68,N_4725,N_4668);
and UO_69 (O_69,N_4769,N_4771);
or UO_70 (O_70,N_4670,N_4671);
nand UO_71 (O_71,N_4751,N_4833);
and UO_72 (O_72,N_4656,N_4537);
nand UO_73 (O_73,N_4531,N_4752);
and UO_74 (O_74,N_4798,N_4673);
nor UO_75 (O_75,N_4755,N_4803);
nor UO_76 (O_76,N_4746,N_4721);
nand UO_77 (O_77,N_4741,N_4972);
and UO_78 (O_78,N_4887,N_4785);
nor UO_79 (O_79,N_4831,N_4948);
nor UO_80 (O_80,N_4913,N_4774);
or UO_81 (O_81,N_4731,N_4888);
nand UO_82 (O_82,N_4994,N_4744);
nand UO_83 (O_83,N_4651,N_4770);
and UO_84 (O_84,N_4524,N_4945);
nor UO_85 (O_85,N_4874,N_4965);
nor UO_86 (O_86,N_4503,N_4908);
nand UO_87 (O_87,N_4688,N_4507);
or UO_88 (O_88,N_4886,N_4858);
nor UO_89 (O_89,N_4736,N_4964);
or UO_90 (O_90,N_4684,N_4513);
nand UO_91 (O_91,N_4742,N_4586);
nor UO_92 (O_92,N_4873,N_4916);
xnor UO_93 (O_93,N_4946,N_4931);
nand UO_94 (O_94,N_4781,N_4800);
or UO_95 (O_95,N_4637,N_4957);
xnor UO_96 (O_96,N_4601,N_4696);
and UO_97 (O_97,N_4909,N_4927);
nand UO_98 (O_98,N_4704,N_4687);
nor UO_99 (O_99,N_4937,N_4911);
nor UO_100 (O_100,N_4573,N_4611);
or UO_101 (O_101,N_4813,N_4852);
or UO_102 (O_102,N_4584,N_4579);
and UO_103 (O_103,N_4628,N_4951);
and UO_104 (O_104,N_4966,N_4664);
or UO_105 (O_105,N_4837,N_4708);
nor UO_106 (O_106,N_4532,N_4677);
and UO_107 (O_107,N_4819,N_4932);
or UO_108 (O_108,N_4828,N_4982);
and UO_109 (O_109,N_4817,N_4968);
and UO_110 (O_110,N_4669,N_4582);
and UO_111 (O_111,N_4614,N_4809);
nor UO_112 (O_112,N_4649,N_4861);
and UO_113 (O_113,N_4639,N_4545);
nor UO_114 (O_114,N_4762,N_4569);
and UO_115 (O_115,N_4949,N_4796);
nor UO_116 (O_116,N_4528,N_4757);
nand UO_117 (O_117,N_4718,N_4756);
nor UO_118 (O_118,N_4959,N_4882);
and UO_119 (O_119,N_4665,N_4950);
or UO_120 (O_120,N_4516,N_4571);
or UO_121 (O_121,N_4553,N_4645);
nand UO_122 (O_122,N_4595,N_4728);
and UO_123 (O_123,N_4971,N_4592);
or UO_124 (O_124,N_4655,N_4635);
and UO_125 (O_125,N_4542,N_4522);
nand UO_126 (O_126,N_4940,N_4783);
nor UO_127 (O_127,N_4697,N_4694);
nor UO_128 (O_128,N_4705,N_4702);
nor UO_129 (O_129,N_4558,N_4647);
nand UO_130 (O_130,N_4506,N_4779);
xor UO_131 (O_131,N_4835,N_4620);
and UO_132 (O_132,N_4901,N_4938);
and UO_133 (O_133,N_4799,N_4789);
nand UO_134 (O_134,N_4777,N_4899);
nand UO_135 (O_135,N_4698,N_4621);
nor UO_136 (O_136,N_4631,N_4682);
nor UO_137 (O_137,N_4608,N_4654);
or UO_138 (O_138,N_4605,N_4603);
and UO_139 (O_139,N_4967,N_4663);
nor UO_140 (O_140,N_4814,N_4985);
nor UO_141 (O_141,N_4818,N_4640);
or UO_142 (O_142,N_4729,N_4685);
or UO_143 (O_143,N_4976,N_4840);
nand UO_144 (O_144,N_4749,N_4501);
or UO_145 (O_145,N_4525,N_4609);
nor UO_146 (O_146,N_4917,N_4926);
and UO_147 (O_147,N_4626,N_4849);
nor UO_148 (O_148,N_4877,N_4561);
xor UO_149 (O_149,N_4678,N_4508);
nor UO_150 (O_150,N_4986,N_4759);
or UO_151 (O_151,N_4839,N_4904);
nand UO_152 (O_152,N_4981,N_4868);
and UO_153 (O_153,N_4987,N_4802);
and UO_154 (O_154,N_4768,N_4934);
or UO_155 (O_155,N_4907,N_4866);
nand UO_156 (O_156,N_4761,N_4879);
nand UO_157 (O_157,N_4845,N_4857);
nor UO_158 (O_158,N_4604,N_4739);
nor UO_159 (O_159,N_4693,N_4748);
and UO_160 (O_160,N_4807,N_4598);
nand UO_161 (O_161,N_4619,N_4500);
nand UO_162 (O_162,N_4962,N_4552);
nor UO_163 (O_163,N_4735,N_4661);
and UO_164 (O_164,N_4653,N_4776);
and UO_165 (O_165,N_4821,N_4546);
or UO_166 (O_166,N_4576,N_4921);
nand UO_167 (O_167,N_4790,N_4832);
nor UO_168 (O_168,N_4692,N_4617);
or UO_169 (O_169,N_4918,N_4935);
and UO_170 (O_170,N_4587,N_4502);
or UO_171 (O_171,N_4559,N_4615);
or UO_172 (O_172,N_4691,N_4509);
or UO_173 (O_173,N_4953,N_4681);
and UO_174 (O_174,N_4606,N_4551);
and UO_175 (O_175,N_4591,N_4529);
and UO_176 (O_176,N_4557,N_4984);
nand UO_177 (O_177,N_4672,N_4969);
and UO_178 (O_178,N_4658,N_4980);
nor UO_179 (O_179,N_4514,N_4910);
and UO_180 (O_180,N_4530,N_4903);
or UO_181 (O_181,N_4709,N_4575);
nand UO_182 (O_182,N_4765,N_4710);
or UO_183 (O_183,N_4690,N_4662);
nor UO_184 (O_184,N_4700,N_4650);
xnor UO_185 (O_185,N_4723,N_4973);
or UO_186 (O_186,N_4997,N_4795);
or UO_187 (O_187,N_4792,N_4750);
nor UO_188 (O_188,N_4701,N_4894);
nor UO_189 (O_189,N_4955,N_4939);
or UO_190 (O_190,N_4518,N_4574);
nand UO_191 (O_191,N_4724,N_4572);
nor UO_192 (O_192,N_4515,N_4811);
nor UO_193 (O_193,N_4775,N_4703);
or UO_194 (O_194,N_4989,N_4505);
nand UO_195 (O_195,N_4747,N_4791);
nand UO_196 (O_196,N_4726,N_4784);
or UO_197 (O_197,N_4780,N_4535);
nand UO_198 (O_198,N_4547,N_4782);
or UO_199 (O_199,N_4855,N_4593);
nor UO_200 (O_200,N_4875,N_4753);
nor UO_201 (O_201,N_4996,N_4827);
and UO_202 (O_202,N_4797,N_4616);
or UO_203 (O_203,N_4536,N_4897);
or UO_204 (O_204,N_4659,N_4589);
nor UO_205 (O_205,N_4517,N_4956);
xnor UO_206 (O_206,N_4998,N_4527);
nand UO_207 (O_207,N_4892,N_4667);
nor UO_208 (O_208,N_4826,N_4834);
nand UO_209 (O_209,N_4550,N_4713);
nand UO_210 (O_210,N_4836,N_4942);
or UO_211 (O_211,N_4995,N_4893);
nor UO_212 (O_212,N_4727,N_4560);
nand UO_213 (O_213,N_4767,N_4680);
nand UO_214 (O_214,N_4847,N_4648);
nor UO_215 (O_215,N_4936,N_4556);
nor UO_216 (O_216,N_4924,N_4856);
or UO_217 (O_217,N_4930,N_4555);
or UO_218 (O_218,N_4679,N_4634);
or UO_219 (O_219,N_4745,N_4754);
or UO_220 (O_220,N_4624,N_4567);
or UO_221 (O_221,N_4999,N_4850);
or UO_222 (O_222,N_4919,N_4979);
and UO_223 (O_223,N_4618,N_4596);
nand UO_224 (O_224,N_4844,N_4541);
nor UO_225 (O_225,N_4534,N_4804);
or UO_226 (O_226,N_4732,N_4715);
nor UO_227 (O_227,N_4943,N_4787);
nand UO_228 (O_228,N_4548,N_4788);
or UO_229 (O_229,N_4961,N_4880);
or UO_230 (O_230,N_4629,N_4578);
nand UO_231 (O_231,N_4906,N_4644);
or UO_232 (O_232,N_4933,N_4613);
and UO_233 (O_233,N_4549,N_4599);
or UO_234 (O_234,N_4865,N_4923);
nand UO_235 (O_235,N_4689,N_4941);
or UO_236 (O_236,N_4707,N_4878);
or UO_237 (O_237,N_4869,N_4607);
nand UO_238 (O_238,N_4988,N_4632);
nand UO_239 (O_239,N_4970,N_4625);
and UO_240 (O_240,N_4870,N_4666);
and UO_241 (O_241,N_4929,N_4872);
nor UO_242 (O_242,N_4674,N_4520);
or UO_243 (O_243,N_4646,N_4838);
nor UO_244 (O_244,N_4612,N_4993);
or UO_245 (O_245,N_4510,N_4896);
nand UO_246 (O_246,N_4643,N_4928);
nand UO_247 (O_247,N_4960,N_4540);
or UO_248 (O_248,N_4519,N_4876);
and UO_249 (O_249,N_4511,N_4623);
or UO_250 (O_250,N_4761,N_4958);
and UO_251 (O_251,N_4667,N_4995);
nand UO_252 (O_252,N_4775,N_4706);
and UO_253 (O_253,N_4587,N_4755);
and UO_254 (O_254,N_4686,N_4823);
nand UO_255 (O_255,N_4834,N_4627);
and UO_256 (O_256,N_4850,N_4510);
and UO_257 (O_257,N_4830,N_4502);
and UO_258 (O_258,N_4802,N_4871);
and UO_259 (O_259,N_4618,N_4630);
nor UO_260 (O_260,N_4844,N_4677);
and UO_261 (O_261,N_4551,N_4774);
nand UO_262 (O_262,N_4761,N_4875);
nand UO_263 (O_263,N_4963,N_4886);
nand UO_264 (O_264,N_4569,N_4604);
nand UO_265 (O_265,N_4825,N_4508);
nand UO_266 (O_266,N_4922,N_4771);
and UO_267 (O_267,N_4648,N_4949);
and UO_268 (O_268,N_4549,N_4670);
nand UO_269 (O_269,N_4808,N_4846);
and UO_270 (O_270,N_4798,N_4849);
or UO_271 (O_271,N_4759,N_4744);
nand UO_272 (O_272,N_4797,N_4883);
or UO_273 (O_273,N_4693,N_4861);
xor UO_274 (O_274,N_4914,N_4693);
or UO_275 (O_275,N_4811,N_4886);
xnor UO_276 (O_276,N_4855,N_4997);
nor UO_277 (O_277,N_4908,N_4753);
nor UO_278 (O_278,N_4530,N_4689);
xor UO_279 (O_279,N_4691,N_4972);
or UO_280 (O_280,N_4897,N_4984);
xnor UO_281 (O_281,N_4787,N_4605);
nand UO_282 (O_282,N_4604,N_4996);
or UO_283 (O_283,N_4880,N_4695);
or UO_284 (O_284,N_4501,N_4813);
and UO_285 (O_285,N_4760,N_4561);
nor UO_286 (O_286,N_4706,N_4694);
nor UO_287 (O_287,N_4929,N_4804);
nor UO_288 (O_288,N_4554,N_4875);
nor UO_289 (O_289,N_4956,N_4918);
xnor UO_290 (O_290,N_4954,N_4836);
nand UO_291 (O_291,N_4819,N_4940);
and UO_292 (O_292,N_4959,N_4510);
or UO_293 (O_293,N_4648,N_4597);
nand UO_294 (O_294,N_4865,N_4946);
and UO_295 (O_295,N_4971,N_4757);
nand UO_296 (O_296,N_4576,N_4825);
and UO_297 (O_297,N_4827,N_4591);
and UO_298 (O_298,N_4991,N_4662);
or UO_299 (O_299,N_4594,N_4662);
nor UO_300 (O_300,N_4993,N_4576);
nand UO_301 (O_301,N_4617,N_4777);
nor UO_302 (O_302,N_4952,N_4653);
or UO_303 (O_303,N_4882,N_4569);
xnor UO_304 (O_304,N_4925,N_4574);
and UO_305 (O_305,N_4802,N_4793);
or UO_306 (O_306,N_4642,N_4790);
or UO_307 (O_307,N_4618,N_4675);
or UO_308 (O_308,N_4737,N_4813);
nand UO_309 (O_309,N_4792,N_4781);
or UO_310 (O_310,N_4537,N_4578);
and UO_311 (O_311,N_4850,N_4957);
or UO_312 (O_312,N_4720,N_4512);
or UO_313 (O_313,N_4665,N_4931);
nor UO_314 (O_314,N_4978,N_4663);
nor UO_315 (O_315,N_4616,N_4780);
nor UO_316 (O_316,N_4735,N_4625);
or UO_317 (O_317,N_4913,N_4602);
or UO_318 (O_318,N_4637,N_4887);
nor UO_319 (O_319,N_4748,N_4904);
or UO_320 (O_320,N_4726,N_4689);
or UO_321 (O_321,N_4537,N_4911);
or UO_322 (O_322,N_4735,N_4972);
and UO_323 (O_323,N_4872,N_4975);
nand UO_324 (O_324,N_4707,N_4530);
and UO_325 (O_325,N_4891,N_4697);
nand UO_326 (O_326,N_4530,N_4879);
nor UO_327 (O_327,N_4781,N_4935);
and UO_328 (O_328,N_4581,N_4921);
and UO_329 (O_329,N_4921,N_4555);
or UO_330 (O_330,N_4629,N_4725);
or UO_331 (O_331,N_4586,N_4868);
and UO_332 (O_332,N_4574,N_4891);
nand UO_333 (O_333,N_4875,N_4572);
or UO_334 (O_334,N_4541,N_4552);
nor UO_335 (O_335,N_4916,N_4882);
and UO_336 (O_336,N_4640,N_4678);
nor UO_337 (O_337,N_4604,N_4925);
or UO_338 (O_338,N_4691,N_4526);
or UO_339 (O_339,N_4551,N_4972);
nand UO_340 (O_340,N_4611,N_4524);
nor UO_341 (O_341,N_4653,N_4548);
nand UO_342 (O_342,N_4922,N_4876);
nand UO_343 (O_343,N_4640,N_4841);
and UO_344 (O_344,N_4658,N_4933);
or UO_345 (O_345,N_4939,N_4682);
and UO_346 (O_346,N_4969,N_4747);
or UO_347 (O_347,N_4992,N_4743);
or UO_348 (O_348,N_4629,N_4561);
and UO_349 (O_349,N_4814,N_4578);
and UO_350 (O_350,N_4877,N_4797);
nand UO_351 (O_351,N_4701,N_4997);
or UO_352 (O_352,N_4872,N_4697);
or UO_353 (O_353,N_4745,N_4699);
and UO_354 (O_354,N_4791,N_4524);
nand UO_355 (O_355,N_4541,N_4625);
and UO_356 (O_356,N_4651,N_4510);
nand UO_357 (O_357,N_4940,N_4510);
xnor UO_358 (O_358,N_4695,N_4564);
nand UO_359 (O_359,N_4523,N_4661);
and UO_360 (O_360,N_4965,N_4716);
nand UO_361 (O_361,N_4734,N_4709);
or UO_362 (O_362,N_4936,N_4928);
or UO_363 (O_363,N_4903,N_4861);
and UO_364 (O_364,N_4553,N_4811);
and UO_365 (O_365,N_4761,N_4977);
nor UO_366 (O_366,N_4675,N_4508);
or UO_367 (O_367,N_4672,N_4718);
or UO_368 (O_368,N_4855,N_4786);
nor UO_369 (O_369,N_4725,N_4926);
or UO_370 (O_370,N_4880,N_4784);
or UO_371 (O_371,N_4525,N_4902);
and UO_372 (O_372,N_4511,N_4823);
and UO_373 (O_373,N_4776,N_4844);
or UO_374 (O_374,N_4972,N_4528);
or UO_375 (O_375,N_4542,N_4669);
nor UO_376 (O_376,N_4606,N_4616);
nor UO_377 (O_377,N_4805,N_4572);
or UO_378 (O_378,N_4591,N_4531);
and UO_379 (O_379,N_4514,N_4617);
nand UO_380 (O_380,N_4742,N_4653);
nand UO_381 (O_381,N_4931,N_4978);
and UO_382 (O_382,N_4524,N_4739);
nor UO_383 (O_383,N_4830,N_4548);
nand UO_384 (O_384,N_4882,N_4615);
or UO_385 (O_385,N_4945,N_4612);
nor UO_386 (O_386,N_4836,N_4511);
nor UO_387 (O_387,N_4674,N_4627);
or UO_388 (O_388,N_4665,N_4633);
or UO_389 (O_389,N_4523,N_4618);
nand UO_390 (O_390,N_4978,N_4816);
and UO_391 (O_391,N_4556,N_4861);
nand UO_392 (O_392,N_4577,N_4668);
nor UO_393 (O_393,N_4657,N_4795);
nand UO_394 (O_394,N_4552,N_4529);
nand UO_395 (O_395,N_4675,N_4826);
or UO_396 (O_396,N_4913,N_4773);
and UO_397 (O_397,N_4685,N_4946);
nand UO_398 (O_398,N_4989,N_4798);
and UO_399 (O_399,N_4912,N_4757);
nor UO_400 (O_400,N_4720,N_4774);
nor UO_401 (O_401,N_4842,N_4851);
xnor UO_402 (O_402,N_4624,N_4890);
nor UO_403 (O_403,N_4745,N_4641);
and UO_404 (O_404,N_4917,N_4523);
and UO_405 (O_405,N_4730,N_4784);
nand UO_406 (O_406,N_4932,N_4775);
and UO_407 (O_407,N_4928,N_4768);
nor UO_408 (O_408,N_4817,N_4601);
nor UO_409 (O_409,N_4770,N_4559);
and UO_410 (O_410,N_4645,N_4551);
or UO_411 (O_411,N_4549,N_4932);
and UO_412 (O_412,N_4651,N_4741);
and UO_413 (O_413,N_4802,N_4997);
nand UO_414 (O_414,N_4859,N_4671);
or UO_415 (O_415,N_4830,N_4562);
and UO_416 (O_416,N_4697,N_4610);
nand UO_417 (O_417,N_4554,N_4699);
or UO_418 (O_418,N_4825,N_4949);
and UO_419 (O_419,N_4923,N_4723);
nand UO_420 (O_420,N_4796,N_4837);
nand UO_421 (O_421,N_4937,N_4578);
xnor UO_422 (O_422,N_4830,N_4590);
or UO_423 (O_423,N_4550,N_4772);
or UO_424 (O_424,N_4618,N_4518);
nand UO_425 (O_425,N_4997,N_4978);
nor UO_426 (O_426,N_4762,N_4991);
nand UO_427 (O_427,N_4850,N_4759);
or UO_428 (O_428,N_4870,N_4980);
and UO_429 (O_429,N_4595,N_4975);
nand UO_430 (O_430,N_4580,N_4538);
and UO_431 (O_431,N_4589,N_4548);
and UO_432 (O_432,N_4694,N_4730);
and UO_433 (O_433,N_4975,N_4717);
or UO_434 (O_434,N_4550,N_4543);
xor UO_435 (O_435,N_4769,N_4956);
or UO_436 (O_436,N_4997,N_4777);
nor UO_437 (O_437,N_4519,N_4594);
or UO_438 (O_438,N_4742,N_4945);
or UO_439 (O_439,N_4873,N_4762);
nand UO_440 (O_440,N_4920,N_4540);
nor UO_441 (O_441,N_4512,N_4766);
and UO_442 (O_442,N_4687,N_4699);
nor UO_443 (O_443,N_4826,N_4653);
or UO_444 (O_444,N_4903,N_4892);
and UO_445 (O_445,N_4588,N_4518);
nor UO_446 (O_446,N_4925,N_4903);
and UO_447 (O_447,N_4543,N_4640);
or UO_448 (O_448,N_4923,N_4798);
and UO_449 (O_449,N_4587,N_4559);
or UO_450 (O_450,N_4543,N_4835);
and UO_451 (O_451,N_4541,N_4696);
and UO_452 (O_452,N_4659,N_4993);
nor UO_453 (O_453,N_4786,N_4880);
or UO_454 (O_454,N_4884,N_4900);
and UO_455 (O_455,N_4828,N_4792);
nand UO_456 (O_456,N_4587,N_4537);
nor UO_457 (O_457,N_4525,N_4516);
nand UO_458 (O_458,N_4503,N_4593);
nor UO_459 (O_459,N_4795,N_4791);
nand UO_460 (O_460,N_4660,N_4937);
or UO_461 (O_461,N_4503,N_4800);
nand UO_462 (O_462,N_4837,N_4682);
or UO_463 (O_463,N_4538,N_4775);
and UO_464 (O_464,N_4558,N_4740);
xor UO_465 (O_465,N_4979,N_4573);
or UO_466 (O_466,N_4876,N_4871);
or UO_467 (O_467,N_4564,N_4690);
nand UO_468 (O_468,N_4607,N_4891);
or UO_469 (O_469,N_4672,N_4962);
or UO_470 (O_470,N_4595,N_4663);
or UO_471 (O_471,N_4917,N_4845);
nor UO_472 (O_472,N_4749,N_4500);
or UO_473 (O_473,N_4656,N_4776);
and UO_474 (O_474,N_4817,N_4679);
nor UO_475 (O_475,N_4503,N_4500);
nor UO_476 (O_476,N_4703,N_4911);
xnor UO_477 (O_477,N_4730,N_4707);
nand UO_478 (O_478,N_4723,N_4519);
or UO_479 (O_479,N_4788,N_4650);
nor UO_480 (O_480,N_4832,N_4841);
or UO_481 (O_481,N_4842,N_4779);
nor UO_482 (O_482,N_4536,N_4755);
nor UO_483 (O_483,N_4828,N_4731);
nor UO_484 (O_484,N_4983,N_4595);
nand UO_485 (O_485,N_4535,N_4823);
nand UO_486 (O_486,N_4517,N_4844);
nand UO_487 (O_487,N_4832,N_4518);
or UO_488 (O_488,N_4695,N_4548);
and UO_489 (O_489,N_4730,N_4791);
nor UO_490 (O_490,N_4501,N_4880);
nand UO_491 (O_491,N_4804,N_4673);
nor UO_492 (O_492,N_4798,N_4602);
nor UO_493 (O_493,N_4726,N_4506);
and UO_494 (O_494,N_4961,N_4659);
xnor UO_495 (O_495,N_4526,N_4734);
and UO_496 (O_496,N_4986,N_4847);
nor UO_497 (O_497,N_4505,N_4537);
or UO_498 (O_498,N_4994,N_4940);
nor UO_499 (O_499,N_4835,N_4661);
nor UO_500 (O_500,N_4715,N_4767);
nand UO_501 (O_501,N_4724,N_4866);
nor UO_502 (O_502,N_4710,N_4797);
and UO_503 (O_503,N_4582,N_4588);
and UO_504 (O_504,N_4921,N_4844);
nand UO_505 (O_505,N_4539,N_4907);
nor UO_506 (O_506,N_4778,N_4589);
or UO_507 (O_507,N_4945,N_4900);
or UO_508 (O_508,N_4843,N_4608);
nand UO_509 (O_509,N_4924,N_4901);
xnor UO_510 (O_510,N_4642,N_4791);
nand UO_511 (O_511,N_4971,N_4640);
nor UO_512 (O_512,N_4753,N_4629);
nor UO_513 (O_513,N_4894,N_4630);
nand UO_514 (O_514,N_4809,N_4538);
nor UO_515 (O_515,N_4844,N_4516);
nor UO_516 (O_516,N_4983,N_4816);
nand UO_517 (O_517,N_4771,N_4640);
and UO_518 (O_518,N_4649,N_4595);
and UO_519 (O_519,N_4771,N_4757);
and UO_520 (O_520,N_4983,N_4531);
nand UO_521 (O_521,N_4933,N_4837);
nor UO_522 (O_522,N_4945,N_4835);
or UO_523 (O_523,N_4554,N_4673);
and UO_524 (O_524,N_4868,N_4689);
nand UO_525 (O_525,N_4704,N_4541);
or UO_526 (O_526,N_4547,N_4694);
and UO_527 (O_527,N_4765,N_4531);
and UO_528 (O_528,N_4692,N_4879);
nor UO_529 (O_529,N_4811,N_4870);
nor UO_530 (O_530,N_4628,N_4725);
and UO_531 (O_531,N_4710,N_4509);
and UO_532 (O_532,N_4782,N_4684);
nand UO_533 (O_533,N_4844,N_4506);
nor UO_534 (O_534,N_4881,N_4748);
or UO_535 (O_535,N_4598,N_4608);
and UO_536 (O_536,N_4899,N_4689);
or UO_537 (O_537,N_4645,N_4803);
nor UO_538 (O_538,N_4753,N_4696);
and UO_539 (O_539,N_4972,N_4937);
and UO_540 (O_540,N_4585,N_4697);
nand UO_541 (O_541,N_4532,N_4827);
or UO_542 (O_542,N_4822,N_4503);
and UO_543 (O_543,N_4632,N_4616);
and UO_544 (O_544,N_4657,N_4734);
and UO_545 (O_545,N_4541,N_4741);
nand UO_546 (O_546,N_4695,N_4893);
or UO_547 (O_547,N_4887,N_4678);
and UO_548 (O_548,N_4655,N_4910);
and UO_549 (O_549,N_4670,N_4692);
nor UO_550 (O_550,N_4914,N_4654);
nor UO_551 (O_551,N_4748,N_4880);
nand UO_552 (O_552,N_4959,N_4511);
nand UO_553 (O_553,N_4868,N_4669);
and UO_554 (O_554,N_4939,N_4753);
and UO_555 (O_555,N_4743,N_4557);
or UO_556 (O_556,N_4732,N_4742);
nor UO_557 (O_557,N_4598,N_4948);
nand UO_558 (O_558,N_4824,N_4828);
xor UO_559 (O_559,N_4957,N_4579);
nand UO_560 (O_560,N_4814,N_4648);
nor UO_561 (O_561,N_4506,N_4957);
nand UO_562 (O_562,N_4919,N_4706);
and UO_563 (O_563,N_4523,N_4727);
and UO_564 (O_564,N_4639,N_4651);
or UO_565 (O_565,N_4564,N_4519);
and UO_566 (O_566,N_4801,N_4588);
and UO_567 (O_567,N_4530,N_4763);
nor UO_568 (O_568,N_4846,N_4633);
or UO_569 (O_569,N_4667,N_4646);
nor UO_570 (O_570,N_4520,N_4831);
and UO_571 (O_571,N_4917,N_4735);
or UO_572 (O_572,N_4590,N_4616);
or UO_573 (O_573,N_4929,N_4918);
and UO_574 (O_574,N_4574,N_4900);
nand UO_575 (O_575,N_4591,N_4620);
and UO_576 (O_576,N_4879,N_4938);
nor UO_577 (O_577,N_4675,N_4521);
and UO_578 (O_578,N_4532,N_4869);
nor UO_579 (O_579,N_4875,N_4743);
and UO_580 (O_580,N_4872,N_4999);
nor UO_581 (O_581,N_4543,N_4711);
nor UO_582 (O_582,N_4760,N_4540);
nor UO_583 (O_583,N_4620,N_4985);
nor UO_584 (O_584,N_4766,N_4933);
nand UO_585 (O_585,N_4678,N_4992);
and UO_586 (O_586,N_4635,N_4582);
and UO_587 (O_587,N_4678,N_4609);
nand UO_588 (O_588,N_4781,N_4957);
nor UO_589 (O_589,N_4544,N_4581);
nor UO_590 (O_590,N_4919,N_4540);
and UO_591 (O_591,N_4574,N_4936);
nor UO_592 (O_592,N_4605,N_4528);
or UO_593 (O_593,N_4962,N_4548);
and UO_594 (O_594,N_4654,N_4630);
and UO_595 (O_595,N_4595,N_4894);
nor UO_596 (O_596,N_4825,N_4932);
and UO_597 (O_597,N_4880,N_4810);
and UO_598 (O_598,N_4507,N_4740);
and UO_599 (O_599,N_4591,N_4603);
and UO_600 (O_600,N_4930,N_4566);
or UO_601 (O_601,N_4998,N_4911);
nor UO_602 (O_602,N_4914,N_4511);
or UO_603 (O_603,N_4906,N_4674);
xnor UO_604 (O_604,N_4504,N_4592);
or UO_605 (O_605,N_4714,N_4592);
nor UO_606 (O_606,N_4919,N_4506);
or UO_607 (O_607,N_4670,N_4508);
nand UO_608 (O_608,N_4773,N_4707);
xnor UO_609 (O_609,N_4791,N_4818);
xnor UO_610 (O_610,N_4685,N_4648);
or UO_611 (O_611,N_4906,N_4528);
nand UO_612 (O_612,N_4807,N_4889);
nand UO_613 (O_613,N_4944,N_4665);
or UO_614 (O_614,N_4617,N_4723);
and UO_615 (O_615,N_4654,N_4911);
nand UO_616 (O_616,N_4670,N_4505);
and UO_617 (O_617,N_4508,N_4911);
nand UO_618 (O_618,N_4606,N_4653);
or UO_619 (O_619,N_4516,N_4614);
nand UO_620 (O_620,N_4734,N_4961);
nand UO_621 (O_621,N_4792,N_4682);
nor UO_622 (O_622,N_4657,N_4598);
nand UO_623 (O_623,N_4873,N_4565);
or UO_624 (O_624,N_4967,N_4772);
nor UO_625 (O_625,N_4625,N_4851);
or UO_626 (O_626,N_4764,N_4732);
and UO_627 (O_627,N_4767,N_4713);
nor UO_628 (O_628,N_4968,N_4807);
nand UO_629 (O_629,N_4662,N_4627);
nor UO_630 (O_630,N_4990,N_4955);
and UO_631 (O_631,N_4862,N_4712);
nor UO_632 (O_632,N_4838,N_4532);
nor UO_633 (O_633,N_4773,N_4579);
or UO_634 (O_634,N_4846,N_4511);
nor UO_635 (O_635,N_4879,N_4931);
and UO_636 (O_636,N_4719,N_4544);
and UO_637 (O_637,N_4508,N_4832);
or UO_638 (O_638,N_4841,N_4724);
and UO_639 (O_639,N_4947,N_4801);
nor UO_640 (O_640,N_4535,N_4526);
nor UO_641 (O_641,N_4839,N_4737);
nor UO_642 (O_642,N_4815,N_4685);
and UO_643 (O_643,N_4581,N_4872);
nand UO_644 (O_644,N_4920,N_4645);
nand UO_645 (O_645,N_4831,N_4756);
or UO_646 (O_646,N_4516,N_4807);
nor UO_647 (O_647,N_4873,N_4504);
and UO_648 (O_648,N_4619,N_4970);
nand UO_649 (O_649,N_4676,N_4648);
or UO_650 (O_650,N_4982,N_4843);
or UO_651 (O_651,N_4669,N_4973);
nor UO_652 (O_652,N_4570,N_4885);
or UO_653 (O_653,N_4613,N_4543);
nand UO_654 (O_654,N_4828,N_4839);
and UO_655 (O_655,N_4785,N_4698);
and UO_656 (O_656,N_4948,N_4588);
nand UO_657 (O_657,N_4827,N_4666);
and UO_658 (O_658,N_4780,N_4970);
nand UO_659 (O_659,N_4608,N_4593);
or UO_660 (O_660,N_4665,N_4865);
or UO_661 (O_661,N_4830,N_4877);
and UO_662 (O_662,N_4615,N_4964);
nor UO_663 (O_663,N_4654,N_4799);
nor UO_664 (O_664,N_4718,N_4707);
nand UO_665 (O_665,N_4650,N_4890);
or UO_666 (O_666,N_4674,N_4551);
or UO_667 (O_667,N_4865,N_4571);
or UO_668 (O_668,N_4831,N_4699);
xnor UO_669 (O_669,N_4733,N_4692);
nor UO_670 (O_670,N_4652,N_4683);
nor UO_671 (O_671,N_4501,N_4782);
or UO_672 (O_672,N_4551,N_4949);
and UO_673 (O_673,N_4558,N_4757);
nand UO_674 (O_674,N_4621,N_4502);
and UO_675 (O_675,N_4967,N_4568);
nand UO_676 (O_676,N_4713,N_4909);
or UO_677 (O_677,N_4639,N_4782);
nor UO_678 (O_678,N_4847,N_4983);
nand UO_679 (O_679,N_4713,N_4921);
nand UO_680 (O_680,N_4732,N_4920);
and UO_681 (O_681,N_4560,N_4651);
nor UO_682 (O_682,N_4579,N_4750);
nand UO_683 (O_683,N_4582,N_4985);
nor UO_684 (O_684,N_4547,N_4599);
nand UO_685 (O_685,N_4628,N_4851);
nand UO_686 (O_686,N_4601,N_4653);
nand UO_687 (O_687,N_4509,N_4569);
nor UO_688 (O_688,N_4788,N_4955);
and UO_689 (O_689,N_4997,N_4547);
nor UO_690 (O_690,N_4657,N_4865);
nand UO_691 (O_691,N_4764,N_4923);
and UO_692 (O_692,N_4638,N_4996);
nand UO_693 (O_693,N_4530,N_4963);
nand UO_694 (O_694,N_4996,N_4667);
nand UO_695 (O_695,N_4567,N_4600);
nor UO_696 (O_696,N_4769,N_4944);
nand UO_697 (O_697,N_4896,N_4751);
and UO_698 (O_698,N_4576,N_4980);
nor UO_699 (O_699,N_4783,N_4797);
and UO_700 (O_700,N_4977,N_4587);
nand UO_701 (O_701,N_4691,N_4597);
nand UO_702 (O_702,N_4541,N_4751);
nand UO_703 (O_703,N_4896,N_4845);
or UO_704 (O_704,N_4843,N_4524);
or UO_705 (O_705,N_4923,N_4647);
and UO_706 (O_706,N_4949,N_4876);
nor UO_707 (O_707,N_4763,N_4939);
and UO_708 (O_708,N_4712,N_4801);
or UO_709 (O_709,N_4593,N_4892);
nand UO_710 (O_710,N_4680,N_4876);
nand UO_711 (O_711,N_4515,N_4736);
nand UO_712 (O_712,N_4691,N_4815);
and UO_713 (O_713,N_4688,N_4715);
and UO_714 (O_714,N_4576,N_4714);
and UO_715 (O_715,N_4754,N_4916);
or UO_716 (O_716,N_4511,N_4512);
and UO_717 (O_717,N_4551,N_4983);
nand UO_718 (O_718,N_4955,N_4509);
xnor UO_719 (O_719,N_4677,N_4583);
or UO_720 (O_720,N_4904,N_4972);
nor UO_721 (O_721,N_4820,N_4671);
nor UO_722 (O_722,N_4613,N_4972);
and UO_723 (O_723,N_4619,N_4954);
nor UO_724 (O_724,N_4920,N_4780);
or UO_725 (O_725,N_4797,N_4853);
and UO_726 (O_726,N_4780,N_4956);
or UO_727 (O_727,N_4688,N_4610);
nand UO_728 (O_728,N_4818,N_4691);
and UO_729 (O_729,N_4532,N_4725);
nand UO_730 (O_730,N_4759,N_4831);
or UO_731 (O_731,N_4780,N_4735);
xor UO_732 (O_732,N_4677,N_4580);
nand UO_733 (O_733,N_4836,N_4626);
nor UO_734 (O_734,N_4983,N_4958);
nor UO_735 (O_735,N_4873,N_4787);
nand UO_736 (O_736,N_4526,N_4505);
nor UO_737 (O_737,N_4924,N_4813);
nor UO_738 (O_738,N_4950,N_4952);
nor UO_739 (O_739,N_4718,N_4974);
nor UO_740 (O_740,N_4571,N_4798);
or UO_741 (O_741,N_4605,N_4738);
or UO_742 (O_742,N_4759,N_4696);
and UO_743 (O_743,N_4959,N_4949);
nand UO_744 (O_744,N_4876,N_4952);
or UO_745 (O_745,N_4787,N_4843);
or UO_746 (O_746,N_4586,N_4722);
nand UO_747 (O_747,N_4530,N_4889);
or UO_748 (O_748,N_4922,N_4967);
nand UO_749 (O_749,N_4894,N_4638);
or UO_750 (O_750,N_4972,N_4919);
and UO_751 (O_751,N_4697,N_4724);
and UO_752 (O_752,N_4875,N_4796);
or UO_753 (O_753,N_4967,N_4549);
nor UO_754 (O_754,N_4704,N_4924);
nand UO_755 (O_755,N_4612,N_4665);
and UO_756 (O_756,N_4718,N_4987);
or UO_757 (O_757,N_4907,N_4917);
xor UO_758 (O_758,N_4697,N_4569);
or UO_759 (O_759,N_4617,N_4730);
nand UO_760 (O_760,N_4526,N_4579);
nor UO_761 (O_761,N_4586,N_4568);
and UO_762 (O_762,N_4617,N_4933);
and UO_763 (O_763,N_4750,N_4696);
nor UO_764 (O_764,N_4568,N_4827);
and UO_765 (O_765,N_4536,N_4736);
or UO_766 (O_766,N_4872,N_4784);
or UO_767 (O_767,N_4910,N_4946);
nand UO_768 (O_768,N_4553,N_4943);
and UO_769 (O_769,N_4567,N_4628);
nor UO_770 (O_770,N_4677,N_4771);
and UO_771 (O_771,N_4867,N_4842);
nor UO_772 (O_772,N_4992,N_4645);
nor UO_773 (O_773,N_4855,N_4842);
nand UO_774 (O_774,N_4680,N_4932);
and UO_775 (O_775,N_4811,N_4835);
and UO_776 (O_776,N_4844,N_4916);
or UO_777 (O_777,N_4615,N_4522);
nand UO_778 (O_778,N_4707,N_4757);
nor UO_779 (O_779,N_4520,N_4525);
nand UO_780 (O_780,N_4564,N_4881);
nand UO_781 (O_781,N_4709,N_4522);
and UO_782 (O_782,N_4900,N_4850);
nor UO_783 (O_783,N_4539,N_4578);
and UO_784 (O_784,N_4526,N_4700);
nand UO_785 (O_785,N_4772,N_4868);
and UO_786 (O_786,N_4961,N_4720);
and UO_787 (O_787,N_4562,N_4550);
or UO_788 (O_788,N_4813,N_4971);
or UO_789 (O_789,N_4878,N_4865);
nor UO_790 (O_790,N_4794,N_4656);
and UO_791 (O_791,N_4851,N_4698);
nand UO_792 (O_792,N_4913,N_4932);
nand UO_793 (O_793,N_4536,N_4601);
or UO_794 (O_794,N_4579,N_4630);
and UO_795 (O_795,N_4501,N_4945);
nor UO_796 (O_796,N_4585,N_4997);
nor UO_797 (O_797,N_4795,N_4868);
and UO_798 (O_798,N_4727,N_4804);
or UO_799 (O_799,N_4679,N_4932);
and UO_800 (O_800,N_4597,N_4565);
or UO_801 (O_801,N_4654,N_4725);
and UO_802 (O_802,N_4984,N_4791);
nor UO_803 (O_803,N_4564,N_4502);
and UO_804 (O_804,N_4946,N_4947);
or UO_805 (O_805,N_4997,N_4842);
or UO_806 (O_806,N_4766,N_4802);
and UO_807 (O_807,N_4826,N_4755);
nand UO_808 (O_808,N_4738,N_4712);
and UO_809 (O_809,N_4874,N_4834);
or UO_810 (O_810,N_4902,N_4529);
and UO_811 (O_811,N_4850,N_4552);
nor UO_812 (O_812,N_4832,N_4713);
and UO_813 (O_813,N_4502,N_4788);
nor UO_814 (O_814,N_4912,N_4523);
and UO_815 (O_815,N_4890,N_4829);
or UO_816 (O_816,N_4876,N_4539);
nor UO_817 (O_817,N_4668,N_4870);
nor UO_818 (O_818,N_4534,N_4873);
nor UO_819 (O_819,N_4571,N_4656);
or UO_820 (O_820,N_4833,N_4912);
or UO_821 (O_821,N_4569,N_4649);
nand UO_822 (O_822,N_4663,N_4840);
and UO_823 (O_823,N_4749,N_4632);
nor UO_824 (O_824,N_4609,N_4829);
nor UO_825 (O_825,N_4559,N_4644);
or UO_826 (O_826,N_4642,N_4861);
xnor UO_827 (O_827,N_4637,N_4687);
or UO_828 (O_828,N_4869,N_4764);
nand UO_829 (O_829,N_4750,N_4590);
nand UO_830 (O_830,N_4567,N_4967);
or UO_831 (O_831,N_4547,N_4876);
nand UO_832 (O_832,N_4746,N_4602);
or UO_833 (O_833,N_4988,N_4754);
nand UO_834 (O_834,N_4509,N_4625);
or UO_835 (O_835,N_4771,N_4842);
or UO_836 (O_836,N_4977,N_4500);
or UO_837 (O_837,N_4931,N_4518);
nand UO_838 (O_838,N_4951,N_4587);
and UO_839 (O_839,N_4922,N_4564);
nor UO_840 (O_840,N_4794,N_4969);
nor UO_841 (O_841,N_4828,N_4797);
or UO_842 (O_842,N_4933,N_4720);
and UO_843 (O_843,N_4761,N_4754);
or UO_844 (O_844,N_4629,N_4917);
nor UO_845 (O_845,N_4588,N_4840);
xor UO_846 (O_846,N_4905,N_4880);
xnor UO_847 (O_847,N_4853,N_4591);
or UO_848 (O_848,N_4555,N_4739);
and UO_849 (O_849,N_4559,N_4591);
or UO_850 (O_850,N_4723,N_4634);
nand UO_851 (O_851,N_4636,N_4524);
or UO_852 (O_852,N_4658,N_4572);
or UO_853 (O_853,N_4895,N_4595);
nor UO_854 (O_854,N_4910,N_4718);
or UO_855 (O_855,N_4954,N_4830);
nor UO_856 (O_856,N_4755,N_4977);
nor UO_857 (O_857,N_4598,N_4717);
or UO_858 (O_858,N_4505,N_4617);
and UO_859 (O_859,N_4901,N_4675);
or UO_860 (O_860,N_4671,N_4848);
or UO_861 (O_861,N_4793,N_4751);
nor UO_862 (O_862,N_4994,N_4988);
nand UO_863 (O_863,N_4942,N_4532);
or UO_864 (O_864,N_4894,N_4541);
xor UO_865 (O_865,N_4596,N_4631);
or UO_866 (O_866,N_4879,N_4835);
and UO_867 (O_867,N_4785,N_4934);
nand UO_868 (O_868,N_4856,N_4917);
nand UO_869 (O_869,N_4530,N_4728);
and UO_870 (O_870,N_4672,N_4573);
nand UO_871 (O_871,N_4581,N_4781);
nand UO_872 (O_872,N_4753,N_4838);
or UO_873 (O_873,N_4882,N_4799);
nor UO_874 (O_874,N_4734,N_4831);
nand UO_875 (O_875,N_4763,N_4985);
nand UO_876 (O_876,N_4682,N_4626);
and UO_877 (O_877,N_4516,N_4550);
nor UO_878 (O_878,N_4726,N_4503);
nor UO_879 (O_879,N_4653,N_4904);
or UO_880 (O_880,N_4845,N_4861);
nand UO_881 (O_881,N_4914,N_4555);
nor UO_882 (O_882,N_4666,N_4603);
nor UO_883 (O_883,N_4576,N_4618);
or UO_884 (O_884,N_4685,N_4910);
and UO_885 (O_885,N_4791,N_4546);
and UO_886 (O_886,N_4701,N_4593);
or UO_887 (O_887,N_4966,N_4624);
and UO_888 (O_888,N_4661,N_4976);
nand UO_889 (O_889,N_4520,N_4647);
nand UO_890 (O_890,N_4578,N_4973);
and UO_891 (O_891,N_4626,N_4687);
nand UO_892 (O_892,N_4605,N_4676);
or UO_893 (O_893,N_4815,N_4507);
and UO_894 (O_894,N_4663,N_4949);
nand UO_895 (O_895,N_4972,N_4888);
and UO_896 (O_896,N_4501,N_4677);
or UO_897 (O_897,N_4779,N_4774);
or UO_898 (O_898,N_4738,N_4923);
nor UO_899 (O_899,N_4624,N_4756);
or UO_900 (O_900,N_4641,N_4990);
and UO_901 (O_901,N_4538,N_4759);
and UO_902 (O_902,N_4524,N_4603);
xnor UO_903 (O_903,N_4851,N_4725);
nand UO_904 (O_904,N_4788,N_4729);
nor UO_905 (O_905,N_4601,N_4849);
nor UO_906 (O_906,N_4589,N_4767);
and UO_907 (O_907,N_4662,N_4557);
or UO_908 (O_908,N_4608,N_4741);
nand UO_909 (O_909,N_4514,N_4813);
or UO_910 (O_910,N_4585,N_4745);
or UO_911 (O_911,N_4978,N_4811);
or UO_912 (O_912,N_4943,N_4884);
and UO_913 (O_913,N_4762,N_4822);
and UO_914 (O_914,N_4685,N_4554);
nand UO_915 (O_915,N_4700,N_4592);
nor UO_916 (O_916,N_4627,N_4777);
nor UO_917 (O_917,N_4514,N_4507);
xor UO_918 (O_918,N_4641,N_4646);
nand UO_919 (O_919,N_4927,N_4602);
or UO_920 (O_920,N_4957,N_4709);
nand UO_921 (O_921,N_4913,N_4848);
nand UO_922 (O_922,N_4729,N_4580);
or UO_923 (O_923,N_4684,N_4523);
nor UO_924 (O_924,N_4503,N_4948);
or UO_925 (O_925,N_4826,N_4983);
nand UO_926 (O_926,N_4974,N_4687);
nor UO_927 (O_927,N_4868,N_4701);
and UO_928 (O_928,N_4906,N_4589);
nor UO_929 (O_929,N_4631,N_4713);
nor UO_930 (O_930,N_4821,N_4853);
and UO_931 (O_931,N_4853,N_4890);
or UO_932 (O_932,N_4660,N_4931);
and UO_933 (O_933,N_4863,N_4653);
nor UO_934 (O_934,N_4743,N_4556);
nor UO_935 (O_935,N_4927,N_4858);
xnor UO_936 (O_936,N_4619,N_4919);
or UO_937 (O_937,N_4991,N_4900);
or UO_938 (O_938,N_4663,N_4525);
nor UO_939 (O_939,N_4523,N_4925);
or UO_940 (O_940,N_4583,N_4828);
or UO_941 (O_941,N_4855,N_4548);
nand UO_942 (O_942,N_4664,N_4702);
or UO_943 (O_943,N_4521,N_4666);
or UO_944 (O_944,N_4746,N_4781);
nand UO_945 (O_945,N_4769,N_4934);
nand UO_946 (O_946,N_4522,N_4617);
nand UO_947 (O_947,N_4918,N_4982);
and UO_948 (O_948,N_4837,N_4663);
and UO_949 (O_949,N_4922,N_4662);
nor UO_950 (O_950,N_4654,N_4628);
or UO_951 (O_951,N_4728,N_4649);
or UO_952 (O_952,N_4629,N_4563);
nand UO_953 (O_953,N_4669,N_4910);
or UO_954 (O_954,N_4680,N_4908);
nor UO_955 (O_955,N_4942,N_4516);
or UO_956 (O_956,N_4746,N_4724);
nor UO_957 (O_957,N_4631,N_4909);
or UO_958 (O_958,N_4901,N_4663);
or UO_959 (O_959,N_4650,N_4915);
or UO_960 (O_960,N_4837,N_4922);
nand UO_961 (O_961,N_4786,N_4906);
nand UO_962 (O_962,N_4619,N_4719);
and UO_963 (O_963,N_4937,N_4875);
or UO_964 (O_964,N_4826,N_4950);
and UO_965 (O_965,N_4829,N_4654);
and UO_966 (O_966,N_4742,N_4957);
or UO_967 (O_967,N_4734,N_4926);
nor UO_968 (O_968,N_4509,N_4956);
or UO_969 (O_969,N_4565,N_4596);
nand UO_970 (O_970,N_4875,N_4992);
or UO_971 (O_971,N_4538,N_4656);
nor UO_972 (O_972,N_4541,N_4853);
nor UO_973 (O_973,N_4975,N_4805);
or UO_974 (O_974,N_4999,N_4895);
nand UO_975 (O_975,N_4867,N_4886);
nand UO_976 (O_976,N_4721,N_4915);
nor UO_977 (O_977,N_4823,N_4500);
and UO_978 (O_978,N_4523,N_4543);
or UO_979 (O_979,N_4623,N_4686);
nor UO_980 (O_980,N_4806,N_4521);
and UO_981 (O_981,N_4526,N_4630);
nand UO_982 (O_982,N_4968,N_4999);
nor UO_983 (O_983,N_4600,N_4671);
and UO_984 (O_984,N_4531,N_4813);
nand UO_985 (O_985,N_4738,N_4974);
xnor UO_986 (O_986,N_4719,N_4773);
nand UO_987 (O_987,N_4685,N_4613);
nor UO_988 (O_988,N_4526,N_4648);
or UO_989 (O_989,N_4628,N_4996);
or UO_990 (O_990,N_4820,N_4997);
nor UO_991 (O_991,N_4667,N_4830);
nand UO_992 (O_992,N_4655,N_4866);
and UO_993 (O_993,N_4512,N_4694);
or UO_994 (O_994,N_4879,N_4636);
nand UO_995 (O_995,N_4715,N_4968);
and UO_996 (O_996,N_4848,N_4749);
and UO_997 (O_997,N_4685,N_4833);
and UO_998 (O_998,N_4521,N_4595);
and UO_999 (O_999,N_4637,N_4507);
endmodule