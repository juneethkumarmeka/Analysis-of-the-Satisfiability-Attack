module basic_2000_20000_2500_100_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_668,In_1553);
nor U1 (N_1,In_756,In_313);
nand U2 (N_2,In_1163,In_356);
nand U3 (N_3,In_804,In_460);
xor U4 (N_4,In_1862,In_1669);
nand U5 (N_5,In_1707,In_321);
nand U6 (N_6,In_1739,In_673);
xor U7 (N_7,In_743,In_108);
or U8 (N_8,In_1458,In_383);
xnor U9 (N_9,In_1251,In_784);
xnor U10 (N_10,In_613,In_975);
and U11 (N_11,In_954,In_1535);
nand U12 (N_12,In_1182,In_652);
xor U13 (N_13,In_646,In_865);
nand U14 (N_14,In_75,In_221);
xor U15 (N_15,In_828,In_1501);
and U16 (N_16,In_366,In_1289);
or U17 (N_17,In_1278,In_1878);
nor U18 (N_18,In_480,In_1870);
nand U19 (N_19,In_1990,In_918);
xnor U20 (N_20,In_22,In_279);
or U21 (N_21,In_1088,In_1113);
or U22 (N_22,In_219,In_380);
or U23 (N_23,In_370,In_821);
and U24 (N_24,In_131,In_1534);
xor U25 (N_25,In_1295,In_1936);
nand U26 (N_26,In_1116,In_361);
and U27 (N_27,In_1581,In_156);
xor U28 (N_28,In_1191,In_116);
or U29 (N_29,In_80,In_708);
and U30 (N_30,In_332,In_850);
or U31 (N_31,In_1793,In_766);
nand U32 (N_32,In_1290,In_642);
nand U33 (N_33,In_1482,In_1008);
nand U34 (N_34,In_189,In_1005);
and U35 (N_35,In_433,In_586);
nor U36 (N_36,In_879,In_76);
nand U37 (N_37,In_495,In_952);
and U38 (N_38,In_1033,In_1966);
and U39 (N_39,In_549,In_62);
and U40 (N_40,In_1179,In_1794);
nand U41 (N_41,In_771,In_1048);
or U42 (N_42,In_883,In_599);
xor U43 (N_43,In_143,In_896);
nand U44 (N_44,In_1331,In_653);
nand U45 (N_45,In_1464,In_1655);
and U46 (N_46,In_1454,In_477);
and U47 (N_47,In_1624,In_1880);
or U48 (N_48,In_364,In_455);
or U49 (N_49,In_1060,In_450);
or U50 (N_50,In_691,In_331);
and U51 (N_51,In_1531,In_1571);
and U52 (N_52,In_1902,In_773);
xnor U53 (N_53,In_163,In_1114);
nor U54 (N_54,In_1888,In_580);
nand U55 (N_55,In_961,In_991);
nor U56 (N_56,In_393,In_1002);
nand U57 (N_57,In_630,In_685);
and U58 (N_58,In_1219,In_1420);
or U59 (N_59,In_248,In_700);
and U60 (N_60,In_1737,In_1968);
and U61 (N_61,In_791,In_699);
and U62 (N_62,In_1627,In_1500);
or U63 (N_63,In_641,In_262);
xor U64 (N_64,In_794,In_768);
or U65 (N_65,In_201,In_1859);
nor U66 (N_66,In_1897,In_1914);
and U67 (N_67,In_1211,In_500);
nand U68 (N_68,In_1233,In_417);
and U69 (N_69,In_396,In_1177);
nand U70 (N_70,In_795,In_144);
xnor U71 (N_71,In_1046,In_1674);
or U72 (N_72,In_1169,In_1073);
and U73 (N_73,In_1195,In_1315);
nor U74 (N_74,In_435,In_1103);
xnor U75 (N_75,In_1619,In_1801);
nor U76 (N_76,In_504,In_1988);
nand U77 (N_77,In_360,In_409);
nor U78 (N_78,In_1323,In_792);
nand U79 (N_79,In_342,In_1369);
xnor U80 (N_80,In_1950,In_899);
nor U81 (N_81,In_245,In_702);
or U82 (N_82,In_114,In_1283);
nor U83 (N_83,In_1330,In_1561);
or U84 (N_84,In_1814,In_538);
xnor U85 (N_85,In_437,In_90);
and U86 (N_86,In_742,In_5);
or U87 (N_87,In_11,In_870);
and U88 (N_88,In_884,In_1221);
or U89 (N_89,In_544,In_1496);
and U90 (N_90,In_1190,In_823);
or U91 (N_91,In_1383,In_929);
xor U92 (N_92,In_927,In_329);
or U93 (N_93,In_166,In_1480);
nor U94 (N_94,In_953,In_634);
and U95 (N_95,In_1151,In_514);
xnor U96 (N_96,In_1587,In_1522);
nand U97 (N_97,In_782,In_434);
nor U98 (N_98,In_1145,In_1997);
xnor U99 (N_99,In_1376,In_1452);
nor U100 (N_100,In_1134,In_1017);
nand U101 (N_101,In_1625,In_1064);
nor U102 (N_102,In_632,In_1717);
nand U103 (N_103,In_923,In_119);
and U104 (N_104,In_1379,In_733);
or U105 (N_105,In_1370,In_1952);
nand U106 (N_106,In_620,In_501);
xnor U107 (N_107,In_1304,In_858);
and U108 (N_108,In_1385,In_150);
and U109 (N_109,In_1319,In_1960);
nand U110 (N_110,In_648,In_415);
and U111 (N_111,In_349,In_1162);
and U112 (N_112,In_1810,In_844);
or U113 (N_113,In_1932,In_604);
nand U114 (N_114,In_1956,In_252);
nor U115 (N_115,In_1300,In_1983);
and U116 (N_116,In_1846,In_1631);
and U117 (N_117,In_1909,In_135);
xnor U118 (N_118,In_1682,In_720);
nor U119 (N_119,In_1549,In_1259);
nand U120 (N_120,In_1779,In_46);
or U121 (N_121,In_1227,In_1636);
nor U122 (N_122,In_461,In_617);
nand U123 (N_123,In_564,In_1099);
or U124 (N_124,In_631,In_511);
nand U125 (N_125,In_32,In_280);
nand U126 (N_126,In_831,In_488);
and U127 (N_127,In_846,In_1509);
or U128 (N_128,In_320,In_1542);
xnor U129 (N_129,In_354,In_519);
nor U130 (N_130,In_1266,In_925);
nand U131 (N_131,In_1071,In_355);
and U132 (N_132,In_340,In_1159);
and U133 (N_133,In_1398,In_1855);
and U134 (N_134,In_23,In_1638);
or U135 (N_135,In_1730,In_573);
xnor U136 (N_136,In_1362,In_161);
xnor U137 (N_137,In_1461,In_471);
and U138 (N_138,In_198,In_203);
nor U139 (N_139,In_1848,In_177);
nand U140 (N_140,In_1132,In_608);
or U141 (N_141,In_148,In_359);
nand U142 (N_142,In_1937,In_1395);
nand U143 (N_143,In_1204,In_1075);
and U144 (N_144,In_1731,In_1070);
xnor U145 (N_145,In_241,In_52);
nand U146 (N_146,In_1170,In_1043);
nor U147 (N_147,In_1945,In_1382);
or U148 (N_148,In_847,In_1757);
nand U149 (N_149,In_1813,In_350);
or U150 (N_150,In_137,In_1506);
and U151 (N_151,In_1441,In_1488);
or U152 (N_152,In_1551,In_1687);
nand U153 (N_153,In_1519,In_1618);
and U154 (N_154,In_226,In_17);
or U155 (N_155,In_81,In_1450);
nand U156 (N_156,In_1883,In_817);
nor U157 (N_157,In_751,In_1664);
nor U158 (N_158,In_1093,In_1605);
nor U159 (N_159,In_659,In_240);
nand U160 (N_160,In_266,In_1746);
or U161 (N_161,In_1372,In_748);
and U162 (N_162,In_338,In_173);
xnor U163 (N_163,In_20,In_315);
xnor U164 (N_164,In_1640,In_272);
xnor U165 (N_165,In_1394,In_346);
nand U166 (N_166,In_1986,In_502);
and U167 (N_167,In_1147,In_717);
nor U168 (N_168,In_1332,In_1063);
nor U169 (N_169,In_1051,In_696);
or U170 (N_170,In_1250,In_1028);
xor U171 (N_171,In_1938,In_1939);
xnor U172 (N_172,In_1342,In_594);
nor U173 (N_173,In_1595,In_664);
or U174 (N_174,In_1146,In_1351);
nor U175 (N_175,In_1041,In_107);
nand U176 (N_176,In_1069,In_440);
and U177 (N_177,In_1807,In_299);
nor U178 (N_178,In_429,In_864);
and U179 (N_179,In_1261,In_302);
or U180 (N_180,In_412,In_1306);
xnor U181 (N_181,In_808,In_209);
nor U182 (N_182,In_1785,In_1107);
xnor U183 (N_183,In_1702,In_1040);
xnor U184 (N_184,In_783,In_935);
xnor U185 (N_185,In_1317,In_420);
or U186 (N_186,In_1431,In_258);
nand U187 (N_187,In_1439,In_405);
or U188 (N_188,In_932,In_1076);
or U189 (N_189,In_1958,In_764);
or U190 (N_190,In_1877,In_97);
or U191 (N_191,In_352,In_1314);
xor U192 (N_192,In_1526,In_1565);
nor U193 (N_193,In_555,In_1856);
or U194 (N_194,In_1733,In_515);
nor U195 (N_195,In_1675,In_138);
or U196 (N_196,In_196,In_1079);
xor U197 (N_197,In_277,In_1769);
and U198 (N_198,In_1035,In_686);
nor U199 (N_199,In_669,In_85);
xor U200 (N_200,In_936,In_543);
and U201 (N_201,In_33,In_164);
xnor U202 (N_202,In_158,In_1156);
or U203 (N_203,N_91,In_224);
or U204 (N_204,In_259,In_275);
nand U205 (N_205,In_1206,In_1894);
nand U206 (N_206,In_183,In_1105);
or U207 (N_207,In_162,In_1131);
or U208 (N_208,N_104,In_176);
xor U209 (N_209,In_1401,In_67);
nor U210 (N_210,In_120,In_180);
or U211 (N_211,In_922,In_1994);
and U212 (N_212,In_368,In_1863);
or U213 (N_213,In_1455,In_997);
nor U214 (N_214,In_1047,N_101);
nor U215 (N_215,In_318,In_1776);
nor U216 (N_216,In_1288,In_799);
or U217 (N_217,In_895,In_944);
nor U218 (N_218,In_6,In_1586);
nor U219 (N_219,In_454,In_1792);
xor U220 (N_220,In_34,N_136);
nand U221 (N_221,In_1951,In_1699);
nor U222 (N_222,In_375,In_1828);
and U223 (N_223,In_1606,In_1973);
xor U224 (N_224,In_1912,In_7);
xor U225 (N_225,In_1826,In_1798);
nor U226 (N_226,In_1343,In_1649);
nand U227 (N_227,In_588,In_778);
and U228 (N_228,In_1641,In_570);
nor U229 (N_229,In_228,In_753);
xnor U230 (N_230,In_449,In_872);
nand U231 (N_231,In_1780,In_1208);
xnor U232 (N_232,N_174,In_339);
nand U233 (N_233,N_76,In_979);
and U234 (N_234,In_760,In_1141);
xor U235 (N_235,N_89,In_47);
nand U236 (N_236,In_45,In_1371);
nor U237 (N_237,In_607,In_1492);
and U238 (N_238,In_1056,N_53);
nor U239 (N_239,N_25,In_55);
and U240 (N_240,In_507,In_692);
and U241 (N_241,N_75,N_44);
or U242 (N_242,In_1505,N_148);
xnor U243 (N_243,In_9,In_1175);
nor U244 (N_244,In_963,In_1192);
xor U245 (N_245,In_1712,In_1767);
nand U246 (N_246,In_1689,In_1039);
xor U247 (N_247,In_1583,In_598);
and U248 (N_248,In_72,In_1822);
xnor U249 (N_249,In_1241,In_1670);
nand U250 (N_250,In_1930,In_1018);
or U251 (N_251,In_13,In_816);
and U252 (N_252,N_7,In_1212);
nand U253 (N_253,In_1710,In_1752);
or U254 (N_254,In_851,In_1965);
and U255 (N_255,In_1165,In_60);
nor U256 (N_256,In_1511,In_1515);
nor U257 (N_257,In_582,In_1708);
nor U258 (N_258,In_862,In_1200);
xor U259 (N_259,In_391,In_660);
xnor U260 (N_260,In_1078,In_1832);
or U261 (N_261,In_818,N_11);
and U262 (N_262,N_156,N_27);
and U263 (N_263,In_955,In_591);
or U264 (N_264,In_1310,In_1218);
nand U265 (N_265,In_242,In_394);
xor U266 (N_266,In_293,In_1836);
xor U267 (N_267,In_1484,In_1921);
nand U268 (N_268,In_1262,In_157);
nor U269 (N_269,In_662,In_466);
xor U270 (N_270,N_150,In_1238);
or U271 (N_271,In_1700,N_186);
xnor U272 (N_272,In_1665,In_348);
nor U273 (N_273,N_124,In_1889);
xor U274 (N_274,In_1612,In_267);
nor U275 (N_275,In_765,N_38);
nor U276 (N_276,In_386,In_64);
nor U277 (N_277,In_551,In_1774);
and U278 (N_278,In_459,In_19);
nor U279 (N_279,N_58,In_1438);
or U280 (N_280,N_151,In_1477);
nor U281 (N_281,N_28,N_179);
nand U282 (N_282,In_1629,In_1718);
nor U283 (N_283,In_644,In_897);
and U284 (N_284,In_210,In_890);
and U285 (N_285,In_1024,In_182);
and U286 (N_286,In_1280,In_188);
and U287 (N_287,In_377,In_1471);
xnor U288 (N_288,In_1235,In_1677);
nand U289 (N_289,In_465,In_129);
and U290 (N_290,N_54,In_898);
and U291 (N_291,N_22,In_1497);
nand U292 (N_292,In_1972,In_1974);
nand U293 (N_293,N_10,In_1337);
xnor U294 (N_294,In_1597,In_1691);
and U295 (N_295,In_635,In_398);
xnor U296 (N_296,In_1946,In_1352);
xnor U297 (N_297,In_1839,In_1916);
and U298 (N_298,N_195,In_1704);
and U299 (N_299,In_1365,In_21);
nand U300 (N_300,N_112,In_1311);
and U301 (N_301,N_52,In_616);
nor U302 (N_302,In_295,In_1536);
nand U303 (N_303,In_1294,In_980);
and U304 (N_304,In_1486,In_117);
xnor U305 (N_305,In_1007,In_841);
or U306 (N_306,In_351,In_1487);
nor U307 (N_307,In_367,N_123);
and U308 (N_308,In_694,N_120);
or U309 (N_309,N_196,In_1812);
or U310 (N_310,In_1264,In_561);
and U311 (N_311,In_1387,In_1281);
nand U312 (N_312,N_90,In_1166);
nor U313 (N_313,In_633,In_1562);
xor U314 (N_314,In_1596,In_1963);
xnor U315 (N_315,In_886,In_618);
nand U316 (N_316,In_880,N_6);
or U317 (N_317,In_655,In_649);
nand U318 (N_318,In_1819,N_184);
nand U319 (N_319,In_1180,In_1899);
xnor U320 (N_320,In_305,N_165);
nor U321 (N_321,N_181,In_1308);
or U322 (N_322,In_1434,In_807);
nor U323 (N_323,In_407,In_1258);
and U324 (N_324,In_1426,In_1396);
xor U325 (N_325,In_1554,N_141);
xor U326 (N_326,In_575,In_423);
nand U327 (N_327,In_727,In_610);
and U328 (N_328,In_571,In_704);
nand U329 (N_329,In_875,N_110);
xor U330 (N_330,In_637,In_413);
or U331 (N_331,In_1592,In_568);
nor U332 (N_332,In_548,In_845);
nand U333 (N_333,In_559,In_436);
and U334 (N_334,In_336,In_710);
or U335 (N_335,In_1891,In_921);
nand U336 (N_336,In_1504,In_110);
and U337 (N_337,In_1547,N_122);
or U338 (N_338,In_181,In_552);
nand U339 (N_339,In_452,N_145);
nand U340 (N_340,In_53,In_1481);
or U341 (N_341,In_913,In_1809);
xor U342 (N_342,In_1725,In_894);
xor U343 (N_343,In_1875,In_572);
and U344 (N_344,In_984,In_1226);
nand U345 (N_345,In_472,In_1789);
nor U346 (N_346,In_1849,In_1011);
xor U347 (N_347,N_100,In_237);
nor U348 (N_348,In_776,In_1908);
xnor U349 (N_349,In_1892,In_1475);
or U350 (N_350,In_546,N_63);
nand U351 (N_351,In_324,N_129);
and U352 (N_352,In_1876,In_214);
nand U353 (N_353,In_1815,In_624);
or U354 (N_354,In_1788,In_438);
nor U355 (N_355,In_1516,In_57);
or U356 (N_356,In_930,In_48);
or U357 (N_357,N_109,In_836);
nand U358 (N_358,In_508,In_1014);
xor U359 (N_359,In_1142,In_1584);
and U360 (N_360,In_1981,In_658);
or U361 (N_361,In_124,In_113);
or U362 (N_362,In_993,N_126);
xor U363 (N_363,In_1777,In_1835);
nand U364 (N_364,In_838,In_726);
nand U365 (N_365,In_1409,In_1045);
xor U366 (N_366,In_1977,In_1913);
xnor U367 (N_367,In_1214,In_1273);
nor U368 (N_368,In_421,N_159);
nand U369 (N_369,In_1265,N_170);
nand U370 (N_370,In_906,In_530);
nand U371 (N_371,In_468,In_1959);
xnor U372 (N_372,N_188,In_1639);
xor U373 (N_373,In_640,In_687);
xnor U374 (N_374,In_283,In_772);
nor U375 (N_375,In_379,In_385);
xnor U376 (N_376,In_1969,In_382);
nor U377 (N_377,In_1507,In_1036);
and U378 (N_378,In_663,In_333);
xnor U379 (N_379,In_65,In_536);
nand U380 (N_380,In_311,In_0);
nor U381 (N_381,In_940,In_1160);
and U382 (N_382,In_969,In_1953);
nand U383 (N_383,In_186,In_1591);
nand U384 (N_384,In_1301,In_523);
xor U385 (N_385,In_612,In_123);
nand U386 (N_386,In_1924,In_244);
nor U387 (N_387,In_408,N_96);
xnor U388 (N_388,In_1736,In_1217);
xnor U389 (N_389,In_312,In_172);
xnor U390 (N_390,In_861,In_672);
or U391 (N_391,In_892,In_1980);
and U392 (N_392,In_681,N_49);
and U393 (N_393,In_948,In_1186);
nand U394 (N_394,In_1422,In_537);
nand U395 (N_395,In_1850,In_199);
nor U396 (N_396,N_133,In_737);
nand U397 (N_397,In_1359,In_558);
nand U398 (N_398,N_24,In_889);
or U399 (N_399,In_1222,In_593);
or U400 (N_400,N_78,N_40);
nand U401 (N_401,N_130,N_378);
xnor U402 (N_402,In_814,In_467);
nand U403 (N_403,In_982,In_645);
xnor U404 (N_404,N_102,In_1582);
xor U405 (N_405,In_1468,In_1628);
xor U406 (N_406,N_376,In_238);
and U407 (N_407,N_237,In_531);
xor U408 (N_408,In_996,In_389);
xor U409 (N_409,In_825,N_62);
xnor U410 (N_410,In_424,In_920);
nand U411 (N_411,N_202,In_1149);
or U412 (N_412,In_943,In_1714);
nor U413 (N_413,In_1987,In_780);
and U414 (N_414,In_1430,In_443);
or U415 (N_415,In_1852,In_1335);
nand U416 (N_416,N_152,In_1292);
nor U417 (N_417,In_724,N_344);
and U418 (N_418,In_1644,In_706);
and U419 (N_419,N_392,In_1513);
and U420 (N_420,In_414,In_956);
xor U421 (N_421,In_1445,In_1599);
xnor U422 (N_422,In_1027,In_1795);
nor U423 (N_423,In_142,In_1000);
xor U424 (N_424,N_36,In_1982);
xnor U425 (N_425,N_268,In_790);
or U426 (N_426,In_1428,In_934);
or U427 (N_427,In_26,N_23);
nor U428 (N_428,In_1216,In_265);
nor U429 (N_429,N_215,N_192);
nor U430 (N_430,In_754,In_1);
nor U431 (N_431,In_521,In_185);
and U432 (N_432,In_1560,In_344);
and U433 (N_433,In_740,In_1962);
nor U434 (N_434,In_584,In_1275);
and U435 (N_435,N_59,In_731);
nor U436 (N_436,In_253,In_474);
nor U437 (N_437,In_852,In_486);
nand U438 (N_438,In_1201,In_1685);
or U439 (N_439,In_247,In_1322);
and U440 (N_440,N_231,In_1555);
nor U441 (N_441,In_1067,In_1282);
and U442 (N_442,In_217,In_758);
nand U443 (N_443,In_650,N_3);
xor U444 (N_444,In_1348,In_235);
nand U445 (N_445,In_1044,In_689);
or U446 (N_446,In_1676,In_1237);
or U447 (N_447,N_332,N_50);
or U448 (N_448,In_1632,In_403);
and U449 (N_449,In_1716,In_713);
and U450 (N_450,In_950,In_1643);
and U451 (N_451,In_651,In_215);
and U452 (N_452,In_1309,In_622);
or U453 (N_453,In_40,N_398);
and U454 (N_454,In_296,In_1646);
or U455 (N_455,In_96,In_1635);
xor U456 (N_456,In_453,In_1589);
xor U457 (N_457,In_1873,In_268);
and U458 (N_458,In_494,N_203);
xnor U459 (N_459,In_1269,In_227);
xor U460 (N_460,N_43,In_767);
nor U461 (N_461,In_1013,In_1747);
xnor U462 (N_462,N_31,N_397);
or U463 (N_463,In_1016,In_307);
nor U464 (N_464,In_1168,In_427);
xnor U465 (N_465,N_118,N_347);
nor U466 (N_466,In_42,In_441);
and U467 (N_467,In_1403,N_206);
and U468 (N_468,In_239,In_1673);
nor U469 (N_469,In_1068,In_1907);
and U470 (N_470,In_1349,N_263);
xor U471 (N_471,In_1101,N_374);
or U472 (N_472,In_1524,In_1900);
nand U473 (N_473,In_1473,In_1413);
xnor U474 (N_474,N_285,N_311);
and U475 (N_475,In_59,In_1844);
or U476 (N_476,In_901,N_352);
nand U477 (N_477,N_72,In_1642);
nand U478 (N_478,N_42,N_337);
xor U479 (N_479,In_392,In_964);
and U480 (N_480,In_960,N_175);
and U481 (N_481,In_1345,In_256);
nor U482 (N_482,In_1660,In_230);
xor U483 (N_483,N_339,N_81);
nand U484 (N_484,In_1726,In_1607);
xor U485 (N_485,In_1630,In_1715);
and U486 (N_486,N_37,N_314);
nand U487 (N_487,In_1459,In_965);
or U488 (N_488,In_1520,In_1249);
xnor U489 (N_489,In_1922,In_657);
nor U490 (N_490,In_966,In_842);
nor U491 (N_491,N_176,In_770);
or U492 (N_492,In_178,In_1927);
nand U493 (N_493,In_1761,In_959);
xnor U494 (N_494,In_503,In_118);
xnor U495 (N_495,In_1463,In_234);
or U496 (N_496,In_1272,In_1820);
or U497 (N_497,In_1246,In_1161);
nor U498 (N_498,In_1502,N_117);
nand U499 (N_499,In_999,In_725);
and U500 (N_500,In_1037,In_1424);
nand U501 (N_501,In_891,In_983);
nor U502 (N_502,In_1532,In_1097);
or U503 (N_503,In_614,In_1961);
and U504 (N_504,In_1548,N_51);
or U505 (N_505,In_1684,In_1979);
xnor U506 (N_506,In_1451,In_824);
nand U507 (N_507,In_29,N_229);
and U508 (N_508,In_1366,In_563);
nor U509 (N_509,In_1029,In_524);
and U510 (N_510,In_802,In_1125);
or U511 (N_511,In_1293,In_1474);
and U512 (N_512,In_1781,In_1566);
nor U513 (N_513,In_539,In_1239);
xor U514 (N_514,N_19,In_998);
nor U515 (N_515,N_334,In_1693);
nor U516 (N_516,N_18,In_775);
nor U517 (N_517,N_57,In_1402);
xor U518 (N_518,In_469,In_1340);
and U519 (N_519,In_600,In_1525);
xnor U520 (N_520,In_1109,In_1442);
or U521 (N_521,In_992,In_746);
and U522 (N_522,N_368,In_1412);
xnor U523 (N_523,In_1893,In_987);
nand U524 (N_524,In_28,In_855);
nor U525 (N_525,In_1658,In_1470);
and U526 (N_526,In_1357,In_1242);
and U527 (N_527,N_227,In_1759);
or U528 (N_528,In_1770,In_1437);
nand U529 (N_529,In_1738,N_381);
or U530 (N_530,N_138,In_1735);
xnor U531 (N_531,In_1128,N_279);
nor U532 (N_532,In_1400,In_1102);
or U533 (N_533,In_626,N_262);
xor U534 (N_534,In_712,N_380);
xor U535 (N_535,N_319,In_309);
nand U536 (N_536,In_512,In_1188);
xnor U537 (N_537,In_1052,In_1032);
and U538 (N_538,In_327,In_1654);
xnor U539 (N_539,In_974,N_209);
and U540 (N_540,In_800,In_881);
or U541 (N_541,In_290,In_325);
and U542 (N_542,In_18,In_222);
nand U543 (N_543,N_322,In_853);
or U544 (N_544,In_136,In_1381);
nand U545 (N_545,In_989,N_217);
nand U546 (N_546,N_281,In_1049);
nor U547 (N_547,In_949,In_1845);
nand U548 (N_548,In_1663,In_1072);
or U549 (N_549,N_234,In_1499);
or U550 (N_550,N_160,In_251);
or U551 (N_551,In_160,In_1457);
nand U552 (N_552,In_1905,In_1144);
or U553 (N_553,In_1783,In_867);
or U554 (N_554,In_431,In_1508);
nor U555 (N_555,In_1847,N_143);
nand U556 (N_556,In_1971,In_1666);
and U557 (N_557,In_1042,In_442);
nor U558 (N_558,In_1833,In_1600);
nor U559 (N_559,In_1346,In_581);
nand U560 (N_560,In_499,In_292);
nand U561 (N_561,In_1485,N_135);
nand U562 (N_562,N_4,In_1518);
and U563 (N_563,In_50,In_388);
nor U564 (N_564,N_253,In_1478);
or U565 (N_565,In_1286,In_1268);
xnor U566 (N_566,In_464,In_15);
and U567 (N_567,In_1421,In_1110);
or U568 (N_568,N_303,N_265);
nor U569 (N_569,N_146,N_257);
and U570 (N_570,In_1967,In_281);
and U571 (N_571,N_121,In_1528);
and U572 (N_572,In_1690,N_320);
xor U573 (N_573,N_167,N_247);
and U574 (N_574,In_1347,In_1098);
nand U575 (N_575,In_422,In_1059);
nand U576 (N_576,In_1806,In_1521);
nand U577 (N_577,In_73,N_35);
nor U578 (N_578,In_1933,N_318);
nand U579 (N_579,In_1248,N_286);
or U580 (N_580,N_189,In_907);
xnor U581 (N_581,N_55,In_106);
or U582 (N_582,In_1827,In_1910);
nand U583 (N_583,In_1816,N_137);
nand U584 (N_584,In_1408,In_542);
nor U585 (N_585,In_211,In_1010);
and U586 (N_586,In_876,In_1012);
xor U587 (N_587,In_1231,In_1920);
nor U588 (N_588,In_1537,In_498);
nand U589 (N_589,N_208,In_456);
nand U590 (N_590,N_399,In_200);
or U591 (N_591,N_114,In_1446);
and U592 (N_592,In_843,N_377);
and U593 (N_593,In_741,In_528);
or U594 (N_594,N_256,In_1709);
xnor U595 (N_595,In_1425,In_788);
nand U596 (N_596,In_1935,In_381);
xor U597 (N_597,In_721,N_224);
or U598 (N_598,In_152,N_331);
and U599 (N_599,In_1616,N_306);
and U600 (N_600,N_105,In_1662);
nand U601 (N_601,N_173,In_516);
nor U602 (N_602,N_157,In_1720);
nor U603 (N_603,In_212,In_1784);
xor U604 (N_604,In_680,N_298);
and U605 (N_605,In_1054,In_1138);
and U606 (N_606,In_871,In_10);
nor U607 (N_607,In_1719,In_1164);
nor U608 (N_608,N_302,N_475);
and U609 (N_609,In_1578,In_1100);
xnor U610 (N_610,In_1975,In_1414);
or U611 (N_611,In_492,In_1608);
nor U612 (N_612,N_364,In_1705);
nor U613 (N_613,In_529,In_87);
and U614 (N_614,In_1853,N_310);
or U615 (N_615,In_714,In_1942);
xnor U616 (N_616,In_291,In_1004);
nor U617 (N_617,In_1298,In_93);
nor U618 (N_618,In_924,In_1498);
nand U619 (N_619,N_115,In_473);
or U620 (N_620,In_207,In_1741);
xnor U621 (N_621,In_1148,In_566);
and U622 (N_622,In_1466,In_1252);
and U623 (N_623,In_153,In_286);
xor U624 (N_624,In_274,N_447);
or U625 (N_625,In_335,N_2);
nand U626 (N_626,In_1659,N_284);
xnor U627 (N_627,N_232,N_563);
and U628 (N_628,N_442,N_382);
xor U629 (N_629,In_1397,In_909);
nand U630 (N_630,In_401,N_597);
nand U631 (N_631,N_363,N_471);
nor U632 (N_632,In_419,In_1080);
or U633 (N_633,N_94,In_1681);
and U634 (N_634,In_656,In_1378);
or U635 (N_635,N_266,N_74);
xnor U636 (N_636,In_1978,In_1399);
or U637 (N_637,In_1577,In_243);
xor U638 (N_638,N_505,In_1223);
nand U639 (N_639,N_367,N_431);
xor U640 (N_640,N_304,In_1620);
xor U641 (N_641,In_1734,N_570);
and U642 (N_642,In_1657,In_1433);
and U643 (N_643,In_1244,N_239);
nor U644 (N_644,In_1647,In_1453);
and U645 (N_645,In_301,In_926);
xor U646 (N_646,In_1171,In_1240);
xor U647 (N_647,In_1364,In_522);
xor U648 (N_648,In_1964,N_69);
nand U649 (N_649,N_521,In_1626);
and U650 (N_650,In_31,In_1559);
nor U651 (N_651,In_981,N_558);
xnor U652 (N_652,In_353,In_451);
or U653 (N_653,N_255,N_585);
nor U654 (N_654,In_1818,In_1768);
or U655 (N_655,In_1544,N_574);
nand U656 (N_656,In_1653,In_534);
nor U657 (N_657,N_204,In_490);
and U658 (N_658,N_271,In_1199);
or U659 (N_659,In_246,In_1567);
xor U660 (N_660,In_809,In_1274);
or U661 (N_661,In_1609,In_112);
xnor U662 (N_662,In_1025,In_595);
nor U663 (N_663,In_175,In_1061);
xnor U664 (N_664,In_962,N_372);
or U665 (N_665,In_479,In_1984);
or U666 (N_666,In_533,In_860);
nor U667 (N_667,N_250,N_87);
xor U668 (N_668,N_321,N_139);
and U669 (N_669,In_66,In_139);
or U670 (N_670,In_390,In_1842);
and U671 (N_671,N_0,In_1743);
or U672 (N_672,N_540,In_1570);
nand U673 (N_673,N_422,In_840);
nor U674 (N_674,In_1183,In_1808);
nor U675 (N_675,In_470,In_1193);
and U676 (N_676,In_1375,In_2);
nand U677 (N_677,N_421,In_229);
or U678 (N_678,In_565,In_1341);
xor U679 (N_679,N_415,N_200);
and U680 (N_680,N_32,N_269);
nor U681 (N_681,N_389,In_1197);
nand U682 (N_682,N_350,In_1755);
and U683 (N_683,In_1533,N_424);
nand U684 (N_684,In_1465,N_267);
nor U685 (N_685,In_1557,In_254);
xnor U686 (N_686,In_127,In_425);
nand U687 (N_687,N_65,In_491);
nand U688 (N_688,In_191,In_105);
nand U689 (N_689,N_577,N_395);
and U690 (N_690,In_376,N_532);
and U691 (N_691,In_1604,In_1296);
or U692 (N_692,N_592,In_1449);
xor U693 (N_693,N_459,In_967);
xor U694 (N_694,In_1136,In_1344);
nor U695 (N_695,N_572,In_30);
and U696 (N_696,In_732,In_358);
and U697 (N_697,In_115,In_1786);
nand U698 (N_698,In_101,N_233);
or U699 (N_699,N_299,In_509);
or U700 (N_700,In_938,N_328);
xor U701 (N_701,In_829,In_1860);
or U702 (N_702,N_457,N_405);
nor U703 (N_703,In_463,In_1205);
or U704 (N_704,In_1901,In_1510);
nor U705 (N_705,N_343,In_1943);
nor U706 (N_706,In_447,In_1800);
nor U707 (N_707,In_1129,In_1215);
nand U708 (N_708,In_854,In_308);
and U709 (N_709,N_477,In_812);
nor U710 (N_710,In_255,In_1260);
and U711 (N_711,N_68,In_1419);
xor U712 (N_712,N_30,In_1751);
nor U713 (N_713,In_1881,In_225);
xnor U714 (N_714,In_1377,In_839);
xor U715 (N_715,N_258,In_1135);
nor U716 (N_716,N_305,N_385);
nand U717 (N_717,In_675,N_323);
xnor U718 (N_718,N_274,In_1722);
xnor U719 (N_719,N_125,In_1001);
nor U720 (N_720,In_1701,N_482);
and U721 (N_721,In_1650,In_1090);
xor U722 (N_722,N_168,N_439);
or U723 (N_723,In_111,In_1084);
or U724 (N_724,In_902,In_1388);
and U725 (N_725,N_226,N_536);
nand U726 (N_726,In_769,In_835);
xnor U727 (N_727,N_409,In_1074);
and U728 (N_728,In_1634,N_243);
nor U729 (N_729,In_1184,N_197);
xor U730 (N_730,N_312,In_126);
nand U731 (N_731,N_503,In_977);
nand U732 (N_732,In_1178,In_317);
and U733 (N_733,In_1447,In_547);
or U734 (N_734,In_868,N_446);
and U735 (N_735,N_449,N_245);
nand U736 (N_736,In_276,N_85);
nand U737 (N_737,In_1579,N_366);
or U738 (N_738,In_1363,In_1837);
or U739 (N_739,In_1527,In_1898);
nand U740 (N_740,In_1778,In_44);
nor U741 (N_741,In_1995,In_1393);
or U742 (N_742,In_1864,N_526);
or U743 (N_743,In_1811,In_1325);
nand U744 (N_744,N_199,In_1955);
or U745 (N_745,In_1834,In_1688);
or U746 (N_746,In_1787,In_579);
nor U747 (N_747,In_583,In_1139);
nor U748 (N_748,N_73,N_163);
nor U749 (N_749,In_1022,In_1749);
and U750 (N_750,In_1460,N_333);
nor U751 (N_751,N_70,N_591);
or U752 (N_752,In_493,N_162);
and U753 (N_753,N_83,In_933);
and U754 (N_754,N_564,In_1489);
nor U755 (N_755,N_66,N_444);
nor U756 (N_756,In_1514,N_492);
or U757 (N_757,N_460,In_1181);
and U758 (N_758,N_153,N_598);
xnor U759 (N_759,In_1763,N_487);
and U760 (N_760,N_433,In_1874);
nand U761 (N_761,In_679,N_441);
and U762 (N_762,In_300,N_512);
nor U763 (N_763,In_1350,In_1115);
nor U764 (N_764,In_147,In_1748);
or U765 (N_765,N_147,N_194);
or U766 (N_766,N_354,N_466);
nor U767 (N_767,In_170,N_565);
nor U768 (N_768,In_155,In_697);
and U769 (N_769,In_1355,In_373);
or U770 (N_770,N_533,In_1610);
xor U771 (N_771,N_1,In_873);
xor U772 (N_772,In_1764,In_89);
xor U773 (N_773,In_1119,In_1993);
nor U774 (N_774,N_236,In_1229);
nand U775 (N_775,N_8,In_122);
and U776 (N_776,In_718,In_1267);
xnor U777 (N_777,In_1989,N_329);
nor U778 (N_778,In_908,N_348);
nand U779 (N_779,In_1585,In_343);
or U780 (N_780,In_1594,In_1305);
and U781 (N_781,In_1360,N_365);
or U782 (N_782,In_446,In_1065);
xnor U783 (N_783,In_1411,In_36);
nor U784 (N_784,In_54,In_8);
and U785 (N_785,In_1802,N_166);
nor U786 (N_786,In_674,N_293);
and U787 (N_787,N_413,In_574);
nand U788 (N_788,In_602,N_556);
nand U789 (N_789,In_345,N_596);
nand U790 (N_790,In_1613,In_1552);
nand U791 (N_791,In_1886,In_903);
xor U792 (N_792,N_404,In_1563);
or U793 (N_793,N_593,N_506);
and U794 (N_794,In_411,In_1117);
nand U795 (N_795,N_92,In_1256);
nor U796 (N_796,N_357,In_785);
or U797 (N_797,In_1415,In_476);
xor U798 (N_798,In_216,In_1652);
nand U799 (N_799,N_288,In_1213);
nor U800 (N_800,N_713,In_1443);
xor U801 (N_801,In_1821,In_1791);
and U802 (N_802,N_17,N_718);
nand U803 (N_803,In_12,N_587);
nand U804 (N_804,In_68,In_1224);
or U805 (N_805,In_1580,N_498);
xor U806 (N_806,N_275,N_60);
nor U807 (N_807,In_16,In_556);
xnor U808 (N_808,In_35,In_1882);
xnor U809 (N_809,In_1885,N_693);
xnor U810 (N_810,N_552,In_1556);
or U811 (N_811,In_79,N_467);
or U812 (N_812,In_285,In_1529);
or U813 (N_813,N_733,In_734);
and U814 (N_814,In_676,N_756);
nand U815 (N_815,N_703,N_220);
nor U816 (N_816,N_691,In_942);
xnor U817 (N_817,In_1324,In_1517);
nor U818 (N_818,In_1187,N_360);
or U819 (N_819,In_1472,In_1573);
or U820 (N_820,In_1368,In_1427);
and U821 (N_821,N_108,In_605);
xnor U822 (N_822,N_681,N_359);
nor U823 (N_823,In_1123,N_644);
and U824 (N_824,In_168,N_662);
or U825 (N_825,N_517,In_395);
and U826 (N_826,N_799,In_95);
nand U827 (N_827,In_223,In_94);
or U828 (N_828,N_649,N_641);
xor U829 (N_829,N_14,In_750);
xor U830 (N_830,N_595,N_426);
or U831 (N_831,N_425,In_1572);
xnor U832 (N_832,N_289,In_905);
or U833 (N_833,N_655,In_562);
or U834 (N_834,In_193,In_863);
nor U835 (N_835,N_346,N_416);
nor U836 (N_836,N_648,In_165);
and U837 (N_837,N_538,N_316);
xnor U838 (N_838,In_39,In_1417);
nand U839 (N_839,In_803,In_1220);
or U840 (N_840,In_1058,In_919);
nor U841 (N_841,In_179,N_155);
or U842 (N_842,N_193,In_1602);
or U843 (N_843,N_185,In_1236);
and U844 (N_844,In_86,N_182);
nand U845 (N_845,N_796,In_1615);
or U846 (N_846,In_786,In_578);
or U847 (N_847,N_93,In_576);
and U848 (N_848,In_1291,N_762);
xor U849 (N_849,In_1569,N_551);
or U850 (N_850,N_676,In_250);
or U851 (N_851,In_1406,In_878);
nand U852 (N_852,N_684,In_1203);
nand U853 (N_853,N_715,N_610);
or U854 (N_854,In_513,N_632);
or U855 (N_855,In_1407,N_722);
nand U856 (N_856,In_1276,N_575);
or U857 (N_857,In_334,N_615);
and U858 (N_858,In_592,N_119);
or U859 (N_859,N_753,N_777);
nor U860 (N_860,In_314,In_1111);
xnor U861 (N_861,In_1328,N_504);
or U862 (N_862,N_29,N_391);
and U863 (N_863,N_480,In_690);
and U864 (N_864,In_1590,In_1353);
or U865 (N_865,N_735,In_707);
nand U866 (N_866,In_1405,In_682);
and U867 (N_867,In_1031,In_208);
and U868 (N_868,In_1198,In_146);
or U869 (N_869,In_1081,N_127);
nor U870 (N_870,N_628,N_455);
and U871 (N_871,In_1970,In_278);
and U872 (N_872,In_970,N_520);
xor U873 (N_873,In_1703,In_722);
nor U874 (N_874,In_1598,In_1637);
nand U875 (N_875,In_1096,In_601);
xnor U876 (N_876,N_34,In_310);
nor U877 (N_877,N_349,In_606);
or U878 (N_878,In_1038,N_625);
xnor U879 (N_879,In_1804,N_680);
nor U880 (N_880,N_573,In_947);
xor U881 (N_881,N_154,In_550);
nand U882 (N_882,N_158,In_1782);
nor U883 (N_883,In_1668,N_402);
nand U884 (N_884,In_994,N_476);
or U885 (N_885,N_531,In_130);
nand U886 (N_886,N_97,In_25);
or U887 (N_887,In_985,In_627);
and U888 (N_888,In_104,In_1817);
nand U889 (N_889,N_307,In_497);
xnor U890 (N_890,N_790,In_735);
or U891 (N_891,In_70,N_412);
nand U892 (N_892,N_9,N_527);
nor U893 (N_893,In_912,In_1077);
nand U894 (N_894,N_774,N_379);
and U895 (N_895,In_3,In_827);
and U896 (N_896,N_423,In_257);
nand U897 (N_897,In_1692,N_786);
nand U898 (N_898,N_210,N_340);
or U899 (N_899,In_709,N_356);
nor U900 (N_900,N_736,N_618);
nor U901 (N_901,In_1336,In_945);
xnor U902 (N_902,In_893,In_793);
or U903 (N_903,N_657,N_580);
nand U904 (N_904,N_16,In_410);
or U905 (N_905,In_1762,N_5);
xnor U906 (N_906,In_1543,N_132);
nand U907 (N_907,N_779,N_671);
xor U908 (N_908,In_51,In_197);
nor U909 (N_909,In_759,In_1172);
and U910 (N_910,In_1122,N_324);
xnor U911 (N_911,In_74,In_98);
nor U912 (N_912,In_82,In_798);
xor U913 (N_913,In_815,N_260);
xnor U914 (N_914,In_887,N_164);
and U915 (N_915,In_1672,In_1380);
nor U916 (N_916,In_729,In_1255);
nor U917 (N_917,N_282,In_1588);
xor U918 (N_918,In_263,In_187);
and U919 (N_919,In_357,N_683);
nand U920 (N_920,N_555,N_605);
or U921 (N_921,In_306,In_1790);
and U922 (N_922,N_261,N_327);
nor U923 (N_923,In_988,In_1155);
nor U924 (N_924,N_702,In_56);
nor U925 (N_925,In_1374,In_1137);
nor U926 (N_926,N_99,In_1243);
and U927 (N_927,In_946,In_1207);
nand U928 (N_928,In_448,In_1742);
nand U929 (N_929,In_859,In_496);
or U930 (N_930,In_92,In_972);
nand U931 (N_931,In_1112,In_931);
nor U932 (N_932,In_457,In_418);
or U933 (N_933,In_1303,N_700);
nand U934 (N_934,In_1623,N_741);
or U935 (N_935,N_524,N_623);
or U936 (N_936,In_69,In_439);
nand U937 (N_937,In_1271,N_39);
and U938 (N_938,In_1277,In_1538);
xor U939 (N_939,N_694,N_643);
nor U940 (N_940,In_1879,In_369);
and U941 (N_941,In_294,N_15);
or U942 (N_942,N_669,In_1176);
nor U943 (N_943,In_233,N_769);
xnor U944 (N_944,N_745,In_1890);
nor U945 (N_945,In_1840,N_218);
or U946 (N_946,In_749,In_347);
nand U947 (N_947,In_526,N_629);
nor U948 (N_948,N_510,In_1085);
or U949 (N_949,N_534,N_513);
xnor U950 (N_950,N_342,In_1418);
nor U951 (N_951,In_915,N_734);
or U952 (N_952,In_744,N_546);
xnor U953 (N_953,In_1270,N_291);
xnor U954 (N_954,In_1721,N_528);
or U955 (N_955,N_583,N_584);
nand U956 (N_956,In_273,N_544);
and U957 (N_957,In_1019,N_468);
nor U958 (N_958,In_1866,In_1575);
xnor U959 (N_959,N_488,N_586);
nand U960 (N_960,N_670,In_326);
nand U961 (N_961,In_882,In_289);
and U962 (N_962,In_834,In_745);
nand U963 (N_963,In_518,N_493);
nor U964 (N_964,In_1941,In_1150);
nor U965 (N_965,In_1389,In_874);
nor U966 (N_966,In_619,N_473);
or U967 (N_967,In_1998,In_1232);
nand U968 (N_968,N_228,In_303);
nand U969 (N_969,N_317,In_1903);
nor U970 (N_970,In_1423,In_596);
or U971 (N_971,N_622,N_485);
and U972 (N_972,In_1354,N_766);
xor U973 (N_973,In_1558,In_848);
xnor U974 (N_974,In_1895,In_1095);
or U975 (N_975,In_1263,N_549);
or U976 (N_976,N_417,In_1771);
xnor U977 (N_977,In_1329,N_726);
or U978 (N_978,N_249,N_252);
xnor U979 (N_979,N_561,In_1838);
or U980 (N_980,In_4,N_752);
xor U981 (N_981,In_484,In_866);
nor U982 (N_982,N_780,N_338);
xor U983 (N_983,In_1823,N_278);
xor U984 (N_984,In_1157,In_917);
nor U985 (N_985,In_1695,In_1210);
nor U986 (N_986,N_666,In_1926);
or U987 (N_987,In_1230,N_47);
xor U988 (N_988,N_207,N_633);
nor U989 (N_989,In_1750,N_499);
nor U990 (N_990,In_1130,N_198);
and U991 (N_991,In_978,In_723);
xor U992 (N_992,In_1949,In_1679);
nor U993 (N_993,N_71,N_754);
or U994 (N_994,In_1234,In_1285);
nor U995 (N_995,N_682,N_113);
nand U996 (N_996,N_205,In_609);
xnor U997 (N_997,In_1392,N_438);
nand U998 (N_998,In_693,N_674);
nand U999 (N_999,In_937,In_957);
nor U1000 (N_1000,N_469,N_812);
or U1001 (N_1001,N_969,N_82);
nor U1002 (N_1002,In_666,N_128);
and U1003 (N_1003,N_880,N_933);
or U1004 (N_1004,N_386,In_1104);
or U1005 (N_1005,In_505,In_41);
nand U1006 (N_1006,In_260,In_297);
and U1007 (N_1007,In_1713,N_495);
and U1008 (N_1008,In_1656,N_984);
nand U1009 (N_1009,N_246,In_1622);
or U1010 (N_1010,N_695,N_839);
nor U1011 (N_1011,In_553,N_867);
or U1012 (N_1012,N_946,N_778);
nand U1013 (N_1013,N_659,N_893);
nand U1014 (N_1014,N_743,In_755);
nor U1015 (N_1015,In_639,In_830);
xor U1016 (N_1016,N_960,In_151);
nand U1017 (N_1017,In_1991,N_191);
and U1018 (N_1018,In_688,In_384);
and U1019 (N_1019,In_973,N_470);
nor U1020 (N_1020,N_248,In_149);
xor U1021 (N_1021,N_362,N_481);
xnor U1022 (N_1022,N_678,In_271);
nor U1023 (N_1023,N_773,In_1678);
xor U1024 (N_1024,N_272,N_761);
and U1025 (N_1025,In_1432,N_437);
and U1026 (N_1026,N_901,N_971);
and U1027 (N_1027,N_111,N_959);
nor U1028 (N_1028,N_180,N_637);
or U1029 (N_1029,In_527,N_353);
xor U1030 (N_1030,N_923,In_475);
and U1031 (N_1031,N_994,N_788);
nand U1032 (N_1032,N_917,N_723);
xor U1033 (N_1033,N_67,In_1476);
xnor U1034 (N_1034,N_223,N_427);
or U1035 (N_1035,N_836,In_1871);
nor U1036 (N_1036,In_1564,N_808);
xor U1037 (N_1037,In_1120,In_1928);
xnor U1038 (N_1038,N_711,In_1797);
xnor U1039 (N_1039,In_1158,N_667);
xor U1040 (N_1040,N_907,N_709);
and U1041 (N_1041,In_1896,In_520);
or U1042 (N_1042,In_387,In_801);
or U1043 (N_1043,N_747,In_703);
nand U1044 (N_1044,N_496,N_647);
nor U1045 (N_1045,N_948,In_372);
nand U1046 (N_1046,N_932,In_1756);
or U1047 (N_1047,N_451,N_95);
or U1048 (N_1048,N_860,N_908);
xnor U1049 (N_1049,N_461,N_991);
nand U1050 (N_1050,In_1066,In_728);
nor U1051 (N_1051,N_749,N_704);
nor U1052 (N_1052,N_483,In_1030);
or U1053 (N_1053,N_730,In_1279);
and U1054 (N_1054,In_145,N_494);
nand U1055 (N_1055,N_842,N_956);
xnor U1056 (N_1056,N_920,In_535);
xnor U1057 (N_1057,N_934,In_154);
xnor U1058 (N_1058,N_751,In_402);
nand U1059 (N_1059,N_484,N_689);
nand U1060 (N_1060,In_1320,In_14);
xor U1061 (N_1061,N_589,N_793);
xnor U1062 (N_1062,N_539,In_805);
xnor U1063 (N_1063,N_77,N_620);
xnor U1064 (N_1064,N_530,In_833);
nand U1065 (N_1065,N_975,In_603);
nor U1066 (N_1066,In_910,N_668);
or U1067 (N_1067,N_296,N_491);
xor U1068 (N_1068,In_171,N_846);
nand U1069 (N_1069,N_898,N_394);
or U1070 (N_1070,In_1062,N_955);
nand U1071 (N_1071,In_1050,In_1667);
xor U1072 (N_1072,In_1851,N_783);
nand U1073 (N_1073,N_813,N_835);
nor U1074 (N_1074,N_336,In_1775);
nor U1075 (N_1075,In_1919,N_732);
nand U1076 (N_1076,N_650,In_1831);
xnor U1077 (N_1077,N_48,In_365);
nor U1078 (N_1078,In_857,N_988);
nand U1079 (N_1079,N_878,N_887);
or U1080 (N_1080,N_914,In_218);
xor U1081 (N_1081,In_397,In_99);
or U1082 (N_1082,N_918,In_1327);
or U1083 (N_1083,N_748,N_962);
xor U1084 (N_1084,N_993,In_1530);
nor U1085 (N_1085,In_730,N_420);
xor U1086 (N_1086,N_183,In_287);
nand U1087 (N_1087,N_864,In_900);
nand U1088 (N_1088,N_807,N_952);
xnor U1089 (N_1089,N_829,In_585);
and U1090 (N_1090,N_213,N_961);
or U1091 (N_1091,In_1829,In_1133);
and U1092 (N_1092,N_817,N_792);
xor U1093 (N_1093,N_140,N_837);
and U1094 (N_1094,In_611,In_37);
xnor U1095 (N_1095,N_631,N_883);
nor U1096 (N_1096,N_844,N_161);
xnor U1097 (N_1097,In_1503,In_489);
or U1098 (N_1098,In_670,N_98);
nand U1099 (N_1099,N_978,N_881);
nand U1100 (N_1100,In_1728,N_937);
xnor U1101 (N_1101,N_222,N_912);
or U1102 (N_1102,In_506,N_760);
xor U1103 (N_1103,In_1985,In_1753);
or U1104 (N_1104,In_1440,In_58);
nand U1105 (N_1105,In_589,N_462);
and U1106 (N_1106,In_517,In_1254);
nand U1107 (N_1107,In_826,N_822);
xor U1108 (N_1108,N_273,In_159);
and U1109 (N_1109,N_612,In_820);
xnor U1110 (N_1110,In_1906,N_560);
nor U1111 (N_1111,N_295,In_1410);
nand U1112 (N_1112,In_194,In_1429);
nor U1113 (N_1113,In_762,N_781);
nor U1114 (N_1114,In_406,In_1338);
nor U1115 (N_1115,In_190,In_298);
and U1116 (N_1116,In_916,In_1824);
nor U1117 (N_1117,In_416,In_1196);
and U1118 (N_1118,N_400,In_1469);
nor U1119 (N_1119,N_985,N_201);
and U1120 (N_1120,N_654,N_64);
xor U1121 (N_1121,In_1911,N_134);
nand U1122 (N_1122,N_982,N_904);
and U1123 (N_1123,In_1284,N_606);
or U1124 (N_1124,N_297,N_673);
nor U1125 (N_1125,N_464,N_885);
xor U1126 (N_1126,In_483,In_739);
and U1127 (N_1127,N_873,N_696);
and U1128 (N_1128,N_672,In_1633);
nand U1129 (N_1129,N_862,In_1386);
nor U1130 (N_1130,N_785,N_568);
or U1131 (N_1131,N_557,In_102);
and U1132 (N_1132,N_708,In_1805);
xnor U1133 (N_1133,N_675,In_341);
and U1134 (N_1134,In_597,N_841);
xor U1135 (N_1135,N_627,In_84);
xnor U1136 (N_1136,In_478,N_906);
nand U1137 (N_1137,N_264,N_519);
nor U1138 (N_1138,N_550,N_225);
nor U1139 (N_1139,In_444,In_1209);
nor U1140 (N_1140,N_945,N_315);
and U1141 (N_1141,N_103,In_1724);
and U1142 (N_1142,In_1384,N_393);
and U1143 (N_1143,In_738,N_686);
nand U1144 (N_1144,In_1540,N_514);
nand U1145 (N_1145,N_621,In_282);
xnor U1146 (N_1146,In_426,In_877);
and U1147 (N_1147,N_953,In_1772);
and U1148 (N_1148,N_782,In_761);
nor U1149 (N_1149,In_789,N_515);
nor U1150 (N_1150,N_106,In_577);
xor U1151 (N_1151,N_891,In_1456);
or U1152 (N_1152,In_49,In_661);
xor U1153 (N_1153,N_770,In_1550);
and U1154 (N_1154,N_849,N_26);
nand U1155 (N_1155,N_803,In_1092);
or U1156 (N_1156,N_635,In_363);
nand U1157 (N_1157,N_501,In_1055);
nor U1158 (N_1158,N_652,In_1754);
nand U1159 (N_1159,In_1091,N_687);
nor U1160 (N_1160,In_1495,N_942);
and U1161 (N_1161,N_924,In_1512);
nand U1162 (N_1162,N_458,N_235);
and U1163 (N_1163,N_905,In_284);
nand U1164 (N_1164,N_931,N_401);
nand U1165 (N_1165,N_868,In_1917);
nor U1166 (N_1166,N_169,In_819);
xnor U1167 (N_1167,N_740,N_679);
xor U1168 (N_1168,N_765,N_802);
xnor U1169 (N_1169,N_848,In_330);
or U1170 (N_1170,In_83,In_1094);
nor U1171 (N_1171,N_634,In_1299);
xnor U1172 (N_1172,N_351,In_1614);
and U1173 (N_1173,N_825,In_1034);
and U1174 (N_1174,In_487,In_1462);
or U1175 (N_1175,N_866,In_554);
and U1176 (N_1176,In_1576,In_1706);
nand U1177 (N_1177,N_986,N_661);
nor U1178 (N_1178,N_877,N_889);
and U1179 (N_1179,In_1391,N_731);
and U1180 (N_1180,N_280,N_916);
nor U1181 (N_1181,In_939,In_1390);
nor U1182 (N_1182,N_214,N_388);
or U1183 (N_1183,N_56,In_1003);
xnor U1184 (N_1184,N_411,N_928);
xnor U1185 (N_1185,N_710,In_557);
or U1186 (N_1186,In_677,In_485);
or U1187 (N_1187,N_525,N_238);
and U1188 (N_1188,N_995,In_796);
nor U1189 (N_1189,N_190,In_1127);
and U1190 (N_1190,In_777,In_911);
xnor U1191 (N_1191,N_358,N_452);
nand U1192 (N_1192,In_667,N_454);
nor U1193 (N_1193,N_576,N_645);
xor U1194 (N_1194,In_458,N_757);
and U1195 (N_1195,N_478,In_220);
nor U1196 (N_1196,N_863,In_623);
nor U1197 (N_1197,In_1611,N_436);
or U1198 (N_1198,N_896,N_996);
nor U1199 (N_1199,In_1603,N_857);
nand U1200 (N_1200,In_264,N_720);
or U1201 (N_1201,In_615,In_1867);
or U1202 (N_1202,In_1493,In_371);
nor U1203 (N_1203,N_1114,N_1142);
xor U1204 (N_1204,In_716,In_1723);
and U1205 (N_1205,N_390,N_1089);
nor U1206 (N_1206,In_1999,In_1825);
xor U1207 (N_1207,N_1141,N_746);
xnor U1208 (N_1208,N_1097,N_888);
xnor U1209 (N_1209,N_1170,N_1162);
nor U1210 (N_1210,N_828,N_1180);
and U1211 (N_1211,N_212,N_479);
xnor U1212 (N_1212,N_716,In_569);
nor U1213 (N_1213,N_1083,N_1165);
nand U1214 (N_1214,In_1661,N_1085);
or U1215 (N_1215,N_1077,N_290);
nor U1216 (N_1216,N_838,In_1861);
nand U1217 (N_1217,N_1066,N_403);
xnor U1218 (N_1218,N_764,In_813);
nor U1219 (N_1219,N_692,N_899);
xor U1220 (N_1220,N_518,N_805);
xnor U1221 (N_1221,N_970,In_1167);
xor U1222 (N_1222,In_128,In_540);
and U1223 (N_1223,N_1185,N_472);
nand U1224 (N_1224,N_859,In_1904);
nor U1225 (N_1225,N_820,N_1020);
nand U1226 (N_1226,In_1416,In_849);
and U1227 (N_1227,N_1104,In_1696);
or U1228 (N_1228,N_972,N_88);
xor U1229 (N_1229,N_1163,N_313);
nand U1230 (N_1230,N_958,N_1171);
or U1231 (N_1231,N_1005,In_1302);
xor U1232 (N_1232,In_141,In_1796);
nor U1233 (N_1233,In_1225,N_1139);
xor U1234 (N_1234,In_1841,N_1011);
nor U1235 (N_1235,In_1307,In_856);
xnor U1236 (N_1236,N_843,N_1055);
nor U1237 (N_1237,N_1183,N_1161);
and U1238 (N_1238,N_784,In_752);
nor U1239 (N_1239,N_992,In_1698);
and U1240 (N_1240,In_231,N_755);
and U1241 (N_1241,N_806,N_1145);
nand U1242 (N_1242,In_78,In_1491);
and U1243 (N_1243,N_432,N_1198);
or U1244 (N_1244,In_1467,In_77);
and U1245 (N_1245,In_1869,In_1023);
nor U1246 (N_1246,N_974,N_856);
or U1247 (N_1247,N_599,N_938);
or U1248 (N_1248,N_345,N_690);
or U1249 (N_1249,N_283,In_1297);
or U1250 (N_1250,In_1057,N_221);
nor U1251 (N_1251,In_914,In_91);
nor U1252 (N_1252,N_759,N_309);
and U1253 (N_1253,In_1593,N_818);
nor U1254 (N_1254,N_142,In_1106);
xnor U1255 (N_1255,N_1111,N_450);
and U1256 (N_1256,N_706,In_103);
nand U1257 (N_1257,In_1929,N_897);
or U1258 (N_1258,In_1318,N_375);
nand U1259 (N_1259,N_816,N_964);
or U1260 (N_1260,N_594,In_958);
nor U1261 (N_1261,N_1025,N_1186);
nand U1262 (N_1262,In_88,N_1168);
nand U1263 (N_1263,N_892,N_537);
xor U1264 (N_1264,N_474,N_832);
xnor U1265 (N_1265,N_172,In_869);
nand U1266 (N_1266,N_913,N_600);
nand U1267 (N_1267,N_1102,N_875);
xor U1268 (N_1268,N_1127,N_727);
nand U1269 (N_1269,N_1043,N_847);
and U1270 (N_1270,N_941,N_1042);
and U1271 (N_1271,In_678,In_701);
xnor U1272 (N_1272,N_511,N_602);
and U1273 (N_1273,In_779,N_369);
or U1274 (N_1274,In_837,N_1175);
nand U1275 (N_1275,N_911,N_1048);
or U1276 (N_1276,N_486,N_719);
or U1277 (N_1277,In_1361,N_601);
nand U1278 (N_1278,N_1080,In_125);
and U1279 (N_1279,N_771,N_824);
and U1280 (N_1280,N_1092,In_629);
nand U1281 (N_1281,In_665,N_639);
and U1282 (N_1282,N_171,N_325);
and U1283 (N_1283,N_815,N_131);
nor U1284 (N_1284,N_1129,In_428);
or U1285 (N_1285,N_187,In_1740);
xor U1286 (N_1286,N_1110,In_38);
nand U1287 (N_1287,N_1156,In_1617);
nand U1288 (N_1288,In_378,In_590);
and U1289 (N_1289,N_614,N_1035);
nor U1290 (N_1290,N_581,In_1976);
and U1291 (N_1291,N_890,In_1568);
xnor U1292 (N_1292,In_316,In_1694);
nand U1293 (N_1293,In_781,N_1063);
and U1294 (N_1294,In_482,N_407);
nor U1295 (N_1295,N_300,In_319);
nand U1296 (N_1296,In_1729,N_604);
xor U1297 (N_1297,N_1000,N_211);
xor U1298 (N_1298,In_1765,N_701);
or U1299 (N_1299,In_1915,In_132);
and U1300 (N_1300,N_1118,N_707);
nor U1301 (N_1301,N_922,In_1448);
nor U1302 (N_1302,N_1182,N_1058);
xnor U1303 (N_1303,N_1086,N_1017);
xor U1304 (N_1304,N_851,In_719);
xnor U1305 (N_1305,N_1027,In_213);
xor U1306 (N_1306,N_638,N_677);
nor U1307 (N_1307,N_1196,N_1113);
nand U1308 (N_1308,N_882,N_1046);
nand U1309 (N_1309,In_643,N_535);
nor U1310 (N_1310,N_950,In_621);
or U1311 (N_1311,In_1082,N_562);
or U1312 (N_1312,N_1140,N_244);
xor U1313 (N_1313,N_1103,N_789);
nor U1314 (N_1314,In_1053,In_1479);
xor U1315 (N_1315,N_1049,In_337);
xor U1316 (N_1316,In_1086,In_510);
or U1317 (N_1317,In_625,N_1194);
and U1318 (N_1318,N_724,N_1169);
nor U1319 (N_1319,In_1940,N_965);
or U1320 (N_1320,In_971,N_590);
nand U1321 (N_1321,N_903,N_737);
nor U1322 (N_1322,In_1947,N_489);
and U1323 (N_1323,N_840,N_1166);
nor U1324 (N_1324,N_456,N_1018);
and U1325 (N_1325,N_1044,N_1052);
nand U1326 (N_1326,N_61,N_981);
xnor U1327 (N_1327,In_1645,In_362);
and U1328 (N_1328,N_714,N_1028);
nand U1329 (N_1329,In_1026,N_1149);
and U1330 (N_1330,In_636,N_254);
nor U1331 (N_1331,N_46,In_1154);
nand U1332 (N_1332,N_1117,N_819);
or U1333 (N_1333,N_1130,In_1152);
nand U1334 (N_1334,In_1287,N_241);
and U1335 (N_1335,In_1621,N_1187);
and U1336 (N_1336,N_144,N_373);
and U1337 (N_1337,In_1546,N_276);
and U1338 (N_1338,In_205,In_1373);
and U1339 (N_1339,N_1034,N_430);
nand U1340 (N_1340,N_301,In_432);
nor U1341 (N_1341,N_418,N_1021);
xor U1342 (N_1342,In_1189,N_588);
xnor U1343 (N_1343,In_757,In_806);
xnor U1344 (N_1344,N_826,N_578);
and U1345 (N_1345,In_1766,In_1745);
or U1346 (N_1346,N_553,N_925);
nand U1347 (N_1347,N_833,N_463);
xor U1348 (N_1348,N_251,N_939);
or U1349 (N_1349,N_980,N_636);
xor U1350 (N_1350,In_628,In_1996);
or U1351 (N_1351,N_915,N_1024);
nor U1352 (N_1352,N_797,N_1096);
nor U1353 (N_1353,In_885,In_797);
nor U1354 (N_1354,N_930,N_651);
xor U1355 (N_1355,N_926,In_1854);
nor U1356 (N_1356,N_1056,N_1015);
xnor U1357 (N_1357,In_1228,In_1857);
xor U1358 (N_1358,N_497,In_1404);
and U1359 (N_1359,N_853,N_1061);
or U1360 (N_1360,N_811,N_1152);
and U1361 (N_1361,In_195,N_640);
and U1362 (N_1362,In_747,N_947);
and U1363 (N_1363,In_481,N_1167);
xor U1364 (N_1364,N_571,N_886);
nand U1365 (N_1365,N_775,In_1760);
or U1366 (N_1366,N_1131,In_206);
nand U1367 (N_1367,In_24,N_1075);
or U1368 (N_1368,In_1173,N_768);
nand U1369 (N_1369,N_617,N_1054);
nand U1370 (N_1370,N_500,N_1125);
nor U1371 (N_1371,N_445,In_1436);
xnor U1372 (N_1372,In_1918,In_1683);
and U1373 (N_1373,N_607,N_435);
and U1374 (N_1374,In_328,In_1858);
xnor U1375 (N_1375,N_979,N_798);
or U1376 (N_1376,N_1122,In_587);
nand U1377 (N_1377,N_943,N_384);
and U1378 (N_1378,N_742,N_408);
nand U1379 (N_1379,In_462,N_750);
and U1380 (N_1380,N_1094,N_902);
xor U1381 (N_1381,N_1007,In_1686);
and U1382 (N_1382,N_1093,N_809);
or U1383 (N_1383,N_20,N_508);
nor U1384 (N_1384,In_1574,N_428);
or U1385 (N_1385,N_1192,In_100);
xor U1386 (N_1386,In_202,N_855);
or U1387 (N_1387,In_1957,In_1174);
and U1388 (N_1388,N_1116,N_1070);
or U1389 (N_1389,In_1015,N_1144);
nand U1390 (N_1390,N_529,N_1159);
nor U1391 (N_1391,N_406,N_725);
nand U1392 (N_1392,In_1153,In_1247);
nor U1393 (N_1393,N_951,N_277);
or U1394 (N_1394,In_968,N_936);
nor U1395 (N_1395,N_795,N_1047);
nor U1396 (N_1396,N_502,N_86);
xnor U1397 (N_1397,N_616,N_976);
nor U1398 (N_1398,In_1887,In_1697);
xor U1399 (N_1399,N_341,In_1830);
xnor U1400 (N_1400,N_1255,N_1115);
and U1401 (N_1401,In_774,In_1185);
xnor U1402 (N_1402,N_383,N_977);
nor U1403 (N_1403,N_1227,N_1076);
or U1404 (N_1404,In_525,N_1349);
or U1405 (N_1405,N_1338,In_671);
or U1406 (N_1406,In_1108,N_1283);
or U1407 (N_1407,N_1385,N_927);
xnor U1408 (N_1408,N_1314,N_1013);
nand U1409 (N_1409,N_1098,N_1304);
xnor U1410 (N_1410,N_1345,N_1164);
nor U1411 (N_1411,N_1189,N_1388);
nor U1412 (N_1412,N_1073,N_688);
or U1413 (N_1413,In_1954,N_1375);
nand U1414 (N_1414,N_1010,N_738);
nor U1415 (N_1415,N_1356,In_1671);
nor U1416 (N_1416,N_1274,N_45);
nor U1417 (N_1417,N_968,N_1151);
nor U1418 (N_1418,N_954,N_1393);
xnor U1419 (N_1419,N_1233,N_810);
nor U1420 (N_1420,In_654,N_998);
and U1421 (N_1421,N_1280,N_1390);
or U1422 (N_1422,N_387,N_1307);
or U1423 (N_1423,N_1135,N_910);
nor U1424 (N_1424,In_1948,N_355);
and U1425 (N_1425,N_1365,N_1259);
and U1426 (N_1426,N_1099,N_603);
or U1427 (N_1427,N_1155,N_653);
or U1428 (N_1428,N_1339,N_794);
nand U1429 (N_1429,N_865,N_1235);
xnor U1430 (N_1430,N_1347,N_1374);
or U1431 (N_1431,N_626,In_763);
or U1432 (N_1432,N_1241,N_1041);
nand U1433 (N_1433,N_1277,N_1380);
xnor U1434 (N_1434,N_1362,In_400);
nand U1435 (N_1435,N_1147,In_1744);
nor U1436 (N_1436,N_712,In_61);
nor U1437 (N_1437,N_13,N_116);
nor U1438 (N_1438,N_1206,N_963);
nor U1439 (N_1439,N_287,N_1353);
nand U1440 (N_1440,N_646,N_944);
or U1441 (N_1441,N_1389,N_1371);
and U1442 (N_1442,N_1224,N_1243);
nor U1443 (N_1443,N_1112,N_1381);
or U1444 (N_1444,N_1294,In_1194);
or U1445 (N_1445,N_1285,N_989);
and U1446 (N_1446,N_569,N_1090);
xor U1447 (N_1447,N_921,N_1337);
nand U1448 (N_1448,In_1944,N_1160);
nor U1449 (N_1449,N_1254,N_791);
or U1450 (N_1450,N_1051,N_1370);
xnor U1451 (N_1451,N_1032,N_1273);
xnor U1452 (N_1452,N_663,N_1306);
and U1453 (N_1453,N_1290,In_1872);
nand U1454 (N_1454,N_1208,In_1923);
or U1455 (N_1455,N_830,N_1324);
nor U1456 (N_1456,N_1313,In_832);
nor U1457 (N_1457,N_656,In_1648);
and U1458 (N_1458,N_1373,N_1137);
xor U1459 (N_1459,In_192,N_1301);
nor U1460 (N_1460,In_705,N_1272);
nand U1461 (N_1461,N_1221,N_1298);
and U1462 (N_1462,N_259,N_219);
nor U1463 (N_1463,N_1226,N_1193);
or U1464 (N_1464,In_1992,N_800);
nor U1465 (N_1465,N_1296,N_1281);
nor U1466 (N_1466,N_21,N_1269);
and U1467 (N_1467,N_1143,In_430);
nor U1468 (N_1468,N_763,N_1002);
and U1469 (N_1469,In_71,N_1211);
and U1470 (N_1470,In_951,N_1246);
nor U1471 (N_1471,N_1326,In_174);
nor U1472 (N_1472,N_1234,N_294);
or U1473 (N_1473,In_1483,N_1240);
or U1474 (N_1474,N_1068,In_27);
nand U1475 (N_1475,In_1339,N_1348);
nor U1476 (N_1476,N_1188,N_1384);
or U1477 (N_1477,In_1545,In_1006);
or U1478 (N_1478,N_270,N_611);
nand U1479 (N_1479,In_1727,N_1217);
and U1480 (N_1480,N_79,N_1209);
nor U1481 (N_1481,N_624,In_822);
or U1482 (N_1482,N_1202,N_1248);
nor U1483 (N_1483,N_1312,In_1934);
or U1484 (N_1484,N_1053,N_1256);
xor U1485 (N_1485,N_1062,N_242);
nor U1486 (N_1486,N_1263,N_861);
nor U1487 (N_1487,N_465,N_559);
nor U1488 (N_1488,N_1333,N_1026);
and U1489 (N_1489,In_736,N_821);
nand U1490 (N_1490,N_1074,In_404);
nand U1491 (N_1491,N_1119,N_999);
nand U1492 (N_1492,N_935,N_1250);
nand U1493 (N_1493,N_1391,In_1732);
and U1494 (N_1494,N_1223,In_1367);
nand U1495 (N_1495,In_232,N_1278);
nand U1496 (N_1496,In_647,N_178);
and U1497 (N_1497,N_1377,N_1214);
or U1498 (N_1498,N_776,N_216);
and U1499 (N_1499,In_249,N_1382);
and U1500 (N_1500,N_1244,N_1030);
xnor U1501 (N_1501,N_1340,In_941);
xnor U1502 (N_1502,In_133,N_894);
or U1503 (N_1503,N_787,N_1264);
and U1504 (N_1504,N_1351,N_361);
nor U1505 (N_1505,N_1123,N_1327);
or U1506 (N_1506,N_1336,N_1060);
and U1507 (N_1507,In_304,N_1343);
xnor U1508 (N_1508,N_1201,N_1105);
or U1509 (N_1509,N_1268,In_1316);
and U1510 (N_1510,N_973,In_1124);
and U1511 (N_1511,In_1202,N_1369);
and U1512 (N_1512,In_1523,N_1237);
and U1513 (N_1513,In_1799,N_1316);
or U1514 (N_1514,N_1203,N_1009);
nand U1515 (N_1515,In_1541,N_1242);
and U1516 (N_1516,N_1078,N_1247);
and U1517 (N_1517,N_414,N_1177);
xnor U1518 (N_1518,N_292,In_1126);
nor U1519 (N_1519,N_1300,N_630);
xnor U1520 (N_1520,N_1216,In_1773);
xor U1521 (N_1521,N_1004,N_1245);
nor U1522 (N_1522,N_1109,N_1395);
or U1523 (N_1523,N_827,In_1021);
xor U1524 (N_1524,N_1219,In_445);
nand U1525 (N_1525,N_1232,N_516);
and U1526 (N_1526,N_1261,In_1083);
or U1527 (N_1527,In_1539,In_63);
and U1528 (N_1528,In_1494,N_767);
nor U1529 (N_1529,N_507,N_1266);
nand U1530 (N_1530,N_326,N_1174);
nand U1531 (N_1531,N_1321,N_1210);
and U1532 (N_1532,N_1039,N_1178);
nand U1533 (N_1533,N_772,N_523);
nand U1534 (N_1534,In_204,N_1108);
xnor U1535 (N_1535,N_1359,In_1313);
nor U1536 (N_1536,In_810,In_1321);
nand U1537 (N_1537,N_1138,N_1236);
xnor U1538 (N_1538,N_1012,N_1069);
nand U1539 (N_1539,N_522,N_1392);
nand U1540 (N_1540,In_1140,N_1265);
xnor U1541 (N_1541,N_1134,N_1372);
xor U1542 (N_1542,N_1368,N_854);
or U1543 (N_1543,N_1229,N_1270);
nor U1544 (N_1544,In_1257,N_1334);
xnor U1545 (N_1545,In_1253,N_1376);
xnor U1546 (N_1546,N_997,N_642);
nor U1547 (N_1547,N_1050,N_330);
or U1548 (N_1548,N_987,In_109);
or U1549 (N_1549,In_1245,In_270);
xor U1550 (N_1550,N_717,N_1342);
nand U1551 (N_1551,N_814,N_1126);
nor U1552 (N_1552,N_1249,N_371);
xnor U1553 (N_1553,N_1038,N_1031);
or U1554 (N_1554,N_1315,N_554);
or U1555 (N_1555,N_1022,N_1332);
nand U1556 (N_1556,N_80,N_1360);
xor U1557 (N_1557,N_1084,N_1215);
xor U1558 (N_1558,In_1118,N_1251);
and U1559 (N_1559,N_850,In_1601);
nand U1560 (N_1560,In_1803,N_1081);
xor U1561 (N_1561,In_1334,In_1680);
nor U1562 (N_1562,N_1225,N_658);
xnor U1563 (N_1563,N_308,N_1016);
nor U1564 (N_1564,N_1146,N_758);
xor U1565 (N_1565,N_966,N_1191);
or U1566 (N_1566,N_1386,In_399);
and U1567 (N_1567,In_541,N_1132);
xnor U1568 (N_1568,In_1358,N_1154);
or U1569 (N_1569,N_1291,N_1218);
or U1570 (N_1570,N_1220,N_1230);
xor U1571 (N_1571,N_490,N_705);
or U1572 (N_1572,N_1346,N_665);
nand U1573 (N_1573,In_1333,N_1195);
or U1574 (N_1574,N_1181,N_1036);
xor U1575 (N_1575,N_541,In_698);
and U1576 (N_1576,N_1019,N_1158);
xor U1577 (N_1577,N_1267,N_1088);
and U1578 (N_1578,In_1925,N_1335);
and U1579 (N_1579,N_1363,N_1253);
nor U1580 (N_1580,N_1354,N_41);
nor U1581 (N_1581,In_269,N_1072);
nand U1582 (N_1582,In_288,N_1258);
or U1583 (N_1583,In_1435,N_1087);
nor U1584 (N_1584,N_12,N_370);
nand U1585 (N_1585,N_1040,N_509);
and U1586 (N_1586,N_869,N_1003);
or U1587 (N_1587,N_1059,N_874);
and U1588 (N_1588,In_1020,In_1312);
xnor U1589 (N_1589,N_1322,N_1200);
and U1590 (N_1590,In_1121,In_322);
nor U1591 (N_1591,N_1399,N_582);
nand U1592 (N_1592,N_440,N_884);
nor U1593 (N_1593,N_1124,N_1325);
xnor U1594 (N_1594,N_1023,N_1101);
and U1595 (N_1595,N_1303,N_579);
xnor U1596 (N_1596,In_976,N_1100);
nor U1597 (N_1597,N_1364,N_967);
or U1598 (N_1598,N_1029,N_858);
nand U1599 (N_1599,N_1320,N_1252);
xnor U1600 (N_1600,N_1456,N_1057);
xor U1601 (N_1601,N_1577,N_1133);
xor U1602 (N_1602,In_184,N_1599);
nand U1603 (N_1603,N_1411,N_1429);
xor U1604 (N_1604,N_1199,N_1582);
nand U1605 (N_1605,N_919,In_169);
or U1606 (N_1606,N_1308,N_1495);
and U1607 (N_1607,N_1425,N_1434);
or U1608 (N_1608,N_1572,N_1554);
nor U1609 (N_1609,N_1006,N_33);
nand U1610 (N_1610,N_1297,In_986);
nand U1611 (N_1611,N_1430,In_1868);
or U1612 (N_1612,N_1379,N_1594);
or U1613 (N_1613,In_43,N_1590);
nand U1614 (N_1614,N_1474,N_1366);
xnor U1615 (N_1615,N_1418,N_1561);
nor U1616 (N_1616,N_1485,N_609);
xnor U1617 (N_1617,N_1541,N_448);
nor U1618 (N_1618,N_1525,N_1568);
xor U1619 (N_1619,N_872,N_990);
nor U1620 (N_1620,N_548,N_608);
nor U1621 (N_1621,N_1504,N_1257);
or U1622 (N_1622,N_1443,In_995);
nand U1623 (N_1623,N_1579,N_1396);
and U1624 (N_1624,N_1421,N_1417);
xor U1625 (N_1625,N_1439,N_1516);
or U1626 (N_1626,N_1444,N_1427);
xor U1627 (N_1627,N_1449,N_1473);
nand U1628 (N_1628,N_1424,N_909);
or U1629 (N_1629,N_804,N_335);
or U1630 (N_1630,N_1262,N_443);
nand U1631 (N_1631,In_1490,N_1287);
and U1632 (N_1632,N_1446,N_410);
nor U1633 (N_1633,N_1292,N_1302);
nor U1634 (N_1634,N_1546,N_1387);
and U1635 (N_1635,N_1534,N_1065);
xor U1636 (N_1636,N_1596,N_1463);
nor U1637 (N_1637,N_1578,In_167);
and U1638 (N_1638,N_1328,N_1518);
or U1639 (N_1639,N_1358,N_1213);
xnor U1640 (N_1640,N_1136,N_1482);
and U1641 (N_1641,N_1148,N_1588);
xnor U1642 (N_1642,N_1498,N_1271);
and U1643 (N_1643,N_1408,N_876);
nand U1644 (N_1644,N_983,N_1079);
or U1645 (N_1645,In_695,N_1423);
and U1646 (N_1646,N_1575,In_1711);
and U1647 (N_1647,N_1414,N_1350);
nor U1648 (N_1648,N_1432,N_1415);
nor U1649 (N_1649,In_1356,N_1573);
xnor U1650 (N_1650,N_1082,N_1515);
nand U1651 (N_1651,N_1555,N_1305);
nor U1652 (N_1652,N_728,In_1651);
nand U1653 (N_1653,N_1467,N_1407);
and U1654 (N_1654,N_1282,N_1576);
or U1655 (N_1655,N_1536,N_1319);
or U1656 (N_1656,N_1491,N_660);
xnor U1657 (N_1657,N_1450,In_1089);
nor U1658 (N_1658,N_1121,N_1526);
and U1659 (N_1659,N_1490,N_1586);
nor U1660 (N_1660,N_1445,N_1564);
or U1661 (N_1661,N_1212,N_1309);
xnor U1662 (N_1662,N_1496,N_1157);
xnor U1663 (N_1663,N_1484,N_1488);
nand U1664 (N_1664,N_107,N_1204);
nand U1665 (N_1665,N_1595,N_1293);
nand U1666 (N_1666,N_567,N_547);
nand U1667 (N_1667,N_1585,N_1317);
and U1668 (N_1668,In_532,N_1583);
and U1669 (N_1669,N_1549,N_1344);
or U1670 (N_1670,N_545,N_434);
nor U1671 (N_1671,N_1487,N_1462);
or U1672 (N_1672,N_1533,N_1436);
xor U1673 (N_1673,N_1501,N_1481);
nand U1674 (N_1674,N_1565,N_1404);
and U1675 (N_1675,N_1514,N_1508);
or U1676 (N_1676,N_1475,N_1402);
and U1677 (N_1677,N_1355,N_1567);
and U1678 (N_1678,N_1571,N_1551);
nor U1679 (N_1679,N_940,N_1431);
and U1680 (N_1680,N_429,N_1091);
nand U1681 (N_1681,In_374,In_811);
nor U1682 (N_1682,N_1548,N_1483);
nand U1683 (N_1683,N_1289,N_1507);
and U1684 (N_1684,N_729,N_1540);
and U1685 (N_1685,N_1420,N_1288);
nor U1686 (N_1686,N_1357,N_685);
or U1687 (N_1687,N_744,N_1410);
xnor U1688 (N_1688,N_1486,N_1400);
or U1689 (N_1689,N_895,N_1447);
and U1690 (N_1690,N_1512,N_1067);
or U1691 (N_1691,N_1464,N_1409);
or U1692 (N_1692,In_1758,N_1465);
nand U1693 (N_1693,N_1497,In_567);
xor U1694 (N_1694,N_929,N_1064);
and U1695 (N_1695,N_1466,N_1383);
xor U1696 (N_1696,N_1560,N_1150);
or U1697 (N_1697,N_1037,N_1428);
nand U1698 (N_1698,N_1557,N_1352);
nand U1699 (N_1699,N_834,N_1520);
or U1700 (N_1700,N_1457,N_1517);
and U1701 (N_1701,N_1598,N_149);
nand U1702 (N_1702,N_1419,In_134);
nand U1703 (N_1703,N_1207,N_1231);
nor U1704 (N_1704,N_1511,N_1239);
nor U1705 (N_1705,N_831,N_1530);
nand U1706 (N_1706,N_1001,N_1422);
xnor U1707 (N_1707,N_1179,N_543);
xnor U1708 (N_1708,N_1503,N_1397);
xnor U1709 (N_1709,N_1597,N_1522);
nor U1710 (N_1710,N_1470,In_638);
nand U1711 (N_1711,N_1506,N_697);
and U1712 (N_1712,N_1437,N_1412);
xor U1713 (N_1713,N_1528,N_1341);
or U1714 (N_1714,N_1532,N_230);
nor U1715 (N_1715,N_1545,N_1562);
nor U1716 (N_1716,N_1558,N_1531);
xnor U1717 (N_1717,In_787,N_1587);
nand U1718 (N_1718,N_1401,N_1279);
or U1719 (N_1719,N_1228,N_1329);
or U1720 (N_1720,In_1444,N_1476);
or U1721 (N_1721,N_1190,N_1547);
and U1722 (N_1722,N_1455,N_1238);
nand U1723 (N_1723,N_1014,N_1406);
nor U1724 (N_1724,N_1524,N_801);
xor U1725 (N_1725,N_1260,In_1087);
or U1726 (N_1726,N_1538,N_84);
xor U1727 (N_1727,N_1435,N_949);
and U1728 (N_1728,N_1071,N_1453);
and U1729 (N_1729,N_1172,N_542);
nor U1730 (N_1730,N_1378,N_1458);
nor U1731 (N_1731,N_1566,N_1323);
xor U1732 (N_1732,In_684,N_1367);
xor U1733 (N_1733,In_1009,N_1550);
xor U1734 (N_1734,N_1438,N_1284);
nand U1735 (N_1735,N_1106,N_1472);
nand U1736 (N_1736,N_1299,N_1563);
or U1737 (N_1737,N_1095,N_1128);
and U1738 (N_1738,N_1153,N_1500);
or U1739 (N_1739,N_1045,N_1361);
nand U1740 (N_1740,N_1295,N_823);
nand U1741 (N_1741,In_1865,In_1143);
xnor U1742 (N_1742,N_1441,In_1326);
xnor U1743 (N_1743,N_1535,N_1176);
nor U1744 (N_1744,In_323,N_1591);
xor U1745 (N_1745,N_240,N_1107);
or U1746 (N_1746,N_1509,N_1584);
and U1747 (N_1747,N_699,N_1480);
xor U1748 (N_1748,N_1460,N_1398);
xnor U1749 (N_1749,N_1494,N_1519);
nand U1750 (N_1750,N_1477,N_870);
nand U1751 (N_1751,N_1033,In_121);
nor U1752 (N_1752,N_1426,N_1433);
and U1753 (N_1753,In_715,N_1454);
nor U1754 (N_1754,N_1394,N_1542);
xnor U1755 (N_1755,N_1403,N_1513);
or U1756 (N_1756,N_1286,N_1440);
nor U1757 (N_1757,N_396,N_1493);
nor U1758 (N_1758,N_1527,N_698);
xnor U1759 (N_1759,N_879,N_1468);
and U1760 (N_1760,N_871,N_1205);
nand U1761 (N_1761,N_1451,N_1537);
xor U1762 (N_1762,N_1521,In_888);
or U1763 (N_1763,N_1120,N_1478);
xnor U1764 (N_1764,N_1276,N_1173);
or U1765 (N_1765,N_1413,N_957);
and U1766 (N_1766,N_1184,N_1552);
nand U1767 (N_1767,In_990,N_1459);
nand U1768 (N_1768,N_1448,N_1553);
or U1769 (N_1769,N_664,In_1931);
nand U1770 (N_1770,N_619,N_1471);
xor U1771 (N_1771,In_236,N_1556);
xor U1772 (N_1772,N_1592,N_1502);
xor U1773 (N_1773,N_1589,N_1008);
xnor U1774 (N_1774,N_1580,N_1405);
nor U1775 (N_1775,N_721,N_1479);
or U1776 (N_1776,N_1318,In_545);
or U1777 (N_1777,N_1544,In_928);
and U1778 (N_1778,In_683,N_1574);
xor U1779 (N_1779,N_1559,N_845);
nand U1780 (N_1780,N_1492,N_1569);
and U1781 (N_1781,N_1593,N_1489);
xor U1782 (N_1782,N_1499,N_1331);
nor U1783 (N_1783,N_1197,N_1581);
and U1784 (N_1784,In_1884,N_177);
and U1785 (N_1785,N_1310,N_1543);
nand U1786 (N_1786,In_904,N_1529);
or U1787 (N_1787,In_1843,N_1222);
and U1788 (N_1788,N_1275,N_739);
nand U1789 (N_1789,N_613,N_1469);
xnor U1790 (N_1790,In_140,In_560);
nor U1791 (N_1791,N_1461,N_1416);
xnor U1792 (N_1792,N_1570,N_453);
nor U1793 (N_1793,N_1442,In_711);
and U1794 (N_1794,In_261,N_1452);
nand U1795 (N_1795,N_1523,N_1510);
nand U1796 (N_1796,N_1539,N_1311);
nand U1797 (N_1797,N_852,N_566);
xnor U1798 (N_1798,N_900,N_1330);
and U1799 (N_1799,N_1505,N_419);
or U1800 (N_1800,N_1732,N_1693);
and U1801 (N_1801,N_1749,N_1615);
and U1802 (N_1802,N_1625,N_1631);
or U1803 (N_1803,N_1629,N_1704);
or U1804 (N_1804,N_1636,N_1602);
xor U1805 (N_1805,N_1705,N_1607);
xor U1806 (N_1806,N_1726,N_1670);
nor U1807 (N_1807,N_1683,N_1765);
nand U1808 (N_1808,N_1622,N_1745);
nand U1809 (N_1809,N_1772,N_1784);
and U1810 (N_1810,N_1734,N_1685);
and U1811 (N_1811,N_1656,N_1603);
nand U1812 (N_1812,N_1623,N_1643);
nor U1813 (N_1813,N_1746,N_1662);
nor U1814 (N_1814,N_1681,N_1616);
xor U1815 (N_1815,N_1678,N_1755);
and U1816 (N_1816,N_1740,N_1692);
nand U1817 (N_1817,N_1761,N_1609);
or U1818 (N_1818,N_1758,N_1727);
nor U1819 (N_1819,N_1613,N_1730);
and U1820 (N_1820,N_1661,N_1788);
nor U1821 (N_1821,N_1669,N_1645);
nand U1822 (N_1822,N_1647,N_1779);
nor U1823 (N_1823,N_1640,N_1757);
or U1824 (N_1824,N_1688,N_1795);
or U1825 (N_1825,N_1697,N_1708);
or U1826 (N_1826,N_1781,N_1687);
xor U1827 (N_1827,N_1780,N_1621);
nor U1828 (N_1828,N_1775,N_1718);
xnor U1829 (N_1829,N_1604,N_1675);
nand U1830 (N_1830,N_1703,N_1762);
xnor U1831 (N_1831,N_1763,N_1699);
or U1832 (N_1832,N_1676,N_1690);
nand U1833 (N_1833,N_1711,N_1619);
or U1834 (N_1834,N_1796,N_1766);
nand U1835 (N_1835,N_1793,N_1709);
xnor U1836 (N_1836,N_1701,N_1728);
nand U1837 (N_1837,N_1677,N_1725);
nand U1838 (N_1838,N_1630,N_1782);
xnor U1839 (N_1839,N_1628,N_1614);
or U1840 (N_1840,N_1664,N_1665);
xnor U1841 (N_1841,N_1611,N_1794);
or U1842 (N_1842,N_1691,N_1663);
nand U1843 (N_1843,N_1741,N_1733);
nor U1844 (N_1844,N_1715,N_1717);
nor U1845 (N_1845,N_1600,N_1658);
nor U1846 (N_1846,N_1632,N_1624);
and U1847 (N_1847,N_1649,N_1798);
nand U1848 (N_1848,N_1689,N_1713);
nor U1849 (N_1849,N_1768,N_1744);
xor U1850 (N_1850,N_1682,N_1627);
or U1851 (N_1851,N_1698,N_1684);
nor U1852 (N_1852,N_1694,N_1799);
nand U1853 (N_1853,N_1738,N_1736);
nand U1854 (N_1854,N_1606,N_1756);
nor U1855 (N_1855,N_1770,N_1743);
xnor U1856 (N_1856,N_1724,N_1617);
or U1857 (N_1857,N_1605,N_1791);
or U1858 (N_1858,N_1633,N_1774);
and U1859 (N_1859,N_1783,N_1680);
xor U1860 (N_1860,N_1773,N_1706);
and U1861 (N_1861,N_1722,N_1660);
and U1862 (N_1862,N_1721,N_1648);
nor U1863 (N_1863,N_1750,N_1635);
nor U1864 (N_1864,N_1618,N_1747);
and U1865 (N_1865,N_1639,N_1612);
nand U1866 (N_1866,N_1769,N_1771);
or U1867 (N_1867,N_1729,N_1737);
nor U1868 (N_1868,N_1641,N_1797);
or U1869 (N_1869,N_1601,N_1686);
nor U1870 (N_1870,N_1716,N_1702);
xor U1871 (N_1871,N_1719,N_1651);
or U1872 (N_1872,N_1785,N_1787);
xnor U1873 (N_1873,N_1735,N_1638);
or U1874 (N_1874,N_1634,N_1748);
nor U1875 (N_1875,N_1778,N_1714);
nor U1876 (N_1876,N_1650,N_1789);
nand U1877 (N_1877,N_1786,N_1751);
or U1878 (N_1878,N_1626,N_1655);
xnor U1879 (N_1879,N_1672,N_1760);
and U1880 (N_1880,N_1654,N_1642);
or U1881 (N_1881,N_1752,N_1608);
and U1882 (N_1882,N_1700,N_1667);
xor U1883 (N_1883,N_1777,N_1671);
nand U1884 (N_1884,N_1790,N_1696);
xor U1885 (N_1885,N_1679,N_1720);
or U1886 (N_1886,N_1739,N_1668);
xnor U1887 (N_1887,N_1742,N_1759);
or U1888 (N_1888,N_1707,N_1754);
or U1889 (N_1889,N_1644,N_1767);
xor U1890 (N_1890,N_1646,N_1712);
nand U1891 (N_1891,N_1695,N_1776);
nand U1892 (N_1892,N_1657,N_1792);
nor U1893 (N_1893,N_1659,N_1710);
or U1894 (N_1894,N_1620,N_1731);
nand U1895 (N_1895,N_1652,N_1753);
and U1896 (N_1896,N_1723,N_1764);
xnor U1897 (N_1897,N_1653,N_1666);
and U1898 (N_1898,N_1610,N_1637);
nand U1899 (N_1899,N_1674,N_1673);
nand U1900 (N_1900,N_1714,N_1635);
and U1901 (N_1901,N_1723,N_1789);
xnor U1902 (N_1902,N_1603,N_1769);
and U1903 (N_1903,N_1600,N_1790);
or U1904 (N_1904,N_1774,N_1634);
nand U1905 (N_1905,N_1655,N_1616);
nor U1906 (N_1906,N_1776,N_1746);
nand U1907 (N_1907,N_1727,N_1712);
or U1908 (N_1908,N_1685,N_1628);
nor U1909 (N_1909,N_1789,N_1677);
or U1910 (N_1910,N_1717,N_1728);
xor U1911 (N_1911,N_1688,N_1651);
and U1912 (N_1912,N_1747,N_1716);
xnor U1913 (N_1913,N_1781,N_1778);
and U1914 (N_1914,N_1731,N_1625);
xor U1915 (N_1915,N_1792,N_1664);
nor U1916 (N_1916,N_1739,N_1630);
nand U1917 (N_1917,N_1696,N_1736);
xor U1918 (N_1918,N_1713,N_1669);
xnor U1919 (N_1919,N_1735,N_1760);
and U1920 (N_1920,N_1723,N_1660);
nand U1921 (N_1921,N_1728,N_1630);
xor U1922 (N_1922,N_1661,N_1748);
xor U1923 (N_1923,N_1789,N_1782);
nor U1924 (N_1924,N_1642,N_1778);
xnor U1925 (N_1925,N_1657,N_1786);
nand U1926 (N_1926,N_1797,N_1691);
and U1927 (N_1927,N_1667,N_1689);
nor U1928 (N_1928,N_1678,N_1668);
xnor U1929 (N_1929,N_1778,N_1770);
nand U1930 (N_1930,N_1760,N_1787);
xor U1931 (N_1931,N_1734,N_1709);
or U1932 (N_1932,N_1761,N_1793);
nor U1933 (N_1933,N_1637,N_1729);
or U1934 (N_1934,N_1617,N_1685);
nor U1935 (N_1935,N_1764,N_1647);
or U1936 (N_1936,N_1685,N_1706);
xnor U1937 (N_1937,N_1745,N_1690);
nor U1938 (N_1938,N_1671,N_1612);
nor U1939 (N_1939,N_1649,N_1665);
nor U1940 (N_1940,N_1701,N_1707);
or U1941 (N_1941,N_1695,N_1747);
and U1942 (N_1942,N_1603,N_1755);
nor U1943 (N_1943,N_1600,N_1617);
nor U1944 (N_1944,N_1622,N_1635);
and U1945 (N_1945,N_1645,N_1757);
nor U1946 (N_1946,N_1701,N_1662);
nand U1947 (N_1947,N_1680,N_1600);
and U1948 (N_1948,N_1665,N_1768);
xor U1949 (N_1949,N_1664,N_1607);
xor U1950 (N_1950,N_1743,N_1740);
nor U1951 (N_1951,N_1711,N_1620);
nand U1952 (N_1952,N_1725,N_1744);
or U1953 (N_1953,N_1660,N_1789);
nor U1954 (N_1954,N_1749,N_1693);
nand U1955 (N_1955,N_1699,N_1611);
xnor U1956 (N_1956,N_1634,N_1741);
or U1957 (N_1957,N_1733,N_1619);
nor U1958 (N_1958,N_1770,N_1751);
and U1959 (N_1959,N_1735,N_1721);
or U1960 (N_1960,N_1711,N_1780);
nand U1961 (N_1961,N_1779,N_1674);
and U1962 (N_1962,N_1734,N_1720);
or U1963 (N_1963,N_1769,N_1748);
or U1964 (N_1964,N_1602,N_1762);
nand U1965 (N_1965,N_1696,N_1602);
nand U1966 (N_1966,N_1628,N_1774);
or U1967 (N_1967,N_1635,N_1727);
or U1968 (N_1968,N_1705,N_1613);
and U1969 (N_1969,N_1613,N_1761);
nand U1970 (N_1970,N_1730,N_1760);
and U1971 (N_1971,N_1722,N_1718);
nand U1972 (N_1972,N_1699,N_1716);
or U1973 (N_1973,N_1732,N_1751);
xor U1974 (N_1974,N_1669,N_1690);
and U1975 (N_1975,N_1742,N_1667);
or U1976 (N_1976,N_1746,N_1735);
nor U1977 (N_1977,N_1718,N_1651);
nor U1978 (N_1978,N_1700,N_1638);
or U1979 (N_1979,N_1654,N_1733);
xnor U1980 (N_1980,N_1717,N_1703);
or U1981 (N_1981,N_1718,N_1734);
or U1982 (N_1982,N_1743,N_1622);
nor U1983 (N_1983,N_1660,N_1609);
xor U1984 (N_1984,N_1767,N_1663);
xnor U1985 (N_1985,N_1750,N_1703);
and U1986 (N_1986,N_1740,N_1684);
or U1987 (N_1987,N_1667,N_1614);
or U1988 (N_1988,N_1755,N_1677);
xor U1989 (N_1989,N_1635,N_1610);
xnor U1990 (N_1990,N_1721,N_1797);
nand U1991 (N_1991,N_1650,N_1658);
xnor U1992 (N_1992,N_1742,N_1710);
xnor U1993 (N_1993,N_1680,N_1656);
or U1994 (N_1994,N_1678,N_1769);
xnor U1995 (N_1995,N_1735,N_1645);
xnor U1996 (N_1996,N_1684,N_1716);
and U1997 (N_1997,N_1739,N_1719);
or U1998 (N_1998,N_1719,N_1671);
xnor U1999 (N_1999,N_1799,N_1792);
xnor U2000 (N_2000,N_1807,N_1881);
nand U2001 (N_2001,N_1983,N_1865);
nor U2002 (N_2002,N_1984,N_1966);
and U2003 (N_2003,N_1872,N_1967);
nor U2004 (N_2004,N_1802,N_1895);
nand U2005 (N_2005,N_1852,N_1862);
nand U2006 (N_2006,N_1943,N_1860);
or U2007 (N_2007,N_1866,N_1937);
nand U2008 (N_2008,N_1936,N_1871);
nor U2009 (N_2009,N_1816,N_1949);
nor U2010 (N_2010,N_1810,N_1854);
xor U2011 (N_2011,N_1896,N_1837);
and U2012 (N_2012,N_1999,N_1976);
nand U2013 (N_2013,N_1844,N_1954);
or U2014 (N_2014,N_1805,N_1817);
and U2015 (N_2015,N_1975,N_1992);
nor U2016 (N_2016,N_1877,N_1888);
and U2017 (N_2017,N_1884,N_1990);
or U2018 (N_2018,N_1820,N_1917);
nand U2019 (N_2019,N_1841,N_1955);
nand U2020 (N_2020,N_1907,N_1809);
nor U2021 (N_2021,N_1869,N_1856);
nand U2022 (N_2022,N_1938,N_1926);
and U2023 (N_2023,N_1977,N_1800);
nor U2024 (N_2024,N_1879,N_1850);
xnor U2025 (N_2025,N_1801,N_1929);
or U2026 (N_2026,N_1913,N_1858);
nor U2027 (N_2027,N_1830,N_1857);
nor U2028 (N_2028,N_1952,N_1935);
xnor U2029 (N_2029,N_1883,N_1867);
nand U2030 (N_2030,N_1873,N_1847);
or U2031 (N_2031,N_1964,N_1996);
nor U2032 (N_2032,N_1875,N_1973);
and U2033 (N_2033,N_1957,N_1928);
nand U2034 (N_2034,N_1988,N_1861);
and U2035 (N_2035,N_1812,N_1918);
xnor U2036 (N_2036,N_1925,N_1835);
or U2037 (N_2037,N_1824,N_1922);
or U2038 (N_2038,N_1985,N_1946);
and U2039 (N_2039,N_1815,N_1961);
or U2040 (N_2040,N_1934,N_1828);
or U2041 (N_2041,N_1890,N_1940);
and U2042 (N_2042,N_1924,N_1995);
nor U2043 (N_2043,N_1930,N_1953);
or U2044 (N_2044,N_1887,N_1829);
nand U2045 (N_2045,N_1838,N_1894);
xor U2046 (N_2046,N_1920,N_1959);
nand U2047 (N_2047,N_1901,N_1944);
xor U2048 (N_2048,N_1904,N_1902);
xor U2049 (N_2049,N_1915,N_1911);
or U2050 (N_2050,N_1803,N_1851);
xor U2051 (N_2051,N_1832,N_1994);
and U2052 (N_2052,N_1876,N_1848);
or U2053 (N_2053,N_1965,N_1956);
nand U2054 (N_2054,N_1827,N_1912);
nor U2055 (N_2055,N_1974,N_1905);
or U2056 (N_2056,N_1921,N_1989);
nor U2057 (N_2057,N_1980,N_1981);
or U2058 (N_2058,N_1997,N_1914);
xnor U2059 (N_2059,N_1826,N_1840);
nand U2060 (N_2060,N_1839,N_1855);
xnor U2061 (N_2061,N_1945,N_1806);
nand U2062 (N_2062,N_1972,N_1853);
or U2063 (N_2063,N_1836,N_1931);
nor U2064 (N_2064,N_1886,N_1843);
xor U2065 (N_2065,N_1960,N_1874);
or U2066 (N_2066,N_1932,N_1822);
nor U2067 (N_2067,N_1948,N_1814);
nand U2068 (N_2068,N_1909,N_1906);
nor U2069 (N_2069,N_1951,N_1947);
xor U2070 (N_2070,N_1979,N_1882);
xnor U2071 (N_2071,N_1991,N_1823);
nand U2072 (N_2072,N_1833,N_1868);
or U2073 (N_2073,N_1933,N_1923);
or U2074 (N_2074,N_1939,N_1880);
nand U2075 (N_2075,N_1885,N_1897);
and U2076 (N_2076,N_1987,N_1962);
nor U2077 (N_2077,N_1900,N_1971);
or U2078 (N_2078,N_1834,N_1893);
and U2079 (N_2079,N_1831,N_1819);
and U2080 (N_2080,N_1908,N_1916);
and U2081 (N_2081,N_1864,N_1993);
nor U2082 (N_2082,N_1808,N_1870);
nor U2083 (N_2083,N_1863,N_1950);
nand U2084 (N_2084,N_1898,N_1813);
and U2085 (N_2085,N_1804,N_1889);
and U2086 (N_2086,N_1878,N_1919);
or U2087 (N_2087,N_1891,N_1982);
or U2088 (N_2088,N_1998,N_1818);
xnor U2089 (N_2089,N_1942,N_1969);
nand U2090 (N_2090,N_1846,N_1859);
or U2091 (N_2091,N_1849,N_1978);
xor U2092 (N_2092,N_1892,N_1958);
nor U2093 (N_2093,N_1899,N_1927);
or U2094 (N_2094,N_1825,N_1968);
nand U2095 (N_2095,N_1821,N_1970);
and U2096 (N_2096,N_1811,N_1903);
or U2097 (N_2097,N_1986,N_1941);
nand U2098 (N_2098,N_1842,N_1845);
nor U2099 (N_2099,N_1910,N_1963);
or U2100 (N_2100,N_1971,N_1865);
nor U2101 (N_2101,N_1847,N_1970);
or U2102 (N_2102,N_1995,N_1845);
nor U2103 (N_2103,N_1937,N_1823);
xor U2104 (N_2104,N_1985,N_1900);
nand U2105 (N_2105,N_1898,N_1887);
or U2106 (N_2106,N_1987,N_1955);
and U2107 (N_2107,N_1830,N_1983);
nand U2108 (N_2108,N_1904,N_1978);
xnor U2109 (N_2109,N_1855,N_1935);
or U2110 (N_2110,N_1836,N_1899);
or U2111 (N_2111,N_1863,N_1960);
or U2112 (N_2112,N_1895,N_1913);
xor U2113 (N_2113,N_1883,N_1941);
nor U2114 (N_2114,N_1863,N_1883);
xor U2115 (N_2115,N_1955,N_1958);
nand U2116 (N_2116,N_1818,N_1834);
nand U2117 (N_2117,N_1834,N_1863);
or U2118 (N_2118,N_1885,N_1925);
nand U2119 (N_2119,N_1866,N_1875);
xor U2120 (N_2120,N_1842,N_1933);
xnor U2121 (N_2121,N_1868,N_1976);
nand U2122 (N_2122,N_1900,N_1980);
nand U2123 (N_2123,N_1964,N_1827);
and U2124 (N_2124,N_1857,N_1890);
xnor U2125 (N_2125,N_1904,N_1881);
nor U2126 (N_2126,N_1813,N_1851);
or U2127 (N_2127,N_1947,N_1845);
and U2128 (N_2128,N_1890,N_1804);
nor U2129 (N_2129,N_1972,N_1833);
nand U2130 (N_2130,N_1917,N_1837);
nand U2131 (N_2131,N_1948,N_1971);
nand U2132 (N_2132,N_1932,N_1865);
nand U2133 (N_2133,N_1869,N_1865);
and U2134 (N_2134,N_1854,N_1894);
xnor U2135 (N_2135,N_1905,N_1815);
nor U2136 (N_2136,N_1856,N_1876);
or U2137 (N_2137,N_1918,N_1977);
nand U2138 (N_2138,N_1921,N_1997);
and U2139 (N_2139,N_1938,N_1857);
or U2140 (N_2140,N_1868,N_1931);
xor U2141 (N_2141,N_1878,N_1977);
nand U2142 (N_2142,N_1967,N_1972);
xor U2143 (N_2143,N_1919,N_1832);
nand U2144 (N_2144,N_1894,N_1986);
and U2145 (N_2145,N_1818,N_1980);
nand U2146 (N_2146,N_1964,N_1893);
xnor U2147 (N_2147,N_1988,N_1973);
nor U2148 (N_2148,N_1956,N_1813);
nor U2149 (N_2149,N_1971,N_1856);
xnor U2150 (N_2150,N_1830,N_1829);
nor U2151 (N_2151,N_1873,N_1958);
nor U2152 (N_2152,N_1902,N_1913);
nor U2153 (N_2153,N_1988,N_1972);
and U2154 (N_2154,N_1843,N_1840);
or U2155 (N_2155,N_1844,N_1846);
and U2156 (N_2156,N_1833,N_1994);
and U2157 (N_2157,N_1848,N_1885);
xor U2158 (N_2158,N_1997,N_1852);
and U2159 (N_2159,N_1854,N_1983);
or U2160 (N_2160,N_1814,N_1847);
xnor U2161 (N_2161,N_1838,N_1877);
or U2162 (N_2162,N_1835,N_1837);
nand U2163 (N_2163,N_1868,N_1960);
or U2164 (N_2164,N_1986,N_1980);
nand U2165 (N_2165,N_1978,N_1885);
xnor U2166 (N_2166,N_1981,N_1815);
or U2167 (N_2167,N_1973,N_1960);
or U2168 (N_2168,N_1838,N_1826);
xor U2169 (N_2169,N_1835,N_1918);
and U2170 (N_2170,N_1928,N_1848);
xor U2171 (N_2171,N_1985,N_1960);
nand U2172 (N_2172,N_1878,N_1908);
and U2173 (N_2173,N_1938,N_1952);
and U2174 (N_2174,N_1819,N_1824);
xor U2175 (N_2175,N_1813,N_1830);
nor U2176 (N_2176,N_1882,N_1936);
or U2177 (N_2177,N_1935,N_1854);
or U2178 (N_2178,N_1876,N_1884);
nand U2179 (N_2179,N_1924,N_1818);
and U2180 (N_2180,N_1811,N_1843);
nor U2181 (N_2181,N_1956,N_1997);
or U2182 (N_2182,N_1977,N_1801);
or U2183 (N_2183,N_1969,N_1946);
and U2184 (N_2184,N_1979,N_1909);
xnor U2185 (N_2185,N_1895,N_1848);
nand U2186 (N_2186,N_1853,N_1913);
nor U2187 (N_2187,N_1883,N_1945);
and U2188 (N_2188,N_1879,N_1960);
or U2189 (N_2189,N_1843,N_1848);
nand U2190 (N_2190,N_1832,N_1924);
or U2191 (N_2191,N_1929,N_1847);
and U2192 (N_2192,N_1981,N_1881);
or U2193 (N_2193,N_1857,N_1952);
or U2194 (N_2194,N_1933,N_1967);
xor U2195 (N_2195,N_1898,N_1948);
xnor U2196 (N_2196,N_1872,N_1867);
nand U2197 (N_2197,N_1943,N_1877);
xor U2198 (N_2198,N_1831,N_1889);
nor U2199 (N_2199,N_1878,N_1904);
or U2200 (N_2200,N_2049,N_2061);
xnor U2201 (N_2201,N_2059,N_2000);
nor U2202 (N_2202,N_2187,N_2137);
nand U2203 (N_2203,N_2180,N_2105);
and U2204 (N_2204,N_2173,N_2077);
xnor U2205 (N_2205,N_2177,N_2151);
or U2206 (N_2206,N_2158,N_2184);
or U2207 (N_2207,N_2074,N_2008);
nand U2208 (N_2208,N_2010,N_2035);
xor U2209 (N_2209,N_2024,N_2178);
xor U2210 (N_2210,N_2139,N_2124);
or U2211 (N_2211,N_2038,N_2018);
and U2212 (N_2212,N_2104,N_2051);
xnor U2213 (N_2213,N_2076,N_2075);
nand U2214 (N_2214,N_2007,N_2050);
xnor U2215 (N_2215,N_2183,N_2153);
and U2216 (N_2216,N_2176,N_2016);
and U2217 (N_2217,N_2055,N_2040);
xnor U2218 (N_2218,N_2067,N_2029);
xnor U2219 (N_2219,N_2172,N_2097);
xor U2220 (N_2220,N_2090,N_2193);
nor U2221 (N_2221,N_2045,N_2140);
xnor U2222 (N_2222,N_2047,N_2156);
or U2223 (N_2223,N_2135,N_2027);
xor U2224 (N_2224,N_2086,N_2098);
and U2225 (N_2225,N_2003,N_2071);
or U2226 (N_2226,N_2006,N_2128);
nor U2227 (N_2227,N_2068,N_2170);
nor U2228 (N_2228,N_2119,N_2033);
and U2229 (N_2229,N_2015,N_2191);
nand U2230 (N_2230,N_2113,N_2188);
nand U2231 (N_2231,N_2083,N_2081);
nor U2232 (N_2232,N_2195,N_2133);
or U2233 (N_2233,N_2123,N_2054);
and U2234 (N_2234,N_2174,N_2100);
or U2235 (N_2235,N_2053,N_2022);
and U2236 (N_2236,N_2002,N_2021);
and U2237 (N_2237,N_2162,N_2044);
nor U2238 (N_2238,N_2186,N_2102);
nor U2239 (N_2239,N_2175,N_2196);
xnor U2240 (N_2240,N_2046,N_2017);
nand U2241 (N_2241,N_2181,N_2080);
nand U2242 (N_2242,N_2088,N_2056);
nor U2243 (N_2243,N_2062,N_2145);
nand U2244 (N_2244,N_2111,N_2108);
and U2245 (N_2245,N_2093,N_2011);
nor U2246 (N_2246,N_2043,N_2060);
nand U2247 (N_2247,N_2157,N_2149);
xor U2248 (N_2248,N_2199,N_2122);
nand U2249 (N_2249,N_2130,N_2118);
nand U2250 (N_2250,N_2036,N_2079);
nand U2251 (N_2251,N_2089,N_2148);
or U2252 (N_2252,N_2095,N_2169);
nand U2253 (N_2253,N_2131,N_2078);
and U2254 (N_2254,N_2120,N_2037);
and U2255 (N_2255,N_2165,N_2161);
xnor U2256 (N_2256,N_2072,N_2099);
nand U2257 (N_2257,N_2185,N_2155);
xnor U2258 (N_2258,N_2144,N_2025);
xor U2259 (N_2259,N_2147,N_2064);
xor U2260 (N_2260,N_2114,N_2032);
or U2261 (N_2261,N_2082,N_2048);
nor U2262 (N_2262,N_2163,N_2063);
nor U2263 (N_2263,N_2031,N_2026);
nand U2264 (N_2264,N_2197,N_2092);
or U2265 (N_2265,N_2052,N_2101);
nand U2266 (N_2266,N_2109,N_2150);
xnor U2267 (N_2267,N_2106,N_2041);
and U2268 (N_2268,N_2009,N_2143);
or U2269 (N_2269,N_2152,N_2004);
or U2270 (N_2270,N_2034,N_2057);
nand U2271 (N_2271,N_2039,N_2073);
xnor U2272 (N_2272,N_2166,N_2091);
and U2273 (N_2273,N_2154,N_2189);
nor U2274 (N_2274,N_2069,N_2110);
or U2275 (N_2275,N_2085,N_2164);
or U2276 (N_2276,N_2117,N_2142);
nor U2277 (N_2277,N_2141,N_2094);
nor U2278 (N_2278,N_2146,N_2182);
or U2279 (N_2279,N_2058,N_2121);
nand U2280 (N_2280,N_2070,N_2013);
nor U2281 (N_2281,N_2160,N_2192);
and U2282 (N_2282,N_2066,N_2065);
xor U2283 (N_2283,N_2167,N_2001);
xor U2284 (N_2284,N_2028,N_2107);
nor U2285 (N_2285,N_2005,N_2136);
and U2286 (N_2286,N_2012,N_2014);
xor U2287 (N_2287,N_2084,N_2019);
nand U2288 (N_2288,N_2179,N_2168);
nor U2289 (N_2289,N_2194,N_2159);
or U2290 (N_2290,N_2126,N_2132);
nand U2291 (N_2291,N_2020,N_2116);
xor U2292 (N_2292,N_2087,N_2023);
xor U2293 (N_2293,N_2042,N_2190);
xnor U2294 (N_2294,N_2129,N_2138);
and U2295 (N_2295,N_2198,N_2112);
xor U2296 (N_2296,N_2103,N_2127);
nor U2297 (N_2297,N_2115,N_2134);
nand U2298 (N_2298,N_2030,N_2096);
nand U2299 (N_2299,N_2125,N_2171);
and U2300 (N_2300,N_2113,N_2155);
nand U2301 (N_2301,N_2101,N_2142);
nand U2302 (N_2302,N_2031,N_2094);
nand U2303 (N_2303,N_2187,N_2120);
and U2304 (N_2304,N_2051,N_2018);
nor U2305 (N_2305,N_2173,N_2135);
nor U2306 (N_2306,N_2171,N_2064);
nand U2307 (N_2307,N_2185,N_2131);
and U2308 (N_2308,N_2115,N_2004);
and U2309 (N_2309,N_2054,N_2103);
xor U2310 (N_2310,N_2059,N_2048);
nand U2311 (N_2311,N_2158,N_2094);
xor U2312 (N_2312,N_2094,N_2075);
nand U2313 (N_2313,N_2013,N_2027);
nor U2314 (N_2314,N_2037,N_2127);
nor U2315 (N_2315,N_2139,N_2134);
nand U2316 (N_2316,N_2101,N_2133);
or U2317 (N_2317,N_2138,N_2054);
xnor U2318 (N_2318,N_2115,N_2000);
nand U2319 (N_2319,N_2168,N_2143);
nor U2320 (N_2320,N_2084,N_2163);
or U2321 (N_2321,N_2190,N_2010);
and U2322 (N_2322,N_2194,N_2004);
and U2323 (N_2323,N_2032,N_2045);
nor U2324 (N_2324,N_2122,N_2144);
xor U2325 (N_2325,N_2006,N_2024);
and U2326 (N_2326,N_2189,N_2059);
nor U2327 (N_2327,N_2180,N_2151);
xnor U2328 (N_2328,N_2092,N_2075);
xor U2329 (N_2329,N_2150,N_2132);
and U2330 (N_2330,N_2113,N_2141);
nor U2331 (N_2331,N_2097,N_2006);
and U2332 (N_2332,N_2079,N_2125);
nand U2333 (N_2333,N_2193,N_2032);
or U2334 (N_2334,N_2035,N_2117);
nand U2335 (N_2335,N_2156,N_2128);
xor U2336 (N_2336,N_2083,N_2178);
nand U2337 (N_2337,N_2159,N_2055);
or U2338 (N_2338,N_2150,N_2143);
nand U2339 (N_2339,N_2025,N_2149);
nand U2340 (N_2340,N_2023,N_2083);
and U2341 (N_2341,N_2117,N_2006);
xor U2342 (N_2342,N_2026,N_2151);
nand U2343 (N_2343,N_2196,N_2015);
nor U2344 (N_2344,N_2152,N_2017);
and U2345 (N_2345,N_2038,N_2172);
or U2346 (N_2346,N_2108,N_2073);
nand U2347 (N_2347,N_2126,N_2016);
xnor U2348 (N_2348,N_2026,N_2023);
nor U2349 (N_2349,N_2016,N_2089);
nor U2350 (N_2350,N_2169,N_2160);
and U2351 (N_2351,N_2183,N_2031);
or U2352 (N_2352,N_2177,N_2133);
and U2353 (N_2353,N_2142,N_2024);
nor U2354 (N_2354,N_2062,N_2196);
and U2355 (N_2355,N_2047,N_2137);
nor U2356 (N_2356,N_2135,N_2105);
nand U2357 (N_2357,N_2019,N_2060);
nand U2358 (N_2358,N_2192,N_2051);
and U2359 (N_2359,N_2139,N_2058);
or U2360 (N_2360,N_2025,N_2125);
xnor U2361 (N_2361,N_2162,N_2065);
and U2362 (N_2362,N_2065,N_2076);
xor U2363 (N_2363,N_2015,N_2194);
nand U2364 (N_2364,N_2133,N_2031);
xor U2365 (N_2365,N_2043,N_2086);
nor U2366 (N_2366,N_2043,N_2092);
xnor U2367 (N_2367,N_2106,N_2144);
or U2368 (N_2368,N_2133,N_2053);
nor U2369 (N_2369,N_2119,N_2138);
nand U2370 (N_2370,N_2179,N_2066);
or U2371 (N_2371,N_2144,N_2183);
xor U2372 (N_2372,N_2151,N_2007);
or U2373 (N_2373,N_2090,N_2178);
or U2374 (N_2374,N_2083,N_2186);
or U2375 (N_2375,N_2137,N_2055);
or U2376 (N_2376,N_2016,N_2040);
nor U2377 (N_2377,N_2187,N_2194);
and U2378 (N_2378,N_2133,N_2139);
or U2379 (N_2379,N_2120,N_2192);
nand U2380 (N_2380,N_2177,N_2119);
or U2381 (N_2381,N_2166,N_2043);
xor U2382 (N_2382,N_2039,N_2097);
and U2383 (N_2383,N_2172,N_2006);
nor U2384 (N_2384,N_2009,N_2113);
nor U2385 (N_2385,N_2163,N_2168);
nand U2386 (N_2386,N_2064,N_2035);
nand U2387 (N_2387,N_2004,N_2104);
xor U2388 (N_2388,N_2117,N_2098);
nor U2389 (N_2389,N_2011,N_2021);
xor U2390 (N_2390,N_2029,N_2081);
and U2391 (N_2391,N_2078,N_2112);
nor U2392 (N_2392,N_2058,N_2191);
nand U2393 (N_2393,N_2196,N_2048);
xnor U2394 (N_2394,N_2162,N_2190);
and U2395 (N_2395,N_2016,N_2066);
nand U2396 (N_2396,N_2183,N_2128);
nor U2397 (N_2397,N_2169,N_2064);
nand U2398 (N_2398,N_2154,N_2068);
xor U2399 (N_2399,N_2026,N_2186);
nor U2400 (N_2400,N_2243,N_2330);
or U2401 (N_2401,N_2312,N_2230);
nand U2402 (N_2402,N_2376,N_2293);
or U2403 (N_2403,N_2358,N_2244);
nand U2404 (N_2404,N_2207,N_2281);
and U2405 (N_2405,N_2300,N_2276);
or U2406 (N_2406,N_2348,N_2394);
nor U2407 (N_2407,N_2211,N_2323);
and U2408 (N_2408,N_2246,N_2256);
nand U2409 (N_2409,N_2272,N_2327);
nand U2410 (N_2410,N_2343,N_2324);
and U2411 (N_2411,N_2236,N_2255);
nor U2412 (N_2412,N_2303,N_2325);
xnor U2413 (N_2413,N_2223,N_2264);
or U2414 (N_2414,N_2310,N_2205);
nor U2415 (N_2415,N_2347,N_2260);
nor U2416 (N_2416,N_2289,N_2284);
or U2417 (N_2417,N_2268,N_2353);
and U2418 (N_2418,N_2209,N_2302);
and U2419 (N_2419,N_2322,N_2228);
xnor U2420 (N_2420,N_2317,N_2235);
xor U2421 (N_2421,N_2263,N_2399);
and U2422 (N_2422,N_2292,N_2380);
nor U2423 (N_2423,N_2231,N_2372);
nand U2424 (N_2424,N_2252,N_2392);
xor U2425 (N_2425,N_2349,N_2378);
xor U2426 (N_2426,N_2237,N_2224);
nor U2427 (N_2427,N_2249,N_2368);
or U2428 (N_2428,N_2297,N_2308);
or U2429 (N_2429,N_2233,N_2200);
or U2430 (N_2430,N_2339,N_2395);
nor U2431 (N_2431,N_2337,N_2332);
or U2432 (N_2432,N_2356,N_2221);
nor U2433 (N_2433,N_2383,N_2393);
xor U2434 (N_2434,N_2258,N_2273);
or U2435 (N_2435,N_2363,N_2384);
xor U2436 (N_2436,N_2329,N_2321);
nor U2437 (N_2437,N_2307,N_2241);
and U2438 (N_2438,N_2288,N_2257);
or U2439 (N_2439,N_2346,N_2261);
or U2440 (N_2440,N_2355,N_2240);
nand U2441 (N_2441,N_2309,N_2374);
xnor U2442 (N_2442,N_2352,N_2301);
or U2443 (N_2443,N_2328,N_2359);
and U2444 (N_2444,N_2253,N_2334);
nor U2445 (N_2445,N_2286,N_2385);
nand U2446 (N_2446,N_2345,N_2280);
nand U2447 (N_2447,N_2217,N_2298);
xor U2448 (N_2448,N_2282,N_2371);
and U2449 (N_2449,N_2215,N_2338);
nor U2450 (N_2450,N_2204,N_2283);
nor U2451 (N_2451,N_2214,N_2262);
nand U2452 (N_2452,N_2396,N_2218);
and U2453 (N_2453,N_2270,N_2340);
xor U2454 (N_2454,N_2361,N_2234);
or U2455 (N_2455,N_2344,N_2266);
and U2456 (N_2456,N_2357,N_2320);
and U2457 (N_2457,N_2203,N_2294);
xnor U2458 (N_2458,N_2222,N_2375);
nand U2459 (N_2459,N_2342,N_2350);
nand U2460 (N_2460,N_2201,N_2202);
nor U2461 (N_2461,N_2387,N_2351);
nand U2462 (N_2462,N_2265,N_2238);
nor U2463 (N_2463,N_2326,N_2366);
nor U2464 (N_2464,N_2239,N_2295);
nor U2465 (N_2465,N_2247,N_2386);
xor U2466 (N_2466,N_2373,N_2269);
or U2467 (N_2467,N_2381,N_2336);
and U2468 (N_2468,N_2274,N_2277);
xnor U2469 (N_2469,N_2227,N_2219);
nor U2470 (N_2470,N_2305,N_2254);
and U2471 (N_2471,N_2341,N_2314);
xor U2472 (N_2472,N_2212,N_2210);
nand U2473 (N_2473,N_2316,N_2291);
nor U2474 (N_2474,N_2206,N_2335);
and U2475 (N_2475,N_2319,N_2331);
and U2476 (N_2476,N_2259,N_2296);
and U2477 (N_2477,N_2354,N_2248);
nor U2478 (N_2478,N_2390,N_2397);
or U2479 (N_2479,N_2232,N_2364);
or U2480 (N_2480,N_2220,N_2365);
and U2481 (N_2481,N_2279,N_2275);
or U2482 (N_2482,N_2290,N_2333);
or U2483 (N_2483,N_2278,N_2318);
nand U2484 (N_2484,N_2267,N_2245);
or U2485 (N_2485,N_2299,N_2391);
nand U2486 (N_2486,N_2377,N_2362);
nand U2487 (N_2487,N_2398,N_2304);
nor U2488 (N_2488,N_2229,N_2287);
and U2489 (N_2489,N_2315,N_2226);
xnor U2490 (N_2490,N_2369,N_2388);
or U2491 (N_2491,N_2379,N_2225);
xnor U2492 (N_2492,N_2313,N_2251);
nand U2493 (N_2493,N_2250,N_2213);
xor U2494 (N_2494,N_2370,N_2360);
and U2495 (N_2495,N_2216,N_2271);
and U2496 (N_2496,N_2208,N_2285);
and U2497 (N_2497,N_2311,N_2242);
nor U2498 (N_2498,N_2306,N_2382);
and U2499 (N_2499,N_2367,N_2389);
or U2500 (N_2500,N_2361,N_2350);
xor U2501 (N_2501,N_2382,N_2284);
nand U2502 (N_2502,N_2300,N_2327);
and U2503 (N_2503,N_2288,N_2237);
nand U2504 (N_2504,N_2264,N_2214);
nand U2505 (N_2505,N_2341,N_2255);
nor U2506 (N_2506,N_2350,N_2366);
or U2507 (N_2507,N_2220,N_2372);
nand U2508 (N_2508,N_2263,N_2256);
or U2509 (N_2509,N_2243,N_2278);
xor U2510 (N_2510,N_2339,N_2382);
nand U2511 (N_2511,N_2228,N_2254);
and U2512 (N_2512,N_2343,N_2252);
and U2513 (N_2513,N_2312,N_2329);
nor U2514 (N_2514,N_2397,N_2298);
and U2515 (N_2515,N_2337,N_2238);
or U2516 (N_2516,N_2246,N_2236);
nand U2517 (N_2517,N_2342,N_2361);
nand U2518 (N_2518,N_2327,N_2285);
and U2519 (N_2519,N_2206,N_2275);
or U2520 (N_2520,N_2208,N_2310);
and U2521 (N_2521,N_2321,N_2268);
nor U2522 (N_2522,N_2230,N_2347);
and U2523 (N_2523,N_2342,N_2209);
nand U2524 (N_2524,N_2278,N_2205);
xnor U2525 (N_2525,N_2313,N_2299);
nor U2526 (N_2526,N_2291,N_2343);
or U2527 (N_2527,N_2237,N_2340);
and U2528 (N_2528,N_2393,N_2205);
nor U2529 (N_2529,N_2245,N_2305);
and U2530 (N_2530,N_2265,N_2213);
nand U2531 (N_2531,N_2322,N_2255);
nor U2532 (N_2532,N_2239,N_2311);
xor U2533 (N_2533,N_2369,N_2206);
nand U2534 (N_2534,N_2340,N_2242);
nand U2535 (N_2535,N_2203,N_2253);
or U2536 (N_2536,N_2254,N_2358);
nor U2537 (N_2537,N_2318,N_2315);
nor U2538 (N_2538,N_2299,N_2379);
and U2539 (N_2539,N_2205,N_2295);
xnor U2540 (N_2540,N_2223,N_2330);
xor U2541 (N_2541,N_2244,N_2368);
xnor U2542 (N_2542,N_2248,N_2332);
nor U2543 (N_2543,N_2297,N_2357);
and U2544 (N_2544,N_2370,N_2206);
and U2545 (N_2545,N_2302,N_2389);
xnor U2546 (N_2546,N_2232,N_2288);
or U2547 (N_2547,N_2310,N_2370);
xnor U2548 (N_2548,N_2250,N_2367);
or U2549 (N_2549,N_2300,N_2282);
xor U2550 (N_2550,N_2393,N_2282);
nand U2551 (N_2551,N_2236,N_2229);
nor U2552 (N_2552,N_2366,N_2338);
nand U2553 (N_2553,N_2232,N_2276);
nor U2554 (N_2554,N_2374,N_2305);
xor U2555 (N_2555,N_2301,N_2387);
nor U2556 (N_2556,N_2304,N_2298);
nand U2557 (N_2557,N_2349,N_2231);
xor U2558 (N_2558,N_2346,N_2332);
xor U2559 (N_2559,N_2302,N_2351);
and U2560 (N_2560,N_2236,N_2288);
xor U2561 (N_2561,N_2287,N_2239);
xor U2562 (N_2562,N_2394,N_2378);
nor U2563 (N_2563,N_2316,N_2200);
and U2564 (N_2564,N_2352,N_2238);
nand U2565 (N_2565,N_2266,N_2214);
xor U2566 (N_2566,N_2364,N_2345);
xor U2567 (N_2567,N_2278,N_2237);
or U2568 (N_2568,N_2365,N_2344);
or U2569 (N_2569,N_2356,N_2286);
nor U2570 (N_2570,N_2219,N_2365);
and U2571 (N_2571,N_2383,N_2281);
and U2572 (N_2572,N_2334,N_2378);
or U2573 (N_2573,N_2313,N_2352);
xnor U2574 (N_2574,N_2365,N_2241);
nand U2575 (N_2575,N_2276,N_2320);
nor U2576 (N_2576,N_2277,N_2315);
nor U2577 (N_2577,N_2259,N_2269);
and U2578 (N_2578,N_2258,N_2226);
and U2579 (N_2579,N_2270,N_2368);
or U2580 (N_2580,N_2232,N_2389);
or U2581 (N_2581,N_2327,N_2227);
nor U2582 (N_2582,N_2265,N_2232);
nand U2583 (N_2583,N_2379,N_2341);
or U2584 (N_2584,N_2393,N_2215);
or U2585 (N_2585,N_2360,N_2201);
or U2586 (N_2586,N_2211,N_2390);
xnor U2587 (N_2587,N_2328,N_2300);
or U2588 (N_2588,N_2253,N_2240);
nor U2589 (N_2589,N_2230,N_2367);
xor U2590 (N_2590,N_2342,N_2313);
or U2591 (N_2591,N_2216,N_2375);
nor U2592 (N_2592,N_2284,N_2387);
or U2593 (N_2593,N_2260,N_2248);
nand U2594 (N_2594,N_2246,N_2350);
and U2595 (N_2595,N_2259,N_2311);
xnor U2596 (N_2596,N_2336,N_2325);
xor U2597 (N_2597,N_2213,N_2298);
nand U2598 (N_2598,N_2304,N_2271);
nor U2599 (N_2599,N_2354,N_2366);
and U2600 (N_2600,N_2423,N_2472);
or U2601 (N_2601,N_2470,N_2494);
and U2602 (N_2602,N_2435,N_2443);
or U2603 (N_2603,N_2580,N_2542);
nand U2604 (N_2604,N_2469,N_2444);
xor U2605 (N_2605,N_2438,N_2520);
and U2606 (N_2606,N_2499,N_2473);
or U2607 (N_2607,N_2552,N_2549);
nor U2608 (N_2608,N_2431,N_2554);
and U2609 (N_2609,N_2433,N_2486);
nand U2610 (N_2610,N_2572,N_2512);
or U2611 (N_2611,N_2418,N_2555);
nand U2612 (N_2612,N_2599,N_2597);
or U2613 (N_2613,N_2461,N_2578);
nand U2614 (N_2614,N_2491,N_2452);
and U2615 (N_2615,N_2592,N_2583);
or U2616 (N_2616,N_2407,N_2574);
nor U2617 (N_2617,N_2403,N_2519);
and U2618 (N_2618,N_2576,N_2485);
and U2619 (N_2619,N_2594,N_2406);
nand U2620 (N_2620,N_2568,N_2563);
or U2621 (N_2621,N_2544,N_2500);
xor U2622 (N_2622,N_2454,N_2510);
and U2623 (N_2623,N_2489,N_2573);
nand U2624 (N_2624,N_2593,N_2532);
nand U2625 (N_2625,N_2577,N_2450);
xor U2626 (N_2626,N_2537,N_2515);
or U2627 (N_2627,N_2547,N_2501);
or U2628 (N_2628,N_2558,N_2527);
nor U2629 (N_2629,N_2458,N_2462);
and U2630 (N_2630,N_2447,N_2405);
nor U2631 (N_2631,N_2587,N_2411);
nand U2632 (N_2632,N_2595,N_2449);
and U2633 (N_2633,N_2508,N_2457);
nor U2634 (N_2634,N_2586,N_2495);
nand U2635 (N_2635,N_2582,N_2585);
or U2636 (N_2636,N_2548,N_2451);
or U2637 (N_2637,N_2562,N_2480);
nor U2638 (N_2638,N_2584,N_2401);
xor U2639 (N_2639,N_2538,N_2456);
xnor U2640 (N_2640,N_2497,N_2476);
nor U2641 (N_2641,N_2565,N_2477);
nor U2642 (N_2642,N_2579,N_2455);
or U2643 (N_2643,N_2517,N_2468);
nor U2644 (N_2644,N_2530,N_2424);
nor U2645 (N_2645,N_2531,N_2509);
xor U2646 (N_2646,N_2536,N_2570);
xor U2647 (N_2647,N_2414,N_2591);
xor U2648 (N_2648,N_2541,N_2463);
or U2649 (N_2649,N_2581,N_2404);
xor U2650 (N_2650,N_2417,N_2483);
or U2651 (N_2651,N_2429,N_2420);
nand U2652 (N_2652,N_2566,N_2409);
nand U2653 (N_2653,N_2416,N_2422);
nand U2654 (N_2654,N_2434,N_2569);
nor U2655 (N_2655,N_2564,N_2419);
and U2656 (N_2656,N_2464,N_2553);
xnor U2657 (N_2657,N_2410,N_2430);
or U2658 (N_2658,N_2557,N_2513);
or U2659 (N_2659,N_2448,N_2493);
or U2660 (N_2660,N_2425,N_2521);
xnor U2661 (N_2661,N_2432,N_2534);
nor U2662 (N_2662,N_2545,N_2488);
nor U2663 (N_2663,N_2441,N_2507);
and U2664 (N_2664,N_2465,N_2487);
nand U2665 (N_2665,N_2561,N_2421);
nor U2666 (N_2666,N_2467,N_2551);
nand U2667 (N_2667,N_2596,N_2540);
nand U2668 (N_2668,N_2475,N_2539);
nand U2669 (N_2669,N_2560,N_2439);
nand U2670 (N_2670,N_2567,N_2484);
and U2671 (N_2671,N_2524,N_2466);
xor U2672 (N_2672,N_2550,N_2498);
nor U2673 (N_2673,N_2529,N_2459);
nand U2674 (N_2674,N_2511,N_2492);
nor U2675 (N_2675,N_2543,N_2479);
nor U2676 (N_2676,N_2481,N_2496);
nor U2677 (N_2677,N_2526,N_2506);
and U2678 (N_2678,N_2598,N_2460);
nor U2679 (N_2679,N_2490,N_2436);
nor U2680 (N_2680,N_2559,N_2535);
nand U2681 (N_2681,N_2525,N_2445);
nand U2682 (N_2682,N_2428,N_2588);
nor U2683 (N_2683,N_2528,N_2590);
or U2684 (N_2684,N_2504,N_2505);
and U2685 (N_2685,N_2402,N_2478);
xor U2686 (N_2686,N_2482,N_2533);
and U2687 (N_2687,N_2412,N_2437);
and U2688 (N_2688,N_2446,N_2503);
nand U2689 (N_2689,N_2589,N_2453);
xor U2690 (N_2690,N_2514,N_2427);
nor U2691 (N_2691,N_2575,N_2518);
and U2692 (N_2692,N_2400,N_2408);
nor U2693 (N_2693,N_2546,N_2523);
nor U2694 (N_2694,N_2442,N_2474);
nor U2695 (N_2695,N_2415,N_2471);
xor U2696 (N_2696,N_2440,N_2556);
xor U2697 (N_2697,N_2413,N_2522);
and U2698 (N_2698,N_2502,N_2571);
xor U2699 (N_2699,N_2516,N_2426);
and U2700 (N_2700,N_2575,N_2431);
nand U2701 (N_2701,N_2586,N_2428);
nand U2702 (N_2702,N_2555,N_2403);
or U2703 (N_2703,N_2406,N_2400);
and U2704 (N_2704,N_2481,N_2508);
or U2705 (N_2705,N_2595,N_2410);
and U2706 (N_2706,N_2460,N_2490);
and U2707 (N_2707,N_2589,N_2513);
nor U2708 (N_2708,N_2558,N_2438);
xor U2709 (N_2709,N_2524,N_2579);
or U2710 (N_2710,N_2507,N_2402);
nand U2711 (N_2711,N_2519,N_2495);
nand U2712 (N_2712,N_2436,N_2523);
xor U2713 (N_2713,N_2438,N_2578);
nand U2714 (N_2714,N_2590,N_2597);
and U2715 (N_2715,N_2411,N_2466);
or U2716 (N_2716,N_2409,N_2591);
or U2717 (N_2717,N_2575,N_2400);
or U2718 (N_2718,N_2475,N_2410);
nand U2719 (N_2719,N_2500,N_2512);
and U2720 (N_2720,N_2427,N_2451);
nor U2721 (N_2721,N_2552,N_2572);
nor U2722 (N_2722,N_2463,N_2529);
or U2723 (N_2723,N_2443,N_2474);
nand U2724 (N_2724,N_2501,N_2471);
xnor U2725 (N_2725,N_2422,N_2575);
or U2726 (N_2726,N_2455,N_2540);
and U2727 (N_2727,N_2474,N_2590);
xnor U2728 (N_2728,N_2494,N_2409);
nand U2729 (N_2729,N_2441,N_2492);
xnor U2730 (N_2730,N_2434,N_2461);
and U2731 (N_2731,N_2472,N_2444);
nand U2732 (N_2732,N_2460,N_2544);
nand U2733 (N_2733,N_2424,N_2486);
or U2734 (N_2734,N_2512,N_2513);
or U2735 (N_2735,N_2498,N_2418);
nor U2736 (N_2736,N_2509,N_2508);
and U2737 (N_2737,N_2429,N_2492);
or U2738 (N_2738,N_2432,N_2516);
nand U2739 (N_2739,N_2540,N_2502);
nand U2740 (N_2740,N_2416,N_2444);
and U2741 (N_2741,N_2498,N_2466);
and U2742 (N_2742,N_2463,N_2570);
xor U2743 (N_2743,N_2495,N_2492);
and U2744 (N_2744,N_2406,N_2550);
or U2745 (N_2745,N_2562,N_2411);
and U2746 (N_2746,N_2438,N_2493);
and U2747 (N_2747,N_2499,N_2523);
nand U2748 (N_2748,N_2464,N_2575);
xor U2749 (N_2749,N_2596,N_2409);
xor U2750 (N_2750,N_2446,N_2534);
xor U2751 (N_2751,N_2532,N_2424);
nor U2752 (N_2752,N_2411,N_2464);
and U2753 (N_2753,N_2534,N_2482);
nand U2754 (N_2754,N_2585,N_2593);
xor U2755 (N_2755,N_2573,N_2567);
xor U2756 (N_2756,N_2554,N_2574);
and U2757 (N_2757,N_2572,N_2539);
or U2758 (N_2758,N_2549,N_2485);
nor U2759 (N_2759,N_2516,N_2465);
nor U2760 (N_2760,N_2555,N_2597);
nor U2761 (N_2761,N_2568,N_2400);
xor U2762 (N_2762,N_2588,N_2537);
or U2763 (N_2763,N_2467,N_2417);
or U2764 (N_2764,N_2556,N_2446);
and U2765 (N_2765,N_2422,N_2424);
xor U2766 (N_2766,N_2529,N_2474);
nand U2767 (N_2767,N_2430,N_2434);
or U2768 (N_2768,N_2590,N_2574);
xor U2769 (N_2769,N_2519,N_2595);
nor U2770 (N_2770,N_2537,N_2582);
or U2771 (N_2771,N_2470,N_2596);
nor U2772 (N_2772,N_2592,N_2507);
or U2773 (N_2773,N_2502,N_2552);
and U2774 (N_2774,N_2520,N_2599);
or U2775 (N_2775,N_2563,N_2573);
nand U2776 (N_2776,N_2437,N_2491);
nor U2777 (N_2777,N_2469,N_2507);
nand U2778 (N_2778,N_2430,N_2545);
or U2779 (N_2779,N_2594,N_2434);
xor U2780 (N_2780,N_2556,N_2439);
nand U2781 (N_2781,N_2575,N_2441);
nor U2782 (N_2782,N_2477,N_2548);
and U2783 (N_2783,N_2590,N_2505);
and U2784 (N_2784,N_2516,N_2538);
xnor U2785 (N_2785,N_2517,N_2525);
nand U2786 (N_2786,N_2551,N_2413);
nor U2787 (N_2787,N_2442,N_2434);
nand U2788 (N_2788,N_2479,N_2434);
and U2789 (N_2789,N_2522,N_2504);
and U2790 (N_2790,N_2504,N_2542);
nand U2791 (N_2791,N_2592,N_2458);
and U2792 (N_2792,N_2534,N_2566);
nand U2793 (N_2793,N_2532,N_2516);
or U2794 (N_2794,N_2587,N_2426);
and U2795 (N_2795,N_2473,N_2563);
and U2796 (N_2796,N_2538,N_2469);
and U2797 (N_2797,N_2445,N_2549);
nor U2798 (N_2798,N_2448,N_2572);
xnor U2799 (N_2799,N_2532,N_2441);
xnor U2800 (N_2800,N_2650,N_2692);
nor U2801 (N_2801,N_2716,N_2701);
and U2802 (N_2802,N_2667,N_2649);
xor U2803 (N_2803,N_2636,N_2628);
xor U2804 (N_2804,N_2654,N_2708);
nand U2805 (N_2805,N_2767,N_2675);
xor U2806 (N_2806,N_2647,N_2691);
and U2807 (N_2807,N_2602,N_2683);
and U2808 (N_2808,N_2601,N_2603);
and U2809 (N_2809,N_2705,N_2612);
nor U2810 (N_2810,N_2702,N_2617);
nor U2811 (N_2811,N_2773,N_2789);
xnor U2812 (N_2812,N_2720,N_2693);
nand U2813 (N_2813,N_2787,N_2726);
and U2814 (N_2814,N_2686,N_2724);
nor U2815 (N_2815,N_2652,N_2729);
nand U2816 (N_2816,N_2673,N_2710);
nand U2817 (N_2817,N_2674,N_2769);
xnor U2818 (N_2818,N_2732,N_2658);
xnor U2819 (N_2819,N_2754,N_2662);
and U2820 (N_2820,N_2608,N_2728);
xor U2821 (N_2821,N_2753,N_2718);
or U2822 (N_2822,N_2605,N_2611);
and U2823 (N_2823,N_2719,N_2661);
and U2824 (N_2824,N_2759,N_2666);
nor U2825 (N_2825,N_2723,N_2743);
xor U2826 (N_2826,N_2788,N_2768);
xor U2827 (N_2827,N_2707,N_2737);
or U2828 (N_2828,N_2755,N_2614);
nor U2829 (N_2829,N_2796,N_2615);
xnor U2830 (N_2830,N_2681,N_2797);
xnor U2831 (N_2831,N_2643,N_2697);
and U2832 (N_2832,N_2688,N_2791);
nand U2833 (N_2833,N_2786,N_2669);
nor U2834 (N_2834,N_2704,N_2727);
and U2835 (N_2835,N_2740,N_2757);
or U2836 (N_2836,N_2607,N_2721);
xor U2837 (N_2837,N_2616,N_2656);
and U2838 (N_2838,N_2741,N_2633);
xnor U2839 (N_2839,N_2785,N_2766);
or U2840 (N_2840,N_2752,N_2709);
nor U2841 (N_2841,N_2635,N_2776);
or U2842 (N_2842,N_2779,N_2792);
and U2843 (N_2843,N_2610,N_2751);
xor U2844 (N_2844,N_2622,N_2657);
and U2845 (N_2845,N_2618,N_2627);
nor U2846 (N_2846,N_2665,N_2745);
nor U2847 (N_2847,N_2749,N_2756);
nand U2848 (N_2848,N_2730,N_2680);
xor U2849 (N_2849,N_2774,N_2638);
and U2850 (N_2850,N_2758,N_2700);
xor U2851 (N_2851,N_2735,N_2762);
and U2852 (N_2852,N_2696,N_2750);
xnor U2853 (N_2853,N_2690,N_2760);
nor U2854 (N_2854,N_2623,N_2703);
nor U2855 (N_2855,N_2670,N_2798);
nor U2856 (N_2856,N_2624,N_2770);
nand U2857 (N_2857,N_2699,N_2793);
nor U2858 (N_2858,N_2712,N_2738);
nand U2859 (N_2859,N_2715,N_2634);
nand U2860 (N_2860,N_2799,N_2604);
and U2861 (N_2861,N_2678,N_2748);
xor U2862 (N_2862,N_2717,N_2777);
nand U2863 (N_2863,N_2668,N_2642);
nor U2864 (N_2864,N_2713,N_2694);
xnor U2865 (N_2865,N_2664,N_2641);
nor U2866 (N_2866,N_2646,N_2653);
nand U2867 (N_2867,N_2706,N_2744);
or U2868 (N_2868,N_2734,N_2725);
and U2869 (N_2869,N_2687,N_2640);
nor U2870 (N_2870,N_2606,N_2763);
or U2871 (N_2871,N_2764,N_2742);
xor U2872 (N_2872,N_2739,N_2682);
xnor U2873 (N_2873,N_2651,N_2600);
or U2874 (N_2874,N_2632,N_2761);
xnor U2875 (N_2875,N_2684,N_2648);
nand U2876 (N_2876,N_2639,N_2689);
and U2877 (N_2877,N_2631,N_2771);
nor U2878 (N_2878,N_2629,N_2626);
nor U2879 (N_2879,N_2772,N_2609);
nor U2880 (N_2880,N_2722,N_2711);
and U2881 (N_2881,N_2677,N_2765);
or U2882 (N_2882,N_2625,N_2795);
xor U2883 (N_2883,N_2731,N_2695);
xnor U2884 (N_2884,N_2794,N_2747);
xnor U2885 (N_2885,N_2676,N_2775);
or U2886 (N_2886,N_2630,N_2746);
nor U2887 (N_2887,N_2679,N_2637);
nand U2888 (N_2888,N_2698,N_2781);
xnor U2889 (N_2889,N_2663,N_2655);
xor U2890 (N_2890,N_2685,N_2671);
and U2891 (N_2891,N_2736,N_2645);
nor U2892 (N_2892,N_2782,N_2672);
nor U2893 (N_2893,N_2644,N_2780);
xnor U2894 (N_2894,N_2778,N_2619);
nand U2895 (N_2895,N_2621,N_2784);
nand U2896 (N_2896,N_2790,N_2620);
nor U2897 (N_2897,N_2714,N_2733);
nand U2898 (N_2898,N_2613,N_2783);
or U2899 (N_2899,N_2660,N_2659);
xor U2900 (N_2900,N_2772,N_2662);
or U2901 (N_2901,N_2612,N_2778);
nor U2902 (N_2902,N_2705,N_2684);
xnor U2903 (N_2903,N_2647,N_2715);
nand U2904 (N_2904,N_2710,N_2625);
and U2905 (N_2905,N_2629,N_2781);
nand U2906 (N_2906,N_2709,N_2753);
and U2907 (N_2907,N_2629,N_2780);
nand U2908 (N_2908,N_2684,N_2729);
or U2909 (N_2909,N_2688,N_2646);
nand U2910 (N_2910,N_2767,N_2793);
nor U2911 (N_2911,N_2622,N_2728);
xnor U2912 (N_2912,N_2665,N_2769);
or U2913 (N_2913,N_2732,N_2760);
nor U2914 (N_2914,N_2651,N_2622);
and U2915 (N_2915,N_2764,N_2781);
nor U2916 (N_2916,N_2671,N_2607);
and U2917 (N_2917,N_2722,N_2643);
and U2918 (N_2918,N_2733,N_2693);
nand U2919 (N_2919,N_2600,N_2729);
and U2920 (N_2920,N_2792,N_2738);
nand U2921 (N_2921,N_2645,N_2795);
nand U2922 (N_2922,N_2687,N_2652);
and U2923 (N_2923,N_2770,N_2721);
or U2924 (N_2924,N_2781,N_2748);
nor U2925 (N_2925,N_2792,N_2734);
nor U2926 (N_2926,N_2644,N_2778);
or U2927 (N_2927,N_2619,N_2615);
xnor U2928 (N_2928,N_2614,N_2600);
and U2929 (N_2929,N_2727,N_2743);
xnor U2930 (N_2930,N_2776,N_2783);
nand U2931 (N_2931,N_2625,N_2684);
xnor U2932 (N_2932,N_2777,N_2781);
or U2933 (N_2933,N_2730,N_2711);
xor U2934 (N_2934,N_2619,N_2621);
and U2935 (N_2935,N_2699,N_2688);
nor U2936 (N_2936,N_2777,N_2656);
and U2937 (N_2937,N_2717,N_2651);
xnor U2938 (N_2938,N_2724,N_2634);
and U2939 (N_2939,N_2642,N_2693);
nand U2940 (N_2940,N_2675,N_2795);
and U2941 (N_2941,N_2648,N_2625);
or U2942 (N_2942,N_2783,N_2625);
nor U2943 (N_2943,N_2635,N_2706);
or U2944 (N_2944,N_2724,N_2640);
nor U2945 (N_2945,N_2733,N_2748);
nor U2946 (N_2946,N_2642,N_2630);
nand U2947 (N_2947,N_2614,N_2677);
or U2948 (N_2948,N_2780,N_2678);
and U2949 (N_2949,N_2745,N_2686);
nor U2950 (N_2950,N_2791,N_2675);
xor U2951 (N_2951,N_2769,N_2627);
nand U2952 (N_2952,N_2779,N_2767);
or U2953 (N_2953,N_2674,N_2795);
xnor U2954 (N_2954,N_2720,N_2677);
and U2955 (N_2955,N_2610,N_2668);
and U2956 (N_2956,N_2748,N_2715);
nand U2957 (N_2957,N_2661,N_2600);
nand U2958 (N_2958,N_2696,N_2717);
and U2959 (N_2959,N_2657,N_2691);
xor U2960 (N_2960,N_2754,N_2683);
or U2961 (N_2961,N_2723,N_2774);
xor U2962 (N_2962,N_2711,N_2647);
and U2963 (N_2963,N_2675,N_2650);
xor U2964 (N_2964,N_2667,N_2618);
or U2965 (N_2965,N_2696,N_2612);
and U2966 (N_2966,N_2645,N_2655);
xor U2967 (N_2967,N_2705,N_2665);
xor U2968 (N_2968,N_2645,N_2783);
nand U2969 (N_2969,N_2637,N_2646);
nand U2970 (N_2970,N_2683,N_2713);
or U2971 (N_2971,N_2697,N_2671);
xor U2972 (N_2972,N_2647,N_2713);
and U2973 (N_2973,N_2711,N_2664);
xor U2974 (N_2974,N_2716,N_2611);
or U2975 (N_2975,N_2768,N_2671);
xnor U2976 (N_2976,N_2659,N_2675);
or U2977 (N_2977,N_2604,N_2728);
and U2978 (N_2978,N_2605,N_2637);
or U2979 (N_2979,N_2716,N_2770);
nand U2980 (N_2980,N_2765,N_2678);
nand U2981 (N_2981,N_2661,N_2702);
xor U2982 (N_2982,N_2607,N_2723);
xnor U2983 (N_2983,N_2616,N_2785);
or U2984 (N_2984,N_2665,N_2724);
nor U2985 (N_2985,N_2618,N_2695);
nand U2986 (N_2986,N_2623,N_2644);
or U2987 (N_2987,N_2699,N_2658);
nor U2988 (N_2988,N_2689,N_2737);
xor U2989 (N_2989,N_2740,N_2703);
nor U2990 (N_2990,N_2735,N_2667);
nor U2991 (N_2991,N_2683,N_2758);
and U2992 (N_2992,N_2672,N_2744);
xor U2993 (N_2993,N_2682,N_2686);
and U2994 (N_2994,N_2639,N_2718);
or U2995 (N_2995,N_2775,N_2751);
and U2996 (N_2996,N_2772,N_2625);
and U2997 (N_2997,N_2690,N_2628);
nand U2998 (N_2998,N_2695,N_2761);
nor U2999 (N_2999,N_2679,N_2629);
xor U3000 (N_3000,N_2990,N_2952);
xnor U3001 (N_3001,N_2951,N_2869);
and U3002 (N_3002,N_2837,N_2859);
nand U3003 (N_3003,N_2899,N_2875);
nor U3004 (N_3004,N_2846,N_2957);
or U3005 (N_3005,N_2840,N_2880);
or U3006 (N_3006,N_2820,N_2913);
and U3007 (N_3007,N_2860,N_2973);
nor U3008 (N_3008,N_2904,N_2924);
nor U3009 (N_3009,N_2809,N_2864);
xnor U3010 (N_3010,N_2877,N_2812);
xor U3011 (N_3011,N_2898,N_2953);
or U3012 (N_3012,N_2964,N_2982);
and U3013 (N_3013,N_2976,N_2802);
nor U3014 (N_3014,N_2863,N_2977);
nand U3015 (N_3015,N_2969,N_2935);
nand U3016 (N_3016,N_2984,N_2878);
or U3017 (N_3017,N_2821,N_2813);
xnor U3018 (N_3018,N_2845,N_2816);
xor U3019 (N_3019,N_2841,N_2865);
nor U3020 (N_3020,N_2942,N_2822);
nor U3021 (N_3021,N_2808,N_2823);
and U3022 (N_3022,N_2858,N_2872);
xnor U3023 (N_3023,N_2893,N_2938);
xnor U3024 (N_3024,N_2826,N_2804);
or U3025 (N_3025,N_2810,N_2932);
nor U3026 (N_3026,N_2896,N_2906);
nand U3027 (N_3027,N_2879,N_2931);
nor U3028 (N_3028,N_2948,N_2834);
and U3029 (N_3029,N_2882,N_2980);
and U3030 (N_3030,N_2881,N_2936);
nor U3031 (N_3031,N_2828,N_2968);
xor U3032 (N_3032,N_2824,N_2836);
and U3033 (N_3033,N_2844,N_2926);
nor U3034 (N_3034,N_2850,N_2832);
and U3035 (N_3035,N_2999,N_2966);
xor U3036 (N_3036,N_2974,N_2944);
and U3037 (N_3037,N_2928,N_2890);
nor U3038 (N_3038,N_2909,N_2993);
or U3039 (N_3039,N_2914,N_2908);
and U3040 (N_3040,N_2815,N_2852);
nand U3041 (N_3041,N_2986,N_2866);
or U3042 (N_3042,N_2918,N_2949);
nand U3043 (N_3043,N_2996,N_2994);
nor U3044 (N_3044,N_2857,N_2922);
xor U3045 (N_3045,N_2870,N_2958);
nand U3046 (N_3046,N_2916,N_2934);
xor U3047 (N_3047,N_2970,N_2997);
xnor U3048 (N_3048,N_2972,N_2847);
or U3049 (N_3049,N_2800,N_2917);
or U3050 (N_3050,N_2983,N_2897);
nand U3051 (N_3051,N_2954,N_2910);
nor U3052 (N_3052,N_2987,N_2831);
xor U3053 (N_3053,N_2874,N_2939);
and U3054 (N_3054,N_2903,N_2923);
xor U3055 (N_3055,N_2825,N_2806);
xor U3056 (N_3056,N_2830,N_2885);
nor U3057 (N_3057,N_2876,N_2895);
xnor U3058 (N_3058,N_2902,N_2839);
and U3059 (N_3059,N_2827,N_2959);
and U3060 (N_3060,N_2961,N_2975);
or U3061 (N_3061,N_2956,N_2985);
nand U3062 (N_3062,N_2979,N_2873);
xnor U3063 (N_3063,N_2955,N_2884);
xnor U3064 (N_3064,N_2921,N_2929);
nor U3065 (N_3065,N_2965,N_2988);
and U3066 (N_3066,N_2886,N_2894);
and U3067 (N_3067,N_2971,N_2843);
and U3068 (N_3068,N_2945,N_2946);
nor U3069 (N_3069,N_2907,N_2941);
nor U3070 (N_3070,N_2887,N_2992);
or U3071 (N_3071,N_2848,N_2892);
xor U3072 (N_3072,N_2801,N_2842);
nand U3073 (N_3073,N_2829,N_2905);
xor U3074 (N_3074,N_2891,N_2807);
nor U3075 (N_3075,N_2818,N_2967);
or U3076 (N_3076,N_2912,N_2838);
or U3077 (N_3077,N_2861,N_2851);
and U3078 (N_3078,N_2814,N_2811);
nand U3079 (N_3079,N_2855,N_2943);
nor U3080 (N_3080,N_2960,N_2849);
nand U3081 (N_3081,N_2963,N_2981);
nor U3082 (N_3082,N_2833,N_2868);
and U3083 (N_3083,N_2888,N_2853);
xnor U3084 (N_3084,N_2805,N_2911);
nand U3085 (N_3085,N_2950,N_2889);
nand U3086 (N_3086,N_2856,N_2854);
and U3087 (N_3087,N_2803,N_2871);
nor U3088 (N_3088,N_2978,N_2819);
or U3089 (N_3089,N_2919,N_2940);
nor U3090 (N_3090,N_2900,N_2883);
xor U3091 (N_3091,N_2933,N_2920);
and U3092 (N_3092,N_2991,N_2937);
nor U3093 (N_3093,N_2867,N_2925);
or U3094 (N_3094,N_2998,N_2835);
and U3095 (N_3095,N_2995,N_2862);
nor U3096 (N_3096,N_2947,N_2817);
or U3097 (N_3097,N_2989,N_2962);
nor U3098 (N_3098,N_2915,N_2901);
or U3099 (N_3099,N_2927,N_2930);
and U3100 (N_3100,N_2957,N_2820);
xor U3101 (N_3101,N_2823,N_2832);
or U3102 (N_3102,N_2992,N_2925);
or U3103 (N_3103,N_2902,N_2972);
or U3104 (N_3104,N_2804,N_2806);
or U3105 (N_3105,N_2899,N_2986);
or U3106 (N_3106,N_2872,N_2905);
nor U3107 (N_3107,N_2992,N_2838);
nand U3108 (N_3108,N_2931,N_2800);
nor U3109 (N_3109,N_2929,N_2963);
nand U3110 (N_3110,N_2911,N_2904);
or U3111 (N_3111,N_2909,N_2818);
nand U3112 (N_3112,N_2887,N_2927);
and U3113 (N_3113,N_2911,N_2890);
xor U3114 (N_3114,N_2913,N_2895);
nand U3115 (N_3115,N_2815,N_2869);
or U3116 (N_3116,N_2867,N_2885);
and U3117 (N_3117,N_2830,N_2981);
nand U3118 (N_3118,N_2851,N_2859);
and U3119 (N_3119,N_2891,N_2935);
nand U3120 (N_3120,N_2969,N_2948);
and U3121 (N_3121,N_2944,N_2938);
nor U3122 (N_3122,N_2986,N_2924);
and U3123 (N_3123,N_2887,N_2942);
nand U3124 (N_3124,N_2801,N_2802);
xor U3125 (N_3125,N_2955,N_2802);
nor U3126 (N_3126,N_2930,N_2874);
and U3127 (N_3127,N_2855,N_2863);
and U3128 (N_3128,N_2999,N_2938);
xnor U3129 (N_3129,N_2841,N_2920);
or U3130 (N_3130,N_2807,N_2854);
or U3131 (N_3131,N_2844,N_2934);
nor U3132 (N_3132,N_2829,N_2926);
or U3133 (N_3133,N_2843,N_2927);
or U3134 (N_3134,N_2852,N_2858);
nand U3135 (N_3135,N_2909,N_2923);
nand U3136 (N_3136,N_2863,N_2982);
nand U3137 (N_3137,N_2956,N_2856);
nand U3138 (N_3138,N_2953,N_2811);
nand U3139 (N_3139,N_2900,N_2872);
nand U3140 (N_3140,N_2855,N_2894);
nor U3141 (N_3141,N_2909,N_2881);
xnor U3142 (N_3142,N_2915,N_2976);
and U3143 (N_3143,N_2895,N_2869);
nor U3144 (N_3144,N_2806,N_2955);
xnor U3145 (N_3145,N_2822,N_2891);
xor U3146 (N_3146,N_2820,N_2939);
and U3147 (N_3147,N_2843,N_2860);
nor U3148 (N_3148,N_2802,N_2911);
nor U3149 (N_3149,N_2827,N_2908);
nand U3150 (N_3150,N_2857,N_2880);
nand U3151 (N_3151,N_2984,N_2938);
nand U3152 (N_3152,N_2830,N_2868);
xor U3153 (N_3153,N_2818,N_2941);
xor U3154 (N_3154,N_2968,N_2935);
or U3155 (N_3155,N_2857,N_2847);
and U3156 (N_3156,N_2808,N_2820);
and U3157 (N_3157,N_2820,N_2834);
nor U3158 (N_3158,N_2867,N_2849);
nand U3159 (N_3159,N_2998,N_2975);
nand U3160 (N_3160,N_2868,N_2892);
xnor U3161 (N_3161,N_2864,N_2868);
and U3162 (N_3162,N_2960,N_2861);
xor U3163 (N_3163,N_2819,N_2882);
or U3164 (N_3164,N_2825,N_2901);
or U3165 (N_3165,N_2844,N_2821);
nor U3166 (N_3166,N_2821,N_2985);
xor U3167 (N_3167,N_2928,N_2972);
and U3168 (N_3168,N_2835,N_2885);
nor U3169 (N_3169,N_2941,N_2870);
xnor U3170 (N_3170,N_2923,N_2865);
nor U3171 (N_3171,N_2832,N_2830);
nand U3172 (N_3172,N_2970,N_2920);
xor U3173 (N_3173,N_2840,N_2989);
nand U3174 (N_3174,N_2919,N_2921);
nand U3175 (N_3175,N_2880,N_2940);
or U3176 (N_3176,N_2988,N_2969);
or U3177 (N_3177,N_2805,N_2980);
nand U3178 (N_3178,N_2922,N_2889);
nand U3179 (N_3179,N_2825,N_2838);
xor U3180 (N_3180,N_2956,N_2839);
and U3181 (N_3181,N_2936,N_2955);
xnor U3182 (N_3182,N_2877,N_2970);
and U3183 (N_3183,N_2804,N_2961);
or U3184 (N_3184,N_2861,N_2963);
nand U3185 (N_3185,N_2921,N_2823);
nor U3186 (N_3186,N_2908,N_2853);
or U3187 (N_3187,N_2878,N_2968);
nand U3188 (N_3188,N_2819,N_2909);
nor U3189 (N_3189,N_2862,N_2842);
and U3190 (N_3190,N_2965,N_2818);
and U3191 (N_3191,N_2871,N_2899);
nor U3192 (N_3192,N_2898,N_2808);
nor U3193 (N_3193,N_2811,N_2936);
nand U3194 (N_3194,N_2941,N_2944);
nor U3195 (N_3195,N_2905,N_2885);
nand U3196 (N_3196,N_2820,N_2962);
and U3197 (N_3197,N_2964,N_2811);
xor U3198 (N_3198,N_2859,N_2944);
or U3199 (N_3199,N_2905,N_2943);
nand U3200 (N_3200,N_3079,N_3164);
xor U3201 (N_3201,N_3047,N_3126);
or U3202 (N_3202,N_3076,N_3194);
nand U3203 (N_3203,N_3121,N_3022);
nor U3204 (N_3204,N_3173,N_3197);
xnor U3205 (N_3205,N_3091,N_3003);
or U3206 (N_3206,N_3016,N_3025);
nor U3207 (N_3207,N_3137,N_3188);
nand U3208 (N_3208,N_3104,N_3138);
or U3209 (N_3209,N_3096,N_3002);
or U3210 (N_3210,N_3008,N_3048);
nand U3211 (N_3211,N_3199,N_3108);
and U3212 (N_3212,N_3097,N_3136);
xor U3213 (N_3213,N_3129,N_3087);
and U3214 (N_3214,N_3105,N_3195);
and U3215 (N_3215,N_3169,N_3049);
or U3216 (N_3216,N_3056,N_3058);
and U3217 (N_3217,N_3122,N_3174);
nand U3218 (N_3218,N_3118,N_3168);
or U3219 (N_3219,N_3123,N_3027);
xnor U3220 (N_3220,N_3190,N_3083);
or U3221 (N_3221,N_3167,N_3141);
xor U3222 (N_3222,N_3117,N_3158);
xnor U3223 (N_3223,N_3040,N_3115);
nor U3224 (N_3224,N_3162,N_3031);
and U3225 (N_3225,N_3156,N_3110);
nor U3226 (N_3226,N_3088,N_3112);
nand U3227 (N_3227,N_3014,N_3103);
or U3228 (N_3228,N_3139,N_3042);
nor U3229 (N_3229,N_3045,N_3033);
nor U3230 (N_3230,N_3142,N_3067);
or U3231 (N_3231,N_3095,N_3052);
nor U3232 (N_3232,N_3070,N_3114);
and U3233 (N_3233,N_3061,N_3145);
and U3234 (N_3234,N_3119,N_3099);
xnor U3235 (N_3235,N_3054,N_3039);
or U3236 (N_3236,N_3128,N_3152);
and U3237 (N_3237,N_3144,N_3155);
or U3238 (N_3238,N_3055,N_3013);
and U3239 (N_3239,N_3113,N_3165);
or U3240 (N_3240,N_3077,N_3018);
xor U3241 (N_3241,N_3090,N_3157);
nor U3242 (N_3242,N_3127,N_3187);
nor U3243 (N_3243,N_3010,N_3130);
xnor U3244 (N_3244,N_3051,N_3044);
or U3245 (N_3245,N_3034,N_3150);
xnor U3246 (N_3246,N_3109,N_3050);
nor U3247 (N_3247,N_3030,N_3021);
or U3248 (N_3248,N_3098,N_3075);
xnor U3249 (N_3249,N_3053,N_3159);
xnor U3250 (N_3250,N_3106,N_3160);
and U3251 (N_3251,N_3180,N_3064);
and U3252 (N_3252,N_3071,N_3149);
and U3253 (N_3253,N_3192,N_3147);
and U3254 (N_3254,N_3132,N_3073);
nor U3255 (N_3255,N_3024,N_3085);
nand U3256 (N_3256,N_3072,N_3125);
nand U3257 (N_3257,N_3111,N_3193);
nor U3258 (N_3258,N_3038,N_3086);
nand U3259 (N_3259,N_3089,N_3166);
nor U3260 (N_3260,N_3029,N_3116);
xor U3261 (N_3261,N_3094,N_3170);
xnor U3262 (N_3262,N_3009,N_3175);
xor U3263 (N_3263,N_3059,N_3081);
or U3264 (N_3264,N_3163,N_3062);
xnor U3265 (N_3265,N_3133,N_3068);
nor U3266 (N_3266,N_3177,N_3146);
and U3267 (N_3267,N_3196,N_3186);
xnor U3268 (N_3268,N_3065,N_3134);
nand U3269 (N_3269,N_3074,N_3035);
and U3270 (N_3270,N_3102,N_3100);
and U3271 (N_3271,N_3006,N_3026);
and U3272 (N_3272,N_3148,N_3161);
nand U3273 (N_3273,N_3046,N_3176);
and U3274 (N_3274,N_3140,N_3041);
xnor U3275 (N_3275,N_3107,N_3066);
or U3276 (N_3276,N_3060,N_3028);
xnor U3277 (N_3277,N_3037,N_3171);
or U3278 (N_3278,N_3005,N_3154);
xnor U3279 (N_3279,N_3124,N_3063);
nor U3280 (N_3280,N_3172,N_3143);
nor U3281 (N_3281,N_3120,N_3183);
xor U3282 (N_3282,N_3185,N_3001);
or U3283 (N_3283,N_3007,N_3084);
nor U3284 (N_3284,N_3182,N_3135);
xor U3285 (N_3285,N_3178,N_3080);
or U3286 (N_3286,N_3153,N_3043);
nand U3287 (N_3287,N_3198,N_3151);
nand U3288 (N_3288,N_3093,N_3000);
or U3289 (N_3289,N_3020,N_3069);
xnor U3290 (N_3290,N_3092,N_3019);
nor U3291 (N_3291,N_3023,N_3011);
xor U3292 (N_3292,N_3082,N_3184);
xnor U3293 (N_3293,N_3057,N_3015);
or U3294 (N_3294,N_3078,N_3101);
and U3295 (N_3295,N_3181,N_3191);
nand U3296 (N_3296,N_3036,N_3131);
nand U3297 (N_3297,N_3189,N_3179);
nand U3298 (N_3298,N_3004,N_3012);
and U3299 (N_3299,N_3032,N_3017);
or U3300 (N_3300,N_3173,N_3049);
nor U3301 (N_3301,N_3000,N_3034);
and U3302 (N_3302,N_3012,N_3071);
and U3303 (N_3303,N_3047,N_3143);
or U3304 (N_3304,N_3076,N_3074);
or U3305 (N_3305,N_3058,N_3119);
nor U3306 (N_3306,N_3031,N_3009);
and U3307 (N_3307,N_3148,N_3124);
and U3308 (N_3308,N_3019,N_3178);
nand U3309 (N_3309,N_3136,N_3159);
and U3310 (N_3310,N_3155,N_3067);
and U3311 (N_3311,N_3039,N_3010);
nor U3312 (N_3312,N_3094,N_3063);
xnor U3313 (N_3313,N_3079,N_3193);
xnor U3314 (N_3314,N_3126,N_3027);
and U3315 (N_3315,N_3031,N_3137);
or U3316 (N_3316,N_3164,N_3034);
and U3317 (N_3317,N_3090,N_3113);
or U3318 (N_3318,N_3003,N_3026);
and U3319 (N_3319,N_3001,N_3060);
nand U3320 (N_3320,N_3134,N_3138);
and U3321 (N_3321,N_3086,N_3070);
nand U3322 (N_3322,N_3150,N_3141);
nand U3323 (N_3323,N_3158,N_3012);
nor U3324 (N_3324,N_3092,N_3051);
xor U3325 (N_3325,N_3011,N_3041);
xnor U3326 (N_3326,N_3107,N_3067);
xor U3327 (N_3327,N_3004,N_3013);
xnor U3328 (N_3328,N_3161,N_3030);
nor U3329 (N_3329,N_3022,N_3089);
xor U3330 (N_3330,N_3110,N_3048);
nor U3331 (N_3331,N_3170,N_3120);
nand U3332 (N_3332,N_3177,N_3073);
nand U3333 (N_3333,N_3061,N_3196);
or U3334 (N_3334,N_3156,N_3137);
nor U3335 (N_3335,N_3022,N_3069);
or U3336 (N_3336,N_3055,N_3125);
or U3337 (N_3337,N_3171,N_3001);
nor U3338 (N_3338,N_3073,N_3117);
and U3339 (N_3339,N_3080,N_3098);
xor U3340 (N_3340,N_3005,N_3086);
or U3341 (N_3341,N_3159,N_3111);
nor U3342 (N_3342,N_3135,N_3153);
nor U3343 (N_3343,N_3193,N_3042);
nor U3344 (N_3344,N_3135,N_3009);
and U3345 (N_3345,N_3107,N_3148);
nor U3346 (N_3346,N_3127,N_3177);
xor U3347 (N_3347,N_3185,N_3140);
nand U3348 (N_3348,N_3066,N_3047);
nand U3349 (N_3349,N_3040,N_3193);
and U3350 (N_3350,N_3043,N_3045);
or U3351 (N_3351,N_3087,N_3194);
xnor U3352 (N_3352,N_3142,N_3131);
nor U3353 (N_3353,N_3045,N_3001);
nand U3354 (N_3354,N_3093,N_3004);
nor U3355 (N_3355,N_3011,N_3121);
or U3356 (N_3356,N_3173,N_3115);
or U3357 (N_3357,N_3142,N_3112);
xnor U3358 (N_3358,N_3105,N_3193);
nand U3359 (N_3359,N_3090,N_3122);
and U3360 (N_3360,N_3043,N_3187);
and U3361 (N_3361,N_3086,N_3065);
nand U3362 (N_3362,N_3125,N_3150);
and U3363 (N_3363,N_3149,N_3130);
and U3364 (N_3364,N_3096,N_3121);
xnor U3365 (N_3365,N_3184,N_3194);
and U3366 (N_3366,N_3092,N_3034);
nor U3367 (N_3367,N_3154,N_3042);
nor U3368 (N_3368,N_3185,N_3132);
and U3369 (N_3369,N_3021,N_3069);
nand U3370 (N_3370,N_3010,N_3015);
nor U3371 (N_3371,N_3135,N_3001);
nor U3372 (N_3372,N_3092,N_3157);
xnor U3373 (N_3373,N_3042,N_3172);
or U3374 (N_3374,N_3158,N_3179);
or U3375 (N_3375,N_3182,N_3067);
xnor U3376 (N_3376,N_3050,N_3160);
nor U3377 (N_3377,N_3075,N_3135);
xor U3378 (N_3378,N_3104,N_3111);
and U3379 (N_3379,N_3001,N_3137);
nor U3380 (N_3380,N_3137,N_3116);
xor U3381 (N_3381,N_3160,N_3023);
or U3382 (N_3382,N_3108,N_3112);
nor U3383 (N_3383,N_3152,N_3018);
and U3384 (N_3384,N_3140,N_3023);
and U3385 (N_3385,N_3043,N_3154);
and U3386 (N_3386,N_3001,N_3092);
nor U3387 (N_3387,N_3080,N_3029);
nand U3388 (N_3388,N_3126,N_3141);
xor U3389 (N_3389,N_3120,N_3002);
nor U3390 (N_3390,N_3121,N_3137);
and U3391 (N_3391,N_3010,N_3083);
xnor U3392 (N_3392,N_3084,N_3161);
nand U3393 (N_3393,N_3103,N_3118);
or U3394 (N_3394,N_3011,N_3125);
nand U3395 (N_3395,N_3122,N_3191);
nand U3396 (N_3396,N_3063,N_3162);
xor U3397 (N_3397,N_3066,N_3078);
or U3398 (N_3398,N_3027,N_3168);
xor U3399 (N_3399,N_3043,N_3074);
xor U3400 (N_3400,N_3313,N_3272);
and U3401 (N_3401,N_3309,N_3293);
nor U3402 (N_3402,N_3326,N_3227);
nor U3403 (N_3403,N_3241,N_3344);
nand U3404 (N_3404,N_3219,N_3332);
nand U3405 (N_3405,N_3233,N_3331);
xor U3406 (N_3406,N_3297,N_3248);
or U3407 (N_3407,N_3240,N_3260);
nand U3408 (N_3408,N_3236,N_3340);
nand U3409 (N_3409,N_3282,N_3257);
nor U3410 (N_3410,N_3203,N_3205);
or U3411 (N_3411,N_3350,N_3376);
nor U3412 (N_3412,N_3342,N_3371);
and U3413 (N_3413,N_3390,N_3379);
nor U3414 (N_3414,N_3298,N_3360);
and U3415 (N_3415,N_3374,N_3206);
nand U3416 (N_3416,N_3354,N_3396);
or U3417 (N_3417,N_3264,N_3391);
nor U3418 (N_3418,N_3259,N_3255);
or U3419 (N_3419,N_3222,N_3202);
xor U3420 (N_3420,N_3372,N_3336);
or U3421 (N_3421,N_3339,N_3279);
nand U3422 (N_3422,N_3212,N_3221);
xnor U3423 (N_3423,N_3277,N_3315);
and U3424 (N_3424,N_3238,N_3213);
nor U3425 (N_3425,N_3303,N_3305);
or U3426 (N_3426,N_3254,N_3366);
nor U3427 (N_3427,N_3209,N_3242);
nor U3428 (N_3428,N_3226,N_3249);
xor U3429 (N_3429,N_3263,N_3224);
or U3430 (N_3430,N_3311,N_3239);
and U3431 (N_3431,N_3268,N_3245);
or U3432 (N_3432,N_3351,N_3211);
nor U3433 (N_3433,N_3365,N_3208);
and U3434 (N_3434,N_3377,N_3285);
or U3435 (N_3435,N_3341,N_3327);
and U3436 (N_3436,N_3333,N_3355);
nand U3437 (N_3437,N_3352,N_3356);
nand U3438 (N_3438,N_3246,N_3232);
nor U3439 (N_3439,N_3393,N_3345);
nand U3440 (N_3440,N_3381,N_3296);
or U3441 (N_3441,N_3317,N_3325);
xor U3442 (N_3442,N_3383,N_3316);
nand U3443 (N_3443,N_3370,N_3382);
and U3444 (N_3444,N_3273,N_3385);
or U3445 (N_3445,N_3284,N_3278);
nand U3446 (N_3446,N_3395,N_3281);
or U3447 (N_3447,N_3274,N_3329);
or U3448 (N_3448,N_3337,N_3247);
nor U3449 (N_3449,N_3266,N_3312);
nor U3450 (N_3450,N_3225,N_3358);
nand U3451 (N_3451,N_3369,N_3320);
nor U3452 (N_3452,N_3322,N_3357);
xor U3453 (N_3453,N_3392,N_3301);
nor U3454 (N_3454,N_3330,N_3307);
and U3455 (N_3455,N_3368,N_3201);
or U3456 (N_3456,N_3314,N_3394);
nand U3457 (N_3457,N_3228,N_3335);
or U3458 (N_3458,N_3270,N_3286);
or U3459 (N_3459,N_3220,N_3265);
nor U3460 (N_3460,N_3218,N_3223);
nand U3461 (N_3461,N_3306,N_3308);
and U3462 (N_3462,N_3328,N_3399);
nand U3463 (N_3463,N_3364,N_3234);
xor U3464 (N_3464,N_3321,N_3304);
xnor U3465 (N_3465,N_3200,N_3210);
nor U3466 (N_3466,N_3388,N_3275);
nor U3467 (N_3467,N_3300,N_3291);
or U3468 (N_3468,N_3318,N_3346);
nor U3469 (N_3469,N_3384,N_3231);
and U3470 (N_3470,N_3290,N_3253);
or U3471 (N_3471,N_3230,N_3204);
nor U3472 (N_3472,N_3386,N_3269);
and U3473 (N_3473,N_3271,N_3295);
nand U3474 (N_3474,N_3243,N_3324);
xor U3475 (N_3475,N_3319,N_3363);
xnor U3476 (N_3476,N_3348,N_3310);
or U3477 (N_3477,N_3256,N_3338);
nor U3478 (N_3478,N_3375,N_3323);
nor U3479 (N_3479,N_3216,N_3289);
or U3480 (N_3480,N_3299,N_3294);
or U3481 (N_3481,N_3214,N_3261);
and U3482 (N_3482,N_3349,N_3217);
or U3483 (N_3483,N_3237,N_3267);
or U3484 (N_3484,N_3258,N_3359);
and U3485 (N_3485,N_3215,N_3250);
nor U3486 (N_3486,N_3343,N_3398);
and U3487 (N_3487,N_3207,N_3276);
or U3488 (N_3488,N_3347,N_3292);
and U3489 (N_3489,N_3389,N_3244);
xnor U3490 (N_3490,N_3235,N_3378);
or U3491 (N_3491,N_3361,N_3353);
nor U3492 (N_3492,N_3280,N_3287);
and U3493 (N_3493,N_3251,N_3334);
or U3494 (N_3494,N_3302,N_3397);
or U3495 (N_3495,N_3283,N_3288);
nor U3496 (N_3496,N_3367,N_3252);
nand U3497 (N_3497,N_3362,N_3380);
nor U3498 (N_3498,N_3229,N_3387);
or U3499 (N_3499,N_3262,N_3373);
nor U3500 (N_3500,N_3285,N_3286);
or U3501 (N_3501,N_3340,N_3394);
nor U3502 (N_3502,N_3367,N_3284);
nand U3503 (N_3503,N_3323,N_3340);
xnor U3504 (N_3504,N_3389,N_3207);
and U3505 (N_3505,N_3259,N_3289);
nor U3506 (N_3506,N_3365,N_3331);
nor U3507 (N_3507,N_3252,N_3270);
or U3508 (N_3508,N_3323,N_3302);
and U3509 (N_3509,N_3248,N_3222);
xnor U3510 (N_3510,N_3292,N_3355);
and U3511 (N_3511,N_3382,N_3302);
nand U3512 (N_3512,N_3363,N_3324);
or U3513 (N_3513,N_3379,N_3279);
nor U3514 (N_3514,N_3296,N_3315);
nand U3515 (N_3515,N_3317,N_3388);
nand U3516 (N_3516,N_3200,N_3296);
or U3517 (N_3517,N_3217,N_3290);
and U3518 (N_3518,N_3388,N_3304);
nand U3519 (N_3519,N_3271,N_3392);
and U3520 (N_3520,N_3286,N_3362);
nor U3521 (N_3521,N_3207,N_3331);
and U3522 (N_3522,N_3365,N_3350);
and U3523 (N_3523,N_3288,N_3350);
and U3524 (N_3524,N_3370,N_3201);
and U3525 (N_3525,N_3388,N_3248);
and U3526 (N_3526,N_3201,N_3306);
nor U3527 (N_3527,N_3227,N_3294);
and U3528 (N_3528,N_3317,N_3253);
nand U3529 (N_3529,N_3362,N_3282);
xnor U3530 (N_3530,N_3314,N_3250);
nor U3531 (N_3531,N_3382,N_3322);
xnor U3532 (N_3532,N_3282,N_3234);
or U3533 (N_3533,N_3323,N_3284);
nand U3534 (N_3534,N_3373,N_3249);
nand U3535 (N_3535,N_3330,N_3264);
nand U3536 (N_3536,N_3219,N_3255);
nor U3537 (N_3537,N_3244,N_3248);
or U3538 (N_3538,N_3227,N_3264);
xor U3539 (N_3539,N_3283,N_3271);
xnor U3540 (N_3540,N_3223,N_3253);
nor U3541 (N_3541,N_3296,N_3394);
or U3542 (N_3542,N_3315,N_3224);
nor U3543 (N_3543,N_3360,N_3307);
nor U3544 (N_3544,N_3350,N_3374);
and U3545 (N_3545,N_3214,N_3333);
and U3546 (N_3546,N_3260,N_3381);
nand U3547 (N_3547,N_3224,N_3330);
xnor U3548 (N_3548,N_3328,N_3335);
nor U3549 (N_3549,N_3276,N_3361);
and U3550 (N_3550,N_3362,N_3395);
nor U3551 (N_3551,N_3361,N_3251);
nor U3552 (N_3552,N_3241,N_3291);
xnor U3553 (N_3553,N_3320,N_3365);
nand U3554 (N_3554,N_3396,N_3258);
and U3555 (N_3555,N_3386,N_3271);
nand U3556 (N_3556,N_3210,N_3260);
and U3557 (N_3557,N_3229,N_3364);
and U3558 (N_3558,N_3273,N_3258);
xor U3559 (N_3559,N_3251,N_3256);
nand U3560 (N_3560,N_3237,N_3253);
xnor U3561 (N_3561,N_3262,N_3235);
and U3562 (N_3562,N_3307,N_3354);
nor U3563 (N_3563,N_3210,N_3304);
and U3564 (N_3564,N_3208,N_3314);
nand U3565 (N_3565,N_3264,N_3327);
and U3566 (N_3566,N_3232,N_3200);
and U3567 (N_3567,N_3289,N_3382);
nor U3568 (N_3568,N_3317,N_3201);
nand U3569 (N_3569,N_3350,N_3394);
and U3570 (N_3570,N_3214,N_3240);
nand U3571 (N_3571,N_3375,N_3359);
xor U3572 (N_3572,N_3388,N_3338);
and U3573 (N_3573,N_3361,N_3227);
nand U3574 (N_3574,N_3334,N_3293);
or U3575 (N_3575,N_3272,N_3323);
nand U3576 (N_3576,N_3371,N_3290);
or U3577 (N_3577,N_3387,N_3236);
xnor U3578 (N_3578,N_3211,N_3229);
nor U3579 (N_3579,N_3394,N_3343);
xor U3580 (N_3580,N_3230,N_3210);
nor U3581 (N_3581,N_3239,N_3204);
and U3582 (N_3582,N_3288,N_3257);
xor U3583 (N_3583,N_3249,N_3316);
xnor U3584 (N_3584,N_3227,N_3248);
nor U3585 (N_3585,N_3316,N_3289);
nand U3586 (N_3586,N_3297,N_3279);
or U3587 (N_3587,N_3296,N_3253);
xor U3588 (N_3588,N_3342,N_3274);
xnor U3589 (N_3589,N_3219,N_3260);
or U3590 (N_3590,N_3222,N_3399);
or U3591 (N_3591,N_3214,N_3234);
xor U3592 (N_3592,N_3248,N_3394);
and U3593 (N_3593,N_3276,N_3349);
xor U3594 (N_3594,N_3283,N_3394);
and U3595 (N_3595,N_3297,N_3385);
or U3596 (N_3596,N_3236,N_3214);
and U3597 (N_3597,N_3270,N_3266);
or U3598 (N_3598,N_3303,N_3293);
and U3599 (N_3599,N_3221,N_3390);
nand U3600 (N_3600,N_3465,N_3566);
nor U3601 (N_3601,N_3445,N_3533);
nor U3602 (N_3602,N_3451,N_3573);
nand U3603 (N_3603,N_3499,N_3491);
nor U3604 (N_3604,N_3590,N_3525);
nor U3605 (N_3605,N_3421,N_3441);
xnor U3606 (N_3606,N_3449,N_3487);
and U3607 (N_3607,N_3505,N_3534);
nor U3608 (N_3608,N_3442,N_3584);
or U3609 (N_3609,N_3524,N_3575);
xnor U3610 (N_3610,N_3532,N_3531);
nor U3611 (N_3611,N_3474,N_3446);
and U3612 (N_3612,N_3429,N_3548);
nand U3613 (N_3613,N_3581,N_3588);
and U3614 (N_3614,N_3472,N_3425);
nor U3615 (N_3615,N_3527,N_3593);
nor U3616 (N_3616,N_3556,N_3520);
nor U3617 (N_3617,N_3550,N_3485);
or U3618 (N_3618,N_3591,N_3511);
nor U3619 (N_3619,N_3435,N_3479);
nor U3620 (N_3620,N_3483,N_3502);
or U3621 (N_3621,N_3419,N_3408);
nand U3622 (N_3622,N_3553,N_3519);
xor U3623 (N_3623,N_3493,N_3565);
and U3624 (N_3624,N_3571,N_3506);
nand U3625 (N_3625,N_3536,N_3557);
nor U3626 (N_3626,N_3495,N_3458);
nor U3627 (N_3627,N_3438,N_3475);
or U3628 (N_3628,N_3522,N_3407);
and U3629 (N_3629,N_3488,N_3521);
nor U3630 (N_3630,N_3587,N_3547);
nand U3631 (N_3631,N_3523,N_3517);
xor U3632 (N_3632,N_3572,N_3529);
nand U3633 (N_3633,N_3447,N_3436);
and U3634 (N_3634,N_3585,N_3539);
nand U3635 (N_3635,N_3486,N_3471);
or U3636 (N_3636,N_3466,N_3481);
or U3637 (N_3637,N_3530,N_3559);
or U3638 (N_3638,N_3583,N_3461);
and U3639 (N_3639,N_3510,N_3450);
or U3640 (N_3640,N_3443,N_3545);
or U3641 (N_3641,N_3453,N_3542);
nor U3642 (N_3642,N_3592,N_3574);
nand U3643 (N_3643,N_3457,N_3526);
and U3644 (N_3644,N_3404,N_3482);
xor U3645 (N_3645,N_3433,N_3444);
or U3646 (N_3646,N_3589,N_3409);
nor U3647 (N_3647,N_3416,N_3504);
xnor U3648 (N_3648,N_3538,N_3518);
or U3649 (N_3649,N_3470,N_3423);
and U3650 (N_3650,N_3498,N_3422);
and U3651 (N_3651,N_3403,N_3512);
or U3652 (N_3652,N_3464,N_3546);
and U3653 (N_3653,N_3417,N_3568);
or U3654 (N_3654,N_3497,N_3543);
xnor U3655 (N_3655,N_3544,N_3406);
nor U3656 (N_3656,N_3469,N_3463);
nor U3657 (N_3657,N_3509,N_3560);
nor U3658 (N_3658,N_3494,N_3595);
and U3659 (N_3659,N_3582,N_3480);
nand U3660 (N_3660,N_3428,N_3551);
xor U3661 (N_3661,N_3555,N_3478);
nand U3662 (N_3662,N_3549,N_3562);
nand U3663 (N_3663,N_3439,N_3578);
xnor U3664 (N_3664,N_3516,N_3434);
xnor U3665 (N_3665,N_3496,N_3460);
or U3666 (N_3666,N_3500,N_3596);
xor U3667 (N_3667,N_3411,N_3456);
nor U3668 (N_3668,N_3431,N_3427);
xnor U3669 (N_3669,N_3569,N_3405);
or U3670 (N_3670,N_3537,N_3437);
nand U3671 (N_3671,N_3594,N_3489);
or U3672 (N_3672,N_3432,N_3528);
and U3673 (N_3673,N_3467,N_3426);
or U3674 (N_3674,N_3490,N_3541);
nor U3675 (N_3675,N_3476,N_3412);
or U3676 (N_3676,N_3473,N_3402);
nor U3677 (N_3677,N_3418,N_3597);
nor U3678 (N_3678,N_3579,N_3576);
and U3679 (N_3679,N_3535,N_3501);
and U3680 (N_3680,N_3503,N_3508);
nor U3681 (N_3681,N_3477,N_3558);
or U3682 (N_3682,N_3599,N_3415);
and U3683 (N_3683,N_3484,N_3580);
xor U3684 (N_3684,N_3414,N_3507);
or U3685 (N_3685,N_3564,N_3413);
xor U3686 (N_3686,N_3452,N_3459);
nor U3687 (N_3687,N_3492,N_3577);
nor U3688 (N_3688,N_3561,N_3563);
xor U3689 (N_3689,N_3514,N_3430);
and U3690 (N_3690,N_3420,N_3552);
or U3691 (N_3691,N_3424,N_3570);
nor U3692 (N_3692,N_3468,N_3586);
or U3693 (N_3693,N_3515,N_3448);
xnor U3694 (N_3694,N_3454,N_3540);
xor U3695 (N_3695,N_3554,N_3598);
xnor U3696 (N_3696,N_3410,N_3513);
nor U3697 (N_3697,N_3400,N_3440);
or U3698 (N_3698,N_3455,N_3462);
xnor U3699 (N_3699,N_3401,N_3567);
nor U3700 (N_3700,N_3590,N_3500);
nand U3701 (N_3701,N_3482,N_3490);
and U3702 (N_3702,N_3535,N_3516);
and U3703 (N_3703,N_3494,N_3506);
nand U3704 (N_3704,N_3409,N_3449);
and U3705 (N_3705,N_3574,N_3430);
and U3706 (N_3706,N_3558,N_3545);
and U3707 (N_3707,N_3479,N_3518);
xnor U3708 (N_3708,N_3434,N_3491);
nand U3709 (N_3709,N_3417,N_3411);
xor U3710 (N_3710,N_3420,N_3469);
or U3711 (N_3711,N_3405,N_3417);
or U3712 (N_3712,N_3572,N_3462);
nor U3713 (N_3713,N_3582,N_3484);
and U3714 (N_3714,N_3553,N_3501);
or U3715 (N_3715,N_3485,N_3446);
or U3716 (N_3716,N_3581,N_3548);
nand U3717 (N_3717,N_3586,N_3587);
nand U3718 (N_3718,N_3517,N_3471);
xnor U3719 (N_3719,N_3459,N_3494);
nand U3720 (N_3720,N_3598,N_3546);
or U3721 (N_3721,N_3484,N_3449);
and U3722 (N_3722,N_3448,N_3409);
or U3723 (N_3723,N_3517,N_3582);
xnor U3724 (N_3724,N_3482,N_3451);
and U3725 (N_3725,N_3427,N_3433);
or U3726 (N_3726,N_3466,N_3509);
and U3727 (N_3727,N_3474,N_3432);
or U3728 (N_3728,N_3579,N_3585);
and U3729 (N_3729,N_3527,N_3447);
and U3730 (N_3730,N_3481,N_3470);
and U3731 (N_3731,N_3566,N_3411);
or U3732 (N_3732,N_3478,N_3461);
or U3733 (N_3733,N_3412,N_3491);
nor U3734 (N_3734,N_3574,N_3426);
and U3735 (N_3735,N_3500,N_3424);
or U3736 (N_3736,N_3599,N_3460);
xnor U3737 (N_3737,N_3483,N_3524);
nor U3738 (N_3738,N_3582,N_3549);
xnor U3739 (N_3739,N_3559,N_3550);
xnor U3740 (N_3740,N_3453,N_3478);
nor U3741 (N_3741,N_3477,N_3468);
nand U3742 (N_3742,N_3447,N_3442);
nor U3743 (N_3743,N_3583,N_3430);
or U3744 (N_3744,N_3449,N_3550);
nand U3745 (N_3745,N_3537,N_3534);
and U3746 (N_3746,N_3447,N_3511);
xor U3747 (N_3747,N_3586,N_3454);
xor U3748 (N_3748,N_3496,N_3400);
nor U3749 (N_3749,N_3513,N_3534);
xnor U3750 (N_3750,N_3544,N_3549);
and U3751 (N_3751,N_3546,N_3453);
nor U3752 (N_3752,N_3577,N_3597);
nor U3753 (N_3753,N_3576,N_3584);
nor U3754 (N_3754,N_3503,N_3494);
nand U3755 (N_3755,N_3533,N_3588);
and U3756 (N_3756,N_3548,N_3457);
nand U3757 (N_3757,N_3511,N_3405);
nor U3758 (N_3758,N_3574,N_3538);
xnor U3759 (N_3759,N_3525,N_3479);
or U3760 (N_3760,N_3427,N_3472);
nor U3761 (N_3761,N_3597,N_3462);
nor U3762 (N_3762,N_3432,N_3548);
and U3763 (N_3763,N_3429,N_3501);
nor U3764 (N_3764,N_3462,N_3496);
and U3765 (N_3765,N_3563,N_3582);
xor U3766 (N_3766,N_3551,N_3521);
xor U3767 (N_3767,N_3402,N_3589);
nor U3768 (N_3768,N_3427,N_3492);
nor U3769 (N_3769,N_3422,N_3470);
or U3770 (N_3770,N_3500,N_3458);
xor U3771 (N_3771,N_3405,N_3582);
and U3772 (N_3772,N_3462,N_3431);
nand U3773 (N_3773,N_3514,N_3495);
xnor U3774 (N_3774,N_3594,N_3549);
xnor U3775 (N_3775,N_3498,N_3597);
nor U3776 (N_3776,N_3432,N_3571);
nor U3777 (N_3777,N_3407,N_3405);
nand U3778 (N_3778,N_3584,N_3444);
or U3779 (N_3779,N_3403,N_3528);
nand U3780 (N_3780,N_3555,N_3468);
xor U3781 (N_3781,N_3560,N_3558);
nand U3782 (N_3782,N_3418,N_3529);
nor U3783 (N_3783,N_3596,N_3497);
nand U3784 (N_3784,N_3554,N_3470);
xor U3785 (N_3785,N_3413,N_3429);
and U3786 (N_3786,N_3463,N_3418);
or U3787 (N_3787,N_3576,N_3411);
or U3788 (N_3788,N_3464,N_3406);
nand U3789 (N_3789,N_3580,N_3491);
or U3790 (N_3790,N_3446,N_3492);
xor U3791 (N_3791,N_3421,N_3575);
nand U3792 (N_3792,N_3459,N_3427);
xor U3793 (N_3793,N_3545,N_3512);
or U3794 (N_3794,N_3541,N_3435);
nor U3795 (N_3795,N_3459,N_3455);
or U3796 (N_3796,N_3547,N_3447);
nor U3797 (N_3797,N_3477,N_3497);
or U3798 (N_3798,N_3467,N_3440);
and U3799 (N_3799,N_3495,N_3550);
xnor U3800 (N_3800,N_3616,N_3739);
or U3801 (N_3801,N_3696,N_3751);
or U3802 (N_3802,N_3767,N_3752);
nor U3803 (N_3803,N_3731,N_3613);
xnor U3804 (N_3804,N_3639,N_3723);
xnor U3805 (N_3805,N_3712,N_3735);
xnor U3806 (N_3806,N_3701,N_3738);
or U3807 (N_3807,N_3663,N_3710);
and U3808 (N_3808,N_3722,N_3730);
nand U3809 (N_3809,N_3636,N_3720);
nor U3810 (N_3810,N_3754,N_3689);
nor U3811 (N_3811,N_3706,N_3627);
nor U3812 (N_3812,N_3733,N_3654);
or U3813 (N_3813,N_3603,N_3615);
and U3814 (N_3814,N_3607,N_3625);
nand U3815 (N_3815,N_3676,N_3747);
xor U3816 (N_3816,N_3624,N_3734);
and U3817 (N_3817,N_3770,N_3737);
and U3818 (N_3818,N_3708,N_3668);
nor U3819 (N_3819,N_3766,N_3764);
nor U3820 (N_3820,N_3640,N_3635);
nand U3821 (N_3821,N_3776,N_3610);
nor U3822 (N_3822,N_3719,N_3728);
nor U3823 (N_3823,N_3688,N_3691);
xnor U3824 (N_3824,N_3662,N_3736);
or U3825 (N_3825,N_3619,N_3727);
and U3826 (N_3826,N_3634,N_3763);
xor U3827 (N_3827,N_3618,N_3681);
or U3828 (N_3828,N_3630,N_3661);
nor U3829 (N_3829,N_3711,N_3784);
nor U3830 (N_3830,N_3673,N_3664);
or U3831 (N_3831,N_3702,N_3601);
or U3832 (N_3832,N_3693,N_3667);
nor U3833 (N_3833,N_3651,N_3791);
and U3834 (N_3834,N_3638,N_3797);
xnor U3835 (N_3835,N_3602,N_3773);
or U3836 (N_3836,N_3718,N_3652);
xor U3837 (N_3837,N_3623,N_3709);
nor U3838 (N_3838,N_3778,N_3682);
nand U3839 (N_3839,N_3740,N_3671);
nor U3840 (N_3840,N_3721,N_3765);
xor U3841 (N_3841,N_3707,N_3694);
xor U3842 (N_3842,N_3724,N_3665);
nand U3843 (N_3843,N_3685,N_3798);
nor U3844 (N_3844,N_3622,N_3726);
or U3845 (N_3845,N_3666,N_3695);
xnor U3846 (N_3846,N_3632,N_3750);
nor U3847 (N_3847,N_3641,N_3692);
and U3848 (N_3848,N_3631,N_3612);
nor U3849 (N_3849,N_3748,N_3698);
nand U3850 (N_3850,N_3606,N_3741);
and U3851 (N_3851,N_3657,N_3787);
nor U3852 (N_3852,N_3658,N_3659);
nand U3853 (N_3853,N_3725,N_3617);
and U3854 (N_3854,N_3604,N_3672);
or U3855 (N_3855,N_3780,N_3793);
and U3856 (N_3856,N_3759,N_3690);
and U3857 (N_3857,N_3675,N_3753);
nand U3858 (N_3858,N_3680,N_3611);
and U3859 (N_3859,N_3628,N_3713);
nor U3860 (N_3860,N_3660,N_3755);
nand U3861 (N_3861,N_3796,N_3669);
or U3862 (N_3862,N_3732,N_3684);
or U3863 (N_3863,N_3783,N_3761);
or U3864 (N_3864,N_3647,N_3794);
or U3865 (N_3865,N_3746,N_3717);
or U3866 (N_3866,N_3792,N_3655);
xnor U3867 (N_3867,N_3789,N_3629);
nor U3868 (N_3868,N_3633,N_3642);
xnor U3869 (N_3869,N_3757,N_3756);
or U3870 (N_3870,N_3677,N_3714);
or U3871 (N_3871,N_3687,N_3790);
nand U3872 (N_3872,N_3645,N_3786);
xor U3873 (N_3873,N_3774,N_3729);
or U3874 (N_3874,N_3626,N_3775);
xor U3875 (N_3875,N_3777,N_3697);
or U3876 (N_3876,N_3614,N_3744);
or U3877 (N_3877,N_3795,N_3700);
nor U3878 (N_3878,N_3621,N_3768);
or U3879 (N_3879,N_3779,N_3760);
nor U3880 (N_3880,N_3743,N_3769);
or U3881 (N_3881,N_3745,N_3749);
xor U3882 (N_3882,N_3678,N_3653);
xnor U3883 (N_3883,N_3785,N_3704);
and U3884 (N_3884,N_3716,N_3799);
or U3885 (N_3885,N_3781,N_3646);
xor U3886 (N_3886,N_3643,N_3605);
or U3887 (N_3887,N_3762,N_3674);
nand U3888 (N_3888,N_3772,N_3705);
nand U3889 (N_3889,N_3683,N_3600);
or U3890 (N_3890,N_3608,N_3703);
and U3891 (N_3891,N_3649,N_3644);
nand U3892 (N_3892,N_3715,N_3782);
nand U3893 (N_3893,N_3771,N_3679);
or U3894 (N_3894,N_3686,N_3758);
xnor U3895 (N_3895,N_3742,N_3609);
and U3896 (N_3896,N_3637,N_3670);
and U3897 (N_3897,N_3620,N_3656);
nand U3898 (N_3898,N_3699,N_3788);
and U3899 (N_3899,N_3650,N_3648);
nand U3900 (N_3900,N_3751,N_3619);
xor U3901 (N_3901,N_3774,N_3611);
nor U3902 (N_3902,N_3796,N_3639);
nor U3903 (N_3903,N_3617,N_3631);
and U3904 (N_3904,N_3641,N_3675);
xor U3905 (N_3905,N_3752,N_3735);
xor U3906 (N_3906,N_3784,N_3700);
or U3907 (N_3907,N_3780,N_3712);
or U3908 (N_3908,N_3625,N_3699);
nand U3909 (N_3909,N_3612,N_3722);
xnor U3910 (N_3910,N_3761,N_3644);
xnor U3911 (N_3911,N_3634,N_3744);
nand U3912 (N_3912,N_3783,N_3768);
nor U3913 (N_3913,N_3674,N_3709);
and U3914 (N_3914,N_3765,N_3619);
and U3915 (N_3915,N_3772,N_3669);
and U3916 (N_3916,N_3628,N_3702);
and U3917 (N_3917,N_3614,N_3726);
xnor U3918 (N_3918,N_3730,N_3782);
nand U3919 (N_3919,N_3687,N_3703);
xor U3920 (N_3920,N_3709,N_3740);
xor U3921 (N_3921,N_3602,N_3657);
nor U3922 (N_3922,N_3703,N_3749);
or U3923 (N_3923,N_3608,N_3639);
xnor U3924 (N_3924,N_3793,N_3601);
and U3925 (N_3925,N_3712,N_3717);
and U3926 (N_3926,N_3786,N_3750);
xor U3927 (N_3927,N_3795,N_3657);
nor U3928 (N_3928,N_3688,N_3669);
nor U3929 (N_3929,N_3612,N_3718);
nor U3930 (N_3930,N_3743,N_3658);
and U3931 (N_3931,N_3606,N_3679);
nor U3932 (N_3932,N_3735,N_3767);
or U3933 (N_3933,N_3766,N_3688);
xor U3934 (N_3934,N_3796,N_3785);
nor U3935 (N_3935,N_3677,N_3710);
nor U3936 (N_3936,N_3643,N_3786);
or U3937 (N_3937,N_3695,N_3628);
nor U3938 (N_3938,N_3737,N_3714);
or U3939 (N_3939,N_3761,N_3779);
or U3940 (N_3940,N_3696,N_3613);
nor U3941 (N_3941,N_3745,N_3621);
nor U3942 (N_3942,N_3715,N_3779);
nor U3943 (N_3943,N_3695,N_3689);
xor U3944 (N_3944,N_3767,N_3641);
or U3945 (N_3945,N_3791,N_3638);
nor U3946 (N_3946,N_3699,N_3655);
and U3947 (N_3947,N_3764,N_3614);
xor U3948 (N_3948,N_3623,N_3710);
nand U3949 (N_3949,N_3677,N_3689);
xor U3950 (N_3950,N_3725,N_3731);
nand U3951 (N_3951,N_3750,N_3630);
nand U3952 (N_3952,N_3715,N_3641);
nand U3953 (N_3953,N_3686,N_3652);
nor U3954 (N_3954,N_3679,N_3668);
nor U3955 (N_3955,N_3759,N_3674);
nor U3956 (N_3956,N_3680,N_3775);
or U3957 (N_3957,N_3641,N_3644);
xnor U3958 (N_3958,N_3748,N_3694);
nand U3959 (N_3959,N_3736,N_3702);
and U3960 (N_3960,N_3604,N_3718);
or U3961 (N_3961,N_3686,N_3664);
nand U3962 (N_3962,N_3773,N_3761);
xnor U3963 (N_3963,N_3774,N_3784);
and U3964 (N_3964,N_3747,N_3703);
nor U3965 (N_3965,N_3659,N_3688);
and U3966 (N_3966,N_3749,N_3761);
nor U3967 (N_3967,N_3762,N_3790);
and U3968 (N_3968,N_3613,N_3624);
nor U3969 (N_3969,N_3704,N_3640);
xor U3970 (N_3970,N_3792,N_3771);
xor U3971 (N_3971,N_3690,N_3610);
nor U3972 (N_3972,N_3724,N_3673);
nand U3973 (N_3973,N_3674,N_3771);
nor U3974 (N_3974,N_3629,N_3729);
and U3975 (N_3975,N_3678,N_3718);
and U3976 (N_3976,N_3750,N_3654);
nor U3977 (N_3977,N_3603,N_3711);
xnor U3978 (N_3978,N_3673,N_3601);
nor U3979 (N_3979,N_3756,N_3643);
xor U3980 (N_3980,N_3620,N_3683);
and U3981 (N_3981,N_3798,N_3625);
xor U3982 (N_3982,N_3624,N_3641);
and U3983 (N_3983,N_3761,N_3785);
nor U3984 (N_3984,N_3729,N_3686);
xor U3985 (N_3985,N_3713,N_3723);
nor U3986 (N_3986,N_3784,N_3793);
and U3987 (N_3987,N_3732,N_3655);
nand U3988 (N_3988,N_3669,N_3675);
xor U3989 (N_3989,N_3796,N_3764);
xnor U3990 (N_3990,N_3715,N_3744);
nor U3991 (N_3991,N_3681,N_3721);
nor U3992 (N_3992,N_3646,N_3754);
xnor U3993 (N_3993,N_3607,N_3782);
nor U3994 (N_3994,N_3714,N_3675);
or U3995 (N_3995,N_3604,N_3686);
nor U3996 (N_3996,N_3788,N_3602);
xnor U3997 (N_3997,N_3688,N_3728);
nor U3998 (N_3998,N_3789,N_3785);
xnor U3999 (N_3999,N_3678,N_3789);
and U4000 (N_4000,N_3944,N_3935);
nor U4001 (N_4001,N_3972,N_3884);
nor U4002 (N_4002,N_3986,N_3918);
nand U4003 (N_4003,N_3949,N_3899);
and U4004 (N_4004,N_3859,N_3874);
or U4005 (N_4005,N_3869,N_3921);
nand U4006 (N_4006,N_3922,N_3805);
and U4007 (N_4007,N_3945,N_3929);
nor U4008 (N_4008,N_3973,N_3821);
and U4009 (N_4009,N_3910,N_3837);
xnor U4010 (N_4010,N_3810,N_3822);
nand U4011 (N_4011,N_3906,N_3917);
nor U4012 (N_4012,N_3872,N_3852);
nor U4013 (N_4013,N_3926,N_3901);
and U4014 (N_4014,N_3824,N_3849);
nand U4015 (N_4015,N_3877,N_3825);
nand U4016 (N_4016,N_3947,N_3826);
nor U4017 (N_4017,N_3955,N_3807);
nor U4018 (N_4018,N_3913,N_3931);
or U4019 (N_4019,N_3943,N_3878);
or U4020 (N_4020,N_3843,N_3881);
nor U4021 (N_4021,N_3948,N_3978);
nor U4022 (N_4022,N_3862,N_3989);
or U4023 (N_4023,N_3924,N_3984);
xnor U4024 (N_4024,N_3836,N_3827);
or U4025 (N_4025,N_3936,N_3971);
xnor U4026 (N_4026,N_3991,N_3806);
and U4027 (N_4027,N_3815,N_3992);
nand U4028 (N_4028,N_3932,N_3856);
and U4029 (N_4029,N_3829,N_3858);
and U4030 (N_4030,N_3867,N_3847);
xor U4031 (N_4031,N_3930,N_3855);
xnor U4032 (N_4032,N_3850,N_3934);
nor U4033 (N_4033,N_3832,N_3817);
xor U4034 (N_4034,N_3960,N_3942);
or U4035 (N_4035,N_3889,N_3959);
nand U4036 (N_4036,N_3893,N_3954);
nand U4037 (N_4037,N_3802,N_3941);
or U4038 (N_4038,N_3903,N_3923);
or U4039 (N_4039,N_3813,N_3896);
and U4040 (N_4040,N_3857,N_3828);
xor U4041 (N_4041,N_3981,N_3995);
and U4042 (N_4042,N_3964,N_3915);
nor U4043 (N_4043,N_3838,N_3839);
nor U4044 (N_4044,N_3808,N_3845);
and U4045 (N_4045,N_3868,N_3844);
and U4046 (N_4046,N_3834,N_3866);
and U4047 (N_4047,N_3979,N_3974);
or U4048 (N_4048,N_3993,N_3916);
nor U4049 (N_4049,N_3909,N_3886);
and U4050 (N_4050,N_3919,N_3871);
xnor U4051 (N_4051,N_3863,N_3880);
or U4052 (N_4052,N_3894,N_3933);
nand U4053 (N_4053,N_3800,N_3983);
nand U4054 (N_4054,N_3883,N_3890);
and U4055 (N_4055,N_3965,N_3908);
or U4056 (N_4056,N_3892,N_3876);
or U4057 (N_4057,N_3968,N_3854);
nor U4058 (N_4058,N_3804,N_3885);
nor U4059 (N_4059,N_3803,N_3996);
nand U4060 (N_4060,N_3814,N_3898);
nand U4061 (N_4061,N_3976,N_3985);
or U4062 (N_4062,N_3879,N_3911);
or U4063 (N_4063,N_3952,N_3953);
nand U4064 (N_4064,N_3994,N_3895);
and U4065 (N_4065,N_3946,N_3870);
nand U4066 (N_4066,N_3820,N_3969);
and U4067 (N_4067,N_3990,N_3835);
xnor U4068 (N_4068,N_3875,N_3816);
nor U4069 (N_4069,N_3887,N_3823);
nand U4070 (N_4070,N_3966,N_3865);
nand U4071 (N_4071,N_3925,N_3891);
or U4072 (N_4072,N_3853,N_3846);
and U4073 (N_4073,N_3961,N_3904);
or U4074 (N_4074,N_3900,N_3998);
or U4075 (N_4075,N_3905,N_3980);
nand U4076 (N_4076,N_3907,N_3956);
xnor U4077 (N_4077,N_3902,N_3848);
nand U4078 (N_4078,N_3975,N_3912);
nor U4079 (N_4079,N_3939,N_3967);
and U4080 (N_4080,N_3819,N_3861);
xnor U4081 (N_4081,N_3833,N_3811);
nor U4082 (N_4082,N_3873,N_3987);
and U4083 (N_4083,N_3982,N_3977);
nor U4084 (N_4084,N_3914,N_3951);
and U4085 (N_4085,N_3927,N_3997);
or U4086 (N_4086,N_3957,N_3864);
xnor U4087 (N_4087,N_3840,N_3958);
xnor U4088 (N_4088,N_3812,N_3938);
nor U4089 (N_4089,N_3801,N_3842);
or U4090 (N_4090,N_3970,N_3963);
or U4091 (N_4091,N_3897,N_3928);
or U4092 (N_4092,N_3830,N_3831);
nor U4093 (N_4093,N_3888,N_3988);
and U4094 (N_4094,N_3818,N_3940);
nand U4095 (N_4095,N_3860,N_3841);
or U4096 (N_4096,N_3882,N_3962);
xor U4097 (N_4097,N_3999,N_3851);
nand U4098 (N_4098,N_3950,N_3920);
and U4099 (N_4099,N_3937,N_3809);
nand U4100 (N_4100,N_3915,N_3806);
or U4101 (N_4101,N_3905,N_3806);
xor U4102 (N_4102,N_3869,N_3957);
nor U4103 (N_4103,N_3961,N_3936);
nand U4104 (N_4104,N_3896,N_3981);
and U4105 (N_4105,N_3882,N_3968);
nand U4106 (N_4106,N_3827,N_3876);
nor U4107 (N_4107,N_3803,N_3819);
and U4108 (N_4108,N_3994,N_3850);
and U4109 (N_4109,N_3995,N_3990);
xor U4110 (N_4110,N_3919,N_3976);
or U4111 (N_4111,N_3991,N_3832);
nand U4112 (N_4112,N_3916,N_3812);
nor U4113 (N_4113,N_3943,N_3986);
xor U4114 (N_4114,N_3944,N_3819);
xnor U4115 (N_4115,N_3936,N_3897);
or U4116 (N_4116,N_3957,N_3832);
or U4117 (N_4117,N_3818,N_3921);
or U4118 (N_4118,N_3839,N_3957);
nand U4119 (N_4119,N_3888,N_3884);
nor U4120 (N_4120,N_3825,N_3964);
nor U4121 (N_4121,N_3833,N_3823);
nand U4122 (N_4122,N_3894,N_3807);
nand U4123 (N_4123,N_3939,N_3855);
nor U4124 (N_4124,N_3953,N_3975);
and U4125 (N_4125,N_3927,N_3966);
or U4126 (N_4126,N_3833,N_3956);
nor U4127 (N_4127,N_3815,N_3879);
nor U4128 (N_4128,N_3924,N_3980);
xnor U4129 (N_4129,N_3901,N_3804);
or U4130 (N_4130,N_3982,N_3888);
nor U4131 (N_4131,N_3829,N_3993);
or U4132 (N_4132,N_3889,N_3902);
and U4133 (N_4133,N_3973,N_3909);
xor U4134 (N_4134,N_3829,N_3850);
or U4135 (N_4135,N_3865,N_3975);
or U4136 (N_4136,N_3947,N_3904);
nor U4137 (N_4137,N_3816,N_3915);
and U4138 (N_4138,N_3814,N_3943);
and U4139 (N_4139,N_3958,N_3990);
xor U4140 (N_4140,N_3931,N_3894);
nand U4141 (N_4141,N_3980,N_3990);
and U4142 (N_4142,N_3943,N_3890);
xnor U4143 (N_4143,N_3808,N_3905);
or U4144 (N_4144,N_3919,N_3928);
xnor U4145 (N_4145,N_3839,N_3962);
nor U4146 (N_4146,N_3882,N_3944);
or U4147 (N_4147,N_3817,N_3889);
nand U4148 (N_4148,N_3948,N_3932);
nand U4149 (N_4149,N_3997,N_3899);
or U4150 (N_4150,N_3913,N_3861);
nand U4151 (N_4151,N_3981,N_3827);
nor U4152 (N_4152,N_3968,N_3894);
or U4153 (N_4153,N_3943,N_3842);
nand U4154 (N_4154,N_3818,N_3881);
nor U4155 (N_4155,N_3829,N_3967);
and U4156 (N_4156,N_3814,N_3890);
nor U4157 (N_4157,N_3959,N_3816);
and U4158 (N_4158,N_3807,N_3988);
nor U4159 (N_4159,N_3843,N_3989);
nand U4160 (N_4160,N_3864,N_3941);
nor U4161 (N_4161,N_3854,N_3974);
nor U4162 (N_4162,N_3988,N_3962);
nor U4163 (N_4163,N_3835,N_3918);
nand U4164 (N_4164,N_3840,N_3839);
or U4165 (N_4165,N_3821,N_3937);
xor U4166 (N_4166,N_3960,N_3913);
and U4167 (N_4167,N_3826,N_3846);
nand U4168 (N_4168,N_3869,N_3903);
nor U4169 (N_4169,N_3986,N_3904);
and U4170 (N_4170,N_3976,N_3837);
xor U4171 (N_4171,N_3982,N_3825);
nor U4172 (N_4172,N_3820,N_3990);
xor U4173 (N_4173,N_3893,N_3897);
and U4174 (N_4174,N_3939,N_3941);
xor U4175 (N_4175,N_3995,N_3914);
xnor U4176 (N_4176,N_3884,N_3849);
nand U4177 (N_4177,N_3811,N_3848);
nor U4178 (N_4178,N_3955,N_3855);
nor U4179 (N_4179,N_3828,N_3939);
xor U4180 (N_4180,N_3877,N_3996);
nor U4181 (N_4181,N_3893,N_3830);
nor U4182 (N_4182,N_3988,N_3918);
or U4183 (N_4183,N_3855,N_3816);
nand U4184 (N_4184,N_3853,N_3875);
xnor U4185 (N_4185,N_3812,N_3872);
and U4186 (N_4186,N_3925,N_3907);
xnor U4187 (N_4187,N_3877,N_3949);
or U4188 (N_4188,N_3828,N_3844);
nand U4189 (N_4189,N_3806,N_3953);
nor U4190 (N_4190,N_3871,N_3895);
xnor U4191 (N_4191,N_3807,N_3801);
or U4192 (N_4192,N_3880,N_3908);
xnor U4193 (N_4193,N_3991,N_3804);
xor U4194 (N_4194,N_3892,N_3842);
nand U4195 (N_4195,N_3943,N_3993);
xor U4196 (N_4196,N_3940,N_3981);
and U4197 (N_4197,N_3937,N_3886);
nor U4198 (N_4198,N_3812,N_3899);
or U4199 (N_4199,N_3902,N_3978);
nand U4200 (N_4200,N_4079,N_4081);
nor U4201 (N_4201,N_4130,N_4008);
and U4202 (N_4202,N_4192,N_4014);
nand U4203 (N_4203,N_4110,N_4027);
nand U4204 (N_4204,N_4120,N_4126);
nor U4205 (N_4205,N_4167,N_4029);
xor U4206 (N_4206,N_4197,N_4077);
or U4207 (N_4207,N_4090,N_4051);
nor U4208 (N_4208,N_4125,N_4164);
or U4209 (N_4209,N_4054,N_4095);
nand U4210 (N_4210,N_4002,N_4046);
xnor U4211 (N_4211,N_4104,N_4086);
nor U4212 (N_4212,N_4025,N_4012);
nand U4213 (N_4213,N_4185,N_4033);
nand U4214 (N_4214,N_4088,N_4039);
and U4215 (N_4215,N_4038,N_4007);
nand U4216 (N_4216,N_4177,N_4028);
xor U4217 (N_4217,N_4063,N_4065);
and U4218 (N_4218,N_4089,N_4070);
or U4219 (N_4219,N_4073,N_4119);
xnor U4220 (N_4220,N_4024,N_4064);
nand U4221 (N_4221,N_4170,N_4022);
nor U4222 (N_4222,N_4092,N_4004);
or U4223 (N_4223,N_4153,N_4032);
or U4224 (N_4224,N_4041,N_4031);
nor U4225 (N_4225,N_4067,N_4140);
nand U4226 (N_4226,N_4159,N_4176);
nor U4227 (N_4227,N_4040,N_4056);
or U4228 (N_4228,N_4163,N_4115);
nand U4229 (N_4229,N_4009,N_4050);
nor U4230 (N_4230,N_4179,N_4103);
xnor U4231 (N_4231,N_4133,N_4048);
nor U4232 (N_4232,N_4053,N_4187);
or U4233 (N_4233,N_4148,N_4193);
nor U4234 (N_4234,N_4047,N_4134);
nand U4235 (N_4235,N_4083,N_4138);
nor U4236 (N_4236,N_4161,N_4108);
or U4237 (N_4237,N_4122,N_4175);
nand U4238 (N_4238,N_4173,N_4144);
xor U4239 (N_4239,N_4107,N_4160);
nor U4240 (N_4240,N_4150,N_4182);
and U4241 (N_4241,N_4172,N_4016);
nand U4242 (N_4242,N_4001,N_4184);
or U4243 (N_4243,N_4093,N_4194);
and U4244 (N_4244,N_4037,N_4174);
xor U4245 (N_4245,N_4074,N_4082);
nor U4246 (N_4246,N_4178,N_4114);
or U4247 (N_4247,N_4106,N_4015);
and U4248 (N_4248,N_4198,N_4034);
xnor U4249 (N_4249,N_4075,N_4141);
and U4250 (N_4250,N_4078,N_4196);
nor U4251 (N_4251,N_4005,N_4019);
xnor U4252 (N_4252,N_4036,N_4100);
or U4253 (N_4253,N_4169,N_4094);
xnor U4254 (N_4254,N_4139,N_4017);
or U4255 (N_4255,N_4098,N_4101);
xor U4256 (N_4256,N_4069,N_4151);
and U4257 (N_4257,N_4066,N_4080);
xnor U4258 (N_4258,N_4146,N_4072);
or U4259 (N_4259,N_4062,N_4155);
nand U4260 (N_4260,N_4044,N_4023);
nand U4261 (N_4261,N_4042,N_4118);
nor U4262 (N_4262,N_4189,N_4030);
xnor U4263 (N_4263,N_4112,N_4097);
and U4264 (N_4264,N_4055,N_4102);
and U4265 (N_4265,N_4128,N_4188);
or U4266 (N_4266,N_4137,N_4035);
nand U4267 (N_4267,N_4010,N_4135);
xor U4268 (N_4268,N_4096,N_4171);
and U4269 (N_4269,N_4149,N_4154);
and U4270 (N_4270,N_4057,N_4156);
xnor U4271 (N_4271,N_4043,N_4168);
nand U4272 (N_4272,N_4180,N_4013);
nand U4273 (N_4273,N_4132,N_4157);
nor U4274 (N_4274,N_4111,N_4116);
nor U4275 (N_4275,N_4026,N_4052);
nand U4276 (N_4276,N_4186,N_4131);
nand U4277 (N_4277,N_4113,N_4045);
or U4278 (N_4278,N_4076,N_4183);
nor U4279 (N_4279,N_4003,N_4021);
nand U4280 (N_4280,N_4006,N_4145);
or U4281 (N_4281,N_4117,N_4147);
nor U4282 (N_4282,N_4124,N_4087);
nand U4283 (N_4283,N_4058,N_4166);
and U4284 (N_4284,N_4091,N_4142);
nand U4285 (N_4285,N_4190,N_4085);
nor U4286 (N_4286,N_4191,N_4195);
nor U4287 (N_4287,N_4121,N_4127);
nor U4288 (N_4288,N_4060,N_4136);
and U4289 (N_4289,N_4158,N_4143);
or U4290 (N_4290,N_4165,N_4049);
and U4291 (N_4291,N_4061,N_4105);
xnor U4292 (N_4292,N_4071,N_4059);
nand U4293 (N_4293,N_4099,N_4018);
or U4294 (N_4294,N_4199,N_4129);
and U4295 (N_4295,N_4162,N_4123);
nand U4296 (N_4296,N_4152,N_4011);
nand U4297 (N_4297,N_4084,N_4181);
or U4298 (N_4298,N_4020,N_4109);
nor U4299 (N_4299,N_4068,N_4000);
nand U4300 (N_4300,N_4163,N_4165);
nand U4301 (N_4301,N_4117,N_4042);
or U4302 (N_4302,N_4197,N_4195);
and U4303 (N_4303,N_4115,N_4181);
or U4304 (N_4304,N_4115,N_4194);
or U4305 (N_4305,N_4088,N_4096);
nor U4306 (N_4306,N_4061,N_4098);
nor U4307 (N_4307,N_4016,N_4166);
xnor U4308 (N_4308,N_4103,N_4064);
nor U4309 (N_4309,N_4094,N_4138);
or U4310 (N_4310,N_4146,N_4185);
xnor U4311 (N_4311,N_4068,N_4171);
or U4312 (N_4312,N_4090,N_4113);
nor U4313 (N_4313,N_4130,N_4019);
nand U4314 (N_4314,N_4093,N_4024);
or U4315 (N_4315,N_4057,N_4095);
or U4316 (N_4316,N_4183,N_4074);
and U4317 (N_4317,N_4121,N_4013);
xor U4318 (N_4318,N_4098,N_4051);
nand U4319 (N_4319,N_4185,N_4152);
xnor U4320 (N_4320,N_4133,N_4023);
xor U4321 (N_4321,N_4146,N_4090);
and U4322 (N_4322,N_4117,N_4077);
and U4323 (N_4323,N_4198,N_4064);
xnor U4324 (N_4324,N_4165,N_4147);
xnor U4325 (N_4325,N_4130,N_4111);
or U4326 (N_4326,N_4188,N_4129);
nand U4327 (N_4327,N_4008,N_4052);
or U4328 (N_4328,N_4153,N_4107);
and U4329 (N_4329,N_4194,N_4123);
or U4330 (N_4330,N_4193,N_4059);
and U4331 (N_4331,N_4140,N_4032);
and U4332 (N_4332,N_4009,N_4163);
and U4333 (N_4333,N_4164,N_4100);
nand U4334 (N_4334,N_4109,N_4037);
or U4335 (N_4335,N_4069,N_4048);
nor U4336 (N_4336,N_4179,N_4092);
nand U4337 (N_4337,N_4060,N_4007);
nor U4338 (N_4338,N_4056,N_4188);
xor U4339 (N_4339,N_4195,N_4188);
nand U4340 (N_4340,N_4056,N_4164);
xor U4341 (N_4341,N_4109,N_4175);
xor U4342 (N_4342,N_4094,N_4047);
nand U4343 (N_4343,N_4123,N_4034);
and U4344 (N_4344,N_4141,N_4006);
or U4345 (N_4345,N_4144,N_4160);
nor U4346 (N_4346,N_4132,N_4067);
xnor U4347 (N_4347,N_4017,N_4167);
xnor U4348 (N_4348,N_4069,N_4169);
xnor U4349 (N_4349,N_4148,N_4106);
nor U4350 (N_4350,N_4087,N_4094);
and U4351 (N_4351,N_4128,N_4016);
and U4352 (N_4352,N_4035,N_4119);
xnor U4353 (N_4353,N_4115,N_4113);
nor U4354 (N_4354,N_4077,N_4091);
nand U4355 (N_4355,N_4044,N_4053);
xnor U4356 (N_4356,N_4030,N_4015);
nand U4357 (N_4357,N_4115,N_4179);
nor U4358 (N_4358,N_4006,N_4110);
nand U4359 (N_4359,N_4018,N_4071);
or U4360 (N_4360,N_4019,N_4020);
or U4361 (N_4361,N_4053,N_4128);
nand U4362 (N_4362,N_4049,N_4001);
nand U4363 (N_4363,N_4140,N_4153);
and U4364 (N_4364,N_4011,N_4139);
xor U4365 (N_4365,N_4096,N_4102);
nand U4366 (N_4366,N_4084,N_4175);
xor U4367 (N_4367,N_4056,N_4045);
xnor U4368 (N_4368,N_4121,N_4061);
and U4369 (N_4369,N_4148,N_4152);
nand U4370 (N_4370,N_4023,N_4015);
nand U4371 (N_4371,N_4037,N_4158);
nand U4372 (N_4372,N_4105,N_4153);
and U4373 (N_4373,N_4053,N_4134);
xor U4374 (N_4374,N_4084,N_4135);
or U4375 (N_4375,N_4037,N_4156);
nor U4376 (N_4376,N_4140,N_4193);
nor U4377 (N_4377,N_4133,N_4078);
and U4378 (N_4378,N_4157,N_4021);
nand U4379 (N_4379,N_4194,N_4141);
xor U4380 (N_4380,N_4128,N_4127);
nor U4381 (N_4381,N_4149,N_4106);
and U4382 (N_4382,N_4023,N_4059);
xor U4383 (N_4383,N_4140,N_4125);
and U4384 (N_4384,N_4002,N_4004);
nor U4385 (N_4385,N_4120,N_4062);
and U4386 (N_4386,N_4031,N_4183);
nand U4387 (N_4387,N_4113,N_4012);
or U4388 (N_4388,N_4109,N_4081);
and U4389 (N_4389,N_4022,N_4005);
xor U4390 (N_4390,N_4036,N_4023);
nor U4391 (N_4391,N_4065,N_4131);
nor U4392 (N_4392,N_4101,N_4173);
and U4393 (N_4393,N_4011,N_4026);
and U4394 (N_4394,N_4116,N_4054);
or U4395 (N_4395,N_4084,N_4164);
and U4396 (N_4396,N_4181,N_4128);
or U4397 (N_4397,N_4147,N_4017);
nor U4398 (N_4398,N_4013,N_4102);
or U4399 (N_4399,N_4058,N_4197);
and U4400 (N_4400,N_4307,N_4251);
xnor U4401 (N_4401,N_4294,N_4396);
and U4402 (N_4402,N_4298,N_4218);
nor U4403 (N_4403,N_4332,N_4375);
or U4404 (N_4404,N_4272,N_4237);
and U4405 (N_4405,N_4327,N_4285);
or U4406 (N_4406,N_4235,N_4341);
nor U4407 (N_4407,N_4348,N_4368);
and U4408 (N_4408,N_4271,N_4270);
nor U4409 (N_4409,N_4395,N_4373);
nand U4410 (N_4410,N_4352,N_4391);
xnor U4411 (N_4411,N_4293,N_4282);
and U4412 (N_4412,N_4369,N_4222);
and U4413 (N_4413,N_4258,N_4220);
and U4414 (N_4414,N_4232,N_4217);
or U4415 (N_4415,N_4339,N_4316);
xor U4416 (N_4416,N_4288,N_4241);
and U4417 (N_4417,N_4228,N_4287);
nor U4418 (N_4418,N_4215,N_4301);
nor U4419 (N_4419,N_4315,N_4336);
and U4420 (N_4420,N_4312,N_4351);
nand U4421 (N_4421,N_4345,N_4299);
nor U4422 (N_4422,N_4381,N_4303);
or U4423 (N_4423,N_4328,N_4394);
and U4424 (N_4424,N_4249,N_4261);
nand U4425 (N_4425,N_4386,N_4234);
or U4426 (N_4426,N_4262,N_4364);
nor U4427 (N_4427,N_4239,N_4275);
nand U4428 (N_4428,N_4240,N_4242);
and U4429 (N_4429,N_4280,N_4384);
nand U4430 (N_4430,N_4357,N_4284);
or U4431 (N_4431,N_4231,N_4319);
or U4432 (N_4432,N_4359,N_4387);
xnor U4433 (N_4433,N_4318,N_4245);
and U4434 (N_4434,N_4211,N_4207);
nand U4435 (N_4435,N_4221,N_4355);
nand U4436 (N_4436,N_4212,N_4233);
xnor U4437 (N_4437,N_4229,N_4246);
or U4438 (N_4438,N_4398,N_4354);
xor U4439 (N_4439,N_4290,N_4252);
xor U4440 (N_4440,N_4302,N_4356);
nor U4441 (N_4441,N_4238,N_4362);
xnor U4442 (N_4442,N_4347,N_4392);
or U4443 (N_4443,N_4291,N_4204);
and U4444 (N_4444,N_4340,N_4297);
or U4445 (N_4445,N_4289,N_4338);
nor U4446 (N_4446,N_4264,N_4324);
or U4447 (N_4447,N_4283,N_4236);
and U4448 (N_4448,N_4334,N_4317);
nand U4449 (N_4449,N_4206,N_4247);
xor U4450 (N_4450,N_4311,N_4276);
nand U4451 (N_4451,N_4329,N_4335);
nand U4452 (N_4452,N_4333,N_4230);
nand U4453 (N_4453,N_4397,N_4343);
xnor U4454 (N_4454,N_4277,N_4265);
xnor U4455 (N_4455,N_4292,N_4380);
nand U4456 (N_4456,N_4323,N_4353);
nor U4457 (N_4457,N_4337,N_4313);
xnor U4458 (N_4458,N_4349,N_4260);
xnor U4459 (N_4459,N_4296,N_4378);
nor U4460 (N_4460,N_4300,N_4366);
nand U4461 (N_4461,N_4320,N_4255);
and U4462 (N_4462,N_4267,N_4205);
or U4463 (N_4463,N_4309,N_4254);
nor U4464 (N_4464,N_4266,N_4304);
nor U4465 (N_4465,N_4393,N_4257);
or U4466 (N_4466,N_4225,N_4379);
nor U4467 (N_4467,N_4216,N_4263);
nor U4468 (N_4468,N_4306,N_4253);
and U4469 (N_4469,N_4259,N_4342);
xor U4470 (N_4470,N_4273,N_4363);
and U4471 (N_4471,N_4269,N_4250);
nand U4472 (N_4472,N_4248,N_4360);
and U4473 (N_4473,N_4202,N_4390);
nand U4474 (N_4474,N_4308,N_4376);
or U4475 (N_4475,N_4344,N_4331);
nor U4476 (N_4476,N_4281,N_4389);
xnor U4477 (N_4477,N_4224,N_4358);
and U4478 (N_4478,N_4322,N_4370);
and U4479 (N_4479,N_4374,N_4382);
and U4480 (N_4480,N_4325,N_4219);
nor U4481 (N_4481,N_4274,N_4209);
nand U4482 (N_4482,N_4244,N_4201);
nor U4483 (N_4483,N_4326,N_4346);
and U4484 (N_4484,N_4321,N_4279);
nand U4485 (N_4485,N_4383,N_4367);
nand U4486 (N_4486,N_4227,N_4243);
and U4487 (N_4487,N_4214,N_4365);
nor U4488 (N_4488,N_4286,N_4226);
xnor U4489 (N_4489,N_4385,N_4305);
or U4490 (N_4490,N_4377,N_4372);
xor U4491 (N_4491,N_4223,N_4361);
and U4492 (N_4492,N_4399,N_4200);
nand U4493 (N_4493,N_4208,N_4256);
or U4494 (N_4494,N_4314,N_4350);
xnor U4495 (N_4495,N_4310,N_4371);
nand U4496 (N_4496,N_4210,N_4295);
and U4497 (N_4497,N_4268,N_4330);
xor U4498 (N_4498,N_4388,N_4213);
xnor U4499 (N_4499,N_4203,N_4278);
nor U4500 (N_4500,N_4374,N_4278);
nand U4501 (N_4501,N_4319,N_4298);
nor U4502 (N_4502,N_4330,N_4201);
and U4503 (N_4503,N_4365,N_4293);
or U4504 (N_4504,N_4243,N_4296);
nor U4505 (N_4505,N_4271,N_4321);
xor U4506 (N_4506,N_4341,N_4381);
and U4507 (N_4507,N_4201,N_4299);
xnor U4508 (N_4508,N_4205,N_4289);
xor U4509 (N_4509,N_4310,N_4390);
nor U4510 (N_4510,N_4274,N_4395);
and U4511 (N_4511,N_4369,N_4295);
nand U4512 (N_4512,N_4278,N_4385);
nand U4513 (N_4513,N_4398,N_4273);
nand U4514 (N_4514,N_4214,N_4355);
or U4515 (N_4515,N_4280,N_4263);
and U4516 (N_4516,N_4297,N_4243);
xnor U4517 (N_4517,N_4322,N_4271);
nand U4518 (N_4518,N_4363,N_4300);
xnor U4519 (N_4519,N_4274,N_4318);
nand U4520 (N_4520,N_4210,N_4271);
or U4521 (N_4521,N_4377,N_4390);
nor U4522 (N_4522,N_4276,N_4281);
nand U4523 (N_4523,N_4288,N_4314);
xor U4524 (N_4524,N_4228,N_4336);
nor U4525 (N_4525,N_4398,N_4201);
and U4526 (N_4526,N_4313,N_4307);
nor U4527 (N_4527,N_4263,N_4365);
xor U4528 (N_4528,N_4201,N_4352);
and U4529 (N_4529,N_4208,N_4292);
nand U4530 (N_4530,N_4352,N_4218);
nand U4531 (N_4531,N_4333,N_4246);
and U4532 (N_4532,N_4228,N_4305);
nand U4533 (N_4533,N_4296,N_4385);
nor U4534 (N_4534,N_4332,N_4369);
nor U4535 (N_4535,N_4285,N_4258);
xnor U4536 (N_4536,N_4363,N_4281);
or U4537 (N_4537,N_4325,N_4205);
nand U4538 (N_4538,N_4353,N_4289);
xnor U4539 (N_4539,N_4244,N_4217);
or U4540 (N_4540,N_4381,N_4256);
and U4541 (N_4541,N_4379,N_4358);
nor U4542 (N_4542,N_4371,N_4314);
nand U4543 (N_4543,N_4241,N_4335);
or U4544 (N_4544,N_4288,N_4293);
xnor U4545 (N_4545,N_4360,N_4264);
and U4546 (N_4546,N_4338,N_4258);
nand U4547 (N_4547,N_4251,N_4380);
nor U4548 (N_4548,N_4343,N_4303);
and U4549 (N_4549,N_4230,N_4209);
nor U4550 (N_4550,N_4333,N_4287);
nor U4551 (N_4551,N_4385,N_4221);
nand U4552 (N_4552,N_4306,N_4337);
nand U4553 (N_4553,N_4292,N_4231);
nand U4554 (N_4554,N_4382,N_4248);
nand U4555 (N_4555,N_4227,N_4383);
nor U4556 (N_4556,N_4358,N_4212);
nor U4557 (N_4557,N_4329,N_4364);
and U4558 (N_4558,N_4234,N_4285);
nor U4559 (N_4559,N_4361,N_4227);
or U4560 (N_4560,N_4362,N_4204);
xnor U4561 (N_4561,N_4213,N_4297);
nand U4562 (N_4562,N_4357,N_4228);
nand U4563 (N_4563,N_4270,N_4309);
and U4564 (N_4564,N_4243,N_4244);
or U4565 (N_4565,N_4314,N_4247);
nand U4566 (N_4566,N_4378,N_4281);
nor U4567 (N_4567,N_4244,N_4327);
xnor U4568 (N_4568,N_4301,N_4380);
and U4569 (N_4569,N_4207,N_4357);
and U4570 (N_4570,N_4327,N_4214);
nand U4571 (N_4571,N_4392,N_4300);
and U4572 (N_4572,N_4220,N_4327);
nand U4573 (N_4573,N_4304,N_4257);
nand U4574 (N_4574,N_4386,N_4327);
nand U4575 (N_4575,N_4270,N_4203);
or U4576 (N_4576,N_4252,N_4211);
nor U4577 (N_4577,N_4388,N_4368);
nor U4578 (N_4578,N_4360,N_4368);
and U4579 (N_4579,N_4322,N_4377);
and U4580 (N_4580,N_4304,N_4273);
and U4581 (N_4581,N_4222,N_4392);
nand U4582 (N_4582,N_4231,N_4379);
xor U4583 (N_4583,N_4366,N_4227);
or U4584 (N_4584,N_4219,N_4327);
nand U4585 (N_4585,N_4232,N_4273);
nand U4586 (N_4586,N_4335,N_4309);
xor U4587 (N_4587,N_4397,N_4203);
or U4588 (N_4588,N_4352,N_4305);
xnor U4589 (N_4589,N_4246,N_4256);
and U4590 (N_4590,N_4346,N_4256);
nor U4591 (N_4591,N_4370,N_4329);
nand U4592 (N_4592,N_4338,N_4329);
nor U4593 (N_4593,N_4232,N_4243);
and U4594 (N_4594,N_4332,N_4319);
or U4595 (N_4595,N_4320,N_4302);
nand U4596 (N_4596,N_4352,N_4368);
nor U4597 (N_4597,N_4266,N_4262);
and U4598 (N_4598,N_4220,N_4237);
nand U4599 (N_4599,N_4200,N_4359);
nand U4600 (N_4600,N_4599,N_4580);
and U4601 (N_4601,N_4473,N_4520);
nand U4602 (N_4602,N_4479,N_4405);
and U4603 (N_4603,N_4558,N_4478);
xor U4604 (N_4604,N_4496,N_4453);
nand U4605 (N_4605,N_4560,N_4494);
nor U4606 (N_4606,N_4505,N_4504);
nand U4607 (N_4607,N_4549,N_4433);
nor U4608 (N_4608,N_4484,N_4528);
nand U4609 (N_4609,N_4537,N_4567);
xnor U4610 (N_4610,N_4446,N_4429);
nand U4611 (N_4611,N_4527,N_4532);
nand U4612 (N_4612,N_4579,N_4559);
nor U4613 (N_4613,N_4465,N_4462);
xnor U4614 (N_4614,N_4404,N_4459);
or U4615 (N_4615,N_4587,N_4486);
and U4616 (N_4616,N_4588,N_4454);
nor U4617 (N_4617,N_4590,N_4416);
xor U4618 (N_4618,N_4447,N_4535);
xor U4619 (N_4619,N_4491,N_4492);
nand U4620 (N_4620,N_4557,N_4452);
and U4621 (N_4621,N_4461,N_4403);
nor U4622 (N_4622,N_4570,N_4544);
and U4623 (N_4623,N_4450,N_4519);
nand U4624 (N_4624,N_4449,N_4583);
nor U4625 (N_4625,N_4445,N_4418);
nor U4626 (N_4626,N_4586,N_4421);
xor U4627 (N_4627,N_4551,N_4594);
xor U4628 (N_4628,N_4460,N_4414);
nand U4629 (N_4629,N_4493,N_4472);
nand U4630 (N_4630,N_4543,N_4555);
or U4631 (N_4631,N_4516,N_4485);
and U4632 (N_4632,N_4408,N_4430);
xor U4633 (N_4633,N_4510,N_4524);
and U4634 (N_4634,N_4565,N_4498);
nand U4635 (N_4635,N_4495,N_4578);
nor U4636 (N_4636,N_4435,N_4471);
and U4637 (N_4637,N_4434,N_4514);
and U4638 (N_4638,N_4584,N_4536);
or U4639 (N_4639,N_4585,N_4523);
or U4640 (N_4640,N_4562,N_4547);
xor U4641 (N_4641,N_4458,N_4515);
xor U4642 (N_4642,N_4553,N_4468);
nor U4643 (N_4643,N_4508,N_4596);
or U4644 (N_4644,N_4542,N_4469);
or U4645 (N_4645,N_4503,N_4406);
and U4646 (N_4646,N_4538,N_4425);
xnor U4647 (N_4647,N_4428,N_4455);
xor U4648 (N_4648,N_4420,N_4534);
and U4649 (N_4649,N_4442,N_4502);
and U4650 (N_4650,N_4439,N_4554);
xnor U4651 (N_4651,N_4499,N_4480);
nor U4652 (N_4652,N_4563,N_4571);
nand U4653 (N_4653,N_4507,N_4598);
xnor U4654 (N_4654,N_4443,N_4540);
or U4655 (N_4655,N_4561,N_4476);
nand U4656 (N_4656,N_4417,N_4566);
nand U4657 (N_4657,N_4556,N_4501);
nor U4658 (N_4658,N_4597,N_4409);
or U4659 (N_4659,N_4474,N_4402);
xor U4660 (N_4660,N_4531,N_4470);
and U4661 (N_4661,N_4546,N_4422);
xnor U4662 (N_4662,N_4483,N_4575);
or U4663 (N_4663,N_4550,N_4545);
nand U4664 (N_4664,N_4490,N_4518);
xnor U4665 (N_4665,N_4463,N_4456);
xor U4666 (N_4666,N_4400,N_4592);
nor U4667 (N_4667,N_4441,N_4477);
and U4668 (N_4668,N_4438,N_4451);
nor U4669 (N_4669,N_4457,N_4407);
xor U4670 (N_4670,N_4552,N_4467);
nor U4671 (N_4671,N_4521,N_4413);
or U4672 (N_4672,N_4436,N_4426);
or U4673 (N_4673,N_4431,N_4424);
xnor U4674 (N_4674,N_4412,N_4512);
nand U4675 (N_4675,N_4589,N_4569);
or U4676 (N_4676,N_4573,N_4432);
nand U4677 (N_4677,N_4509,N_4574);
or U4678 (N_4678,N_4577,N_4482);
nor U4679 (N_4679,N_4410,N_4437);
nand U4680 (N_4680,N_4481,N_4564);
xnor U4681 (N_4681,N_4541,N_4440);
or U4682 (N_4682,N_4464,N_4530);
or U4683 (N_4683,N_4411,N_4593);
xor U4684 (N_4684,N_4513,N_4582);
nand U4685 (N_4685,N_4591,N_4595);
xor U4686 (N_4686,N_4475,N_4497);
nand U4687 (N_4687,N_4568,N_4522);
and U4688 (N_4688,N_4427,N_4506);
or U4689 (N_4689,N_4444,N_4489);
or U4690 (N_4690,N_4525,N_4401);
and U4691 (N_4691,N_4500,N_4517);
and U4692 (N_4692,N_4415,N_4539);
nand U4693 (N_4693,N_4548,N_4526);
and U4694 (N_4694,N_4448,N_4487);
nand U4695 (N_4695,N_4423,N_4488);
nand U4696 (N_4696,N_4511,N_4466);
nor U4697 (N_4697,N_4533,N_4576);
or U4698 (N_4698,N_4419,N_4572);
and U4699 (N_4699,N_4581,N_4529);
and U4700 (N_4700,N_4579,N_4464);
nor U4701 (N_4701,N_4441,N_4545);
and U4702 (N_4702,N_4457,N_4439);
and U4703 (N_4703,N_4579,N_4571);
xnor U4704 (N_4704,N_4498,N_4444);
xnor U4705 (N_4705,N_4462,N_4527);
or U4706 (N_4706,N_4555,N_4407);
nor U4707 (N_4707,N_4414,N_4409);
and U4708 (N_4708,N_4571,N_4459);
nand U4709 (N_4709,N_4592,N_4489);
and U4710 (N_4710,N_4578,N_4423);
nor U4711 (N_4711,N_4431,N_4523);
nand U4712 (N_4712,N_4478,N_4564);
nor U4713 (N_4713,N_4437,N_4433);
xor U4714 (N_4714,N_4555,N_4557);
or U4715 (N_4715,N_4567,N_4418);
nor U4716 (N_4716,N_4477,N_4459);
xnor U4717 (N_4717,N_4428,N_4531);
xnor U4718 (N_4718,N_4585,N_4512);
and U4719 (N_4719,N_4571,N_4536);
or U4720 (N_4720,N_4511,N_4407);
nor U4721 (N_4721,N_4547,N_4574);
nand U4722 (N_4722,N_4598,N_4458);
nand U4723 (N_4723,N_4518,N_4542);
or U4724 (N_4724,N_4475,N_4523);
or U4725 (N_4725,N_4592,N_4408);
xor U4726 (N_4726,N_4403,N_4405);
or U4727 (N_4727,N_4565,N_4526);
nand U4728 (N_4728,N_4583,N_4432);
nand U4729 (N_4729,N_4579,N_4536);
or U4730 (N_4730,N_4449,N_4488);
nand U4731 (N_4731,N_4561,N_4589);
xor U4732 (N_4732,N_4505,N_4547);
nand U4733 (N_4733,N_4409,N_4503);
nand U4734 (N_4734,N_4466,N_4563);
nand U4735 (N_4735,N_4462,N_4480);
or U4736 (N_4736,N_4586,N_4477);
nor U4737 (N_4737,N_4560,N_4566);
nand U4738 (N_4738,N_4485,N_4586);
and U4739 (N_4739,N_4573,N_4555);
xnor U4740 (N_4740,N_4469,N_4439);
xor U4741 (N_4741,N_4449,N_4419);
nand U4742 (N_4742,N_4508,N_4438);
xnor U4743 (N_4743,N_4421,N_4501);
and U4744 (N_4744,N_4532,N_4503);
nor U4745 (N_4745,N_4584,N_4470);
xnor U4746 (N_4746,N_4477,N_4561);
nand U4747 (N_4747,N_4544,N_4598);
xor U4748 (N_4748,N_4578,N_4559);
nor U4749 (N_4749,N_4584,N_4453);
xnor U4750 (N_4750,N_4501,N_4544);
xor U4751 (N_4751,N_4470,N_4485);
nand U4752 (N_4752,N_4589,N_4526);
or U4753 (N_4753,N_4456,N_4547);
or U4754 (N_4754,N_4522,N_4564);
nand U4755 (N_4755,N_4469,N_4597);
or U4756 (N_4756,N_4439,N_4419);
nor U4757 (N_4757,N_4538,N_4588);
xnor U4758 (N_4758,N_4519,N_4484);
or U4759 (N_4759,N_4444,N_4561);
or U4760 (N_4760,N_4552,N_4514);
nor U4761 (N_4761,N_4530,N_4532);
nand U4762 (N_4762,N_4560,N_4421);
and U4763 (N_4763,N_4472,N_4467);
or U4764 (N_4764,N_4555,N_4454);
xnor U4765 (N_4765,N_4474,N_4440);
or U4766 (N_4766,N_4437,N_4413);
nand U4767 (N_4767,N_4576,N_4596);
or U4768 (N_4768,N_4474,N_4565);
nor U4769 (N_4769,N_4599,N_4487);
or U4770 (N_4770,N_4473,N_4407);
and U4771 (N_4771,N_4491,N_4451);
nor U4772 (N_4772,N_4436,N_4548);
nand U4773 (N_4773,N_4427,N_4569);
nor U4774 (N_4774,N_4409,N_4554);
and U4775 (N_4775,N_4414,N_4477);
nand U4776 (N_4776,N_4509,N_4428);
xor U4777 (N_4777,N_4580,N_4512);
nand U4778 (N_4778,N_4542,N_4423);
or U4779 (N_4779,N_4583,N_4510);
xor U4780 (N_4780,N_4512,N_4436);
nor U4781 (N_4781,N_4420,N_4444);
xnor U4782 (N_4782,N_4411,N_4564);
xor U4783 (N_4783,N_4582,N_4447);
and U4784 (N_4784,N_4584,N_4594);
or U4785 (N_4785,N_4480,N_4542);
or U4786 (N_4786,N_4588,N_4470);
xnor U4787 (N_4787,N_4552,N_4578);
and U4788 (N_4788,N_4520,N_4541);
xnor U4789 (N_4789,N_4585,N_4482);
nor U4790 (N_4790,N_4448,N_4413);
and U4791 (N_4791,N_4434,N_4573);
xnor U4792 (N_4792,N_4489,N_4521);
xor U4793 (N_4793,N_4471,N_4501);
nor U4794 (N_4794,N_4425,N_4540);
and U4795 (N_4795,N_4534,N_4580);
and U4796 (N_4796,N_4581,N_4580);
and U4797 (N_4797,N_4485,N_4557);
nand U4798 (N_4798,N_4464,N_4485);
and U4799 (N_4799,N_4432,N_4430);
and U4800 (N_4800,N_4780,N_4649);
and U4801 (N_4801,N_4746,N_4630);
or U4802 (N_4802,N_4617,N_4654);
nand U4803 (N_4803,N_4657,N_4639);
nor U4804 (N_4804,N_4619,N_4641);
or U4805 (N_4805,N_4632,N_4683);
xnor U4806 (N_4806,N_4756,N_4603);
nor U4807 (N_4807,N_4796,N_4627);
nor U4808 (N_4808,N_4610,N_4607);
or U4809 (N_4809,N_4682,N_4601);
or U4810 (N_4810,N_4661,N_4676);
or U4811 (N_4811,N_4737,N_4717);
xnor U4812 (N_4812,N_4602,N_4622);
nand U4813 (N_4813,N_4700,N_4776);
xor U4814 (N_4814,N_4604,N_4653);
nor U4815 (N_4815,N_4742,N_4624);
or U4816 (N_4816,N_4788,N_4696);
xnor U4817 (N_4817,N_4690,N_4795);
or U4818 (N_4818,N_4783,N_4763);
xnor U4819 (N_4819,N_4613,N_4723);
or U4820 (N_4820,N_4640,N_4659);
nand U4821 (N_4821,N_4773,N_4600);
nand U4822 (N_4822,N_4771,N_4638);
xor U4823 (N_4823,N_4710,N_4711);
nor U4824 (N_4824,N_4799,N_4626);
nor U4825 (N_4825,N_4618,N_4716);
and U4826 (N_4826,N_4736,N_4793);
or U4827 (N_4827,N_4655,N_4787);
nor U4828 (N_4828,N_4757,N_4731);
nor U4829 (N_4829,N_4652,N_4615);
nor U4830 (N_4830,N_4608,N_4688);
nor U4831 (N_4831,N_4747,N_4735);
and U4832 (N_4832,N_4645,N_4671);
nor U4833 (N_4833,N_4673,N_4754);
or U4834 (N_4834,N_4797,N_4663);
nor U4835 (N_4835,N_4621,N_4770);
or U4836 (N_4836,N_4666,N_4634);
xor U4837 (N_4837,N_4702,N_4753);
xnor U4838 (N_4838,N_4705,N_4628);
and U4839 (N_4839,N_4761,N_4719);
and U4840 (N_4840,N_4679,N_4740);
nand U4841 (N_4841,N_4733,N_4636);
and U4842 (N_4842,N_4744,N_4739);
nor U4843 (N_4843,N_4790,N_4693);
or U4844 (N_4844,N_4772,N_4726);
xnor U4845 (N_4845,N_4703,N_4779);
xnor U4846 (N_4846,N_4785,N_4662);
nand U4847 (N_4847,N_4701,N_4714);
xnor U4848 (N_4848,N_4758,N_4727);
nand U4849 (N_4849,N_4794,N_4750);
or U4850 (N_4850,N_4633,N_4698);
nand U4851 (N_4851,N_4620,N_4665);
or U4852 (N_4852,N_4791,N_4616);
and U4853 (N_4853,N_4730,N_4670);
nor U4854 (N_4854,N_4672,N_4721);
or U4855 (N_4855,N_4775,N_4781);
xor U4856 (N_4856,N_4692,N_4729);
nor U4857 (N_4857,N_4689,N_4715);
xnor U4858 (N_4858,N_4612,N_4678);
nor U4859 (N_4859,N_4675,N_4748);
and U4860 (N_4860,N_4647,N_4722);
nor U4861 (N_4861,N_4764,N_4668);
nor U4862 (N_4862,N_4743,N_4691);
nand U4863 (N_4863,N_4784,N_4642);
nand U4864 (N_4864,N_4686,N_4732);
or U4865 (N_4865,N_4725,N_4694);
nand U4866 (N_4866,N_4708,N_4681);
xnor U4867 (N_4867,N_4745,N_4786);
xor U4868 (N_4868,N_4765,N_4611);
nand U4869 (N_4869,N_4749,N_4774);
nand U4870 (N_4870,N_4685,N_4769);
nand U4871 (N_4871,N_4658,N_4656);
or U4872 (N_4872,N_4741,N_4789);
xnor U4873 (N_4873,N_4720,N_4635);
xor U4874 (N_4874,N_4629,N_4777);
and U4875 (N_4875,N_4631,N_4643);
nand U4876 (N_4876,N_4646,N_4759);
xor U4877 (N_4877,N_4724,N_4782);
nand U4878 (N_4878,N_4752,N_4792);
or U4879 (N_4879,N_4709,N_4718);
or U4880 (N_4880,N_4778,N_4664);
or U4881 (N_4881,N_4760,N_4684);
nor U4882 (N_4882,N_4614,N_4755);
or U4883 (N_4883,N_4674,N_4707);
or U4884 (N_4884,N_4625,N_4767);
nor U4885 (N_4885,N_4699,N_4704);
or U4886 (N_4886,N_4644,N_4606);
nor U4887 (N_4887,N_4766,N_4734);
xor U4888 (N_4888,N_4713,N_4712);
nor U4889 (N_4889,N_4697,N_4762);
nor U4890 (N_4890,N_4751,N_4623);
and U4891 (N_4891,N_4609,N_4738);
or U4892 (N_4892,N_4768,N_4728);
nor U4893 (N_4893,N_4637,N_4605);
nand U4894 (N_4894,N_4695,N_4706);
xnor U4895 (N_4895,N_4667,N_4680);
nor U4896 (N_4896,N_4651,N_4660);
nand U4897 (N_4897,N_4687,N_4669);
nand U4898 (N_4898,N_4677,N_4798);
nand U4899 (N_4899,N_4648,N_4650);
xnor U4900 (N_4900,N_4623,N_4664);
xor U4901 (N_4901,N_4765,N_4746);
nor U4902 (N_4902,N_4665,N_4763);
xnor U4903 (N_4903,N_4671,N_4776);
nor U4904 (N_4904,N_4797,N_4782);
nor U4905 (N_4905,N_4669,N_4709);
nand U4906 (N_4906,N_4780,N_4646);
nor U4907 (N_4907,N_4625,N_4781);
nor U4908 (N_4908,N_4651,N_4766);
or U4909 (N_4909,N_4629,N_4742);
nor U4910 (N_4910,N_4775,N_4766);
nand U4911 (N_4911,N_4724,N_4638);
and U4912 (N_4912,N_4703,N_4634);
xnor U4913 (N_4913,N_4682,N_4730);
nand U4914 (N_4914,N_4700,N_4610);
or U4915 (N_4915,N_4737,N_4742);
nand U4916 (N_4916,N_4795,N_4683);
and U4917 (N_4917,N_4706,N_4688);
or U4918 (N_4918,N_4664,N_4634);
xnor U4919 (N_4919,N_4636,N_4681);
nor U4920 (N_4920,N_4763,N_4648);
and U4921 (N_4921,N_4779,N_4611);
nor U4922 (N_4922,N_4616,N_4680);
or U4923 (N_4923,N_4611,N_4770);
xnor U4924 (N_4924,N_4716,N_4797);
nor U4925 (N_4925,N_4713,N_4663);
nor U4926 (N_4926,N_4675,N_4611);
or U4927 (N_4927,N_4767,N_4697);
xnor U4928 (N_4928,N_4623,N_4782);
xor U4929 (N_4929,N_4663,N_4795);
and U4930 (N_4930,N_4773,N_4621);
nand U4931 (N_4931,N_4661,N_4668);
and U4932 (N_4932,N_4750,N_4761);
or U4933 (N_4933,N_4680,N_4765);
or U4934 (N_4934,N_4708,N_4750);
or U4935 (N_4935,N_4634,N_4693);
or U4936 (N_4936,N_4740,N_4728);
and U4937 (N_4937,N_4702,N_4740);
xnor U4938 (N_4938,N_4670,N_4742);
nor U4939 (N_4939,N_4638,N_4661);
nor U4940 (N_4940,N_4773,N_4681);
nand U4941 (N_4941,N_4724,N_4654);
nand U4942 (N_4942,N_4602,N_4740);
xor U4943 (N_4943,N_4770,N_4736);
xnor U4944 (N_4944,N_4641,N_4707);
and U4945 (N_4945,N_4603,N_4671);
and U4946 (N_4946,N_4636,N_4774);
and U4947 (N_4947,N_4705,N_4745);
nand U4948 (N_4948,N_4757,N_4680);
xnor U4949 (N_4949,N_4741,N_4747);
and U4950 (N_4950,N_4610,N_4719);
nand U4951 (N_4951,N_4732,N_4619);
xnor U4952 (N_4952,N_4672,N_4631);
nor U4953 (N_4953,N_4681,N_4642);
and U4954 (N_4954,N_4629,N_4744);
nand U4955 (N_4955,N_4655,N_4642);
xor U4956 (N_4956,N_4625,N_4765);
nand U4957 (N_4957,N_4600,N_4691);
or U4958 (N_4958,N_4621,N_4789);
nor U4959 (N_4959,N_4762,N_4772);
xor U4960 (N_4960,N_4736,N_4686);
nand U4961 (N_4961,N_4778,N_4659);
xor U4962 (N_4962,N_4625,N_4621);
nor U4963 (N_4963,N_4728,N_4792);
or U4964 (N_4964,N_4730,N_4643);
xor U4965 (N_4965,N_4750,N_4649);
and U4966 (N_4966,N_4797,N_4724);
or U4967 (N_4967,N_4661,N_4658);
or U4968 (N_4968,N_4651,N_4600);
and U4969 (N_4969,N_4607,N_4617);
nor U4970 (N_4970,N_4771,N_4604);
and U4971 (N_4971,N_4797,N_4722);
or U4972 (N_4972,N_4636,N_4736);
xnor U4973 (N_4973,N_4601,N_4616);
nand U4974 (N_4974,N_4633,N_4744);
and U4975 (N_4975,N_4764,N_4650);
nand U4976 (N_4976,N_4724,N_4747);
or U4977 (N_4977,N_4785,N_4722);
xnor U4978 (N_4978,N_4704,N_4721);
nor U4979 (N_4979,N_4761,N_4672);
and U4980 (N_4980,N_4702,N_4778);
nor U4981 (N_4981,N_4783,N_4655);
and U4982 (N_4982,N_4704,N_4720);
xnor U4983 (N_4983,N_4634,N_4769);
nand U4984 (N_4984,N_4742,N_4617);
nand U4985 (N_4985,N_4785,N_4608);
xnor U4986 (N_4986,N_4768,N_4629);
and U4987 (N_4987,N_4631,N_4696);
or U4988 (N_4988,N_4621,N_4642);
and U4989 (N_4989,N_4742,N_4730);
xor U4990 (N_4990,N_4709,N_4771);
xnor U4991 (N_4991,N_4691,N_4667);
or U4992 (N_4992,N_4633,N_4717);
nor U4993 (N_4993,N_4745,N_4690);
and U4994 (N_4994,N_4759,N_4710);
and U4995 (N_4995,N_4617,N_4761);
and U4996 (N_4996,N_4694,N_4709);
nor U4997 (N_4997,N_4754,N_4791);
nand U4998 (N_4998,N_4763,N_4650);
xnor U4999 (N_4999,N_4653,N_4767);
nor U5000 (N_5000,N_4925,N_4956);
nand U5001 (N_5001,N_4823,N_4931);
nor U5002 (N_5002,N_4876,N_4829);
nor U5003 (N_5003,N_4968,N_4949);
nor U5004 (N_5004,N_4984,N_4918);
xor U5005 (N_5005,N_4962,N_4814);
nand U5006 (N_5006,N_4980,N_4878);
nor U5007 (N_5007,N_4974,N_4977);
xnor U5008 (N_5008,N_4887,N_4946);
nor U5009 (N_5009,N_4948,N_4899);
or U5010 (N_5010,N_4831,N_4819);
nand U5011 (N_5011,N_4882,N_4902);
xnor U5012 (N_5012,N_4842,N_4989);
and U5013 (N_5013,N_4896,N_4843);
nand U5014 (N_5014,N_4802,N_4862);
nand U5015 (N_5015,N_4839,N_4860);
nor U5016 (N_5016,N_4930,N_4990);
nor U5017 (N_5017,N_4986,N_4967);
or U5018 (N_5018,N_4982,N_4915);
and U5019 (N_5019,N_4816,N_4972);
xor U5020 (N_5020,N_4957,N_4863);
or U5021 (N_5021,N_4805,N_4922);
xor U5022 (N_5022,N_4952,N_4826);
xor U5023 (N_5023,N_4848,N_4824);
and U5024 (N_5024,N_4847,N_4870);
and U5025 (N_5025,N_4961,N_4813);
nand U5026 (N_5026,N_4940,N_4886);
nand U5027 (N_5027,N_4893,N_4871);
xnor U5028 (N_5028,N_4992,N_4907);
xor U5029 (N_5029,N_4912,N_4937);
xnor U5030 (N_5030,N_4801,N_4945);
or U5031 (N_5031,N_4923,N_4810);
nor U5032 (N_5032,N_4869,N_4865);
or U5033 (N_5033,N_4854,N_4808);
nand U5034 (N_5034,N_4935,N_4856);
nand U5035 (N_5035,N_4908,N_4951);
nand U5036 (N_5036,N_4881,N_4909);
nor U5037 (N_5037,N_4874,N_4832);
or U5038 (N_5038,N_4944,N_4913);
xor U5039 (N_5039,N_4890,N_4966);
or U5040 (N_5040,N_4836,N_4894);
nand U5041 (N_5041,N_4807,N_4970);
and U5042 (N_5042,N_4845,N_4861);
xnor U5043 (N_5043,N_4818,N_4809);
or U5044 (N_5044,N_4994,N_4963);
xor U5045 (N_5045,N_4958,N_4934);
and U5046 (N_5046,N_4924,N_4891);
xor U5047 (N_5047,N_4892,N_4927);
nor U5048 (N_5048,N_4827,N_4837);
nand U5049 (N_5049,N_4953,N_4914);
xnor U5050 (N_5050,N_4866,N_4910);
or U5051 (N_5051,N_4825,N_4985);
and U5052 (N_5052,N_4959,N_4853);
or U5053 (N_5053,N_4841,N_4997);
xor U5054 (N_5054,N_4857,N_4975);
nand U5055 (N_5055,N_4875,N_4916);
and U5056 (N_5056,N_4877,N_4901);
and U5057 (N_5057,N_4898,N_4955);
and U5058 (N_5058,N_4942,N_4999);
xor U5059 (N_5059,N_4996,N_4904);
nor U5060 (N_5060,N_4821,N_4838);
or U5061 (N_5061,N_4965,N_4833);
nor U5062 (N_5062,N_4976,N_4888);
nand U5063 (N_5063,N_4903,N_4979);
and U5064 (N_5064,N_4828,N_4983);
nand U5065 (N_5065,N_4921,N_4905);
nand U5066 (N_5066,N_4993,N_4803);
nor U5067 (N_5067,N_4830,N_4969);
xnor U5068 (N_5068,N_4895,N_4806);
and U5069 (N_5069,N_4954,N_4947);
or U5070 (N_5070,N_4868,N_4987);
nor U5071 (N_5071,N_4858,N_4851);
nand U5072 (N_5072,N_4919,N_4822);
xnor U5073 (N_5073,N_4900,N_4846);
xnor U5074 (N_5074,N_4800,N_4812);
nor U5075 (N_5075,N_4995,N_4873);
xor U5076 (N_5076,N_4815,N_4883);
xor U5077 (N_5077,N_4804,N_4835);
xnor U5078 (N_5078,N_4840,N_4981);
or U5079 (N_5079,N_4911,N_4817);
xor U5080 (N_5080,N_4906,N_4932);
and U5081 (N_5081,N_4964,N_4943);
nand U5082 (N_5082,N_4897,N_4973);
nor U5083 (N_5083,N_4889,N_4917);
or U5084 (N_5084,N_4926,N_4879);
and U5085 (N_5085,N_4885,N_4933);
and U5086 (N_5086,N_4920,N_4939);
or U5087 (N_5087,N_4880,N_4864);
or U5088 (N_5088,N_4991,N_4811);
or U5089 (N_5089,N_4941,N_4850);
nand U5090 (N_5090,N_4820,N_4971);
nand U5091 (N_5091,N_4928,N_4849);
and U5092 (N_5092,N_4936,N_4844);
and U5093 (N_5093,N_4859,N_4872);
nor U5094 (N_5094,N_4998,N_4960);
xnor U5095 (N_5095,N_4938,N_4834);
xor U5096 (N_5096,N_4852,N_4867);
nand U5097 (N_5097,N_4855,N_4950);
nand U5098 (N_5098,N_4988,N_4884);
nor U5099 (N_5099,N_4978,N_4929);
and U5100 (N_5100,N_4969,N_4936);
and U5101 (N_5101,N_4949,N_4981);
or U5102 (N_5102,N_4805,N_4923);
nor U5103 (N_5103,N_4982,N_4867);
and U5104 (N_5104,N_4887,N_4917);
xor U5105 (N_5105,N_4880,N_4997);
nor U5106 (N_5106,N_4915,N_4994);
nor U5107 (N_5107,N_4953,N_4969);
or U5108 (N_5108,N_4841,N_4891);
and U5109 (N_5109,N_4898,N_4862);
or U5110 (N_5110,N_4820,N_4981);
xnor U5111 (N_5111,N_4907,N_4819);
or U5112 (N_5112,N_4978,N_4883);
xor U5113 (N_5113,N_4925,N_4919);
or U5114 (N_5114,N_4815,N_4814);
nor U5115 (N_5115,N_4976,N_4951);
xnor U5116 (N_5116,N_4873,N_4920);
nor U5117 (N_5117,N_4836,N_4807);
or U5118 (N_5118,N_4808,N_4825);
xnor U5119 (N_5119,N_4827,N_4875);
nor U5120 (N_5120,N_4813,N_4912);
nand U5121 (N_5121,N_4873,N_4950);
nor U5122 (N_5122,N_4914,N_4823);
nor U5123 (N_5123,N_4849,N_4979);
xor U5124 (N_5124,N_4817,N_4866);
nand U5125 (N_5125,N_4919,N_4968);
nand U5126 (N_5126,N_4813,N_4874);
xnor U5127 (N_5127,N_4872,N_4850);
nor U5128 (N_5128,N_4852,N_4822);
xnor U5129 (N_5129,N_4886,N_4881);
xor U5130 (N_5130,N_4966,N_4967);
or U5131 (N_5131,N_4827,N_4864);
or U5132 (N_5132,N_4945,N_4880);
nor U5133 (N_5133,N_4907,N_4997);
xnor U5134 (N_5134,N_4854,N_4912);
nand U5135 (N_5135,N_4881,N_4998);
and U5136 (N_5136,N_4924,N_4861);
xor U5137 (N_5137,N_4991,N_4823);
or U5138 (N_5138,N_4879,N_4831);
nor U5139 (N_5139,N_4858,N_4906);
xnor U5140 (N_5140,N_4856,N_4803);
xnor U5141 (N_5141,N_4993,N_4973);
nand U5142 (N_5142,N_4919,N_4909);
or U5143 (N_5143,N_4922,N_4873);
nand U5144 (N_5144,N_4981,N_4992);
nor U5145 (N_5145,N_4990,N_4801);
nand U5146 (N_5146,N_4930,N_4977);
or U5147 (N_5147,N_4837,N_4939);
or U5148 (N_5148,N_4851,N_4884);
or U5149 (N_5149,N_4899,N_4816);
nor U5150 (N_5150,N_4823,N_4840);
or U5151 (N_5151,N_4937,N_4884);
nand U5152 (N_5152,N_4906,N_4976);
or U5153 (N_5153,N_4884,N_4904);
and U5154 (N_5154,N_4804,N_4851);
nor U5155 (N_5155,N_4924,N_4906);
nand U5156 (N_5156,N_4848,N_4953);
nand U5157 (N_5157,N_4836,N_4993);
nand U5158 (N_5158,N_4935,N_4834);
or U5159 (N_5159,N_4806,N_4944);
nor U5160 (N_5160,N_4971,N_4816);
and U5161 (N_5161,N_4892,N_4885);
xor U5162 (N_5162,N_4823,N_4888);
xor U5163 (N_5163,N_4816,N_4946);
or U5164 (N_5164,N_4941,N_4947);
or U5165 (N_5165,N_4884,N_4845);
or U5166 (N_5166,N_4808,N_4994);
or U5167 (N_5167,N_4807,N_4856);
or U5168 (N_5168,N_4986,N_4821);
xor U5169 (N_5169,N_4839,N_4952);
nand U5170 (N_5170,N_4889,N_4804);
or U5171 (N_5171,N_4960,N_4869);
or U5172 (N_5172,N_4896,N_4880);
nand U5173 (N_5173,N_4958,N_4920);
nor U5174 (N_5174,N_4886,N_4802);
and U5175 (N_5175,N_4879,N_4989);
xor U5176 (N_5176,N_4984,N_4956);
xor U5177 (N_5177,N_4820,N_4968);
nand U5178 (N_5178,N_4917,N_4822);
and U5179 (N_5179,N_4941,N_4992);
nand U5180 (N_5180,N_4919,N_4841);
xnor U5181 (N_5181,N_4948,N_4962);
nand U5182 (N_5182,N_4826,N_4951);
nor U5183 (N_5183,N_4802,N_4923);
and U5184 (N_5184,N_4807,N_4942);
or U5185 (N_5185,N_4919,N_4949);
nand U5186 (N_5186,N_4800,N_4831);
nor U5187 (N_5187,N_4970,N_4876);
nand U5188 (N_5188,N_4851,N_4912);
nand U5189 (N_5189,N_4954,N_4822);
or U5190 (N_5190,N_4966,N_4935);
xnor U5191 (N_5191,N_4979,N_4932);
xor U5192 (N_5192,N_4890,N_4837);
nor U5193 (N_5193,N_4876,N_4891);
nor U5194 (N_5194,N_4926,N_4803);
nor U5195 (N_5195,N_4930,N_4874);
nor U5196 (N_5196,N_4893,N_4948);
nor U5197 (N_5197,N_4868,N_4870);
nand U5198 (N_5198,N_4811,N_4943);
xnor U5199 (N_5199,N_4876,N_4802);
xnor U5200 (N_5200,N_5186,N_5113);
and U5201 (N_5201,N_5046,N_5188);
and U5202 (N_5202,N_5061,N_5037);
xor U5203 (N_5203,N_5114,N_5051);
nor U5204 (N_5204,N_5162,N_5116);
or U5205 (N_5205,N_5104,N_5137);
xnor U5206 (N_5206,N_5183,N_5055);
nor U5207 (N_5207,N_5194,N_5014);
or U5208 (N_5208,N_5089,N_5050);
nor U5209 (N_5209,N_5158,N_5086);
or U5210 (N_5210,N_5049,N_5005);
nor U5211 (N_5211,N_5144,N_5142);
xor U5212 (N_5212,N_5063,N_5112);
nand U5213 (N_5213,N_5131,N_5146);
nor U5214 (N_5214,N_5066,N_5048);
nor U5215 (N_5215,N_5199,N_5011);
or U5216 (N_5216,N_5178,N_5039);
or U5217 (N_5217,N_5175,N_5052);
xnor U5218 (N_5218,N_5187,N_5138);
and U5219 (N_5219,N_5090,N_5099);
and U5220 (N_5220,N_5134,N_5191);
and U5221 (N_5221,N_5044,N_5043);
nand U5222 (N_5222,N_5076,N_5130);
or U5223 (N_5223,N_5079,N_5125);
xor U5224 (N_5224,N_5070,N_5082);
or U5225 (N_5225,N_5108,N_5163);
nor U5226 (N_5226,N_5042,N_5150);
xor U5227 (N_5227,N_5083,N_5197);
nor U5228 (N_5228,N_5006,N_5028);
or U5229 (N_5229,N_5034,N_5075);
xnor U5230 (N_5230,N_5153,N_5102);
nand U5231 (N_5231,N_5151,N_5120);
and U5232 (N_5232,N_5007,N_5156);
nor U5233 (N_5233,N_5110,N_5121);
nor U5234 (N_5234,N_5073,N_5000);
xor U5235 (N_5235,N_5016,N_5184);
nand U5236 (N_5236,N_5004,N_5025);
and U5237 (N_5237,N_5088,N_5077);
nand U5238 (N_5238,N_5038,N_5032);
xor U5239 (N_5239,N_5103,N_5094);
nor U5240 (N_5240,N_5035,N_5095);
xor U5241 (N_5241,N_5129,N_5020);
and U5242 (N_5242,N_5115,N_5097);
nor U5243 (N_5243,N_5109,N_5118);
nand U5244 (N_5244,N_5068,N_5133);
xnor U5245 (N_5245,N_5045,N_5054);
nand U5246 (N_5246,N_5023,N_5193);
nor U5247 (N_5247,N_5056,N_5093);
or U5248 (N_5248,N_5064,N_5026);
xnor U5249 (N_5249,N_5182,N_5124);
and U5250 (N_5250,N_5015,N_5096);
or U5251 (N_5251,N_5003,N_5018);
nand U5252 (N_5252,N_5053,N_5081);
or U5253 (N_5253,N_5008,N_5195);
and U5254 (N_5254,N_5069,N_5179);
and U5255 (N_5255,N_5084,N_5117);
and U5256 (N_5256,N_5141,N_5196);
xor U5257 (N_5257,N_5128,N_5027);
nand U5258 (N_5258,N_5165,N_5019);
nor U5259 (N_5259,N_5148,N_5009);
nor U5260 (N_5260,N_5161,N_5181);
xnor U5261 (N_5261,N_5135,N_5145);
or U5262 (N_5262,N_5036,N_5013);
xor U5263 (N_5263,N_5157,N_5170);
xnor U5264 (N_5264,N_5127,N_5155);
and U5265 (N_5265,N_5167,N_5171);
nor U5266 (N_5266,N_5085,N_5098);
or U5267 (N_5267,N_5074,N_5172);
nor U5268 (N_5268,N_5149,N_5072);
or U5269 (N_5269,N_5143,N_5198);
and U5270 (N_5270,N_5107,N_5101);
nand U5271 (N_5271,N_5062,N_5185);
nand U5272 (N_5272,N_5078,N_5060);
nor U5273 (N_5273,N_5106,N_5168);
xor U5274 (N_5274,N_5057,N_5017);
nor U5275 (N_5275,N_5091,N_5040);
nand U5276 (N_5276,N_5126,N_5164);
and U5277 (N_5277,N_5010,N_5058);
xor U5278 (N_5278,N_5029,N_5136);
nand U5279 (N_5279,N_5002,N_5100);
xor U5280 (N_5280,N_5024,N_5123);
nand U5281 (N_5281,N_5047,N_5067);
xor U5282 (N_5282,N_5152,N_5166);
nand U5283 (N_5283,N_5159,N_5176);
or U5284 (N_5284,N_5190,N_5147);
xor U5285 (N_5285,N_5041,N_5174);
xor U5286 (N_5286,N_5105,N_5012);
and U5287 (N_5287,N_5160,N_5173);
xnor U5288 (N_5288,N_5119,N_5031);
xor U5289 (N_5289,N_5140,N_5154);
and U5290 (N_5290,N_5071,N_5033);
nand U5291 (N_5291,N_5111,N_5080);
or U5292 (N_5292,N_5001,N_5189);
and U5293 (N_5293,N_5021,N_5030);
or U5294 (N_5294,N_5180,N_5132);
and U5295 (N_5295,N_5139,N_5022);
xnor U5296 (N_5296,N_5192,N_5092);
or U5297 (N_5297,N_5122,N_5177);
or U5298 (N_5298,N_5065,N_5169);
or U5299 (N_5299,N_5059,N_5087);
or U5300 (N_5300,N_5193,N_5003);
and U5301 (N_5301,N_5163,N_5038);
nor U5302 (N_5302,N_5009,N_5006);
and U5303 (N_5303,N_5102,N_5061);
nor U5304 (N_5304,N_5094,N_5049);
or U5305 (N_5305,N_5036,N_5153);
xnor U5306 (N_5306,N_5195,N_5095);
and U5307 (N_5307,N_5030,N_5159);
nand U5308 (N_5308,N_5047,N_5107);
or U5309 (N_5309,N_5035,N_5123);
nor U5310 (N_5310,N_5091,N_5059);
xor U5311 (N_5311,N_5051,N_5055);
nor U5312 (N_5312,N_5040,N_5194);
or U5313 (N_5313,N_5106,N_5163);
or U5314 (N_5314,N_5136,N_5014);
or U5315 (N_5315,N_5006,N_5074);
nor U5316 (N_5316,N_5142,N_5174);
xnor U5317 (N_5317,N_5050,N_5020);
and U5318 (N_5318,N_5152,N_5073);
nand U5319 (N_5319,N_5084,N_5072);
or U5320 (N_5320,N_5051,N_5113);
and U5321 (N_5321,N_5192,N_5088);
or U5322 (N_5322,N_5069,N_5064);
and U5323 (N_5323,N_5094,N_5077);
nor U5324 (N_5324,N_5128,N_5106);
and U5325 (N_5325,N_5017,N_5034);
xnor U5326 (N_5326,N_5187,N_5156);
or U5327 (N_5327,N_5103,N_5033);
xor U5328 (N_5328,N_5166,N_5154);
nand U5329 (N_5329,N_5172,N_5031);
or U5330 (N_5330,N_5067,N_5134);
nor U5331 (N_5331,N_5114,N_5039);
xnor U5332 (N_5332,N_5097,N_5085);
nand U5333 (N_5333,N_5023,N_5171);
xor U5334 (N_5334,N_5017,N_5152);
and U5335 (N_5335,N_5010,N_5033);
nor U5336 (N_5336,N_5115,N_5045);
xor U5337 (N_5337,N_5168,N_5038);
and U5338 (N_5338,N_5180,N_5131);
or U5339 (N_5339,N_5130,N_5096);
nor U5340 (N_5340,N_5001,N_5085);
nor U5341 (N_5341,N_5119,N_5052);
xor U5342 (N_5342,N_5038,N_5056);
xor U5343 (N_5343,N_5168,N_5022);
xor U5344 (N_5344,N_5056,N_5186);
or U5345 (N_5345,N_5116,N_5040);
nor U5346 (N_5346,N_5011,N_5197);
and U5347 (N_5347,N_5009,N_5158);
or U5348 (N_5348,N_5049,N_5084);
or U5349 (N_5349,N_5151,N_5137);
or U5350 (N_5350,N_5032,N_5103);
and U5351 (N_5351,N_5080,N_5160);
and U5352 (N_5352,N_5080,N_5060);
nand U5353 (N_5353,N_5157,N_5115);
nand U5354 (N_5354,N_5154,N_5090);
nor U5355 (N_5355,N_5014,N_5106);
or U5356 (N_5356,N_5167,N_5050);
nor U5357 (N_5357,N_5083,N_5089);
nor U5358 (N_5358,N_5049,N_5001);
and U5359 (N_5359,N_5013,N_5073);
and U5360 (N_5360,N_5088,N_5008);
nor U5361 (N_5361,N_5199,N_5104);
or U5362 (N_5362,N_5012,N_5024);
or U5363 (N_5363,N_5109,N_5155);
and U5364 (N_5364,N_5136,N_5051);
and U5365 (N_5365,N_5193,N_5108);
and U5366 (N_5366,N_5111,N_5105);
xor U5367 (N_5367,N_5159,N_5081);
xnor U5368 (N_5368,N_5086,N_5032);
xnor U5369 (N_5369,N_5087,N_5029);
xnor U5370 (N_5370,N_5023,N_5072);
xnor U5371 (N_5371,N_5110,N_5050);
nor U5372 (N_5372,N_5047,N_5122);
xnor U5373 (N_5373,N_5137,N_5165);
xor U5374 (N_5374,N_5194,N_5156);
or U5375 (N_5375,N_5152,N_5095);
nand U5376 (N_5376,N_5105,N_5078);
or U5377 (N_5377,N_5072,N_5073);
nand U5378 (N_5378,N_5085,N_5179);
and U5379 (N_5379,N_5089,N_5053);
and U5380 (N_5380,N_5024,N_5131);
xnor U5381 (N_5381,N_5009,N_5077);
nand U5382 (N_5382,N_5161,N_5017);
nor U5383 (N_5383,N_5161,N_5120);
or U5384 (N_5384,N_5109,N_5170);
nand U5385 (N_5385,N_5071,N_5160);
nor U5386 (N_5386,N_5100,N_5007);
and U5387 (N_5387,N_5116,N_5100);
and U5388 (N_5388,N_5060,N_5097);
nand U5389 (N_5389,N_5170,N_5185);
nor U5390 (N_5390,N_5061,N_5165);
nor U5391 (N_5391,N_5154,N_5035);
or U5392 (N_5392,N_5157,N_5074);
nor U5393 (N_5393,N_5155,N_5183);
nor U5394 (N_5394,N_5196,N_5192);
nand U5395 (N_5395,N_5033,N_5098);
and U5396 (N_5396,N_5163,N_5056);
and U5397 (N_5397,N_5171,N_5009);
or U5398 (N_5398,N_5136,N_5141);
and U5399 (N_5399,N_5174,N_5054);
or U5400 (N_5400,N_5268,N_5265);
xnor U5401 (N_5401,N_5295,N_5312);
nor U5402 (N_5402,N_5306,N_5207);
and U5403 (N_5403,N_5227,N_5240);
and U5404 (N_5404,N_5392,N_5230);
and U5405 (N_5405,N_5283,N_5334);
and U5406 (N_5406,N_5250,N_5277);
and U5407 (N_5407,N_5260,N_5378);
or U5408 (N_5408,N_5363,N_5318);
nand U5409 (N_5409,N_5337,N_5221);
xnor U5410 (N_5410,N_5242,N_5220);
nand U5411 (N_5411,N_5259,N_5310);
nor U5412 (N_5412,N_5302,N_5369);
or U5413 (N_5413,N_5288,N_5313);
or U5414 (N_5414,N_5280,N_5261);
or U5415 (N_5415,N_5203,N_5211);
nand U5416 (N_5416,N_5238,N_5380);
nand U5417 (N_5417,N_5370,N_5274);
nor U5418 (N_5418,N_5309,N_5388);
or U5419 (N_5419,N_5285,N_5258);
or U5420 (N_5420,N_5225,N_5212);
xor U5421 (N_5421,N_5264,N_5224);
or U5422 (N_5422,N_5291,N_5299);
xnor U5423 (N_5423,N_5209,N_5279);
nor U5424 (N_5424,N_5353,N_5335);
nand U5425 (N_5425,N_5204,N_5373);
nand U5426 (N_5426,N_5216,N_5282);
nand U5427 (N_5427,N_5348,N_5367);
nand U5428 (N_5428,N_5303,N_5322);
and U5429 (N_5429,N_5248,N_5243);
and U5430 (N_5430,N_5390,N_5394);
or U5431 (N_5431,N_5293,N_5254);
or U5432 (N_5432,N_5346,N_5389);
and U5433 (N_5433,N_5201,N_5397);
or U5434 (N_5434,N_5252,N_5287);
nor U5435 (N_5435,N_5251,N_5368);
xnor U5436 (N_5436,N_5253,N_5358);
xnor U5437 (N_5437,N_5231,N_5338);
or U5438 (N_5438,N_5342,N_5266);
or U5439 (N_5439,N_5304,N_5355);
and U5440 (N_5440,N_5239,N_5255);
nor U5441 (N_5441,N_5256,N_5249);
and U5442 (N_5442,N_5272,N_5343);
nor U5443 (N_5443,N_5215,N_5233);
nand U5444 (N_5444,N_5317,N_5321);
and U5445 (N_5445,N_5381,N_5340);
and U5446 (N_5446,N_5314,N_5360);
nand U5447 (N_5447,N_5396,N_5359);
xor U5448 (N_5448,N_5226,N_5361);
and U5449 (N_5449,N_5289,N_5270);
xor U5450 (N_5450,N_5333,N_5329);
and U5451 (N_5451,N_5382,N_5281);
nor U5452 (N_5452,N_5214,N_5349);
or U5453 (N_5453,N_5323,N_5324);
or U5454 (N_5454,N_5296,N_5362);
xor U5455 (N_5455,N_5327,N_5300);
nor U5456 (N_5456,N_5395,N_5365);
xor U5457 (N_5457,N_5237,N_5357);
or U5458 (N_5458,N_5319,N_5352);
or U5459 (N_5459,N_5244,N_5301);
or U5460 (N_5460,N_5391,N_5377);
xor U5461 (N_5461,N_5372,N_5305);
or U5462 (N_5462,N_5200,N_5241);
nor U5463 (N_5463,N_5217,N_5383);
or U5464 (N_5464,N_5278,N_5234);
or U5465 (N_5465,N_5292,N_5315);
xor U5466 (N_5466,N_5245,N_5236);
and U5467 (N_5467,N_5208,N_5222);
xnor U5468 (N_5468,N_5386,N_5320);
or U5469 (N_5469,N_5276,N_5262);
or U5470 (N_5470,N_5247,N_5284);
or U5471 (N_5471,N_5311,N_5206);
xor U5472 (N_5472,N_5347,N_5316);
and U5473 (N_5473,N_5351,N_5375);
and U5474 (N_5474,N_5356,N_5218);
xnor U5475 (N_5475,N_5232,N_5345);
or U5476 (N_5476,N_5366,N_5275);
and U5477 (N_5477,N_5325,N_5205);
or U5478 (N_5478,N_5399,N_5269);
nand U5479 (N_5479,N_5393,N_5344);
xnor U5480 (N_5480,N_5297,N_5398);
and U5481 (N_5481,N_5213,N_5364);
xnor U5482 (N_5482,N_5219,N_5331);
nor U5483 (N_5483,N_5371,N_5350);
nand U5484 (N_5484,N_5290,N_5235);
nand U5485 (N_5485,N_5326,N_5379);
nor U5486 (N_5486,N_5229,N_5228);
or U5487 (N_5487,N_5271,N_5330);
nor U5488 (N_5488,N_5257,N_5286);
and U5489 (N_5489,N_5341,N_5308);
nor U5490 (N_5490,N_5298,N_5202);
and U5491 (N_5491,N_5273,N_5294);
nand U5492 (N_5492,N_5263,N_5223);
nand U5493 (N_5493,N_5332,N_5376);
or U5494 (N_5494,N_5374,N_5267);
or U5495 (N_5495,N_5384,N_5328);
nand U5496 (N_5496,N_5246,N_5339);
and U5497 (N_5497,N_5307,N_5336);
or U5498 (N_5498,N_5210,N_5354);
xor U5499 (N_5499,N_5385,N_5387);
nor U5500 (N_5500,N_5220,N_5329);
nor U5501 (N_5501,N_5220,N_5374);
or U5502 (N_5502,N_5278,N_5384);
nor U5503 (N_5503,N_5207,N_5228);
nand U5504 (N_5504,N_5218,N_5361);
or U5505 (N_5505,N_5282,N_5265);
nand U5506 (N_5506,N_5379,N_5397);
or U5507 (N_5507,N_5351,N_5394);
or U5508 (N_5508,N_5276,N_5317);
and U5509 (N_5509,N_5340,N_5224);
nor U5510 (N_5510,N_5209,N_5313);
and U5511 (N_5511,N_5379,N_5200);
and U5512 (N_5512,N_5346,N_5256);
or U5513 (N_5513,N_5338,N_5334);
nand U5514 (N_5514,N_5287,N_5283);
and U5515 (N_5515,N_5396,N_5360);
nand U5516 (N_5516,N_5321,N_5268);
or U5517 (N_5517,N_5232,N_5250);
nor U5518 (N_5518,N_5395,N_5309);
or U5519 (N_5519,N_5374,N_5262);
or U5520 (N_5520,N_5221,N_5324);
xnor U5521 (N_5521,N_5284,N_5326);
or U5522 (N_5522,N_5345,N_5312);
nor U5523 (N_5523,N_5347,N_5372);
xnor U5524 (N_5524,N_5278,N_5213);
xnor U5525 (N_5525,N_5350,N_5256);
or U5526 (N_5526,N_5302,N_5266);
xnor U5527 (N_5527,N_5344,N_5362);
or U5528 (N_5528,N_5391,N_5278);
nor U5529 (N_5529,N_5260,N_5387);
xor U5530 (N_5530,N_5280,N_5312);
xor U5531 (N_5531,N_5204,N_5396);
xnor U5532 (N_5532,N_5254,N_5362);
nor U5533 (N_5533,N_5374,N_5223);
or U5534 (N_5534,N_5298,N_5338);
or U5535 (N_5535,N_5200,N_5288);
nand U5536 (N_5536,N_5375,N_5276);
xnor U5537 (N_5537,N_5320,N_5247);
nand U5538 (N_5538,N_5300,N_5368);
xor U5539 (N_5539,N_5302,N_5236);
nor U5540 (N_5540,N_5342,N_5382);
nor U5541 (N_5541,N_5288,N_5368);
nor U5542 (N_5542,N_5358,N_5365);
or U5543 (N_5543,N_5395,N_5331);
and U5544 (N_5544,N_5280,N_5203);
nand U5545 (N_5545,N_5312,N_5390);
nand U5546 (N_5546,N_5369,N_5220);
xnor U5547 (N_5547,N_5288,N_5260);
nor U5548 (N_5548,N_5271,N_5257);
xnor U5549 (N_5549,N_5355,N_5358);
nor U5550 (N_5550,N_5244,N_5262);
nor U5551 (N_5551,N_5381,N_5254);
nor U5552 (N_5552,N_5277,N_5247);
or U5553 (N_5553,N_5286,N_5265);
or U5554 (N_5554,N_5316,N_5257);
or U5555 (N_5555,N_5372,N_5217);
nand U5556 (N_5556,N_5327,N_5274);
and U5557 (N_5557,N_5394,N_5300);
and U5558 (N_5558,N_5241,N_5283);
nand U5559 (N_5559,N_5295,N_5210);
xor U5560 (N_5560,N_5254,N_5251);
or U5561 (N_5561,N_5227,N_5371);
and U5562 (N_5562,N_5243,N_5326);
or U5563 (N_5563,N_5273,N_5386);
nand U5564 (N_5564,N_5324,N_5395);
xor U5565 (N_5565,N_5213,N_5384);
or U5566 (N_5566,N_5209,N_5308);
xnor U5567 (N_5567,N_5215,N_5263);
and U5568 (N_5568,N_5221,N_5298);
nand U5569 (N_5569,N_5358,N_5371);
xor U5570 (N_5570,N_5328,N_5367);
xor U5571 (N_5571,N_5339,N_5263);
nor U5572 (N_5572,N_5223,N_5308);
nor U5573 (N_5573,N_5273,N_5359);
nor U5574 (N_5574,N_5332,N_5205);
xnor U5575 (N_5575,N_5252,N_5224);
or U5576 (N_5576,N_5329,N_5308);
or U5577 (N_5577,N_5235,N_5212);
or U5578 (N_5578,N_5397,N_5303);
nand U5579 (N_5579,N_5368,N_5265);
nor U5580 (N_5580,N_5392,N_5357);
xnor U5581 (N_5581,N_5383,N_5241);
or U5582 (N_5582,N_5293,N_5317);
nand U5583 (N_5583,N_5242,N_5376);
or U5584 (N_5584,N_5340,N_5294);
nand U5585 (N_5585,N_5281,N_5296);
xor U5586 (N_5586,N_5203,N_5337);
and U5587 (N_5587,N_5386,N_5237);
and U5588 (N_5588,N_5303,N_5242);
nor U5589 (N_5589,N_5243,N_5335);
and U5590 (N_5590,N_5214,N_5261);
xor U5591 (N_5591,N_5208,N_5394);
xnor U5592 (N_5592,N_5260,N_5208);
nor U5593 (N_5593,N_5329,N_5263);
or U5594 (N_5594,N_5265,N_5245);
or U5595 (N_5595,N_5208,N_5387);
nor U5596 (N_5596,N_5398,N_5321);
xor U5597 (N_5597,N_5263,N_5290);
and U5598 (N_5598,N_5383,N_5243);
and U5599 (N_5599,N_5201,N_5344);
and U5600 (N_5600,N_5548,N_5407);
nand U5601 (N_5601,N_5557,N_5406);
and U5602 (N_5602,N_5504,N_5487);
or U5603 (N_5603,N_5498,N_5518);
and U5604 (N_5604,N_5490,N_5563);
nor U5605 (N_5605,N_5560,N_5484);
and U5606 (N_5606,N_5467,N_5497);
nor U5607 (N_5607,N_5469,N_5567);
xor U5608 (N_5608,N_5551,N_5447);
and U5609 (N_5609,N_5438,N_5522);
or U5610 (N_5610,N_5499,N_5482);
xnor U5611 (N_5611,N_5565,N_5587);
and U5612 (N_5612,N_5411,N_5479);
nand U5613 (N_5613,N_5480,N_5453);
nor U5614 (N_5614,N_5478,N_5405);
xnor U5615 (N_5615,N_5568,N_5594);
nand U5616 (N_5616,N_5413,N_5496);
xnor U5617 (N_5617,N_5416,N_5425);
xnor U5618 (N_5618,N_5597,N_5439);
and U5619 (N_5619,N_5468,N_5515);
or U5620 (N_5620,N_5502,N_5473);
nor U5621 (N_5621,N_5431,N_5595);
and U5622 (N_5622,N_5542,N_5593);
xor U5623 (N_5623,N_5506,N_5520);
or U5624 (N_5624,N_5538,N_5562);
and U5625 (N_5625,N_5474,N_5500);
xnor U5626 (N_5626,N_5466,N_5546);
nor U5627 (N_5627,N_5476,N_5489);
nor U5628 (N_5628,N_5402,N_5417);
or U5629 (N_5629,N_5461,N_5537);
or U5630 (N_5630,N_5420,N_5539);
and U5631 (N_5631,N_5552,N_5460);
and U5632 (N_5632,N_5401,N_5588);
xnor U5633 (N_5633,N_5592,N_5450);
nand U5634 (N_5634,N_5579,N_5483);
nor U5635 (N_5635,N_5519,N_5509);
and U5636 (N_5636,N_5458,N_5533);
nor U5637 (N_5637,N_5530,N_5571);
nand U5638 (N_5638,N_5550,N_5400);
or U5639 (N_5639,N_5514,N_5589);
or U5640 (N_5640,N_5404,N_5532);
and U5641 (N_5641,N_5582,N_5513);
nand U5642 (N_5642,N_5491,N_5516);
xor U5643 (N_5643,N_5575,N_5536);
or U5644 (N_5644,N_5572,N_5555);
nand U5645 (N_5645,N_5449,N_5403);
or U5646 (N_5646,N_5523,N_5451);
nand U5647 (N_5647,N_5507,N_5554);
or U5648 (N_5648,N_5547,N_5493);
xor U5649 (N_5649,N_5412,N_5418);
nor U5650 (N_5650,N_5486,N_5511);
or U5651 (N_5651,N_5505,N_5591);
or U5652 (N_5652,N_5508,N_5445);
or U5653 (N_5653,N_5529,N_5434);
xor U5654 (N_5654,N_5426,N_5524);
and U5655 (N_5655,N_5424,N_5495);
nor U5656 (N_5656,N_5590,N_5477);
xor U5657 (N_5657,N_5570,N_5446);
xnor U5658 (N_5658,N_5540,N_5430);
or U5659 (N_5659,N_5442,N_5423);
xor U5660 (N_5660,N_5471,N_5528);
or U5661 (N_5661,N_5585,N_5421);
nand U5662 (N_5662,N_5429,N_5566);
and U5663 (N_5663,N_5472,N_5517);
or U5664 (N_5664,N_5553,N_5414);
or U5665 (N_5665,N_5462,N_5432);
nand U5666 (N_5666,N_5456,N_5428);
nor U5667 (N_5667,N_5544,N_5526);
xor U5668 (N_5668,N_5475,N_5457);
and U5669 (N_5669,N_5598,N_5501);
nor U5670 (N_5670,N_5427,N_5559);
and U5671 (N_5671,N_5556,N_5535);
and U5672 (N_5672,N_5581,N_5580);
nand U5673 (N_5673,N_5578,N_5564);
xnor U5674 (N_5674,N_5415,N_5422);
or U5675 (N_5675,N_5436,N_5510);
nand U5676 (N_5676,N_5527,N_5576);
xor U5677 (N_5677,N_5463,N_5573);
and U5678 (N_5678,N_5561,N_5419);
nor U5679 (N_5679,N_5409,N_5569);
nor U5680 (N_5680,N_5454,N_5433);
xnor U5681 (N_5681,N_5583,N_5464);
or U5682 (N_5682,N_5534,N_5494);
or U5683 (N_5683,N_5410,N_5465);
xnor U5684 (N_5684,N_5459,N_5437);
nand U5685 (N_5685,N_5435,N_5543);
xnor U5686 (N_5686,N_5485,N_5481);
xnor U5687 (N_5687,N_5586,N_5558);
or U5688 (N_5688,N_5512,N_5441);
nor U5689 (N_5689,N_5408,N_5599);
xor U5690 (N_5690,N_5549,N_5443);
and U5691 (N_5691,N_5577,N_5596);
or U5692 (N_5692,N_5448,N_5455);
and U5693 (N_5693,N_5541,N_5444);
nor U5694 (N_5694,N_5584,N_5492);
and U5695 (N_5695,N_5574,N_5488);
nor U5696 (N_5696,N_5452,N_5470);
nand U5697 (N_5697,N_5440,N_5521);
or U5698 (N_5698,N_5525,N_5503);
nor U5699 (N_5699,N_5545,N_5531);
xor U5700 (N_5700,N_5426,N_5564);
or U5701 (N_5701,N_5479,N_5403);
or U5702 (N_5702,N_5567,N_5453);
and U5703 (N_5703,N_5554,N_5508);
and U5704 (N_5704,N_5472,N_5511);
nand U5705 (N_5705,N_5424,N_5571);
xnor U5706 (N_5706,N_5463,N_5515);
nor U5707 (N_5707,N_5587,N_5503);
or U5708 (N_5708,N_5489,N_5482);
and U5709 (N_5709,N_5414,N_5594);
nor U5710 (N_5710,N_5420,N_5561);
nor U5711 (N_5711,N_5404,N_5464);
nor U5712 (N_5712,N_5466,N_5478);
and U5713 (N_5713,N_5533,N_5475);
nand U5714 (N_5714,N_5420,N_5493);
xnor U5715 (N_5715,N_5492,N_5591);
nor U5716 (N_5716,N_5478,N_5443);
nand U5717 (N_5717,N_5466,N_5525);
nand U5718 (N_5718,N_5581,N_5545);
nand U5719 (N_5719,N_5534,N_5420);
xor U5720 (N_5720,N_5455,N_5444);
and U5721 (N_5721,N_5438,N_5498);
nand U5722 (N_5722,N_5442,N_5445);
nor U5723 (N_5723,N_5435,N_5583);
and U5724 (N_5724,N_5411,N_5430);
and U5725 (N_5725,N_5400,N_5412);
xor U5726 (N_5726,N_5454,N_5430);
and U5727 (N_5727,N_5574,N_5447);
and U5728 (N_5728,N_5499,N_5469);
nand U5729 (N_5729,N_5561,N_5569);
nor U5730 (N_5730,N_5450,N_5586);
and U5731 (N_5731,N_5593,N_5536);
and U5732 (N_5732,N_5432,N_5574);
and U5733 (N_5733,N_5563,N_5474);
or U5734 (N_5734,N_5552,N_5497);
or U5735 (N_5735,N_5519,N_5435);
or U5736 (N_5736,N_5468,N_5480);
nand U5737 (N_5737,N_5431,N_5413);
or U5738 (N_5738,N_5527,N_5584);
nand U5739 (N_5739,N_5401,N_5454);
nand U5740 (N_5740,N_5494,N_5460);
nand U5741 (N_5741,N_5535,N_5543);
or U5742 (N_5742,N_5507,N_5531);
xnor U5743 (N_5743,N_5556,N_5526);
or U5744 (N_5744,N_5405,N_5568);
xor U5745 (N_5745,N_5551,N_5448);
or U5746 (N_5746,N_5595,N_5508);
nor U5747 (N_5747,N_5425,N_5539);
or U5748 (N_5748,N_5456,N_5541);
or U5749 (N_5749,N_5583,N_5469);
nand U5750 (N_5750,N_5499,N_5470);
and U5751 (N_5751,N_5526,N_5442);
xor U5752 (N_5752,N_5425,N_5520);
nor U5753 (N_5753,N_5565,N_5475);
nand U5754 (N_5754,N_5585,N_5514);
or U5755 (N_5755,N_5577,N_5489);
nor U5756 (N_5756,N_5584,N_5536);
or U5757 (N_5757,N_5570,N_5456);
and U5758 (N_5758,N_5560,N_5435);
and U5759 (N_5759,N_5520,N_5539);
nor U5760 (N_5760,N_5407,N_5463);
and U5761 (N_5761,N_5525,N_5502);
and U5762 (N_5762,N_5544,N_5458);
or U5763 (N_5763,N_5580,N_5462);
nor U5764 (N_5764,N_5599,N_5553);
nor U5765 (N_5765,N_5407,N_5409);
nor U5766 (N_5766,N_5488,N_5440);
xnor U5767 (N_5767,N_5570,N_5402);
nand U5768 (N_5768,N_5444,N_5404);
xnor U5769 (N_5769,N_5542,N_5467);
nor U5770 (N_5770,N_5471,N_5503);
or U5771 (N_5771,N_5588,N_5554);
or U5772 (N_5772,N_5517,N_5551);
nand U5773 (N_5773,N_5410,N_5451);
nor U5774 (N_5774,N_5485,N_5462);
nand U5775 (N_5775,N_5486,N_5562);
nor U5776 (N_5776,N_5474,N_5556);
xor U5777 (N_5777,N_5430,N_5410);
xnor U5778 (N_5778,N_5469,N_5440);
nand U5779 (N_5779,N_5403,N_5497);
or U5780 (N_5780,N_5545,N_5484);
or U5781 (N_5781,N_5463,N_5478);
or U5782 (N_5782,N_5470,N_5564);
nand U5783 (N_5783,N_5512,N_5586);
nor U5784 (N_5784,N_5531,N_5594);
nor U5785 (N_5785,N_5492,N_5442);
nor U5786 (N_5786,N_5541,N_5457);
nor U5787 (N_5787,N_5572,N_5596);
nand U5788 (N_5788,N_5560,N_5542);
nor U5789 (N_5789,N_5511,N_5431);
xor U5790 (N_5790,N_5472,N_5515);
xnor U5791 (N_5791,N_5441,N_5503);
nor U5792 (N_5792,N_5415,N_5471);
and U5793 (N_5793,N_5428,N_5492);
or U5794 (N_5794,N_5437,N_5424);
xor U5795 (N_5795,N_5439,N_5430);
xor U5796 (N_5796,N_5416,N_5412);
nor U5797 (N_5797,N_5551,N_5590);
xor U5798 (N_5798,N_5551,N_5441);
and U5799 (N_5799,N_5402,N_5512);
xor U5800 (N_5800,N_5780,N_5737);
and U5801 (N_5801,N_5690,N_5756);
nand U5802 (N_5802,N_5699,N_5747);
and U5803 (N_5803,N_5625,N_5734);
or U5804 (N_5804,N_5637,N_5604);
and U5805 (N_5805,N_5755,N_5790);
nand U5806 (N_5806,N_5698,N_5675);
nand U5807 (N_5807,N_5605,N_5719);
or U5808 (N_5808,N_5705,N_5706);
xnor U5809 (N_5809,N_5680,N_5651);
nand U5810 (N_5810,N_5621,N_5703);
or U5811 (N_5811,N_5634,N_5669);
or U5812 (N_5812,N_5733,N_5682);
or U5813 (N_5813,N_5765,N_5723);
xnor U5814 (N_5814,N_5693,N_5662);
and U5815 (N_5815,N_5670,N_5798);
and U5816 (N_5816,N_5764,N_5683);
nand U5817 (N_5817,N_5758,N_5794);
and U5818 (N_5818,N_5781,N_5799);
nand U5819 (N_5819,N_5766,N_5636);
nor U5820 (N_5820,N_5762,N_5668);
nand U5821 (N_5821,N_5757,N_5784);
or U5822 (N_5822,N_5676,N_5612);
xnor U5823 (N_5823,N_5633,N_5717);
xnor U5824 (N_5824,N_5639,N_5769);
nand U5825 (N_5825,N_5797,N_5660);
nor U5826 (N_5826,N_5772,N_5646);
xnor U5827 (N_5827,N_5736,N_5614);
xor U5828 (N_5828,N_5617,N_5658);
xor U5829 (N_5829,N_5759,N_5628);
nand U5830 (N_5830,N_5691,N_5722);
xor U5831 (N_5831,N_5602,N_5749);
nand U5832 (N_5832,N_5709,N_5638);
xor U5833 (N_5833,N_5674,N_5782);
nor U5834 (N_5834,N_5650,N_5725);
and U5835 (N_5835,N_5624,N_5620);
and U5836 (N_5836,N_5778,N_5629);
nor U5837 (N_5837,N_5679,N_5632);
nor U5838 (N_5838,N_5641,N_5652);
nand U5839 (N_5839,N_5731,N_5730);
and U5840 (N_5840,N_5788,N_5729);
and U5841 (N_5841,N_5754,N_5716);
xnor U5842 (N_5842,N_5649,N_5622);
or U5843 (N_5843,N_5606,N_5783);
or U5844 (N_5844,N_5746,N_5609);
or U5845 (N_5845,N_5603,N_5656);
and U5846 (N_5846,N_5607,N_5694);
nand U5847 (N_5847,N_5713,N_5702);
nand U5848 (N_5848,N_5710,N_5745);
or U5849 (N_5849,N_5750,N_5696);
nand U5850 (N_5850,N_5714,N_5777);
and U5851 (N_5851,N_5600,N_5791);
nor U5852 (N_5852,N_5684,N_5771);
xor U5853 (N_5853,N_5678,N_5647);
xor U5854 (N_5854,N_5643,N_5654);
nor U5855 (N_5855,N_5763,N_5775);
or U5856 (N_5856,N_5672,N_5664);
xor U5857 (N_5857,N_5613,N_5626);
xor U5858 (N_5858,N_5739,N_5774);
and U5859 (N_5859,N_5718,N_5740);
nor U5860 (N_5860,N_5751,N_5655);
xor U5861 (N_5861,N_5789,N_5610);
nand U5862 (N_5862,N_5735,N_5692);
nor U5863 (N_5863,N_5619,N_5695);
nand U5864 (N_5864,N_5688,N_5615);
nor U5865 (N_5865,N_5657,N_5689);
nand U5866 (N_5866,N_5732,N_5648);
nand U5867 (N_5867,N_5707,N_5738);
nand U5868 (N_5868,N_5792,N_5685);
or U5869 (N_5869,N_5700,N_5642);
nor U5870 (N_5870,N_5760,N_5770);
xor U5871 (N_5871,N_5616,N_5779);
xnor U5872 (N_5872,N_5761,N_5673);
xnor U5873 (N_5873,N_5666,N_5653);
nand U5874 (N_5874,N_5667,N_5708);
nand U5875 (N_5875,N_5724,N_5601);
and U5876 (N_5876,N_5630,N_5711);
nor U5877 (N_5877,N_5786,N_5742);
nand U5878 (N_5878,N_5785,N_5787);
nand U5879 (N_5879,N_5773,N_5767);
or U5880 (N_5880,N_5726,N_5795);
nor U5881 (N_5881,N_5721,N_5681);
nand U5882 (N_5882,N_5748,N_5635);
nand U5883 (N_5883,N_5712,N_5697);
or U5884 (N_5884,N_5704,N_5623);
nand U5885 (N_5885,N_5753,N_5728);
or U5886 (N_5886,N_5752,N_5663);
xnor U5887 (N_5887,N_5608,N_5645);
or U5888 (N_5888,N_5776,N_5720);
xnor U5889 (N_5889,N_5741,N_5687);
xor U5890 (N_5890,N_5618,N_5727);
xor U5891 (N_5891,N_5611,N_5644);
and U5892 (N_5892,N_5768,N_5743);
nand U5893 (N_5893,N_5659,N_5793);
nand U5894 (N_5894,N_5701,N_5677);
or U5895 (N_5895,N_5671,N_5627);
or U5896 (N_5896,N_5796,N_5665);
xor U5897 (N_5897,N_5640,N_5744);
nand U5898 (N_5898,N_5631,N_5715);
and U5899 (N_5899,N_5661,N_5686);
nor U5900 (N_5900,N_5746,N_5780);
or U5901 (N_5901,N_5640,N_5686);
xor U5902 (N_5902,N_5634,N_5706);
xor U5903 (N_5903,N_5691,N_5736);
xnor U5904 (N_5904,N_5632,N_5790);
nand U5905 (N_5905,N_5698,N_5724);
nand U5906 (N_5906,N_5606,N_5619);
and U5907 (N_5907,N_5659,N_5708);
and U5908 (N_5908,N_5754,N_5786);
nand U5909 (N_5909,N_5630,N_5745);
or U5910 (N_5910,N_5734,N_5749);
nor U5911 (N_5911,N_5647,N_5725);
and U5912 (N_5912,N_5609,N_5641);
or U5913 (N_5913,N_5694,N_5664);
xnor U5914 (N_5914,N_5616,N_5796);
nor U5915 (N_5915,N_5629,N_5708);
nor U5916 (N_5916,N_5677,N_5602);
nand U5917 (N_5917,N_5676,N_5632);
xor U5918 (N_5918,N_5764,N_5651);
xor U5919 (N_5919,N_5651,N_5678);
xor U5920 (N_5920,N_5604,N_5701);
nand U5921 (N_5921,N_5657,N_5746);
xor U5922 (N_5922,N_5766,N_5738);
nand U5923 (N_5923,N_5761,N_5685);
nand U5924 (N_5924,N_5680,N_5627);
nor U5925 (N_5925,N_5677,N_5770);
and U5926 (N_5926,N_5727,N_5625);
or U5927 (N_5927,N_5738,N_5742);
nor U5928 (N_5928,N_5765,N_5775);
or U5929 (N_5929,N_5703,N_5790);
or U5930 (N_5930,N_5671,N_5651);
or U5931 (N_5931,N_5717,N_5738);
nand U5932 (N_5932,N_5652,N_5720);
or U5933 (N_5933,N_5704,N_5734);
nand U5934 (N_5934,N_5614,N_5604);
nand U5935 (N_5935,N_5729,N_5664);
or U5936 (N_5936,N_5675,N_5706);
nand U5937 (N_5937,N_5634,N_5601);
nor U5938 (N_5938,N_5674,N_5645);
and U5939 (N_5939,N_5678,N_5673);
nor U5940 (N_5940,N_5759,N_5618);
nor U5941 (N_5941,N_5709,N_5695);
xor U5942 (N_5942,N_5645,N_5773);
nand U5943 (N_5943,N_5698,N_5772);
xor U5944 (N_5944,N_5771,N_5723);
and U5945 (N_5945,N_5757,N_5764);
nand U5946 (N_5946,N_5741,N_5601);
nor U5947 (N_5947,N_5609,N_5655);
or U5948 (N_5948,N_5673,N_5704);
nor U5949 (N_5949,N_5622,N_5744);
nand U5950 (N_5950,N_5749,N_5780);
nand U5951 (N_5951,N_5791,N_5696);
or U5952 (N_5952,N_5707,N_5650);
nand U5953 (N_5953,N_5724,N_5799);
and U5954 (N_5954,N_5781,N_5640);
nand U5955 (N_5955,N_5781,N_5750);
nand U5956 (N_5956,N_5606,N_5700);
nand U5957 (N_5957,N_5653,N_5787);
nand U5958 (N_5958,N_5697,N_5672);
and U5959 (N_5959,N_5650,N_5632);
nor U5960 (N_5960,N_5683,N_5744);
xor U5961 (N_5961,N_5661,N_5764);
nand U5962 (N_5962,N_5737,N_5656);
and U5963 (N_5963,N_5624,N_5729);
nor U5964 (N_5964,N_5725,N_5738);
or U5965 (N_5965,N_5650,N_5751);
and U5966 (N_5966,N_5785,N_5796);
or U5967 (N_5967,N_5701,N_5770);
or U5968 (N_5968,N_5698,N_5749);
nor U5969 (N_5969,N_5783,N_5702);
xor U5970 (N_5970,N_5650,N_5655);
nand U5971 (N_5971,N_5750,N_5702);
and U5972 (N_5972,N_5760,N_5773);
xnor U5973 (N_5973,N_5725,N_5643);
or U5974 (N_5974,N_5610,N_5770);
xnor U5975 (N_5975,N_5673,N_5646);
nand U5976 (N_5976,N_5775,N_5629);
xor U5977 (N_5977,N_5752,N_5711);
or U5978 (N_5978,N_5748,N_5643);
or U5979 (N_5979,N_5709,N_5684);
nand U5980 (N_5980,N_5656,N_5680);
nor U5981 (N_5981,N_5761,N_5776);
and U5982 (N_5982,N_5665,N_5780);
or U5983 (N_5983,N_5752,N_5691);
nand U5984 (N_5984,N_5656,N_5746);
nor U5985 (N_5985,N_5693,N_5673);
nor U5986 (N_5986,N_5727,N_5660);
nand U5987 (N_5987,N_5784,N_5625);
nand U5988 (N_5988,N_5707,N_5606);
and U5989 (N_5989,N_5691,N_5670);
nand U5990 (N_5990,N_5718,N_5729);
nor U5991 (N_5991,N_5634,N_5666);
and U5992 (N_5992,N_5779,N_5652);
and U5993 (N_5993,N_5723,N_5615);
and U5994 (N_5994,N_5727,N_5763);
and U5995 (N_5995,N_5780,N_5759);
xor U5996 (N_5996,N_5622,N_5741);
or U5997 (N_5997,N_5796,N_5632);
or U5998 (N_5998,N_5686,N_5628);
and U5999 (N_5999,N_5619,N_5614);
xor U6000 (N_6000,N_5883,N_5974);
xor U6001 (N_6001,N_5951,N_5966);
and U6002 (N_6002,N_5829,N_5871);
or U6003 (N_6003,N_5858,N_5999);
nor U6004 (N_6004,N_5996,N_5806);
and U6005 (N_6005,N_5949,N_5846);
nand U6006 (N_6006,N_5833,N_5895);
and U6007 (N_6007,N_5983,N_5811);
xor U6008 (N_6008,N_5938,N_5837);
xor U6009 (N_6009,N_5934,N_5845);
nor U6010 (N_6010,N_5960,N_5828);
xor U6011 (N_6011,N_5916,N_5852);
and U6012 (N_6012,N_5802,N_5910);
xnor U6013 (N_6013,N_5979,N_5939);
or U6014 (N_6014,N_5851,N_5968);
nor U6015 (N_6015,N_5900,N_5942);
and U6016 (N_6016,N_5997,N_5943);
xor U6017 (N_6017,N_5959,N_5918);
or U6018 (N_6018,N_5844,N_5957);
xor U6019 (N_6019,N_5923,N_5867);
or U6020 (N_6020,N_5931,N_5922);
nor U6021 (N_6021,N_5807,N_5946);
nor U6022 (N_6022,N_5855,N_5885);
and U6023 (N_6023,N_5898,N_5897);
nand U6024 (N_6024,N_5834,N_5995);
nor U6025 (N_6025,N_5813,N_5869);
xnor U6026 (N_6026,N_5809,N_5816);
nand U6027 (N_6027,N_5821,N_5849);
nand U6028 (N_6028,N_5964,N_5861);
or U6029 (N_6029,N_5884,N_5808);
or U6030 (N_6030,N_5881,N_5840);
and U6031 (N_6031,N_5892,N_5902);
and U6032 (N_6032,N_5819,N_5945);
nand U6033 (N_6033,N_5894,N_5986);
or U6034 (N_6034,N_5973,N_5929);
xor U6035 (N_6035,N_5870,N_5830);
nand U6036 (N_6036,N_5904,N_5928);
nand U6037 (N_6037,N_5803,N_5927);
and U6038 (N_6038,N_5952,N_5853);
xor U6039 (N_6039,N_5969,N_5890);
nor U6040 (N_6040,N_5914,N_5924);
or U6041 (N_6041,N_5956,N_5825);
or U6042 (N_6042,N_5843,N_5933);
and U6043 (N_6043,N_5990,N_5981);
nand U6044 (N_6044,N_5842,N_5859);
nand U6045 (N_6045,N_5925,N_5822);
and U6046 (N_6046,N_5972,N_5800);
nor U6047 (N_6047,N_5935,N_5814);
nor U6048 (N_6048,N_5866,N_5984);
nand U6049 (N_6049,N_5989,N_5886);
nand U6050 (N_6050,N_5907,N_5919);
or U6051 (N_6051,N_5891,N_5838);
xnor U6052 (N_6052,N_5991,N_5877);
nor U6053 (N_6053,N_5937,N_5970);
and U6054 (N_6054,N_5831,N_5947);
nor U6055 (N_6055,N_5988,N_5824);
and U6056 (N_6056,N_5889,N_5860);
nor U6057 (N_6057,N_5953,N_5868);
xnor U6058 (N_6058,N_5909,N_5872);
xor U6059 (N_6059,N_5976,N_5963);
xor U6060 (N_6060,N_5882,N_5998);
and U6061 (N_6061,N_5815,N_5926);
xnor U6062 (N_6062,N_5812,N_5874);
and U6063 (N_6063,N_5804,N_5823);
nor U6064 (N_6064,N_5832,N_5850);
nand U6065 (N_6065,N_5875,N_5917);
and U6066 (N_6066,N_5920,N_5836);
nand U6067 (N_6067,N_5805,N_5955);
nor U6068 (N_6068,N_5878,N_5978);
or U6069 (N_6069,N_5948,N_5965);
nor U6070 (N_6070,N_5985,N_5993);
or U6071 (N_6071,N_5827,N_5994);
nand U6072 (N_6072,N_5893,N_5954);
or U6073 (N_6073,N_5967,N_5908);
xnor U6074 (N_6074,N_5835,N_5899);
nor U6075 (N_6075,N_5847,N_5854);
or U6076 (N_6076,N_5839,N_5913);
xor U6077 (N_6077,N_5962,N_5876);
nand U6078 (N_6078,N_5896,N_5944);
and U6079 (N_6079,N_5941,N_5958);
nor U6080 (N_6080,N_5915,N_5903);
or U6081 (N_6081,N_5810,N_5879);
nor U6082 (N_6082,N_5950,N_5857);
or U6083 (N_6083,N_5992,N_5865);
and U6084 (N_6084,N_5930,N_5888);
nand U6085 (N_6085,N_5901,N_5864);
and U6086 (N_6086,N_5982,N_5980);
and U6087 (N_6087,N_5921,N_5940);
nand U6088 (N_6088,N_5880,N_5906);
and U6089 (N_6089,N_5905,N_5818);
nand U6090 (N_6090,N_5863,N_5826);
nand U6091 (N_6091,N_5862,N_5911);
xnor U6092 (N_6092,N_5912,N_5801);
and U6093 (N_6093,N_5987,N_5856);
or U6094 (N_6094,N_5932,N_5977);
or U6095 (N_6095,N_5975,N_5887);
nand U6096 (N_6096,N_5873,N_5936);
and U6097 (N_6097,N_5817,N_5961);
and U6098 (N_6098,N_5848,N_5820);
xor U6099 (N_6099,N_5841,N_5971);
or U6100 (N_6100,N_5870,N_5904);
nand U6101 (N_6101,N_5822,N_5868);
and U6102 (N_6102,N_5948,N_5832);
nand U6103 (N_6103,N_5824,N_5853);
and U6104 (N_6104,N_5933,N_5810);
nand U6105 (N_6105,N_5854,N_5989);
or U6106 (N_6106,N_5864,N_5947);
nand U6107 (N_6107,N_5913,N_5935);
xor U6108 (N_6108,N_5933,N_5873);
or U6109 (N_6109,N_5808,N_5926);
xor U6110 (N_6110,N_5912,N_5870);
nand U6111 (N_6111,N_5802,N_5863);
xor U6112 (N_6112,N_5839,N_5908);
and U6113 (N_6113,N_5954,N_5849);
and U6114 (N_6114,N_5813,N_5870);
nor U6115 (N_6115,N_5886,N_5915);
xnor U6116 (N_6116,N_5888,N_5880);
xor U6117 (N_6117,N_5891,N_5962);
nor U6118 (N_6118,N_5845,N_5978);
nand U6119 (N_6119,N_5871,N_5800);
nor U6120 (N_6120,N_5987,N_5958);
xor U6121 (N_6121,N_5809,N_5819);
or U6122 (N_6122,N_5970,N_5922);
or U6123 (N_6123,N_5922,N_5920);
and U6124 (N_6124,N_5876,N_5837);
or U6125 (N_6125,N_5877,N_5910);
xor U6126 (N_6126,N_5809,N_5932);
nand U6127 (N_6127,N_5807,N_5985);
nand U6128 (N_6128,N_5833,N_5965);
nor U6129 (N_6129,N_5805,N_5870);
nand U6130 (N_6130,N_5994,N_5887);
nand U6131 (N_6131,N_5967,N_5952);
and U6132 (N_6132,N_5916,N_5874);
nand U6133 (N_6133,N_5839,N_5914);
nand U6134 (N_6134,N_5970,N_5911);
xnor U6135 (N_6135,N_5930,N_5860);
xor U6136 (N_6136,N_5993,N_5921);
xor U6137 (N_6137,N_5952,N_5911);
nor U6138 (N_6138,N_5870,N_5941);
xnor U6139 (N_6139,N_5946,N_5968);
nor U6140 (N_6140,N_5823,N_5968);
xor U6141 (N_6141,N_5987,N_5936);
or U6142 (N_6142,N_5827,N_5842);
and U6143 (N_6143,N_5921,N_5970);
and U6144 (N_6144,N_5922,N_5910);
xnor U6145 (N_6145,N_5810,N_5860);
nand U6146 (N_6146,N_5968,N_5935);
xnor U6147 (N_6147,N_5942,N_5955);
and U6148 (N_6148,N_5881,N_5821);
nand U6149 (N_6149,N_5933,N_5848);
or U6150 (N_6150,N_5994,N_5886);
and U6151 (N_6151,N_5918,N_5841);
and U6152 (N_6152,N_5981,N_5842);
xor U6153 (N_6153,N_5954,N_5900);
xor U6154 (N_6154,N_5880,N_5977);
and U6155 (N_6155,N_5815,N_5835);
and U6156 (N_6156,N_5839,N_5910);
nand U6157 (N_6157,N_5992,N_5879);
and U6158 (N_6158,N_5925,N_5900);
nand U6159 (N_6159,N_5980,N_5817);
xor U6160 (N_6160,N_5953,N_5938);
or U6161 (N_6161,N_5801,N_5961);
nand U6162 (N_6162,N_5982,N_5818);
and U6163 (N_6163,N_5960,N_5987);
nor U6164 (N_6164,N_5824,N_5871);
and U6165 (N_6165,N_5819,N_5804);
nor U6166 (N_6166,N_5839,N_5990);
or U6167 (N_6167,N_5914,N_5958);
xor U6168 (N_6168,N_5919,N_5981);
or U6169 (N_6169,N_5865,N_5979);
nand U6170 (N_6170,N_5977,N_5959);
nand U6171 (N_6171,N_5950,N_5873);
xnor U6172 (N_6172,N_5933,N_5979);
nor U6173 (N_6173,N_5881,N_5910);
xnor U6174 (N_6174,N_5930,N_5855);
or U6175 (N_6175,N_5896,N_5893);
nand U6176 (N_6176,N_5904,N_5982);
xnor U6177 (N_6177,N_5976,N_5813);
nand U6178 (N_6178,N_5840,N_5938);
nor U6179 (N_6179,N_5985,N_5805);
or U6180 (N_6180,N_5974,N_5922);
xnor U6181 (N_6181,N_5813,N_5943);
nor U6182 (N_6182,N_5939,N_5951);
or U6183 (N_6183,N_5838,N_5806);
and U6184 (N_6184,N_5959,N_5932);
or U6185 (N_6185,N_5916,N_5868);
or U6186 (N_6186,N_5904,N_5873);
nand U6187 (N_6187,N_5834,N_5800);
or U6188 (N_6188,N_5901,N_5815);
xnor U6189 (N_6189,N_5869,N_5944);
xor U6190 (N_6190,N_5898,N_5857);
and U6191 (N_6191,N_5929,N_5931);
and U6192 (N_6192,N_5906,N_5806);
nor U6193 (N_6193,N_5916,N_5966);
nor U6194 (N_6194,N_5935,N_5879);
xor U6195 (N_6195,N_5877,N_5889);
or U6196 (N_6196,N_5978,N_5871);
or U6197 (N_6197,N_5855,N_5822);
or U6198 (N_6198,N_5877,N_5847);
nor U6199 (N_6199,N_5849,N_5991);
or U6200 (N_6200,N_6125,N_6148);
or U6201 (N_6201,N_6174,N_6138);
xor U6202 (N_6202,N_6112,N_6071);
nor U6203 (N_6203,N_6189,N_6085);
and U6204 (N_6204,N_6041,N_6113);
nand U6205 (N_6205,N_6039,N_6199);
nor U6206 (N_6206,N_6183,N_6172);
xor U6207 (N_6207,N_6015,N_6171);
nand U6208 (N_6208,N_6154,N_6118);
or U6209 (N_6209,N_6038,N_6068);
or U6210 (N_6210,N_6197,N_6117);
nand U6211 (N_6211,N_6175,N_6051);
nand U6212 (N_6212,N_6002,N_6170);
xor U6213 (N_6213,N_6100,N_6067);
or U6214 (N_6214,N_6110,N_6106);
and U6215 (N_6215,N_6089,N_6070);
and U6216 (N_6216,N_6166,N_6178);
nand U6217 (N_6217,N_6181,N_6021);
and U6218 (N_6218,N_6044,N_6008);
xnor U6219 (N_6219,N_6077,N_6017);
and U6220 (N_6220,N_6101,N_6005);
and U6221 (N_6221,N_6156,N_6095);
nor U6222 (N_6222,N_6091,N_6099);
xnor U6223 (N_6223,N_6130,N_6050);
nand U6224 (N_6224,N_6129,N_6014);
or U6225 (N_6225,N_6103,N_6078);
nand U6226 (N_6226,N_6036,N_6122);
nor U6227 (N_6227,N_6123,N_6093);
nor U6228 (N_6228,N_6164,N_6163);
or U6229 (N_6229,N_6132,N_6165);
nand U6230 (N_6230,N_6075,N_6143);
nor U6231 (N_6231,N_6094,N_6040);
xor U6232 (N_6232,N_6062,N_6074);
nor U6233 (N_6233,N_6114,N_6065);
or U6234 (N_6234,N_6059,N_6022);
or U6235 (N_6235,N_6063,N_6079);
and U6236 (N_6236,N_6003,N_6142);
or U6237 (N_6237,N_6058,N_6127);
nand U6238 (N_6238,N_6153,N_6048);
xor U6239 (N_6239,N_6134,N_6046);
xor U6240 (N_6240,N_6064,N_6098);
and U6241 (N_6241,N_6188,N_6032);
nand U6242 (N_6242,N_6076,N_6045);
xnor U6243 (N_6243,N_6029,N_6028);
nor U6244 (N_6244,N_6084,N_6155);
nor U6245 (N_6245,N_6157,N_6069);
and U6246 (N_6246,N_6019,N_6033);
nand U6247 (N_6247,N_6081,N_6073);
and U6248 (N_6248,N_6124,N_6027);
nand U6249 (N_6249,N_6092,N_6047);
and U6250 (N_6250,N_6140,N_6115);
nor U6251 (N_6251,N_6111,N_6147);
and U6252 (N_6252,N_6120,N_6086);
nor U6253 (N_6253,N_6090,N_6011);
or U6254 (N_6254,N_6010,N_6042);
or U6255 (N_6255,N_6168,N_6121);
and U6256 (N_6256,N_6016,N_6052);
nand U6257 (N_6257,N_6144,N_6054);
nor U6258 (N_6258,N_6167,N_6177);
and U6259 (N_6259,N_6128,N_6133);
and U6260 (N_6260,N_6191,N_6088);
and U6261 (N_6261,N_6018,N_6192);
or U6262 (N_6262,N_6026,N_6056);
and U6263 (N_6263,N_6107,N_6031);
or U6264 (N_6264,N_6173,N_6083);
xor U6265 (N_6265,N_6160,N_6151);
and U6266 (N_6266,N_6116,N_6024);
or U6267 (N_6267,N_6080,N_6158);
nor U6268 (N_6268,N_6087,N_6119);
and U6269 (N_6269,N_6061,N_6159);
nor U6270 (N_6270,N_6145,N_6057);
or U6271 (N_6271,N_6169,N_6007);
xor U6272 (N_6272,N_6072,N_6013);
xor U6273 (N_6273,N_6012,N_6187);
nor U6274 (N_6274,N_6037,N_6097);
nor U6275 (N_6275,N_6161,N_6136);
xor U6276 (N_6276,N_6135,N_6034);
nor U6277 (N_6277,N_6001,N_6198);
nor U6278 (N_6278,N_6043,N_6049);
xor U6279 (N_6279,N_6179,N_6104);
nand U6280 (N_6280,N_6146,N_6185);
xor U6281 (N_6281,N_6066,N_6162);
and U6282 (N_6282,N_6186,N_6194);
or U6283 (N_6283,N_6180,N_6195);
xor U6284 (N_6284,N_6152,N_6096);
xor U6285 (N_6285,N_6141,N_6131);
xor U6286 (N_6286,N_6139,N_6190);
or U6287 (N_6287,N_6009,N_6055);
and U6288 (N_6288,N_6108,N_6126);
nor U6289 (N_6289,N_6196,N_6184);
xor U6290 (N_6290,N_6035,N_6137);
nor U6291 (N_6291,N_6193,N_6182);
and U6292 (N_6292,N_6023,N_6004);
nor U6293 (N_6293,N_6176,N_6109);
nand U6294 (N_6294,N_6082,N_6025);
nor U6295 (N_6295,N_6006,N_6150);
nor U6296 (N_6296,N_6060,N_6053);
nor U6297 (N_6297,N_6000,N_6102);
and U6298 (N_6298,N_6020,N_6030);
or U6299 (N_6299,N_6105,N_6149);
nand U6300 (N_6300,N_6116,N_6160);
nor U6301 (N_6301,N_6013,N_6095);
and U6302 (N_6302,N_6121,N_6017);
xor U6303 (N_6303,N_6019,N_6187);
nor U6304 (N_6304,N_6156,N_6043);
nor U6305 (N_6305,N_6075,N_6152);
or U6306 (N_6306,N_6002,N_6179);
xor U6307 (N_6307,N_6167,N_6122);
or U6308 (N_6308,N_6178,N_6089);
nor U6309 (N_6309,N_6122,N_6132);
nand U6310 (N_6310,N_6137,N_6026);
and U6311 (N_6311,N_6107,N_6077);
and U6312 (N_6312,N_6155,N_6126);
nor U6313 (N_6313,N_6001,N_6141);
and U6314 (N_6314,N_6046,N_6047);
or U6315 (N_6315,N_6010,N_6182);
xor U6316 (N_6316,N_6186,N_6121);
nand U6317 (N_6317,N_6116,N_6166);
xnor U6318 (N_6318,N_6164,N_6055);
nand U6319 (N_6319,N_6006,N_6101);
and U6320 (N_6320,N_6050,N_6124);
xor U6321 (N_6321,N_6141,N_6086);
xor U6322 (N_6322,N_6017,N_6068);
nand U6323 (N_6323,N_6059,N_6080);
nand U6324 (N_6324,N_6069,N_6046);
or U6325 (N_6325,N_6020,N_6093);
and U6326 (N_6326,N_6192,N_6186);
xnor U6327 (N_6327,N_6056,N_6000);
nor U6328 (N_6328,N_6009,N_6082);
and U6329 (N_6329,N_6025,N_6095);
nand U6330 (N_6330,N_6054,N_6077);
or U6331 (N_6331,N_6120,N_6146);
nor U6332 (N_6332,N_6062,N_6096);
or U6333 (N_6333,N_6131,N_6124);
nand U6334 (N_6334,N_6010,N_6099);
or U6335 (N_6335,N_6149,N_6119);
and U6336 (N_6336,N_6105,N_6024);
nor U6337 (N_6337,N_6052,N_6046);
and U6338 (N_6338,N_6194,N_6112);
nor U6339 (N_6339,N_6079,N_6162);
nand U6340 (N_6340,N_6185,N_6081);
nor U6341 (N_6341,N_6062,N_6072);
nand U6342 (N_6342,N_6082,N_6133);
and U6343 (N_6343,N_6093,N_6111);
nand U6344 (N_6344,N_6140,N_6147);
nand U6345 (N_6345,N_6120,N_6015);
nand U6346 (N_6346,N_6047,N_6071);
or U6347 (N_6347,N_6169,N_6166);
xor U6348 (N_6348,N_6122,N_6041);
and U6349 (N_6349,N_6020,N_6148);
nor U6350 (N_6350,N_6106,N_6046);
xor U6351 (N_6351,N_6111,N_6098);
nor U6352 (N_6352,N_6171,N_6039);
xnor U6353 (N_6353,N_6050,N_6139);
xnor U6354 (N_6354,N_6081,N_6104);
xor U6355 (N_6355,N_6162,N_6052);
and U6356 (N_6356,N_6188,N_6154);
nor U6357 (N_6357,N_6155,N_6095);
nor U6358 (N_6358,N_6167,N_6110);
or U6359 (N_6359,N_6018,N_6077);
xor U6360 (N_6360,N_6102,N_6137);
nand U6361 (N_6361,N_6176,N_6145);
nor U6362 (N_6362,N_6053,N_6076);
or U6363 (N_6363,N_6037,N_6036);
xnor U6364 (N_6364,N_6086,N_6149);
nor U6365 (N_6365,N_6086,N_6020);
xnor U6366 (N_6366,N_6195,N_6068);
xnor U6367 (N_6367,N_6068,N_6067);
or U6368 (N_6368,N_6197,N_6157);
nor U6369 (N_6369,N_6029,N_6067);
xor U6370 (N_6370,N_6096,N_6045);
nor U6371 (N_6371,N_6043,N_6166);
nand U6372 (N_6372,N_6054,N_6068);
nand U6373 (N_6373,N_6055,N_6148);
xor U6374 (N_6374,N_6077,N_6171);
or U6375 (N_6375,N_6034,N_6118);
and U6376 (N_6376,N_6121,N_6036);
xnor U6377 (N_6377,N_6185,N_6067);
xnor U6378 (N_6378,N_6110,N_6055);
xor U6379 (N_6379,N_6126,N_6112);
and U6380 (N_6380,N_6174,N_6117);
or U6381 (N_6381,N_6157,N_6191);
and U6382 (N_6382,N_6027,N_6196);
xor U6383 (N_6383,N_6029,N_6161);
nand U6384 (N_6384,N_6071,N_6136);
or U6385 (N_6385,N_6121,N_6080);
and U6386 (N_6386,N_6157,N_6045);
nor U6387 (N_6387,N_6078,N_6030);
and U6388 (N_6388,N_6148,N_6145);
and U6389 (N_6389,N_6050,N_6126);
xor U6390 (N_6390,N_6062,N_6131);
nand U6391 (N_6391,N_6146,N_6086);
xor U6392 (N_6392,N_6014,N_6055);
xor U6393 (N_6393,N_6156,N_6070);
xnor U6394 (N_6394,N_6014,N_6124);
nor U6395 (N_6395,N_6057,N_6149);
xnor U6396 (N_6396,N_6109,N_6023);
nand U6397 (N_6397,N_6164,N_6107);
nand U6398 (N_6398,N_6131,N_6066);
xnor U6399 (N_6399,N_6110,N_6010);
xor U6400 (N_6400,N_6212,N_6297);
xor U6401 (N_6401,N_6291,N_6215);
nor U6402 (N_6402,N_6306,N_6271);
nand U6403 (N_6403,N_6221,N_6294);
or U6404 (N_6404,N_6227,N_6396);
xor U6405 (N_6405,N_6246,N_6357);
nor U6406 (N_6406,N_6207,N_6243);
nand U6407 (N_6407,N_6301,N_6398);
xnor U6408 (N_6408,N_6372,N_6392);
xnor U6409 (N_6409,N_6397,N_6364);
nand U6410 (N_6410,N_6395,N_6314);
nor U6411 (N_6411,N_6210,N_6299);
nand U6412 (N_6412,N_6278,N_6265);
nand U6413 (N_6413,N_6322,N_6348);
nand U6414 (N_6414,N_6262,N_6270);
nand U6415 (N_6415,N_6283,N_6237);
xnor U6416 (N_6416,N_6287,N_6379);
nand U6417 (N_6417,N_6341,N_6374);
or U6418 (N_6418,N_6268,N_6228);
nand U6419 (N_6419,N_6368,N_6276);
and U6420 (N_6420,N_6361,N_6393);
or U6421 (N_6421,N_6277,N_6256);
nand U6422 (N_6422,N_6209,N_6344);
nor U6423 (N_6423,N_6318,N_6376);
and U6424 (N_6424,N_6213,N_6273);
nand U6425 (N_6425,N_6390,N_6244);
nand U6426 (N_6426,N_6319,N_6292);
and U6427 (N_6427,N_6369,N_6308);
nor U6428 (N_6428,N_6231,N_6248);
and U6429 (N_6429,N_6229,N_6388);
nand U6430 (N_6430,N_6206,N_6238);
nor U6431 (N_6431,N_6370,N_6387);
nand U6432 (N_6432,N_6200,N_6326);
and U6433 (N_6433,N_6303,N_6208);
or U6434 (N_6434,N_6226,N_6217);
nand U6435 (N_6435,N_6358,N_6317);
and U6436 (N_6436,N_6340,N_6331);
or U6437 (N_6437,N_6345,N_6293);
or U6438 (N_6438,N_6282,N_6320);
nand U6439 (N_6439,N_6281,N_6383);
and U6440 (N_6440,N_6360,N_6218);
or U6441 (N_6441,N_6362,N_6295);
nand U6442 (N_6442,N_6216,N_6359);
nand U6443 (N_6443,N_6343,N_6381);
nor U6444 (N_6444,N_6384,N_6353);
xor U6445 (N_6445,N_6267,N_6234);
xor U6446 (N_6446,N_6236,N_6219);
xnor U6447 (N_6447,N_6252,N_6300);
and U6448 (N_6448,N_6366,N_6241);
and U6449 (N_6449,N_6272,N_6230);
nor U6450 (N_6450,N_6232,N_6264);
nand U6451 (N_6451,N_6222,N_6355);
or U6452 (N_6452,N_6202,N_6380);
xnor U6453 (N_6453,N_6205,N_6332);
xor U6454 (N_6454,N_6335,N_6255);
xnor U6455 (N_6455,N_6338,N_6240);
nand U6456 (N_6456,N_6346,N_6214);
or U6457 (N_6457,N_6328,N_6285);
and U6458 (N_6458,N_6349,N_6224);
and U6459 (N_6459,N_6286,N_6352);
nor U6460 (N_6460,N_6251,N_6254);
xor U6461 (N_6461,N_6225,N_6223);
xor U6462 (N_6462,N_6263,N_6249);
or U6463 (N_6463,N_6288,N_6324);
xor U6464 (N_6464,N_6310,N_6386);
and U6465 (N_6465,N_6356,N_6329);
or U6466 (N_6466,N_6367,N_6375);
or U6467 (N_6467,N_6347,N_6305);
nor U6468 (N_6468,N_6258,N_6253);
or U6469 (N_6469,N_6257,N_6284);
xnor U6470 (N_6470,N_6204,N_6203);
or U6471 (N_6471,N_6269,N_6337);
or U6472 (N_6472,N_6309,N_6350);
and U6473 (N_6473,N_6321,N_6260);
nor U6474 (N_6474,N_6354,N_6266);
or U6475 (N_6475,N_6327,N_6211);
nor U6476 (N_6476,N_6336,N_6298);
nor U6477 (N_6477,N_6399,N_6242);
nand U6478 (N_6478,N_6261,N_6233);
nor U6479 (N_6479,N_6296,N_6325);
nor U6480 (N_6480,N_6279,N_6290);
and U6481 (N_6481,N_6259,N_6311);
or U6482 (N_6482,N_6365,N_6389);
nand U6483 (N_6483,N_6312,N_6247);
nor U6484 (N_6484,N_6373,N_6201);
or U6485 (N_6485,N_6385,N_6235);
nand U6486 (N_6486,N_6334,N_6289);
nor U6487 (N_6487,N_6378,N_6363);
or U6488 (N_6488,N_6316,N_6323);
or U6489 (N_6489,N_6351,N_6391);
nand U6490 (N_6490,N_6339,N_6313);
and U6491 (N_6491,N_6330,N_6307);
or U6492 (N_6492,N_6394,N_6250);
nor U6493 (N_6493,N_6371,N_6342);
and U6494 (N_6494,N_6220,N_6280);
or U6495 (N_6495,N_6274,N_6245);
or U6496 (N_6496,N_6275,N_6304);
or U6497 (N_6497,N_6382,N_6315);
or U6498 (N_6498,N_6239,N_6333);
nor U6499 (N_6499,N_6377,N_6302);
nor U6500 (N_6500,N_6298,N_6308);
nand U6501 (N_6501,N_6202,N_6358);
or U6502 (N_6502,N_6275,N_6386);
nor U6503 (N_6503,N_6368,N_6337);
nor U6504 (N_6504,N_6395,N_6227);
nor U6505 (N_6505,N_6366,N_6353);
xor U6506 (N_6506,N_6275,N_6237);
and U6507 (N_6507,N_6212,N_6249);
nor U6508 (N_6508,N_6254,N_6292);
or U6509 (N_6509,N_6382,N_6225);
nand U6510 (N_6510,N_6388,N_6329);
nand U6511 (N_6511,N_6347,N_6277);
nand U6512 (N_6512,N_6349,N_6303);
xnor U6513 (N_6513,N_6394,N_6348);
nand U6514 (N_6514,N_6243,N_6337);
or U6515 (N_6515,N_6237,N_6327);
nor U6516 (N_6516,N_6293,N_6202);
nand U6517 (N_6517,N_6314,N_6216);
and U6518 (N_6518,N_6200,N_6251);
and U6519 (N_6519,N_6310,N_6200);
nor U6520 (N_6520,N_6348,N_6204);
nor U6521 (N_6521,N_6247,N_6354);
nor U6522 (N_6522,N_6307,N_6217);
xnor U6523 (N_6523,N_6274,N_6242);
nand U6524 (N_6524,N_6386,N_6364);
and U6525 (N_6525,N_6212,N_6263);
and U6526 (N_6526,N_6331,N_6342);
xnor U6527 (N_6527,N_6315,N_6323);
nand U6528 (N_6528,N_6241,N_6264);
and U6529 (N_6529,N_6354,N_6252);
xnor U6530 (N_6530,N_6398,N_6286);
nor U6531 (N_6531,N_6267,N_6298);
and U6532 (N_6532,N_6382,N_6246);
nand U6533 (N_6533,N_6390,N_6335);
or U6534 (N_6534,N_6249,N_6353);
xor U6535 (N_6535,N_6214,N_6281);
and U6536 (N_6536,N_6350,N_6337);
xnor U6537 (N_6537,N_6392,N_6323);
and U6538 (N_6538,N_6326,N_6357);
and U6539 (N_6539,N_6297,N_6315);
and U6540 (N_6540,N_6264,N_6375);
or U6541 (N_6541,N_6288,N_6244);
nand U6542 (N_6542,N_6375,N_6332);
or U6543 (N_6543,N_6208,N_6216);
nand U6544 (N_6544,N_6266,N_6274);
xor U6545 (N_6545,N_6234,N_6312);
or U6546 (N_6546,N_6358,N_6307);
or U6547 (N_6547,N_6341,N_6246);
xor U6548 (N_6548,N_6225,N_6211);
nor U6549 (N_6549,N_6341,N_6233);
xnor U6550 (N_6550,N_6242,N_6211);
nor U6551 (N_6551,N_6213,N_6350);
or U6552 (N_6552,N_6389,N_6287);
xnor U6553 (N_6553,N_6396,N_6235);
nor U6554 (N_6554,N_6317,N_6316);
and U6555 (N_6555,N_6236,N_6280);
nand U6556 (N_6556,N_6363,N_6223);
nor U6557 (N_6557,N_6385,N_6397);
or U6558 (N_6558,N_6338,N_6372);
nand U6559 (N_6559,N_6221,N_6318);
nand U6560 (N_6560,N_6219,N_6364);
and U6561 (N_6561,N_6245,N_6310);
xor U6562 (N_6562,N_6264,N_6389);
nor U6563 (N_6563,N_6284,N_6238);
or U6564 (N_6564,N_6266,N_6299);
nand U6565 (N_6565,N_6270,N_6217);
nand U6566 (N_6566,N_6343,N_6204);
or U6567 (N_6567,N_6217,N_6353);
and U6568 (N_6568,N_6304,N_6286);
and U6569 (N_6569,N_6389,N_6216);
nor U6570 (N_6570,N_6231,N_6360);
nand U6571 (N_6571,N_6364,N_6376);
and U6572 (N_6572,N_6213,N_6295);
and U6573 (N_6573,N_6293,N_6347);
or U6574 (N_6574,N_6320,N_6341);
nor U6575 (N_6575,N_6368,N_6363);
and U6576 (N_6576,N_6232,N_6281);
nand U6577 (N_6577,N_6278,N_6243);
nor U6578 (N_6578,N_6351,N_6212);
nor U6579 (N_6579,N_6397,N_6289);
nor U6580 (N_6580,N_6342,N_6381);
nor U6581 (N_6581,N_6389,N_6344);
nor U6582 (N_6582,N_6263,N_6347);
and U6583 (N_6583,N_6278,N_6210);
nand U6584 (N_6584,N_6204,N_6243);
and U6585 (N_6585,N_6298,N_6213);
xnor U6586 (N_6586,N_6295,N_6207);
xnor U6587 (N_6587,N_6229,N_6343);
nand U6588 (N_6588,N_6208,N_6329);
xnor U6589 (N_6589,N_6340,N_6202);
and U6590 (N_6590,N_6309,N_6346);
xor U6591 (N_6591,N_6315,N_6309);
nor U6592 (N_6592,N_6386,N_6239);
nand U6593 (N_6593,N_6358,N_6361);
xnor U6594 (N_6594,N_6376,N_6325);
xnor U6595 (N_6595,N_6375,N_6243);
nor U6596 (N_6596,N_6353,N_6381);
nand U6597 (N_6597,N_6287,N_6233);
nand U6598 (N_6598,N_6325,N_6274);
xor U6599 (N_6599,N_6289,N_6387);
nand U6600 (N_6600,N_6534,N_6500);
and U6601 (N_6601,N_6514,N_6456);
xor U6602 (N_6602,N_6441,N_6538);
nor U6603 (N_6603,N_6458,N_6584);
and U6604 (N_6604,N_6505,N_6537);
and U6605 (N_6605,N_6546,N_6472);
xnor U6606 (N_6606,N_6560,N_6501);
or U6607 (N_6607,N_6433,N_6462);
xor U6608 (N_6608,N_6585,N_6450);
and U6609 (N_6609,N_6463,N_6571);
nand U6610 (N_6610,N_6561,N_6454);
or U6611 (N_6611,N_6532,N_6528);
xor U6612 (N_6612,N_6429,N_6564);
or U6613 (N_6613,N_6540,N_6521);
xnor U6614 (N_6614,N_6533,N_6597);
nand U6615 (N_6615,N_6555,N_6594);
nor U6616 (N_6616,N_6440,N_6490);
or U6617 (N_6617,N_6581,N_6599);
xnor U6618 (N_6618,N_6495,N_6474);
and U6619 (N_6619,N_6436,N_6575);
nand U6620 (N_6620,N_6460,N_6589);
nor U6621 (N_6621,N_6475,N_6570);
or U6622 (N_6622,N_6576,N_6473);
or U6623 (N_6623,N_6497,N_6542);
nor U6624 (N_6624,N_6574,N_6545);
nand U6625 (N_6625,N_6554,N_6407);
nand U6626 (N_6626,N_6579,N_6493);
nor U6627 (N_6627,N_6513,N_6481);
xnor U6628 (N_6628,N_6419,N_6479);
nor U6629 (N_6629,N_6519,N_6438);
nor U6630 (N_6630,N_6518,N_6544);
and U6631 (N_6631,N_6583,N_6580);
nor U6632 (N_6632,N_6443,N_6411);
nand U6633 (N_6633,N_6476,N_6483);
and U6634 (N_6634,N_6509,N_6435);
or U6635 (N_6635,N_6568,N_6563);
and U6636 (N_6636,N_6428,N_6515);
nand U6637 (N_6637,N_6426,N_6502);
and U6638 (N_6638,N_6551,N_6437);
or U6639 (N_6639,N_6446,N_6427);
nor U6640 (N_6640,N_6447,N_6491);
xor U6641 (N_6641,N_6558,N_6482);
xnor U6642 (N_6642,N_6452,N_6413);
and U6643 (N_6643,N_6531,N_6567);
and U6644 (N_6644,N_6402,N_6480);
nor U6645 (N_6645,N_6424,N_6525);
or U6646 (N_6646,N_6586,N_6477);
nor U6647 (N_6647,N_6569,N_6582);
xor U6648 (N_6648,N_6592,N_6549);
nor U6649 (N_6649,N_6595,N_6489);
xnor U6650 (N_6650,N_6449,N_6520);
or U6651 (N_6651,N_6448,N_6539);
nand U6652 (N_6652,N_6425,N_6457);
xor U6653 (N_6653,N_6529,N_6504);
or U6654 (N_6654,N_6503,N_6562);
nand U6655 (N_6655,N_6484,N_6400);
or U6656 (N_6656,N_6578,N_6530);
nor U6657 (N_6657,N_6598,N_6478);
and U6658 (N_6658,N_6432,N_6535);
nand U6659 (N_6659,N_6418,N_6403);
nand U6660 (N_6660,N_6445,N_6467);
nor U6661 (N_6661,N_6593,N_6486);
and U6662 (N_6662,N_6557,N_6414);
xnor U6663 (N_6663,N_6439,N_6409);
or U6664 (N_6664,N_6408,N_6485);
and U6665 (N_6665,N_6469,N_6421);
xnor U6666 (N_6666,N_6417,N_6517);
or U6667 (N_6667,N_6526,N_6543);
or U6668 (N_6668,N_6512,N_6487);
nand U6669 (N_6669,N_6524,N_6455);
xor U6670 (N_6670,N_6412,N_6466);
nand U6671 (N_6671,N_6494,N_6507);
and U6672 (N_6672,N_6415,N_6550);
or U6673 (N_6673,N_6465,N_6488);
nor U6674 (N_6674,N_6468,N_6566);
xor U6675 (N_6675,N_6552,N_6461);
nand U6676 (N_6676,N_6508,N_6434);
or U6677 (N_6677,N_6511,N_6470);
and U6678 (N_6678,N_6516,N_6565);
xor U6679 (N_6679,N_6577,N_6523);
and U6680 (N_6680,N_6406,N_6587);
and U6681 (N_6681,N_6453,N_6553);
xor U6682 (N_6682,N_6401,N_6591);
and U6683 (N_6683,N_6590,N_6442);
nor U6684 (N_6684,N_6405,N_6559);
or U6685 (N_6685,N_6510,N_6536);
and U6686 (N_6686,N_6423,N_6506);
xnor U6687 (N_6687,N_6459,N_6588);
or U6688 (N_6688,N_6451,N_6464);
and U6689 (N_6689,N_6444,N_6430);
xnor U6690 (N_6690,N_6471,N_6431);
xnor U6691 (N_6691,N_6499,N_6527);
or U6692 (N_6692,N_6596,N_6496);
and U6693 (N_6693,N_6548,N_6410);
and U6694 (N_6694,N_6404,N_6556);
xnor U6695 (N_6695,N_6420,N_6422);
nand U6696 (N_6696,N_6547,N_6541);
or U6697 (N_6697,N_6492,N_6573);
nor U6698 (N_6698,N_6572,N_6498);
nand U6699 (N_6699,N_6522,N_6416);
xnor U6700 (N_6700,N_6419,N_6527);
nor U6701 (N_6701,N_6584,N_6439);
and U6702 (N_6702,N_6514,N_6440);
xnor U6703 (N_6703,N_6510,N_6539);
or U6704 (N_6704,N_6474,N_6531);
nand U6705 (N_6705,N_6596,N_6599);
nand U6706 (N_6706,N_6444,N_6545);
xnor U6707 (N_6707,N_6552,N_6481);
xor U6708 (N_6708,N_6499,N_6503);
nand U6709 (N_6709,N_6564,N_6557);
and U6710 (N_6710,N_6532,N_6444);
nand U6711 (N_6711,N_6558,N_6486);
or U6712 (N_6712,N_6449,N_6475);
nor U6713 (N_6713,N_6441,N_6571);
xnor U6714 (N_6714,N_6446,N_6574);
nor U6715 (N_6715,N_6544,N_6498);
nand U6716 (N_6716,N_6579,N_6542);
or U6717 (N_6717,N_6457,N_6476);
nand U6718 (N_6718,N_6499,N_6538);
or U6719 (N_6719,N_6517,N_6443);
nor U6720 (N_6720,N_6472,N_6436);
nor U6721 (N_6721,N_6551,N_6534);
and U6722 (N_6722,N_6576,N_6590);
nand U6723 (N_6723,N_6537,N_6528);
nor U6724 (N_6724,N_6486,N_6475);
or U6725 (N_6725,N_6456,N_6427);
or U6726 (N_6726,N_6569,N_6521);
or U6727 (N_6727,N_6488,N_6420);
or U6728 (N_6728,N_6410,N_6403);
and U6729 (N_6729,N_6427,N_6550);
nor U6730 (N_6730,N_6476,N_6489);
or U6731 (N_6731,N_6455,N_6471);
xor U6732 (N_6732,N_6532,N_6494);
or U6733 (N_6733,N_6479,N_6412);
and U6734 (N_6734,N_6596,N_6415);
nor U6735 (N_6735,N_6474,N_6519);
xor U6736 (N_6736,N_6516,N_6457);
xor U6737 (N_6737,N_6492,N_6400);
xnor U6738 (N_6738,N_6563,N_6418);
nor U6739 (N_6739,N_6410,N_6468);
xor U6740 (N_6740,N_6592,N_6418);
nor U6741 (N_6741,N_6534,N_6457);
nor U6742 (N_6742,N_6451,N_6585);
xor U6743 (N_6743,N_6576,N_6462);
xnor U6744 (N_6744,N_6514,N_6444);
nand U6745 (N_6745,N_6483,N_6566);
xnor U6746 (N_6746,N_6572,N_6566);
nor U6747 (N_6747,N_6456,N_6562);
xnor U6748 (N_6748,N_6522,N_6566);
or U6749 (N_6749,N_6568,N_6492);
and U6750 (N_6750,N_6544,N_6550);
nor U6751 (N_6751,N_6559,N_6421);
or U6752 (N_6752,N_6577,N_6563);
xor U6753 (N_6753,N_6581,N_6402);
nor U6754 (N_6754,N_6453,N_6447);
and U6755 (N_6755,N_6513,N_6476);
nand U6756 (N_6756,N_6586,N_6472);
or U6757 (N_6757,N_6458,N_6425);
nor U6758 (N_6758,N_6415,N_6434);
nand U6759 (N_6759,N_6460,N_6480);
nor U6760 (N_6760,N_6581,N_6596);
or U6761 (N_6761,N_6591,N_6510);
nor U6762 (N_6762,N_6405,N_6546);
nor U6763 (N_6763,N_6512,N_6546);
and U6764 (N_6764,N_6477,N_6551);
xnor U6765 (N_6765,N_6558,N_6542);
and U6766 (N_6766,N_6529,N_6596);
nor U6767 (N_6767,N_6548,N_6539);
nand U6768 (N_6768,N_6537,N_6532);
xor U6769 (N_6769,N_6550,N_6473);
or U6770 (N_6770,N_6485,N_6538);
nand U6771 (N_6771,N_6477,N_6516);
nand U6772 (N_6772,N_6575,N_6442);
nor U6773 (N_6773,N_6497,N_6455);
or U6774 (N_6774,N_6483,N_6443);
nand U6775 (N_6775,N_6451,N_6481);
nor U6776 (N_6776,N_6410,N_6494);
nor U6777 (N_6777,N_6508,N_6420);
or U6778 (N_6778,N_6569,N_6531);
or U6779 (N_6779,N_6497,N_6456);
nor U6780 (N_6780,N_6432,N_6481);
nand U6781 (N_6781,N_6446,N_6442);
nand U6782 (N_6782,N_6500,N_6549);
and U6783 (N_6783,N_6400,N_6594);
and U6784 (N_6784,N_6428,N_6512);
or U6785 (N_6785,N_6423,N_6489);
nor U6786 (N_6786,N_6503,N_6474);
or U6787 (N_6787,N_6569,N_6517);
or U6788 (N_6788,N_6466,N_6591);
nand U6789 (N_6789,N_6456,N_6459);
or U6790 (N_6790,N_6594,N_6564);
and U6791 (N_6791,N_6583,N_6410);
nand U6792 (N_6792,N_6483,N_6543);
or U6793 (N_6793,N_6528,N_6591);
nor U6794 (N_6794,N_6512,N_6575);
xor U6795 (N_6795,N_6596,N_6409);
nand U6796 (N_6796,N_6407,N_6421);
nor U6797 (N_6797,N_6559,N_6512);
or U6798 (N_6798,N_6448,N_6438);
or U6799 (N_6799,N_6589,N_6572);
or U6800 (N_6800,N_6727,N_6773);
nand U6801 (N_6801,N_6637,N_6781);
xor U6802 (N_6802,N_6624,N_6605);
xnor U6803 (N_6803,N_6627,N_6797);
and U6804 (N_6804,N_6633,N_6775);
and U6805 (N_6805,N_6607,N_6794);
xor U6806 (N_6806,N_6748,N_6740);
nor U6807 (N_6807,N_6616,N_6666);
or U6808 (N_6808,N_6609,N_6745);
nand U6809 (N_6809,N_6723,N_6789);
or U6810 (N_6810,N_6731,N_6758);
nor U6811 (N_6811,N_6643,N_6612);
nor U6812 (N_6812,N_6790,N_6788);
nand U6813 (N_6813,N_6630,N_6702);
nor U6814 (N_6814,N_6747,N_6683);
xnor U6815 (N_6815,N_6680,N_6645);
and U6816 (N_6816,N_6783,N_6736);
nand U6817 (N_6817,N_6777,N_6686);
or U6818 (N_6818,N_6798,N_6741);
nor U6819 (N_6819,N_6614,N_6765);
nor U6820 (N_6820,N_6682,N_6601);
xor U6821 (N_6821,N_6655,N_6664);
nand U6822 (N_6822,N_6779,N_6722);
xnor U6823 (N_6823,N_6674,N_6752);
and U6824 (N_6824,N_6638,N_6795);
nor U6825 (N_6825,N_6690,N_6688);
nand U6826 (N_6826,N_6749,N_6782);
and U6827 (N_6827,N_6687,N_6753);
or U6828 (N_6828,N_6604,N_6620);
xor U6829 (N_6829,N_6689,N_6778);
and U6830 (N_6830,N_6771,N_6712);
or U6831 (N_6831,N_6654,N_6634);
and U6832 (N_6832,N_6673,N_6720);
nand U6833 (N_6833,N_6754,N_6602);
and U6834 (N_6834,N_6791,N_6663);
nand U6835 (N_6835,N_6713,N_6640);
and U6836 (N_6836,N_6715,N_6792);
xor U6837 (N_6837,N_6606,N_6732);
or U6838 (N_6838,N_6608,N_6691);
nand U6839 (N_6839,N_6636,N_6676);
and U6840 (N_6840,N_6632,N_6668);
and U6841 (N_6841,N_6684,N_6737);
xor U6842 (N_6842,N_6610,N_6649);
or U6843 (N_6843,N_6743,N_6685);
xor U6844 (N_6844,N_6787,N_6717);
nand U6845 (N_6845,N_6639,N_6660);
nand U6846 (N_6846,N_6622,N_6796);
nand U6847 (N_6847,N_6770,N_6619);
or U6848 (N_6848,N_6651,N_6644);
nor U6849 (N_6849,N_6729,N_6657);
xnor U6850 (N_6850,N_6780,N_6628);
nor U6851 (N_6851,N_6603,N_6786);
nand U6852 (N_6852,N_6709,N_6793);
or U6853 (N_6853,N_6653,N_6799);
nand U6854 (N_6854,N_6719,N_6652);
nand U6855 (N_6855,N_6725,N_6623);
nor U6856 (N_6856,N_6751,N_6726);
nor U6857 (N_6857,N_6759,N_6734);
or U6858 (N_6858,N_6744,N_6647);
xor U6859 (N_6859,N_6703,N_6648);
nand U6860 (N_6860,N_6711,N_6698);
or U6861 (N_6861,N_6662,N_6667);
and U6862 (N_6862,N_6710,N_6700);
or U6863 (N_6863,N_6728,N_6738);
or U6864 (N_6864,N_6769,N_6707);
nand U6865 (N_6865,N_6646,N_6768);
or U6866 (N_6866,N_6661,N_6762);
or U6867 (N_6867,N_6739,N_6756);
nand U6868 (N_6868,N_6656,N_6600);
nor U6869 (N_6869,N_6699,N_6642);
xor U6870 (N_6870,N_6716,N_6692);
xnor U6871 (N_6871,N_6615,N_6681);
nor U6872 (N_6872,N_6705,N_6650);
nand U6873 (N_6873,N_6733,N_6735);
and U6874 (N_6874,N_6697,N_6761);
xor U6875 (N_6875,N_6704,N_6658);
nand U6876 (N_6876,N_6669,N_6613);
nor U6877 (N_6877,N_6678,N_6672);
nor U6878 (N_6878,N_6665,N_6784);
nand U6879 (N_6879,N_6631,N_6695);
nor U6880 (N_6880,N_6785,N_6696);
and U6881 (N_6881,N_6763,N_6659);
xnor U6882 (N_6882,N_6679,N_6635);
nor U6883 (N_6883,N_6746,N_6776);
or U6884 (N_6884,N_6706,N_6757);
nand U6885 (N_6885,N_6701,N_6764);
and U6886 (N_6886,N_6670,N_6625);
xnor U6887 (N_6887,N_6694,N_6772);
or U6888 (N_6888,N_6611,N_6714);
nand U6889 (N_6889,N_6730,N_6693);
nand U6890 (N_6890,N_6617,N_6675);
xor U6891 (N_6891,N_6755,N_6767);
nand U6892 (N_6892,N_6621,N_6718);
nor U6893 (N_6893,N_6629,N_6750);
xnor U6894 (N_6894,N_6742,N_6766);
nand U6895 (N_6895,N_6618,N_6677);
nand U6896 (N_6896,N_6641,N_6721);
xor U6897 (N_6897,N_6708,N_6671);
and U6898 (N_6898,N_6626,N_6774);
or U6899 (N_6899,N_6724,N_6760);
nand U6900 (N_6900,N_6631,N_6727);
and U6901 (N_6901,N_6746,N_6672);
xnor U6902 (N_6902,N_6644,N_6764);
nor U6903 (N_6903,N_6780,N_6602);
xnor U6904 (N_6904,N_6662,N_6604);
nand U6905 (N_6905,N_6704,N_6626);
nand U6906 (N_6906,N_6706,N_6796);
xnor U6907 (N_6907,N_6744,N_6760);
or U6908 (N_6908,N_6609,N_6601);
and U6909 (N_6909,N_6690,N_6694);
nand U6910 (N_6910,N_6760,N_6637);
and U6911 (N_6911,N_6693,N_6685);
nand U6912 (N_6912,N_6676,N_6668);
and U6913 (N_6913,N_6603,N_6789);
nor U6914 (N_6914,N_6616,N_6626);
nor U6915 (N_6915,N_6653,N_6623);
nor U6916 (N_6916,N_6762,N_6765);
and U6917 (N_6917,N_6765,N_6729);
or U6918 (N_6918,N_6643,N_6757);
nor U6919 (N_6919,N_6727,N_6703);
and U6920 (N_6920,N_6720,N_6649);
nand U6921 (N_6921,N_6601,N_6600);
nand U6922 (N_6922,N_6646,N_6676);
xor U6923 (N_6923,N_6795,N_6634);
nand U6924 (N_6924,N_6715,N_6617);
xnor U6925 (N_6925,N_6728,N_6696);
xnor U6926 (N_6926,N_6611,N_6647);
xnor U6927 (N_6927,N_6649,N_6707);
nor U6928 (N_6928,N_6778,N_6729);
nand U6929 (N_6929,N_6691,N_6634);
nor U6930 (N_6930,N_6635,N_6753);
and U6931 (N_6931,N_6629,N_6625);
nand U6932 (N_6932,N_6791,N_6761);
nor U6933 (N_6933,N_6626,N_6799);
and U6934 (N_6934,N_6790,N_6763);
or U6935 (N_6935,N_6690,N_6735);
xor U6936 (N_6936,N_6611,N_6777);
nand U6937 (N_6937,N_6606,N_6738);
or U6938 (N_6938,N_6687,N_6669);
and U6939 (N_6939,N_6689,N_6713);
nand U6940 (N_6940,N_6787,N_6668);
or U6941 (N_6941,N_6688,N_6610);
or U6942 (N_6942,N_6734,N_6676);
nand U6943 (N_6943,N_6687,N_6793);
nor U6944 (N_6944,N_6680,N_6617);
and U6945 (N_6945,N_6767,N_6716);
nand U6946 (N_6946,N_6669,N_6748);
and U6947 (N_6947,N_6693,N_6656);
and U6948 (N_6948,N_6771,N_6656);
nor U6949 (N_6949,N_6641,N_6659);
or U6950 (N_6950,N_6655,N_6685);
and U6951 (N_6951,N_6755,N_6717);
or U6952 (N_6952,N_6708,N_6667);
and U6953 (N_6953,N_6690,N_6754);
xor U6954 (N_6954,N_6788,N_6686);
xor U6955 (N_6955,N_6636,N_6708);
nand U6956 (N_6956,N_6792,N_6788);
or U6957 (N_6957,N_6727,N_6661);
nand U6958 (N_6958,N_6652,N_6797);
xnor U6959 (N_6959,N_6606,N_6681);
or U6960 (N_6960,N_6628,N_6718);
or U6961 (N_6961,N_6736,N_6799);
nand U6962 (N_6962,N_6731,N_6772);
xnor U6963 (N_6963,N_6621,N_6673);
and U6964 (N_6964,N_6688,N_6627);
and U6965 (N_6965,N_6745,N_6731);
or U6966 (N_6966,N_6619,N_6602);
xnor U6967 (N_6967,N_6795,N_6792);
or U6968 (N_6968,N_6684,N_6672);
and U6969 (N_6969,N_6632,N_6793);
xor U6970 (N_6970,N_6771,N_6739);
and U6971 (N_6971,N_6600,N_6703);
and U6972 (N_6972,N_6746,N_6651);
xor U6973 (N_6973,N_6626,N_6796);
and U6974 (N_6974,N_6703,N_6782);
or U6975 (N_6975,N_6616,N_6611);
xnor U6976 (N_6976,N_6710,N_6757);
or U6977 (N_6977,N_6612,N_6609);
or U6978 (N_6978,N_6763,N_6628);
and U6979 (N_6979,N_6799,N_6604);
and U6980 (N_6980,N_6799,N_6694);
xnor U6981 (N_6981,N_6682,N_6640);
or U6982 (N_6982,N_6655,N_6702);
and U6983 (N_6983,N_6711,N_6789);
or U6984 (N_6984,N_6666,N_6771);
and U6985 (N_6985,N_6626,N_6700);
nor U6986 (N_6986,N_6706,N_6733);
nor U6987 (N_6987,N_6615,N_6732);
xor U6988 (N_6988,N_6616,N_6745);
nor U6989 (N_6989,N_6742,N_6738);
xor U6990 (N_6990,N_6704,N_6725);
or U6991 (N_6991,N_6696,N_6629);
or U6992 (N_6992,N_6766,N_6796);
and U6993 (N_6993,N_6795,N_6641);
and U6994 (N_6994,N_6797,N_6752);
nor U6995 (N_6995,N_6658,N_6760);
or U6996 (N_6996,N_6664,N_6602);
or U6997 (N_6997,N_6788,N_6665);
and U6998 (N_6998,N_6791,N_6711);
nor U6999 (N_6999,N_6768,N_6679);
xnor U7000 (N_7000,N_6899,N_6871);
or U7001 (N_7001,N_6810,N_6975);
and U7002 (N_7002,N_6992,N_6894);
nor U7003 (N_7003,N_6932,N_6843);
nor U7004 (N_7004,N_6970,N_6953);
nor U7005 (N_7005,N_6910,N_6919);
xnor U7006 (N_7006,N_6837,N_6951);
xnor U7007 (N_7007,N_6859,N_6920);
xor U7008 (N_7008,N_6940,N_6842);
nor U7009 (N_7009,N_6979,N_6998);
nand U7010 (N_7010,N_6873,N_6972);
xor U7011 (N_7011,N_6862,N_6918);
and U7012 (N_7012,N_6961,N_6808);
nand U7013 (N_7013,N_6895,N_6946);
nor U7014 (N_7014,N_6870,N_6921);
nor U7015 (N_7015,N_6902,N_6849);
xor U7016 (N_7016,N_6876,N_6924);
nor U7017 (N_7017,N_6993,N_6944);
or U7018 (N_7018,N_6957,N_6877);
or U7019 (N_7019,N_6996,N_6826);
and U7020 (N_7020,N_6904,N_6955);
nand U7021 (N_7021,N_6836,N_6860);
and U7022 (N_7022,N_6855,N_6863);
and U7023 (N_7023,N_6880,N_6817);
nand U7024 (N_7024,N_6847,N_6980);
or U7025 (N_7025,N_6867,N_6938);
or U7026 (N_7026,N_6988,N_6890);
nand U7027 (N_7027,N_6911,N_6948);
xnor U7028 (N_7028,N_6884,N_6881);
xnor U7029 (N_7029,N_6845,N_6936);
xor U7030 (N_7030,N_6827,N_6815);
and U7031 (N_7031,N_6858,N_6941);
nand U7032 (N_7032,N_6971,N_6907);
and U7033 (N_7033,N_6829,N_6973);
xnor U7034 (N_7034,N_6925,N_6833);
xor U7035 (N_7035,N_6805,N_6825);
xor U7036 (N_7036,N_6822,N_6802);
or U7037 (N_7037,N_6933,N_6928);
xor U7038 (N_7038,N_6886,N_6875);
or U7039 (N_7039,N_6912,N_6831);
nor U7040 (N_7040,N_6991,N_6964);
and U7041 (N_7041,N_6927,N_6987);
xor U7042 (N_7042,N_6814,N_6995);
or U7043 (N_7043,N_6956,N_6986);
xor U7044 (N_7044,N_6967,N_6950);
nor U7045 (N_7045,N_6968,N_6824);
nor U7046 (N_7046,N_6906,N_6821);
or U7047 (N_7047,N_6931,N_6811);
nor U7048 (N_7048,N_6851,N_6801);
xor U7049 (N_7049,N_6901,N_6848);
and U7050 (N_7050,N_6954,N_6854);
xnor U7051 (N_7051,N_6830,N_6889);
and U7052 (N_7052,N_6838,N_6866);
nor U7053 (N_7053,N_6868,N_6903);
xnor U7054 (N_7054,N_6943,N_6905);
and U7055 (N_7055,N_6909,N_6959);
or U7056 (N_7056,N_6977,N_6828);
and U7057 (N_7057,N_6879,N_6963);
or U7058 (N_7058,N_6929,N_6994);
xor U7059 (N_7059,N_6989,N_6806);
or U7060 (N_7060,N_6878,N_6913);
nand U7061 (N_7061,N_6981,N_6856);
nand U7062 (N_7062,N_6839,N_6804);
or U7063 (N_7063,N_6835,N_6976);
or U7064 (N_7064,N_6897,N_6844);
nand U7065 (N_7065,N_6985,N_6900);
xor U7066 (N_7066,N_6816,N_6893);
or U7067 (N_7067,N_6945,N_6952);
and U7068 (N_7068,N_6869,N_6926);
and U7069 (N_7069,N_6908,N_6803);
nor U7070 (N_7070,N_6984,N_6809);
nor U7071 (N_7071,N_6813,N_6852);
xor U7072 (N_7072,N_6917,N_6960);
and U7073 (N_7073,N_6846,N_6841);
nand U7074 (N_7074,N_6865,N_6883);
nor U7075 (N_7075,N_6914,N_6882);
xnor U7076 (N_7076,N_6888,N_6896);
xnor U7077 (N_7077,N_6978,N_6872);
nor U7078 (N_7078,N_6898,N_6958);
xnor U7079 (N_7079,N_6999,N_6891);
xor U7080 (N_7080,N_6887,N_6937);
nand U7081 (N_7081,N_6922,N_6832);
nand U7082 (N_7082,N_6974,N_6853);
nor U7083 (N_7083,N_6800,N_6861);
xor U7084 (N_7084,N_6812,N_6949);
nor U7085 (N_7085,N_6982,N_6820);
and U7086 (N_7086,N_6823,N_6997);
nand U7087 (N_7087,N_6962,N_6990);
xor U7088 (N_7088,N_6834,N_6930);
xnor U7089 (N_7089,N_6892,N_6965);
xor U7090 (N_7090,N_6850,N_6934);
nor U7091 (N_7091,N_6915,N_6939);
xor U7092 (N_7092,N_6818,N_6885);
nor U7093 (N_7093,N_6916,N_6935);
nand U7094 (N_7094,N_6942,N_6807);
nor U7095 (N_7095,N_6864,N_6874);
nor U7096 (N_7096,N_6857,N_6983);
xor U7097 (N_7097,N_6947,N_6969);
or U7098 (N_7098,N_6819,N_6923);
nand U7099 (N_7099,N_6840,N_6966);
nor U7100 (N_7100,N_6825,N_6965);
and U7101 (N_7101,N_6878,N_6912);
and U7102 (N_7102,N_6927,N_6985);
xnor U7103 (N_7103,N_6866,N_6885);
and U7104 (N_7104,N_6849,N_6856);
xor U7105 (N_7105,N_6915,N_6970);
xnor U7106 (N_7106,N_6837,N_6943);
xor U7107 (N_7107,N_6985,N_6951);
nand U7108 (N_7108,N_6981,N_6809);
and U7109 (N_7109,N_6979,N_6940);
nor U7110 (N_7110,N_6860,N_6914);
xor U7111 (N_7111,N_6806,N_6986);
nand U7112 (N_7112,N_6891,N_6916);
and U7113 (N_7113,N_6971,N_6827);
xor U7114 (N_7114,N_6820,N_6916);
xnor U7115 (N_7115,N_6825,N_6904);
xor U7116 (N_7116,N_6821,N_6999);
or U7117 (N_7117,N_6826,N_6988);
xnor U7118 (N_7118,N_6878,N_6959);
nand U7119 (N_7119,N_6957,N_6813);
nand U7120 (N_7120,N_6976,N_6894);
or U7121 (N_7121,N_6998,N_6853);
nand U7122 (N_7122,N_6868,N_6986);
xnor U7123 (N_7123,N_6911,N_6910);
nand U7124 (N_7124,N_6851,N_6836);
nand U7125 (N_7125,N_6978,N_6972);
nor U7126 (N_7126,N_6946,N_6947);
xor U7127 (N_7127,N_6935,N_6938);
and U7128 (N_7128,N_6972,N_6875);
xnor U7129 (N_7129,N_6866,N_6991);
or U7130 (N_7130,N_6910,N_6938);
nor U7131 (N_7131,N_6925,N_6901);
xnor U7132 (N_7132,N_6825,N_6804);
nand U7133 (N_7133,N_6912,N_6901);
and U7134 (N_7134,N_6824,N_6855);
or U7135 (N_7135,N_6900,N_6869);
xnor U7136 (N_7136,N_6937,N_6915);
and U7137 (N_7137,N_6845,N_6884);
xor U7138 (N_7138,N_6860,N_6837);
xnor U7139 (N_7139,N_6897,N_6847);
nand U7140 (N_7140,N_6900,N_6979);
nor U7141 (N_7141,N_6925,N_6886);
nor U7142 (N_7142,N_6914,N_6884);
xnor U7143 (N_7143,N_6865,N_6815);
xor U7144 (N_7144,N_6854,N_6991);
nand U7145 (N_7145,N_6812,N_6879);
and U7146 (N_7146,N_6975,N_6821);
and U7147 (N_7147,N_6885,N_6858);
nor U7148 (N_7148,N_6909,N_6944);
nand U7149 (N_7149,N_6963,N_6881);
nand U7150 (N_7150,N_6921,N_6937);
or U7151 (N_7151,N_6961,N_6818);
or U7152 (N_7152,N_6999,N_6878);
nand U7153 (N_7153,N_6831,N_6979);
nand U7154 (N_7154,N_6905,N_6945);
and U7155 (N_7155,N_6806,N_6915);
nor U7156 (N_7156,N_6891,N_6990);
nor U7157 (N_7157,N_6834,N_6996);
or U7158 (N_7158,N_6859,N_6956);
and U7159 (N_7159,N_6906,N_6994);
nor U7160 (N_7160,N_6992,N_6967);
and U7161 (N_7161,N_6854,N_6878);
or U7162 (N_7162,N_6851,N_6906);
and U7163 (N_7163,N_6815,N_6810);
or U7164 (N_7164,N_6806,N_6933);
and U7165 (N_7165,N_6951,N_6846);
and U7166 (N_7166,N_6814,N_6942);
nand U7167 (N_7167,N_6852,N_6911);
nand U7168 (N_7168,N_6940,N_6993);
and U7169 (N_7169,N_6925,N_6914);
nor U7170 (N_7170,N_6881,N_6820);
and U7171 (N_7171,N_6881,N_6962);
and U7172 (N_7172,N_6974,N_6832);
and U7173 (N_7173,N_6896,N_6834);
nand U7174 (N_7174,N_6850,N_6893);
and U7175 (N_7175,N_6915,N_6968);
xnor U7176 (N_7176,N_6988,N_6894);
or U7177 (N_7177,N_6967,N_6880);
and U7178 (N_7178,N_6907,N_6896);
and U7179 (N_7179,N_6844,N_6827);
nor U7180 (N_7180,N_6937,N_6861);
or U7181 (N_7181,N_6846,N_6829);
nor U7182 (N_7182,N_6938,N_6965);
xor U7183 (N_7183,N_6888,N_6879);
nand U7184 (N_7184,N_6967,N_6901);
xnor U7185 (N_7185,N_6974,N_6945);
nor U7186 (N_7186,N_6884,N_6873);
and U7187 (N_7187,N_6962,N_6992);
nand U7188 (N_7188,N_6898,N_6853);
xnor U7189 (N_7189,N_6872,N_6995);
or U7190 (N_7190,N_6965,N_6899);
nor U7191 (N_7191,N_6940,N_6883);
or U7192 (N_7192,N_6849,N_6932);
nand U7193 (N_7193,N_6853,N_6818);
xnor U7194 (N_7194,N_6802,N_6895);
xnor U7195 (N_7195,N_6924,N_6872);
nand U7196 (N_7196,N_6842,N_6933);
xnor U7197 (N_7197,N_6808,N_6975);
nand U7198 (N_7198,N_6857,N_6950);
xnor U7199 (N_7199,N_6866,N_6816);
or U7200 (N_7200,N_7086,N_7117);
and U7201 (N_7201,N_7130,N_7078);
nand U7202 (N_7202,N_7102,N_7115);
xor U7203 (N_7203,N_7107,N_7141);
nor U7204 (N_7204,N_7110,N_7177);
nor U7205 (N_7205,N_7093,N_7166);
and U7206 (N_7206,N_7004,N_7082);
nor U7207 (N_7207,N_7173,N_7125);
and U7208 (N_7208,N_7074,N_7135);
nand U7209 (N_7209,N_7094,N_7076);
or U7210 (N_7210,N_7008,N_7099);
nand U7211 (N_7211,N_7030,N_7090);
nand U7212 (N_7212,N_7187,N_7192);
and U7213 (N_7213,N_7118,N_7167);
nor U7214 (N_7214,N_7198,N_7052);
nand U7215 (N_7215,N_7023,N_7010);
nor U7216 (N_7216,N_7084,N_7066);
nand U7217 (N_7217,N_7026,N_7053);
and U7218 (N_7218,N_7028,N_7180);
xor U7219 (N_7219,N_7161,N_7137);
xnor U7220 (N_7220,N_7088,N_7016);
and U7221 (N_7221,N_7001,N_7055);
xor U7222 (N_7222,N_7159,N_7185);
nor U7223 (N_7223,N_7191,N_7059);
xor U7224 (N_7224,N_7062,N_7120);
xor U7225 (N_7225,N_7148,N_7140);
or U7226 (N_7226,N_7119,N_7005);
xnor U7227 (N_7227,N_7064,N_7105);
and U7228 (N_7228,N_7146,N_7077);
xor U7229 (N_7229,N_7024,N_7111);
xnor U7230 (N_7230,N_7170,N_7035);
and U7231 (N_7231,N_7155,N_7020);
and U7232 (N_7232,N_7089,N_7101);
nand U7233 (N_7233,N_7091,N_7129);
and U7234 (N_7234,N_7081,N_7179);
nor U7235 (N_7235,N_7040,N_7065);
nor U7236 (N_7236,N_7070,N_7038);
nand U7237 (N_7237,N_7197,N_7142);
and U7238 (N_7238,N_7048,N_7171);
and U7239 (N_7239,N_7046,N_7156);
nor U7240 (N_7240,N_7182,N_7193);
nor U7241 (N_7241,N_7054,N_7098);
xor U7242 (N_7242,N_7139,N_7196);
or U7243 (N_7243,N_7178,N_7104);
nand U7244 (N_7244,N_7181,N_7083);
xnor U7245 (N_7245,N_7009,N_7061);
xnor U7246 (N_7246,N_7121,N_7163);
nand U7247 (N_7247,N_7122,N_7022);
or U7248 (N_7248,N_7131,N_7034);
xor U7249 (N_7249,N_7186,N_7075);
nand U7250 (N_7250,N_7049,N_7143);
or U7251 (N_7251,N_7013,N_7147);
and U7252 (N_7252,N_7051,N_7073);
nor U7253 (N_7253,N_7144,N_7079);
nor U7254 (N_7254,N_7194,N_7044);
nand U7255 (N_7255,N_7067,N_7095);
nand U7256 (N_7256,N_7056,N_7087);
xor U7257 (N_7257,N_7190,N_7157);
xnor U7258 (N_7258,N_7133,N_7199);
nor U7259 (N_7259,N_7162,N_7006);
or U7260 (N_7260,N_7189,N_7145);
or U7261 (N_7261,N_7195,N_7154);
nor U7262 (N_7262,N_7176,N_7031);
and U7263 (N_7263,N_7114,N_7036);
nor U7264 (N_7264,N_7108,N_7168);
or U7265 (N_7265,N_7175,N_7032);
or U7266 (N_7266,N_7127,N_7136);
and U7267 (N_7267,N_7039,N_7134);
nand U7268 (N_7268,N_7183,N_7007);
xnor U7269 (N_7269,N_7097,N_7164);
or U7270 (N_7270,N_7069,N_7169);
and U7271 (N_7271,N_7126,N_7096);
nor U7272 (N_7272,N_7151,N_7138);
nand U7273 (N_7273,N_7158,N_7050);
or U7274 (N_7274,N_7149,N_7085);
and U7275 (N_7275,N_7058,N_7041);
or U7276 (N_7276,N_7000,N_7172);
or U7277 (N_7277,N_7015,N_7174);
nand U7278 (N_7278,N_7160,N_7021);
nor U7279 (N_7279,N_7152,N_7068);
nand U7280 (N_7280,N_7103,N_7165);
nand U7281 (N_7281,N_7025,N_7042);
and U7282 (N_7282,N_7188,N_7123);
xor U7283 (N_7283,N_7011,N_7113);
nand U7284 (N_7284,N_7150,N_7072);
xor U7285 (N_7285,N_7047,N_7153);
nor U7286 (N_7286,N_7124,N_7043);
xor U7287 (N_7287,N_7029,N_7027);
nand U7288 (N_7288,N_7037,N_7071);
xnor U7289 (N_7289,N_7092,N_7003);
nor U7290 (N_7290,N_7063,N_7002);
nand U7291 (N_7291,N_7109,N_7018);
nand U7292 (N_7292,N_7017,N_7019);
xor U7293 (N_7293,N_7012,N_7100);
nor U7294 (N_7294,N_7184,N_7112);
and U7295 (N_7295,N_7080,N_7014);
and U7296 (N_7296,N_7033,N_7060);
nor U7297 (N_7297,N_7057,N_7132);
or U7298 (N_7298,N_7106,N_7116);
nand U7299 (N_7299,N_7128,N_7045);
nor U7300 (N_7300,N_7060,N_7111);
nor U7301 (N_7301,N_7160,N_7177);
nor U7302 (N_7302,N_7002,N_7066);
or U7303 (N_7303,N_7018,N_7096);
nand U7304 (N_7304,N_7118,N_7036);
nand U7305 (N_7305,N_7117,N_7171);
and U7306 (N_7306,N_7022,N_7159);
nor U7307 (N_7307,N_7016,N_7047);
or U7308 (N_7308,N_7002,N_7106);
xnor U7309 (N_7309,N_7039,N_7073);
and U7310 (N_7310,N_7137,N_7034);
nor U7311 (N_7311,N_7020,N_7163);
nor U7312 (N_7312,N_7017,N_7078);
xnor U7313 (N_7313,N_7184,N_7155);
and U7314 (N_7314,N_7009,N_7075);
nand U7315 (N_7315,N_7065,N_7187);
nor U7316 (N_7316,N_7116,N_7141);
nand U7317 (N_7317,N_7122,N_7177);
or U7318 (N_7318,N_7048,N_7169);
xor U7319 (N_7319,N_7008,N_7095);
xor U7320 (N_7320,N_7192,N_7092);
or U7321 (N_7321,N_7041,N_7136);
nand U7322 (N_7322,N_7197,N_7065);
xnor U7323 (N_7323,N_7048,N_7122);
xnor U7324 (N_7324,N_7097,N_7055);
xnor U7325 (N_7325,N_7058,N_7107);
and U7326 (N_7326,N_7020,N_7116);
or U7327 (N_7327,N_7106,N_7010);
nor U7328 (N_7328,N_7077,N_7153);
xor U7329 (N_7329,N_7124,N_7102);
and U7330 (N_7330,N_7183,N_7124);
xnor U7331 (N_7331,N_7170,N_7188);
nand U7332 (N_7332,N_7003,N_7140);
and U7333 (N_7333,N_7170,N_7051);
and U7334 (N_7334,N_7034,N_7045);
or U7335 (N_7335,N_7062,N_7092);
or U7336 (N_7336,N_7042,N_7145);
nand U7337 (N_7337,N_7098,N_7115);
nor U7338 (N_7338,N_7130,N_7110);
nor U7339 (N_7339,N_7136,N_7163);
and U7340 (N_7340,N_7182,N_7080);
nor U7341 (N_7341,N_7153,N_7113);
nor U7342 (N_7342,N_7041,N_7008);
nor U7343 (N_7343,N_7135,N_7154);
nand U7344 (N_7344,N_7162,N_7149);
or U7345 (N_7345,N_7167,N_7081);
nand U7346 (N_7346,N_7160,N_7145);
nand U7347 (N_7347,N_7144,N_7126);
and U7348 (N_7348,N_7054,N_7067);
xnor U7349 (N_7349,N_7158,N_7151);
xor U7350 (N_7350,N_7170,N_7133);
or U7351 (N_7351,N_7008,N_7001);
nand U7352 (N_7352,N_7137,N_7094);
xor U7353 (N_7353,N_7122,N_7183);
nand U7354 (N_7354,N_7026,N_7165);
nand U7355 (N_7355,N_7115,N_7148);
nor U7356 (N_7356,N_7032,N_7105);
and U7357 (N_7357,N_7039,N_7180);
and U7358 (N_7358,N_7124,N_7128);
nand U7359 (N_7359,N_7194,N_7173);
xor U7360 (N_7360,N_7082,N_7096);
and U7361 (N_7361,N_7116,N_7180);
nor U7362 (N_7362,N_7184,N_7083);
nand U7363 (N_7363,N_7022,N_7127);
or U7364 (N_7364,N_7187,N_7023);
xnor U7365 (N_7365,N_7012,N_7082);
or U7366 (N_7366,N_7104,N_7121);
nor U7367 (N_7367,N_7085,N_7000);
nor U7368 (N_7368,N_7052,N_7094);
or U7369 (N_7369,N_7184,N_7153);
or U7370 (N_7370,N_7135,N_7071);
nand U7371 (N_7371,N_7190,N_7153);
nand U7372 (N_7372,N_7180,N_7037);
nor U7373 (N_7373,N_7189,N_7124);
nand U7374 (N_7374,N_7007,N_7072);
nand U7375 (N_7375,N_7067,N_7061);
nand U7376 (N_7376,N_7136,N_7080);
nand U7377 (N_7377,N_7076,N_7173);
nand U7378 (N_7378,N_7182,N_7082);
and U7379 (N_7379,N_7134,N_7182);
nand U7380 (N_7380,N_7055,N_7017);
xor U7381 (N_7381,N_7111,N_7106);
or U7382 (N_7382,N_7152,N_7008);
and U7383 (N_7383,N_7036,N_7132);
and U7384 (N_7384,N_7079,N_7046);
nand U7385 (N_7385,N_7056,N_7176);
xnor U7386 (N_7386,N_7106,N_7195);
nor U7387 (N_7387,N_7124,N_7098);
nor U7388 (N_7388,N_7021,N_7050);
nor U7389 (N_7389,N_7031,N_7189);
xnor U7390 (N_7390,N_7115,N_7105);
nand U7391 (N_7391,N_7035,N_7101);
nor U7392 (N_7392,N_7053,N_7095);
nor U7393 (N_7393,N_7103,N_7035);
nand U7394 (N_7394,N_7190,N_7132);
nor U7395 (N_7395,N_7048,N_7028);
and U7396 (N_7396,N_7157,N_7137);
or U7397 (N_7397,N_7090,N_7034);
nand U7398 (N_7398,N_7101,N_7153);
nor U7399 (N_7399,N_7083,N_7148);
and U7400 (N_7400,N_7232,N_7200);
nor U7401 (N_7401,N_7266,N_7273);
or U7402 (N_7402,N_7318,N_7315);
and U7403 (N_7403,N_7388,N_7387);
and U7404 (N_7404,N_7209,N_7243);
or U7405 (N_7405,N_7299,N_7220);
and U7406 (N_7406,N_7280,N_7355);
and U7407 (N_7407,N_7398,N_7221);
nor U7408 (N_7408,N_7338,N_7262);
xor U7409 (N_7409,N_7206,N_7389);
and U7410 (N_7410,N_7228,N_7374);
nor U7411 (N_7411,N_7380,N_7247);
nor U7412 (N_7412,N_7361,N_7274);
nand U7413 (N_7413,N_7393,N_7254);
nand U7414 (N_7414,N_7275,N_7351);
and U7415 (N_7415,N_7233,N_7287);
xor U7416 (N_7416,N_7288,N_7252);
and U7417 (N_7417,N_7371,N_7271);
and U7418 (N_7418,N_7353,N_7316);
and U7419 (N_7419,N_7310,N_7330);
nor U7420 (N_7420,N_7261,N_7281);
nor U7421 (N_7421,N_7336,N_7334);
xnor U7422 (N_7422,N_7352,N_7379);
xor U7423 (N_7423,N_7385,N_7240);
and U7424 (N_7424,N_7207,N_7313);
and U7425 (N_7425,N_7296,N_7358);
xnor U7426 (N_7426,N_7203,N_7391);
nand U7427 (N_7427,N_7225,N_7369);
or U7428 (N_7428,N_7293,N_7276);
nor U7429 (N_7429,N_7255,N_7345);
nand U7430 (N_7430,N_7267,N_7249);
nor U7431 (N_7431,N_7308,N_7348);
xnor U7432 (N_7432,N_7363,N_7282);
nand U7433 (N_7433,N_7314,N_7251);
and U7434 (N_7434,N_7223,N_7238);
nand U7435 (N_7435,N_7226,N_7324);
nand U7436 (N_7436,N_7285,N_7272);
or U7437 (N_7437,N_7264,N_7215);
nand U7438 (N_7438,N_7268,N_7214);
nor U7439 (N_7439,N_7202,N_7331);
nor U7440 (N_7440,N_7381,N_7284);
nand U7441 (N_7441,N_7359,N_7392);
or U7442 (N_7442,N_7295,N_7303);
xnor U7443 (N_7443,N_7399,N_7219);
nor U7444 (N_7444,N_7372,N_7269);
nand U7445 (N_7445,N_7257,N_7246);
or U7446 (N_7446,N_7337,N_7395);
or U7447 (N_7447,N_7224,N_7366);
or U7448 (N_7448,N_7213,N_7290);
xor U7449 (N_7449,N_7297,N_7248);
nor U7450 (N_7450,N_7253,N_7367);
nand U7451 (N_7451,N_7218,N_7386);
and U7452 (N_7452,N_7377,N_7364);
and U7453 (N_7453,N_7333,N_7210);
xnor U7454 (N_7454,N_7289,N_7365);
nor U7455 (N_7455,N_7305,N_7394);
nand U7456 (N_7456,N_7217,N_7375);
nor U7457 (N_7457,N_7321,N_7263);
xor U7458 (N_7458,N_7343,N_7292);
and U7459 (N_7459,N_7319,N_7279);
nand U7460 (N_7460,N_7236,N_7328);
and U7461 (N_7461,N_7317,N_7329);
or U7462 (N_7462,N_7384,N_7241);
xor U7463 (N_7463,N_7304,N_7231);
nand U7464 (N_7464,N_7357,N_7309);
nand U7465 (N_7465,N_7346,N_7349);
nand U7466 (N_7466,N_7301,N_7239);
or U7467 (N_7467,N_7307,N_7283);
nor U7468 (N_7468,N_7270,N_7383);
nand U7469 (N_7469,N_7373,N_7370);
xor U7470 (N_7470,N_7312,N_7242);
or U7471 (N_7471,N_7390,N_7212);
xnor U7472 (N_7472,N_7306,N_7347);
xor U7473 (N_7473,N_7234,N_7291);
or U7474 (N_7474,N_7204,N_7201);
nor U7475 (N_7475,N_7211,N_7302);
nand U7476 (N_7476,N_7227,N_7335);
xor U7477 (N_7477,N_7354,N_7286);
xnor U7478 (N_7478,N_7382,N_7360);
nor U7479 (N_7479,N_7294,N_7229);
or U7480 (N_7480,N_7342,N_7356);
nor U7481 (N_7481,N_7244,N_7378);
or U7482 (N_7482,N_7322,N_7320);
xor U7483 (N_7483,N_7300,N_7376);
and U7484 (N_7484,N_7350,N_7237);
and U7485 (N_7485,N_7208,N_7362);
nand U7486 (N_7486,N_7230,N_7258);
or U7487 (N_7487,N_7277,N_7323);
nand U7488 (N_7488,N_7396,N_7397);
and U7489 (N_7489,N_7344,N_7205);
xor U7490 (N_7490,N_7325,N_7216);
or U7491 (N_7491,N_7250,N_7368);
or U7492 (N_7492,N_7311,N_7332);
nor U7493 (N_7493,N_7298,N_7260);
nor U7494 (N_7494,N_7341,N_7256);
and U7495 (N_7495,N_7340,N_7245);
nor U7496 (N_7496,N_7327,N_7259);
and U7497 (N_7497,N_7339,N_7265);
or U7498 (N_7498,N_7235,N_7278);
xor U7499 (N_7499,N_7222,N_7326);
nor U7500 (N_7500,N_7218,N_7316);
and U7501 (N_7501,N_7347,N_7378);
xnor U7502 (N_7502,N_7246,N_7251);
or U7503 (N_7503,N_7389,N_7286);
nand U7504 (N_7504,N_7328,N_7296);
nor U7505 (N_7505,N_7263,N_7277);
and U7506 (N_7506,N_7335,N_7282);
nand U7507 (N_7507,N_7389,N_7291);
xor U7508 (N_7508,N_7258,N_7317);
nor U7509 (N_7509,N_7343,N_7314);
or U7510 (N_7510,N_7395,N_7356);
and U7511 (N_7511,N_7373,N_7221);
and U7512 (N_7512,N_7274,N_7304);
nor U7513 (N_7513,N_7306,N_7328);
nor U7514 (N_7514,N_7227,N_7269);
or U7515 (N_7515,N_7315,N_7336);
or U7516 (N_7516,N_7320,N_7330);
and U7517 (N_7517,N_7216,N_7386);
and U7518 (N_7518,N_7269,N_7383);
xor U7519 (N_7519,N_7247,N_7354);
and U7520 (N_7520,N_7262,N_7388);
or U7521 (N_7521,N_7391,N_7316);
xor U7522 (N_7522,N_7364,N_7329);
nor U7523 (N_7523,N_7376,N_7289);
xnor U7524 (N_7524,N_7213,N_7374);
nor U7525 (N_7525,N_7269,N_7371);
and U7526 (N_7526,N_7316,N_7378);
nand U7527 (N_7527,N_7236,N_7208);
nand U7528 (N_7528,N_7238,N_7326);
and U7529 (N_7529,N_7201,N_7211);
or U7530 (N_7530,N_7388,N_7248);
nor U7531 (N_7531,N_7223,N_7372);
nor U7532 (N_7532,N_7290,N_7204);
nand U7533 (N_7533,N_7397,N_7255);
or U7534 (N_7534,N_7302,N_7337);
or U7535 (N_7535,N_7218,N_7230);
nor U7536 (N_7536,N_7232,N_7264);
or U7537 (N_7537,N_7240,N_7291);
xor U7538 (N_7538,N_7374,N_7398);
nand U7539 (N_7539,N_7200,N_7233);
nand U7540 (N_7540,N_7270,N_7287);
nand U7541 (N_7541,N_7255,N_7358);
nor U7542 (N_7542,N_7336,N_7374);
and U7543 (N_7543,N_7355,N_7267);
nor U7544 (N_7544,N_7217,N_7238);
nor U7545 (N_7545,N_7237,N_7201);
or U7546 (N_7546,N_7300,N_7324);
and U7547 (N_7547,N_7287,N_7343);
nor U7548 (N_7548,N_7265,N_7379);
nand U7549 (N_7549,N_7347,N_7263);
nand U7550 (N_7550,N_7303,N_7257);
or U7551 (N_7551,N_7339,N_7349);
nor U7552 (N_7552,N_7278,N_7216);
nor U7553 (N_7553,N_7307,N_7362);
or U7554 (N_7554,N_7249,N_7285);
and U7555 (N_7555,N_7368,N_7340);
xnor U7556 (N_7556,N_7337,N_7214);
nor U7557 (N_7557,N_7325,N_7215);
xnor U7558 (N_7558,N_7211,N_7392);
or U7559 (N_7559,N_7396,N_7268);
and U7560 (N_7560,N_7254,N_7344);
nor U7561 (N_7561,N_7366,N_7248);
nand U7562 (N_7562,N_7264,N_7351);
xor U7563 (N_7563,N_7322,N_7250);
or U7564 (N_7564,N_7216,N_7306);
xnor U7565 (N_7565,N_7346,N_7290);
and U7566 (N_7566,N_7217,N_7389);
nor U7567 (N_7567,N_7379,N_7338);
xor U7568 (N_7568,N_7378,N_7390);
xor U7569 (N_7569,N_7246,N_7272);
nor U7570 (N_7570,N_7232,N_7219);
nand U7571 (N_7571,N_7269,N_7351);
or U7572 (N_7572,N_7300,N_7283);
nand U7573 (N_7573,N_7207,N_7341);
or U7574 (N_7574,N_7292,N_7271);
nor U7575 (N_7575,N_7331,N_7319);
nor U7576 (N_7576,N_7342,N_7338);
nor U7577 (N_7577,N_7300,N_7239);
nor U7578 (N_7578,N_7335,N_7274);
nor U7579 (N_7579,N_7235,N_7271);
or U7580 (N_7580,N_7280,N_7207);
xnor U7581 (N_7581,N_7223,N_7341);
and U7582 (N_7582,N_7381,N_7299);
or U7583 (N_7583,N_7272,N_7347);
or U7584 (N_7584,N_7281,N_7377);
or U7585 (N_7585,N_7375,N_7379);
nand U7586 (N_7586,N_7364,N_7321);
nor U7587 (N_7587,N_7213,N_7211);
nor U7588 (N_7588,N_7241,N_7330);
or U7589 (N_7589,N_7379,N_7281);
nand U7590 (N_7590,N_7211,N_7271);
nand U7591 (N_7591,N_7278,N_7222);
or U7592 (N_7592,N_7247,N_7364);
nand U7593 (N_7593,N_7378,N_7322);
or U7594 (N_7594,N_7338,N_7294);
nand U7595 (N_7595,N_7261,N_7370);
xor U7596 (N_7596,N_7259,N_7247);
nor U7597 (N_7597,N_7305,N_7376);
nand U7598 (N_7598,N_7390,N_7352);
and U7599 (N_7599,N_7286,N_7262);
and U7600 (N_7600,N_7554,N_7493);
nor U7601 (N_7601,N_7524,N_7407);
or U7602 (N_7602,N_7409,N_7561);
and U7603 (N_7603,N_7544,N_7509);
nor U7604 (N_7604,N_7503,N_7496);
nand U7605 (N_7605,N_7534,N_7430);
nand U7606 (N_7606,N_7596,N_7416);
and U7607 (N_7607,N_7477,N_7460);
xor U7608 (N_7608,N_7568,N_7419);
nand U7609 (N_7609,N_7445,N_7523);
and U7610 (N_7610,N_7589,N_7470);
xor U7611 (N_7611,N_7533,N_7490);
or U7612 (N_7612,N_7482,N_7569);
xor U7613 (N_7613,N_7437,N_7444);
or U7614 (N_7614,N_7473,N_7476);
or U7615 (N_7615,N_7506,N_7462);
nand U7616 (N_7616,N_7467,N_7433);
nor U7617 (N_7617,N_7572,N_7519);
or U7618 (N_7618,N_7406,N_7510);
nor U7619 (N_7619,N_7464,N_7570);
and U7620 (N_7620,N_7483,N_7469);
nand U7621 (N_7621,N_7425,N_7559);
xnor U7622 (N_7622,N_7587,N_7576);
nor U7623 (N_7623,N_7537,N_7441);
and U7624 (N_7624,N_7439,N_7578);
xor U7625 (N_7625,N_7507,N_7586);
or U7626 (N_7626,N_7597,N_7549);
xnor U7627 (N_7627,N_7598,N_7424);
xnor U7628 (N_7628,N_7551,N_7436);
and U7629 (N_7629,N_7417,N_7501);
or U7630 (N_7630,N_7465,N_7508);
or U7631 (N_7631,N_7426,N_7530);
or U7632 (N_7632,N_7573,N_7492);
and U7633 (N_7633,N_7432,N_7491);
or U7634 (N_7634,N_7481,N_7429);
and U7635 (N_7635,N_7498,N_7431);
xnor U7636 (N_7636,N_7427,N_7539);
nor U7637 (N_7637,N_7420,N_7435);
nand U7638 (N_7638,N_7438,N_7457);
nor U7639 (N_7639,N_7422,N_7563);
or U7640 (N_7640,N_7423,N_7562);
nand U7641 (N_7641,N_7455,N_7531);
nor U7642 (N_7642,N_7582,N_7548);
and U7643 (N_7643,N_7487,N_7522);
or U7644 (N_7644,N_7413,N_7564);
nor U7645 (N_7645,N_7471,N_7453);
nand U7646 (N_7646,N_7532,N_7478);
nand U7647 (N_7647,N_7547,N_7517);
or U7648 (N_7648,N_7542,N_7520);
xnor U7649 (N_7649,N_7415,N_7536);
nor U7650 (N_7650,N_7401,N_7412);
xor U7651 (N_7651,N_7553,N_7588);
nor U7652 (N_7652,N_7528,N_7405);
or U7653 (N_7653,N_7583,N_7468);
or U7654 (N_7654,N_7592,N_7514);
and U7655 (N_7655,N_7552,N_7474);
xnor U7656 (N_7656,N_7511,N_7585);
nor U7657 (N_7657,N_7565,N_7489);
or U7658 (N_7658,N_7546,N_7518);
xor U7659 (N_7659,N_7595,N_7408);
nand U7660 (N_7660,N_7504,N_7485);
nand U7661 (N_7661,N_7560,N_7502);
nor U7662 (N_7662,N_7557,N_7590);
xnor U7663 (N_7663,N_7421,N_7512);
nor U7664 (N_7664,N_7410,N_7411);
nor U7665 (N_7665,N_7574,N_7540);
xor U7666 (N_7666,N_7480,N_7494);
nand U7667 (N_7667,N_7486,N_7526);
or U7668 (N_7668,N_7521,N_7525);
and U7669 (N_7669,N_7456,N_7571);
nand U7670 (N_7670,N_7447,N_7529);
nor U7671 (N_7671,N_7575,N_7440);
or U7672 (N_7672,N_7472,N_7599);
nor U7673 (N_7673,N_7400,N_7579);
or U7674 (N_7674,N_7403,N_7558);
and U7675 (N_7675,N_7543,N_7591);
nor U7676 (N_7676,N_7499,N_7449);
nor U7677 (N_7677,N_7545,N_7475);
xnor U7678 (N_7678,N_7567,N_7446);
xor U7679 (N_7679,N_7404,N_7458);
nor U7680 (N_7680,N_7450,N_7555);
nor U7681 (N_7681,N_7556,N_7581);
and U7682 (N_7682,N_7479,N_7488);
or U7683 (N_7683,N_7535,N_7434);
or U7684 (N_7684,N_7428,N_7541);
nor U7685 (N_7685,N_7461,N_7497);
nor U7686 (N_7686,N_7448,N_7495);
or U7687 (N_7687,N_7515,N_7513);
xnor U7688 (N_7688,N_7593,N_7402);
nor U7689 (N_7689,N_7566,N_7580);
nor U7690 (N_7690,N_7442,N_7577);
or U7691 (N_7691,N_7463,N_7484);
or U7692 (N_7692,N_7414,N_7443);
and U7693 (N_7693,N_7516,N_7584);
nor U7694 (N_7694,N_7550,N_7505);
nand U7695 (N_7695,N_7459,N_7451);
or U7696 (N_7696,N_7500,N_7527);
or U7697 (N_7697,N_7418,N_7452);
and U7698 (N_7698,N_7454,N_7538);
xor U7699 (N_7699,N_7466,N_7594);
xnor U7700 (N_7700,N_7496,N_7576);
xnor U7701 (N_7701,N_7428,N_7452);
nand U7702 (N_7702,N_7526,N_7489);
nor U7703 (N_7703,N_7525,N_7504);
nand U7704 (N_7704,N_7470,N_7435);
nor U7705 (N_7705,N_7403,N_7587);
nand U7706 (N_7706,N_7573,N_7424);
or U7707 (N_7707,N_7422,N_7522);
and U7708 (N_7708,N_7467,N_7548);
nor U7709 (N_7709,N_7525,N_7404);
nand U7710 (N_7710,N_7449,N_7571);
nand U7711 (N_7711,N_7593,N_7425);
xor U7712 (N_7712,N_7548,N_7421);
and U7713 (N_7713,N_7430,N_7486);
and U7714 (N_7714,N_7549,N_7560);
or U7715 (N_7715,N_7589,N_7550);
and U7716 (N_7716,N_7572,N_7526);
and U7717 (N_7717,N_7507,N_7517);
xor U7718 (N_7718,N_7509,N_7466);
xnor U7719 (N_7719,N_7530,N_7460);
nor U7720 (N_7720,N_7591,N_7579);
nand U7721 (N_7721,N_7530,N_7592);
nor U7722 (N_7722,N_7478,N_7581);
or U7723 (N_7723,N_7408,N_7549);
nor U7724 (N_7724,N_7444,N_7547);
nor U7725 (N_7725,N_7429,N_7502);
nand U7726 (N_7726,N_7490,N_7488);
and U7727 (N_7727,N_7414,N_7541);
xor U7728 (N_7728,N_7478,N_7534);
xnor U7729 (N_7729,N_7529,N_7435);
xnor U7730 (N_7730,N_7543,N_7498);
nand U7731 (N_7731,N_7527,N_7505);
nand U7732 (N_7732,N_7460,N_7454);
or U7733 (N_7733,N_7452,N_7415);
xnor U7734 (N_7734,N_7463,N_7592);
or U7735 (N_7735,N_7554,N_7480);
xor U7736 (N_7736,N_7497,N_7579);
nor U7737 (N_7737,N_7409,N_7467);
or U7738 (N_7738,N_7508,N_7414);
or U7739 (N_7739,N_7482,N_7423);
or U7740 (N_7740,N_7410,N_7506);
and U7741 (N_7741,N_7518,N_7454);
nor U7742 (N_7742,N_7533,N_7593);
nor U7743 (N_7743,N_7401,N_7530);
and U7744 (N_7744,N_7435,N_7476);
nand U7745 (N_7745,N_7409,N_7404);
and U7746 (N_7746,N_7546,N_7561);
nor U7747 (N_7747,N_7562,N_7482);
and U7748 (N_7748,N_7597,N_7580);
xor U7749 (N_7749,N_7467,N_7560);
nand U7750 (N_7750,N_7525,N_7598);
xor U7751 (N_7751,N_7452,N_7445);
nor U7752 (N_7752,N_7409,N_7509);
and U7753 (N_7753,N_7463,N_7462);
or U7754 (N_7754,N_7474,N_7581);
or U7755 (N_7755,N_7401,N_7400);
or U7756 (N_7756,N_7454,N_7524);
nand U7757 (N_7757,N_7457,N_7444);
nand U7758 (N_7758,N_7475,N_7454);
or U7759 (N_7759,N_7427,N_7505);
nor U7760 (N_7760,N_7463,N_7417);
xor U7761 (N_7761,N_7434,N_7492);
or U7762 (N_7762,N_7534,N_7476);
or U7763 (N_7763,N_7568,N_7405);
nor U7764 (N_7764,N_7506,N_7570);
nand U7765 (N_7765,N_7505,N_7511);
nand U7766 (N_7766,N_7525,N_7508);
nor U7767 (N_7767,N_7487,N_7596);
and U7768 (N_7768,N_7431,N_7587);
or U7769 (N_7769,N_7494,N_7444);
nor U7770 (N_7770,N_7492,N_7414);
or U7771 (N_7771,N_7504,N_7409);
nor U7772 (N_7772,N_7546,N_7572);
nand U7773 (N_7773,N_7450,N_7585);
nand U7774 (N_7774,N_7554,N_7575);
or U7775 (N_7775,N_7468,N_7485);
nand U7776 (N_7776,N_7567,N_7572);
nand U7777 (N_7777,N_7439,N_7597);
xnor U7778 (N_7778,N_7589,N_7516);
and U7779 (N_7779,N_7569,N_7563);
nor U7780 (N_7780,N_7465,N_7567);
xnor U7781 (N_7781,N_7564,N_7443);
nor U7782 (N_7782,N_7512,N_7597);
and U7783 (N_7783,N_7410,N_7433);
and U7784 (N_7784,N_7499,N_7550);
and U7785 (N_7785,N_7582,N_7449);
nand U7786 (N_7786,N_7481,N_7587);
nor U7787 (N_7787,N_7405,N_7461);
or U7788 (N_7788,N_7588,N_7468);
and U7789 (N_7789,N_7584,N_7438);
nand U7790 (N_7790,N_7403,N_7571);
and U7791 (N_7791,N_7513,N_7533);
and U7792 (N_7792,N_7463,N_7460);
nor U7793 (N_7793,N_7404,N_7425);
nand U7794 (N_7794,N_7548,N_7452);
nor U7795 (N_7795,N_7516,N_7474);
nand U7796 (N_7796,N_7493,N_7450);
nor U7797 (N_7797,N_7586,N_7575);
or U7798 (N_7798,N_7540,N_7517);
nand U7799 (N_7799,N_7444,N_7580);
xor U7800 (N_7800,N_7765,N_7756);
xor U7801 (N_7801,N_7707,N_7683);
xor U7802 (N_7802,N_7685,N_7733);
and U7803 (N_7803,N_7672,N_7757);
xnor U7804 (N_7804,N_7729,N_7734);
and U7805 (N_7805,N_7758,N_7721);
or U7806 (N_7806,N_7782,N_7762);
nand U7807 (N_7807,N_7678,N_7657);
and U7808 (N_7808,N_7725,N_7772);
or U7809 (N_7809,N_7670,N_7710);
and U7810 (N_7810,N_7711,N_7748);
xor U7811 (N_7811,N_7664,N_7619);
or U7812 (N_7812,N_7737,N_7776);
nand U7813 (N_7813,N_7736,N_7720);
xor U7814 (N_7814,N_7618,N_7615);
nor U7815 (N_7815,N_7616,N_7724);
xor U7816 (N_7816,N_7605,N_7642);
or U7817 (N_7817,N_7728,N_7699);
xor U7818 (N_7818,N_7676,N_7785);
and U7819 (N_7819,N_7708,N_7744);
xor U7820 (N_7820,N_7633,N_7655);
nor U7821 (N_7821,N_7622,N_7740);
and U7822 (N_7822,N_7671,N_7624);
or U7823 (N_7823,N_7600,N_7726);
nor U7824 (N_7824,N_7639,N_7775);
and U7825 (N_7825,N_7627,N_7634);
and U7826 (N_7826,N_7787,N_7673);
nor U7827 (N_7827,N_7742,N_7743);
or U7828 (N_7828,N_7709,N_7794);
nand U7829 (N_7829,N_7656,N_7735);
nand U7830 (N_7830,N_7768,N_7698);
nand U7831 (N_7831,N_7652,N_7693);
nor U7832 (N_7832,N_7754,N_7688);
or U7833 (N_7833,N_7637,N_7675);
and U7834 (N_7834,N_7704,N_7769);
xnor U7835 (N_7835,N_7774,N_7783);
or U7836 (N_7836,N_7629,N_7695);
and U7837 (N_7837,N_7705,N_7755);
xnor U7838 (N_7838,N_7613,N_7682);
and U7839 (N_7839,N_7749,N_7648);
or U7840 (N_7840,N_7770,N_7674);
and U7841 (N_7841,N_7631,N_7617);
nor U7842 (N_7842,N_7790,N_7692);
and U7843 (N_7843,N_7714,N_7643);
or U7844 (N_7844,N_7786,N_7779);
and U7845 (N_7845,N_7623,N_7793);
nor U7846 (N_7846,N_7750,N_7681);
xnor U7847 (N_7847,N_7628,N_7690);
nand U7848 (N_7848,N_7650,N_7632);
xnor U7849 (N_7849,N_7732,N_7689);
or U7850 (N_7850,N_7646,N_7784);
nand U7851 (N_7851,N_7687,N_7715);
and U7852 (N_7852,N_7649,N_7760);
and U7853 (N_7853,N_7665,N_7752);
nor U7854 (N_7854,N_7700,N_7791);
and U7855 (N_7855,N_7697,N_7792);
nand U7856 (N_7856,N_7799,N_7666);
nor U7857 (N_7857,N_7645,N_7753);
xnor U7858 (N_7858,N_7723,N_7701);
xor U7859 (N_7859,N_7747,N_7761);
xor U7860 (N_7860,N_7612,N_7660);
nand U7861 (N_7861,N_7796,N_7669);
and U7862 (N_7862,N_7778,N_7713);
xnor U7863 (N_7863,N_7731,N_7763);
xor U7864 (N_7864,N_7702,N_7647);
and U7865 (N_7865,N_7626,N_7686);
and U7866 (N_7866,N_7777,N_7625);
nor U7867 (N_7867,N_7767,N_7773);
xnor U7868 (N_7868,N_7780,N_7722);
and U7869 (N_7869,N_7730,N_7653);
nand U7870 (N_7870,N_7659,N_7641);
xnor U7871 (N_7871,N_7604,N_7620);
nor U7872 (N_7872,N_7703,N_7788);
xnor U7873 (N_7873,N_7717,N_7606);
or U7874 (N_7874,N_7798,N_7630);
xor U7875 (N_7875,N_7746,N_7781);
nand U7876 (N_7876,N_7644,N_7667);
or U7877 (N_7877,N_7603,N_7739);
nand U7878 (N_7878,N_7797,N_7759);
nand U7879 (N_7879,N_7694,N_7745);
or U7880 (N_7880,N_7771,N_7795);
xor U7881 (N_7881,N_7663,N_7608);
nand U7882 (N_7882,N_7738,N_7601);
nor U7883 (N_7883,N_7716,N_7712);
nand U7884 (N_7884,N_7621,N_7610);
and U7885 (N_7885,N_7662,N_7602);
or U7886 (N_7886,N_7635,N_7679);
and U7887 (N_7887,N_7609,N_7727);
nor U7888 (N_7888,N_7607,N_7764);
nor U7889 (N_7889,N_7680,N_7751);
or U7890 (N_7890,N_7614,N_7651);
and U7891 (N_7891,N_7696,N_7654);
or U7892 (N_7892,N_7668,N_7789);
and U7893 (N_7893,N_7719,N_7684);
nor U7894 (N_7894,N_7638,N_7706);
or U7895 (N_7895,N_7658,N_7677);
xor U7896 (N_7896,N_7691,N_7718);
and U7897 (N_7897,N_7661,N_7766);
nor U7898 (N_7898,N_7640,N_7636);
and U7899 (N_7899,N_7611,N_7741);
nand U7900 (N_7900,N_7676,N_7796);
nand U7901 (N_7901,N_7689,N_7793);
nand U7902 (N_7902,N_7657,N_7793);
nand U7903 (N_7903,N_7707,N_7664);
or U7904 (N_7904,N_7798,N_7706);
or U7905 (N_7905,N_7706,N_7671);
nor U7906 (N_7906,N_7781,N_7741);
nand U7907 (N_7907,N_7717,N_7794);
xor U7908 (N_7908,N_7637,N_7715);
nor U7909 (N_7909,N_7619,N_7630);
nand U7910 (N_7910,N_7716,N_7634);
nor U7911 (N_7911,N_7642,N_7789);
and U7912 (N_7912,N_7797,N_7616);
xnor U7913 (N_7913,N_7632,N_7628);
nand U7914 (N_7914,N_7681,N_7736);
nand U7915 (N_7915,N_7718,N_7792);
nor U7916 (N_7916,N_7670,N_7600);
nand U7917 (N_7917,N_7698,N_7638);
nor U7918 (N_7918,N_7717,N_7790);
or U7919 (N_7919,N_7766,N_7709);
nand U7920 (N_7920,N_7765,N_7710);
nand U7921 (N_7921,N_7681,N_7757);
nor U7922 (N_7922,N_7606,N_7614);
or U7923 (N_7923,N_7794,N_7789);
or U7924 (N_7924,N_7783,N_7750);
nand U7925 (N_7925,N_7723,N_7761);
or U7926 (N_7926,N_7642,N_7755);
or U7927 (N_7927,N_7749,N_7612);
nand U7928 (N_7928,N_7674,N_7695);
xnor U7929 (N_7929,N_7688,N_7692);
and U7930 (N_7930,N_7681,N_7754);
nor U7931 (N_7931,N_7785,N_7621);
nand U7932 (N_7932,N_7629,N_7650);
or U7933 (N_7933,N_7610,N_7701);
nand U7934 (N_7934,N_7606,N_7783);
xor U7935 (N_7935,N_7792,N_7706);
nor U7936 (N_7936,N_7635,N_7669);
nand U7937 (N_7937,N_7714,N_7604);
xnor U7938 (N_7938,N_7745,N_7674);
nand U7939 (N_7939,N_7799,N_7643);
or U7940 (N_7940,N_7658,N_7739);
nand U7941 (N_7941,N_7763,N_7742);
nand U7942 (N_7942,N_7674,N_7796);
and U7943 (N_7943,N_7739,N_7602);
and U7944 (N_7944,N_7709,N_7705);
nor U7945 (N_7945,N_7730,N_7602);
or U7946 (N_7946,N_7606,N_7796);
nand U7947 (N_7947,N_7699,N_7675);
nand U7948 (N_7948,N_7721,N_7785);
and U7949 (N_7949,N_7729,N_7708);
or U7950 (N_7950,N_7737,N_7712);
and U7951 (N_7951,N_7759,N_7630);
and U7952 (N_7952,N_7762,N_7677);
xnor U7953 (N_7953,N_7696,N_7739);
and U7954 (N_7954,N_7611,N_7785);
or U7955 (N_7955,N_7663,N_7781);
and U7956 (N_7956,N_7646,N_7639);
nor U7957 (N_7957,N_7768,N_7673);
nand U7958 (N_7958,N_7627,N_7677);
nor U7959 (N_7959,N_7693,N_7658);
nor U7960 (N_7960,N_7716,N_7660);
xor U7961 (N_7961,N_7731,N_7661);
nor U7962 (N_7962,N_7667,N_7724);
or U7963 (N_7963,N_7697,N_7728);
nor U7964 (N_7964,N_7755,N_7694);
and U7965 (N_7965,N_7779,N_7605);
nor U7966 (N_7966,N_7749,N_7671);
xnor U7967 (N_7967,N_7701,N_7634);
xnor U7968 (N_7968,N_7721,N_7610);
nor U7969 (N_7969,N_7613,N_7648);
nor U7970 (N_7970,N_7659,N_7782);
xor U7971 (N_7971,N_7616,N_7753);
nand U7972 (N_7972,N_7616,N_7719);
nor U7973 (N_7973,N_7666,N_7761);
or U7974 (N_7974,N_7663,N_7766);
and U7975 (N_7975,N_7677,N_7640);
xnor U7976 (N_7976,N_7780,N_7693);
and U7977 (N_7977,N_7699,N_7724);
nand U7978 (N_7978,N_7736,N_7686);
and U7979 (N_7979,N_7745,N_7634);
and U7980 (N_7980,N_7637,N_7704);
and U7981 (N_7981,N_7770,N_7777);
xor U7982 (N_7982,N_7646,N_7609);
or U7983 (N_7983,N_7777,N_7660);
and U7984 (N_7984,N_7621,N_7736);
nor U7985 (N_7985,N_7779,N_7733);
and U7986 (N_7986,N_7773,N_7629);
nand U7987 (N_7987,N_7790,N_7731);
nand U7988 (N_7988,N_7611,N_7658);
nand U7989 (N_7989,N_7797,N_7738);
nand U7990 (N_7990,N_7632,N_7678);
nand U7991 (N_7991,N_7648,N_7797);
or U7992 (N_7992,N_7668,N_7642);
and U7993 (N_7993,N_7728,N_7724);
nand U7994 (N_7994,N_7702,N_7666);
and U7995 (N_7995,N_7663,N_7768);
nand U7996 (N_7996,N_7603,N_7679);
and U7997 (N_7997,N_7686,N_7723);
nand U7998 (N_7998,N_7606,N_7730);
nor U7999 (N_7999,N_7632,N_7704);
nand U8000 (N_8000,N_7862,N_7863);
or U8001 (N_8001,N_7979,N_7910);
xnor U8002 (N_8002,N_7825,N_7940);
and U8003 (N_8003,N_7885,N_7931);
and U8004 (N_8004,N_7800,N_7982);
or U8005 (N_8005,N_7962,N_7941);
xnor U8006 (N_8006,N_7945,N_7999);
and U8007 (N_8007,N_7967,N_7916);
xnor U8008 (N_8008,N_7832,N_7856);
nand U8009 (N_8009,N_7835,N_7838);
or U8010 (N_8010,N_7874,N_7829);
or U8011 (N_8011,N_7927,N_7840);
or U8012 (N_8012,N_7958,N_7852);
nor U8013 (N_8013,N_7913,N_7834);
and U8014 (N_8014,N_7954,N_7802);
and U8015 (N_8015,N_7892,N_7801);
nand U8016 (N_8016,N_7998,N_7975);
nand U8017 (N_8017,N_7907,N_7837);
and U8018 (N_8018,N_7983,N_7971);
or U8019 (N_8019,N_7974,N_7972);
and U8020 (N_8020,N_7996,N_7928);
and U8021 (N_8021,N_7957,N_7878);
and U8022 (N_8022,N_7803,N_7981);
or U8023 (N_8023,N_7884,N_7893);
or U8024 (N_8024,N_7827,N_7994);
or U8025 (N_8025,N_7929,N_7897);
nand U8026 (N_8026,N_7953,N_7948);
xor U8027 (N_8027,N_7891,N_7848);
or U8028 (N_8028,N_7811,N_7881);
nand U8029 (N_8029,N_7807,N_7944);
xnor U8030 (N_8030,N_7993,N_7877);
nor U8031 (N_8031,N_7926,N_7858);
nor U8032 (N_8032,N_7809,N_7896);
and U8033 (N_8033,N_7933,N_7966);
or U8034 (N_8034,N_7826,N_7908);
or U8035 (N_8035,N_7960,N_7831);
nor U8036 (N_8036,N_7860,N_7869);
xor U8037 (N_8037,N_7977,N_7894);
nor U8038 (N_8038,N_7816,N_7871);
or U8039 (N_8039,N_7951,N_7905);
nand U8040 (N_8040,N_7854,N_7855);
xor U8041 (N_8041,N_7989,N_7900);
or U8042 (N_8042,N_7880,N_7812);
xor U8043 (N_8043,N_7901,N_7959);
or U8044 (N_8044,N_7818,N_7919);
or U8045 (N_8045,N_7946,N_7875);
xor U8046 (N_8046,N_7925,N_7845);
or U8047 (N_8047,N_7824,N_7970);
or U8048 (N_8048,N_7984,N_7911);
xnor U8049 (N_8049,N_7922,N_7844);
and U8050 (N_8050,N_7805,N_7868);
nand U8051 (N_8051,N_7904,N_7853);
nand U8052 (N_8052,N_7997,N_7899);
xnor U8053 (N_8053,N_7846,N_7980);
and U8054 (N_8054,N_7976,N_7820);
and U8055 (N_8055,N_7986,N_7806);
or U8056 (N_8056,N_7920,N_7849);
nor U8057 (N_8057,N_7851,N_7902);
xor U8058 (N_8058,N_7867,N_7889);
and U8059 (N_8059,N_7859,N_7847);
nor U8060 (N_8060,N_7833,N_7823);
nand U8061 (N_8061,N_7836,N_7898);
nor U8062 (N_8062,N_7879,N_7808);
and U8063 (N_8063,N_7887,N_7864);
xnor U8064 (N_8064,N_7850,N_7906);
xor U8065 (N_8065,N_7950,N_7828);
or U8066 (N_8066,N_7866,N_7861);
or U8067 (N_8067,N_7949,N_7810);
nand U8068 (N_8068,N_7990,N_7963);
xor U8069 (N_8069,N_7842,N_7924);
and U8070 (N_8070,N_7938,N_7964);
or U8071 (N_8071,N_7886,N_7813);
nand U8072 (N_8072,N_7985,N_7955);
and U8073 (N_8073,N_7839,N_7921);
and U8074 (N_8074,N_7988,N_7915);
or U8075 (N_8075,N_7969,N_7873);
and U8076 (N_8076,N_7817,N_7947);
xor U8077 (N_8077,N_7987,N_7943);
or U8078 (N_8078,N_7934,N_7843);
nand U8079 (N_8079,N_7952,N_7923);
or U8080 (N_8080,N_7822,N_7882);
xnor U8081 (N_8081,N_7909,N_7841);
nor U8082 (N_8082,N_7895,N_7872);
or U8083 (N_8083,N_7939,N_7956);
or U8084 (N_8084,N_7821,N_7888);
nand U8085 (N_8085,N_7914,N_7936);
xnor U8086 (N_8086,N_7965,N_7992);
and U8087 (N_8087,N_7890,N_7814);
nor U8088 (N_8088,N_7968,N_7961);
and U8089 (N_8089,N_7991,N_7930);
and U8090 (N_8090,N_7973,N_7815);
nand U8091 (N_8091,N_7935,N_7883);
or U8092 (N_8092,N_7937,N_7830);
nand U8093 (N_8093,N_7995,N_7865);
nand U8094 (N_8094,N_7819,N_7942);
xor U8095 (N_8095,N_7876,N_7918);
nor U8096 (N_8096,N_7870,N_7932);
and U8097 (N_8097,N_7857,N_7978);
or U8098 (N_8098,N_7804,N_7903);
or U8099 (N_8099,N_7917,N_7912);
xnor U8100 (N_8100,N_7925,N_7804);
xnor U8101 (N_8101,N_7969,N_7935);
xnor U8102 (N_8102,N_7871,N_7933);
nor U8103 (N_8103,N_7982,N_7821);
or U8104 (N_8104,N_7929,N_7862);
or U8105 (N_8105,N_7883,N_7893);
xnor U8106 (N_8106,N_7887,N_7942);
xnor U8107 (N_8107,N_7876,N_7890);
nor U8108 (N_8108,N_7836,N_7935);
xor U8109 (N_8109,N_7806,N_7800);
nand U8110 (N_8110,N_7970,N_7889);
nand U8111 (N_8111,N_7970,N_7884);
nand U8112 (N_8112,N_7988,N_7845);
and U8113 (N_8113,N_7894,N_7989);
nor U8114 (N_8114,N_7833,N_7927);
or U8115 (N_8115,N_7945,N_7917);
and U8116 (N_8116,N_7912,N_7981);
nand U8117 (N_8117,N_7853,N_7825);
xnor U8118 (N_8118,N_7863,N_7946);
and U8119 (N_8119,N_7933,N_7857);
nand U8120 (N_8120,N_7891,N_7843);
nand U8121 (N_8121,N_7810,N_7956);
or U8122 (N_8122,N_7895,N_7957);
nand U8123 (N_8123,N_7868,N_7827);
nor U8124 (N_8124,N_7806,N_7965);
or U8125 (N_8125,N_7992,N_7877);
xnor U8126 (N_8126,N_7963,N_7906);
xnor U8127 (N_8127,N_7842,N_7921);
nand U8128 (N_8128,N_7801,N_7884);
xor U8129 (N_8129,N_7820,N_7922);
or U8130 (N_8130,N_7858,N_7996);
xor U8131 (N_8131,N_7870,N_7824);
and U8132 (N_8132,N_7873,N_7986);
nor U8133 (N_8133,N_7821,N_7956);
nand U8134 (N_8134,N_7811,N_7977);
nand U8135 (N_8135,N_7895,N_7877);
nor U8136 (N_8136,N_7878,N_7851);
nor U8137 (N_8137,N_7974,N_7851);
and U8138 (N_8138,N_7993,N_7854);
or U8139 (N_8139,N_7808,N_7967);
and U8140 (N_8140,N_7824,N_7832);
or U8141 (N_8141,N_7810,N_7804);
and U8142 (N_8142,N_7838,N_7960);
nand U8143 (N_8143,N_7823,N_7839);
nand U8144 (N_8144,N_7808,N_7826);
and U8145 (N_8145,N_7814,N_7958);
nand U8146 (N_8146,N_7848,N_7828);
or U8147 (N_8147,N_7924,N_7832);
nor U8148 (N_8148,N_7865,N_7960);
or U8149 (N_8149,N_7906,N_7863);
xnor U8150 (N_8150,N_7844,N_7983);
nand U8151 (N_8151,N_7959,N_7864);
and U8152 (N_8152,N_7998,N_7867);
nor U8153 (N_8153,N_7955,N_7883);
or U8154 (N_8154,N_7974,N_7906);
or U8155 (N_8155,N_7924,N_7962);
xnor U8156 (N_8156,N_7983,N_7875);
and U8157 (N_8157,N_7963,N_7991);
xnor U8158 (N_8158,N_7875,N_7955);
nand U8159 (N_8159,N_7878,N_7869);
nand U8160 (N_8160,N_7848,N_7837);
xor U8161 (N_8161,N_7922,N_7803);
or U8162 (N_8162,N_7892,N_7906);
and U8163 (N_8163,N_7806,N_7955);
or U8164 (N_8164,N_7843,N_7894);
nor U8165 (N_8165,N_7918,N_7980);
xor U8166 (N_8166,N_7850,N_7891);
or U8167 (N_8167,N_7888,N_7856);
and U8168 (N_8168,N_7838,N_7903);
xnor U8169 (N_8169,N_7823,N_7933);
nor U8170 (N_8170,N_7835,N_7941);
and U8171 (N_8171,N_7975,N_7977);
xnor U8172 (N_8172,N_7962,N_7925);
and U8173 (N_8173,N_7961,N_7837);
and U8174 (N_8174,N_7878,N_7800);
nand U8175 (N_8175,N_7942,N_7855);
or U8176 (N_8176,N_7859,N_7939);
nand U8177 (N_8177,N_7834,N_7924);
and U8178 (N_8178,N_7877,N_7976);
and U8179 (N_8179,N_7833,N_7940);
and U8180 (N_8180,N_7811,N_7866);
xnor U8181 (N_8181,N_7904,N_7973);
xor U8182 (N_8182,N_7990,N_7861);
nand U8183 (N_8183,N_7854,N_7878);
nor U8184 (N_8184,N_7875,N_7862);
xor U8185 (N_8185,N_7835,N_7883);
or U8186 (N_8186,N_7952,N_7880);
xnor U8187 (N_8187,N_7903,N_7972);
xnor U8188 (N_8188,N_7916,N_7935);
or U8189 (N_8189,N_7806,N_7856);
nand U8190 (N_8190,N_7943,N_7812);
xnor U8191 (N_8191,N_7849,N_7895);
or U8192 (N_8192,N_7875,N_7887);
and U8193 (N_8193,N_7918,N_7810);
xnor U8194 (N_8194,N_7913,N_7937);
nand U8195 (N_8195,N_7826,N_7910);
and U8196 (N_8196,N_7913,N_7954);
nand U8197 (N_8197,N_7876,N_7951);
nand U8198 (N_8198,N_7879,N_7939);
and U8199 (N_8199,N_7980,N_7861);
or U8200 (N_8200,N_8179,N_8129);
and U8201 (N_8201,N_8163,N_8116);
and U8202 (N_8202,N_8151,N_8166);
and U8203 (N_8203,N_8100,N_8128);
nand U8204 (N_8204,N_8119,N_8037);
nor U8205 (N_8205,N_8124,N_8141);
and U8206 (N_8206,N_8011,N_8149);
and U8207 (N_8207,N_8107,N_8028);
nor U8208 (N_8208,N_8016,N_8004);
nor U8209 (N_8209,N_8044,N_8103);
nor U8210 (N_8210,N_8073,N_8019);
and U8211 (N_8211,N_8056,N_8197);
and U8212 (N_8212,N_8130,N_8068);
xor U8213 (N_8213,N_8160,N_8140);
and U8214 (N_8214,N_8136,N_8125);
nor U8215 (N_8215,N_8168,N_8143);
or U8216 (N_8216,N_8185,N_8194);
and U8217 (N_8217,N_8165,N_8075);
nand U8218 (N_8218,N_8024,N_8031);
or U8219 (N_8219,N_8117,N_8034);
or U8220 (N_8220,N_8007,N_8001);
nand U8221 (N_8221,N_8071,N_8155);
or U8222 (N_8222,N_8150,N_8190);
or U8223 (N_8223,N_8181,N_8018);
xnor U8224 (N_8224,N_8041,N_8076);
xor U8225 (N_8225,N_8159,N_8192);
xor U8226 (N_8226,N_8088,N_8000);
or U8227 (N_8227,N_8005,N_8067);
and U8228 (N_8228,N_8058,N_8086);
nand U8229 (N_8229,N_8013,N_8052);
nand U8230 (N_8230,N_8083,N_8180);
nand U8231 (N_8231,N_8137,N_8131);
nor U8232 (N_8232,N_8026,N_8035);
and U8233 (N_8233,N_8081,N_8047);
nand U8234 (N_8234,N_8064,N_8112);
nor U8235 (N_8235,N_8101,N_8142);
nand U8236 (N_8236,N_8033,N_8084);
nand U8237 (N_8237,N_8186,N_8111);
or U8238 (N_8238,N_8030,N_8175);
nand U8239 (N_8239,N_8170,N_8049);
nand U8240 (N_8240,N_8043,N_8147);
xor U8241 (N_8241,N_8182,N_8139);
or U8242 (N_8242,N_8091,N_8072);
or U8243 (N_8243,N_8014,N_8109);
xnor U8244 (N_8244,N_8020,N_8176);
nand U8245 (N_8245,N_8110,N_8187);
or U8246 (N_8246,N_8161,N_8032);
nor U8247 (N_8247,N_8178,N_8177);
nor U8248 (N_8248,N_8120,N_8021);
nand U8249 (N_8249,N_8174,N_8148);
nand U8250 (N_8250,N_8060,N_8118);
xnor U8251 (N_8251,N_8092,N_8055);
and U8252 (N_8252,N_8189,N_8115);
nand U8253 (N_8253,N_8046,N_8054);
nor U8254 (N_8254,N_8114,N_8063);
or U8255 (N_8255,N_8126,N_8123);
or U8256 (N_8256,N_8134,N_8069);
or U8257 (N_8257,N_8015,N_8085);
or U8258 (N_8258,N_8199,N_8006);
xor U8259 (N_8259,N_8195,N_8045);
nand U8260 (N_8260,N_8017,N_8089);
and U8261 (N_8261,N_8051,N_8138);
nor U8262 (N_8262,N_8053,N_8029);
nand U8263 (N_8263,N_8003,N_8087);
or U8264 (N_8264,N_8074,N_8062);
nor U8265 (N_8265,N_8184,N_8162);
and U8266 (N_8266,N_8070,N_8191);
and U8267 (N_8267,N_8121,N_8106);
nand U8268 (N_8268,N_8171,N_8144);
nor U8269 (N_8269,N_8145,N_8152);
xnor U8270 (N_8270,N_8164,N_8036);
nor U8271 (N_8271,N_8048,N_8158);
nand U8272 (N_8272,N_8097,N_8153);
and U8273 (N_8273,N_8057,N_8133);
and U8274 (N_8274,N_8173,N_8094);
nand U8275 (N_8275,N_8113,N_8108);
and U8276 (N_8276,N_8104,N_8132);
and U8277 (N_8277,N_8157,N_8167);
xor U8278 (N_8278,N_8183,N_8154);
nand U8279 (N_8279,N_8009,N_8098);
xor U8280 (N_8280,N_8078,N_8146);
or U8281 (N_8281,N_8065,N_8077);
xor U8282 (N_8282,N_8188,N_8061);
and U8283 (N_8283,N_8039,N_8066);
nor U8284 (N_8284,N_8156,N_8040);
and U8285 (N_8285,N_8012,N_8193);
nand U8286 (N_8286,N_8196,N_8008);
nor U8287 (N_8287,N_8093,N_8080);
xor U8288 (N_8288,N_8102,N_8042);
nand U8289 (N_8289,N_8122,N_8050);
nand U8290 (N_8290,N_8090,N_8079);
nand U8291 (N_8291,N_8025,N_8002);
xor U8292 (N_8292,N_8172,N_8010);
xnor U8293 (N_8293,N_8082,N_8099);
nand U8294 (N_8294,N_8095,N_8169);
xnor U8295 (N_8295,N_8198,N_8105);
xor U8296 (N_8296,N_8096,N_8027);
and U8297 (N_8297,N_8127,N_8022);
and U8298 (N_8298,N_8038,N_8023);
and U8299 (N_8299,N_8135,N_8059);
or U8300 (N_8300,N_8007,N_8166);
or U8301 (N_8301,N_8091,N_8143);
nand U8302 (N_8302,N_8122,N_8164);
xor U8303 (N_8303,N_8040,N_8159);
xnor U8304 (N_8304,N_8031,N_8177);
nor U8305 (N_8305,N_8050,N_8061);
nor U8306 (N_8306,N_8103,N_8040);
nor U8307 (N_8307,N_8153,N_8025);
or U8308 (N_8308,N_8083,N_8015);
and U8309 (N_8309,N_8100,N_8060);
or U8310 (N_8310,N_8054,N_8081);
nor U8311 (N_8311,N_8077,N_8124);
and U8312 (N_8312,N_8016,N_8098);
or U8313 (N_8313,N_8089,N_8157);
nor U8314 (N_8314,N_8142,N_8093);
and U8315 (N_8315,N_8065,N_8192);
or U8316 (N_8316,N_8156,N_8010);
or U8317 (N_8317,N_8099,N_8141);
nand U8318 (N_8318,N_8152,N_8012);
and U8319 (N_8319,N_8020,N_8050);
xnor U8320 (N_8320,N_8069,N_8070);
and U8321 (N_8321,N_8196,N_8159);
or U8322 (N_8322,N_8050,N_8036);
xor U8323 (N_8323,N_8157,N_8099);
or U8324 (N_8324,N_8068,N_8003);
nor U8325 (N_8325,N_8178,N_8023);
or U8326 (N_8326,N_8161,N_8106);
nor U8327 (N_8327,N_8113,N_8111);
nand U8328 (N_8328,N_8195,N_8176);
nand U8329 (N_8329,N_8112,N_8015);
or U8330 (N_8330,N_8170,N_8088);
and U8331 (N_8331,N_8188,N_8173);
and U8332 (N_8332,N_8142,N_8177);
xnor U8333 (N_8333,N_8074,N_8106);
and U8334 (N_8334,N_8017,N_8090);
and U8335 (N_8335,N_8170,N_8092);
nor U8336 (N_8336,N_8100,N_8075);
or U8337 (N_8337,N_8157,N_8037);
nor U8338 (N_8338,N_8104,N_8041);
nor U8339 (N_8339,N_8183,N_8138);
nor U8340 (N_8340,N_8019,N_8107);
xor U8341 (N_8341,N_8096,N_8073);
nor U8342 (N_8342,N_8118,N_8189);
or U8343 (N_8343,N_8043,N_8167);
and U8344 (N_8344,N_8111,N_8136);
or U8345 (N_8345,N_8151,N_8152);
nand U8346 (N_8346,N_8107,N_8175);
xnor U8347 (N_8347,N_8008,N_8083);
or U8348 (N_8348,N_8120,N_8129);
or U8349 (N_8349,N_8099,N_8123);
and U8350 (N_8350,N_8184,N_8012);
or U8351 (N_8351,N_8132,N_8114);
nand U8352 (N_8352,N_8167,N_8086);
nand U8353 (N_8353,N_8096,N_8028);
and U8354 (N_8354,N_8196,N_8176);
nand U8355 (N_8355,N_8149,N_8164);
xor U8356 (N_8356,N_8065,N_8157);
xor U8357 (N_8357,N_8119,N_8066);
nand U8358 (N_8358,N_8194,N_8163);
nor U8359 (N_8359,N_8190,N_8001);
nor U8360 (N_8360,N_8032,N_8141);
nor U8361 (N_8361,N_8021,N_8181);
xnor U8362 (N_8362,N_8032,N_8014);
or U8363 (N_8363,N_8106,N_8042);
nand U8364 (N_8364,N_8080,N_8180);
and U8365 (N_8365,N_8014,N_8163);
nor U8366 (N_8366,N_8112,N_8018);
nand U8367 (N_8367,N_8069,N_8049);
xnor U8368 (N_8368,N_8071,N_8103);
nor U8369 (N_8369,N_8163,N_8142);
and U8370 (N_8370,N_8135,N_8010);
xor U8371 (N_8371,N_8018,N_8019);
xnor U8372 (N_8372,N_8063,N_8181);
nor U8373 (N_8373,N_8033,N_8139);
nor U8374 (N_8374,N_8190,N_8080);
xor U8375 (N_8375,N_8163,N_8050);
xor U8376 (N_8376,N_8066,N_8128);
xor U8377 (N_8377,N_8148,N_8193);
xnor U8378 (N_8378,N_8140,N_8147);
nor U8379 (N_8379,N_8183,N_8089);
and U8380 (N_8380,N_8143,N_8135);
nand U8381 (N_8381,N_8012,N_8146);
and U8382 (N_8382,N_8179,N_8133);
nand U8383 (N_8383,N_8151,N_8096);
nand U8384 (N_8384,N_8115,N_8187);
nand U8385 (N_8385,N_8177,N_8076);
nand U8386 (N_8386,N_8095,N_8036);
nand U8387 (N_8387,N_8199,N_8184);
xnor U8388 (N_8388,N_8190,N_8144);
nand U8389 (N_8389,N_8067,N_8183);
or U8390 (N_8390,N_8113,N_8018);
nand U8391 (N_8391,N_8101,N_8172);
or U8392 (N_8392,N_8146,N_8154);
nor U8393 (N_8393,N_8162,N_8066);
and U8394 (N_8394,N_8104,N_8030);
nand U8395 (N_8395,N_8175,N_8002);
xor U8396 (N_8396,N_8156,N_8021);
or U8397 (N_8397,N_8117,N_8168);
nand U8398 (N_8398,N_8178,N_8067);
nand U8399 (N_8399,N_8061,N_8027);
nor U8400 (N_8400,N_8314,N_8323);
nand U8401 (N_8401,N_8372,N_8344);
nor U8402 (N_8402,N_8378,N_8292);
and U8403 (N_8403,N_8346,N_8353);
nor U8404 (N_8404,N_8262,N_8270);
xor U8405 (N_8405,N_8399,N_8200);
or U8406 (N_8406,N_8364,N_8218);
or U8407 (N_8407,N_8361,N_8360);
or U8408 (N_8408,N_8391,N_8311);
and U8409 (N_8409,N_8339,N_8351);
and U8410 (N_8410,N_8374,N_8260);
and U8411 (N_8411,N_8219,N_8377);
and U8412 (N_8412,N_8368,N_8301);
nand U8413 (N_8413,N_8261,N_8388);
xor U8414 (N_8414,N_8296,N_8357);
and U8415 (N_8415,N_8225,N_8303);
xor U8416 (N_8416,N_8216,N_8226);
and U8417 (N_8417,N_8386,N_8389);
nand U8418 (N_8418,N_8204,N_8205);
or U8419 (N_8419,N_8355,N_8217);
nand U8420 (N_8420,N_8288,N_8320);
nor U8421 (N_8421,N_8274,N_8245);
nand U8422 (N_8422,N_8327,N_8359);
nor U8423 (N_8423,N_8330,N_8257);
xnor U8424 (N_8424,N_8304,N_8211);
and U8425 (N_8425,N_8318,N_8209);
nor U8426 (N_8426,N_8390,N_8367);
nand U8427 (N_8427,N_8221,N_8309);
nor U8428 (N_8428,N_8233,N_8242);
xor U8429 (N_8429,N_8232,N_8237);
xnor U8430 (N_8430,N_8281,N_8235);
xor U8431 (N_8431,N_8285,N_8278);
or U8432 (N_8432,N_8250,N_8263);
and U8433 (N_8433,N_8380,N_8238);
xor U8434 (N_8434,N_8315,N_8295);
nor U8435 (N_8435,N_8332,N_8207);
or U8436 (N_8436,N_8326,N_8338);
nand U8437 (N_8437,N_8383,N_8275);
or U8438 (N_8438,N_8271,N_8228);
xor U8439 (N_8439,N_8306,N_8329);
nor U8440 (N_8440,N_8243,N_8231);
xnor U8441 (N_8441,N_8259,N_8279);
or U8442 (N_8442,N_8381,N_8253);
nand U8443 (N_8443,N_8206,N_8387);
nor U8444 (N_8444,N_8308,N_8341);
xor U8445 (N_8445,N_8283,N_8310);
or U8446 (N_8446,N_8297,N_8363);
and U8447 (N_8447,N_8299,N_8294);
nand U8448 (N_8448,N_8258,N_8349);
and U8449 (N_8449,N_8316,N_8289);
or U8450 (N_8450,N_8254,N_8203);
nor U8451 (N_8451,N_8234,N_8334);
and U8452 (N_8452,N_8291,N_8215);
and U8453 (N_8453,N_8331,N_8251);
and U8454 (N_8454,N_8264,N_8246);
nand U8455 (N_8455,N_8300,N_8248);
and U8456 (N_8456,N_8220,N_8328);
nand U8457 (N_8457,N_8385,N_8373);
xnor U8458 (N_8458,N_8350,N_8201);
and U8459 (N_8459,N_8394,N_8336);
nor U8460 (N_8460,N_8324,N_8282);
and U8461 (N_8461,N_8256,N_8398);
and U8462 (N_8462,N_8319,N_8348);
xnor U8463 (N_8463,N_8210,N_8236);
nand U8464 (N_8464,N_8290,N_8396);
and U8465 (N_8465,N_8202,N_8272);
and U8466 (N_8466,N_8268,N_8375);
and U8467 (N_8467,N_8392,N_8347);
nand U8468 (N_8468,N_8342,N_8255);
nor U8469 (N_8469,N_8273,N_8277);
and U8470 (N_8470,N_8365,N_8333);
nand U8471 (N_8471,N_8239,N_8269);
nor U8472 (N_8472,N_8240,N_8312);
or U8473 (N_8473,N_8343,N_8358);
nor U8474 (N_8474,N_8340,N_8214);
nand U8475 (N_8475,N_8395,N_8213);
and U8476 (N_8476,N_8335,N_8287);
or U8477 (N_8477,N_8230,N_8252);
and U8478 (N_8478,N_8227,N_8371);
or U8479 (N_8479,N_8325,N_8223);
xor U8480 (N_8480,N_8298,N_8352);
nor U8481 (N_8481,N_8313,N_8305);
or U8482 (N_8482,N_8345,N_8247);
nand U8483 (N_8483,N_8307,N_8302);
or U8484 (N_8484,N_8265,N_8241);
and U8485 (N_8485,N_8370,N_8397);
or U8486 (N_8486,N_8224,N_8376);
or U8487 (N_8487,N_8244,N_8384);
nor U8488 (N_8488,N_8293,N_8354);
nor U8489 (N_8489,N_8280,N_8321);
and U8490 (N_8490,N_8369,N_8337);
nand U8491 (N_8491,N_8356,N_8379);
or U8492 (N_8492,N_8229,N_8222);
or U8493 (N_8493,N_8208,N_8284);
nand U8494 (N_8494,N_8212,N_8266);
nand U8495 (N_8495,N_8267,N_8276);
nand U8496 (N_8496,N_8249,N_8317);
nand U8497 (N_8497,N_8362,N_8322);
nor U8498 (N_8498,N_8286,N_8366);
nor U8499 (N_8499,N_8382,N_8393);
and U8500 (N_8500,N_8217,N_8236);
nor U8501 (N_8501,N_8309,N_8241);
nor U8502 (N_8502,N_8324,N_8221);
nor U8503 (N_8503,N_8219,N_8352);
xnor U8504 (N_8504,N_8316,N_8302);
and U8505 (N_8505,N_8321,N_8276);
and U8506 (N_8506,N_8300,N_8239);
nor U8507 (N_8507,N_8368,N_8326);
nand U8508 (N_8508,N_8253,N_8237);
or U8509 (N_8509,N_8309,N_8393);
xnor U8510 (N_8510,N_8331,N_8349);
or U8511 (N_8511,N_8229,N_8329);
nand U8512 (N_8512,N_8256,N_8253);
nand U8513 (N_8513,N_8237,N_8319);
and U8514 (N_8514,N_8378,N_8299);
or U8515 (N_8515,N_8297,N_8388);
or U8516 (N_8516,N_8213,N_8227);
nor U8517 (N_8517,N_8375,N_8331);
xor U8518 (N_8518,N_8235,N_8218);
and U8519 (N_8519,N_8355,N_8230);
xor U8520 (N_8520,N_8390,N_8389);
nor U8521 (N_8521,N_8293,N_8215);
nor U8522 (N_8522,N_8393,N_8304);
nor U8523 (N_8523,N_8304,N_8394);
nor U8524 (N_8524,N_8319,N_8326);
xnor U8525 (N_8525,N_8253,N_8374);
nand U8526 (N_8526,N_8313,N_8317);
xnor U8527 (N_8527,N_8299,N_8292);
nand U8528 (N_8528,N_8279,N_8251);
nand U8529 (N_8529,N_8271,N_8368);
or U8530 (N_8530,N_8352,N_8337);
nand U8531 (N_8531,N_8260,N_8282);
xnor U8532 (N_8532,N_8315,N_8384);
and U8533 (N_8533,N_8329,N_8395);
xor U8534 (N_8534,N_8282,N_8392);
or U8535 (N_8535,N_8307,N_8299);
xnor U8536 (N_8536,N_8231,N_8219);
nand U8537 (N_8537,N_8396,N_8202);
nor U8538 (N_8538,N_8358,N_8250);
xnor U8539 (N_8539,N_8326,N_8278);
xor U8540 (N_8540,N_8220,N_8382);
and U8541 (N_8541,N_8235,N_8367);
and U8542 (N_8542,N_8344,N_8353);
nor U8543 (N_8543,N_8311,N_8220);
nor U8544 (N_8544,N_8267,N_8257);
nor U8545 (N_8545,N_8397,N_8350);
or U8546 (N_8546,N_8353,N_8241);
nand U8547 (N_8547,N_8304,N_8209);
and U8548 (N_8548,N_8341,N_8217);
xnor U8549 (N_8549,N_8237,N_8335);
or U8550 (N_8550,N_8296,N_8359);
xor U8551 (N_8551,N_8263,N_8324);
nor U8552 (N_8552,N_8222,N_8278);
xor U8553 (N_8553,N_8263,N_8218);
nor U8554 (N_8554,N_8208,N_8291);
nor U8555 (N_8555,N_8372,N_8271);
nor U8556 (N_8556,N_8385,N_8295);
nand U8557 (N_8557,N_8230,N_8338);
nor U8558 (N_8558,N_8204,N_8319);
nand U8559 (N_8559,N_8261,N_8205);
nor U8560 (N_8560,N_8308,N_8368);
and U8561 (N_8561,N_8279,N_8366);
and U8562 (N_8562,N_8238,N_8222);
nor U8563 (N_8563,N_8211,N_8338);
nand U8564 (N_8564,N_8309,N_8346);
nand U8565 (N_8565,N_8213,N_8292);
xnor U8566 (N_8566,N_8262,N_8261);
nand U8567 (N_8567,N_8236,N_8235);
and U8568 (N_8568,N_8341,N_8222);
xor U8569 (N_8569,N_8392,N_8298);
and U8570 (N_8570,N_8320,N_8355);
and U8571 (N_8571,N_8264,N_8398);
or U8572 (N_8572,N_8331,N_8323);
and U8573 (N_8573,N_8267,N_8350);
nand U8574 (N_8574,N_8349,N_8222);
and U8575 (N_8575,N_8362,N_8305);
or U8576 (N_8576,N_8207,N_8375);
and U8577 (N_8577,N_8257,N_8217);
and U8578 (N_8578,N_8275,N_8310);
and U8579 (N_8579,N_8335,N_8354);
and U8580 (N_8580,N_8281,N_8204);
xor U8581 (N_8581,N_8312,N_8344);
xor U8582 (N_8582,N_8343,N_8338);
nand U8583 (N_8583,N_8226,N_8342);
nand U8584 (N_8584,N_8279,N_8376);
xnor U8585 (N_8585,N_8257,N_8225);
nor U8586 (N_8586,N_8204,N_8287);
xor U8587 (N_8587,N_8252,N_8368);
or U8588 (N_8588,N_8254,N_8205);
nor U8589 (N_8589,N_8244,N_8236);
nor U8590 (N_8590,N_8214,N_8375);
and U8591 (N_8591,N_8280,N_8206);
and U8592 (N_8592,N_8378,N_8276);
or U8593 (N_8593,N_8397,N_8203);
nor U8594 (N_8594,N_8340,N_8288);
and U8595 (N_8595,N_8397,N_8239);
and U8596 (N_8596,N_8260,N_8293);
nor U8597 (N_8597,N_8285,N_8368);
or U8598 (N_8598,N_8328,N_8378);
nand U8599 (N_8599,N_8349,N_8242);
nor U8600 (N_8600,N_8425,N_8554);
or U8601 (N_8601,N_8497,N_8501);
and U8602 (N_8602,N_8500,N_8457);
or U8603 (N_8603,N_8506,N_8434);
and U8604 (N_8604,N_8541,N_8507);
xor U8605 (N_8605,N_8558,N_8591);
nor U8606 (N_8606,N_8513,N_8413);
nand U8607 (N_8607,N_8402,N_8551);
and U8608 (N_8608,N_8552,N_8414);
or U8609 (N_8609,N_8480,N_8411);
nor U8610 (N_8610,N_8423,N_8407);
nand U8611 (N_8611,N_8536,N_8589);
xor U8612 (N_8612,N_8486,N_8508);
nand U8613 (N_8613,N_8468,N_8509);
nand U8614 (N_8614,N_8467,N_8475);
nand U8615 (N_8615,N_8473,N_8460);
and U8616 (N_8616,N_8422,N_8531);
or U8617 (N_8617,N_8462,N_8491);
and U8618 (N_8618,N_8489,N_8561);
nand U8619 (N_8619,N_8590,N_8474);
or U8620 (N_8620,N_8446,N_8530);
xor U8621 (N_8621,N_8597,N_8592);
xnor U8622 (N_8622,N_8432,N_8450);
nor U8623 (N_8623,N_8424,N_8463);
and U8624 (N_8624,N_8503,N_8569);
or U8625 (N_8625,N_8499,N_8431);
and U8626 (N_8626,N_8504,N_8576);
nor U8627 (N_8627,N_8459,N_8524);
nand U8628 (N_8628,N_8427,N_8525);
and U8629 (N_8629,N_8581,N_8546);
nor U8630 (N_8630,N_8540,N_8488);
xnor U8631 (N_8631,N_8415,N_8417);
and U8632 (N_8632,N_8485,N_8492);
nand U8633 (N_8633,N_8573,N_8498);
or U8634 (N_8634,N_8555,N_8547);
nor U8635 (N_8635,N_8449,N_8527);
xnor U8636 (N_8636,N_8409,N_8584);
nor U8637 (N_8637,N_8585,N_8443);
nand U8638 (N_8638,N_8571,N_8545);
nand U8639 (N_8639,N_8521,N_8563);
and U8640 (N_8640,N_8448,N_8549);
xor U8641 (N_8641,N_8494,N_8440);
xor U8642 (N_8642,N_8511,N_8428);
or U8643 (N_8643,N_8534,N_8567);
and U8644 (N_8644,N_8582,N_8520);
xor U8645 (N_8645,N_8514,N_8502);
nand U8646 (N_8646,N_8442,N_8532);
nand U8647 (N_8647,N_8518,N_8533);
and U8648 (N_8648,N_8564,N_8483);
and U8649 (N_8649,N_8400,N_8481);
or U8650 (N_8650,N_8416,N_8566);
nand U8651 (N_8651,N_8542,N_8410);
and U8652 (N_8652,N_8444,N_8577);
xnor U8653 (N_8653,N_8505,N_8418);
nand U8654 (N_8654,N_8437,N_8470);
nand U8655 (N_8655,N_8593,N_8478);
xor U8656 (N_8656,N_8512,N_8438);
xnor U8657 (N_8657,N_8515,N_8565);
and U8658 (N_8658,N_8535,N_8430);
or U8659 (N_8659,N_8496,N_8404);
nand U8660 (N_8660,N_8594,N_8465);
or U8661 (N_8661,N_8575,N_8447);
xor U8662 (N_8662,N_8516,N_8445);
and U8663 (N_8663,N_8408,N_8439);
nand U8664 (N_8664,N_8403,N_8586);
and U8665 (N_8665,N_8529,N_8405);
nand U8666 (N_8666,N_8433,N_8487);
nand U8667 (N_8667,N_8557,N_8537);
nor U8668 (N_8668,N_8490,N_8493);
and U8669 (N_8669,N_8596,N_8495);
nand U8670 (N_8670,N_8543,N_8570);
or U8671 (N_8671,N_8560,N_8472);
nor U8672 (N_8672,N_8466,N_8401);
or U8673 (N_8673,N_8484,N_8598);
xor U8674 (N_8674,N_8482,N_8526);
and U8675 (N_8675,N_8538,N_8559);
and U8676 (N_8676,N_8588,N_8455);
and U8677 (N_8677,N_8572,N_8464);
xor U8678 (N_8678,N_8587,N_8579);
xnor U8679 (N_8679,N_8406,N_8469);
nand U8680 (N_8680,N_8441,N_8574);
nand U8681 (N_8681,N_8454,N_8580);
xnor U8682 (N_8682,N_8519,N_8528);
xnor U8683 (N_8683,N_8436,N_8429);
nor U8684 (N_8684,N_8451,N_8578);
xnor U8685 (N_8685,N_8435,N_8419);
xnor U8686 (N_8686,N_8562,N_8426);
nor U8687 (N_8687,N_8522,N_8556);
nor U8688 (N_8688,N_8523,N_8583);
and U8689 (N_8689,N_8595,N_8548);
and U8690 (N_8690,N_8471,N_8599);
nand U8691 (N_8691,N_8477,N_8544);
and U8692 (N_8692,N_8458,N_8456);
nand U8693 (N_8693,N_8568,N_8420);
or U8694 (N_8694,N_8421,N_8550);
nand U8695 (N_8695,N_8412,N_8553);
nor U8696 (N_8696,N_8461,N_8510);
nand U8697 (N_8697,N_8517,N_8452);
xnor U8698 (N_8698,N_8539,N_8479);
xnor U8699 (N_8699,N_8476,N_8453);
or U8700 (N_8700,N_8568,N_8589);
nor U8701 (N_8701,N_8579,N_8403);
nor U8702 (N_8702,N_8495,N_8458);
xnor U8703 (N_8703,N_8520,N_8496);
nor U8704 (N_8704,N_8523,N_8591);
or U8705 (N_8705,N_8561,N_8586);
nor U8706 (N_8706,N_8451,N_8506);
or U8707 (N_8707,N_8554,N_8499);
nor U8708 (N_8708,N_8599,N_8401);
nor U8709 (N_8709,N_8528,N_8417);
xor U8710 (N_8710,N_8450,N_8404);
xnor U8711 (N_8711,N_8473,N_8534);
and U8712 (N_8712,N_8426,N_8466);
nand U8713 (N_8713,N_8541,N_8492);
or U8714 (N_8714,N_8425,N_8512);
nand U8715 (N_8715,N_8504,N_8596);
and U8716 (N_8716,N_8476,N_8466);
or U8717 (N_8717,N_8503,N_8417);
and U8718 (N_8718,N_8599,N_8580);
nand U8719 (N_8719,N_8434,N_8491);
xor U8720 (N_8720,N_8475,N_8458);
xnor U8721 (N_8721,N_8574,N_8440);
nor U8722 (N_8722,N_8548,N_8474);
nand U8723 (N_8723,N_8439,N_8415);
nand U8724 (N_8724,N_8528,N_8461);
nand U8725 (N_8725,N_8417,N_8476);
nor U8726 (N_8726,N_8505,N_8514);
xnor U8727 (N_8727,N_8521,N_8514);
and U8728 (N_8728,N_8513,N_8510);
xor U8729 (N_8729,N_8497,N_8476);
and U8730 (N_8730,N_8456,N_8492);
nor U8731 (N_8731,N_8462,N_8562);
or U8732 (N_8732,N_8567,N_8411);
nand U8733 (N_8733,N_8560,N_8568);
or U8734 (N_8734,N_8581,N_8493);
nand U8735 (N_8735,N_8476,N_8517);
and U8736 (N_8736,N_8403,N_8421);
and U8737 (N_8737,N_8567,N_8522);
xnor U8738 (N_8738,N_8555,N_8495);
or U8739 (N_8739,N_8461,N_8447);
xnor U8740 (N_8740,N_8462,N_8490);
and U8741 (N_8741,N_8578,N_8484);
and U8742 (N_8742,N_8405,N_8457);
nor U8743 (N_8743,N_8523,N_8559);
and U8744 (N_8744,N_8577,N_8561);
nor U8745 (N_8745,N_8573,N_8413);
or U8746 (N_8746,N_8401,N_8486);
or U8747 (N_8747,N_8512,N_8568);
and U8748 (N_8748,N_8432,N_8558);
nand U8749 (N_8749,N_8536,N_8467);
nor U8750 (N_8750,N_8463,N_8419);
nand U8751 (N_8751,N_8421,N_8451);
and U8752 (N_8752,N_8509,N_8472);
nand U8753 (N_8753,N_8598,N_8474);
or U8754 (N_8754,N_8466,N_8564);
nand U8755 (N_8755,N_8467,N_8553);
or U8756 (N_8756,N_8510,N_8465);
and U8757 (N_8757,N_8451,N_8539);
nor U8758 (N_8758,N_8528,N_8591);
nand U8759 (N_8759,N_8541,N_8456);
nor U8760 (N_8760,N_8591,N_8406);
xor U8761 (N_8761,N_8598,N_8445);
nor U8762 (N_8762,N_8419,N_8411);
and U8763 (N_8763,N_8416,N_8550);
xnor U8764 (N_8764,N_8530,N_8549);
and U8765 (N_8765,N_8405,N_8586);
nor U8766 (N_8766,N_8415,N_8452);
or U8767 (N_8767,N_8436,N_8400);
or U8768 (N_8768,N_8452,N_8511);
or U8769 (N_8769,N_8500,N_8431);
or U8770 (N_8770,N_8417,N_8592);
xnor U8771 (N_8771,N_8427,N_8462);
nor U8772 (N_8772,N_8435,N_8553);
nor U8773 (N_8773,N_8446,N_8437);
nor U8774 (N_8774,N_8538,N_8411);
nand U8775 (N_8775,N_8591,N_8451);
nand U8776 (N_8776,N_8531,N_8439);
nor U8777 (N_8777,N_8549,N_8493);
nor U8778 (N_8778,N_8542,N_8593);
or U8779 (N_8779,N_8566,N_8435);
nor U8780 (N_8780,N_8416,N_8498);
xor U8781 (N_8781,N_8583,N_8538);
nand U8782 (N_8782,N_8485,N_8537);
nand U8783 (N_8783,N_8521,N_8493);
nand U8784 (N_8784,N_8435,N_8420);
nor U8785 (N_8785,N_8471,N_8504);
or U8786 (N_8786,N_8450,N_8462);
nand U8787 (N_8787,N_8547,N_8447);
nand U8788 (N_8788,N_8564,N_8431);
nor U8789 (N_8789,N_8428,N_8487);
xor U8790 (N_8790,N_8470,N_8573);
and U8791 (N_8791,N_8573,N_8476);
nand U8792 (N_8792,N_8518,N_8525);
and U8793 (N_8793,N_8569,N_8514);
nor U8794 (N_8794,N_8422,N_8421);
nand U8795 (N_8795,N_8566,N_8494);
or U8796 (N_8796,N_8554,N_8440);
nand U8797 (N_8797,N_8494,N_8584);
or U8798 (N_8798,N_8575,N_8445);
nor U8799 (N_8799,N_8467,N_8583);
xor U8800 (N_8800,N_8740,N_8713);
nor U8801 (N_8801,N_8655,N_8645);
and U8802 (N_8802,N_8635,N_8772);
nand U8803 (N_8803,N_8735,N_8756);
xor U8804 (N_8804,N_8720,N_8656);
nand U8805 (N_8805,N_8642,N_8691);
nor U8806 (N_8806,N_8777,N_8702);
nor U8807 (N_8807,N_8640,N_8705);
or U8808 (N_8808,N_8738,N_8664);
xor U8809 (N_8809,N_8616,N_8725);
xor U8810 (N_8810,N_8753,N_8650);
xor U8811 (N_8811,N_8674,N_8629);
nand U8812 (N_8812,N_8663,N_8763);
xor U8813 (N_8813,N_8697,N_8701);
or U8814 (N_8814,N_8637,N_8641);
and U8815 (N_8815,N_8610,N_8728);
xor U8816 (N_8816,N_8638,N_8647);
xor U8817 (N_8817,N_8631,N_8758);
and U8818 (N_8818,N_8613,N_8748);
xor U8819 (N_8819,N_8709,N_8694);
or U8820 (N_8820,N_8632,N_8741);
and U8821 (N_8821,N_8700,N_8754);
nand U8822 (N_8822,N_8606,N_8743);
xor U8823 (N_8823,N_8770,N_8611);
or U8824 (N_8824,N_8734,N_8752);
xnor U8825 (N_8825,N_8687,N_8727);
xnor U8826 (N_8826,N_8711,N_8786);
and U8827 (N_8827,N_8677,N_8775);
or U8828 (N_8828,N_8757,N_8712);
or U8829 (N_8829,N_8744,N_8685);
or U8830 (N_8830,N_8779,N_8760);
and U8831 (N_8831,N_8612,N_8704);
and U8832 (N_8832,N_8755,N_8733);
and U8833 (N_8833,N_8790,N_8659);
and U8834 (N_8834,N_8710,N_8789);
and U8835 (N_8835,N_8716,N_8771);
xor U8836 (N_8836,N_8633,N_8667);
and U8837 (N_8837,N_8739,N_8676);
or U8838 (N_8838,N_8796,N_8601);
or U8839 (N_8839,N_8722,N_8695);
or U8840 (N_8840,N_8699,N_8785);
or U8841 (N_8841,N_8729,N_8762);
and U8842 (N_8842,N_8609,N_8604);
nor U8843 (N_8843,N_8683,N_8692);
nand U8844 (N_8844,N_8792,N_8723);
xnor U8845 (N_8845,N_8788,N_8780);
xor U8846 (N_8846,N_8634,N_8767);
nand U8847 (N_8847,N_8718,N_8681);
xor U8848 (N_8848,N_8773,N_8736);
xnor U8849 (N_8849,N_8668,N_8665);
nand U8850 (N_8850,N_8628,N_8625);
xor U8851 (N_8851,N_8776,N_8615);
nor U8852 (N_8852,N_8791,N_8660);
or U8853 (N_8853,N_8781,N_8620);
nand U8854 (N_8854,N_8782,N_8795);
or U8855 (N_8855,N_8707,N_8658);
and U8856 (N_8856,N_8602,N_8747);
xnor U8857 (N_8857,N_8666,N_8639);
nand U8858 (N_8858,N_8759,N_8670);
nor U8859 (N_8859,N_8769,N_8689);
or U8860 (N_8860,N_8693,N_8732);
nand U8861 (N_8861,N_8652,N_8717);
and U8862 (N_8862,N_8746,N_8797);
nand U8863 (N_8863,N_8643,N_8799);
xor U8864 (N_8864,N_8731,N_8794);
xor U8865 (N_8865,N_8706,N_8624);
nor U8866 (N_8866,N_8672,N_8646);
nor U8867 (N_8867,N_8793,N_8686);
xnor U8868 (N_8868,N_8688,N_8654);
nor U8869 (N_8869,N_8698,N_8675);
nand U8870 (N_8870,N_8766,N_8648);
xnor U8871 (N_8871,N_8764,N_8607);
xor U8872 (N_8872,N_8798,N_8614);
and U8873 (N_8873,N_8679,N_8630);
or U8874 (N_8874,N_8626,N_8730);
or U8875 (N_8875,N_8708,N_8726);
xor U8876 (N_8876,N_8715,N_8608);
or U8877 (N_8877,N_8605,N_8644);
nor U8878 (N_8878,N_8600,N_8703);
xor U8879 (N_8879,N_8680,N_8742);
or U8880 (N_8880,N_8774,N_8678);
or U8881 (N_8881,N_8719,N_8673);
or U8882 (N_8882,N_8749,N_8669);
nor U8883 (N_8883,N_8783,N_8778);
nand U8884 (N_8884,N_8684,N_8657);
nand U8885 (N_8885,N_8617,N_8721);
and U8886 (N_8886,N_8627,N_8623);
or U8887 (N_8887,N_8750,N_8651);
xnor U8888 (N_8888,N_8603,N_8768);
nor U8889 (N_8889,N_8765,N_8745);
xnor U8890 (N_8890,N_8714,N_8696);
xnor U8891 (N_8891,N_8690,N_8682);
or U8892 (N_8892,N_8671,N_8724);
nand U8893 (N_8893,N_8761,N_8622);
nand U8894 (N_8894,N_8787,N_8653);
and U8895 (N_8895,N_8662,N_8619);
or U8896 (N_8896,N_8661,N_8618);
or U8897 (N_8897,N_8784,N_8737);
or U8898 (N_8898,N_8621,N_8751);
or U8899 (N_8899,N_8636,N_8649);
xor U8900 (N_8900,N_8762,N_8661);
or U8901 (N_8901,N_8644,N_8752);
nand U8902 (N_8902,N_8685,N_8728);
or U8903 (N_8903,N_8679,N_8697);
and U8904 (N_8904,N_8643,N_8777);
nor U8905 (N_8905,N_8605,N_8663);
nor U8906 (N_8906,N_8623,N_8743);
xor U8907 (N_8907,N_8645,N_8697);
nor U8908 (N_8908,N_8605,N_8676);
xnor U8909 (N_8909,N_8779,N_8769);
nand U8910 (N_8910,N_8609,N_8605);
xnor U8911 (N_8911,N_8771,N_8754);
nor U8912 (N_8912,N_8722,N_8631);
nand U8913 (N_8913,N_8640,N_8605);
nor U8914 (N_8914,N_8656,N_8775);
or U8915 (N_8915,N_8627,N_8701);
nand U8916 (N_8916,N_8709,N_8691);
and U8917 (N_8917,N_8733,N_8633);
or U8918 (N_8918,N_8719,N_8648);
nor U8919 (N_8919,N_8670,N_8664);
nor U8920 (N_8920,N_8639,N_8795);
nand U8921 (N_8921,N_8700,N_8657);
nor U8922 (N_8922,N_8668,N_8753);
or U8923 (N_8923,N_8782,N_8623);
xor U8924 (N_8924,N_8789,N_8695);
and U8925 (N_8925,N_8696,N_8649);
xnor U8926 (N_8926,N_8608,N_8796);
nand U8927 (N_8927,N_8739,N_8643);
xnor U8928 (N_8928,N_8651,N_8606);
and U8929 (N_8929,N_8716,N_8780);
nand U8930 (N_8930,N_8644,N_8763);
and U8931 (N_8931,N_8692,N_8738);
and U8932 (N_8932,N_8609,N_8603);
nand U8933 (N_8933,N_8792,N_8766);
and U8934 (N_8934,N_8704,N_8631);
and U8935 (N_8935,N_8647,N_8742);
or U8936 (N_8936,N_8784,N_8691);
and U8937 (N_8937,N_8773,N_8753);
nor U8938 (N_8938,N_8750,N_8773);
or U8939 (N_8939,N_8736,N_8637);
nor U8940 (N_8940,N_8685,N_8734);
nor U8941 (N_8941,N_8690,N_8754);
and U8942 (N_8942,N_8650,N_8639);
nor U8943 (N_8943,N_8698,N_8652);
and U8944 (N_8944,N_8607,N_8659);
nand U8945 (N_8945,N_8613,N_8747);
xor U8946 (N_8946,N_8680,N_8758);
xor U8947 (N_8947,N_8710,N_8788);
nand U8948 (N_8948,N_8752,N_8725);
nor U8949 (N_8949,N_8665,N_8705);
nand U8950 (N_8950,N_8647,N_8789);
nand U8951 (N_8951,N_8671,N_8705);
xnor U8952 (N_8952,N_8736,N_8748);
nor U8953 (N_8953,N_8713,N_8733);
nor U8954 (N_8954,N_8753,N_8758);
nor U8955 (N_8955,N_8771,N_8626);
and U8956 (N_8956,N_8790,N_8766);
nor U8957 (N_8957,N_8699,N_8787);
nand U8958 (N_8958,N_8706,N_8707);
or U8959 (N_8959,N_8679,N_8758);
and U8960 (N_8960,N_8656,N_8664);
or U8961 (N_8961,N_8655,N_8685);
xnor U8962 (N_8962,N_8601,N_8733);
and U8963 (N_8963,N_8603,N_8702);
nor U8964 (N_8964,N_8763,N_8772);
and U8965 (N_8965,N_8742,N_8703);
xor U8966 (N_8966,N_8692,N_8731);
xnor U8967 (N_8967,N_8613,N_8637);
nand U8968 (N_8968,N_8762,N_8784);
and U8969 (N_8969,N_8782,N_8638);
nor U8970 (N_8970,N_8720,N_8626);
nor U8971 (N_8971,N_8674,N_8613);
nor U8972 (N_8972,N_8694,N_8623);
nand U8973 (N_8973,N_8656,N_8708);
nor U8974 (N_8974,N_8781,N_8733);
xor U8975 (N_8975,N_8792,N_8728);
nand U8976 (N_8976,N_8717,N_8613);
and U8977 (N_8977,N_8635,N_8639);
xor U8978 (N_8978,N_8627,N_8775);
and U8979 (N_8979,N_8695,N_8706);
and U8980 (N_8980,N_8762,N_8605);
and U8981 (N_8981,N_8712,N_8636);
or U8982 (N_8982,N_8764,N_8755);
or U8983 (N_8983,N_8794,N_8622);
xor U8984 (N_8984,N_8758,N_8709);
xnor U8985 (N_8985,N_8682,N_8748);
xor U8986 (N_8986,N_8682,N_8717);
and U8987 (N_8987,N_8641,N_8704);
or U8988 (N_8988,N_8700,N_8612);
xnor U8989 (N_8989,N_8688,N_8793);
nand U8990 (N_8990,N_8662,N_8681);
xnor U8991 (N_8991,N_8731,N_8755);
or U8992 (N_8992,N_8798,N_8700);
nor U8993 (N_8993,N_8631,N_8657);
and U8994 (N_8994,N_8764,N_8776);
and U8995 (N_8995,N_8665,N_8681);
nand U8996 (N_8996,N_8766,N_8612);
nor U8997 (N_8997,N_8663,N_8767);
nand U8998 (N_8998,N_8701,N_8606);
nor U8999 (N_8999,N_8671,N_8773);
xnor U9000 (N_9000,N_8928,N_8894);
nor U9001 (N_9001,N_8879,N_8972);
nor U9002 (N_9002,N_8938,N_8874);
nor U9003 (N_9003,N_8968,N_8833);
and U9004 (N_9004,N_8843,N_8876);
nor U9005 (N_9005,N_8808,N_8924);
nor U9006 (N_9006,N_8906,N_8957);
or U9007 (N_9007,N_8918,N_8820);
nand U9008 (N_9008,N_8971,N_8909);
and U9009 (N_9009,N_8884,N_8885);
nor U9010 (N_9010,N_8907,N_8853);
and U9011 (N_9011,N_8966,N_8826);
and U9012 (N_9012,N_8866,N_8806);
nand U9013 (N_9013,N_8814,N_8996);
nand U9014 (N_9014,N_8877,N_8855);
xor U9015 (N_9015,N_8954,N_8913);
xnor U9016 (N_9016,N_8872,N_8847);
or U9017 (N_9017,N_8893,N_8807);
and U9018 (N_9018,N_8922,N_8976);
nor U9019 (N_9019,N_8825,N_8989);
and U9020 (N_9020,N_8811,N_8816);
nor U9021 (N_9021,N_8994,N_8952);
xor U9022 (N_9022,N_8871,N_8870);
nand U9023 (N_9023,N_8956,N_8849);
or U9024 (N_9024,N_8867,N_8882);
and U9025 (N_9025,N_8945,N_8891);
or U9026 (N_9026,N_8995,N_8939);
nand U9027 (N_9027,N_8819,N_8915);
xnor U9028 (N_9028,N_8813,N_8959);
and U9029 (N_9029,N_8979,N_8930);
nand U9030 (N_9030,N_8982,N_8887);
and U9031 (N_9031,N_8969,N_8852);
nor U9032 (N_9032,N_8933,N_8932);
and U9033 (N_9033,N_8821,N_8862);
nor U9034 (N_9034,N_8985,N_8836);
and U9035 (N_9035,N_8993,N_8828);
or U9036 (N_9036,N_8801,N_8898);
or U9037 (N_9037,N_8838,N_8981);
or U9038 (N_9038,N_8953,N_8896);
xnor U9039 (N_9039,N_8992,N_8990);
xor U9040 (N_9040,N_8960,N_8889);
and U9041 (N_9041,N_8958,N_8944);
and U9042 (N_9042,N_8842,N_8840);
xnor U9043 (N_9043,N_8931,N_8991);
nor U9044 (N_9044,N_8817,N_8858);
xnor U9045 (N_9045,N_8947,N_8927);
or U9046 (N_9046,N_8875,N_8926);
nand U9047 (N_9047,N_8940,N_8845);
or U9048 (N_9048,N_8835,N_8805);
xor U9049 (N_9049,N_8834,N_8935);
nor U9050 (N_9050,N_8941,N_8902);
or U9051 (N_9051,N_8897,N_8937);
or U9052 (N_9052,N_8873,N_8934);
xor U9053 (N_9053,N_8854,N_8892);
xor U9054 (N_9054,N_8802,N_8977);
and U9055 (N_9055,N_8949,N_8943);
and U9056 (N_9056,N_8865,N_8839);
and U9057 (N_9057,N_8946,N_8970);
or U9058 (N_9058,N_8963,N_8987);
and U9059 (N_9059,N_8832,N_8905);
and U9060 (N_9060,N_8859,N_8880);
or U9061 (N_9061,N_8851,N_8878);
or U9062 (N_9062,N_8844,N_8864);
and U9063 (N_9063,N_8974,N_8950);
nor U9064 (N_9064,N_8883,N_8923);
nor U9065 (N_9065,N_8964,N_8965);
nor U9066 (N_9066,N_8860,N_8888);
nand U9067 (N_9067,N_8948,N_8986);
nand U9068 (N_9068,N_8978,N_8973);
and U9069 (N_9069,N_8830,N_8929);
or U9070 (N_9070,N_8857,N_8908);
xor U9071 (N_9071,N_8810,N_8856);
nor U9072 (N_9072,N_8812,N_8881);
and U9073 (N_9073,N_8975,N_8967);
nand U9074 (N_9074,N_8921,N_8900);
xor U9075 (N_9075,N_8848,N_8822);
or U9076 (N_9076,N_8868,N_8831);
xor U9077 (N_9077,N_8999,N_8997);
nor U9078 (N_9078,N_8912,N_8818);
nor U9079 (N_9079,N_8829,N_8827);
nand U9080 (N_9080,N_8942,N_8804);
and U9081 (N_9081,N_8988,N_8823);
xnor U9082 (N_9082,N_8850,N_8899);
xnor U9083 (N_9083,N_8951,N_8984);
xnor U9084 (N_9084,N_8936,N_8890);
nor U9085 (N_9085,N_8886,N_8914);
nand U9086 (N_9086,N_8919,N_8809);
xnor U9087 (N_9087,N_8815,N_8916);
and U9088 (N_9088,N_8920,N_8846);
xor U9089 (N_9089,N_8925,N_8955);
nand U9090 (N_9090,N_8962,N_8961);
and U9091 (N_9091,N_8861,N_8910);
nand U9092 (N_9092,N_8904,N_8895);
xnor U9093 (N_9093,N_8980,N_8983);
xnor U9094 (N_9094,N_8903,N_8917);
or U9095 (N_9095,N_8841,N_8998);
nand U9096 (N_9096,N_8869,N_8803);
xnor U9097 (N_9097,N_8800,N_8837);
xor U9098 (N_9098,N_8824,N_8911);
nand U9099 (N_9099,N_8863,N_8901);
or U9100 (N_9100,N_8850,N_8970);
and U9101 (N_9101,N_8837,N_8816);
or U9102 (N_9102,N_8862,N_8878);
xor U9103 (N_9103,N_8927,N_8998);
and U9104 (N_9104,N_8972,N_8980);
nor U9105 (N_9105,N_8875,N_8886);
and U9106 (N_9106,N_8937,N_8976);
xor U9107 (N_9107,N_8831,N_8928);
nor U9108 (N_9108,N_8956,N_8979);
nand U9109 (N_9109,N_8823,N_8804);
nand U9110 (N_9110,N_8998,N_8839);
xor U9111 (N_9111,N_8864,N_8829);
xor U9112 (N_9112,N_8963,N_8854);
nand U9113 (N_9113,N_8811,N_8809);
nor U9114 (N_9114,N_8986,N_8849);
xor U9115 (N_9115,N_8952,N_8884);
nor U9116 (N_9116,N_8813,N_8921);
and U9117 (N_9117,N_8969,N_8978);
nor U9118 (N_9118,N_8885,N_8805);
or U9119 (N_9119,N_8944,N_8997);
nand U9120 (N_9120,N_8827,N_8805);
nand U9121 (N_9121,N_8803,N_8930);
or U9122 (N_9122,N_8848,N_8963);
nand U9123 (N_9123,N_8871,N_8970);
nand U9124 (N_9124,N_8871,N_8899);
nor U9125 (N_9125,N_8933,N_8837);
and U9126 (N_9126,N_8916,N_8809);
nor U9127 (N_9127,N_8842,N_8817);
nand U9128 (N_9128,N_8805,N_8947);
nand U9129 (N_9129,N_8875,N_8830);
nand U9130 (N_9130,N_8922,N_8982);
nor U9131 (N_9131,N_8801,N_8916);
xnor U9132 (N_9132,N_8967,N_8981);
nand U9133 (N_9133,N_8878,N_8875);
or U9134 (N_9134,N_8853,N_8879);
or U9135 (N_9135,N_8840,N_8921);
or U9136 (N_9136,N_8819,N_8858);
nand U9137 (N_9137,N_8961,N_8820);
and U9138 (N_9138,N_8825,N_8901);
and U9139 (N_9139,N_8991,N_8862);
and U9140 (N_9140,N_8931,N_8964);
nor U9141 (N_9141,N_8945,N_8885);
nand U9142 (N_9142,N_8921,N_8997);
nor U9143 (N_9143,N_8925,N_8832);
or U9144 (N_9144,N_8805,N_8936);
nand U9145 (N_9145,N_8935,N_8915);
xnor U9146 (N_9146,N_8902,N_8925);
nand U9147 (N_9147,N_8956,N_8870);
nand U9148 (N_9148,N_8846,N_8922);
nor U9149 (N_9149,N_8812,N_8959);
xnor U9150 (N_9150,N_8966,N_8835);
nor U9151 (N_9151,N_8838,N_8927);
nand U9152 (N_9152,N_8838,N_8961);
nand U9153 (N_9153,N_8915,N_8885);
xnor U9154 (N_9154,N_8898,N_8915);
and U9155 (N_9155,N_8875,N_8946);
xor U9156 (N_9156,N_8912,N_8802);
xor U9157 (N_9157,N_8882,N_8965);
nor U9158 (N_9158,N_8966,N_8909);
nand U9159 (N_9159,N_8975,N_8953);
xor U9160 (N_9160,N_8805,N_8953);
nand U9161 (N_9161,N_8976,N_8845);
nand U9162 (N_9162,N_8979,N_8946);
nor U9163 (N_9163,N_8953,N_8841);
nand U9164 (N_9164,N_8878,N_8810);
and U9165 (N_9165,N_8846,N_8829);
and U9166 (N_9166,N_8882,N_8984);
nor U9167 (N_9167,N_8880,N_8934);
or U9168 (N_9168,N_8896,N_8856);
xnor U9169 (N_9169,N_8833,N_8812);
xnor U9170 (N_9170,N_8982,N_8990);
xnor U9171 (N_9171,N_8914,N_8962);
and U9172 (N_9172,N_8981,N_8848);
or U9173 (N_9173,N_8881,N_8944);
and U9174 (N_9174,N_8979,N_8885);
and U9175 (N_9175,N_8863,N_8924);
or U9176 (N_9176,N_8912,N_8971);
nand U9177 (N_9177,N_8926,N_8957);
and U9178 (N_9178,N_8911,N_8965);
and U9179 (N_9179,N_8952,N_8849);
nand U9180 (N_9180,N_8967,N_8854);
or U9181 (N_9181,N_8859,N_8845);
nand U9182 (N_9182,N_8931,N_8870);
nor U9183 (N_9183,N_8913,N_8965);
or U9184 (N_9184,N_8800,N_8833);
and U9185 (N_9185,N_8892,N_8802);
and U9186 (N_9186,N_8947,N_8819);
or U9187 (N_9187,N_8866,N_8915);
and U9188 (N_9188,N_8980,N_8913);
nand U9189 (N_9189,N_8943,N_8934);
or U9190 (N_9190,N_8959,N_8926);
nand U9191 (N_9191,N_8810,N_8916);
nor U9192 (N_9192,N_8989,N_8945);
nand U9193 (N_9193,N_8813,N_8906);
nor U9194 (N_9194,N_8850,N_8861);
or U9195 (N_9195,N_8974,N_8867);
xor U9196 (N_9196,N_8981,N_8951);
or U9197 (N_9197,N_8911,N_8871);
xor U9198 (N_9198,N_8984,N_8801);
and U9199 (N_9199,N_8999,N_8965);
nand U9200 (N_9200,N_9181,N_9005);
nor U9201 (N_9201,N_9179,N_9155);
and U9202 (N_9202,N_9017,N_9031);
and U9203 (N_9203,N_9089,N_9189);
nor U9204 (N_9204,N_9078,N_9093);
and U9205 (N_9205,N_9166,N_9053);
nor U9206 (N_9206,N_9185,N_9020);
xor U9207 (N_9207,N_9000,N_9038);
xnor U9208 (N_9208,N_9195,N_9150);
nand U9209 (N_9209,N_9070,N_9036);
or U9210 (N_9210,N_9127,N_9001);
nor U9211 (N_9211,N_9123,N_9035);
xnor U9212 (N_9212,N_9197,N_9033);
xor U9213 (N_9213,N_9016,N_9113);
nand U9214 (N_9214,N_9096,N_9061);
nand U9215 (N_9215,N_9073,N_9129);
xnor U9216 (N_9216,N_9182,N_9046);
nand U9217 (N_9217,N_9173,N_9190);
nand U9218 (N_9218,N_9074,N_9007);
xor U9219 (N_9219,N_9135,N_9076);
nor U9220 (N_9220,N_9171,N_9006);
and U9221 (N_9221,N_9002,N_9041);
or U9222 (N_9222,N_9065,N_9178);
nor U9223 (N_9223,N_9130,N_9092);
and U9224 (N_9224,N_9163,N_9151);
or U9225 (N_9225,N_9160,N_9121);
or U9226 (N_9226,N_9167,N_9013);
or U9227 (N_9227,N_9192,N_9146);
nor U9228 (N_9228,N_9148,N_9102);
and U9229 (N_9229,N_9100,N_9083);
xnor U9230 (N_9230,N_9153,N_9091);
or U9231 (N_9231,N_9126,N_9060);
and U9232 (N_9232,N_9198,N_9186);
nand U9233 (N_9233,N_9169,N_9072);
nand U9234 (N_9234,N_9047,N_9177);
nor U9235 (N_9235,N_9018,N_9188);
or U9236 (N_9236,N_9012,N_9042);
xor U9237 (N_9237,N_9176,N_9152);
or U9238 (N_9238,N_9030,N_9164);
xor U9239 (N_9239,N_9117,N_9084);
nand U9240 (N_9240,N_9106,N_9099);
xnor U9241 (N_9241,N_9194,N_9043);
nand U9242 (N_9242,N_9141,N_9142);
or U9243 (N_9243,N_9116,N_9157);
xor U9244 (N_9244,N_9094,N_9097);
and U9245 (N_9245,N_9087,N_9162);
nand U9246 (N_9246,N_9023,N_9052);
or U9247 (N_9247,N_9128,N_9156);
nand U9248 (N_9248,N_9086,N_9193);
or U9249 (N_9249,N_9137,N_9079);
nand U9250 (N_9250,N_9080,N_9004);
nand U9251 (N_9251,N_9191,N_9075);
nor U9252 (N_9252,N_9124,N_9048);
and U9253 (N_9253,N_9066,N_9067);
nand U9254 (N_9254,N_9132,N_9054);
and U9255 (N_9255,N_9105,N_9139);
or U9256 (N_9256,N_9056,N_9120);
xnor U9257 (N_9257,N_9122,N_9085);
or U9258 (N_9258,N_9021,N_9104);
or U9259 (N_9259,N_9140,N_9098);
nor U9260 (N_9260,N_9088,N_9071);
nor U9261 (N_9261,N_9170,N_9009);
nor U9262 (N_9262,N_9183,N_9119);
nand U9263 (N_9263,N_9057,N_9109);
nand U9264 (N_9264,N_9045,N_9040);
and U9265 (N_9265,N_9022,N_9026);
or U9266 (N_9266,N_9008,N_9154);
xor U9267 (N_9267,N_9159,N_9103);
and U9268 (N_9268,N_9051,N_9138);
or U9269 (N_9269,N_9187,N_9108);
nor U9270 (N_9270,N_9069,N_9158);
nor U9271 (N_9271,N_9165,N_9118);
nor U9272 (N_9272,N_9050,N_9077);
nor U9273 (N_9273,N_9136,N_9028);
xnor U9274 (N_9274,N_9027,N_9032);
and U9275 (N_9275,N_9111,N_9029);
or U9276 (N_9276,N_9145,N_9003);
nand U9277 (N_9277,N_9039,N_9064);
or U9278 (N_9278,N_9112,N_9147);
or U9279 (N_9279,N_9010,N_9044);
nand U9280 (N_9280,N_9174,N_9144);
or U9281 (N_9281,N_9082,N_9101);
nand U9282 (N_9282,N_9011,N_9175);
nor U9283 (N_9283,N_9172,N_9125);
nor U9284 (N_9284,N_9095,N_9134);
or U9285 (N_9285,N_9058,N_9062);
xnor U9286 (N_9286,N_9014,N_9184);
or U9287 (N_9287,N_9115,N_9055);
or U9288 (N_9288,N_9068,N_9110);
or U9289 (N_9289,N_9131,N_9015);
or U9290 (N_9290,N_9196,N_9149);
and U9291 (N_9291,N_9133,N_9114);
or U9292 (N_9292,N_9161,N_9143);
and U9293 (N_9293,N_9049,N_9034);
nor U9294 (N_9294,N_9059,N_9107);
nor U9295 (N_9295,N_9025,N_9180);
nand U9296 (N_9296,N_9168,N_9199);
nand U9297 (N_9297,N_9063,N_9081);
or U9298 (N_9298,N_9024,N_9019);
or U9299 (N_9299,N_9037,N_9090);
and U9300 (N_9300,N_9078,N_9000);
nand U9301 (N_9301,N_9071,N_9113);
or U9302 (N_9302,N_9112,N_9071);
nor U9303 (N_9303,N_9112,N_9068);
nor U9304 (N_9304,N_9067,N_9117);
or U9305 (N_9305,N_9024,N_9114);
nor U9306 (N_9306,N_9021,N_9198);
nor U9307 (N_9307,N_9028,N_9193);
or U9308 (N_9308,N_9054,N_9197);
and U9309 (N_9309,N_9100,N_9014);
nor U9310 (N_9310,N_9018,N_9019);
nand U9311 (N_9311,N_9154,N_9051);
xor U9312 (N_9312,N_9090,N_9113);
or U9313 (N_9313,N_9123,N_9122);
nand U9314 (N_9314,N_9088,N_9181);
nor U9315 (N_9315,N_9035,N_9112);
xnor U9316 (N_9316,N_9038,N_9147);
and U9317 (N_9317,N_9193,N_9037);
or U9318 (N_9318,N_9174,N_9127);
and U9319 (N_9319,N_9183,N_9022);
nand U9320 (N_9320,N_9136,N_9041);
nor U9321 (N_9321,N_9107,N_9106);
nor U9322 (N_9322,N_9158,N_9105);
xor U9323 (N_9323,N_9017,N_9139);
xnor U9324 (N_9324,N_9178,N_9044);
or U9325 (N_9325,N_9070,N_9034);
xor U9326 (N_9326,N_9116,N_9049);
nor U9327 (N_9327,N_9110,N_9115);
nor U9328 (N_9328,N_9183,N_9122);
and U9329 (N_9329,N_9065,N_9016);
and U9330 (N_9330,N_9101,N_9076);
nand U9331 (N_9331,N_9013,N_9056);
xor U9332 (N_9332,N_9122,N_9057);
nand U9333 (N_9333,N_9115,N_9088);
nand U9334 (N_9334,N_9127,N_9193);
nand U9335 (N_9335,N_9049,N_9090);
nand U9336 (N_9336,N_9133,N_9029);
nor U9337 (N_9337,N_9121,N_9077);
nor U9338 (N_9338,N_9175,N_9116);
and U9339 (N_9339,N_9100,N_9166);
and U9340 (N_9340,N_9034,N_9075);
nor U9341 (N_9341,N_9067,N_9100);
nand U9342 (N_9342,N_9191,N_9044);
xnor U9343 (N_9343,N_9007,N_9115);
nor U9344 (N_9344,N_9038,N_9041);
or U9345 (N_9345,N_9105,N_9075);
nand U9346 (N_9346,N_9013,N_9119);
xnor U9347 (N_9347,N_9190,N_9087);
or U9348 (N_9348,N_9031,N_9136);
nand U9349 (N_9349,N_9000,N_9170);
nand U9350 (N_9350,N_9103,N_9006);
nand U9351 (N_9351,N_9149,N_9184);
or U9352 (N_9352,N_9056,N_9119);
nor U9353 (N_9353,N_9077,N_9115);
xnor U9354 (N_9354,N_9020,N_9023);
nor U9355 (N_9355,N_9068,N_9018);
nor U9356 (N_9356,N_9083,N_9167);
and U9357 (N_9357,N_9197,N_9142);
xnor U9358 (N_9358,N_9187,N_9015);
or U9359 (N_9359,N_9056,N_9045);
nand U9360 (N_9360,N_9120,N_9071);
or U9361 (N_9361,N_9102,N_9010);
xnor U9362 (N_9362,N_9030,N_9031);
nand U9363 (N_9363,N_9155,N_9113);
xor U9364 (N_9364,N_9077,N_9079);
and U9365 (N_9365,N_9073,N_9059);
or U9366 (N_9366,N_9164,N_9065);
and U9367 (N_9367,N_9081,N_9001);
nand U9368 (N_9368,N_9101,N_9148);
xnor U9369 (N_9369,N_9186,N_9189);
xnor U9370 (N_9370,N_9016,N_9017);
or U9371 (N_9371,N_9114,N_9145);
or U9372 (N_9372,N_9096,N_9070);
nand U9373 (N_9373,N_9155,N_9118);
nor U9374 (N_9374,N_9039,N_9143);
nand U9375 (N_9375,N_9072,N_9196);
nand U9376 (N_9376,N_9147,N_9014);
nor U9377 (N_9377,N_9046,N_9012);
nand U9378 (N_9378,N_9090,N_9075);
nand U9379 (N_9379,N_9078,N_9072);
xor U9380 (N_9380,N_9135,N_9112);
and U9381 (N_9381,N_9089,N_9108);
xor U9382 (N_9382,N_9110,N_9020);
or U9383 (N_9383,N_9161,N_9090);
nor U9384 (N_9384,N_9090,N_9067);
or U9385 (N_9385,N_9044,N_9165);
nand U9386 (N_9386,N_9003,N_9109);
or U9387 (N_9387,N_9174,N_9128);
nor U9388 (N_9388,N_9115,N_9045);
nor U9389 (N_9389,N_9123,N_9156);
nand U9390 (N_9390,N_9096,N_9044);
nor U9391 (N_9391,N_9027,N_9171);
or U9392 (N_9392,N_9012,N_9076);
nor U9393 (N_9393,N_9036,N_9194);
or U9394 (N_9394,N_9096,N_9036);
nor U9395 (N_9395,N_9136,N_9096);
or U9396 (N_9396,N_9146,N_9094);
nand U9397 (N_9397,N_9115,N_9036);
xor U9398 (N_9398,N_9046,N_9038);
and U9399 (N_9399,N_9126,N_9195);
nand U9400 (N_9400,N_9242,N_9209);
or U9401 (N_9401,N_9219,N_9390);
or U9402 (N_9402,N_9270,N_9366);
nand U9403 (N_9403,N_9393,N_9202);
nor U9404 (N_9404,N_9326,N_9200);
or U9405 (N_9405,N_9260,N_9205);
nand U9406 (N_9406,N_9216,N_9322);
xnor U9407 (N_9407,N_9340,N_9259);
xor U9408 (N_9408,N_9271,N_9212);
and U9409 (N_9409,N_9309,N_9374);
nor U9410 (N_9410,N_9308,N_9223);
xnor U9411 (N_9411,N_9354,N_9389);
xnor U9412 (N_9412,N_9349,N_9249);
nand U9413 (N_9413,N_9336,N_9352);
nand U9414 (N_9414,N_9284,N_9338);
or U9415 (N_9415,N_9207,N_9386);
and U9416 (N_9416,N_9300,N_9225);
and U9417 (N_9417,N_9224,N_9321);
nor U9418 (N_9418,N_9359,N_9360);
and U9419 (N_9419,N_9283,N_9245);
or U9420 (N_9420,N_9337,N_9262);
and U9421 (N_9421,N_9278,N_9233);
nand U9422 (N_9422,N_9380,N_9320);
or U9423 (N_9423,N_9214,N_9281);
xnor U9424 (N_9424,N_9327,N_9215);
or U9425 (N_9425,N_9381,N_9232);
nand U9426 (N_9426,N_9286,N_9294);
or U9427 (N_9427,N_9398,N_9290);
xor U9428 (N_9428,N_9237,N_9251);
or U9429 (N_9429,N_9310,N_9288);
or U9430 (N_9430,N_9276,N_9228);
xor U9431 (N_9431,N_9285,N_9333);
nor U9432 (N_9432,N_9341,N_9235);
nand U9433 (N_9433,N_9234,N_9229);
xor U9434 (N_9434,N_9355,N_9350);
nor U9435 (N_9435,N_9268,N_9396);
nand U9436 (N_9436,N_9206,N_9247);
nor U9437 (N_9437,N_9365,N_9246);
nand U9438 (N_9438,N_9346,N_9343);
xor U9439 (N_9439,N_9287,N_9267);
and U9440 (N_9440,N_9264,N_9213);
nor U9441 (N_9441,N_9369,N_9339);
nand U9442 (N_9442,N_9208,N_9221);
nor U9443 (N_9443,N_9377,N_9266);
xnor U9444 (N_9444,N_9201,N_9238);
or U9445 (N_9445,N_9303,N_9344);
and U9446 (N_9446,N_9204,N_9399);
nor U9447 (N_9447,N_9311,N_9368);
nand U9448 (N_9448,N_9272,N_9296);
nand U9449 (N_9449,N_9301,N_9241);
and U9450 (N_9450,N_9392,N_9356);
or U9451 (N_9451,N_9370,N_9265);
xnor U9452 (N_9452,N_9319,N_9330);
and U9453 (N_9453,N_9334,N_9351);
or U9454 (N_9454,N_9302,N_9275);
nor U9455 (N_9455,N_9227,N_9314);
nand U9456 (N_9456,N_9277,N_9255);
nand U9457 (N_9457,N_9306,N_9280);
nand U9458 (N_9458,N_9388,N_9361);
nor U9459 (N_9459,N_9331,N_9293);
nor U9460 (N_9460,N_9307,N_9243);
nand U9461 (N_9461,N_9317,N_9394);
xnor U9462 (N_9462,N_9289,N_9328);
and U9463 (N_9463,N_9376,N_9323);
or U9464 (N_9464,N_9282,N_9304);
or U9465 (N_9465,N_9305,N_9312);
and U9466 (N_9466,N_9387,N_9373);
nor U9467 (N_9467,N_9353,N_9298);
and U9468 (N_9468,N_9342,N_9203);
or U9469 (N_9469,N_9291,N_9378);
or U9470 (N_9470,N_9332,N_9250);
and U9471 (N_9471,N_9274,N_9222);
nor U9472 (N_9472,N_9318,N_9297);
nor U9473 (N_9473,N_9347,N_9217);
xor U9474 (N_9474,N_9364,N_9231);
nor U9475 (N_9475,N_9218,N_9220);
or U9476 (N_9476,N_9295,N_9375);
nor U9477 (N_9477,N_9329,N_9382);
nand U9478 (N_9478,N_9335,N_9357);
and U9479 (N_9479,N_9367,N_9345);
nand U9480 (N_9480,N_9324,N_9256);
and U9481 (N_9481,N_9397,N_9379);
nor U9482 (N_9482,N_9313,N_9372);
xor U9483 (N_9483,N_9348,N_9211);
or U9484 (N_9484,N_9239,N_9385);
and U9485 (N_9485,N_9315,N_9240);
nor U9486 (N_9486,N_9244,N_9362);
xnor U9487 (N_9487,N_9292,N_9226);
nand U9488 (N_9488,N_9358,N_9363);
nand U9489 (N_9489,N_9230,N_9279);
or U9490 (N_9490,N_9261,N_9273);
nand U9491 (N_9491,N_9253,N_9371);
and U9492 (N_9492,N_9299,N_9236);
nand U9493 (N_9493,N_9395,N_9263);
and U9494 (N_9494,N_9316,N_9254);
and U9495 (N_9495,N_9384,N_9257);
xnor U9496 (N_9496,N_9391,N_9258);
and U9497 (N_9497,N_9210,N_9252);
nand U9498 (N_9498,N_9383,N_9325);
and U9499 (N_9499,N_9269,N_9248);
or U9500 (N_9500,N_9352,N_9263);
nand U9501 (N_9501,N_9306,N_9225);
nand U9502 (N_9502,N_9220,N_9358);
or U9503 (N_9503,N_9344,N_9227);
and U9504 (N_9504,N_9334,N_9335);
xor U9505 (N_9505,N_9305,N_9347);
nor U9506 (N_9506,N_9200,N_9330);
nor U9507 (N_9507,N_9255,N_9244);
nor U9508 (N_9508,N_9265,N_9297);
nor U9509 (N_9509,N_9393,N_9275);
nor U9510 (N_9510,N_9239,N_9386);
xor U9511 (N_9511,N_9206,N_9216);
and U9512 (N_9512,N_9264,N_9238);
nor U9513 (N_9513,N_9331,N_9357);
xnor U9514 (N_9514,N_9216,N_9315);
and U9515 (N_9515,N_9373,N_9362);
nand U9516 (N_9516,N_9255,N_9390);
or U9517 (N_9517,N_9363,N_9392);
xor U9518 (N_9518,N_9327,N_9209);
xor U9519 (N_9519,N_9322,N_9283);
nor U9520 (N_9520,N_9207,N_9228);
and U9521 (N_9521,N_9368,N_9338);
xnor U9522 (N_9522,N_9358,N_9373);
nand U9523 (N_9523,N_9355,N_9299);
or U9524 (N_9524,N_9298,N_9309);
nand U9525 (N_9525,N_9318,N_9273);
xor U9526 (N_9526,N_9264,N_9233);
xnor U9527 (N_9527,N_9215,N_9202);
xnor U9528 (N_9528,N_9283,N_9279);
or U9529 (N_9529,N_9312,N_9396);
nor U9530 (N_9530,N_9275,N_9280);
or U9531 (N_9531,N_9267,N_9245);
xor U9532 (N_9532,N_9345,N_9281);
xnor U9533 (N_9533,N_9218,N_9246);
nand U9534 (N_9534,N_9360,N_9301);
xor U9535 (N_9535,N_9346,N_9275);
nand U9536 (N_9536,N_9234,N_9220);
nor U9537 (N_9537,N_9312,N_9268);
and U9538 (N_9538,N_9389,N_9209);
or U9539 (N_9539,N_9399,N_9252);
or U9540 (N_9540,N_9398,N_9326);
nor U9541 (N_9541,N_9382,N_9280);
xor U9542 (N_9542,N_9358,N_9313);
nand U9543 (N_9543,N_9301,N_9204);
or U9544 (N_9544,N_9315,N_9227);
nand U9545 (N_9545,N_9360,N_9328);
xor U9546 (N_9546,N_9337,N_9273);
xnor U9547 (N_9547,N_9341,N_9238);
nand U9548 (N_9548,N_9369,N_9210);
nor U9549 (N_9549,N_9298,N_9294);
or U9550 (N_9550,N_9360,N_9259);
nand U9551 (N_9551,N_9266,N_9255);
xnor U9552 (N_9552,N_9219,N_9253);
or U9553 (N_9553,N_9297,N_9203);
or U9554 (N_9554,N_9313,N_9297);
and U9555 (N_9555,N_9322,N_9244);
nor U9556 (N_9556,N_9371,N_9342);
xnor U9557 (N_9557,N_9312,N_9353);
nor U9558 (N_9558,N_9257,N_9352);
xnor U9559 (N_9559,N_9320,N_9378);
and U9560 (N_9560,N_9272,N_9321);
or U9561 (N_9561,N_9358,N_9384);
and U9562 (N_9562,N_9272,N_9292);
nand U9563 (N_9563,N_9235,N_9223);
or U9564 (N_9564,N_9361,N_9269);
xnor U9565 (N_9565,N_9336,N_9290);
or U9566 (N_9566,N_9276,N_9270);
or U9567 (N_9567,N_9259,N_9394);
xnor U9568 (N_9568,N_9315,N_9239);
nor U9569 (N_9569,N_9289,N_9225);
or U9570 (N_9570,N_9265,N_9255);
nand U9571 (N_9571,N_9264,N_9361);
nor U9572 (N_9572,N_9302,N_9319);
and U9573 (N_9573,N_9391,N_9221);
nand U9574 (N_9574,N_9339,N_9344);
and U9575 (N_9575,N_9303,N_9233);
or U9576 (N_9576,N_9224,N_9218);
nor U9577 (N_9577,N_9389,N_9246);
nand U9578 (N_9578,N_9355,N_9351);
nand U9579 (N_9579,N_9305,N_9220);
xor U9580 (N_9580,N_9253,N_9246);
and U9581 (N_9581,N_9345,N_9328);
xor U9582 (N_9582,N_9306,N_9345);
nand U9583 (N_9583,N_9241,N_9367);
nor U9584 (N_9584,N_9359,N_9267);
or U9585 (N_9585,N_9277,N_9315);
nand U9586 (N_9586,N_9331,N_9298);
and U9587 (N_9587,N_9251,N_9214);
or U9588 (N_9588,N_9285,N_9298);
or U9589 (N_9589,N_9389,N_9285);
xnor U9590 (N_9590,N_9275,N_9266);
nand U9591 (N_9591,N_9334,N_9376);
or U9592 (N_9592,N_9201,N_9287);
nand U9593 (N_9593,N_9382,N_9222);
or U9594 (N_9594,N_9244,N_9321);
and U9595 (N_9595,N_9328,N_9317);
nor U9596 (N_9596,N_9343,N_9314);
nand U9597 (N_9597,N_9288,N_9298);
xnor U9598 (N_9598,N_9361,N_9329);
nand U9599 (N_9599,N_9265,N_9220);
xor U9600 (N_9600,N_9412,N_9526);
nor U9601 (N_9601,N_9535,N_9599);
nand U9602 (N_9602,N_9588,N_9544);
or U9603 (N_9603,N_9420,N_9576);
nand U9604 (N_9604,N_9435,N_9414);
nand U9605 (N_9605,N_9453,N_9490);
and U9606 (N_9606,N_9468,N_9426);
nand U9607 (N_9607,N_9474,N_9569);
xnor U9608 (N_9608,N_9579,N_9571);
nand U9609 (N_9609,N_9597,N_9587);
or U9610 (N_9610,N_9523,N_9424);
nand U9611 (N_9611,N_9473,N_9447);
nand U9612 (N_9612,N_9520,N_9545);
nand U9613 (N_9613,N_9409,N_9596);
xnor U9614 (N_9614,N_9512,N_9431);
nor U9615 (N_9615,N_9527,N_9491);
or U9616 (N_9616,N_9427,N_9481);
nor U9617 (N_9617,N_9561,N_9593);
or U9618 (N_9618,N_9476,N_9539);
and U9619 (N_9619,N_9483,N_9438);
nand U9620 (N_9620,N_9470,N_9408);
xnor U9621 (N_9621,N_9556,N_9584);
nor U9622 (N_9622,N_9421,N_9585);
or U9623 (N_9623,N_9560,N_9485);
xor U9624 (N_9624,N_9482,N_9546);
nand U9625 (N_9625,N_9404,N_9402);
xnor U9626 (N_9626,N_9501,N_9416);
xnor U9627 (N_9627,N_9439,N_9507);
or U9628 (N_9628,N_9595,N_9513);
xnor U9629 (N_9629,N_9542,N_9417);
nand U9630 (N_9630,N_9541,N_9466);
nor U9631 (N_9631,N_9573,N_9515);
and U9632 (N_9632,N_9534,N_9423);
or U9633 (N_9633,N_9455,N_9403);
nand U9634 (N_9634,N_9503,N_9458);
nor U9635 (N_9635,N_9457,N_9500);
and U9636 (N_9636,N_9567,N_9449);
xnor U9637 (N_9637,N_9415,N_9442);
nor U9638 (N_9638,N_9492,N_9405);
nor U9639 (N_9639,N_9574,N_9422);
nor U9640 (N_9640,N_9570,N_9496);
nand U9641 (N_9641,N_9552,N_9589);
xnor U9642 (N_9642,N_9484,N_9428);
xnor U9643 (N_9643,N_9499,N_9452);
xor U9644 (N_9644,N_9598,N_9462);
nor U9645 (N_9645,N_9537,N_9592);
xor U9646 (N_9646,N_9559,N_9448);
nand U9647 (N_9647,N_9531,N_9495);
or U9648 (N_9648,N_9510,N_9555);
nor U9649 (N_9649,N_9434,N_9437);
xnor U9650 (N_9650,N_9430,N_9443);
xnor U9651 (N_9651,N_9451,N_9400);
xor U9652 (N_9652,N_9410,N_9553);
and U9653 (N_9653,N_9538,N_9425);
and U9654 (N_9654,N_9548,N_9557);
and U9655 (N_9655,N_9480,N_9488);
nor U9656 (N_9656,N_9497,N_9464);
nand U9657 (N_9657,N_9407,N_9508);
or U9658 (N_9658,N_9540,N_9519);
nor U9659 (N_9659,N_9440,N_9493);
and U9660 (N_9660,N_9433,N_9578);
and U9661 (N_9661,N_9516,N_9459);
and U9662 (N_9662,N_9518,N_9562);
and U9663 (N_9663,N_9532,N_9401);
nand U9664 (N_9664,N_9465,N_9486);
xor U9665 (N_9665,N_9554,N_9517);
and U9666 (N_9666,N_9471,N_9536);
nor U9667 (N_9667,N_9446,N_9411);
and U9668 (N_9668,N_9472,N_9575);
nand U9669 (N_9669,N_9505,N_9547);
and U9670 (N_9670,N_9583,N_9502);
nor U9671 (N_9671,N_9564,N_9550);
nor U9672 (N_9672,N_9504,N_9525);
or U9673 (N_9673,N_9591,N_9477);
nand U9674 (N_9674,N_9582,N_9524);
and U9675 (N_9675,N_9568,N_9450);
xnor U9676 (N_9676,N_9586,N_9577);
xor U9677 (N_9677,N_9413,N_9436);
or U9678 (N_9678,N_9514,N_9498);
and U9679 (N_9679,N_9419,N_9521);
nand U9680 (N_9680,N_9489,N_9590);
and U9681 (N_9681,N_9487,N_9549);
xnor U9682 (N_9682,N_9511,N_9581);
nor U9683 (N_9683,N_9580,N_9429);
nor U9684 (N_9684,N_9529,N_9543);
or U9685 (N_9685,N_9522,N_9551);
or U9686 (N_9686,N_9444,N_9563);
or U9687 (N_9687,N_9456,N_9445);
xor U9688 (N_9688,N_9406,N_9461);
xor U9689 (N_9689,N_9475,N_9566);
nor U9690 (N_9690,N_9533,N_9478);
and U9691 (N_9691,N_9467,N_9469);
or U9692 (N_9692,N_9528,N_9530);
or U9693 (N_9693,N_9479,N_9454);
xnor U9694 (N_9694,N_9494,N_9565);
nand U9695 (N_9695,N_9432,N_9506);
nor U9696 (N_9696,N_9441,N_9509);
xnor U9697 (N_9697,N_9463,N_9558);
xnor U9698 (N_9698,N_9572,N_9418);
or U9699 (N_9699,N_9460,N_9594);
xor U9700 (N_9700,N_9556,N_9548);
nor U9701 (N_9701,N_9500,N_9502);
nand U9702 (N_9702,N_9478,N_9592);
nand U9703 (N_9703,N_9453,N_9417);
xor U9704 (N_9704,N_9475,N_9428);
xor U9705 (N_9705,N_9522,N_9534);
nand U9706 (N_9706,N_9554,N_9591);
and U9707 (N_9707,N_9434,N_9527);
nor U9708 (N_9708,N_9594,N_9425);
or U9709 (N_9709,N_9500,N_9568);
or U9710 (N_9710,N_9488,N_9468);
and U9711 (N_9711,N_9416,N_9453);
xor U9712 (N_9712,N_9543,N_9598);
and U9713 (N_9713,N_9535,N_9554);
nand U9714 (N_9714,N_9539,N_9598);
and U9715 (N_9715,N_9524,N_9478);
xnor U9716 (N_9716,N_9442,N_9479);
or U9717 (N_9717,N_9441,N_9472);
xor U9718 (N_9718,N_9503,N_9491);
xnor U9719 (N_9719,N_9553,N_9517);
nand U9720 (N_9720,N_9588,N_9476);
nor U9721 (N_9721,N_9533,N_9447);
nor U9722 (N_9722,N_9537,N_9413);
nand U9723 (N_9723,N_9461,N_9500);
nor U9724 (N_9724,N_9485,N_9525);
or U9725 (N_9725,N_9598,N_9578);
nand U9726 (N_9726,N_9514,N_9599);
xnor U9727 (N_9727,N_9575,N_9481);
nor U9728 (N_9728,N_9468,N_9497);
nand U9729 (N_9729,N_9540,N_9417);
nor U9730 (N_9730,N_9515,N_9424);
nor U9731 (N_9731,N_9484,N_9521);
nor U9732 (N_9732,N_9480,N_9493);
and U9733 (N_9733,N_9521,N_9464);
nand U9734 (N_9734,N_9580,N_9576);
nor U9735 (N_9735,N_9490,N_9491);
and U9736 (N_9736,N_9563,N_9474);
or U9737 (N_9737,N_9418,N_9510);
and U9738 (N_9738,N_9483,N_9507);
or U9739 (N_9739,N_9511,N_9432);
and U9740 (N_9740,N_9545,N_9547);
xor U9741 (N_9741,N_9476,N_9423);
or U9742 (N_9742,N_9591,N_9537);
nand U9743 (N_9743,N_9456,N_9506);
or U9744 (N_9744,N_9512,N_9549);
nand U9745 (N_9745,N_9424,N_9501);
nand U9746 (N_9746,N_9526,N_9421);
or U9747 (N_9747,N_9406,N_9574);
xnor U9748 (N_9748,N_9520,N_9473);
nor U9749 (N_9749,N_9576,N_9542);
xor U9750 (N_9750,N_9544,N_9552);
or U9751 (N_9751,N_9571,N_9448);
nor U9752 (N_9752,N_9548,N_9497);
nor U9753 (N_9753,N_9503,N_9481);
and U9754 (N_9754,N_9471,N_9571);
nand U9755 (N_9755,N_9400,N_9489);
and U9756 (N_9756,N_9448,N_9427);
or U9757 (N_9757,N_9458,N_9419);
or U9758 (N_9758,N_9565,N_9559);
xnor U9759 (N_9759,N_9471,N_9469);
xor U9760 (N_9760,N_9403,N_9413);
nor U9761 (N_9761,N_9587,N_9433);
nand U9762 (N_9762,N_9466,N_9527);
xnor U9763 (N_9763,N_9506,N_9524);
xnor U9764 (N_9764,N_9569,N_9572);
xor U9765 (N_9765,N_9425,N_9529);
xor U9766 (N_9766,N_9510,N_9527);
nand U9767 (N_9767,N_9417,N_9483);
or U9768 (N_9768,N_9457,N_9546);
and U9769 (N_9769,N_9582,N_9496);
or U9770 (N_9770,N_9581,N_9584);
or U9771 (N_9771,N_9450,N_9565);
or U9772 (N_9772,N_9509,N_9592);
xnor U9773 (N_9773,N_9490,N_9541);
and U9774 (N_9774,N_9403,N_9562);
nand U9775 (N_9775,N_9471,N_9522);
or U9776 (N_9776,N_9568,N_9472);
or U9777 (N_9777,N_9537,N_9573);
nor U9778 (N_9778,N_9576,N_9535);
nand U9779 (N_9779,N_9407,N_9559);
nor U9780 (N_9780,N_9410,N_9594);
nor U9781 (N_9781,N_9447,N_9589);
or U9782 (N_9782,N_9580,N_9402);
nor U9783 (N_9783,N_9542,N_9589);
nor U9784 (N_9784,N_9467,N_9433);
nand U9785 (N_9785,N_9488,N_9582);
xnor U9786 (N_9786,N_9506,N_9556);
xor U9787 (N_9787,N_9554,N_9573);
and U9788 (N_9788,N_9511,N_9518);
nor U9789 (N_9789,N_9403,N_9420);
nor U9790 (N_9790,N_9405,N_9484);
nand U9791 (N_9791,N_9486,N_9435);
nor U9792 (N_9792,N_9483,N_9557);
or U9793 (N_9793,N_9597,N_9565);
nor U9794 (N_9794,N_9520,N_9535);
nor U9795 (N_9795,N_9420,N_9518);
or U9796 (N_9796,N_9423,N_9556);
nand U9797 (N_9797,N_9477,N_9428);
nor U9798 (N_9798,N_9403,N_9508);
or U9799 (N_9799,N_9433,N_9450);
or U9800 (N_9800,N_9627,N_9795);
and U9801 (N_9801,N_9693,N_9680);
and U9802 (N_9802,N_9729,N_9790);
and U9803 (N_9803,N_9759,N_9740);
or U9804 (N_9804,N_9768,N_9771);
or U9805 (N_9805,N_9727,N_9610);
xnor U9806 (N_9806,N_9754,N_9648);
nand U9807 (N_9807,N_9682,N_9644);
nor U9808 (N_9808,N_9684,N_9751);
xor U9809 (N_9809,N_9666,N_9755);
nand U9810 (N_9810,N_9690,N_9641);
and U9811 (N_9811,N_9647,N_9619);
nor U9812 (N_9812,N_9658,N_9654);
and U9813 (N_9813,N_9659,N_9633);
nand U9814 (N_9814,N_9700,N_9718);
xor U9815 (N_9815,N_9672,N_9750);
or U9816 (N_9816,N_9667,N_9653);
nand U9817 (N_9817,N_9786,N_9652);
nor U9818 (N_9818,N_9605,N_9630);
nand U9819 (N_9819,N_9760,N_9770);
and U9820 (N_9820,N_9702,N_9797);
xor U9821 (N_9821,N_9618,N_9695);
or U9822 (N_9822,N_9634,N_9613);
and U9823 (N_9823,N_9642,N_9776);
nor U9824 (N_9824,N_9712,N_9792);
or U9825 (N_9825,N_9688,N_9791);
nand U9826 (N_9826,N_9753,N_9701);
nor U9827 (N_9827,N_9663,N_9748);
nor U9828 (N_9828,N_9721,N_9779);
nand U9829 (N_9829,N_9628,N_9625);
nor U9830 (N_9830,N_9780,N_9762);
or U9831 (N_9831,N_9621,N_9720);
or U9832 (N_9832,N_9631,N_9725);
and U9833 (N_9833,N_9743,N_9734);
and U9834 (N_9834,N_9703,N_9774);
xor U9835 (N_9835,N_9739,N_9664);
nand U9836 (N_9836,N_9685,N_9752);
and U9837 (N_9837,N_9707,N_9675);
and U9838 (N_9838,N_9668,N_9655);
nor U9839 (N_9839,N_9607,N_9719);
and U9840 (N_9840,N_9717,N_9794);
xor U9841 (N_9841,N_9635,N_9710);
or U9842 (N_9842,N_9705,N_9784);
and U9843 (N_9843,N_9764,N_9636);
and U9844 (N_9844,N_9724,N_9761);
or U9845 (N_9845,N_9765,N_9670);
xnor U9846 (N_9846,N_9726,N_9772);
and U9847 (N_9847,N_9778,N_9715);
nor U9848 (N_9848,N_9669,N_9747);
nand U9849 (N_9849,N_9650,N_9601);
xor U9850 (N_9850,N_9713,N_9632);
xor U9851 (N_9851,N_9783,N_9741);
nand U9852 (N_9852,N_9602,N_9620);
xnor U9853 (N_9853,N_9671,N_9657);
and U9854 (N_9854,N_9709,N_9678);
and U9855 (N_9855,N_9656,N_9617);
or U9856 (N_9856,N_9733,N_9732);
or U9857 (N_9857,N_9694,N_9766);
or U9858 (N_9858,N_9683,N_9612);
nor U9859 (N_9859,N_9745,N_9638);
xnor U9860 (N_9860,N_9735,N_9603);
and U9861 (N_9861,N_9737,N_9640);
xnor U9862 (N_9862,N_9742,N_9689);
xnor U9863 (N_9863,N_9781,N_9676);
xor U9864 (N_9864,N_9738,N_9660);
or U9865 (N_9865,N_9787,N_9758);
xor U9866 (N_9866,N_9637,N_9622);
xnor U9867 (N_9867,N_9763,N_9645);
or U9868 (N_9868,N_9639,N_9757);
or U9869 (N_9869,N_9796,N_9608);
and U9870 (N_9870,N_9600,N_9651);
xor U9871 (N_9871,N_9646,N_9699);
and U9872 (N_9872,N_9606,N_9691);
and U9873 (N_9873,N_9736,N_9611);
or U9874 (N_9874,N_9785,N_9687);
and U9875 (N_9875,N_9696,N_9775);
and U9876 (N_9876,N_9769,N_9626);
nor U9877 (N_9877,N_9662,N_9777);
nor U9878 (N_9878,N_9679,N_9698);
nor U9879 (N_9879,N_9623,N_9731);
nor U9880 (N_9880,N_9773,N_9756);
nand U9881 (N_9881,N_9728,N_9624);
nand U9882 (N_9882,N_9681,N_9604);
xor U9883 (N_9883,N_9704,N_9673);
nor U9884 (N_9884,N_9706,N_9714);
xor U9885 (N_9885,N_9686,N_9744);
or U9886 (N_9886,N_9798,N_9782);
and U9887 (N_9887,N_9616,N_9749);
or U9888 (N_9888,N_9789,N_9799);
xnor U9889 (N_9889,N_9674,N_9614);
and U9890 (N_9890,N_9629,N_9649);
nand U9891 (N_9891,N_9767,N_9723);
or U9892 (N_9892,N_9697,N_9722);
nand U9893 (N_9893,N_9643,N_9692);
nor U9894 (N_9894,N_9615,N_9793);
nor U9895 (N_9895,N_9711,N_9665);
nor U9896 (N_9896,N_9746,N_9677);
or U9897 (N_9897,N_9661,N_9708);
nand U9898 (N_9898,N_9730,N_9716);
nor U9899 (N_9899,N_9609,N_9788);
and U9900 (N_9900,N_9646,N_9602);
and U9901 (N_9901,N_9688,N_9654);
or U9902 (N_9902,N_9624,N_9691);
xor U9903 (N_9903,N_9708,N_9605);
xnor U9904 (N_9904,N_9670,N_9654);
nor U9905 (N_9905,N_9713,N_9760);
nand U9906 (N_9906,N_9721,N_9725);
xor U9907 (N_9907,N_9623,N_9685);
nand U9908 (N_9908,N_9607,N_9695);
xnor U9909 (N_9909,N_9763,N_9699);
nor U9910 (N_9910,N_9714,N_9645);
nor U9911 (N_9911,N_9607,N_9654);
xor U9912 (N_9912,N_9603,N_9646);
and U9913 (N_9913,N_9613,N_9644);
or U9914 (N_9914,N_9628,N_9685);
xor U9915 (N_9915,N_9692,N_9728);
and U9916 (N_9916,N_9613,N_9625);
or U9917 (N_9917,N_9717,N_9783);
nand U9918 (N_9918,N_9687,N_9742);
xor U9919 (N_9919,N_9655,N_9693);
nand U9920 (N_9920,N_9677,N_9747);
xnor U9921 (N_9921,N_9693,N_9670);
nor U9922 (N_9922,N_9699,N_9727);
xnor U9923 (N_9923,N_9695,N_9671);
nor U9924 (N_9924,N_9620,N_9692);
and U9925 (N_9925,N_9723,N_9649);
nand U9926 (N_9926,N_9653,N_9763);
or U9927 (N_9927,N_9683,N_9747);
nand U9928 (N_9928,N_9668,N_9658);
or U9929 (N_9929,N_9717,N_9762);
xnor U9930 (N_9930,N_9662,N_9778);
nor U9931 (N_9931,N_9744,N_9781);
and U9932 (N_9932,N_9654,N_9792);
nor U9933 (N_9933,N_9626,N_9759);
or U9934 (N_9934,N_9616,N_9773);
nand U9935 (N_9935,N_9723,N_9644);
or U9936 (N_9936,N_9719,N_9786);
and U9937 (N_9937,N_9780,N_9797);
nor U9938 (N_9938,N_9748,N_9644);
nand U9939 (N_9939,N_9787,N_9704);
nand U9940 (N_9940,N_9790,N_9631);
or U9941 (N_9941,N_9604,N_9633);
nor U9942 (N_9942,N_9642,N_9774);
nor U9943 (N_9943,N_9670,N_9759);
xnor U9944 (N_9944,N_9629,N_9782);
and U9945 (N_9945,N_9672,N_9754);
or U9946 (N_9946,N_9621,N_9733);
or U9947 (N_9947,N_9747,N_9742);
and U9948 (N_9948,N_9738,N_9773);
and U9949 (N_9949,N_9612,N_9777);
nor U9950 (N_9950,N_9796,N_9667);
or U9951 (N_9951,N_9735,N_9643);
or U9952 (N_9952,N_9694,N_9752);
nor U9953 (N_9953,N_9625,N_9731);
nor U9954 (N_9954,N_9612,N_9687);
and U9955 (N_9955,N_9674,N_9789);
nand U9956 (N_9956,N_9627,N_9767);
xnor U9957 (N_9957,N_9773,N_9609);
xnor U9958 (N_9958,N_9663,N_9639);
xor U9959 (N_9959,N_9603,N_9610);
and U9960 (N_9960,N_9686,N_9693);
xnor U9961 (N_9961,N_9699,N_9621);
and U9962 (N_9962,N_9756,N_9722);
xor U9963 (N_9963,N_9729,N_9673);
nor U9964 (N_9964,N_9776,N_9795);
and U9965 (N_9965,N_9754,N_9736);
and U9966 (N_9966,N_9675,N_9781);
nand U9967 (N_9967,N_9700,N_9795);
or U9968 (N_9968,N_9696,N_9714);
nand U9969 (N_9969,N_9604,N_9799);
nor U9970 (N_9970,N_9636,N_9792);
nand U9971 (N_9971,N_9761,N_9646);
or U9972 (N_9972,N_9697,N_9657);
nand U9973 (N_9973,N_9697,N_9665);
xnor U9974 (N_9974,N_9767,N_9605);
and U9975 (N_9975,N_9704,N_9654);
nor U9976 (N_9976,N_9749,N_9769);
xnor U9977 (N_9977,N_9650,N_9645);
nand U9978 (N_9978,N_9683,N_9769);
nand U9979 (N_9979,N_9712,N_9632);
xor U9980 (N_9980,N_9660,N_9636);
nand U9981 (N_9981,N_9777,N_9689);
xor U9982 (N_9982,N_9644,N_9740);
and U9983 (N_9983,N_9726,N_9695);
and U9984 (N_9984,N_9758,N_9686);
nand U9985 (N_9985,N_9675,N_9717);
nand U9986 (N_9986,N_9759,N_9646);
and U9987 (N_9987,N_9624,N_9773);
nor U9988 (N_9988,N_9686,N_9793);
xnor U9989 (N_9989,N_9740,N_9645);
and U9990 (N_9990,N_9769,N_9680);
or U9991 (N_9991,N_9685,N_9607);
nor U9992 (N_9992,N_9720,N_9682);
or U9993 (N_9993,N_9659,N_9770);
nand U9994 (N_9994,N_9658,N_9758);
or U9995 (N_9995,N_9796,N_9648);
nand U9996 (N_9996,N_9716,N_9645);
or U9997 (N_9997,N_9674,N_9773);
and U9998 (N_9998,N_9651,N_9627);
nand U9999 (N_9999,N_9650,N_9639);
nand U10000 (N_10000,N_9953,N_9834);
or U10001 (N_10001,N_9827,N_9946);
or U10002 (N_10002,N_9940,N_9842);
and U10003 (N_10003,N_9902,N_9811);
nor U10004 (N_10004,N_9813,N_9990);
xnor U10005 (N_10005,N_9839,N_9890);
and U10006 (N_10006,N_9830,N_9911);
xnor U10007 (N_10007,N_9966,N_9944);
or U10008 (N_10008,N_9992,N_9910);
nand U10009 (N_10009,N_9958,N_9879);
nor U10010 (N_10010,N_9818,N_9980);
xnor U10011 (N_10011,N_9820,N_9851);
and U10012 (N_10012,N_9939,N_9878);
nor U10013 (N_10013,N_9871,N_9885);
and U10014 (N_10014,N_9826,N_9899);
nor U10015 (N_10015,N_9805,N_9965);
and U10016 (N_10016,N_9912,N_9845);
nand U10017 (N_10017,N_9840,N_9947);
xnor U10018 (N_10018,N_9831,N_9859);
or U10019 (N_10019,N_9926,N_9846);
nand U10020 (N_10020,N_9988,N_9861);
and U10021 (N_10021,N_9867,N_9967);
nor U10022 (N_10022,N_9886,N_9882);
and U10023 (N_10023,N_9987,N_9907);
and U10024 (N_10024,N_9961,N_9956);
xor U10025 (N_10025,N_9924,N_9994);
nor U10026 (N_10026,N_9815,N_9962);
nand U10027 (N_10027,N_9986,N_9854);
xnor U10028 (N_10028,N_9989,N_9853);
nor U10029 (N_10029,N_9875,N_9841);
xor U10030 (N_10030,N_9898,N_9801);
or U10031 (N_10031,N_9909,N_9933);
xnor U10032 (N_10032,N_9937,N_9825);
xor U10033 (N_10033,N_9971,N_9935);
or U10034 (N_10034,N_9881,N_9900);
nand U10035 (N_10035,N_9888,N_9968);
xor U10036 (N_10036,N_9873,N_9970);
nand U10037 (N_10037,N_9903,N_9942);
and U10038 (N_10038,N_9856,N_9915);
nor U10039 (N_10039,N_9951,N_9809);
nand U10040 (N_10040,N_9857,N_9802);
and U10041 (N_10041,N_9869,N_9976);
nand U10042 (N_10042,N_9877,N_9804);
or U10043 (N_10043,N_9897,N_9983);
nor U10044 (N_10044,N_9978,N_9998);
xor U10045 (N_10045,N_9810,N_9843);
or U10046 (N_10046,N_9932,N_9922);
nand U10047 (N_10047,N_9829,N_9838);
xor U10048 (N_10048,N_9808,N_9923);
or U10049 (N_10049,N_9862,N_9930);
xor U10050 (N_10050,N_9889,N_9925);
and U10051 (N_10051,N_9814,N_9884);
nand U10052 (N_10052,N_9858,N_9863);
nand U10053 (N_10053,N_9936,N_9816);
xor U10054 (N_10054,N_9918,N_9905);
xor U10055 (N_10055,N_9849,N_9864);
nand U10056 (N_10056,N_9913,N_9904);
or U10057 (N_10057,N_9806,N_9945);
nand U10058 (N_10058,N_9824,N_9921);
and U10059 (N_10059,N_9927,N_9895);
and U10060 (N_10060,N_9835,N_9916);
and U10061 (N_10061,N_9959,N_9821);
and U10062 (N_10062,N_9828,N_9969);
or U10063 (N_10063,N_9952,N_9974);
nor U10064 (N_10064,N_9844,N_9876);
nand U10065 (N_10065,N_9896,N_9880);
or U10066 (N_10066,N_9991,N_9865);
xnor U10067 (N_10067,N_9914,N_9800);
xor U10068 (N_10068,N_9872,N_9931);
or U10069 (N_10069,N_9855,N_9850);
nor U10070 (N_10070,N_9929,N_9997);
and U10071 (N_10071,N_9948,N_9891);
nand U10072 (N_10072,N_9906,N_9860);
or U10073 (N_10073,N_9870,N_9938);
nor U10074 (N_10074,N_9848,N_9999);
nor U10075 (N_10075,N_9972,N_9837);
nor U10076 (N_10076,N_9981,N_9985);
and U10077 (N_10077,N_9893,N_9934);
nor U10078 (N_10078,N_9955,N_9812);
xor U10079 (N_10079,N_9819,N_9977);
xor U10080 (N_10080,N_9887,N_9917);
xor U10081 (N_10081,N_9847,N_9852);
nand U10082 (N_10082,N_9964,N_9822);
xnor U10083 (N_10083,N_9979,N_9949);
nor U10084 (N_10084,N_9996,N_9807);
or U10085 (N_10085,N_9883,N_9993);
and U10086 (N_10086,N_9894,N_9973);
xor U10087 (N_10087,N_9919,N_9803);
nor U10088 (N_10088,N_9874,N_9963);
or U10089 (N_10089,N_9908,N_9984);
nor U10090 (N_10090,N_9833,N_9868);
nand U10091 (N_10091,N_9817,N_9954);
or U10092 (N_10092,N_9957,N_9995);
nor U10093 (N_10093,N_9866,N_9836);
xor U10094 (N_10094,N_9960,N_9975);
and U10095 (N_10095,N_9943,N_9832);
xor U10096 (N_10096,N_9901,N_9892);
and U10097 (N_10097,N_9823,N_9950);
and U10098 (N_10098,N_9928,N_9982);
and U10099 (N_10099,N_9920,N_9941);
and U10100 (N_10100,N_9968,N_9971);
xnor U10101 (N_10101,N_9974,N_9886);
nand U10102 (N_10102,N_9899,N_9834);
nand U10103 (N_10103,N_9937,N_9843);
nand U10104 (N_10104,N_9930,N_9962);
or U10105 (N_10105,N_9959,N_9974);
nor U10106 (N_10106,N_9876,N_9867);
xnor U10107 (N_10107,N_9960,N_9936);
nand U10108 (N_10108,N_9857,N_9968);
xor U10109 (N_10109,N_9959,N_9826);
nand U10110 (N_10110,N_9926,N_9818);
xnor U10111 (N_10111,N_9852,N_9973);
xor U10112 (N_10112,N_9959,N_9886);
nor U10113 (N_10113,N_9954,N_9838);
xnor U10114 (N_10114,N_9976,N_9865);
and U10115 (N_10115,N_9930,N_9965);
or U10116 (N_10116,N_9806,N_9850);
or U10117 (N_10117,N_9972,N_9817);
nor U10118 (N_10118,N_9881,N_9805);
or U10119 (N_10119,N_9967,N_9913);
or U10120 (N_10120,N_9914,N_9997);
nand U10121 (N_10121,N_9871,N_9802);
nor U10122 (N_10122,N_9940,N_9897);
xor U10123 (N_10123,N_9890,N_9918);
or U10124 (N_10124,N_9913,N_9987);
nor U10125 (N_10125,N_9806,N_9936);
nand U10126 (N_10126,N_9953,N_9832);
or U10127 (N_10127,N_9814,N_9878);
or U10128 (N_10128,N_9964,N_9862);
nand U10129 (N_10129,N_9869,N_9827);
nand U10130 (N_10130,N_9948,N_9803);
xor U10131 (N_10131,N_9838,N_9885);
xnor U10132 (N_10132,N_9845,N_9891);
nor U10133 (N_10133,N_9806,N_9961);
nor U10134 (N_10134,N_9968,N_9924);
or U10135 (N_10135,N_9822,N_9932);
and U10136 (N_10136,N_9955,N_9915);
xor U10137 (N_10137,N_9837,N_9839);
xnor U10138 (N_10138,N_9915,N_9902);
nor U10139 (N_10139,N_9928,N_9863);
or U10140 (N_10140,N_9965,N_9990);
nand U10141 (N_10141,N_9961,N_9902);
xnor U10142 (N_10142,N_9944,N_9870);
nand U10143 (N_10143,N_9963,N_9853);
or U10144 (N_10144,N_9866,N_9968);
and U10145 (N_10145,N_9963,N_9886);
nand U10146 (N_10146,N_9836,N_9837);
xnor U10147 (N_10147,N_9947,N_9870);
and U10148 (N_10148,N_9971,N_9970);
nor U10149 (N_10149,N_9851,N_9859);
and U10150 (N_10150,N_9966,N_9940);
xnor U10151 (N_10151,N_9902,N_9868);
nor U10152 (N_10152,N_9836,N_9879);
and U10153 (N_10153,N_9810,N_9901);
nor U10154 (N_10154,N_9890,N_9844);
or U10155 (N_10155,N_9981,N_9906);
or U10156 (N_10156,N_9908,N_9850);
xor U10157 (N_10157,N_9976,N_9845);
nor U10158 (N_10158,N_9919,N_9900);
or U10159 (N_10159,N_9804,N_9846);
xnor U10160 (N_10160,N_9948,N_9932);
or U10161 (N_10161,N_9835,N_9905);
nand U10162 (N_10162,N_9999,N_9825);
or U10163 (N_10163,N_9827,N_9851);
xor U10164 (N_10164,N_9840,N_9862);
and U10165 (N_10165,N_9811,N_9948);
xor U10166 (N_10166,N_9875,N_9989);
nor U10167 (N_10167,N_9998,N_9932);
nand U10168 (N_10168,N_9868,N_9807);
xnor U10169 (N_10169,N_9925,N_9877);
nand U10170 (N_10170,N_9897,N_9939);
and U10171 (N_10171,N_9989,N_9920);
nand U10172 (N_10172,N_9965,N_9925);
or U10173 (N_10173,N_9901,N_9824);
or U10174 (N_10174,N_9852,N_9867);
and U10175 (N_10175,N_9832,N_9937);
or U10176 (N_10176,N_9976,N_9989);
nor U10177 (N_10177,N_9900,N_9878);
nand U10178 (N_10178,N_9998,N_9881);
and U10179 (N_10179,N_9929,N_9894);
nor U10180 (N_10180,N_9839,N_9947);
or U10181 (N_10181,N_9832,N_9958);
nand U10182 (N_10182,N_9943,N_9920);
nor U10183 (N_10183,N_9817,N_9876);
xor U10184 (N_10184,N_9824,N_9808);
nand U10185 (N_10185,N_9906,N_9874);
xor U10186 (N_10186,N_9933,N_9938);
xor U10187 (N_10187,N_9835,N_9946);
xnor U10188 (N_10188,N_9851,N_9912);
and U10189 (N_10189,N_9930,N_9953);
and U10190 (N_10190,N_9868,N_9806);
nor U10191 (N_10191,N_9929,N_9813);
xor U10192 (N_10192,N_9864,N_9858);
and U10193 (N_10193,N_9959,N_9957);
xnor U10194 (N_10194,N_9905,N_9927);
xnor U10195 (N_10195,N_9830,N_9836);
nand U10196 (N_10196,N_9975,N_9845);
and U10197 (N_10197,N_9829,N_9920);
nor U10198 (N_10198,N_9989,N_9848);
or U10199 (N_10199,N_9815,N_9877);
xnor U10200 (N_10200,N_10081,N_10157);
xor U10201 (N_10201,N_10188,N_10073);
xnor U10202 (N_10202,N_10022,N_10044);
nand U10203 (N_10203,N_10153,N_10050);
or U10204 (N_10204,N_10111,N_10100);
nor U10205 (N_10205,N_10065,N_10159);
xor U10206 (N_10206,N_10162,N_10094);
nor U10207 (N_10207,N_10057,N_10142);
nand U10208 (N_10208,N_10064,N_10008);
nand U10209 (N_10209,N_10087,N_10123);
and U10210 (N_10210,N_10071,N_10067);
and U10211 (N_10211,N_10000,N_10038);
and U10212 (N_10212,N_10131,N_10060);
and U10213 (N_10213,N_10175,N_10069);
nor U10214 (N_10214,N_10035,N_10105);
nand U10215 (N_10215,N_10079,N_10075);
nand U10216 (N_10216,N_10037,N_10156);
xor U10217 (N_10217,N_10195,N_10063);
or U10218 (N_10218,N_10090,N_10102);
nand U10219 (N_10219,N_10164,N_10154);
xnor U10220 (N_10220,N_10146,N_10034);
and U10221 (N_10221,N_10169,N_10119);
nor U10222 (N_10222,N_10137,N_10092);
nand U10223 (N_10223,N_10017,N_10026);
nor U10224 (N_10224,N_10056,N_10132);
or U10225 (N_10225,N_10055,N_10061);
and U10226 (N_10226,N_10014,N_10040);
nand U10227 (N_10227,N_10187,N_10047);
nor U10228 (N_10228,N_10011,N_10193);
xnor U10229 (N_10229,N_10015,N_10160);
and U10230 (N_10230,N_10128,N_10088);
xor U10231 (N_10231,N_10190,N_10178);
xnor U10232 (N_10232,N_10167,N_10096);
nor U10233 (N_10233,N_10165,N_10024);
xor U10234 (N_10234,N_10140,N_10077);
nor U10235 (N_10235,N_10052,N_10023);
or U10236 (N_10236,N_10103,N_10145);
or U10237 (N_10237,N_10019,N_10054);
or U10238 (N_10238,N_10120,N_10149);
nand U10239 (N_10239,N_10152,N_10184);
xnor U10240 (N_10240,N_10138,N_10173);
xnor U10241 (N_10241,N_10002,N_10136);
xnor U10242 (N_10242,N_10084,N_10158);
and U10243 (N_10243,N_10194,N_10174);
and U10244 (N_10244,N_10036,N_10021);
nor U10245 (N_10245,N_10179,N_10127);
xor U10246 (N_10246,N_10106,N_10129);
and U10247 (N_10247,N_10001,N_10101);
nor U10248 (N_10248,N_10112,N_10150);
nor U10249 (N_10249,N_10176,N_10141);
xnor U10250 (N_10250,N_10130,N_10161);
nand U10251 (N_10251,N_10041,N_10196);
nor U10252 (N_10252,N_10029,N_10076);
xor U10253 (N_10253,N_10007,N_10010);
nand U10254 (N_10254,N_10147,N_10108);
xnor U10255 (N_10255,N_10125,N_10181);
and U10256 (N_10256,N_10030,N_10185);
or U10257 (N_10257,N_10114,N_10171);
nand U10258 (N_10258,N_10006,N_10025);
nor U10259 (N_10259,N_10099,N_10072);
and U10260 (N_10260,N_10139,N_10033);
and U10261 (N_10261,N_10113,N_10104);
and U10262 (N_10262,N_10197,N_10083);
and U10263 (N_10263,N_10070,N_10048);
or U10264 (N_10264,N_10039,N_10004);
xnor U10265 (N_10265,N_10163,N_10031);
or U10266 (N_10266,N_10049,N_10199);
nor U10267 (N_10267,N_10170,N_10045);
and U10268 (N_10268,N_10080,N_10180);
nor U10269 (N_10269,N_10134,N_10122);
nor U10270 (N_10270,N_10148,N_10097);
nor U10271 (N_10271,N_10177,N_10110);
xnor U10272 (N_10272,N_10192,N_10124);
and U10273 (N_10273,N_10089,N_10155);
xnor U10274 (N_10274,N_10143,N_10003);
nor U10275 (N_10275,N_10117,N_10068);
nand U10276 (N_10276,N_10109,N_10053);
nor U10277 (N_10277,N_10085,N_10166);
nand U10278 (N_10278,N_10093,N_10098);
xnor U10279 (N_10279,N_10043,N_10183);
or U10280 (N_10280,N_10172,N_10121);
nand U10281 (N_10281,N_10133,N_10046);
and U10282 (N_10282,N_10078,N_10107);
or U10283 (N_10283,N_10115,N_10012);
nor U10284 (N_10284,N_10198,N_10042);
or U10285 (N_10285,N_10151,N_10066);
and U10286 (N_10286,N_10189,N_10062);
and U10287 (N_10287,N_10126,N_10051);
xor U10288 (N_10288,N_10095,N_10082);
nand U10289 (N_10289,N_10186,N_10009);
or U10290 (N_10290,N_10116,N_10086);
and U10291 (N_10291,N_10058,N_10182);
and U10292 (N_10292,N_10013,N_10144);
nand U10293 (N_10293,N_10168,N_10027);
or U10294 (N_10294,N_10059,N_10018);
nor U10295 (N_10295,N_10091,N_10135);
xor U10296 (N_10296,N_10005,N_10032);
or U10297 (N_10297,N_10020,N_10191);
xnor U10298 (N_10298,N_10118,N_10016);
or U10299 (N_10299,N_10028,N_10074);
or U10300 (N_10300,N_10091,N_10160);
nor U10301 (N_10301,N_10103,N_10150);
nor U10302 (N_10302,N_10040,N_10067);
nand U10303 (N_10303,N_10122,N_10171);
xor U10304 (N_10304,N_10102,N_10020);
or U10305 (N_10305,N_10105,N_10089);
xor U10306 (N_10306,N_10000,N_10154);
nand U10307 (N_10307,N_10189,N_10097);
or U10308 (N_10308,N_10082,N_10022);
xnor U10309 (N_10309,N_10097,N_10173);
or U10310 (N_10310,N_10070,N_10084);
nor U10311 (N_10311,N_10091,N_10143);
nand U10312 (N_10312,N_10136,N_10008);
and U10313 (N_10313,N_10087,N_10112);
xnor U10314 (N_10314,N_10161,N_10107);
and U10315 (N_10315,N_10036,N_10112);
nand U10316 (N_10316,N_10035,N_10151);
nor U10317 (N_10317,N_10092,N_10001);
nand U10318 (N_10318,N_10104,N_10099);
nand U10319 (N_10319,N_10159,N_10096);
xnor U10320 (N_10320,N_10104,N_10160);
nand U10321 (N_10321,N_10174,N_10010);
nor U10322 (N_10322,N_10140,N_10047);
nand U10323 (N_10323,N_10163,N_10150);
nand U10324 (N_10324,N_10123,N_10148);
nand U10325 (N_10325,N_10113,N_10176);
and U10326 (N_10326,N_10025,N_10059);
or U10327 (N_10327,N_10140,N_10132);
and U10328 (N_10328,N_10103,N_10122);
nand U10329 (N_10329,N_10165,N_10127);
xnor U10330 (N_10330,N_10030,N_10191);
nor U10331 (N_10331,N_10153,N_10154);
xnor U10332 (N_10332,N_10069,N_10187);
nand U10333 (N_10333,N_10066,N_10037);
xor U10334 (N_10334,N_10164,N_10029);
or U10335 (N_10335,N_10097,N_10165);
nor U10336 (N_10336,N_10127,N_10146);
and U10337 (N_10337,N_10012,N_10008);
nor U10338 (N_10338,N_10071,N_10171);
and U10339 (N_10339,N_10028,N_10006);
nand U10340 (N_10340,N_10097,N_10035);
nor U10341 (N_10341,N_10184,N_10062);
xor U10342 (N_10342,N_10175,N_10037);
xor U10343 (N_10343,N_10019,N_10088);
nor U10344 (N_10344,N_10128,N_10031);
nor U10345 (N_10345,N_10105,N_10041);
and U10346 (N_10346,N_10131,N_10094);
and U10347 (N_10347,N_10020,N_10024);
nand U10348 (N_10348,N_10011,N_10148);
nor U10349 (N_10349,N_10172,N_10171);
or U10350 (N_10350,N_10122,N_10077);
nand U10351 (N_10351,N_10057,N_10008);
nand U10352 (N_10352,N_10016,N_10104);
nand U10353 (N_10353,N_10081,N_10171);
and U10354 (N_10354,N_10088,N_10176);
nor U10355 (N_10355,N_10128,N_10062);
xor U10356 (N_10356,N_10184,N_10123);
and U10357 (N_10357,N_10120,N_10099);
or U10358 (N_10358,N_10087,N_10194);
nor U10359 (N_10359,N_10062,N_10086);
nand U10360 (N_10360,N_10016,N_10042);
or U10361 (N_10361,N_10024,N_10109);
nand U10362 (N_10362,N_10039,N_10124);
or U10363 (N_10363,N_10170,N_10123);
or U10364 (N_10364,N_10104,N_10098);
and U10365 (N_10365,N_10134,N_10060);
or U10366 (N_10366,N_10198,N_10181);
and U10367 (N_10367,N_10078,N_10062);
nand U10368 (N_10368,N_10123,N_10063);
or U10369 (N_10369,N_10154,N_10126);
and U10370 (N_10370,N_10021,N_10089);
nand U10371 (N_10371,N_10092,N_10080);
and U10372 (N_10372,N_10035,N_10149);
nand U10373 (N_10373,N_10120,N_10050);
nor U10374 (N_10374,N_10047,N_10115);
nor U10375 (N_10375,N_10036,N_10069);
and U10376 (N_10376,N_10017,N_10103);
and U10377 (N_10377,N_10074,N_10033);
or U10378 (N_10378,N_10059,N_10009);
nand U10379 (N_10379,N_10014,N_10030);
and U10380 (N_10380,N_10102,N_10130);
nor U10381 (N_10381,N_10146,N_10082);
nand U10382 (N_10382,N_10017,N_10165);
xnor U10383 (N_10383,N_10054,N_10061);
nor U10384 (N_10384,N_10071,N_10132);
or U10385 (N_10385,N_10196,N_10106);
nor U10386 (N_10386,N_10075,N_10083);
nand U10387 (N_10387,N_10089,N_10064);
or U10388 (N_10388,N_10098,N_10145);
or U10389 (N_10389,N_10121,N_10127);
nand U10390 (N_10390,N_10092,N_10122);
and U10391 (N_10391,N_10109,N_10043);
nor U10392 (N_10392,N_10194,N_10158);
or U10393 (N_10393,N_10173,N_10031);
xor U10394 (N_10394,N_10058,N_10152);
or U10395 (N_10395,N_10076,N_10185);
xor U10396 (N_10396,N_10186,N_10160);
xor U10397 (N_10397,N_10189,N_10104);
xnor U10398 (N_10398,N_10010,N_10018);
or U10399 (N_10399,N_10150,N_10194);
xor U10400 (N_10400,N_10240,N_10366);
and U10401 (N_10401,N_10320,N_10297);
xnor U10402 (N_10402,N_10383,N_10245);
nor U10403 (N_10403,N_10347,N_10292);
and U10404 (N_10404,N_10284,N_10214);
or U10405 (N_10405,N_10231,N_10340);
xor U10406 (N_10406,N_10215,N_10211);
or U10407 (N_10407,N_10207,N_10316);
nand U10408 (N_10408,N_10296,N_10308);
nand U10409 (N_10409,N_10398,N_10326);
xor U10410 (N_10410,N_10254,N_10218);
xor U10411 (N_10411,N_10270,N_10362);
and U10412 (N_10412,N_10235,N_10293);
xor U10413 (N_10413,N_10222,N_10229);
or U10414 (N_10414,N_10336,N_10375);
xor U10415 (N_10415,N_10325,N_10249);
and U10416 (N_10416,N_10247,N_10387);
and U10417 (N_10417,N_10321,N_10312);
and U10418 (N_10418,N_10352,N_10223);
xor U10419 (N_10419,N_10232,N_10217);
xnor U10420 (N_10420,N_10390,N_10323);
or U10421 (N_10421,N_10210,N_10283);
xor U10422 (N_10422,N_10230,N_10276);
nor U10423 (N_10423,N_10313,N_10342);
xnor U10424 (N_10424,N_10286,N_10318);
and U10425 (N_10425,N_10365,N_10274);
nand U10426 (N_10426,N_10327,N_10275);
nor U10427 (N_10427,N_10324,N_10343);
and U10428 (N_10428,N_10392,N_10221);
nor U10429 (N_10429,N_10259,N_10373);
and U10430 (N_10430,N_10379,N_10268);
and U10431 (N_10431,N_10309,N_10233);
and U10432 (N_10432,N_10302,N_10315);
or U10433 (N_10433,N_10278,N_10306);
nor U10434 (N_10434,N_10220,N_10279);
nand U10435 (N_10435,N_10380,N_10291);
nand U10436 (N_10436,N_10359,N_10317);
xor U10437 (N_10437,N_10346,N_10310);
and U10438 (N_10438,N_10290,N_10258);
xor U10439 (N_10439,N_10226,N_10260);
and U10440 (N_10440,N_10396,N_10386);
nor U10441 (N_10441,N_10267,N_10202);
nand U10442 (N_10442,N_10227,N_10266);
and U10443 (N_10443,N_10394,N_10225);
and U10444 (N_10444,N_10397,N_10388);
nor U10445 (N_10445,N_10361,N_10219);
nand U10446 (N_10446,N_10355,N_10305);
nor U10447 (N_10447,N_10204,N_10332);
nand U10448 (N_10448,N_10206,N_10234);
nor U10449 (N_10449,N_10261,N_10281);
and U10450 (N_10450,N_10263,N_10289);
and U10451 (N_10451,N_10333,N_10307);
xor U10452 (N_10452,N_10213,N_10371);
xor U10453 (N_10453,N_10212,N_10242);
xnor U10454 (N_10454,N_10354,N_10244);
and U10455 (N_10455,N_10271,N_10304);
nand U10456 (N_10456,N_10282,N_10228);
and U10457 (N_10457,N_10369,N_10368);
nor U10458 (N_10458,N_10294,N_10395);
nand U10459 (N_10459,N_10350,N_10280);
nand U10460 (N_10460,N_10273,N_10262);
nand U10461 (N_10461,N_10248,N_10328);
nor U10462 (N_10462,N_10377,N_10238);
nand U10463 (N_10463,N_10358,N_10364);
nand U10464 (N_10464,N_10237,N_10329);
nand U10465 (N_10465,N_10356,N_10295);
and U10466 (N_10466,N_10391,N_10341);
or U10467 (N_10467,N_10224,N_10251);
nand U10468 (N_10468,N_10385,N_10250);
or U10469 (N_10469,N_10301,N_10216);
nor U10470 (N_10470,N_10298,N_10209);
nand U10471 (N_10471,N_10239,N_10393);
nand U10472 (N_10472,N_10338,N_10353);
or U10473 (N_10473,N_10330,N_10372);
nor U10474 (N_10474,N_10264,N_10288);
and U10475 (N_10475,N_10208,N_10370);
and U10476 (N_10476,N_10272,N_10382);
nor U10477 (N_10477,N_10335,N_10265);
nor U10478 (N_10478,N_10381,N_10351);
nor U10479 (N_10479,N_10389,N_10331);
and U10480 (N_10480,N_10344,N_10201);
xor U10481 (N_10481,N_10256,N_10399);
or U10482 (N_10482,N_10334,N_10339);
or U10483 (N_10483,N_10205,N_10374);
and U10484 (N_10484,N_10243,N_10348);
nor U10485 (N_10485,N_10303,N_10314);
nand U10486 (N_10486,N_10378,N_10285);
and U10487 (N_10487,N_10277,N_10300);
nor U10488 (N_10488,N_10246,N_10269);
nor U10489 (N_10489,N_10357,N_10376);
and U10490 (N_10490,N_10363,N_10253);
nor U10491 (N_10491,N_10257,N_10319);
and U10492 (N_10492,N_10384,N_10322);
nor U10493 (N_10493,N_10311,N_10252);
or U10494 (N_10494,N_10345,N_10241);
nor U10495 (N_10495,N_10360,N_10200);
xor U10496 (N_10496,N_10349,N_10236);
nand U10497 (N_10497,N_10287,N_10337);
nand U10498 (N_10498,N_10203,N_10255);
nor U10499 (N_10499,N_10367,N_10299);
and U10500 (N_10500,N_10286,N_10338);
xnor U10501 (N_10501,N_10233,N_10228);
or U10502 (N_10502,N_10361,N_10267);
or U10503 (N_10503,N_10364,N_10338);
and U10504 (N_10504,N_10248,N_10259);
and U10505 (N_10505,N_10305,N_10233);
nand U10506 (N_10506,N_10305,N_10368);
or U10507 (N_10507,N_10353,N_10394);
xor U10508 (N_10508,N_10234,N_10369);
xor U10509 (N_10509,N_10374,N_10207);
or U10510 (N_10510,N_10235,N_10328);
nor U10511 (N_10511,N_10273,N_10224);
and U10512 (N_10512,N_10241,N_10272);
or U10513 (N_10513,N_10256,N_10254);
nor U10514 (N_10514,N_10381,N_10253);
xnor U10515 (N_10515,N_10377,N_10354);
xor U10516 (N_10516,N_10263,N_10250);
and U10517 (N_10517,N_10398,N_10282);
or U10518 (N_10518,N_10306,N_10284);
xnor U10519 (N_10519,N_10309,N_10323);
xor U10520 (N_10520,N_10242,N_10231);
nor U10521 (N_10521,N_10240,N_10312);
nand U10522 (N_10522,N_10316,N_10349);
xor U10523 (N_10523,N_10206,N_10225);
nor U10524 (N_10524,N_10297,N_10235);
nor U10525 (N_10525,N_10315,N_10325);
nor U10526 (N_10526,N_10244,N_10239);
xor U10527 (N_10527,N_10311,N_10207);
and U10528 (N_10528,N_10266,N_10259);
nor U10529 (N_10529,N_10332,N_10291);
xnor U10530 (N_10530,N_10339,N_10275);
nor U10531 (N_10531,N_10298,N_10293);
xor U10532 (N_10532,N_10348,N_10278);
nand U10533 (N_10533,N_10304,N_10204);
nand U10534 (N_10534,N_10266,N_10356);
or U10535 (N_10535,N_10362,N_10200);
and U10536 (N_10536,N_10248,N_10296);
and U10537 (N_10537,N_10274,N_10289);
or U10538 (N_10538,N_10344,N_10215);
nor U10539 (N_10539,N_10224,N_10287);
nor U10540 (N_10540,N_10239,N_10353);
and U10541 (N_10541,N_10289,N_10331);
or U10542 (N_10542,N_10272,N_10307);
nor U10543 (N_10543,N_10367,N_10276);
xor U10544 (N_10544,N_10212,N_10279);
nand U10545 (N_10545,N_10340,N_10398);
nand U10546 (N_10546,N_10370,N_10323);
nand U10547 (N_10547,N_10263,N_10312);
xor U10548 (N_10548,N_10237,N_10305);
and U10549 (N_10549,N_10327,N_10263);
or U10550 (N_10550,N_10247,N_10253);
or U10551 (N_10551,N_10227,N_10348);
or U10552 (N_10552,N_10271,N_10398);
and U10553 (N_10553,N_10252,N_10359);
xnor U10554 (N_10554,N_10319,N_10348);
or U10555 (N_10555,N_10343,N_10237);
nand U10556 (N_10556,N_10385,N_10234);
and U10557 (N_10557,N_10292,N_10287);
or U10558 (N_10558,N_10284,N_10366);
or U10559 (N_10559,N_10349,N_10232);
nand U10560 (N_10560,N_10324,N_10364);
nor U10561 (N_10561,N_10372,N_10365);
nor U10562 (N_10562,N_10323,N_10235);
nand U10563 (N_10563,N_10372,N_10229);
and U10564 (N_10564,N_10231,N_10309);
and U10565 (N_10565,N_10209,N_10332);
nand U10566 (N_10566,N_10315,N_10337);
or U10567 (N_10567,N_10216,N_10351);
xnor U10568 (N_10568,N_10272,N_10341);
xor U10569 (N_10569,N_10276,N_10237);
xnor U10570 (N_10570,N_10212,N_10382);
xor U10571 (N_10571,N_10366,N_10390);
nor U10572 (N_10572,N_10295,N_10336);
nand U10573 (N_10573,N_10202,N_10254);
or U10574 (N_10574,N_10364,N_10297);
xnor U10575 (N_10575,N_10245,N_10315);
nor U10576 (N_10576,N_10372,N_10219);
nand U10577 (N_10577,N_10213,N_10386);
nor U10578 (N_10578,N_10382,N_10265);
xnor U10579 (N_10579,N_10230,N_10298);
xnor U10580 (N_10580,N_10303,N_10322);
or U10581 (N_10581,N_10377,N_10274);
xor U10582 (N_10582,N_10269,N_10309);
and U10583 (N_10583,N_10231,N_10355);
xnor U10584 (N_10584,N_10313,N_10378);
xnor U10585 (N_10585,N_10334,N_10307);
nand U10586 (N_10586,N_10256,N_10336);
nor U10587 (N_10587,N_10326,N_10284);
nand U10588 (N_10588,N_10381,N_10341);
nor U10589 (N_10589,N_10396,N_10289);
and U10590 (N_10590,N_10386,N_10352);
xnor U10591 (N_10591,N_10372,N_10215);
nand U10592 (N_10592,N_10290,N_10233);
and U10593 (N_10593,N_10283,N_10234);
nand U10594 (N_10594,N_10201,N_10367);
nand U10595 (N_10595,N_10223,N_10302);
nor U10596 (N_10596,N_10393,N_10329);
nand U10597 (N_10597,N_10381,N_10302);
nor U10598 (N_10598,N_10200,N_10240);
and U10599 (N_10599,N_10210,N_10205);
nand U10600 (N_10600,N_10438,N_10542);
and U10601 (N_10601,N_10441,N_10589);
nand U10602 (N_10602,N_10491,N_10577);
or U10603 (N_10603,N_10567,N_10562);
nand U10604 (N_10604,N_10578,N_10476);
nor U10605 (N_10605,N_10473,N_10457);
and U10606 (N_10606,N_10581,N_10512);
nor U10607 (N_10607,N_10454,N_10549);
nand U10608 (N_10608,N_10516,N_10499);
xnor U10609 (N_10609,N_10488,N_10430);
nand U10610 (N_10610,N_10460,N_10530);
xnor U10611 (N_10611,N_10495,N_10422);
or U10612 (N_10612,N_10467,N_10547);
nor U10613 (N_10613,N_10555,N_10568);
nor U10614 (N_10614,N_10481,N_10558);
and U10615 (N_10615,N_10545,N_10400);
nor U10616 (N_10616,N_10576,N_10415);
and U10617 (N_10617,N_10543,N_10424);
or U10618 (N_10618,N_10406,N_10446);
xor U10619 (N_10619,N_10437,N_10518);
nor U10620 (N_10620,N_10540,N_10408);
or U10621 (N_10621,N_10557,N_10447);
nand U10622 (N_10622,N_10469,N_10486);
or U10623 (N_10623,N_10598,N_10405);
nand U10624 (N_10624,N_10500,N_10551);
and U10625 (N_10625,N_10592,N_10514);
nor U10626 (N_10626,N_10421,N_10480);
xor U10627 (N_10627,N_10450,N_10556);
and U10628 (N_10628,N_10490,N_10536);
nand U10629 (N_10629,N_10564,N_10599);
xor U10630 (N_10630,N_10523,N_10475);
nand U10631 (N_10631,N_10501,N_10432);
nand U10632 (N_10632,N_10413,N_10487);
nor U10633 (N_10633,N_10571,N_10485);
nor U10634 (N_10634,N_10559,N_10489);
or U10635 (N_10635,N_10584,N_10456);
nand U10636 (N_10636,N_10449,N_10402);
nand U10637 (N_10637,N_10409,N_10461);
nor U10638 (N_10638,N_10496,N_10515);
or U10639 (N_10639,N_10570,N_10572);
nand U10640 (N_10640,N_10426,N_10463);
or U10641 (N_10641,N_10580,N_10579);
nand U10642 (N_10642,N_10539,N_10504);
xor U10643 (N_10643,N_10428,N_10417);
or U10644 (N_10644,N_10464,N_10586);
nor U10645 (N_10645,N_10513,N_10484);
and U10646 (N_10646,N_10565,N_10596);
xor U10647 (N_10647,N_10458,N_10591);
xor U10648 (N_10648,N_10433,N_10595);
nor U10649 (N_10649,N_10535,N_10552);
or U10650 (N_10650,N_10532,N_10472);
xnor U10651 (N_10651,N_10493,N_10478);
and U10652 (N_10652,N_10597,N_10548);
xor U10653 (N_10653,N_10554,N_10416);
xnor U10654 (N_10654,N_10550,N_10507);
and U10655 (N_10655,N_10404,N_10560);
xor U10656 (N_10656,N_10418,N_10414);
xnor U10657 (N_10657,N_10519,N_10517);
and U10658 (N_10658,N_10455,N_10590);
nor U10659 (N_10659,N_10511,N_10588);
nand U10660 (N_10660,N_10401,N_10462);
and U10661 (N_10661,N_10498,N_10444);
or U10662 (N_10662,N_10448,N_10453);
xnor U10663 (N_10663,N_10582,N_10510);
or U10664 (N_10664,N_10520,N_10420);
nor U10665 (N_10665,N_10429,N_10479);
nor U10666 (N_10666,N_10522,N_10587);
or U10667 (N_10667,N_10427,N_10583);
xnor U10668 (N_10668,N_10497,N_10492);
or U10669 (N_10669,N_10412,N_10440);
nor U10670 (N_10670,N_10419,N_10544);
or U10671 (N_10671,N_10494,N_10435);
xnor U10672 (N_10672,N_10573,N_10431);
or U10673 (N_10673,N_10531,N_10533);
and U10674 (N_10674,N_10529,N_10509);
and U10675 (N_10675,N_10541,N_10527);
nand U10676 (N_10676,N_10521,N_10425);
xnor U10677 (N_10677,N_10575,N_10526);
or U10678 (N_10678,N_10483,N_10525);
nor U10679 (N_10679,N_10471,N_10445);
nand U10680 (N_10680,N_10411,N_10434);
nor U10681 (N_10681,N_10561,N_10534);
and U10682 (N_10682,N_10403,N_10442);
nor U10683 (N_10683,N_10528,N_10436);
nand U10684 (N_10684,N_10506,N_10466);
xnor U10685 (N_10685,N_10593,N_10574);
and U10686 (N_10686,N_10470,N_10474);
and U10687 (N_10687,N_10594,N_10566);
and U10688 (N_10688,N_10537,N_10505);
and U10689 (N_10689,N_10407,N_10443);
nor U10690 (N_10690,N_10503,N_10451);
nand U10691 (N_10691,N_10563,N_10439);
nor U10692 (N_10692,N_10468,N_10569);
or U10693 (N_10693,N_10546,N_10538);
and U10694 (N_10694,N_10423,N_10482);
xor U10695 (N_10695,N_10508,N_10452);
and U10696 (N_10696,N_10477,N_10459);
nor U10697 (N_10697,N_10465,N_10585);
or U10698 (N_10698,N_10524,N_10502);
or U10699 (N_10699,N_10553,N_10410);
nand U10700 (N_10700,N_10424,N_10563);
nand U10701 (N_10701,N_10568,N_10419);
xnor U10702 (N_10702,N_10458,N_10413);
xor U10703 (N_10703,N_10464,N_10414);
nand U10704 (N_10704,N_10516,N_10557);
nand U10705 (N_10705,N_10533,N_10443);
nand U10706 (N_10706,N_10448,N_10545);
or U10707 (N_10707,N_10449,N_10556);
nand U10708 (N_10708,N_10506,N_10553);
xor U10709 (N_10709,N_10473,N_10437);
nand U10710 (N_10710,N_10429,N_10461);
nand U10711 (N_10711,N_10589,N_10536);
nor U10712 (N_10712,N_10464,N_10584);
or U10713 (N_10713,N_10506,N_10426);
nand U10714 (N_10714,N_10531,N_10484);
and U10715 (N_10715,N_10517,N_10560);
or U10716 (N_10716,N_10562,N_10457);
nor U10717 (N_10717,N_10545,N_10470);
xor U10718 (N_10718,N_10473,N_10477);
xor U10719 (N_10719,N_10481,N_10598);
nand U10720 (N_10720,N_10421,N_10588);
and U10721 (N_10721,N_10524,N_10493);
xnor U10722 (N_10722,N_10488,N_10483);
and U10723 (N_10723,N_10595,N_10493);
and U10724 (N_10724,N_10580,N_10457);
xnor U10725 (N_10725,N_10448,N_10598);
xnor U10726 (N_10726,N_10544,N_10506);
nand U10727 (N_10727,N_10422,N_10526);
or U10728 (N_10728,N_10487,N_10560);
xor U10729 (N_10729,N_10475,N_10443);
nor U10730 (N_10730,N_10572,N_10533);
nor U10731 (N_10731,N_10472,N_10486);
nor U10732 (N_10732,N_10547,N_10587);
or U10733 (N_10733,N_10564,N_10443);
or U10734 (N_10734,N_10541,N_10592);
or U10735 (N_10735,N_10485,N_10531);
and U10736 (N_10736,N_10587,N_10579);
or U10737 (N_10737,N_10578,N_10565);
nand U10738 (N_10738,N_10516,N_10476);
xnor U10739 (N_10739,N_10438,N_10509);
xnor U10740 (N_10740,N_10561,N_10526);
xnor U10741 (N_10741,N_10505,N_10535);
xor U10742 (N_10742,N_10533,N_10535);
or U10743 (N_10743,N_10532,N_10599);
or U10744 (N_10744,N_10466,N_10437);
nor U10745 (N_10745,N_10520,N_10576);
nand U10746 (N_10746,N_10451,N_10559);
nor U10747 (N_10747,N_10402,N_10590);
nor U10748 (N_10748,N_10407,N_10496);
or U10749 (N_10749,N_10575,N_10492);
xnor U10750 (N_10750,N_10422,N_10508);
nor U10751 (N_10751,N_10468,N_10527);
xnor U10752 (N_10752,N_10543,N_10531);
or U10753 (N_10753,N_10470,N_10468);
and U10754 (N_10754,N_10473,N_10495);
xnor U10755 (N_10755,N_10499,N_10461);
nor U10756 (N_10756,N_10589,N_10534);
nor U10757 (N_10757,N_10490,N_10483);
and U10758 (N_10758,N_10597,N_10465);
nand U10759 (N_10759,N_10407,N_10540);
nand U10760 (N_10760,N_10510,N_10470);
nor U10761 (N_10761,N_10554,N_10598);
and U10762 (N_10762,N_10538,N_10553);
nor U10763 (N_10763,N_10543,N_10528);
or U10764 (N_10764,N_10461,N_10465);
or U10765 (N_10765,N_10509,N_10440);
and U10766 (N_10766,N_10430,N_10478);
nand U10767 (N_10767,N_10511,N_10522);
or U10768 (N_10768,N_10536,N_10415);
or U10769 (N_10769,N_10433,N_10459);
and U10770 (N_10770,N_10500,N_10517);
nor U10771 (N_10771,N_10578,N_10518);
or U10772 (N_10772,N_10485,N_10460);
nor U10773 (N_10773,N_10566,N_10439);
or U10774 (N_10774,N_10480,N_10531);
or U10775 (N_10775,N_10449,N_10401);
and U10776 (N_10776,N_10547,N_10525);
nand U10777 (N_10777,N_10468,N_10402);
nand U10778 (N_10778,N_10496,N_10454);
xor U10779 (N_10779,N_10446,N_10561);
nand U10780 (N_10780,N_10430,N_10577);
nor U10781 (N_10781,N_10517,N_10486);
and U10782 (N_10782,N_10453,N_10597);
or U10783 (N_10783,N_10401,N_10591);
or U10784 (N_10784,N_10436,N_10521);
or U10785 (N_10785,N_10568,N_10436);
nor U10786 (N_10786,N_10530,N_10432);
nand U10787 (N_10787,N_10447,N_10506);
and U10788 (N_10788,N_10460,N_10473);
nand U10789 (N_10789,N_10570,N_10561);
nand U10790 (N_10790,N_10517,N_10451);
nor U10791 (N_10791,N_10420,N_10595);
nor U10792 (N_10792,N_10459,N_10460);
nor U10793 (N_10793,N_10556,N_10486);
and U10794 (N_10794,N_10470,N_10475);
nand U10795 (N_10795,N_10482,N_10522);
nor U10796 (N_10796,N_10434,N_10522);
nor U10797 (N_10797,N_10448,N_10435);
nand U10798 (N_10798,N_10529,N_10401);
or U10799 (N_10799,N_10550,N_10455);
nand U10800 (N_10800,N_10664,N_10675);
xnor U10801 (N_10801,N_10603,N_10642);
nand U10802 (N_10802,N_10606,N_10608);
or U10803 (N_10803,N_10754,N_10689);
xnor U10804 (N_10804,N_10637,N_10601);
and U10805 (N_10805,N_10784,N_10658);
xnor U10806 (N_10806,N_10772,N_10654);
or U10807 (N_10807,N_10697,N_10794);
or U10808 (N_10808,N_10778,N_10727);
xor U10809 (N_10809,N_10706,N_10635);
nor U10810 (N_10810,N_10692,N_10752);
or U10811 (N_10811,N_10701,N_10634);
or U10812 (N_10812,N_10703,N_10735);
and U10813 (N_10813,N_10653,N_10681);
nor U10814 (N_10814,N_10788,N_10655);
nand U10815 (N_10815,N_10704,N_10650);
and U10816 (N_10816,N_10748,N_10696);
nand U10817 (N_10817,N_10728,N_10607);
nor U10818 (N_10818,N_10707,N_10604);
xor U10819 (N_10819,N_10764,N_10737);
or U10820 (N_10820,N_10734,N_10739);
and U10821 (N_10821,N_10765,N_10649);
nand U10822 (N_10822,N_10648,N_10633);
xnor U10823 (N_10823,N_10729,N_10796);
nand U10824 (N_10824,N_10719,N_10717);
xor U10825 (N_10825,N_10647,N_10676);
nor U10826 (N_10826,N_10611,N_10720);
nand U10827 (N_10827,N_10627,N_10759);
nand U10828 (N_10828,N_10741,N_10605);
or U10829 (N_10829,N_10708,N_10693);
or U10830 (N_10830,N_10685,N_10745);
nand U10831 (N_10831,N_10652,N_10700);
xor U10832 (N_10832,N_10631,N_10698);
or U10833 (N_10833,N_10711,N_10666);
and U10834 (N_10834,N_10699,N_10616);
nand U10835 (N_10835,N_10623,N_10638);
and U10836 (N_10836,N_10673,N_10686);
or U10837 (N_10837,N_10758,N_10755);
nand U10838 (N_10838,N_10742,N_10746);
or U10839 (N_10839,N_10756,N_10643);
xor U10840 (N_10840,N_10640,N_10690);
nand U10841 (N_10841,N_10731,N_10750);
or U10842 (N_10842,N_10799,N_10789);
xor U10843 (N_10843,N_10667,N_10702);
nor U10844 (N_10844,N_10757,N_10776);
xnor U10845 (N_10845,N_10663,N_10782);
xnor U10846 (N_10846,N_10670,N_10783);
nand U10847 (N_10847,N_10730,N_10678);
nor U10848 (N_10848,N_10715,N_10680);
nand U10849 (N_10849,N_10695,N_10621);
and U10850 (N_10850,N_10618,N_10726);
or U10851 (N_10851,N_10786,N_10614);
and U10852 (N_10852,N_10682,N_10615);
xor U10853 (N_10853,N_10645,N_10660);
xnor U10854 (N_10854,N_10798,N_10684);
and U10855 (N_10855,N_10629,N_10723);
or U10856 (N_10856,N_10749,N_10716);
nand U10857 (N_10857,N_10795,N_10714);
or U10858 (N_10858,N_10722,N_10612);
or U10859 (N_10859,N_10777,N_10761);
xnor U10860 (N_10860,N_10600,N_10767);
nand U10861 (N_10861,N_10733,N_10773);
or U10862 (N_10862,N_10781,N_10792);
nand U10863 (N_10863,N_10641,N_10713);
xnor U10864 (N_10864,N_10646,N_10787);
or U10865 (N_10865,N_10766,N_10768);
nand U10866 (N_10866,N_10677,N_10724);
and U10867 (N_10867,N_10740,N_10628);
xor U10868 (N_10868,N_10625,N_10622);
nor U10869 (N_10869,N_10718,N_10738);
and U10870 (N_10870,N_10709,N_10639);
nor U10871 (N_10871,N_10705,N_10632);
nor U10872 (N_10872,N_10657,N_10797);
or U10873 (N_10873,N_10683,N_10617);
nand U10874 (N_10874,N_10785,N_10774);
xnor U10875 (N_10875,N_10779,N_10688);
or U10876 (N_10876,N_10602,N_10791);
xor U10877 (N_10877,N_10636,N_10669);
nand U10878 (N_10878,N_10651,N_10644);
or U10879 (N_10879,N_10775,N_10736);
and U10880 (N_10880,N_10674,N_10610);
or U10881 (N_10881,N_10626,N_10656);
or U10882 (N_10882,N_10762,N_10747);
and U10883 (N_10883,N_10790,N_10620);
nor U10884 (N_10884,N_10694,N_10712);
nor U10885 (N_10885,N_10793,N_10609);
nor U10886 (N_10886,N_10721,N_10671);
nor U10887 (N_10887,N_10662,N_10630);
nor U10888 (N_10888,N_10624,N_10691);
and U10889 (N_10889,N_10751,N_10770);
and U10890 (N_10890,N_10771,N_10753);
xor U10891 (N_10891,N_10659,N_10668);
xor U10892 (N_10892,N_10613,N_10710);
or U10893 (N_10893,N_10665,N_10760);
nor U10894 (N_10894,N_10661,N_10769);
or U10895 (N_10895,N_10687,N_10679);
xor U10896 (N_10896,N_10763,N_10780);
or U10897 (N_10897,N_10672,N_10619);
xor U10898 (N_10898,N_10725,N_10743);
nor U10899 (N_10899,N_10744,N_10732);
or U10900 (N_10900,N_10732,N_10606);
nor U10901 (N_10901,N_10652,N_10750);
or U10902 (N_10902,N_10628,N_10696);
nor U10903 (N_10903,N_10674,N_10777);
or U10904 (N_10904,N_10697,N_10618);
nand U10905 (N_10905,N_10625,N_10740);
xnor U10906 (N_10906,N_10671,N_10698);
xor U10907 (N_10907,N_10706,N_10792);
or U10908 (N_10908,N_10795,N_10685);
nor U10909 (N_10909,N_10632,N_10778);
or U10910 (N_10910,N_10688,N_10773);
nand U10911 (N_10911,N_10671,N_10752);
or U10912 (N_10912,N_10701,N_10792);
nor U10913 (N_10913,N_10634,N_10650);
nor U10914 (N_10914,N_10621,N_10629);
nand U10915 (N_10915,N_10686,N_10741);
nand U10916 (N_10916,N_10740,N_10626);
and U10917 (N_10917,N_10745,N_10698);
nand U10918 (N_10918,N_10759,N_10793);
nand U10919 (N_10919,N_10680,N_10698);
nand U10920 (N_10920,N_10715,N_10756);
nor U10921 (N_10921,N_10622,N_10668);
and U10922 (N_10922,N_10614,N_10646);
or U10923 (N_10923,N_10619,N_10674);
or U10924 (N_10924,N_10789,N_10795);
and U10925 (N_10925,N_10677,N_10668);
and U10926 (N_10926,N_10638,N_10676);
xor U10927 (N_10927,N_10742,N_10759);
nor U10928 (N_10928,N_10656,N_10667);
xor U10929 (N_10929,N_10715,N_10656);
xor U10930 (N_10930,N_10748,N_10698);
nor U10931 (N_10931,N_10736,N_10604);
and U10932 (N_10932,N_10766,N_10608);
nand U10933 (N_10933,N_10721,N_10606);
nand U10934 (N_10934,N_10679,N_10730);
and U10935 (N_10935,N_10645,N_10729);
nor U10936 (N_10936,N_10702,N_10618);
xor U10937 (N_10937,N_10798,N_10729);
or U10938 (N_10938,N_10744,N_10702);
and U10939 (N_10939,N_10616,N_10775);
and U10940 (N_10940,N_10645,N_10603);
and U10941 (N_10941,N_10739,N_10747);
nor U10942 (N_10942,N_10681,N_10680);
and U10943 (N_10943,N_10698,N_10791);
nor U10944 (N_10944,N_10696,N_10772);
and U10945 (N_10945,N_10653,N_10624);
and U10946 (N_10946,N_10616,N_10683);
and U10947 (N_10947,N_10798,N_10788);
nand U10948 (N_10948,N_10678,N_10600);
nand U10949 (N_10949,N_10768,N_10729);
xnor U10950 (N_10950,N_10771,N_10653);
nand U10951 (N_10951,N_10751,N_10708);
nor U10952 (N_10952,N_10604,N_10621);
nor U10953 (N_10953,N_10738,N_10695);
nand U10954 (N_10954,N_10742,N_10779);
or U10955 (N_10955,N_10756,N_10772);
or U10956 (N_10956,N_10663,N_10778);
and U10957 (N_10957,N_10665,N_10612);
or U10958 (N_10958,N_10614,N_10706);
nor U10959 (N_10959,N_10791,N_10651);
and U10960 (N_10960,N_10734,N_10752);
or U10961 (N_10961,N_10693,N_10746);
nand U10962 (N_10962,N_10648,N_10614);
nand U10963 (N_10963,N_10666,N_10776);
or U10964 (N_10964,N_10791,N_10694);
or U10965 (N_10965,N_10692,N_10741);
nor U10966 (N_10966,N_10788,N_10708);
and U10967 (N_10967,N_10771,N_10605);
nand U10968 (N_10968,N_10643,N_10702);
and U10969 (N_10969,N_10619,N_10709);
nand U10970 (N_10970,N_10715,N_10604);
nand U10971 (N_10971,N_10723,N_10666);
and U10972 (N_10972,N_10629,N_10743);
nand U10973 (N_10973,N_10700,N_10603);
or U10974 (N_10974,N_10679,N_10688);
or U10975 (N_10975,N_10776,N_10739);
nor U10976 (N_10976,N_10613,N_10658);
or U10977 (N_10977,N_10748,N_10745);
xnor U10978 (N_10978,N_10716,N_10731);
xnor U10979 (N_10979,N_10742,N_10639);
nand U10980 (N_10980,N_10790,N_10616);
and U10981 (N_10981,N_10735,N_10794);
xnor U10982 (N_10982,N_10650,N_10703);
nor U10983 (N_10983,N_10688,N_10770);
nand U10984 (N_10984,N_10756,N_10776);
nand U10985 (N_10985,N_10657,N_10775);
nand U10986 (N_10986,N_10799,N_10780);
nor U10987 (N_10987,N_10667,N_10661);
or U10988 (N_10988,N_10771,N_10739);
xor U10989 (N_10989,N_10630,N_10764);
and U10990 (N_10990,N_10642,N_10744);
nand U10991 (N_10991,N_10788,N_10755);
or U10992 (N_10992,N_10693,N_10658);
or U10993 (N_10993,N_10655,N_10757);
nor U10994 (N_10994,N_10603,N_10776);
or U10995 (N_10995,N_10692,N_10781);
and U10996 (N_10996,N_10699,N_10673);
xnor U10997 (N_10997,N_10649,N_10676);
nor U10998 (N_10998,N_10612,N_10756);
nand U10999 (N_10999,N_10713,N_10780);
and U11000 (N_11000,N_10912,N_10986);
nor U11001 (N_11001,N_10960,N_10946);
or U11002 (N_11002,N_10950,N_10804);
nand U11003 (N_11003,N_10840,N_10987);
and U11004 (N_11004,N_10883,N_10981);
xnor U11005 (N_11005,N_10969,N_10818);
xnor U11006 (N_11006,N_10976,N_10909);
nand U11007 (N_11007,N_10989,N_10983);
nor U11008 (N_11008,N_10951,N_10801);
nor U11009 (N_11009,N_10964,N_10844);
xnor U11010 (N_11010,N_10957,N_10884);
xnor U11011 (N_11011,N_10933,N_10822);
xor U11012 (N_11012,N_10811,N_10938);
xnor U11013 (N_11013,N_10955,N_10902);
and U11014 (N_11014,N_10854,N_10991);
or U11015 (N_11015,N_10891,N_10843);
or U11016 (N_11016,N_10863,N_10813);
and U11017 (N_11017,N_10887,N_10925);
or U11018 (N_11018,N_10966,N_10929);
nand U11019 (N_11019,N_10921,N_10927);
nand U11020 (N_11020,N_10807,N_10920);
or U11021 (N_11021,N_10875,N_10958);
and U11022 (N_11022,N_10905,N_10837);
nand U11023 (N_11023,N_10815,N_10903);
and U11024 (N_11024,N_10817,N_10823);
xor U11025 (N_11025,N_10864,N_10900);
and U11026 (N_11026,N_10857,N_10993);
or U11027 (N_11027,N_10935,N_10995);
xnor U11028 (N_11028,N_10810,N_10849);
and U11029 (N_11029,N_10914,N_10972);
nor U11030 (N_11030,N_10835,N_10866);
nor U11031 (N_11031,N_10963,N_10959);
xnor U11032 (N_11032,N_10992,N_10937);
xnor U11033 (N_11033,N_10990,N_10885);
and U11034 (N_11034,N_10907,N_10802);
or U11035 (N_11035,N_10882,N_10880);
nor U11036 (N_11036,N_10994,N_10936);
nor U11037 (N_11037,N_10978,N_10838);
and U11038 (N_11038,N_10879,N_10997);
xnor U11039 (N_11039,N_10824,N_10979);
and U11040 (N_11040,N_10996,N_10839);
nor U11041 (N_11041,N_10834,N_10919);
and U11042 (N_11042,N_10998,N_10874);
xor U11043 (N_11043,N_10825,N_10812);
nor U11044 (N_11044,N_10999,N_10913);
and U11045 (N_11045,N_10806,N_10831);
nor U11046 (N_11046,N_10939,N_10895);
nand U11047 (N_11047,N_10906,N_10865);
nand U11048 (N_11048,N_10872,N_10974);
and U11049 (N_11049,N_10859,N_10856);
xnor U11050 (N_11050,N_10800,N_10878);
xnor U11051 (N_11051,N_10973,N_10977);
and U11052 (N_11052,N_10848,N_10908);
nor U11053 (N_11053,N_10821,N_10982);
nand U11054 (N_11054,N_10965,N_10853);
or U11055 (N_11055,N_10868,N_10949);
nand U11056 (N_11056,N_10968,N_10881);
xnor U11057 (N_11057,N_10894,N_10956);
nand U11058 (N_11058,N_10803,N_10877);
nor U11059 (N_11059,N_10899,N_10918);
or U11060 (N_11060,N_10873,N_10855);
and U11061 (N_11061,N_10869,N_10886);
and U11062 (N_11062,N_10829,N_10952);
nand U11063 (N_11063,N_10941,N_10970);
xor U11064 (N_11064,N_10947,N_10858);
and U11065 (N_11065,N_10985,N_10917);
nand U11066 (N_11066,N_10888,N_10876);
nand U11067 (N_11067,N_10841,N_10861);
and U11068 (N_11068,N_10826,N_10842);
nor U11069 (N_11069,N_10820,N_10961);
nor U11070 (N_11070,N_10836,N_10847);
nor U11071 (N_11071,N_10896,N_10808);
nand U11072 (N_11072,N_10928,N_10945);
nor U11073 (N_11073,N_10984,N_10910);
or U11074 (N_11074,N_10851,N_10860);
and U11075 (N_11075,N_10828,N_10892);
or U11076 (N_11076,N_10809,N_10942);
and U11077 (N_11077,N_10819,N_10922);
nor U11078 (N_11078,N_10830,N_10805);
or U11079 (N_11079,N_10850,N_10980);
nor U11080 (N_11080,N_10871,N_10924);
nor U11081 (N_11081,N_10845,N_10988);
or U11082 (N_11082,N_10862,N_10816);
and U11083 (N_11083,N_10890,N_10954);
nor U11084 (N_11084,N_10846,N_10898);
nor U11085 (N_11085,N_10827,N_10971);
xor U11086 (N_11086,N_10867,N_10948);
or U11087 (N_11087,N_10934,N_10916);
xnor U11088 (N_11088,N_10975,N_10901);
nor U11089 (N_11089,N_10930,N_10967);
nand U11090 (N_11090,N_10931,N_10852);
nand U11091 (N_11091,N_10932,N_10832);
nor U11092 (N_11092,N_10943,N_10926);
and U11093 (N_11093,N_10814,N_10915);
nand U11094 (N_11094,N_10911,N_10923);
nor U11095 (N_11095,N_10893,N_10962);
and U11096 (N_11096,N_10944,N_10897);
or U11097 (N_11097,N_10870,N_10940);
and U11098 (N_11098,N_10904,N_10889);
nor U11099 (N_11099,N_10953,N_10833);
nor U11100 (N_11100,N_10824,N_10990);
or U11101 (N_11101,N_10996,N_10805);
or U11102 (N_11102,N_10960,N_10854);
or U11103 (N_11103,N_10867,N_10919);
nand U11104 (N_11104,N_10916,N_10864);
nand U11105 (N_11105,N_10966,N_10908);
nand U11106 (N_11106,N_10887,N_10881);
or U11107 (N_11107,N_10941,N_10902);
xor U11108 (N_11108,N_10936,N_10905);
nor U11109 (N_11109,N_10990,N_10830);
xor U11110 (N_11110,N_10843,N_10975);
nand U11111 (N_11111,N_10967,N_10932);
nand U11112 (N_11112,N_10869,N_10913);
nor U11113 (N_11113,N_10916,N_10800);
or U11114 (N_11114,N_10949,N_10902);
nand U11115 (N_11115,N_10993,N_10920);
or U11116 (N_11116,N_10881,N_10879);
nand U11117 (N_11117,N_10809,N_10882);
and U11118 (N_11118,N_10894,N_10892);
nand U11119 (N_11119,N_10825,N_10855);
nor U11120 (N_11120,N_10809,N_10908);
nor U11121 (N_11121,N_10958,N_10967);
or U11122 (N_11122,N_10904,N_10946);
xor U11123 (N_11123,N_10938,N_10925);
xnor U11124 (N_11124,N_10825,N_10851);
nor U11125 (N_11125,N_10802,N_10870);
nor U11126 (N_11126,N_10822,N_10834);
and U11127 (N_11127,N_10805,N_10869);
nor U11128 (N_11128,N_10804,N_10848);
and U11129 (N_11129,N_10890,N_10903);
nor U11130 (N_11130,N_10810,N_10911);
and U11131 (N_11131,N_10844,N_10948);
nand U11132 (N_11132,N_10893,N_10819);
or U11133 (N_11133,N_10808,N_10994);
xor U11134 (N_11134,N_10958,N_10943);
and U11135 (N_11135,N_10839,N_10995);
and U11136 (N_11136,N_10914,N_10871);
nor U11137 (N_11137,N_10959,N_10853);
nand U11138 (N_11138,N_10832,N_10853);
nor U11139 (N_11139,N_10852,N_10994);
and U11140 (N_11140,N_10835,N_10991);
nor U11141 (N_11141,N_10878,N_10887);
nor U11142 (N_11142,N_10950,N_10834);
and U11143 (N_11143,N_10820,N_10898);
nand U11144 (N_11144,N_10874,N_10993);
nand U11145 (N_11145,N_10916,N_10914);
nor U11146 (N_11146,N_10926,N_10996);
xnor U11147 (N_11147,N_10834,N_10939);
nor U11148 (N_11148,N_10844,N_10904);
and U11149 (N_11149,N_10957,N_10935);
or U11150 (N_11150,N_10978,N_10883);
nor U11151 (N_11151,N_10913,N_10851);
and U11152 (N_11152,N_10815,N_10883);
nand U11153 (N_11153,N_10802,N_10860);
and U11154 (N_11154,N_10932,N_10920);
and U11155 (N_11155,N_10938,N_10899);
nor U11156 (N_11156,N_10940,N_10828);
nand U11157 (N_11157,N_10863,N_10881);
nor U11158 (N_11158,N_10867,N_10841);
or U11159 (N_11159,N_10838,N_10923);
nor U11160 (N_11160,N_10930,N_10903);
xnor U11161 (N_11161,N_10904,N_10879);
or U11162 (N_11162,N_10824,N_10879);
xor U11163 (N_11163,N_10969,N_10972);
nor U11164 (N_11164,N_10962,N_10923);
xnor U11165 (N_11165,N_10867,N_10977);
nor U11166 (N_11166,N_10952,N_10985);
nand U11167 (N_11167,N_10817,N_10864);
and U11168 (N_11168,N_10874,N_10953);
and U11169 (N_11169,N_10985,N_10999);
xnor U11170 (N_11170,N_10963,N_10867);
nor U11171 (N_11171,N_10995,N_10817);
nand U11172 (N_11172,N_10921,N_10882);
xnor U11173 (N_11173,N_10931,N_10884);
nand U11174 (N_11174,N_10924,N_10882);
xnor U11175 (N_11175,N_10877,N_10837);
xor U11176 (N_11176,N_10817,N_10978);
nand U11177 (N_11177,N_10858,N_10976);
nand U11178 (N_11178,N_10916,N_10919);
or U11179 (N_11179,N_10922,N_10979);
nand U11180 (N_11180,N_10872,N_10875);
and U11181 (N_11181,N_10826,N_10835);
xnor U11182 (N_11182,N_10926,N_10805);
or U11183 (N_11183,N_10838,N_10814);
nand U11184 (N_11184,N_10898,N_10953);
or U11185 (N_11185,N_10867,N_10976);
or U11186 (N_11186,N_10840,N_10964);
nand U11187 (N_11187,N_10871,N_10892);
and U11188 (N_11188,N_10839,N_10820);
nand U11189 (N_11189,N_10991,N_10932);
nand U11190 (N_11190,N_10889,N_10836);
or U11191 (N_11191,N_10976,N_10938);
xor U11192 (N_11192,N_10926,N_10993);
and U11193 (N_11193,N_10850,N_10969);
nor U11194 (N_11194,N_10853,N_10841);
nand U11195 (N_11195,N_10898,N_10848);
nor U11196 (N_11196,N_10960,N_10917);
or U11197 (N_11197,N_10832,N_10920);
nand U11198 (N_11198,N_10805,N_10999);
nor U11199 (N_11199,N_10865,N_10803);
nor U11200 (N_11200,N_11119,N_11079);
nand U11201 (N_11201,N_11137,N_11197);
nand U11202 (N_11202,N_11054,N_11061);
xnor U11203 (N_11203,N_11142,N_11006);
nor U11204 (N_11204,N_11138,N_11180);
or U11205 (N_11205,N_11120,N_11179);
nor U11206 (N_11206,N_11190,N_11086);
nand U11207 (N_11207,N_11044,N_11192);
xor U11208 (N_11208,N_11011,N_11058);
xnor U11209 (N_11209,N_11130,N_11004);
nand U11210 (N_11210,N_11195,N_11060);
or U11211 (N_11211,N_11113,N_11123);
and U11212 (N_11212,N_11152,N_11189);
nand U11213 (N_11213,N_11172,N_11104);
and U11214 (N_11214,N_11096,N_11048);
nor U11215 (N_11215,N_11045,N_11154);
nor U11216 (N_11216,N_11052,N_11077);
and U11217 (N_11217,N_11013,N_11078);
or U11218 (N_11218,N_11017,N_11056);
and U11219 (N_11219,N_11005,N_11143);
and U11220 (N_11220,N_11187,N_11173);
nand U11221 (N_11221,N_11016,N_11162);
nor U11222 (N_11222,N_11121,N_11170);
nor U11223 (N_11223,N_11183,N_11194);
and U11224 (N_11224,N_11181,N_11031);
nor U11225 (N_11225,N_11102,N_11167);
nor U11226 (N_11226,N_11027,N_11186);
or U11227 (N_11227,N_11047,N_11097);
xor U11228 (N_11228,N_11133,N_11127);
nor U11229 (N_11229,N_11026,N_11043);
and U11230 (N_11230,N_11020,N_11002);
nand U11231 (N_11231,N_11168,N_11038);
nand U11232 (N_11232,N_11111,N_11141);
and U11233 (N_11233,N_11191,N_11064);
or U11234 (N_11234,N_11080,N_11144);
and U11235 (N_11235,N_11018,N_11176);
xnor U11236 (N_11236,N_11035,N_11057);
nor U11237 (N_11237,N_11110,N_11131);
or U11238 (N_11238,N_11065,N_11073);
xnor U11239 (N_11239,N_11101,N_11160);
or U11240 (N_11240,N_11166,N_11030);
xor U11241 (N_11241,N_11075,N_11157);
or U11242 (N_11242,N_11126,N_11029);
xor U11243 (N_11243,N_11128,N_11069);
or U11244 (N_11244,N_11093,N_11023);
and U11245 (N_11245,N_11107,N_11147);
or U11246 (N_11246,N_11178,N_11037);
xnor U11247 (N_11247,N_11053,N_11024);
or U11248 (N_11248,N_11041,N_11182);
nor U11249 (N_11249,N_11169,N_11090);
nand U11250 (N_11250,N_11028,N_11034);
and U11251 (N_11251,N_11100,N_11001);
xnor U11252 (N_11252,N_11066,N_11000);
or U11253 (N_11253,N_11136,N_11049);
or U11254 (N_11254,N_11174,N_11116);
nor U11255 (N_11255,N_11055,N_11040);
and U11256 (N_11256,N_11145,N_11033);
nor U11257 (N_11257,N_11199,N_11067);
xnor U11258 (N_11258,N_11095,N_11140);
xor U11259 (N_11259,N_11087,N_11106);
and U11260 (N_11260,N_11085,N_11149);
and U11261 (N_11261,N_11171,N_11129);
xnor U11262 (N_11262,N_11159,N_11021);
xor U11263 (N_11263,N_11177,N_11135);
nand U11264 (N_11264,N_11155,N_11051);
xor U11265 (N_11265,N_11132,N_11099);
nand U11266 (N_11266,N_11070,N_11025);
nand U11267 (N_11267,N_11165,N_11124);
or U11268 (N_11268,N_11084,N_11042);
and U11269 (N_11269,N_11083,N_11059);
nand U11270 (N_11270,N_11071,N_11117);
xnor U11271 (N_11271,N_11063,N_11007);
and U11272 (N_11272,N_11146,N_11134);
xnor U11273 (N_11273,N_11003,N_11032);
nand U11274 (N_11274,N_11161,N_11118);
nor U11275 (N_11275,N_11188,N_11039);
and U11276 (N_11276,N_11009,N_11164);
and U11277 (N_11277,N_11148,N_11112);
and U11278 (N_11278,N_11156,N_11103);
nor U11279 (N_11279,N_11012,N_11050);
nand U11280 (N_11280,N_11151,N_11098);
nand U11281 (N_11281,N_11122,N_11114);
xnor U11282 (N_11282,N_11105,N_11082);
and U11283 (N_11283,N_11108,N_11185);
xnor U11284 (N_11284,N_11046,N_11081);
xor U11285 (N_11285,N_11198,N_11019);
nand U11286 (N_11286,N_11175,N_11163);
nor U11287 (N_11287,N_11139,N_11158);
nor U11288 (N_11288,N_11014,N_11153);
nand U11289 (N_11289,N_11062,N_11092);
nand U11290 (N_11290,N_11036,N_11184);
xnor U11291 (N_11291,N_11115,N_11094);
xor U11292 (N_11292,N_11150,N_11076);
nand U11293 (N_11293,N_11109,N_11196);
xnor U11294 (N_11294,N_11089,N_11125);
xnor U11295 (N_11295,N_11074,N_11010);
and U11296 (N_11296,N_11091,N_11193);
nor U11297 (N_11297,N_11068,N_11022);
nor U11298 (N_11298,N_11072,N_11015);
or U11299 (N_11299,N_11088,N_11008);
and U11300 (N_11300,N_11189,N_11126);
xor U11301 (N_11301,N_11145,N_11043);
or U11302 (N_11302,N_11086,N_11119);
xor U11303 (N_11303,N_11177,N_11178);
nor U11304 (N_11304,N_11010,N_11164);
nand U11305 (N_11305,N_11146,N_11018);
or U11306 (N_11306,N_11006,N_11189);
nor U11307 (N_11307,N_11049,N_11173);
nand U11308 (N_11308,N_11017,N_11144);
nor U11309 (N_11309,N_11119,N_11029);
nand U11310 (N_11310,N_11135,N_11046);
or U11311 (N_11311,N_11159,N_11108);
and U11312 (N_11312,N_11025,N_11177);
xor U11313 (N_11313,N_11160,N_11059);
nand U11314 (N_11314,N_11038,N_11073);
and U11315 (N_11315,N_11143,N_11042);
nand U11316 (N_11316,N_11145,N_11088);
and U11317 (N_11317,N_11064,N_11146);
nand U11318 (N_11318,N_11047,N_11131);
or U11319 (N_11319,N_11012,N_11057);
xor U11320 (N_11320,N_11174,N_11009);
nand U11321 (N_11321,N_11197,N_11104);
or U11322 (N_11322,N_11092,N_11168);
and U11323 (N_11323,N_11149,N_11059);
xnor U11324 (N_11324,N_11189,N_11195);
nand U11325 (N_11325,N_11043,N_11115);
xor U11326 (N_11326,N_11177,N_11047);
or U11327 (N_11327,N_11114,N_11037);
and U11328 (N_11328,N_11001,N_11137);
xnor U11329 (N_11329,N_11136,N_11138);
nand U11330 (N_11330,N_11149,N_11133);
or U11331 (N_11331,N_11002,N_11072);
or U11332 (N_11332,N_11109,N_11067);
or U11333 (N_11333,N_11109,N_11144);
and U11334 (N_11334,N_11032,N_11103);
or U11335 (N_11335,N_11074,N_11075);
xnor U11336 (N_11336,N_11187,N_11030);
nor U11337 (N_11337,N_11019,N_11075);
or U11338 (N_11338,N_11148,N_11062);
xor U11339 (N_11339,N_11111,N_11135);
nor U11340 (N_11340,N_11169,N_11118);
xor U11341 (N_11341,N_11009,N_11077);
nand U11342 (N_11342,N_11122,N_11165);
and U11343 (N_11343,N_11087,N_11167);
and U11344 (N_11344,N_11066,N_11113);
nand U11345 (N_11345,N_11176,N_11142);
xor U11346 (N_11346,N_11170,N_11007);
xnor U11347 (N_11347,N_11086,N_11114);
xnor U11348 (N_11348,N_11174,N_11168);
or U11349 (N_11349,N_11087,N_11001);
nand U11350 (N_11350,N_11138,N_11110);
xor U11351 (N_11351,N_11089,N_11065);
xor U11352 (N_11352,N_11027,N_11167);
nor U11353 (N_11353,N_11177,N_11038);
nand U11354 (N_11354,N_11171,N_11079);
or U11355 (N_11355,N_11086,N_11009);
nor U11356 (N_11356,N_11039,N_11165);
and U11357 (N_11357,N_11144,N_11062);
and U11358 (N_11358,N_11069,N_11041);
xor U11359 (N_11359,N_11151,N_11142);
and U11360 (N_11360,N_11117,N_11061);
xor U11361 (N_11361,N_11117,N_11144);
or U11362 (N_11362,N_11194,N_11155);
nor U11363 (N_11363,N_11050,N_11194);
nor U11364 (N_11364,N_11174,N_11028);
nor U11365 (N_11365,N_11183,N_11004);
or U11366 (N_11366,N_11106,N_11047);
nand U11367 (N_11367,N_11058,N_11043);
and U11368 (N_11368,N_11012,N_11054);
or U11369 (N_11369,N_11057,N_11193);
nor U11370 (N_11370,N_11021,N_11073);
and U11371 (N_11371,N_11174,N_11179);
or U11372 (N_11372,N_11015,N_11036);
or U11373 (N_11373,N_11066,N_11179);
nor U11374 (N_11374,N_11059,N_11179);
or U11375 (N_11375,N_11051,N_11139);
and U11376 (N_11376,N_11072,N_11020);
nand U11377 (N_11377,N_11095,N_11013);
or U11378 (N_11378,N_11058,N_11187);
nand U11379 (N_11379,N_11083,N_11139);
nor U11380 (N_11380,N_11158,N_11176);
or U11381 (N_11381,N_11109,N_11173);
xnor U11382 (N_11382,N_11066,N_11174);
and U11383 (N_11383,N_11190,N_11033);
or U11384 (N_11384,N_11016,N_11072);
nand U11385 (N_11385,N_11080,N_11012);
and U11386 (N_11386,N_11146,N_11154);
or U11387 (N_11387,N_11084,N_11060);
nor U11388 (N_11388,N_11062,N_11125);
or U11389 (N_11389,N_11135,N_11125);
and U11390 (N_11390,N_11004,N_11052);
nor U11391 (N_11391,N_11101,N_11173);
nand U11392 (N_11392,N_11117,N_11121);
or U11393 (N_11393,N_11187,N_11071);
or U11394 (N_11394,N_11093,N_11081);
xnor U11395 (N_11395,N_11109,N_11141);
and U11396 (N_11396,N_11167,N_11028);
nor U11397 (N_11397,N_11030,N_11075);
and U11398 (N_11398,N_11197,N_11025);
or U11399 (N_11399,N_11096,N_11126);
nor U11400 (N_11400,N_11224,N_11262);
and U11401 (N_11401,N_11371,N_11299);
nor U11402 (N_11402,N_11390,N_11227);
xnor U11403 (N_11403,N_11347,N_11304);
or U11404 (N_11404,N_11216,N_11375);
or U11405 (N_11405,N_11367,N_11248);
or U11406 (N_11406,N_11255,N_11240);
nor U11407 (N_11407,N_11238,N_11206);
and U11408 (N_11408,N_11338,N_11201);
or U11409 (N_11409,N_11277,N_11320);
nand U11410 (N_11410,N_11392,N_11245);
xor U11411 (N_11411,N_11391,N_11334);
nand U11412 (N_11412,N_11272,N_11373);
or U11413 (N_11413,N_11268,N_11399);
nor U11414 (N_11414,N_11340,N_11329);
nand U11415 (N_11415,N_11203,N_11280);
and U11416 (N_11416,N_11351,N_11247);
and U11417 (N_11417,N_11376,N_11353);
nand U11418 (N_11418,N_11349,N_11225);
or U11419 (N_11419,N_11208,N_11316);
xor U11420 (N_11420,N_11327,N_11237);
xor U11421 (N_11421,N_11275,N_11253);
and U11422 (N_11422,N_11374,N_11305);
nand U11423 (N_11423,N_11241,N_11362);
xor U11424 (N_11424,N_11310,N_11243);
xor U11425 (N_11425,N_11239,N_11257);
nand U11426 (N_11426,N_11372,N_11378);
xor U11427 (N_11427,N_11383,N_11330);
or U11428 (N_11428,N_11267,N_11301);
nand U11429 (N_11429,N_11321,N_11252);
nor U11430 (N_11430,N_11302,N_11274);
nand U11431 (N_11431,N_11346,N_11235);
or U11432 (N_11432,N_11335,N_11395);
nor U11433 (N_11433,N_11264,N_11314);
nand U11434 (N_11434,N_11328,N_11290);
and U11435 (N_11435,N_11251,N_11219);
and U11436 (N_11436,N_11270,N_11218);
and U11437 (N_11437,N_11344,N_11356);
or U11438 (N_11438,N_11322,N_11229);
or U11439 (N_11439,N_11387,N_11363);
xor U11440 (N_11440,N_11369,N_11209);
or U11441 (N_11441,N_11359,N_11307);
nor U11442 (N_11442,N_11331,N_11318);
or U11443 (N_11443,N_11337,N_11360);
nor U11444 (N_11444,N_11273,N_11271);
nor U11445 (N_11445,N_11233,N_11386);
xnor U11446 (N_11446,N_11396,N_11249);
nor U11447 (N_11447,N_11308,N_11291);
or U11448 (N_11448,N_11244,N_11293);
or U11449 (N_11449,N_11236,N_11295);
or U11450 (N_11450,N_11370,N_11232);
and U11451 (N_11451,N_11341,N_11368);
or U11452 (N_11452,N_11254,N_11300);
nand U11453 (N_11453,N_11296,N_11297);
xor U11454 (N_11454,N_11250,N_11364);
and U11455 (N_11455,N_11246,N_11213);
nor U11456 (N_11456,N_11382,N_11388);
xnor U11457 (N_11457,N_11377,N_11207);
nand U11458 (N_11458,N_11398,N_11289);
nor U11459 (N_11459,N_11343,N_11294);
xor U11460 (N_11460,N_11352,N_11228);
xor U11461 (N_11461,N_11278,N_11279);
xor U11462 (N_11462,N_11269,N_11357);
xor U11463 (N_11463,N_11220,N_11205);
nor U11464 (N_11464,N_11265,N_11309);
nor U11465 (N_11465,N_11266,N_11214);
xor U11466 (N_11466,N_11223,N_11389);
and U11467 (N_11467,N_11355,N_11324);
or U11468 (N_11468,N_11215,N_11380);
nor U11469 (N_11469,N_11221,N_11306);
and U11470 (N_11470,N_11385,N_11282);
or U11471 (N_11471,N_11261,N_11312);
nor U11472 (N_11472,N_11281,N_11339);
xor U11473 (N_11473,N_11298,N_11394);
nor U11474 (N_11474,N_11287,N_11292);
xnor U11475 (N_11475,N_11345,N_11354);
nand U11476 (N_11476,N_11258,N_11283);
and U11477 (N_11477,N_11212,N_11332);
xor U11478 (N_11478,N_11222,N_11397);
nor U11479 (N_11479,N_11285,N_11313);
or U11480 (N_11480,N_11204,N_11234);
nor U11481 (N_11481,N_11384,N_11200);
nand U11482 (N_11482,N_11226,N_11288);
or U11483 (N_11483,N_11230,N_11323);
or U11484 (N_11484,N_11348,N_11210);
and U11485 (N_11485,N_11211,N_11315);
and U11486 (N_11486,N_11381,N_11263);
nor U11487 (N_11487,N_11217,N_11365);
nand U11488 (N_11488,N_11202,N_11242);
nand U11489 (N_11489,N_11336,N_11311);
nand U11490 (N_11490,N_11319,N_11333);
and U11491 (N_11491,N_11379,N_11350);
and U11492 (N_11492,N_11358,N_11366);
xor U11493 (N_11493,N_11393,N_11284);
xor U11494 (N_11494,N_11303,N_11326);
and U11495 (N_11495,N_11231,N_11260);
nor U11496 (N_11496,N_11361,N_11317);
or U11497 (N_11497,N_11256,N_11259);
and U11498 (N_11498,N_11276,N_11342);
xnor U11499 (N_11499,N_11286,N_11325);
xor U11500 (N_11500,N_11307,N_11266);
and U11501 (N_11501,N_11257,N_11235);
xor U11502 (N_11502,N_11217,N_11262);
nor U11503 (N_11503,N_11234,N_11324);
xor U11504 (N_11504,N_11388,N_11227);
nand U11505 (N_11505,N_11202,N_11347);
nand U11506 (N_11506,N_11270,N_11265);
xor U11507 (N_11507,N_11293,N_11235);
nand U11508 (N_11508,N_11262,N_11249);
or U11509 (N_11509,N_11374,N_11254);
and U11510 (N_11510,N_11360,N_11244);
or U11511 (N_11511,N_11384,N_11227);
xor U11512 (N_11512,N_11310,N_11369);
xor U11513 (N_11513,N_11236,N_11324);
or U11514 (N_11514,N_11332,N_11220);
nor U11515 (N_11515,N_11388,N_11333);
nand U11516 (N_11516,N_11356,N_11202);
xor U11517 (N_11517,N_11322,N_11366);
and U11518 (N_11518,N_11301,N_11270);
or U11519 (N_11519,N_11395,N_11243);
and U11520 (N_11520,N_11282,N_11331);
or U11521 (N_11521,N_11346,N_11201);
nand U11522 (N_11522,N_11297,N_11236);
nand U11523 (N_11523,N_11324,N_11360);
and U11524 (N_11524,N_11319,N_11399);
and U11525 (N_11525,N_11238,N_11334);
and U11526 (N_11526,N_11269,N_11292);
xor U11527 (N_11527,N_11251,N_11248);
nor U11528 (N_11528,N_11271,N_11384);
and U11529 (N_11529,N_11291,N_11389);
xor U11530 (N_11530,N_11238,N_11229);
or U11531 (N_11531,N_11246,N_11227);
nand U11532 (N_11532,N_11265,N_11392);
nor U11533 (N_11533,N_11261,N_11354);
and U11534 (N_11534,N_11396,N_11298);
and U11535 (N_11535,N_11296,N_11274);
or U11536 (N_11536,N_11231,N_11273);
or U11537 (N_11537,N_11221,N_11234);
xor U11538 (N_11538,N_11215,N_11356);
nand U11539 (N_11539,N_11266,N_11249);
or U11540 (N_11540,N_11355,N_11248);
and U11541 (N_11541,N_11232,N_11346);
or U11542 (N_11542,N_11203,N_11369);
xor U11543 (N_11543,N_11367,N_11259);
or U11544 (N_11544,N_11254,N_11252);
nor U11545 (N_11545,N_11231,N_11358);
or U11546 (N_11546,N_11253,N_11306);
nor U11547 (N_11547,N_11398,N_11288);
nor U11548 (N_11548,N_11285,N_11332);
nor U11549 (N_11549,N_11368,N_11325);
and U11550 (N_11550,N_11256,N_11204);
or U11551 (N_11551,N_11341,N_11382);
and U11552 (N_11552,N_11262,N_11239);
xnor U11553 (N_11553,N_11278,N_11223);
nor U11554 (N_11554,N_11364,N_11248);
nor U11555 (N_11555,N_11387,N_11380);
nand U11556 (N_11556,N_11310,N_11348);
and U11557 (N_11557,N_11390,N_11359);
nor U11558 (N_11558,N_11244,N_11335);
and U11559 (N_11559,N_11274,N_11341);
or U11560 (N_11560,N_11250,N_11288);
and U11561 (N_11561,N_11207,N_11225);
nand U11562 (N_11562,N_11389,N_11237);
xnor U11563 (N_11563,N_11276,N_11231);
nand U11564 (N_11564,N_11231,N_11376);
nand U11565 (N_11565,N_11395,N_11262);
nand U11566 (N_11566,N_11353,N_11368);
nand U11567 (N_11567,N_11279,N_11329);
nand U11568 (N_11568,N_11398,N_11322);
and U11569 (N_11569,N_11274,N_11371);
and U11570 (N_11570,N_11324,N_11245);
nor U11571 (N_11571,N_11358,N_11337);
or U11572 (N_11572,N_11326,N_11327);
and U11573 (N_11573,N_11298,N_11363);
xor U11574 (N_11574,N_11307,N_11387);
nand U11575 (N_11575,N_11370,N_11283);
nand U11576 (N_11576,N_11319,N_11378);
and U11577 (N_11577,N_11207,N_11235);
xnor U11578 (N_11578,N_11313,N_11342);
or U11579 (N_11579,N_11285,N_11239);
and U11580 (N_11580,N_11213,N_11327);
nor U11581 (N_11581,N_11267,N_11316);
nor U11582 (N_11582,N_11301,N_11215);
nand U11583 (N_11583,N_11243,N_11397);
nor U11584 (N_11584,N_11390,N_11329);
xnor U11585 (N_11585,N_11386,N_11330);
xnor U11586 (N_11586,N_11305,N_11301);
xnor U11587 (N_11587,N_11325,N_11390);
xnor U11588 (N_11588,N_11267,N_11278);
nor U11589 (N_11589,N_11398,N_11399);
or U11590 (N_11590,N_11390,N_11298);
nand U11591 (N_11591,N_11325,N_11231);
nand U11592 (N_11592,N_11346,N_11318);
nand U11593 (N_11593,N_11262,N_11294);
or U11594 (N_11594,N_11391,N_11331);
and U11595 (N_11595,N_11228,N_11246);
or U11596 (N_11596,N_11331,N_11295);
or U11597 (N_11597,N_11260,N_11297);
or U11598 (N_11598,N_11266,N_11217);
or U11599 (N_11599,N_11269,N_11391);
nor U11600 (N_11600,N_11503,N_11470);
nand U11601 (N_11601,N_11558,N_11413);
nand U11602 (N_11602,N_11482,N_11435);
and U11603 (N_11603,N_11593,N_11466);
or U11604 (N_11604,N_11425,N_11513);
or U11605 (N_11605,N_11449,N_11401);
nor U11606 (N_11606,N_11578,N_11576);
xnor U11607 (N_11607,N_11548,N_11434);
or U11608 (N_11608,N_11537,N_11440);
nor U11609 (N_11609,N_11564,N_11517);
or U11610 (N_11610,N_11584,N_11567);
xnor U11611 (N_11611,N_11444,N_11533);
xor U11612 (N_11612,N_11455,N_11439);
or U11613 (N_11613,N_11500,N_11492);
xnor U11614 (N_11614,N_11471,N_11411);
and U11615 (N_11615,N_11595,N_11546);
or U11616 (N_11616,N_11424,N_11536);
and U11617 (N_11617,N_11501,N_11510);
nand U11618 (N_11618,N_11462,N_11436);
nor U11619 (N_11619,N_11549,N_11532);
and U11620 (N_11620,N_11485,N_11502);
xnor U11621 (N_11621,N_11402,N_11465);
and U11622 (N_11622,N_11438,N_11433);
nor U11623 (N_11623,N_11540,N_11582);
xor U11624 (N_11624,N_11598,N_11423);
xor U11625 (N_11625,N_11431,N_11539);
nor U11626 (N_11626,N_11432,N_11543);
xnor U11627 (N_11627,N_11426,N_11474);
nand U11628 (N_11628,N_11562,N_11448);
xor U11629 (N_11629,N_11407,N_11568);
or U11630 (N_11630,N_11592,N_11491);
nand U11631 (N_11631,N_11530,N_11415);
or U11632 (N_11632,N_11475,N_11556);
nand U11633 (N_11633,N_11490,N_11538);
or U11634 (N_11634,N_11486,N_11515);
and U11635 (N_11635,N_11479,N_11428);
xnor U11636 (N_11636,N_11561,N_11450);
or U11637 (N_11637,N_11585,N_11419);
nor U11638 (N_11638,N_11569,N_11454);
nor U11639 (N_11639,N_11406,N_11520);
or U11640 (N_11640,N_11575,N_11463);
or U11641 (N_11641,N_11544,N_11400);
and U11642 (N_11642,N_11487,N_11464);
and U11643 (N_11643,N_11557,N_11480);
and U11644 (N_11644,N_11506,N_11405);
xnor U11645 (N_11645,N_11408,N_11523);
nand U11646 (N_11646,N_11551,N_11467);
nand U11647 (N_11647,N_11511,N_11519);
or U11648 (N_11648,N_11553,N_11514);
nand U11649 (N_11649,N_11473,N_11573);
nand U11650 (N_11650,N_11458,N_11550);
xor U11651 (N_11651,N_11498,N_11521);
nand U11652 (N_11652,N_11484,N_11478);
xnor U11653 (N_11653,N_11403,N_11504);
and U11654 (N_11654,N_11468,N_11518);
or U11655 (N_11655,N_11497,N_11509);
xnor U11656 (N_11656,N_11421,N_11446);
nor U11657 (N_11657,N_11531,N_11429);
and U11658 (N_11658,N_11545,N_11445);
and U11659 (N_11659,N_11404,N_11591);
nor U11660 (N_11660,N_11499,N_11451);
nor U11661 (N_11661,N_11422,N_11427);
xnor U11662 (N_11662,N_11589,N_11507);
xnor U11663 (N_11663,N_11547,N_11508);
xnor U11664 (N_11664,N_11409,N_11457);
nand U11665 (N_11665,N_11541,N_11418);
nor U11666 (N_11666,N_11442,N_11460);
xnor U11667 (N_11667,N_11472,N_11443);
nor U11668 (N_11668,N_11489,N_11483);
nand U11669 (N_11669,N_11441,N_11493);
nand U11670 (N_11670,N_11453,N_11412);
nand U11671 (N_11671,N_11488,N_11528);
and U11672 (N_11672,N_11525,N_11452);
or U11673 (N_11673,N_11566,N_11577);
nand U11674 (N_11674,N_11524,N_11459);
or U11675 (N_11675,N_11430,N_11586);
nor U11676 (N_11676,N_11416,N_11522);
xnor U11677 (N_11677,N_11420,N_11588);
nand U11678 (N_11678,N_11481,N_11552);
and U11679 (N_11679,N_11565,N_11599);
nand U11680 (N_11680,N_11560,N_11596);
nand U11681 (N_11681,N_11559,N_11594);
nor U11682 (N_11682,N_11417,N_11461);
nand U11683 (N_11683,N_11495,N_11414);
or U11684 (N_11684,N_11456,N_11571);
xnor U11685 (N_11685,N_11535,N_11527);
nor U11686 (N_11686,N_11554,N_11526);
nand U11687 (N_11687,N_11581,N_11555);
and U11688 (N_11688,N_11590,N_11580);
or U11689 (N_11689,N_11587,N_11447);
nor U11690 (N_11690,N_11529,N_11494);
or U11691 (N_11691,N_11505,N_11572);
nor U11692 (N_11692,N_11583,N_11410);
or U11693 (N_11693,N_11437,N_11512);
and U11694 (N_11694,N_11574,N_11563);
nand U11695 (N_11695,N_11496,N_11542);
nand U11696 (N_11696,N_11469,N_11570);
nand U11697 (N_11697,N_11579,N_11476);
xor U11698 (N_11698,N_11534,N_11597);
nor U11699 (N_11699,N_11516,N_11477);
xor U11700 (N_11700,N_11423,N_11485);
nor U11701 (N_11701,N_11474,N_11491);
xnor U11702 (N_11702,N_11597,N_11448);
nor U11703 (N_11703,N_11405,N_11497);
xnor U11704 (N_11704,N_11420,N_11511);
and U11705 (N_11705,N_11465,N_11493);
or U11706 (N_11706,N_11515,N_11458);
xnor U11707 (N_11707,N_11400,N_11553);
xnor U11708 (N_11708,N_11487,N_11581);
xnor U11709 (N_11709,N_11518,N_11422);
or U11710 (N_11710,N_11565,N_11419);
xor U11711 (N_11711,N_11560,N_11425);
and U11712 (N_11712,N_11538,N_11485);
and U11713 (N_11713,N_11555,N_11549);
nor U11714 (N_11714,N_11552,N_11444);
xnor U11715 (N_11715,N_11440,N_11590);
nor U11716 (N_11716,N_11465,N_11401);
and U11717 (N_11717,N_11537,N_11508);
nor U11718 (N_11718,N_11537,N_11434);
and U11719 (N_11719,N_11564,N_11490);
nand U11720 (N_11720,N_11491,N_11494);
and U11721 (N_11721,N_11466,N_11436);
nor U11722 (N_11722,N_11503,N_11480);
and U11723 (N_11723,N_11439,N_11492);
or U11724 (N_11724,N_11542,N_11495);
nand U11725 (N_11725,N_11596,N_11485);
nor U11726 (N_11726,N_11554,N_11517);
xnor U11727 (N_11727,N_11459,N_11504);
xor U11728 (N_11728,N_11457,N_11557);
and U11729 (N_11729,N_11407,N_11442);
and U11730 (N_11730,N_11527,N_11420);
xor U11731 (N_11731,N_11554,N_11464);
and U11732 (N_11732,N_11596,N_11549);
nand U11733 (N_11733,N_11489,N_11585);
or U11734 (N_11734,N_11566,N_11573);
nor U11735 (N_11735,N_11470,N_11484);
nor U11736 (N_11736,N_11482,N_11494);
xor U11737 (N_11737,N_11423,N_11441);
or U11738 (N_11738,N_11401,N_11587);
nand U11739 (N_11739,N_11496,N_11528);
nand U11740 (N_11740,N_11572,N_11583);
and U11741 (N_11741,N_11416,N_11404);
or U11742 (N_11742,N_11467,N_11406);
and U11743 (N_11743,N_11583,N_11597);
or U11744 (N_11744,N_11496,N_11569);
xnor U11745 (N_11745,N_11507,N_11491);
nor U11746 (N_11746,N_11408,N_11445);
xnor U11747 (N_11747,N_11451,N_11430);
xor U11748 (N_11748,N_11406,N_11474);
xnor U11749 (N_11749,N_11408,N_11491);
xor U11750 (N_11750,N_11465,N_11495);
and U11751 (N_11751,N_11497,N_11575);
xor U11752 (N_11752,N_11420,N_11478);
nor U11753 (N_11753,N_11498,N_11501);
or U11754 (N_11754,N_11530,N_11591);
xnor U11755 (N_11755,N_11547,N_11474);
xnor U11756 (N_11756,N_11505,N_11592);
or U11757 (N_11757,N_11537,N_11560);
and U11758 (N_11758,N_11505,N_11480);
nand U11759 (N_11759,N_11587,N_11584);
nand U11760 (N_11760,N_11419,N_11457);
xor U11761 (N_11761,N_11561,N_11411);
and U11762 (N_11762,N_11474,N_11427);
or U11763 (N_11763,N_11585,N_11447);
or U11764 (N_11764,N_11563,N_11426);
or U11765 (N_11765,N_11561,N_11503);
nand U11766 (N_11766,N_11480,N_11485);
nand U11767 (N_11767,N_11478,N_11532);
or U11768 (N_11768,N_11484,N_11577);
nor U11769 (N_11769,N_11418,N_11447);
or U11770 (N_11770,N_11545,N_11536);
and U11771 (N_11771,N_11579,N_11562);
or U11772 (N_11772,N_11463,N_11477);
or U11773 (N_11773,N_11490,N_11588);
or U11774 (N_11774,N_11483,N_11576);
and U11775 (N_11775,N_11553,N_11567);
nor U11776 (N_11776,N_11568,N_11406);
xnor U11777 (N_11777,N_11526,N_11438);
xnor U11778 (N_11778,N_11501,N_11529);
or U11779 (N_11779,N_11534,N_11543);
nand U11780 (N_11780,N_11568,N_11543);
nand U11781 (N_11781,N_11573,N_11463);
nand U11782 (N_11782,N_11441,N_11444);
xnor U11783 (N_11783,N_11553,N_11413);
xnor U11784 (N_11784,N_11568,N_11437);
nand U11785 (N_11785,N_11482,N_11571);
and U11786 (N_11786,N_11519,N_11523);
xnor U11787 (N_11787,N_11479,N_11562);
nor U11788 (N_11788,N_11505,N_11529);
nand U11789 (N_11789,N_11511,N_11542);
and U11790 (N_11790,N_11595,N_11531);
or U11791 (N_11791,N_11467,N_11522);
or U11792 (N_11792,N_11524,N_11411);
or U11793 (N_11793,N_11509,N_11434);
nand U11794 (N_11794,N_11404,N_11502);
nand U11795 (N_11795,N_11585,N_11471);
and U11796 (N_11796,N_11504,N_11587);
nor U11797 (N_11797,N_11463,N_11441);
xnor U11798 (N_11798,N_11402,N_11538);
xnor U11799 (N_11799,N_11596,N_11569);
and U11800 (N_11800,N_11767,N_11631);
nor U11801 (N_11801,N_11740,N_11612);
or U11802 (N_11802,N_11755,N_11735);
xnor U11803 (N_11803,N_11791,N_11657);
nand U11804 (N_11804,N_11701,N_11643);
and U11805 (N_11805,N_11748,N_11694);
nor U11806 (N_11806,N_11655,N_11733);
nor U11807 (N_11807,N_11609,N_11670);
and U11808 (N_11808,N_11610,N_11667);
and U11809 (N_11809,N_11703,N_11676);
or U11810 (N_11810,N_11615,N_11659);
or U11811 (N_11811,N_11674,N_11605);
or U11812 (N_11812,N_11663,N_11705);
nand U11813 (N_11813,N_11603,N_11601);
nand U11814 (N_11814,N_11710,N_11725);
nand U11815 (N_11815,N_11649,N_11633);
and U11816 (N_11816,N_11696,N_11709);
nor U11817 (N_11817,N_11744,N_11789);
or U11818 (N_11818,N_11766,N_11666);
or U11819 (N_11819,N_11621,N_11752);
and U11820 (N_11820,N_11677,N_11765);
nor U11821 (N_11821,N_11698,N_11626);
nand U11822 (N_11822,N_11632,N_11792);
xnor U11823 (N_11823,N_11793,N_11680);
and U11824 (N_11824,N_11684,N_11736);
and U11825 (N_11825,N_11624,N_11784);
or U11826 (N_11826,N_11687,N_11719);
and U11827 (N_11827,N_11679,N_11753);
nor U11828 (N_11828,N_11742,N_11786);
and U11829 (N_11829,N_11781,N_11754);
xor U11830 (N_11830,N_11718,N_11652);
nand U11831 (N_11831,N_11737,N_11651);
nand U11832 (N_11832,N_11650,N_11717);
or U11833 (N_11833,N_11797,N_11660);
and U11834 (N_11834,N_11714,N_11762);
nor U11835 (N_11835,N_11611,N_11732);
or U11836 (N_11836,N_11630,N_11770);
nand U11837 (N_11837,N_11727,N_11749);
or U11838 (N_11838,N_11706,N_11665);
nand U11839 (N_11839,N_11618,N_11774);
nor U11840 (N_11840,N_11600,N_11691);
xnor U11841 (N_11841,N_11757,N_11734);
and U11842 (N_11842,N_11614,N_11640);
and U11843 (N_11843,N_11627,N_11654);
nor U11844 (N_11844,N_11722,N_11639);
xor U11845 (N_11845,N_11697,N_11606);
nor U11846 (N_11846,N_11708,N_11695);
xor U11847 (N_11847,N_11712,N_11799);
or U11848 (N_11848,N_11685,N_11661);
or U11849 (N_11849,N_11634,N_11636);
nand U11850 (N_11850,N_11700,N_11794);
or U11851 (N_11851,N_11731,N_11750);
or U11852 (N_11852,N_11681,N_11656);
or U11853 (N_11853,N_11760,N_11769);
xnor U11854 (N_11854,N_11662,N_11798);
xnor U11855 (N_11855,N_11646,N_11642);
nand U11856 (N_11856,N_11692,N_11778);
nor U11857 (N_11857,N_11653,N_11773);
and U11858 (N_11858,N_11777,N_11788);
xnor U11859 (N_11859,N_11625,N_11716);
xor U11860 (N_11860,N_11720,N_11616);
nand U11861 (N_11861,N_11673,N_11604);
xnor U11862 (N_11862,N_11613,N_11723);
nand U11863 (N_11863,N_11739,N_11758);
or U11864 (N_11864,N_11738,N_11768);
nand U11865 (N_11865,N_11678,N_11729);
nor U11866 (N_11866,N_11771,N_11782);
or U11867 (N_11867,N_11775,N_11751);
nand U11868 (N_11868,N_11726,N_11672);
nand U11869 (N_11869,N_11629,N_11772);
and U11870 (N_11870,N_11713,N_11686);
nand U11871 (N_11871,N_11658,N_11635);
or U11872 (N_11872,N_11780,N_11707);
nand U11873 (N_11873,N_11641,N_11617);
xor U11874 (N_11874,N_11724,N_11647);
nor U11875 (N_11875,N_11623,N_11747);
and U11876 (N_11876,N_11730,N_11648);
xor U11877 (N_11877,N_11622,N_11787);
nor U11878 (N_11878,N_11759,N_11699);
xor U11879 (N_11879,N_11702,N_11728);
and U11880 (N_11880,N_11675,N_11608);
nand U11881 (N_11881,N_11790,N_11682);
xnor U11882 (N_11882,N_11721,N_11620);
nor U11883 (N_11883,N_11756,N_11602);
xor U11884 (N_11884,N_11628,N_11764);
nand U11885 (N_11885,N_11671,N_11743);
and U11886 (N_11886,N_11795,N_11779);
nor U11887 (N_11887,N_11669,N_11637);
xnor U11888 (N_11888,N_11607,N_11796);
and U11889 (N_11889,N_11683,N_11783);
nor U11890 (N_11890,N_11776,N_11704);
or U11891 (N_11891,N_11715,N_11644);
nor U11892 (N_11892,N_11688,N_11746);
nor U11893 (N_11893,N_11711,N_11664);
and U11894 (N_11894,N_11693,N_11638);
or U11895 (N_11895,N_11668,N_11785);
nor U11896 (N_11896,N_11690,N_11761);
and U11897 (N_11897,N_11741,N_11689);
nor U11898 (N_11898,N_11745,N_11619);
or U11899 (N_11899,N_11645,N_11763);
nand U11900 (N_11900,N_11681,N_11663);
or U11901 (N_11901,N_11632,N_11605);
nor U11902 (N_11902,N_11680,N_11711);
and U11903 (N_11903,N_11664,N_11659);
nand U11904 (N_11904,N_11694,N_11690);
xor U11905 (N_11905,N_11710,N_11744);
nand U11906 (N_11906,N_11752,N_11628);
nor U11907 (N_11907,N_11700,N_11637);
nand U11908 (N_11908,N_11698,N_11674);
nor U11909 (N_11909,N_11619,N_11603);
or U11910 (N_11910,N_11794,N_11696);
and U11911 (N_11911,N_11751,N_11682);
or U11912 (N_11912,N_11784,N_11750);
nand U11913 (N_11913,N_11760,N_11695);
nand U11914 (N_11914,N_11772,N_11620);
and U11915 (N_11915,N_11673,N_11711);
nor U11916 (N_11916,N_11701,N_11648);
or U11917 (N_11917,N_11674,N_11782);
nor U11918 (N_11918,N_11725,N_11647);
nor U11919 (N_11919,N_11698,N_11785);
and U11920 (N_11920,N_11611,N_11659);
nand U11921 (N_11921,N_11654,N_11745);
and U11922 (N_11922,N_11622,N_11643);
or U11923 (N_11923,N_11645,N_11635);
nand U11924 (N_11924,N_11672,N_11639);
xnor U11925 (N_11925,N_11781,N_11750);
nand U11926 (N_11926,N_11790,N_11660);
nor U11927 (N_11927,N_11638,N_11773);
nand U11928 (N_11928,N_11765,N_11641);
nor U11929 (N_11929,N_11777,N_11789);
nor U11930 (N_11930,N_11602,N_11709);
nand U11931 (N_11931,N_11780,N_11752);
xnor U11932 (N_11932,N_11780,N_11798);
nand U11933 (N_11933,N_11704,N_11728);
xnor U11934 (N_11934,N_11689,N_11715);
nor U11935 (N_11935,N_11636,N_11639);
nand U11936 (N_11936,N_11615,N_11689);
and U11937 (N_11937,N_11697,N_11609);
and U11938 (N_11938,N_11793,N_11639);
or U11939 (N_11939,N_11795,N_11636);
xnor U11940 (N_11940,N_11731,N_11758);
nor U11941 (N_11941,N_11623,N_11727);
nor U11942 (N_11942,N_11798,N_11609);
nand U11943 (N_11943,N_11645,N_11784);
xnor U11944 (N_11944,N_11738,N_11754);
and U11945 (N_11945,N_11758,N_11716);
xnor U11946 (N_11946,N_11773,N_11705);
xnor U11947 (N_11947,N_11763,N_11742);
nand U11948 (N_11948,N_11604,N_11626);
or U11949 (N_11949,N_11653,N_11779);
or U11950 (N_11950,N_11688,N_11733);
or U11951 (N_11951,N_11606,N_11751);
nor U11952 (N_11952,N_11791,N_11719);
nand U11953 (N_11953,N_11632,N_11601);
xor U11954 (N_11954,N_11635,N_11694);
or U11955 (N_11955,N_11723,N_11640);
xnor U11956 (N_11956,N_11648,N_11683);
nor U11957 (N_11957,N_11740,N_11714);
nand U11958 (N_11958,N_11636,N_11729);
and U11959 (N_11959,N_11705,N_11682);
nand U11960 (N_11960,N_11780,N_11759);
xor U11961 (N_11961,N_11774,N_11666);
nor U11962 (N_11962,N_11739,N_11707);
or U11963 (N_11963,N_11752,N_11661);
and U11964 (N_11964,N_11685,N_11679);
and U11965 (N_11965,N_11670,N_11623);
or U11966 (N_11966,N_11673,N_11671);
and U11967 (N_11967,N_11724,N_11723);
nor U11968 (N_11968,N_11799,N_11675);
nand U11969 (N_11969,N_11793,N_11695);
xnor U11970 (N_11970,N_11741,N_11603);
and U11971 (N_11971,N_11750,N_11719);
or U11972 (N_11972,N_11780,N_11790);
xor U11973 (N_11973,N_11601,N_11657);
xnor U11974 (N_11974,N_11625,N_11699);
nor U11975 (N_11975,N_11786,N_11642);
nand U11976 (N_11976,N_11627,N_11774);
nor U11977 (N_11977,N_11765,N_11774);
or U11978 (N_11978,N_11763,N_11708);
nor U11979 (N_11979,N_11633,N_11667);
nor U11980 (N_11980,N_11663,N_11674);
and U11981 (N_11981,N_11787,N_11680);
nand U11982 (N_11982,N_11641,N_11708);
or U11983 (N_11983,N_11663,N_11678);
nor U11984 (N_11984,N_11660,N_11731);
and U11985 (N_11985,N_11708,N_11739);
nand U11986 (N_11986,N_11605,N_11649);
nor U11987 (N_11987,N_11714,N_11711);
and U11988 (N_11988,N_11603,N_11714);
nor U11989 (N_11989,N_11742,N_11605);
xor U11990 (N_11990,N_11614,N_11695);
xor U11991 (N_11991,N_11673,N_11726);
nor U11992 (N_11992,N_11758,N_11637);
and U11993 (N_11993,N_11646,N_11688);
nor U11994 (N_11994,N_11795,N_11744);
nand U11995 (N_11995,N_11671,N_11797);
nor U11996 (N_11996,N_11697,N_11629);
or U11997 (N_11997,N_11792,N_11723);
nand U11998 (N_11998,N_11717,N_11785);
nor U11999 (N_11999,N_11746,N_11796);
nand U12000 (N_12000,N_11834,N_11840);
and U12001 (N_12001,N_11884,N_11958);
xnor U12002 (N_12002,N_11838,N_11855);
nor U12003 (N_12003,N_11868,N_11954);
xor U12004 (N_12004,N_11897,N_11896);
and U12005 (N_12005,N_11883,N_11909);
and U12006 (N_12006,N_11807,N_11942);
or U12007 (N_12007,N_11910,N_11922);
and U12008 (N_12008,N_11945,N_11949);
nor U12009 (N_12009,N_11819,N_11981);
or U12010 (N_12010,N_11972,N_11940);
xor U12011 (N_12011,N_11933,N_11913);
xnor U12012 (N_12012,N_11995,N_11965);
xor U12013 (N_12013,N_11917,N_11823);
nand U12014 (N_12014,N_11912,N_11944);
xor U12015 (N_12015,N_11880,N_11815);
xor U12016 (N_12016,N_11962,N_11953);
and U12017 (N_12017,N_11964,N_11980);
or U12018 (N_12018,N_11975,N_11996);
or U12019 (N_12019,N_11876,N_11899);
and U12020 (N_12020,N_11930,N_11820);
xnor U12021 (N_12021,N_11875,N_11803);
xor U12022 (N_12022,N_11984,N_11852);
or U12023 (N_12023,N_11987,N_11890);
xor U12024 (N_12024,N_11990,N_11902);
nor U12025 (N_12025,N_11998,N_11821);
or U12026 (N_12026,N_11889,N_11854);
nand U12027 (N_12027,N_11828,N_11918);
and U12028 (N_12028,N_11986,N_11825);
xor U12029 (N_12029,N_11859,N_11830);
and U12030 (N_12030,N_11991,N_11905);
or U12031 (N_12031,N_11911,N_11816);
nand U12032 (N_12032,N_11961,N_11812);
xor U12033 (N_12033,N_11814,N_11831);
and U12034 (N_12034,N_11973,N_11860);
and U12035 (N_12035,N_11824,N_11943);
nor U12036 (N_12036,N_11914,N_11806);
nand U12037 (N_12037,N_11841,N_11849);
xor U12038 (N_12038,N_11992,N_11866);
nor U12039 (N_12039,N_11861,N_11867);
nor U12040 (N_12040,N_11931,N_11941);
nand U12041 (N_12041,N_11809,N_11994);
and U12042 (N_12042,N_11808,N_11857);
nor U12043 (N_12043,N_11850,N_11811);
nand U12044 (N_12044,N_11813,N_11887);
nand U12045 (N_12045,N_11948,N_11862);
nor U12046 (N_12046,N_11937,N_11871);
and U12047 (N_12047,N_11983,N_11999);
and U12048 (N_12048,N_11919,N_11817);
or U12049 (N_12049,N_11835,N_11842);
nand U12050 (N_12050,N_11977,N_11951);
nand U12051 (N_12051,N_11960,N_11869);
or U12052 (N_12052,N_11970,N_11845);
xor U12053 (N_12053,N_11873,N_11928);
or U12054 (N_12054,N_11938,N_11870);
xnor U12055 (N_12055,N_11872,N_11885);
nand U12056 (N_12056,N_11847,N_11920);
and U12057 (N_12057,N_11935,N_11967);
nor U12058 (N_12058,N_11800,N_11924);
or U12059 (N_12059,N_11853,N_11959);
or U12060 (N_12060,N_11926,N_11929);
or U12061 (N_12061,N_11947,N_11925);
xnor U12062 (N_12062,N_11895,N_11974);
nand U12063 (N_12063,N_11907,N_11908);
nand U12064 (N_12064,N_11843,N_11955);
xnor U12065 (N_12065,N_11969,N_11879);
nand U12066 (N_12066,N_11985,N_11901);
nor U12067 (N_12067,N_11863,N_11932);
xnor U12068 (N_12068,N_11878,N_11968);
xnor U12069 (N_12069,N_11837,N_11833);
xnor U12070 (N_12070,N_11822,N_11978);
or U12071 (N_12071,N_11956,N_11818);
and U12072 (N_12072,N_11997,N_11939);
or U12073 (N_12073,N_11858,N_11946);
or U12074 (N_12074,N_11886,N_11971);
nor U12075 (N_12075,N_11810,N_11916);
xor U12076 (N_12076,N_11950,N_11856);
and U12077 (N_12077,N_11900,N_11952);
and U12078 (N_12078,N_11923,N_11836);
nand U12079 (N_12079,N_11826,N_11829);
nand U12080 (N_12080,N_11839,N_11851);
or U12081 (N_12081,N_11966,N_11846);
and U12082 (N_12082,N_11963,N_11874);
nand U12083 (N_12083,N_11934,N_11804);
and U12084 (N_12084,N_11898,N_11877);
xor U12085 (N_12085,N_11976,N_11805);
or U12086 (N_12086,N_11864,N_11891);
nand U12087 (N_12087,N_11848,N_11865);
or U12088 (N_12088,N_11903,N_11801);
xor U12089 (N_12089,N_11904,N_11936);
nand U12090 (N_12090,N_11993,N_11988);
or U12091 (N_12091,N_11893,N_11802);
and U12092 (N_12092,N_11989,N_11906);
xor U12093 (N_12093,N_11957,N_11892);
or U12094 (N_12094,N_11832,N_11888);
nand U12095 (N_12095,N_11882,N_11894);
and U12096 (N_12096,N_11982,N_11827);
xnor U12097 (N_12097,N_11979,N_11881);
nor U12098 (N_12098,N_11927,N_11921);
and U12099 (N_12099,N_11844,N_11915);
nor U12100 (N_12100,N_11886,N_11842);
xor U12101 (N_12101,N_11931,N_11864);
nand U12102 (N_12102,N_11991,N_11873);
and U12103 (N_12103,N_11919,N_11971);
nor U12104 (N_12104,N_11908,N_11800);
nor U12105 (N_12105,N_11848,N_11869);
or U12106 (N_12106,N_11891,N_11906);
nand U12107 (N_12107,N_11895,N_11832);
xor U12108 (N_12108,N_11975,N_11985);
or U12109 (N_12109,N_11962,N_11927);
and U12110 (N_12110,N_11918,N_11901);
nor U12111 (N_12111,N_11865,N_11949);
and U12112 (N_12112,N_11945,N_11814);
nand U12113 (N_12113,N_11957,N_11990);
nor U12114 (N_12114,N_11911,N_11886);
nor U12115 (N_12115,N_11865,N_11896);
xnor U12116 (N_12116,N_11809,N_11801);
or U12117 (N_12117,N_11880,N_11934);
or U12118 (N_12118,N_11908,N_11851);
and U12119 (N_12119,N_11808,N_11841);
nand U12120 (N_12120,N_11801,N_11963);
or U12121 (N_12121,N_11808,N_11815);
nor U12122 (N_12122,N_11807,N_11902);
xnor U12123 (N_12123,N_11867,N_11878);
nand U12124 (N_12124,N_11864,N_11947);
nor U12125 (N_12125,N_11970,N_11881);
or U12126 (N_12126,N_11935,N_11924);
nand U12127 (N_12127,N_11980,N_11804);
or U12128 (N_12128,N_11831,N_11829);
xnor U12129 (N_12129,N_11922,N_11987);
or U12130 (N_12130,N_11821,N_11972);
and U12131 (N_12131,N_11852,N_11949);
and U12132 (N_12132,N_11804,N_11955);
xnor U12133 (N_12133,N_11987,N_11995);
or U12134 (N_12134,N_11838,N_11800);
nand U12135 (N_12135,N_11950,N_11918);
and U12136 (N_12136,N_11951,N_11846);
nand U12137 (N_12137,N_11886,N_11838);
and U12138 (N_12138,N_11979,N_11880);
or U12139 (N_12139,N_11881,N_11991);
xnor U12140 (N_12140,N_11890,N_11939);
and U12141 (N_12141,N_11804,N_11886);
nor U12142 (N_12142,N_11877,N_11800);
nor U12143 (N_12143,N_11898,N_11917);
xnor U12144 (N_12144,N_11881,N_11833);
nand U12145 (N_12145,N_11890,N_11828);
xor U12146 (N_12146,N_11825,N_11951);
or U12147 (N_12147,N_11852,N_11933);
nor U12148 (N_12148,N_11828,N_11938);
nand U12149 (N_12149,N_11846,N_11827);
xor U12150 (N_12150,N_11961,N_11944);
or U12151 (N_12151,N_11811,N_11938);
and U12152 (N_12152,N_11973,N_11984);
or U12153 (N_12153,N_11819,N_11970);
nand U12154 (N_12154,N_11838,N_11873);
and U12155 (N_12155,N_11833,N_11887);
and U12156 (N_12156,N_11935,N_11989);
and U12157 (N_12157,N_11852,N_11886);
xor U12158 (N_12158,N_11875,N_11956);
nand U12159 (N_12159,N_11836,N_11956);
and U12160 (N_12160,N_11931,N_11844);
nand U12161 (N_12161,N_11942,N_11864);
and U12162 (N_12162,N_11909,N_11920);
nand U12163 (N_12163,N_11966,N_11882);
or U12164 (N_12164,N_11964,N_11901);
nand U12165 (N_12165,N_11999,N_11923);
or U12166 (N_12166,N_11932,N_11916);
nand U12167 (N_12167,N_11883,N_11803);
xor U12168 (N_12168,N_11884,N_11946);
nand U12169 (N_12169,N_11958,N_11983);
and U12170 (N_12170,N_11956,N_11940);
nor U12171 (N_12171,N_11814,N_11865);
and U12172 (N_12172,N_11924,N_11958);
nand U12173 (N_12173,N_11900,N_11813);
nor U12174 (N_12174,N_11941,N_11800);
and U12175 (N_12175,N_11812,N_11936);
nor U12176 (N_12176,N_11956,N_11800);
and U12177 (N_12177,N_11812,N_11869);
or U12178 (N_12178,N_11923,N_11888);
xnor U12179 (N_12179,N_11935,N_11821);
nand U12180 (N_12180,N_11949,N_11972);
nor U12181 (N_12181,N_11948,N_11930);
nand U12182 (N_12182,N_11924,N_11962);
or U12183 (N_12183,N_11982,N_11952);
nand U12184 (N_12184,N_11819,N_11900);
nor U12185 (N_12185,N_11802,N_11934);
xor U12186 (N_12186,N_11946,N_11970);
or U12187 (N_12187,N_11864,N_11923);
or U12188 (N_12188,N_11960,N_11975);
nand U12189 (N_12189,N_11974,N_11890);
nand U12190 (N_12190,N_11806,N_11985);
nand U12191 (N_12191,N_11844,N_11925);
or U12192 (N_12192,N_11961,N_11843);
or U12193 (N_12193,N_11925,N_11839);
nand U12194 (N_12194,N_11930,N_11894);
nor U12195 (N_12195,N_11931,N_11897);
nand U12196 (N_12196,N_11932,N_11841);
and U12197 (N_12197,N_11954,N_11953);
nand U12198 (N_12198,N_11808,N_11954);
xnor U12199 (N_12199,N_11862,N_11892);
nand U12200 (N_12200,N_12192,N_12150);
or U12201 (N_12201,N_12089,N_12051);
nand U12202 (N_12202,N_12030,N_12121);
or U12203 (N_12203,N_12129,N_12189);
or U12204 (N_12204,N_12055,N_12184);
and U12205 (N_12205,N_12146,N_12154);
and U12206 (N_12206,N_12163,N_12132);
or U12207 (N_12207,N_12080,N_12024);
nand U12208 (N_12208,N_12152,N_12036);
and U12209 (N_12209,N_12149,N_12137);
nand U12210 (N_12210,N_12028,N_12167);
nand U12211 (N_12211,N_12186,N_12006);
nand U12212 (N_12212,N_12044,N_12148);
and U12213 (N_12213,N_12175,N_12065);
or U12214 (N_12214,N_12013,N_12074);
nand U12215 (N_12215,N_12077,N_12156);
nand U12216 (N_12216,N_12011,N_12164);
and U12217 (N_12217,N_12101,N_12159);
and U12218 (N_12218,N_12168,N_12115);
and U12219 (N_12219,N_12079,N_12139);
nor U12220 (N_12220,N_12123,N_12086);
nor U12221 (N_12221,N_12094,N_12161);
nor U12222 (N_12222,N_12179,N_12068);
and U12223 (N_12223,N_12124,N_12076);
nor U12224 (N_12224,N_12185,N_12191);
nand U12225 (N_12225,N_12140,N_12003);
or U12226 (N_12226,N_12049,N_12022);
xor U12227 (N_12227,N_12195,N_12165);
or U12228 (N_12228,N_12048,N_12128);
or U12229 (N_12229,N_12045,N_12020);
nand U12230 (N_12230,N_12091,N_12016);
nor U12231 (N_12231,N_12052,N_12158);
nor U12232 (N_12232,N_12166,N_12078);
xor U12233 (N_12233,N_12084,N_12099);
and U12234 (N_12234,N_12176,N_12043);
xor U12235 (N_12235,N_12160,N_12182);
xor U12236 (N_12236,N_12112,N_12114);
and U12237 (N_12237,N_12180,N_12040);
or U12238 (N_12238,N_12187,N_12100);
or U12239 (N_12239,N_12083,N_12197);
or U12240 (N_12240,N_12183,N_12174);
xnor U12241 (N_12241,N_12014,N_12090);
nand U12242 (N_12242,N_12062,N_12023);
or U12243 (N_12243,N_12035,N_12029);
and U12244 (N_12244,N_12096,N_12144);
and U12245 (N_12245,N_12116,N_12178);
or U12246 (N_12246,N_12025,N_12138);
or U12247 (N_12247,N_12169,N_12073);
xnor U12248 (N_12248,N_12194,N_12153);
or U12249 (N_12249,N_12133,N_12075);
and U12250 (N_12250,N_12008,N_12193);
or U12251 (N_12251,N_12042,N_12041);
and U12252 (N_12252,N_12039,N_12111);
and U12253 (N_12253,N_12017,N_12050);
or U12254 (N_12254,N_12177,N_12059);
and U12255 (N_12255,N_12047,N_12000);
or U12256 (N_12256,N_12093,N_12141);
and U12257 (N_12257,N_12054,N_12012);
nor U12258 (N_12258,N_12001,N_12033);
nor U12259 (N_12259,N_12199,N_12102);
xor U12260 (N_12260,N_12151,N_12085);
nand U12261 (N_12261,N_12157,N_12155);
nand U12262 (N_12262,N_12097,N_12173);
xor U12263 (N_12263,N_12058,N_12119);
or U12264 (N_12264,N_12004,N_12181);
or U12265 (N_12265,N_12118,N_12147);
nand U12266 (N_12266,N_12027,N_12038);
nand U12267 (N_12267,N_12005,N_12127);
xor U12268 (N_12268,N_12057,N_12095);
xor U12269 (N_12269,N_12136,N_12046);
nand U12270 (N_12270,N_12130,N_12067);
or U12271 (N_12271,N_12108,N_12110);
and U12272 (N_12272,N_12010,N_12126);
or U12273 (N_12273,N_12103,N_12082);
nand U12274 (N_12274,N_12019,N_12092);
nor U12275 (N_12275,N_12117,N_12107);
xor U12276 (N_12276,N_12120,N_12190);
nor U12277 (N_12277,N_12125,N_12145);
nand U12278 (N_12278,N_12122,N_12134);
and U12279 (N_12279,N_12061,N_12071);
xnor U12280 (N_12280,N_12162,N_12081);
nor U12281 (N_12281,N_12198,N_12060);
xor U12282 (N_12282,N_12015,N_12069);
and U12283 (N_12283,N_12143,N_12172);
xnor U12284 (N_12284,N_12106,N_12018);
nand U12285 (N_12285,N_12188,N_12135);
nor U12286 (N_12286,N_12142,N_12105);
xor U12287 (N_12287,N_12064,N_12034);
xor U12288 (N_12288,N_12056,N_12170);
or U12289 (N_12289,N_12171,N_12026);
nand U12290 (N_12290,N_12037,N_12196);
and U12291 (N_12291,N_12072,N_12066);
xor U12292 (N_12292,N_12007,N_12032);
and U12293 (N_12293,N_12009,N_12113);
or U12294 (N_12294,N_12070,N_12021);
or U12295 (N_12295,N_12053,N_12002);
nand U12296 (N_12296,N_12088,N_12098);
nor U12297 (N_12297,N_12087,N_12104);
and U12298 (N_12298,N_12109,N_12063);
nand U12299 (N_12299,N_12131,N_12031);
nand U12300 (N_12300,N_12060,N_12071);
and U12301 (N_12301,N_12001,N_12096);
nor U12302 (N_12302,N_12084,N_12053);
nor U12303 (N_12303,N_12097,N_12019);
or U12304 (N_12304,N_12024,N_12123);
nand U12305 (N_12305,N_12184,N_12174);
xor U12306 (N_12306,N_12023,N_12122);
or U12307 (N_12307,N_12073,N_12072);
and U12308 (N_12308,N_12083,N_12134);
nand U12309 (N_12309,N_12118,N_12146);
nor U12310 (N_12310,N_12185,N_12173);
nand U12311 (N_12311,N_12091,N_12083);
nor U12312 (N_12312,N_12152,N_12176);
xor U12313 (N_12313,N_12079,N_12058);
xnor U12314 (N_12314,N_12121,N_12125);
xor U12315 (N_12315,N_12131,N_12160);
or U12316 (N_12316,N_12030,N_12064);
or U12317 (N_12317,N_12152,N_12114);
nand U12318 (N_12318,N_12152,N_12147);
nand U12319 (N_12319,N_12156,N_12009);
nand U12320 (N_12320,N_12094,N_12003);
or U12321 (N_12321,N_12019,N_12046);
and U12322 (N_12322,N_12154,N_12173);
nor U12323 (N_12323,N_12078,N_12115);
and U12324 (N_12324,N_12133,N_12073);
or U12325 (N_12325,N_12088,N_12029);
xor U12326 (N_12326,N_12078,N_12029);
nor U12327 (N_12327,N_12181,N_12029);
and U12328 (N_12328,N_12114,N_12186);
nor U12329 (N_12329,N_12002,N_12015);
and U12330 (N_12330,N_12189,N_12172);
and U12331 (N_12331,N_12131,N_12149);
nand U12332 (N_12332,N_12076,N_12053);
nand U12333 (N_12333,N_12051,N_12157);
nor U12334 (N_12334,N_12195,N_12051);
xnor U12335 (N_12335,N_12199,N_12076);
nor U12336 (N_12336,N_12184,N_12118);
nand U12337 (N_12337,N_12041,N_12169);
or U12338 (N_12338,N_12015,N_12129);
nand U12339 (N_12339,N_12085,N_12182);
xor U12340 (N_12340,N_12159,N_12183);
xnor U12341 (N_12341,N_12066,N_12149);
xnor U12342 (N_12342,N_12134,N_12073);
xor U12343 (N_12343,N_12136,N_12157);
or U12344 (N_12344,N_12152,N_12018);
nor U12345 (N_12345,N_12037,N_12166);
nand U12346 (N_12346,N_12127,N_12168);
and U12347 (N_12347,N_12195,N_12131);
and U12348 (N_12348,N_12031,N_12126);
or U12349 (N_12349,N_12004,N_12027);
and U12350 (N_12350,N_12093,N_12162);
or U12351 (N_12351,N_12006,N_12183);
xnor U12352 (N_12352,N_12140,N_12119);
nor U12353 (N_12353,N_12053,N_12117);
nand U12354 (N_12354,N_12004,N_12129);
xnor U12355 (N_12355,N_12096,N_12135);
or U12356 (N_12356,N_12158,N_12022);
and U12357 (N_12357,N_12032,N_12052);
or U12358 (N_12358,N_12067,N_12030);
nand U12359 (N_12359,N_12111,N_12003);
or U12360 (N_12360,N_12182,N_12178);
xor U12361 (N_12361,N_12034,N_12075);
or U12362 (N_12362,N_12153,N_12184);
nand U12363 (N_12363,N_12193,N_12125);
nand U12364 (N_12364,N_12146,N_12128);
xor U12365 (N_12365,N_12024,N_12151);
xor U12366 (N_12366,N_12092,N_12125);
nor U12367 (N_12367,N_12198,N_12037);
xor U12368 (N_12368,N_12018,N_12125);
xnor U12369 (N_12369,N_12007,N_12082);
or U12370 (N_12370,N_12141,N_12134);
and U12371 (N_12371,N_12125,N_12028);
xor U12372 (N_12372,N_12146,N_12055);
and U12373 (N_12373,N_12038,N_12156);
and U12374 (N_12374,N_12133,N_12155);
xnor U12375 (N_12375,N_12051,N_12098);
nor U12376 (N_12376,N_12065,N_12034);
and U12377 (N_12377,N_12140,N_12020);
nand U12378 (N_12378,N_12162,N_12198);
nand U12379 (N_12379,N_12154,N_12002);
nand U12380 (N_12380,N_12146,N_12125);
nor U12381 (N_12381,N_12175,N_12189);
xor U12382 (N_12382,N_12124,N_12002);
or U12383 (N_12383,N_12195,N_12008);
or U12384 (N_12384,N_12153,N_12185);
nor U12385 (N_12385,N_12053,N_12074);
nand U12386 (N_12386,N_12063,N_12166);
nand U12387 (N_12387,N_12158,N_12004);
nor U12388 (N_12388,N_12120,N_12189);
or U12389 (N_12389,N_12057,N_12016);
nand U12390 (N_12390,N_12190,N_12088);
nor U12391 (N_12391,N_12065,N_12137);
xnor U12392 (N_12392,N_12139,N_12119);
nor U12393 (N_12393,N_12102,N_12006);
xnor U12394 (N_12394,N_12053,N_12152);
or U12395 (N_12395,N_12127,N_12030);
and U12396 (N_12396,N_12162,N_12034);
xnor U12397 (N_12397,N_12125,N_12057);
xor U12398 (N_12398,N_12026,N_12043);
nor U12399 (N_12399,N_12012,N_12122);
xor U12400 (N_12400,N_12334,N_12318);
and U12401 (N_12401,N_12361,N_12202);
xor U12402 (N_12402,N_12223,N_12354);
xor U12403 (N_12403,N_12364,N_12211);
xnor U12404 (N_12404,N_12221,N_12250);
or U12405 (N_12405,N_12344,N_12206);
or U12406 (N_12406,N_12231,N_12262);
xnor U12407 (N_12407,N_12340,N_12298);
or U12408 (N_12408,N_12321,N_12357);
and U12409 (N_12409,N_12247,N_12261);
or U12410 (N_12410,N_12280,N_12390);
nor U12411 (N_12411,N_12311,N_12320);
xor U12412 (N_12412,N_12270,N_12382);
nand U12413 (N_12413,N_12315,N_12360);
nor U12414 (N_12414,N_12212,N_12260);
and U12415 (N_12415,N_12378,N_12345);
or U12416 (N_12416,N_12368,N_12338);
or U12417 (N_12417,N_12271,N_12233);
nor U12418 (N_12418,N_12375,N_12281);
nand U12419 (N_12419,N_12369,N_12241);
nand U12420 (N_12420,N_12339,N_12376);
nand U12421 (N_12421,N_12277,N_12331);
xnor U12422 (N_12422,N_12371,N_12297);
nor U12423 (N_12423,N_12324,N_12377);
xor U12424 (N_12424,N_12322,N_12227);
or U12425 (N_12425,N_12243,N_12294);
nand U12426 (N_12426,N_12356,N_12395);
or U12427 (N_12427,N_12259,N_12257);
and U12428 (N_12428,N_12200,N_12386);
or U12429 (N_12429,N_12353,N_12396);
xnor U12430 (N_12430,N_12374,N_12385);
or U12431 (N_12431,N_12240,N_12254);
nor U12432 (N_12432,N_12367,N_12303);
and U12433 (N_12433,N_12251,N_12279);
and U12434 (N_12434,N_12252,N_12319);
nor U12435 (N_12435,N_12235,N_12373);
nor U12436 (N_12436,N_12245,N_12276);
or U12437 (N_12437,N_12208,N_12226);
or U12438 (N_12438,N_12342,N_12236);
nor U12439 (N_12439,N_12242,N_12372);
or U12440 (N_12440,N_12292,N_12220);
nand U12441 (N_12441,N_12358,N_12238);
xor U12442 (N_12442,N_12326,N_12380);
xnor U12443 (N_12443,N_12268,N_12325);
and U12444 (N_12444,N_12203,N_12265);
and U12445 (N_12445,N_12218,N_12300);
and U12446 (N_12446,N_12215,N_12224);
nand U12447 (N_12447,N_12341,N_12228);
or U12448 (N_12448,N_12391,N_12316);
xnor U12449 (N_12449,N_12392,N_12301);
xor U12450 (N_12450,N_12350,N_12232);
and U12451 (N_12451,N_12327,N_12222);
xnor U12452 (N_12452,N_12379,N_12399);
xnor U12453 (N_12453,N_12388,N_12355);
nor U12454 (N_12454,N_12328,N_12216);
or U12455 (N_12455,N_12295,N_12349);
xnor U12456 (N_12456,N_12266,N_12205);
nand U12457 (N_12457,N_12393,N_12304);
nor U12458 (N_12458,N_12337,N_12230);
xnor U12459 (N_12459,N_12309,N_12217);
nor U12460 (N_12460,N_12283,N_12347);
xnor U12461 (N_12461,N_12397,N_12272);
xor U12462 (N_12462,N_12343,N_12201);
and U12463 (N_12463,N_12308,N_12351);
nand U12464 (N_12464,N_12306,N_12210);
nor U12465 (N_12465,N_12317,N_12290);
nand U12466 (N_12466,N_12287,N_12299);
or U12467 (N_12467,N_12264,N_12267);
or U12468 (N_12468,N_12313,N_12275);
or U12469 (N_12469,N_12307,N_12296);
nand U12470 (N_12470,N_12365,N_12282);
xor U12471 (N_12471,N_12381,N_12248);
xnor U12472 (N_12472,N_12293,N_12263);
nand U12473 (N_12473,N_12310,N_12289);
xnor U12474 (N_12474,N_12204,N_12219);
nor U12475 (N_12475,N_12366,N_12383);
and U12476 (N_12476,N_12305,N_12274);
nand U12477 (N_12477,N_12387,N_12255);
or U12478 (N_12478,N_12384,N_12323);
nor U12479 (N_12479,N_12285,N_12249);
and U12480 (N_12480,N_12346,N_12336);
nor U12481 (N_12481,N_12398,N_12253);
or U12482 (N_12482,N_12288,N_12237);
xnor U12483 (N_12483,N_12291,N_12362);
nand U12484 (N_12484,N_12225,N_12284);
xor U12485 (N_12485,N_12239,N_12269);
or U12486 (N_12486,N_12246,N_12335);
nand U12487 (N_12487,N_12359,N_12213);
nor U12488 (N_12488,N_12314,N_12286);
xnor U12489 (N_12489,N_12273,N_12394);
or U12490 (N_12490,N_12312,N_12209);
or U12491 (N_12491,N_12302,N_12348);
xnor U12492 (N_12492,N_12258,N_12370);
or U12493 (N_12493,N_12329,N_12244);
nor U12494 (N_12494,N_12352,N_12333);
nor U12495 (N_12495,N_12234,N_12207);
or U12496 (N_12496,N_12278,N_12389);
nor U12497 (N_12497,N_12332,N_12363);
nor U12498 (N_12498,N_12214,N_12229);
or U12499 (N_12499,N_12256,N_12330);
xor U12500 (N_12500,N_12290,N_12244);
nor U12501 (N_12501,N_12336,N_12304);
nor U12502 (N_12502,N_12357,N_12396);
and U12503 (N_12503,N_12246,N_12392);
nand U12504 (N_12504,N_12373,N_12399);
nand U12505 (N_12505,N_12220,N_12310);
or U12506 (N_12506,N_12292,N_12213);
nor U12507 (N_12507,N_12292,N_12377);
xor U12508 (N_12508,N_12293,N_12281);
and U12509 (N_12509,N_12367,N_12310);
nor U12510 (N_12510,N_12329,N_12379);
xnor U12511 (N_12511,N_12307,N_12237);
or U12512 (N_12512,N_12236,N_12270);
nand U12513 (N_12513,N_12367,N_12359);
xnor U12514 (N_12514,N_12345,N_12306);
nor U12515 (N_12515,N_12216,N_12332);
nor U12516 (N_12516,N_12309,N_12244);
or U12517 (N_12517,N_12315,N_12383);
nor U12518 (N_12518,N_12265,N_12309);
xor U12519 (N_12519,N_12300,N_12310);
and U12520 (N_12520,N_12259,N_12395);
xnor U12521 (N_12521,N_12225,N_12229);
xnor U12522 (N_12522,N_12229,N_12218);
nand U12523 (N_12523,N_12212,N_12217);
xnor U12524 (N_12524,N_12285,N_12261);
and U12525 (N_12525,N_12224,N_12323);
nand U12526 (N_12526,N_12228,N_12224);
and U12527 (N_12527,N_12380,N_12307);
nor U12528 (N_12528,N_12238,N_12373);
or U12529 (N_12529,N_12246,N_12339);
and U12530 (N_12530,N_12263,N_12267);
or U12531 (N_12531,N_12334,N_12217);
nor U12532 (N_12532,N_12292,N_12234);
and U12533 (N_12533,N_12205,N_12399);
nor U12534 (N_12534,N_12381,N_12269);
nor U12535 (N_12535,N_12368,N_12202);
xor U12536 (N_12536,N_12352,N_12358);
or U12537 (N_12537,N_12367,N_12364);
nor U12538 (N_12538,N_12363,N_12294);
xor U12539 (N_12539,N_12221,N_12397);
nand U12540 (N_12540,N_12270,N_12218);
nor U12541 (N_12541,N_12375,N_12283);
or U12542 (N_12542,N_12306,N_12215);
or U12543 (N_12543,N_12367,N_12211);
nand U12544 (N_12544,N_12200,N_12321);
and U12545 (N_12545,N_12336,N_12247);
or U12546 (N_12546,N_12242,N_12295);
nand U12547 (N_12547,N_12399,N_12285);
or U12548 (N_12548,N_12310,N_12282);
nor U12549 (N_12549,N_12275,N_12234);
and U12550 (N_12550,N_12272,N_12295);
or U12551 (N_12551,N_12326,N_12348);
or U12552 (N_12552,N_12359,N_12305);
xnor U12553 (N_12553,N_12290,N_12394);
nand U12554 (N_12554,N_12210,N_12227);
xor U12555 (N_12555,N_12237,N_12238);
xnor U12556 (N_12556,N_12231,N_12395);
nand U12557 (N_12557,N_12237,N_12244);
or U12558 (N_12558,N_12377,N_12274);
or U12559 (N_12559,N_12219,N_12291);
and U12560 (N_12560,N_12283,N_12298);
and U12561 (N_12561,N_12295,N_12285);
nand U12562 (N_12562,N_12337,N_12214);
or U12563 (N_12563,N_12255,N_12279);
or U12564 (N_12564,N_12219,N_12363);
and U12565 (N_12565,N_12274,N_12340);
nand U12566 (N_12566,N_12226,N_12326);
nor U12567 (N_12567,N_12381,N_12326);
nand U12568 (N_12568,N_12286,N_12307);
nand U12569 (N_12569,N_12303,N_12347);
nor U12570 (N_12570,N_12351,N_12361);
and U12571 (N_12571,N_12220,N_12396);
nor U12572 (N_12572,N_12218,N_12364);
and U12573 (N_12573,N_12257,N_12222);
or U12574 (N_12574,N_12339,N_12240);
or U12575 (N_12575,N_12379,N_12297);
or U12576 (N_12576,N_12278,N_12393);
nand U12577 (N_12577,N_12382,N_12241);
or U12578 (N_12578,N_12337,N_12360);
and U12579 (N_12579,N_12227,N_12361);
xor U12580 (N_12580,N_12288,N_12372);
nand U12581 (N_12581,N_12339,N_12218);
or U12582 (N_12582,N_12345,N_12308);
nand U12583 (N_12583,N_12235,N_12250);
nand U12584 (N_12584,N_12265,N_12325);
nand U12585 (N_12585,N_12354,N_12343);
and U12586 (N_12586,N_12214,N_12297);
nand U12587 (N_12587,N_12263,N_12336);
and U12588 (N_12588,N_12271,N_12397);
nor U12589 (N_12589,N_12348,N_12300);
nor U12590 (N_12590,N_12215,N_12216);
or U12591 (N_12591,N_12316,N_12348);
or U12592 (N_12592,N_12300,N_12220);
or U12593 (N_12593,N_12303,N_12255);
nor U12594 (N_12594,N_12341,N_12238);
xnor U12595 (N_12595,N_12398,N_12374);
and U12596 (N_12596,N_12262,N_12322);
nor U12597 (N_12597,N_12365,N_12217);
and U12598 (N_12598,N_12369,N_12269);
nor U12599 (N_12599,N_12398,N_12336);
nor U12600 (N_12600,N_12564,N_12419);
and U12601 (N_12601,N_12593,N_12576);
nand U12602 (N_12602,N_12490,N_12502);
xor U12603 (N_12603,N_12413,N_12529);
nand U12604 (N_12604,N_12483,N_12405);
and U12605 (N_12605,N_12526,N_12414);
and U12606 (N_12606,N_12591,N_12418);
and U12607 (N_12607,N_12474,N_12563);
or U12608 (N_12608,N_12545,N_12550);
nor U12609 (N_12609,N_12525,N_12470);
nand U12610 (N_12610,N_12507,N_12448);
nor U12611 (N_12611,N_12570,N_12439);
or U12612 (N_12612,N_12503,N_12513);
nor U12613 (N_12613,N_12595,N_12561);
nand U12614 (N_12614,N_12583,N_12520);
and U12615 (N_12615,N_12555,N_12530);
nor U12616 (N_12616,N_12435,N_12493);
xnor U12617 (N_12617,N_12572,N_12473);
nand U12618 (N_12618,N_12415,N_12598);
or U12619 (N_12619,N_12543,N_12592);
xor U12620 (N_12620,N_12425,N_12539);
and U12621 (N_12621,N_12577,N_12532);
or U12622 (N_12622,N_12587,N_12519);
and U12623 (N_12623,N_12417,N_12504);
xnor U12624 (N_12624,N_12581,N_12586);
nand U12625 (N_12625,N_12508,N_12452);
xor U12626 (N_12626,N_12449,N_12431);
nor U12627 (N_12627,N_12458,N_12516);
and U12628 (N_12628,N_12575,N_12485);
or U12629 (N_12629,N_12585,N_12552);
nor U12630 (N_12630,N_12498,N_12527);
xnor U12631 (N_12631,N_12544,N_12421);
nor U12632 (N_12632,N_12434,N_12432);
or U12633 (N_12633,N_12541,N_12588);
or U12634 (N_12634,N_12409,N_12487);
nor U12635 (N_12635,N_12565,N_12422);
nor U12636 (N_12636,N_12410,N_12568);
or U12637 (N_12637,N_12534,N_12590);
nor U12638 (N_12638,N_12482,N_12472);
nand U12639 (N_12639,N_12571,N_12496);
or U12640 (N_12640,N_12433,N_12535);
nand U12641 (N_12641,N_12491,N_12596);
and U12642 (N_12642,N_12465,N_12506);
nand U12643 (N_12643,N_12406,N_12478);
and U12644 (N_12644,N_12428,N_12430);
xnor U12645 (N_12645,N_12510,N_12479);
and U12646 (N_12646,N_12549,N_12408);
or U12647 (N_12647,N_12567,N_12492);
nand U12648 (N_12648,N_12521,N_12538);
and U12649 (N_12649,N_12442,N_12480);
or U12650 (N_12650,N_12411,N_12500);
nand U12651 (N_12651,N_12559,N_12443);
nand U12652 (N_12652,N_12468,N_12579);
nand U12653 (N_12653,N_12461,N_12589);
xor U12654 (N_12654,N_12540,N_12554);
xor U12655 (N_12655,N_12512,N_12416);
nor U12656 (N_12656,N_12584,N_12445);
nand U12657 (N_12657,N_12522,N_12558);
nand U12658 (N_12658,N_12488,N_12505);
and U12659 (N_12659,N_12412,N_12533);
nand U12660 (N_12660,N_12401,N_12489);
nor U12661 (N_12661,N_12517,N_12597);
and U12662 (N_12662,N_12569,N_12451);
nor U12663 (N_12663,N_12562,N_12573);
nand U12664 (N_12664,N_12557,N_12599);
nand U12665 (N_12665,N_12531,N_12536);
and U12666 (N_12666,N_12429,N_12481);
xor U12667 (N_12667,N_12440,N_12437);
nor U12668 (N_12668,N_12511,N_12403);
nand U12669 (N_12669,N_12537,N_12515);
nand U12670 (N_12670,N_12438,N_12464);
nor U12671 (N_12671,N_12453,N_12523);
xnor U12672 (N_12672,N_12466,N_12441);
or U12673 (N_12673,N_12594,N_12450);
nand U12674 (N_12674,N_12580,N_12444);
nor U12675 (N_12675,N_12475,N_12404);
xnor U12676 (N_12676,N_12547,N_12456);
and U12677 (N_12677,N_12518,N_12467);
xor U12678 (N_12678,N_12427,N_12524);
and U12679 (N_12679,N_12407,N_12497);
nor U12680 (N_12680,N_12471,N_12424);
or U12681 (N_12681,N_12454,N_12556);
nor U12682 (N_12682,N_12462,N_12566);
or U12683 (N_12683,N_12455,N_12426);
or U12684 (N_12684,N_12546,N_12423);
xor U12685 (N_12685,N_12463,N_12446);
xor U12686 (N_12686,N_12459,N_12551);
nand U12687 (N_12687,N_12476,N_12578);
and U12688 (N_12688,N_12484,N_12574);
nor U12689 (N_12689,N_12486,N_12499);
and U12690 (N_12690,N_12400,N_12460);
and U12691 (N_12691,N_12436,N_12528);
nor U12692 (N_12692,N_12501,N_12494);
nand U12693 (N_12693,N_12477,N_12560);
or U12694 (N_12694,N_12514,N_12469);
nand U12695 (N_12695,N_12457,N_12509);
and U12696 (N_12696,N_12548,N_12402);
xor U12697 (N_12697,N_12447,N_12542);
nand U12698 (N_12698,N_12420,N_12495);
or U12699 (N_12699,N_12582,N_12553);
xor U12700 (N_12700,N_12495,N_12570);
xor U12701 (N_12701,N_12594,N_12543);
or U12702 (N_12702,N_12547,N_12583);
or U12703 (N_12703,N_12433,N_12447);
nor U12704 (N_12704,N_12550,N_12534);
nor U12705 (N_12705,N_12424,N_12545);
xor U12706 (N_12706,N_12543,N_12544);
nor U12707 (N_12707,N_12593,N_12444);
nor U12708 (N_12708,N_12482,N_12438);
or U12709 (N_12709,N_12463,N_12543);
and U12710 (N_12710,N_12404,N_12572);
and U12711 (N_12711,N_12411,N_12459);
nor U12712 (N_12712,N_12527,N_12418);
xor U12713 (N_12713,N_12509,N_12521);
xor U12714 (N_12714,N_12484,N_12582);
or U12715 (N_12715,N_12466,N_12533);
xor U12716 (N_12716,N_12504,N_12405);
or U12717 (N_12717,N_12489,N_12481);
nand U12718 (N_12718,N_12544,N_12417);
or U12719 (N_12719,N_12555,N_12407);
nand U12720 (N_12720,N_12512,N_12425);
or U12721 (N_12721,N_12542,N_12442);
nor U12722 (N_12722,N_12519,N_12418);
or U12723 (N_12723,N_12441,N_12500);
nand U12724 (N_12724,N_12494,N_12446);
or U12725 (N_12725,N_12502,N_12575);
nor U12726 (N_12726,N_12416,N_12571);
nand U12727 (N_12727,N_12456,N_12494);
and U12728 (N_12728,N_12496,N_12594);
and U12729 (N_12729,N_12468,N_12557);
xnor U12730 (N_12730,N_12566,N_12400);
nor U12731 (N_12731,N_12453,N_12403);
nand U12732 (N_12732,N_12432,N_12429);
and U12733 (N_12733,N_12505,N_12471);
or U12734 (N_12734,N_12541,N_12510);
nand U12735 (N_12735,N_12570,N_12402);
nor U12736 (N_12736,N_12414,N_12418);
or U12737 (N_12737,N_12463,N_12529);
nor U12738 (N_12738,N_12422,N_12498);
or U12739 (N_12739,N_12500,N_12542);
xor U12740 (N_12740,N_12586,N_12429);
xnor U12741 (N_12741,N_12437,N_12590);
xor U12742 (N_12742,N_12444,N_12528);
or U12743 (N_12743,N_12518,N_12456);
xor U12744 (N_12744,N_12457,N_12503);
nor U12745 (N_12745,N_12542,N_12591);
nand U12746 (N_12746,N_12541,N_12527);
nor U12747 (N_12747,N_12529,N_12485);
nor U12748 (N_12748,N_12458,N_12594);
nand U12749 (N_12749,N_12432,N_12500);
and U12750 (N_12750,N_12446,N_12542);
xnor U12751 (N_12751,N_12401,N_12535);
nor U12752 (N_12752,N_12575,N_12524);
and U12753 (N_12753,N_12520,N_12591);
nand U12754 (N_12754,N_12525,N_12467);
xor U12755 (N_12755,N_12589,N_12433);
nand U12756 (N_12756,N_12577,N_12556);
nand U12757 (N_12757,N_12419,N_12453);
nor U12758 (N_12758,N_12527,N_12446);
nand U12759 (N_12759,N_12407,N_12459);
nor U12760 (N_12760,N_12564,N_12435);
xor U12761 (N_12761,N_12575,N_12514);
or U12762 (N_12762,N_12456,N_12402);
and U12763 (N_12763,N_12494,N_12556);
and U12764 (N_12764,N_12532,N_12417);
xor U12765 (N_12765,N_12587,N_12590);
and U12766 (N_12766,N_12562,N_12446);
or U12767 (N_12767,N_12504,N_12582);
xor U12768 (N_12768,N_12572,N_12577);
xor U12769 (N_12769,N_12568,N_12555);
or U12770 (N_12770,N_12410,N_12536);
xor U12771 (N_12771,N_12516,N_12597);
and U12772 (N_12772,N_12472,N_12411);
and U12773 (N_12773,N_12538,N_12440);
and U12774 (N_12774,N_12576,N_12415);
and U12775 (N_12775,N_12496,N_12588);
and U12776 (N_12776,N_12556,N_12549);
or U12777 (N_12777,N_12585,N_12529);
xor U12778 (N_12778,N_12558,N_12423);
or U12779 (N_12779,N_12590,N_12568);
xnor U12780 (N_12780,N_12562,N_12454);
nand U12781 (N_12781,N_12506,N_12565);
and U12782 (N_12782,N_12595,N_12479);
and U12783 (N_12783,N_12588,N_12563);
xnor U12784 (N_12784,N_12468,N_12452);
xnor U12785 (N_12785,N_12479,N_12412);
xnor U12786 (N_12786,N_12550,N_12540);
nor U12787 (N_12787,N_12486,N_12489);
nor U12788 (N_12788,N_12552,N_12447);
and U12789 (N_12789,N_12588,N_12527);
nand U12790 (N_12790,N_12480,N_12573);
xnor U12791 (N_12791,N_12487,N_12573);
nand U12792 (N_12792,N_12598,N_12503);
xnor U12793 (N_12793,N_12417,N_12596);
or U12794 (N_12794,N_12563,N_12448);
xnor U12795 (N_12795,N_12451,N_12496);
or U12796 (N_12796,N_12437,N_12581);
or U12797 (N_12797,N_12445,N_12459);
nor U12798 (N_12798,N_12456,N_12507);
and U12799 (N_12799,N_12417,N_12441);
nor U12800 (N_12800,N_12627,N_12691);
nand U12801 (N_12801,N_12726,N_12768);
or U12802 (N_12802,N_12723,N_12666);
nor U12803 (N_12803,N_12622,N_12614);
nand U12804 (N_12804,N_12668,N_12780);
nor U12805 (N_12805,N_12672,N_12739);
nor U12806 (N_12806,N_12718,N_12659);
xnor U12807 (N_12807,N_12655,N_12654);
nor U12808 (N_12808,N_12745,N_12634);
or U12809 (N_12809,N_12642,N_12651);
nand U12810 (N_12810,N_12727,N_12774);
or U12811 (N_12811,N_12664,N_12631);
nand U12812 (N_12812,N_12716,N_12736);
and U12813 (N_12813,N_12650,N_12677);
nand U12814 (N_12814,N_12725,N_12710);
nand U12815 (N_12815,N_12757,N_12635);
nand U12816 (N_12816,N_12630,N_12708);
nand U12817 (N_12817,N_12613,N_12619);
nor U12818 (N_12818,N_12660,N_12612);
nor U12819 (N_12819,N_12746,N_12738);
and U12820 (N_12820,N_12674,N_12759);
nor U12821 (N_12821,N_12706,N_12671);
xnor U12822 (N_12822,N_12724,N_12714);
or U12823 (N_12823,N_12741,N_12689);
or U12824 (N_12824,N_12644,N_12798);
nand U12825 (N_12825,N_12751,N_12643);
and U12826 (N_12826,N_12740,N_12719);
xor U12827 (N_12827,N_12787,N_12742);
or U12828 (N_12828,N_12600,N_12703);
nand U12829 (N_12829,N_12688,N_12624);
nor U12830 (N_12830,N_12779,N_12775);
xnor U12831 (N_12831,N_12670,N_12778);
nor U12832 (N_12832,N_12676,N_12784);
xnor U12833 (N_12833,N_12781,N_12733);
or U12834 (N_12834,N_12617,N_12653);
and U12835 (N_12835,N_12709,N_12734);
and U12836 (N_12836,N_12783,N_12773);
nand U12837 (N_12837,N_12683,N_12770);
xnor U12838 (N_12838,N_12645,N_12638);
nand U12839 (N_12839,N_12731,N_12662);
nor U12840 (N_12840,N_12648,N_12609);
or U12841 (N_12841,N_12762,N_12690);
and U12842 (N_12842,N_12789,N_12603);
nand U12843 (N_12843,N_12767,N_12754);
nor U12844 (N_12844,N_12712,N_12679);
nand U12845 (N_12845,N_12737,N_12799);
nor U12846 (N_12846,N_12607,N_12637);
nor U12847 (N_12847,N_12735,N_12615);
xor U12848 (N_12848,N_12728,N_12639);
nor U12849 (N_12849,N_12629,N_12702);
and U12850 (N_12850,N_12772,N_12658);
nand U12851 (N_12851,N_12730,N_12667);
and U12852 (N_12852,N_12608,N_12752);
or U12853 (N_12853,N_12663,N_12625);
nor U12854 (N_12854,N_12758,N_12766);
xor U12855 (N_12855,N_12685,N_12687);
nand U12856 (N_12856,N_12711,N_12753);
nor U12857 (N_12857,N_12649,N_12760);
and U12858 (N_12858,N_12755,N_12606);
or U12859 (N_12859,N_12701,N_12729);
or U12860 (N_12860,N_12682,N_12747);
and U12861 (N_12861,N_12678,N_12681);
xnor U12862 (N_12862,N_12626,N_12633);
nor U12863 (N_12863,N_12704,N_12748);
and U12864 (N_12864,N_12669,N_12697);
nor U12865 (N_12865,N_12769,N_12623);
nand U12866 (N_12866,N_12698,N_12761);
and U12867 (N_12867,N_12616,N_12610);
or U12868 (N_12868,N_12700,N_12797);
nand U12869 (N_12869,N_12665,N_12791);
or U12870 (N_12870,N_12652,N_12602);
nor U12871 (N_12871,N_12765,N_12796);
or U12872 (N_12872,N_12722,N_12713);
nor U12873 (N_12873,N_12686,N_12720);
nand U12874 (N_12874,N_12777,N_12661);
nand U12875 (N_12875,N_12657,N_12794);
nand U12876 (N_12876,N_12786,N_12771);
nand U12877 (N_12877,N_12605,N_12715);
nor U12878 (N_12878,N_12750,N_12707);
and U12879 (N_12879,N_12788,N_12695);
nor U12880 (N_12880,N_12620,N_12647);
or U12881 (N_12881,N_12749,N_12611);
xor U12882 (N_12882,N_12744,N_12705);
nor U12883 (N_12883,N_12776,N_12636);
xnor U12884 (N_12884,N_12721,N_12717);
xor U12885 (N_12885,N_12694,N_12792);
or U12886 (N_12886,N_12782,N_12628);
xor U12887 (N_12887,N_12696,N_12675);
nand U12888 (N_12888,N_12673,N_12646);
nand U12889 (N_12889,N_12732,N_12601);
or U12890 (N_12890,N_12656,N_12684);
nand U12891 (N_12891,N_12790,N_12618);
nor U12892 (N_12892,N_12699,N_12756);
nand U12893 (N_12893,N_12795,N_12621);
and U12894 (N_12894,N_12764,N_12680);
xor U12895 (N_12895,N_12632,N_12763);
and U12896 (N_12896,N_12693,N_12793);
nor U12897 (N_12897,N_12785,N_12692);
nor U12898 (N_12898,N_12640,N_12641);
or U12899 (N_12899,N_12604,N_12743);
xnor U12900 (N_12900,N_12630,N_12676);
or U12901 (N_12901,N_12733,N_12751);
and U12902 (N_12902,N_12673,N_12702);
nand U12903 (N_12903,N_12653,N_12695);
nand U12904 (N_12904,N_12712,N_12780);
nor U12905 (N_12905,N_12720,N_12659);
xor U12906 (N_12906,N_12605,N_12770);
xnor U12907 (N_12907,N_12645,N_12655);
or U12908 (N_12908,N_12735,N_12671);
or U12909 (N_12909,N_12767,N_12657);
nand U12910 (N_12910,N_12637,N_12688);
nor U12911 (N_12911,N_12635,N_12639);
nor U12912 (N_12912,N_12760,N_12720);
nand U12913 (N_12913,N_12600,N_12700);
or U12914 (N_12914,N_12713,N_12728);
nand U12915 (N_12915,N_12627,N_12719);
or U12916 (N_12916,N_12775,N_12748);
nor U12917 (N_12917,N_12726,N_12624);
nand U12918 (N_12918,N_12779,N_12786);
and U12919 (N_12919,N_12714,N_12779);
and U12920 (N_12920,N_12669,N_12632);
xor U12921 (N_12921,N_12780,N_12789);
or U12922 (N_12922,N_12714,N_12782);
and U12923 (N_12923,N_12711,N_12600);
nor U12924 (N_12924,N_12781,N_12798);
nand U12925 (N_12925,N_12765,N_12632);
nor U12926 (N_12926,N_12778,N_12748);
or U12927 (N_12927,N_12755,N_12711);
xnor U12928 (N_12928,N_12727,N_12688);
nor U12929 (N_12929,N_12616,N_12698);
or U12930 (N_12930,N_12715,N_12709);
nor U12931 (N_12931,N_12740,N_12662);
or U12932 (N_12932,N_12680,N_12612);
xor U12933 (N_12933,N_12787,N_12762);
nand U12934 (N_12934,N_12705,N_12723);
nand U12935 (N_12935,N_12774,N_12689);
xnor U12936 (N_12936,N_12620,N_12762);
and U12937 (N_12937,N_12683,N_12697);
nor U12938 (N_12938,N_12601,N_12603);
or U12939 (N_12939,N_12611,N_12632);
and U12940 (N_12940,N_12712,N_12655);
and U12941 (N_12941,N_12773,N_12645);
and U12942 (N_12942,N_12642,N_12772);
xor U12943 (N_12943,N_12739,N_12767);
and U12944 (N_12944,N_12698,N_12671);
nor U12945 (N_12945,N_12696,N_12617);
and U12946 (N_12946,N_12745,N_12736);
nor U12947 (N_12947,N_12680,N_12683);
xnor U12948 (N_12948,N_12689,N_12634);
or U12949 (N_12949,N_12740,N_12669);
nand U12950 (N_12950,N_12612,N_12609);
or U12951 (N_12951,N_12621,N_12758);
or U12952 (N_12952,N_12760,N_12767);
xnor U12953 (N_12953,N_12636,N_12648);
or U12954 (N_12954,N_12798,N_12776);
nand U12955 (N_12955,N_12714,N_12614);
xnor U12956 (N_12956,N_12639,N_12722);
nor U12957 (N_12957,N_12617,N_12639);
nor U12958 (N_12958,N_12751,N_12731);
nand U12959 (N_12959,N_12601,N_12735);
nor U12960 (N_12960,N_12641,N_12675);
and U12961 (N_12961,N_12706,N_12602);
and U12962 (N_12962,N_12782,N_12613);
xnor U12963 (N_12963,N_12773,N_12754);
and U12964 (N_12964,N_12731,N_12645);
and U12965 (N_12965,N_12716,N_12766);
or U12966 (N_12966,N_12732,N_12785);
nor U12967 (N_12967,N_12773,N_12621);
and U12968 (N_12968,N_12735,N_12644);
and U12969 (N_12969,N_12768,N_12692);
or U12970 (N_12970,N_12768,N_12646);
and U12971 (N_12971,N_12682,N_12744);
nand U12972 (N_12972,N_12659,N_12615);
or U12973 (N_12973,N_12606,N_12703);
nand U12974 (N_12974,N_12704,N_12607);
xnor U12975 (N_12975,N_12602,N_12603);
nor U12976 (N_12976,N_12622,N_12681);
xnor U12977 (N_12977,N_12686,N_12729);
or U12978 (N_12978,N_12739,N_12697);
nand U12979 (N_12979,N_12718,N_12668);
xor U12980 (N_12980,N_12761,N_12655);
and U12981 (N_12981,N_12643,N_12633);
nand U12982 (N_12982,N_12751,N_12715);
or U12983 (N_12983,N_12793,N_12771);
nor U12984 (N_12984,N_12784,N_12731);
xnor U12985 (N_12985,N_12704,N_12686);
nor U12986 (N_12986,N_12629,N_12618);
nand U12987 (N_12987,N_12624,N_12606);
and U12988 (N_12988,N_12715,N_12717);
and U12989 (N_12989,N_12788,N_12771);
xnor U12990 (N_12990,N_12626,N_12643);
and U12991 (N_12991,N_12730,N_12622);
or U12992 (N_12992,N_12698,N_12680);
and U12993 (N_12993,N_12676,N_12604);
or U12994 (N_12994,N_12634,N_12619);
and U12995 (N_12995,N_12766,N_12749);
or U12996 (N_12996,N_12627,N_12713);
and U12997 (N_12997,N_12704,N_12608);
xnor U12998 (N_12998,N_12692,N_12601);
nor U12999 (N_12999,N_12610,N_12777);
and U13000 (N_13000,N_12880,N_12892);
and U13001 (N_13001,N_12853,N_12976);
or U13002 (N_13002,N_12820,N_12850);
xnor U13003 (N_13003,N_12920,N_12837);
xor U13004 (N_13004,N_12848,N_12942);
or U13005 (N_13005,N_12830,N_12899);
nand U13006 (N_13006,N_12808,N_12861);
nand U13007 (N_13007,N_12987,N_12950);
nor U13008 (N_13008,N_12862,N_12944);
xnor U13009 (N_13009,N_12904,N_12824);
nand U13010 (N_13010,N_12891,N_12969);
nand U13011 (N_13011,N_12878,N_12807);
nand U13012 (N_13012,N_12858,N_12919);
xor U13013 (N_13013,N_12970,N_12887);
nor U13014 (N_13014,N_12903,N_12957);
nand U13015 (N_13015,N_12869,N_12995);
and U13016 (N_13016,N_12872,N_12800);
or U13017 (N_13017,N_12963,N_12962);
or U13018 (N_13018,N_12926,N_12803);
nand U13019 (N_13019,N_12985,N_12849);
nand U13020 (N_13020,N_12817,N_12806);
and U13021 (N_13021,N_12843,N_12916);
and U13022 (N_13022,N_12941,N_12959);
and U13023 (N_13023,N_12825,N_12992);
and U13024 (N_13024,N_12874,N_12998);
or U13025 (N_13025,N_12821,N_12993);
nor U13026 (N_13026,N_12945,N_12988);
and U13027 (N_13027,N_12936,N_12871);
nand U13028 (N_13028,N_12822,N_12917);
nand U13029 (N_13029,N_12990,N_12951);
or U13030 (N_13030,N_12881,N_12828);
nor U13031 (N_13031,N_12896,N_12938);
nand U13032 (N_13032,N_12856,N_12816);
or U13033 (N_13033,N_12986,N_12860);
nor U13034 (N_13034,N_12973,N_12956);
nor U13035 (N_13035,N_12996,N_12979);
or U13036 (N_13036,N_12894,N_12876);
and U13037 (N_13037,N_12929,N_12813);
and U13038 (N_13038,N_12935,N_12922);
xnor U13039 (N_13039,N_12905,N_12918);
and U13040 (N_13040,N_12831,N_12930);
nand U13041 (N_13041,N_12826,N_12984);
or U13042 (N_13042,N_12863,N_12840);
or U13043 (N_13043,N_12931,N_12851);
xor U13044 (N_13044,N_12827,N_12835);
or U13045 (N_13045,N_12818,N_12964);
xor U13046 (N_13046,N_12801,N_12805);
or U13047 (N_13047,N_12940,N_12909);
nand U13048 (N_13048,N_12804,N_12855);
nand U13049 (N_13049,N_12847,N_12983);
nor U13050 (N_13050,N_12997,N_12852);
and U13051 (N_13051,N_12972,N_12939);
nor U13052 (N_13052,N_12921,N_12839);
and U13053 (N_13053,N_12955,N_12902);
nor U13054 (N_13054,N_12865,N_12967);
and U13055 (N_13055,N_12927,N_12980);
nor U13056 (N_13056,N_12923,N_12906);
or U13057 (N_13057,N_12991,N_12974);
xnor U13058 (N_13058,N_12836,N_12965);
xnor U13059 (N_13059,N_12867,N_12932);
nor U13060 (N_13060,N_12802,N_12908);
and U13061 (N_13061,N_12833,N_12966);
nand U13062 (N_13062,N_12947,N_12819);
xor U13063 (N_13063,N_12900,N_12933);
nand U13064 (N_13064,N_12829,N_12814);
nand U13065 (N_13065,N_12961,N_12893);
or U13066 (N_13066,N_12994,N_12924);
or U13067 (N_13067,N_12915,N_12968);
xor U13068 (N_13068,N_12913,N_12890);
nand U13069 (N_13069,N_12879,N_12812);
nand U13070 (N_13070,N_12999,N_12884);
or U13071 (N_13071,N_12832,N_12885);
and U13072 (N_13072,N_12857,N_12907);
nor U13073 (N_13073,N_12886,N_12977);
nor U13074 (N_13074,N_12834,N_12952);
nor U13075 (N_13075,N_12859,N_12889);
or U13076 (N_13076,N_12911,N_12982);
xnor U13077 (N_13077,N_12888,N_12989);
or U13078 (N_13078,N_12811,N_12910);
and U13079 (N_13079,N_12971,N_12866);
or U13080 (N_13080,N_12958,N_12914);
and U13081 (N_13081,N_12875,N_12841);
nand U13082 (N_13082,N_12912,N_12953);
nand U13083 (N_13083,N_12895,N_12810);
or U13084 (N_13084,N_12901,N_12838);
and U13085 (N_13085,N_12960,N_12897);
and U13086 (N_13086,N_12949,N_12873);
and U13087 (N_13087,N_12868,N_12975);
xor U13088 (N_13088,N_12870,N_12934);
nor U13089 (N_13089,N_12978,N_12815);
or U13090 (N_13090,N_12823,N_12954);
nand U13091 (N_13091,N_12943,N_12898);
xor U13092 (N_13092,N_12809,N_12846);
nor U13093 (N_13093,N_12864,N_12928);
nor U13094 (N_13094,N_12948,N_12844);
and U13095 (N_13095,N_12877,N_12937);
or U13096 (N_13096,N_12981,N_12882);
nor U13097 (N_13097,N_12854,N_12883);
nand U13098 (N_13098,N_12842,N_12946);
or U13099 (N_13099,N_12925,N_12845);
or U13100 (N_13100,N_12899,N_12901);
nand U13101 (N_13101,N_12966,N_12940);
or U13102 (N_13102,N_12963,N_12821);
or U13103 (N_13103,N_12978,N_12895);
or U13104 (N_13104,N_12961,N_12875);
nor U13105 (N_13105,N_12960,N_12890);
nor U13106 (N_13106,N_12827,N_12833);
or U13107 (N_13107,N_12940,N_12834);
and U13108 (N_13108,N_12854,N_12824);
nand U13109 (N_13109,N_12919,N_12941);
xnor U13110 (N_13110,N_12887,N_12938);
xor U13111 (N_13111,N_12916,N_12815);
nand U13112 (N_13112,N_12912,N_12914);
and U13113 (N_13113,N_12851,N_12999);
nor U13114 (N_13114,N_12873,N_12839);
xnor U13115 (N_13115,N_12960,N_12984);
xnor U13116 (N_13116,N_12926,N_12896);
and U13117 (N_13117,N_12972,N_12867);
nand U13118 (N_13118,N_12969,N_12883);
nand U13119 (N_13119,N_12955,N_12891);
or U13120 (N_13120,N_12951,N_12903);
nand U13121 (N_13121,N_12918,N_12928);
xor U13122 (N_13122,N_12819,N_12918);
xnor U13123 (N_13123,N_12815,N_12804);
or U13124 (N_13124,N_12991,N_12927);
nand U13125 (N_13125,N_12991,N_12841);
or U13126 (N_13126,N_12936,N_12948);
nor U13127 (N_13127,N_12982,N_12869);
or U13128 (N_13128,N_12880,N_12916);
and U13129 (N_13129,N_12944,N_12884);
and U13130 (N_13130,N_12984,N_12875);
nor U13131 (N_13131,N_12875,N_12903);
xor U13132 (N_13132,N_12860,N_12952);
and U13133 (N_13133,N_12945,N_12883);
nand U13134 (N_13134,N_12988,N_12875);
xnor U13135 (N_13135,N_12838,N_12869);
or U13136 (N_13136,N_12807,N_12816);
xnor U13137 (N_13137,N_12822,N_12958);
xor U13138 (N_13138,N_12889,N_12918);
and U13139 (N_13139,N_12893,N_12805);
nand U13140 (N_13140,N_12948,N_12801);
or U13141 (N_13141,N_12859,N_12802);
or U13142 (N_13142,N_12891,N_12972);
nor U13143 (N_13143,N_12995,N_12887);
or U13144 (N_13144,N_12812,N_12942);
nand U13145 (N_13145,N_12987,N_12973);
xor U13146 (N_13146,N_12870,N_12988);
xor U13147 (N_13147,N_12936,N_12865);
nand U13148 (N_13148,N_12808,N_12959);
or U13149 (N_13149,N_12916,N_12937);
and U13150 (N_13150,N_12907,N_12975);
nand U13151 (N_13151,N_12812,N_12821);
and U13152 (N_13152,N_12880,N_12962);
nand U13153 (N_13153,N_12941,N_12991);
or U13154 (N_13154,N_12848,N_12819);
xnor U13155 (N_13155,N_12978,N_12951);
xor U13156 (N_13156,N_12955,N_12992);
or U13157 (N_13157,N_12927,N_12998);
nand U13158 (N_13158,N_12999,N_12804);
nand U13159 (N_13159,N_12808,N_12851);
nor U13160 (N_13160,N_12826,N_12999);
nand U13161 (N_13161,N_12828,N_12929);
or U13162 (N_13162,N_12971,N_12943);
xor U13163 (N_13163,N_12810,N_12952);
xnor U13164 (N_13164,N_12937,N_12810);
xnor U13165 (N_13165,N_12965,N_12875);
xnor U13166 (N_13166,N_12858,N_12930);
or U13167 (N_13167,N_12852,N_12902);
xnor U13168 (N_13168,N_12833,N_12995);
nor U13169 (N_13169,N_12820,N_12812);
or U13170 (N_13170,N_12910,N_12882);
nand U13171 (N_13171,N_12955,N_12810);
nor U13172 (N_13172,N_12890,N_12984);
xor U13173 (N_13173,N_12914,N_12943);
and U13174 (N_13174,N_12823,N_12806);
nand U13175 (N_13175,N_12990,N_12894);
nor U13176 (N_13176,N_12800,N_12819);
and U13177 (N_13177,N_12897,N_12912);
nand U13178 (N_13178,N_12951,N_12976);
or U13179 (N_13179,N_12904,N_12927);
nand U13180 (N_13180,N_12984,N_12801);
or U13181 (N_13181,N_12938,N_12870);
or U13182 (N_13182,N_12864,N_12926);
or U13183 (N_13183,N_12838,N_12801);
and U13184 (N_13184,N_12804,N_12988);
nand U13185 (N_13185,N_12864,N_12851);
or U13186 (N_13186,N_12872,N_12804);
nor U13187 (N_13187,N_12816,N_12980);
nand U13188 (N_13188,N_12849,N_12851);
or U13189 (N_13189,N_12933,N_12885);
xnor U13190 (N_13190,N_12985,N_12809);
xor U13191 (N_13191,N_12996,N_12993);
and U13192 (N_13192,N_12896,N_12839);
and U13193 (N_13193,N_12984,N_12971);
nor U13194 (N_13194,N_12919,N_12864);
nor U13195 (N_13195,N_12893,N_12836);
nand U13196 (N_13196,N_12989,N_12912);
nand U13197 (N_13197,N_12820,N_12860);
or U13198 (N_13198,N_12802,N_12810);
xor U13199 (N_13199,N_12828,N_12801);
nor U13200 (N_13200,N_13126,N_13013);
xor U13201 (N_13201,N_13174,N_13106);
nand U13202 (N_13202,N_13093,N_13070);
xor U13203 (N_13203,N_13137,N_13143);
xnor U13204 (N_13204,N_13109,N_13132);
nand U13205 (N_13205,N_13134,N_13122);
and U13206 (N_13206,N_13120,N_13113);
or U13207 (N_13207,N_13035,N_13087);
nor U13208 (N_13208,N_13052,N_13107);
xnor U13209 (N_13209,N_13181,N_13004);
nor U13210 (N_13210,N_13007,N_13168);
nor U13211 (N_13211,N_13149,N_13179);
or U13212 (N_13212,N_13001,N_13102);
nand U13213 (N_13213,N_13025,N_13034);
or U13214 (N_13214,N_13196,N_13129);
xnor U13215 (N_13215,N_13154,N_13145);
nor U13216 (N_13216,N_13158,N_13095);
and U13217 (N_13217,N_13119,N_13186);
xnor U13218 (N_13218,N_13063,N_13199);
nor U13219 (N_13219,N_13178,N_13116);
and U13220 (N_13220,N_13036,N_13068);
or U13221 (N_13221,N_13131,N_13051);
or U13222 (N_13222,N_13194,N_13108);
nor U13223 (N_13223,N_13096,N_13086);
xnor U13224 (N_13224,N_13053,N_13138);
xor U13225 (N_13225,N_13136,N_13082);
and U13226 (N_13226,N_13188,N_13163);
nand U13227 (N_13227,N_13049,N_13077);
xnor U13228 (N_13228,N_13110,N_13187);
xor U13229 (N_13229,N_13060,N_13080);
or U13230 (N_13230,N_13084,N_13130);
and U13231 (N_13231,N_13005,N_13081);
nand U13232 (N_13232,N_13159,N_13195);
or U13233 (N_13233,N_13198,N_13044);
nand U13234 (N_13234,N_13105,N_13073);
and U13235 (N_13235,N_13020,N_13016);
nor U13236 (N_13236,N_13160,N_13058);
nor U13237 (N_13237,N_13041,N_13065);
and U13238 (N_13238,N_13114,N_13164);
xor U13239 (N_13239,N_13031,N_13165);
xor U13240 (N_13240,N_13040,N_13103);
nand U13241 (N_13241,N_13062,N_13017);
nand U13242 (N_13242,N_13072,N_13183);
nor U13243 (N_13243,N_13182,N_13140);
nor U13244 (N_13244,N_13150,N_13184);
xor U13245 (N_13245,N_13045,N_13144);
nand U13246 (N_13246,N_13047,N_13028);
nand U13247 (N_13247,N_13043,N_13000);
nor U13248 (N_13248,N_13092,N_13046);
or U13249 (N_13249,N_13173,N_13079);
or U13250 (N_13250,N_13139,N_13148);
nand U13251 (N_13251,N_13177,N_13094);
nor U13252 (N_13252,N_13078,N_13147);
or U13253 (N_13253,N_13191,N_13112);
and U13254 (N_13254,N_13115,N_13010);
nor U13255 (N_13255,N_13076,N_13056);
and U13256 (N_13256,N_13161,N_13142);
nand U13257 (N_13257,N_13064,N_13111);
or U13258 (N_13258,N_13071,N_13155);
nor U13259 (N_13259,N_13097,N_13133);
nor U13260 (N_13260,N_13170,N_13121);
or U13261 (N_13261,N_13128,N_13171);
or U13262 (N_13262,N_13037,N_13029);
nor U13263 (N_13263,N_13015,N_13061);
or U13264 (N_13264,N_13156,N_13185);
and U13265 (N_13265,N_13011,N_13176);
nor U13266 (N_13266,N_13162,N_13033);
nand U13267 (N_13267,N_13090,N_13039);
xor U13268 (N_13268,N_13098,N_13002);
nor U13269 (N_13269,N_13172,N_13153);
or U13270 (N_13270,N_13123,N_13009);
nor U13271 (N_13271,N_13069,N_13151);
and U13272 (N_13272,N_13019,N_13021);
nor U13273 (N_13273,N_13124,N_13135);
xnor U13274 (N_13274,N_13038,N_13030);
xor U13275 (N_13275,N_13193,N_13085);
and U13276 (N_13276,N_13166,N_13101);
or U13277 (N_13277,N_13104,N_13057);
nand U13278 (N_13278,N_13175,N_13008);
or U13279 (N_13279,N_13088,N_13190);
nor U13280 (N_13280,N_13012,N_13167);
or U13281 (N_13281,N_13023,N_13024);
or U13282 (N_13282,N_13146,N_13022);
xnor U13283 (N_13283,N_13066,N_13055);
nand U13284 (N_13284,N_13026,N_13075);
nor U13285 (N_13285,N_13192,N_13042);
xnor U13286 (N_13286,N_13048,N_13127);
and U13287 (N_13287,N_13018,N_13054);
nand U13288 (N_13288,N_13091,N_13100);
and U13289 (N_13289,N_13074,N_13067);
nand U13290 (N_13290,N_13180,N_13089);
xnor U13291 (N_13291,N_13125,N_13083);
or U13292 (N_13292,N_13059,N_13003);
or U13293 (N_13293,N_13197,N_13099);
xnor U13294 (N_13294,N_13169,N_13027);
and U13295 (N_13295,N_13050,N_13014);
or U13296 (N_13296,N_13032,N_13118);
and U13297 (N_13297,N_13117,N_13141);
nand U13298 (N_13298,N_13006,N_13157);
nand U13299 (N_13299,N_13152,N_13189);
nor U13300 (N_13300,N_13107,N_13174);
xnor U13301 (N_13301,N_13014,N_13185);
xnor U13302 (N_13302,N_13026,N_13129);
or U13303 (N_13303,N_13189,N_13097);
and U13304 (N_13304,N_13069,N_13053);
and U13305 (N_13305,N_13037,N_13146);
nand U13306 (N_13306,N_13187,N_13132);
or U13307 (N_13307,N_13084,N_13153);
and U13308 (N_13308,N_13075,N_13125);
or U13309 (N_13309,N_13057,N_13012);
nor U13310 (N_13310,N_13157,N_13165);
or U13311 (N_13311,N_13198,N_13064);
nor U13312 (N_13312,N_13077,N_13000);
and U13313 (N_13313,N_13159,N_13128);
or U13314 (N_13314,N_13027,N_13124);
nand U13315 (N_13315,N_13163,N_13004);
or U13316 (N_13316,N_13163,N_13140);
or U13317 (N_13317,N_13044,N_13160);
and U13318 (N_13318,N_13033,N_13198);
or U13319 (N_13319,N_13087,N_13107);
nand U13320 (N_13320,N_13079,N_13100);
nand U13321 (N_13321,N_13086,N_13072);
nand U13322 (N_13322,N_13008,N_13002);
or U13323 (N_13323,N_13028,N_13144);
nor U13324 (N_13324,N_13176,N_13151);
nand U13325 (N_13325,N_13012,N_13160);
nand U13326 (N_13326,N_13114,N_13156);
xor U13327 (N_13327,N_13105,N_13180);
nand U13328 (N_13328,N_13194,N_13012);
and U13329 (N_13329,N_13003,N_13035);
nor U13330 (N_13330,N_13071,N_13009);
or U13331 (N_13331,N_13099,N_13111);
nor U13332 (N_13332,N_13048,N_13038);
nor U13333 (N_13333,N_13085,N_13135);
xor U13334 (N_13334,N_13191,N_13002);
nand U13335 (N_13335,N_13189,N_13050);
nor U13336 (N_13336,N_13136,N_13183);
xor U13337 (N_13337,N_13097,N_13047);
and U13338 (N_13338,N_13043,N_13034);
nor U13339 (N_13339,N_13101,N_13165);
or U13340 (N_13340,N_13086,N_13133);
and U13341 (N_13341,N_13176,N_13024);
or U13342 (N_13342,N_13060,N_13138);
nand U13343 (N_13343,N_13006,N_13029);
xnor U13344 (N_13344,N_13016,N_13087);
nor U13345 (N_13345,N_13079,N_13072);
or U13346 (N_13346,N_13194,N_13150);
or U13347 (N_13347,N_13128,N_13007);
nand U13348 (N_13348,N_13074,N_13109);
and U13349 (N_13349,N_13087,N_13102);
or U13350 (N_13350,N_13130,N_13192);
nand U13351 (N_13351,N_13082,N_13193);
or U13352 (N_13352,N_13078,N_13066);
nor U13353 (N_13353,N_13195,N_13167);
xnor U13354 (N_13354,N_13111,N_13090);
nor U13355 (N_13355,N_13067,N_13003);
nand U13356 (N_13356,N_13049,N_13154);
or U13357 (N_13357,N_13042,N_13156);
or U13358 (N_13358,N_13156,N_13075);
nor U13359 (N_13359,N_13063,N_13178);
xnor U13360 (N_13360,N_13102,N_13017);
or U13361 (N_13361,N_13027,N_13197);
nand U13362 (N_13362,N_13016,N_13021);
xnor U13363 (N_13363,N_13115,N_13116);
xor U13364 (N_13364,N_13061,N_13040);
or U13365 (N_13365,N_13186,N_13038);
xnor U13366 (N_13366,N_13023,N_13176);
nor U13367 (N_13367,N_13153,N_13123);
or U13368 (N_13368,N_13037,N_13148);
xnor U13369 (N_13369,N_13049,N_13124);
or U13370 (N_13370,N_13068,N_13172);
nor U13371 (N_13371,N_13072,N_13088);
xnor U13372 (N_13372,N_13094,N_13163);
xor U13373 (N_13373,N_13052,N_13157);
and U13374 (N_13374,N_13194,N_13133);
nand U13375 (N_13375,N_13195,N_13026);
or U13376 (N_13376,N_13030,N_13113);
nand U13377 (N_13377,N_13137,N_13148);
and U13378 (N_13378,N_13146,N_13158);
xnor U13379 (N_13379,N_13079,N_13154);
nor U13380 (N_13380,N_13186,N_13132);
and U13381 (N_13381,N_13022,N_13165);
nor U13382 (N_13382,N_13166,N_13145);
or U13383 (N_13383,N_13177,N_13095);
nand U13384 (N_13384,N_13166,N_13057);
nor U13385 (N_13385,N_13017,N_13034);
nor U13386 (N_13386,N_13097,N_13135);
xnor U13387 (N_13387,N_13169,N_13004);
nor U13388 (N_13388,N_13139,N_13084);
nand U13389 (N_13389,N_13183,N_13196);
and U13390 (N_13390,N_13167,N_13157);
or U13391 (N_13391,N_13050,N_13036);
xnor U13392 (N_13392,N_13004,N_13015);
nor U13393 (N_13393,N_13174,N_13023);
and U13394 (N_13394,N_13065,N_13187);
xor U13395 (N_13395,N_13034,N_13131);
or U13396 (N_13396,N_13004,N_13093);
xnor U13397 (N_13397,N_13082,N_13124);
nor U13398 (N_13398,N_13128,N_13030);
or U13399 (N_13399,N_13044,N_13137);
nand U13400 (N_13400,N_13287,N_13212);
nand U13401 (N_13401,N_13293,N_13319);
nand U13402 (N_13402,N_13234,N_13239);
nand U13403 (N_13403,N_13269,N_13289);
and U13404 (N_13404,N_13205,N_13291);
nor U13405 (N_13405,N_13273,N_13245);
or U13406 (N_13406,N_13310,N_13301);
nor U13407 (N_13407,N_13224,N_13201);
and U13408 (N_13408,N_13252,N_13389);
and U13409 (N_13409,N_13267,N_13263);
xor U13410 (N_13410,N_13315,N_13371);
or U13411 (N_13411,N_13238,N_13312);
or U13412 (N_13412,N_13327,N_13272);
xor U13413 (N_13413,N_13334,N_13226);
nor U13414 (N_13414,N_13214,N_13206);
nand U13415 (N_13415,N_13352,N_13225);
nor U13416 (N_13416,N_13242,N_13229);
nand U13417 (N_13417,N_13391,N_13345);
or U13418 (N_13418,N_13298,N_13309);
xor U13419 (N_13419,N_13337,N_13221);
nor U13420 (N_13420,N_13326,N_13395);
xnor U13421 (N_13421,N_13207,N_13203);
or U13422 (N_13422,N_13220,N_13254);
nand U13423 (N_13423,N_13330,N_13368);
and U13424 (N_13424,N_13303,N_13204);
nand U13425 (N_13425,N_13347,N_13250);
or U13426 (N_13426,N_13283,N_13235);
nor U13427 (N_13427,N_13260,N_13359);
nor U13428 (N_13428,N_13350,N_13339);
and U13429 (N_13429,N_13280,N_13241);
nor U13430 (N_13430,N_13300,N_13304);
xnor U13431 (N_13431,N_13357,N_13286);
nand U13432 (N_13432,N_13213,N_13266);
xor U13433 (N_13433,N_13256,N_13227);
or U13434 (N_13434,N_13305,N_13349);
nand U13435 (N_13435,N_13222,N_13353);
xor U13436 (N_13436,N_13320,N_13306);
nor U13437 (N_13437,N_13248,N_13296);
nor U13438 (N_13438,N_13380,N_13323);
nand U13439 (N_13439,N_13228,N_13311);
and U13440 (N_13440,N_13277,N_13377);
nor U13441 (N_13441,N_13336,N_13346);
nand U13442 (N_13442,N_13322,N_13397);
xnor U13443 (N_13443,N_13384,N_13365);
nand U13444 (N_13444,N_13386,N_13216);
nor U13445 (N_13445,N_13247,N_13297);
nor U13446 (N_13446,N_13275,N_13262);
nand U13447 (N_13447,N_13215,N_13369);
and U13448 (N_13448,N_13351,N_13202);
nor U13449 (N_13449,N_13385,N_13344);
nor U13450 (N_13450,N_13370,N_13209);
xor U13451 (N_13451,N_13268,N_13328);
and U13452 (N_13452,N_13278,N_13233);
and U13453 (N_13453,N_13302,N_13210);
nor U13454 (N_13454,N_13294,N_13279);
nor U13455 (N_13455,N_13374,N_13246);
xnor U13456 (N_13456,N_13354,N_13276);
nor U13457 (N_13457,N_13265,N_13363);
xor U13458 (N_13458,N_13362,N_13398);
and U13459 (N_13459,N_13223,N_13316);
nor U13460 (N_13460,N_13387,N_13390);
and U13461 (N_13461,N_13360,N_13366);
or U13462 (N_13462,N_13314,N_13299);
and U13463 (N_13463,N_13394,N_13324);
xor U13464 (N_13464,N_13393,N_13274);
or U13465 (N_13465,N_13378,N_13249);
or U13466 (N_13466,N_13329,N_13392);
xnor U13467 (N_13467,N_13240,N_13376);
xor U13468 (N_13468,N_13264,N_13208);
or U13469 (N_13469,N_13243,N_13230);
xor U13470 (N_13470,N_13355,N_13321);
nand U13471 (N_13471,N_13341,N_13271);
nand U13472 (N_13472,N_13335,N_13281);
xnor U13473 (N_13473,N_13259,N_13258);
or U13474 (N_13474,N_13307,N_13325);
xor U13475 (N_13475,N_13382,N_13340);
xnor U13476 (N_13476,N_13285,N_13218);
xor U13477 (N_13477,N_13373,N_13217);
nor U13478 (N_13478,N_13290,N_13270);
nor U13479 (N_13479,N_13211,N_13343);
or U13480 (N_13480,N_13348,N_13284);
or U13481 (N_13481,N_13379,N_13383);
nand U13482 (N_13482,N_13372,N_13253);
and U13483 (N_13483,N_13381,N_13338);
nand U13484 (N_13484,N_13333,N_13282);
or U13485 (N_13485,N_13237,N_13388);
or U13486 (N_13486,N_13356,N_13396);
xnor U13487 (N_13487,N_13399,N_13288);
xnor U13488 (N_13488,N_13295,N_13317);
xnor U13489 (N_13489,N_13308,N_13367);
and U13490 (N_13490,N_13236,N_13361);
xor U13491 (N_13491,N_13364,N_13261);
nand U13492 (N_13492,N_13231,N_13292);
nand U13493 (N_13493,N_13200,N_13251);
xor U13494 (N_13494,N_13332,N_13342);
and U13495 (N_13495,N_13255,N_13244);
xor U13496 (N_13496,N_13313,N_13375);
xor U13497 (N_13497,N_13219,N_13358);
nor U13498 (N_13498,N_13232,N_13257);
nand U13499 (N_13499,N_13318,N_13331);
nand U13500 (N_13500,N_13304,N_13251);
xnor U13501 (N_13501,N_13293,N_13374);
or U13502 (N_13502,N_13398,N_13259);
and U13503 (N_13503,N_13215,N_13308);
and U13504 (N_13504,N_13351,N_13377);
or U13505 (N_13505,N_13270,N_13300);
or U13506 (N_13506,N_13346,N_13355);
nand U13507 (N_13507,N_13378,N_13266);
and U13508 (N_13508,N_13389,N_13394);
nor U13509 (N_13509,N_13218,N_13317);
xor U13510 (N_13510,N_13236,N_13258);
nand U13511 (N_13511,N_13226,N_13252);
nor U13512 (N_13512,N_13229,N_13332);
xnor U13513 (N_13513,N_13399,N_13270);
or U13514 (N_13514,N_13350,N_13384);
nand U13515 (N_13515,N_13237,N_13250);
nand U13516 (N_13516,N_13300,N_13234);
and U13517 (N_13517,N_13207,N_13267);
or U13518 (N_13518,N_13378,N_13343);
nor U13519 (N_13519,N_13290,N_13220);
nor U13520 (N_13520,N_13325,N_13203);
nor U13521 (N_13521,N_13384,N_13338);
and U13522 (N_13522,N_13359,N_13269);
xor U13523 (N_13523,N_13261,N_13265);
and U13524 (N_13524,N_13280,N_13398);
nor U13525 (N_13525,N_13362,N_13205);
or U13526 (N_13526,N_13210,N_13203);
nor U13527 (N_13527,N_13382,N_13392);
or U13528 (N_13528,N_13284,N_13208);
nand U13529 (N_13529,N_13338,N_13228);
nand U13530 (N_13530,N_13267,N_13292);
nand U13531 (N_13531,N_13392,N_13376);
nand U13532 (N_13532,N_13329,N_13254);
or U13533 (N_13533,N_13246,N_13292);
nand U13534 (N_13534,N_13387,N_13284);
nor U13535 (N_13535,N_13260,N_13274);
or U13536 (N_13536,N_13240,N_13242);
xor U13537 (N_13537,N_13324,N_13310);
nor U13538 (N_13538,N_13227,N_13367);
xnor U13539 (N_13539,N_13370,N_13386);
nand U13540 (N_13540,N_13378,N_13369);
nand U13541 (N_13541,N_13210,N_13238);
and U13542 (N_13542,N_13336,N_13397);
nor U13543 (N_13543,N_13397,N_13396);
nor U13544 (N_13544,N_13340,N_13385);
and U13545 (N_13545,N_13272,N_13239);
nand U13546 (N_13546,N_13204,N_13391);
nor U13547 (N_13547,N_13272,N_13281);
and U13548 (N_13548,N_13243,N_13200);
and U13549 (N_13549,N_13334,N_13386);
and U13550 (N_13550,N_13216,N_13297);
and U13551 (N_13551,N_13343,N_13296);
xor U13552 (N_13552,N_13291,N_13370);
or U13553 (N_13553,N_13311,N_13249);
xor U13554 (N_13554,N_13304,N_13221);
and U13555 (N_13555,N_13312,N_13326);
nor U13556 (N_13556,N_13219,N_13389);
and U13557 (N_13557,N_13237,N_13310);
nand U13558 (N_13558,N_13257,N_13373);
and U13559 (N_13559,N_13286,N_13340);
xnor U13560 (N_13560,N_13356,N_13265);
nor U13561 (N_13561,N_13313,N_13206);
and U13562 (N_13562,N_13311,N_13355);
xnor U13563 (N_13563,N_13245,N_13393);
or U13564 (N_13564,N_13341,N_13225);
nand U13565 (N_13565,N_13334,N_13370);
or U13566 (N_13566,N_13371,N_13242);
xnor U13567 (N_13567,N_13334,N_13248);
or U13568 (N_13568,N_13297,N_13398);
nor U13569 (N_13569,N_13344,N_13228);
nor U13570 (N_13570,N_13284,N_13361);
or U13571 (N_13571,N_13245,N_13227);
nand U13572 (N_13572,N_13284,N_13382);
xor U13573 (N_13573,N_13389,N_13233);
xnor U13574 (N_13574,N_13360,N_13327);
nor U13575 (N_13575,N_13321,N_13361);
nor U13576 (N_13576,N_13368,N_13399);
and U13577 (N_13577,N_13268,N_13289);
xor U13578 (N_13578,N_13364,N_13311);
nand U13579 (N_13579,N_13385,N_13257);
nor U13580 (N_13580,N_13332,N_13324);
and U13581 (N_13581,N_13220,N_13278);
nand U13582 (N_13582,N_13306,N_13270);
or U13583 (N_13583,N_13243,N_13238);
or U13584 (N_13584,N_13265,N_13274);
and U13585 (N_13585,N_13301,N_13217);
nand U13586 (N_13586,N_13273,N_13332);
or U13587 (N_13587,N_13298,N_13280);
or U13588 (N_13588,N_13216,N_13384);
nand U13589 (N_13589,N_13301,N_13258);
or U13590 (N_13590,N_13331,N_13291);
and U13591 (N_13591,N_13321,N_13278);
and U13592 (N_13592,N_13340,N_13368);
and U13593 (N_13593,N_13349,N_13234);
xor U13594 (N_13594,N_13273,N_13275);
xnor U13595 (N_13595,N_13258,N_13216);
xnor U13596 (N_13596,N_13342,N_13350);
nor U13597 (N_13597,N_13381,N_13388);
nor U13598 (N_13598,N_13283,N_13373);
and U13599 (N_13599,N_13223,N_13280);
or U13600 (N_13600,N_13501,N_13426);
xor U13601 (N_13601,N_13489,N_13532);
xor U13602 (N_13602,N_13575,N_13549);
or U13603 (N_13603,N_13599,N_13416);
and U13604 (N_13604,N_13476,N_13591);
nand U13605 (N_13605,N_13477,N_13504);
nor U13606 (N_13606,N_13482,N_13540);
nor U13607 (N_13607,N_13487,N_13514);
nand U13608 (N_13608,N_13497,N_13502);
or U13609 (N_13609,N_13475,N_13560);
or U13610 (N_13610,N_13576,N_13467);
or U13611 (N_13611,N_13592,N_13431);
or U13612 (N_13612,N_13574,N_13438);
xnor U13613 (N_13613,N_13568,N_13400);
xnor U13614 (N_13614,N_13542,N_13493);
nand U13615 (N_13615,N_13562,N_13443);
xnor U13616 (N_13616,N_13509,N_13454);
nor U13617 (N_13617,N_13480,N_13544);
nor U13618 (N_13618,N_13516,N_13458);
nand U13619 (N_13619,N_13447,N_13573);
or U13620 (N_13620,N_13495,N_13596);
nor U13621 (N_13621,N_13558,N_13430);
xnor U13622 (N_13622,N_13541,N_13524);
and U13623 (N_13623,N_13427,N_13584);
nand U13624 (N_13624,N_13408,N_13434);
nand U13625 (N_13625,N_13419,N_13435);
nand U13626 (N_13626,N_13450,N_13571);
and U13627 (N_13627,N_13559,N_13554);
xor U13628 (N_13628,N_13413,N_13572);
and U13629 (N_13629,N_13452,N_13404);
and U13630 (N_13630,N_13507,N_13481);
or U13631 (N_13631,N_13453,N_13553);
and U13632 (N_13632,N_13456,N_13582);
or U13633 (N_13633,N_13531,N_13439);
xnor U13634 (N_13634,N_13445,N_13523);
nand U13635 (N_13635,N_13498,N_13536);
nand U13636 (N_13636,N_13521,N_13513);
nor U13637 (N_13637,N_13520,N_13537);
xor U13638 (N_13638,N_13593,N_13579);
and U13639 (N_13639,N_13551,N_13429);
nor U13640 (N_13640,N_13457,N_13423);
nor U13641 (N_13641,N_13566,N_13422);
and U13642 (N_13642,N_13526,N_13484);
nand U13643 (N_13643,N_13570,N_13449);
nand U13644 (N_13644,N_13417,N_13412);
xor U13645 (N_13645,N_13451,N_13471);
nor U13646 (N_13646,N_13403,N_13527);
or U13647 (N_13647,N_13469,N_13444);
and U13648 (N_13648,N_13539,N_13468);
xor U13649 (N_13649,N_13581,N_13496);
xnor U13650 (N_13650,N_13485,N_13410);
or U13651 (N_13651,N_13577,N_13595);
and U13652 (N_13652,N_13500,N_13561);
or U13653 (N_13653,N_13491,N_13428);
and U13654 (N_13654,N_13519,N_13545);
and U13655 (N_13655,N_13508,N_13486);
and U13656 (N_13656,N_13437,N_13550);
nand U13657 (N_13657,N_13406,N_13483);
nor U13658 (N_13658,N_13518,N_13436);
nor U13659 (N_13659,N_13563,N_13465);
and U13660 (N_13660,N_13478,N_13505);
and U13661 (N_13661,N_13580,N_13440);
and U13662 (N_13662,N_13474,N_13548);
nor U13663 (N_13663,N_13512,N_13506);
xor U13664 (N_13664,N_13587,N_13511);
or U13665 (N_13665,N_13555,N_13473);
nor U13666 (N_13666,N_13578,N_13530);
nor U13667 (N_13667,N_13499,N_13488);
or U13668 (N_13668,N_13425,N_13433);
nor U13669 (N_13669,N_13462,N_13589);
xor U13670 (N_13670,N_13586,N_13535);
and U13671 (N_13671,N_13466,N_13522);
nor U13672 (N_13672,N_13598,N_13533);
xnor U13673 (N_13673,N_13597,N_13588);
xor U13674 (N_13674,N_13441,N_13552);
xnor U13675 (N_13675,N_13464,N_13546);
or U13676 (N_13676,N_13564,N_13414);
and U13677 (N_13677,N_13503,N_13494);
and U13678 (N_13678,N_13448,N_13432);
nor U13679 (N_13679,N_13407,N_13569);
nand U13680 (N_13680,N_13547,N_13567);
xor U13681 (N_13681,N_13517,N_13415);
or U13682 (N_13682,N_13583,N_13461);
nor U13683 (N_13683,N_13529,N_13565);
nand U13684 (N_13684,N_13515,N_13421);
xnor U13685 (N_13685,N_13402,N_13460);
xnor U13686 (N_13686,N_13446,N_13472);
and U13687 (N_13687,N_13442,N_13411);
xnor U13688 (N_13688,N_13538,N_13528);
or U13689 (N_13689,N_13525,N_13463);
or U13690 (N_13690,N_13492,N_13510);
and U13691 (N_13691,N_13401,N_13418);
or U13692 (N_13692,N_13556,N_13543);
xor U13693 (N_13693,N_13590,N_13479);
nor U13694 (N_13694,N_13470,N_13490);
xnor U13695 (N_13695,N_13557,N_13409);
xnor U13696 (N_13696,N_13455,N_13534);
xor U13697 (N_13697,N_13420,N_13594);
and U13698 (N_13698,N_13405,N_13459);
xnor U13699 (N_13699,N_13424,N_13585);
nor U13700 (N_13700,N_13409,N_13524);
nor U13701 (N_13701,N_13544,N_13479);
nand U13702 (N_13702,N_13531,N_13448);
or U13703 (N_13703,N_13563,N_13523);
nand U13704 (N_13704,N_13495,N_13566);
or U13705 (N_13705,N_13574,N_13476);
or U13706 (N_13706,N_13560,N_13493);
nor U13707 (N_13707,N_13470,N_13564);
xnor U13708 (N_13708,N_13543,N_13520);
nand U13709 (N_13709,N_13587,N_13524);
xnor U13710 (N_13710,N_13585,N_13584);
nor U13711 (N_13711,N_13416,N_13407);
nand U13712 (N_13712,N_13498,N_13590);
xor U13713 (N_13713,N_13543,N_13539);
or U13714 (N_13714,N_13401,N_13519);
xor U13715 (N_13715,N_13568,N_13472);
and U13716 (N_13716,N_13551,N_13467);
xnor U13717 (N_13717,N_13529,N_13593);
or U13718 (N_13718,N_13591,N_13441);
xor U13719 (N_13719,N_13500,N_13469);
and U13720 (N_13720,N_13521,N_13406);
xnor U13721 (N_13721,N_13565,N_13560);
xnor U13722 (N_13722,N_13462,N_13492);
nor U13723 (N_13723,N_13519,N_13466);
or U13724 (N_13724,N_13572,N_13576);
and U13725 (N_13725,N_13469,N_13545);
or U13726 (N_13726,N_13589,N_13425);
xor U13727 (N_13727,N_13535,N_13406);
or U13728 (N_13728,N_13571,N_13499);
xnor U13729 (N_13729,N_13452,N_13523);
nor U13730 (N_13730,N_13422,N_13501);
nor U13731 (N_13731,N_13582,N_13423);
nor U13732 (N_13732,N_13540,N_13537);
xnor U13733 (N_13733,N_13598,N_13465);
nand U13734 (N_13734,N_13562,N_13425);
and U13735 (N_13735,N_13464,N_13592);
and U13736 (N_13736,N_13415,N_13418);
nor U13737 (N_13737,N_13508,N_13595);
or U13738 (N_13738,N_13536,N_13410);
or U13739 (N_13739,N_13402,N_13436);
nor U13740 (N_13740,N_13428,N_13485);
nor U13741 (N_13741,N_13592,N_13525);
nor U13742 (N_13742,N_13546,N_13593);
nor U13743 (N_13743,N_13519,N_13428);
or U13744 (N_13744,N_13544,N_13539);
and U13745 (N_13745,N_13432,N_13417);
nor U13746 (N_13746,N_13486,N_13403);
xnor U13747 (N_13747,N_13596,N_13567);
xnor U13748 (N_13748,N_13540,N_13571);
xnor U13749 (N_13749,N_13464,N_13420);
nor U13750 (N_13750,N_13430,N_13496);
nand U13751 (N_13751,N_13482,N_13534);
nand U13752 (N_13752,N_13516,N_13525);
or U13753 (N_13753,N_13532,N_13475);
and U13754 (N_13754,N_13589,N_13554);
and U13755 (N_13755,N_13402,N_13452);
or U13756 (N_13756,N_13535,N_13480);
nor U13757 (N_13757,N_13511,N_13581);
or U13758 (N_13758,N_13507,N_13570);
xnor U13759 (N_13759,N_13536,N_13435);
nand U13760 (N_13760,N_13561,N_13592);
or U13761 (N_13761,N_13511,N_13413);
nand U13762 (N_13762,N_13462,N_13596);
xor U13763 (N_13763,N_13480,N_13583);
or U13764 (N_13764,N_13519,N_13437);
or U13765 (N_13765,N_13416,N_13481);
or U13766 (N_13766,N_13548,N_13402);
or U13767 (N_13767,N_13405,N_13569);
nand U13768 (N_13768,N_13533,N_13528);
or U13769 (N_13769,N_13451,N_13560);
and U13770 (N_13770,N_13403,N_13532);
nor U13771 (N_13771,N_13475,N_13434);
or U13772 (N_13772,N_13563,N_13586);
or U13773 (N_13773,N_13581,N_13557);
nor U13774 (N_13774,N_13484,N_13548);
and U13775 (N_13775,N_13589,N_13486);
nor U13776 (N_13776,N_13542,N_13436);
nand U13777 (N_13777,N_13551,N_13556);
nand U13778 (N_13778,N_13580,N_13538);
or U13779 (N_13779,N_13443,N_13469);
nand U13780 (N_13780,N_13471,N_13492);
xor U13781 (N_13781,N_13500,N_13550);
or U13782 (N_13782,N_13538,N_13471);
nor U13783 (N_13783,N_13481,N_13411);
or U13784 (N_13784,N_13591,N_13551);
nand U13785 (N_13785,N_13595,N_13449);
or U13786 (N_13786,N_13428,N_13526);
nor U13787 (N_13787,N_13542,N_13461);
nand U13788 (N_13788,N_13489,N_13496);
nor U13789 (N_13789,N_13453,N_13551);
or U13790 (N_13790,N_13578,N_13596);
nand U13791 (N_13791,N_13425,N_13444);
nand U13792 (N_13792,N_13579,N_13471);
and U13793 (N_13793,N_13496,N_13557);
nand U13794 (N_13794,N_13559,N_13542);
nor U13795 (N_13795,N_13517,N_13441);
xor U13796 (N_13796,N_13538,N_13446);
nand U13797 (N_13797,N_13538,N_13505);
and U13798 (N_13798,N_13457,N_13468);
nand U13799 (N_13799,N_13428,N_13520);
nor U13800 (N_13800,N_13783,N_13715);
nand U13801 (N_13801,N_13714,N_13725);
nor U13802 (N_13802,N_13786,N_13704);
nand U13803 (N_13803,N_13627,N_13709);
nand U13804 (N_13804,N_13609,N_13700);
xnor U13805 (N_13805,N_13773,N_13647);
and U13806 (N_13806,N_13744,N_13658);
and U13807 (N_13807,N_13677,N_13689);
nand U13808 (N_13808,N_13799,N_13784);
and U13809 (N_13809,N_13612,N_13674);
nand U13810 (N_13810,N_13630,N_13743);
and U13811 (N_13811,N_13777,N_13653);
and U13812 (N_13812,N_13641,N_13602);
and U13813 (N_13813,N_13755,N_13718);
xnor U13814 (N_13814,N_13633,N_13672);
nor U13815 (N_13815,N_13617,N_13679);
or U13816 (N_13816,N_13606,N_13635);
and U13817 (N_13817,N_13705,N_13615);
nor U13818 (N_13818,N_13798,N_13662);
or U13819 (N_13819,N_13703,N_13789);
and U13820 (N_13820,N_13797,N_13735);
xor U13821 (N_13821,N_13697,N_13721);
and U13822 (N_13822,N_13708,N_13754);
xnor U13823 (N_13823,N_13681,N_13608);
and U13824 (N_13824,N_13722,N_13655);
or U13825 (N_13825,N_13753,N_13650);
or U13826 (N_13826,N_13739,N_13688);
nor U13827 (N_13827,N_13699,N_13669);
nand U13828 (N_13828,N_13770,N_13769);
nor U13829 (N_13829,N_13775,N_13696);
and U13830 (N_13830,N_13724,N_13774);
or U13831 (N_13831,N_13778,N_13643);
xor U13832 (N_13832,N_13772,N_13684);
nand U13833 (N_13833,N_13741,N_13651);
nor U13834 (N_13834,N_13748,N_13624);
xnor U13835 (N_13835,N_13657,N_13761);
and U13836 (N_13836,N_13678,N_13629);
nand U13837 (N_13837,N_13675,N_13791);
nand U13838 (N_13838,N_13640,N_13713);
and U13839 (N_13839,N_13636,N_13654);
or U13840 (N_13840,N_13690,N_13613);
nand U13841 (N_13841,N_13779,N_13719);
nand U13842 (N_13842,N_13746,N_13680);
and U13843 (N_13843,N_13623,N_13666);
xor U13844 (N_13844,N_13659,N_13692);
xor U13845 (N_13845,N_13733,N_13625);
xor U13846 (N_13846,N_13691,N_13747);
nand U13847 (N_13847,N_13729,N_13790);
nor U13848 (N_13848,N_13607,N_13736);
or U13849 (N_13849,N_13695,N_13610);
or U13850 (N_13850,N_13781,N_13734);
nor U13851 (N_13851,N_13639,N_13792);
and U13852 (N_13852,N_13620,N_13614);
and U13853 (N_13853,N_13767,N_13710);
and U13854 (N_13854,N_13600,N_13687);
nand U13855 (N_13855,N_13782,N_13634);
nor U13856 (N_13856,N_13619,N_13763);
and U13857 (N_13857,N_13707,N_13771);
and U13858 (N_13858,N_13702,N_13706);
nand U13859 (N_13859,N_13665,N_13693);
xnor U13860 (N_13860,N_13622,N_13765);
nor U13861 (N_13861,N_13757,N_13793);
xnor U13862 (N_13862,N_13618,N_13723);
nand U13863 (N_13863,N_13712,N_13732);
and U13864 (N_13864,N_13728,N_13648);
xnor U13865 (N_13865,N_13738,N_13605);
or U13866 (N_13866,N_13780,N_13694);
xnor U13867 (N_13867,N_13676,N_13628);
nor U13868 (N_13868,N_13751,N_13632);
or U13869 (N_13869,N_13698,N_13768);
nand U13870 (N_13870,N_13720,N_13776);
nand U13871 (N_13871,N_13711,N_13762);
nor U13872 (N_13872,N_13626,N_13758);
nor U13873 (N_13873,N_13701,N_13742);
xor U13874 (N_13874,N_13656,N_13631);
xnor U13875 (N_13875,N_13785,N_13759);
nor U13876 (N_13876,N_13717,N_13664);
or U13877 (N_13877,N_13740,N_13730);
or U13878 (N_13878,N_13660,N_13644);
and U13879 (N_13879,N_13787,N_13737);
nand U13880 (N_13880,N_13603,N_13621);
nor U13881 (N_13881,N_13745,N_13727);
and U13882 (N_13882,N_13649,N_13716);
and U13883 (N_13883,N_13685,N_13670);
and U13884 (N_13884,N_13642,N_13752);
and U13885 (N_13885,N_13686,N_13749);
nand U13886 (N_13886,N_13663,N_13788);
and U13887 (N_13887,N_13760,N_13604);
or U13888 (N_13888,N_13637,N_13726);
and U13889 (N_13889,N_13756,N_13794);
and U13890 (N_13890,N_13673,N_13671);
and U13891 (N_13891,N_13683,N_13682);
and U13892 (N_13892,N_13731,N_13661);
nor U13893 (N_13893,N_13764,N_13795);
nand U13894 (N_13894,N_13667,N_13616);
nand U13895 (N_13895,N_13766,N_13750);
xnor U13896 (N_13896,N_13652,N_13645);
xor U13897 (N_13897,N_13601,N_13796);
and U13898 (N_13898,N_13668,N_13611);
nand U13899 (N_13899,N_13646,N_13638);
and U13900 (N_13900,N_13609,N_13626);
xnor U13901 (N_13901,N_13692,N_13740);
xor U13902 (N_13902,N_13684,N_13658);
nand U13903 (N_13903,N_13782,N_13695);
xor U13904 (N_13904,N_13641,N_13674);
xor U13905 (N_13905,N_13621,N_13676);
nor U13906 (N_13906,N_13664,N_13734);
xnor U13907 (N_13907,N_13772,N_13798);
nor U13908 (N_13908,N_13614,N_13738);
xnor U13909 (N_13909,N_13722,N_13665);
and U13910 (N_13910,N_13669,N_13799);
nor U13911 (N_13911,N_13716,N_13715);
and U13912 (N_13912,N_13763,N_13622);
nand U13913 (N_13913,N_13732,N_13759);
xnor U13914 (N_13914,N_13753,N_13787);
or U13915 (N_13915,N_13676,N_13745);
and U13916 (N_13916,N_13762,N_13676);
nand U13917 (N_13917,N_13632,N_13648);
xnor U13918 (N_13918,N_13651,N_13700);
and U13919 (N_13919,N_13719,N_13646);
nor U13920 (N_13920,N_13770,N_13785);
xnor U13921 (N_13921,N_13782,N_13781);
and U13922 (N_13922,N_13638,N_13705);
and U13923 (N_13923,N_13734,N_13793);
nor U13924 (N_13924,N_13606,N_13603);
xor U13925 (N_13925,N_13700,N_13755);
xnor U13926 (N_13926,N_13616,N_13737);
and U13927 (N_13927,N_13784,N_13709);
or U13928 (N_13928,N_13764,N_13674);
xor U13929 (N_13929,N_13771,N_13774);
or U13930 (N_13930,N_13685,N_13692);
or U13931 (N_13931,N_13682,N_13684);
nor U13932 (N_13932,N_13638,N_13684);
or U13933 (N_13933,N_13718,N_13782);
nand U13934 (N_13934,N_13713,N_13740);
xnor U13935 (N_13935,N_13782,N_13780);
or U13936 (N_13936,N_13723,N_13691);
or U13937 (N_13937,N_13737,N_13772);
nand U13938 (N_13938,N_13692,N_13739);
xor U13939 (N_13939,N_13745,N_13686);
nor U13940 (N_13940,N_13691,N_13752);
or U13941 (N_13941,N_13704,N_13602);
xnor U13942 (N_13942,N_13671,N_13714);
and U13943 (N_13943,N_13788,N_13692);
and U13944 (N_13944,N_13798,N_13694);
xor U13945 (N_13945,N_13729,N_13675);
and U13946 (N_13946,N_13621,N_13785);
nor U13947 (N_13947,N_13648,N_13601);
and U13948 (N_13948,N_13731,N_13714);
or U13949 (N_13949,N_13737,N_13742);
nand U13950 (N_13950,N_13722,N_13642);
or U13951 (N_13951,N_13787,N_13769);
nor U13952 (N_13952,N_13757,N_13762);
nor U13953 (N_13953,N_13795,N_13705);
or U13954 (N_13954,N_13661,N_13616);
nand U13955 (N_13955,N_13738,N_13700);
or U13956 (N_13956,N_13752,N_13744);
nand U13957 (N_13957,N_13695,N_13707);
and U13958 (N_13958,N_13736,N_13649);
nor U13959 (N_13959,N_13623,N_13653);
and U13960 (N_13960,N_13612,N_13739);
nor U13961 (N_13961,N_13779,N_13601);
nand U13962 (N_13962,N_13773,N_13629);
or U13963 (N_13963,N_13652,N_13666);
or U13964 (N_13964,N_13608,N_13719);
nand U13965 (N_13965,N_13628,N_13660);
nor U13966 (N_13966,N_13669,N_13793);
or U13967 (N_13967,N_13729,N_13617);
or U13968 (N_13968,N_13742,N_13723);
nand U13969 (N_13969,N_13608,N_13676);
xnor U13970 (N_13970,N_13684,N_13612);
nor U13971 (N_13971,N_13654,N_13682);
and U13972 (N_13972,N_13739,N_13793);
nor U13973 (N_13973,N_13732,N_13791);
xor U13974 (N_13974,N_13659,N_13741);
or U13975 (N_13975,N_13707,N_13734);
xor U13976 (N_13976,N_13776,N_13651);
or U13977 (N_13977,N_13702,N_13763);
nor U13978 (N_13978,N_13778,N_13716);
nor U13979 (N_13979,N_13704,N_13723);
and U13980 (N_13980,N_13600,N_13725);
or U13981 (N_13981,N_13609,N_13614);
or U13982 (N_13982,N_13630,N_13737);
or U13983 (N_13983,N_13794,N_13686);
and U13984 (N_13984,N_13638,N_13778);
nand U13985 (N_13985,N_13710,N_13713);
and U13986 (N_13986,N_13716,N_13679);
and U13987 (N_13987,N_13771,N_13716);
xor U13988 (N_13988,N_13762,N_13778);
xnor U13989 (N_13989,N_13616,N_13708);
xor U13990 (N_13990,N_13788,N_13733);
or U13991 (N_13991,N_13612,N_13628);
and U13992 (N_13992,N_13701,N_13679);
nor U13993 (N_13993,N_13739,N_13776);
and U13994 (N_13994,N_13799,N_13617);
or U13995 (N_13995,N_13794,N_13788);
or U13996 (N_13996,N_13615,N_13712);
nand U13997 (N_13997,N_13610,N_13631);
nor U13998 (N_13998,N_13768,N_13726);
xor U13999 (N_13999,N_13629,N_13762);
nand U14000 (N_14000,N_13877,N_13964);
xor U14001 (N_14001,N_13885,N_13898);
and U14002 (N_14002,N_13848,N_13982);
and U14003 (N_14003,N_13908,N_13858);
and U14004 (N_14004,N_13840,N_13828);
nand U14005 (N_14005,N_13892,N_13865);
nand U14006 (N_14006,N_13862,N_13850);
nor U14007 (N_14007,N_13953,N_13811);
or U14008 (N_14008,N_13956,N_13866);
nand U14009 (N_14009,N_13932,N_13938);
and U14010 (N_14010,N_13921,N_13965);
nor U14011 (N_14011,N_13802,N_13816);
nor U14012 (N_14012,N_13970,N_13920);
xnor U14013 (N_14013,N_13940,N_13824);
xor U14014 (N_14014,N_13882,N_13957);
and U14015 (N_14015,N_13911,N_13826);
and U14016 (N_14016,N_13926,N_13919);
and U14017 (N_14017,N_13918,N_13827);
or U14018 (N_14018,N_13843,N_13894);
xnor U14019 (N_14019,N_13949,N_13975);
nand U14020 (N_14020,N_13896,N_13805);
nand U14021 (N_14021,N_13913,N_13856);
nor U14022 (N_14022,N_13985,N_13886);
or U14023 (N_14023,N_13814,N_13976);
nor U14024 (N_14024,N_13854,N_13928);
nor U14025 (N_14025,N_13933,N_13984);
and U14026 (N_14026,N_13838,N_13948);
or U14027 (N_14027,N_13813,N_13800);
and U14028 (N_14028,N_13845,N_13951);
or U14029 (N_14029,N_13869,N_13804);
xnor U14030 (N_14030,N_13995,N_13925);
xor U14031 (N_14031,N_13914,N_13966);
and U14032 (N_14032,N_13955,N_13842);
nor U14033 (N_14033,N_13884,N_13971);
xnor U14034 (N_14034,N_13815,N_13998);
and U14035 (N_14035,N_13929,N_13943);
or U14036 (N_14036,N_13855,N_13915);
nor U14037 (N_14037,N_13830,N_13988);
and U14038 (N_14038,N_13857,N_13909);
and U14039 (N_14039,N_13907,N_13962);
or U14040 (N_14040,N_13978,N_13991);
and U14041 (N_14041,N_13963,N_13844);
xor U14042 (N_14042,N_13801,N_13979);
nand U14043 (N_14043,N_13903,N_13968);
nand U14044 (N_14044,N_13952,N_13977);
and U14045 (N_14045,N_13859,N_13868);
and U14046 (N_14046,N_13846,N_13852);
and U14047 (N_14047,N_13883,N_13853);
or U14048 (N_14048,N_13829,N_13969);
nor U14049 (N_14049,N_13939,N_13992);
nand U14050 (N_14050,N_13916,N_13847);
and U14051 (N_14051,N_13950,N_13822);
and U14052 (N_14052,N_13861,N_13841);
nand U14053 (N_14053,N_13833,N_13931);
nand U14054 (N_14054,N_13936,N_13910);
or U14055 (N_14055,N_13806,N_13810);
xor U14056 (N_14056,N_13895,N_13961);
and U14057 (N_14057,N_13876,N_13818);
nor U14058 (N_14058,N_13820,N_13987);
nor U14059 (N_14059,N_13879,N_13942);
or U14060 (N_14060,N_13904,N_13867);
or U14061 (N_14061,N_13812,N_13807);
xnor U14062 (N_14062,N_13983,N_13905);
nand U14063 (N_14063,N_13878,N_13923);
nand U14064 (N_14064,N_13986,N_13873);
xnor U14065 (N_14065,N_13872,N_13817);
or U14066 (N_14066,N_13863,N_13870);
or U14067 (N_14067,N_13808,N_13990);
nand U14068 (N_14068,N_13941,N_13954);
nand U14069 (N_14069,N_13947,N_13906);
or U14070 (N_14070,N_13912,N_13851);
and U14071 (N_14071,N_13924,N_13831);
nand U14072 (N_14072,N_13881,N_13960);
nand U14073 (N_14073,N_13934,N_13945);
nor U14074 (N_14074,N_13821,N_13917);
nand U14075 (N_14075,N_13902,N_13997);
or U14076 (N_14076,N_13874,N_13922);
xnor U14077 (N_14077,N_13839,N_13819);
nor U14078 (N_14078,N_13888,N_13999);
nand U14079 (N_14079,N_13837,N_13849);
xnor U14080 (N_14080,N_13836,N_13823);
nand U14081 (N_14081,N_13893,N_13875);
and U14082 (N_14082,N_13871,N_13937);
nor U14083 (N_14083,N_13989,N_13900);
and U14084 (N_14084,N_13880,N_13946);
and U14085 (N_14085,N_13887,N_13930);
and U14086 (N_14086,N_13935,N_13891);
nor U14087 (N_14087,N_13944,N_13901);
nand U14088 (N_14088,N_13803,N_13994);
or U14089 (N_14089,N_13889,N_13897);
nor U14090 (N_14090,N_13835,N_13967);
xnor U14091 (N_14091,N_13959,N_13973);
and U14092 (N_14092,N_13981,N_13899);
xnor U14093 (N_14093,N_13974,N_13809);
nor U14094 (N_14094,N_13825,N_13996);
or U14095 (N_14095,N_13890,N_13972);
and U14096 (N_14096,N_13958,N_13864);
nor U14097 (N_14097,N_13834,N_13832);
nor U14098 (N_14098,N_13980,N_13993);
and U14099 (N_14099,N_13927,N_13860);
xor U14100 (N_14100,N_13821,N_13902);
and U14101 (N_14101,N_13984,N_13963);
nor U14102 (N_14102,N_13803,N_13901);
or U14103 (N_14103,N_13813,N_13836);
xor U14104 (N_14104,N_13998,N_13932);
xnor U14105 (N_14105,N_13806,N_13968);
and U14106 (N_14106,N_13946,N_13973);
nand U14107 (N_14107,N_13891,N_13813);
nor U14108 (N_14108,N_13898,N_13830);
or U14109 (N_14109,N_13822,N_13901);
and U14110 (N_14110,N_13856,N_13964);
xnor U14111 (N_14111,N_13843,N_13859);
nor U14112 (N_14112,N_13970,N_13899);
nor U14113 (N_14113,N_13933,N_13836);
or U14114 (N_14114,N_13857,N_13818);
nand U14115 (N_14115,N_13861,N_13899);
nand U14116 (N_14116,N_13932,N_13874);
xor U14117 (N_14117,N_13854,N_13899);
or U14118 (N_14118,N_13894,N_13953);
and U14119 (N_14119,N_13818,N_13971);
nor U14120 (N_14120,N_13984,N_13994);
nand U14121 (N_14121,N_13829,N_13955);
or U14122 (N_14122,N_13813,N_13966);
xnor U14123 (N_14123,N_13953,N_13849);
and U14124 (N_14124,N_13831,N_13972);
nor U14125 (N_14125,N_13819,N_13910);
and U14126 (N_14126,N_13831,N_13884);
or U14127 (N_14127,N_13829,N_13982);
and U14128 (N_14128,N_13832,N_13831);
nor U14129 (N_14129,N_13947,N_13830);
or U14130 (N_14130,N_13949,N_13989);
nor U14131 (N_14131,N_13881,N_13883);
xor U14132 (N_14132,N_13952,N_13999);
or U14133 (N_14133,N_13864,N_13954);
and U14134 (N_14134,N_13918,N_13967);
or U14135 (N_14135,N_13957,N_13877);
or U14136 (N_14136,N_13964,N_13816);
or U14137 (N_14137,N_13957,N_13804);
nand U14138 (N_14138,N_13848,N_13859);
nor U14139 (N_14139,N_13842,N_13981);
xnor U14140 (N_14140,N_13860,N_13888);
xnor U14141 (N_14141,N_13981,N_13995);
and U14142 (N_14142,N_13843,N_13912);
nor U14143 (N_14143,N_13881,N_13810);
xnor U14144 (N_14144,N_13929,N_13826);
and U14145 (N_14145,N_13816,N_13922);
and U14146 (N_14146,N_13869,N_13800);
and U14147 (N_14147,N_13834,N_13843);
nand U14148 (N_14148,N_13904,N_13884);
xor U14149 (N_14149,N_13959,N_13800);
nor U14150 (N_14150,N_13883,N_13819);
nor U14151 (N_14151,N_13862,N_13864);
xnor U14152 (N_14152,N_13866,N_13975);
and U14153 (N_14153,N_13959,N_13949);
nand U14154 (N_14154,N_13909,N_13842);
nand U14155 (N_14155,N_13965,N_13939);
xnor U14156 (N_14156,N_13998,N_13974);
and U14157 (N_14157,N_13950,N_13872);
or U14158 (N_14158,N_13860,N_13966);
nand U14159 (N_14159,N_13941,N_13833);
or U14160 (N_14160,N_13985,N_13930);
and U14161 (N_14161,N_13873,N_13851);
or U14162 (N_14162,N_13840,N_13862);
or U14163 (N_14163,N_13875,N_13838);
nor U14164 (N_14164,N_13822,N_13977);
xor U14165 (N_14165,N_13881,N_13973);
and U14166 (N_14166,N_13883,N_13919);
nand U14167 (N_14167,N_13867,N_13925);
nand U14168 (N_14168,N_13929,N_13880);
or U14169 (N_14169,N_13916,N_13956);
or U14170 (N_14170,N_13984,N_13810);
xnor U14171 (N_14171,N_13800,N_13935);
xnor U14172 (N_14172,N_13988,N_13811);
or U14173 (N_14173,N_13944,N_13860);
and U14174 (N_14174,N_13831,N_13825);
xnor U14175 (N_14175,N_13967,N_13825);
nor U14176 (N_14176,N_13812,N_13879);
and U14177 (N_14177,N_13829,N_13831);
xnor U14178 (N_14178,N_13931,N_13808);
nand U14179 (N_14179,N_13972,N_13973);
nand U14180 (N_14180,N_13830,N_13805);
nand U14181 (N_14181,N_13988,N_13823);
and U14182 (N_14182,N_13985,N_13870);
and U14183 (N_14183,N_13984,N_13986);
and U14184 (N_14184,N_13948,N_13872);
and U14185 (N_14185,N_13958,N_13917);
xor U14186 (N_14186,N_13952,N_13892);
or U14187 (N_14187,N_13884,N_13927);
or U14188 (N_14188,N_13843,N_13919);
and U14189 (N_14189,N_13958,N_13935);
or U14190 (N_14190,N_13922,N_13946);
and U14191 (N_14191,N_13824,N_13879);
nor U14192 (N_14192,N_13820,N_13977);
xnor U14193 (N_14193,N_13971,N_13951);
nor U14194 (N_14194,N_13925,N_13870);
or U14195 (N_14195,N_13801,N_13842);
and U14196 (N_14196,N_13930,N_13953);
nor U14197 (N_14197,N_13829,N_13812);
nor U14198 (N_14198,N_13928,N_13810);
nor U14199 (N_14199,N_13803,N_13969);
or U14200 (N_14200,N_14116,N_14041);
xnor U14201 (N_14201,N_14151,N_14000);
or U14202 (N_14202,N_14052,N_14001);
nor U14203 (N_14203,N_14112,N_14119);
or U14204 (N_14204,N_14020,N_14171);
xor U14205 (N_14205,N_14016,N_14071);
and U14206 (N_14206,N_14093,N_14197);
nand U14207 (N_14207,N_14135,N_14146);
nor U14208 (N_14208,N_14011,N_14130);
or U14209 (N_14209,N_14189,N_14094);
nor U14210 (N_14210,N_14057,N_14061);
nand U14211 (N_14211,N_14046,N_14034);
nor U14212 (N_14212,N_14168,N_14113);
nor U14213 (N_14213,N_14162,N_14107);
or U14214 (N_14214,N_14199,N_14062);
and U14215 (N_14215,N_14076,N_14184);
nor U14216 (N_14216,N_14147,N_14185);
nor U14217 (N_14217,N_14164,N_14152);
xnor U14218 (N_14218,N_14031,N_14072);
and U14219 (N_14219,N_14126,N_14095);
nand U14220 (N_14220,N_14121,N_14100);
nand U14221 (N_14221,N_14044,N_14170);
nand U14222 (N_14222,N_14102,N_14056);
nor U14223 (N_14223,N_14087,N_14086);
or U14224 (N_14224,N_14160,N_14172);
xnor U14225 (N_14225,N_14132,N_14081);
or U14226 (N_14226,N_14165,N_14192);
nand U14227 (N_14227,N_14048,N_14144);
and U14228 (N_14228,N_14058,N_14035);
or U14229 (N_14229,N_14090,N_14068);
xnor U14230 (N_14230,N_14045,N_14059);
xnor U14231 (N_14231,N_14036,N_14003);
nand U14232 (N_14232,N_14033,N_14064);
or U14233 (N_14233,N_14024,N_14115);
and U14234 (N_14234,N_14104,N_14149);
or U14235 (N_14235,N_14118,N_14133);
nand U14236 (N_14236,N_14155,N_14088);
nand U14237 (N_14237,N_14008,N_14142);
nor U14238 (N_14238,N_14021,N_14049);
nand U14239 (N_14239,N_14137,N_14140);
nor U14240 (N_14240,N_14109,N_14037);
and U14241 (N_14241,N_14099,N_14025);
xnor U14242 (N_14242,N_14191,N_14026);
nand U14243 (N_14243,N_14156,N_14154);
or U14244 (N_14244,N_14174,N_14131);
and U14245 (N_14245,N_14089,N_14120);
nand U14246 (N_14246,N_14158,N_14091);
or U14247 (N_14247,N_14069,N_14040);
nor U14248 (N_14248,N_14010,N_14009);
xor U14249 (N_14249,N_14176,N_14015);
nor U14250 (N_14250,N_14128,N_14006);
and U14251 (N_14251,N_14123,N_14080);
nand U14252 (N_14252,N_14043,N_14012);
nand U14253 (N_14253,N_14178,N_14007);
xor U14254 (N_14254,N_14042,N_14183);
xnor U14255 (N_14255,N_14098,N_14150);
nor U14256 (N_14256,N_14078,N_14047);
nor U14257 (N_14257,N_14194,N_14163);
nand U14258 (N_14258,N_14075,N_14103);
nor U14259 (N_14259,N_14055,N_14028);
or U14260 (N_14260,N_14084,N_14079);
nor U14261 (N_14261,N_14063,N_14114);
nor U14262 (N_14262,N_14129,N_14198);
xnor U14263 (N_14263,N_14054,N_14182);
nand U14264 (N_14264,N_14125,N_14097);
nor U14265 (N_14265,N_14005,N_14105);
xnor U14266 (N_14266,N_14193,N_14077);
and U14267 (N_14267,N_14085,N_14032);
xnor U14268 (N_14268,N_14067,N_14111);
nor U14269 (N_14269,N_14023,N_14179);
or U14270 (N_14270,N_14108,N_14141);
xor U14271 (N_14271,N_14074,N_14195);
nor U14272 (N_14272,N_14002,N_14188);
or U14273 (N_14273,N_14004,N_14180);
nor U14274 (N_14274,N_14019,N_14190);
nor U14275 (N_14275,N_14014,N_14017);
nor U14276 (N_14276,N_14117,N_14029);
nor U14277 (N_14277,N_14101,N_14138);
or U14278 (N_14278,N_14145,N_14039);
nand U14279 (N_14279,N_14073,N_14177);
nand U14280 (N_14280,N_14173,N_14122);
and U14281 (N_14281,N_14175,N_14092);
and U14282 (N_14282,N_14181,N_14110);
and U14283 (N_14283,N_14083,N_14127);
and U14284 (N_14284,N_14096,N_14169);
xnor U14285 (N_14285,N_14134,N_14161);
nand U14286 (N_14286,N_14065,N_14136);
nand U14287 (N_14287,N_14013,N_14027);
or U14288 (N_14288,N_14106,N_14060);
nor U14289 (N_14289,N_14066,N_14187);
xnor U14290 (N_14290,N_14143,N_14070);
and U14291 (N_14291,N_14186,N_14167);
nand U14292 (N_14292,N_14159,N_14196);
nand U14293 (N_14293,N_14166,N_14018);
and U14294 (N_14294,N_14038,N_14030);
xor U14295 (N_14295,N_14053,N_14022);
and U14296 (N_14296,N_14153,N_14157);
or U14297 (N_14297,N_14148,N_14082);
or U14298 (N_14298,N_14124,N_14139);
nand U14299 (N_14299,N_14050,N_14051);
nand U14300 (N_14300,N_14000,N_14026);
and U14301 (N_14301,N_14073,N_14067);
nor U14302 (N_14302,N_14029,N_14014);
and U14303 (N_14303,N_14014,N_14018);
nor U14304 (N_14304,N_14008,N_14063);
nand U14305 (N_14305,N_14199,N_14001);
nor U14306 (N_14306,N_14018,N_14026);
and U14307 (N_14307,N_14091,N_14031);
or U14308 (N_14308,N_14049,N_14176);
nor U14309 (N_14309,N_14060,N_14010);
nor U14310 (N_14310,N_14145,N_14169);
nand U14311 (N_14311,N_14180,N_14143);
or U14312 (N_14312,N_14130,N_14170);
nand U14313 (N_14313,N_14171,N_14042);
nand U14314 (N_14314,N_14127,N_14048);
xor U14315 (N_14315,N_14187,N_14197);
and U14316 (N_14316,N_14151,N_14164);
xor U14317 (N_14317,N_14082,N_14104);
xnor U14318 (N_14318,N_14064,N_14121);
xnor U14319 (N_14319,N_14009,N_14165);
nor U14320 (N_14320,N_14187,N_14059);
and U14321 (N_14321,N_14198,N_14162);
nor U14322 (N_14322,N_14024,N_14076);
or U14323 (N_14323,N_14089,N_14091);
xor U14324 (N_14324,N_14141,N_14037);
or U14325 (N_14325,N_14001,N_14057);
nor U14326 (N_14326,N_14181,N_14053);
or U14327 (N_14327,N_14089,N_14159);
nor U14328 (N_14328,N_14188,N_14025);
xor U14329 (N_14329,N_14143,N_14146);
or U14330 (N_14330,N_14149,N_14134);
xor U14331 (N_14331,N_14083,N_14153);
nor U14332 (N_14332,N_14174,N_14122);
or U14333 (N_14333,N_14153,N_14146);
xor U14334 (N_14334,N_14042,N_14079);
and U14335 (N_14335,N_14021,N_14113);
xor U14336 (N_14336,N_14176,N_14042);
xor U14337 (N_14337,N_14150,N_14186);
nand U14338 (N_14338,N_14083,N_14113);
and U14339 (N_14339,N_14165,N_14039);
nor U14340 (N_14340,N_14143,N_14184);
nor U14341 (N_14341,N_14088,N_14139);
nand U14342 (N_14342,N_14169,N_14062);
nand U14343 (N_14343,N_14062,N_14014);
nor U14344 (N_14344,N_14000,N_14019);
and U14345 (N_14345,N_14027,N_14116);
or U14346 (N_14346,N_14130,N_14083);
nor U14347 (N_14347,N_14142,N_14121);
nor U14348 (N_14348,N_14051,N_14177);
xor U14349 (N_14349,N_14066,N_14064);
nand U14350 (N_14350,N_14175,N_14181);
or U14351 (N_14351,N_14059,N_14049);
nand U14352 (N_14352,N_14192,N_14125);
nor U14353 (N_14353,N_14155,N_14038);
nor U14354 (N_14354,N_14073,N_14166);
and U14355 (N_14355,N_14173,N_14155);
and U14356 (N_14356,N_14169,N_14049);
or U14357 (N_14357,N_14076,N_14081);
and U14358 (N_14358,N_14078,N_14087);
or U14359 (N_14359,N_14186,N_14022);
and U14360 (N_14360,N_14143,N_14151);
nand U14361 (N_14361,N_14196,N_14078);
nor U14362 (N_14362,N_14027,N_14170);
nor U14363 (N_14363,N_14085,N_14178);
xor U14364 (N_14364,N_14183,N_14161);
xnor U14365 (N_14365,N_14088,N_14053);
nor U14366 (N_14366,N_14021,N_14133);
nor U14367 (N_14367,N_14090,N_14142);
nor U14368 (N_14368,N_14125,N_14069);
xnor U14369 (N_14369,N_14094,N_14118);
xnor U14370 (N_14370,N_14189,N_14069);
nand U14371 (N_14371,N_14115,N_14041);
nand U14372 (N_14372,N_14166,N_14078);
nand U14373 (N_14373,N_14007,N_14042);
and U14374 (N_14374,N_14105,N_14136);
or U14375 (N_14375,N_14093,N_14097);
and U14376 (N_14376,N_14133,N_14159);
nand U14377 (N_14377,N_14006,N_14125);
nor U14378 (N_14378,N_14183,N_14135);
nor U14379 (N_14379,N_14160,N_14032);
nor U14380 (N_14380,N_14122,N_14060);
xnor U14381 (N_14381,N_14157,N_14195);
or U14382 (N_14382,N_14004,N_14114);
nand U14383 (N_14383,N_14126,N_14061);
xnor U14384 (N_14384,N_14060,N_14146);
and U14385 (N_14385,N_14044,N_14072);
xnor U14386 (N_14386,N_14196,N_14118);
or U14387 (N_14387,N_14059,N_14012);
or U14388 (N_14388,N_14166,N_14170);
xnor U14389 (N_14389,N_14043,N_14109);
or U14390 (N_14390,N_14150,N_14013);
nor U14391 (N_14391,N_14064,N_14184);
nand U14392 (N_14392,N_14009,N_14146);
nand U14393 (N_14393,N_14057,N_14076);
nor U14394 (N_14394,N_14164,N_14021);
nor U14395 (N_14395,N_14130,N_14034);
xnor U14396 (N_14396,N_14016,N_14174);
and U14397 (N_14397,N_14074,N_14170);
nor U14398 (N_14398,N_14106,N_14124);
nor U14399 (N_14399,N_14151,N_14180);
nor U14400 (N_14400,N_14283,N_14250);
nor U14401 (N_14401,N_14356,N_14355);
nor U14402 (N_14402,N_14270,N_14298);
and U14403 (N_14403,N_14302,N_14216);
nor U14404 (N_14404,N_14230,N_14366);
xor U14405 (N_14405,N_14204,N_14310);
and U14406 (N_14406,N_14200,N_14398);
and U14407 (N_14407,N_14397,N_14215);
or U14408 (N_14408,N_14333,N_14324);
xnor U14409 (N_14409,N_14295,N_14307);
nand U14410 (N_14410,N_14218,N_14316);
xnor U14411 (N_14411,N_14344,N_14282);
or U14412 (N_14412,N_14217,N_14321);
xnor U14413 (N_14413,N_14374,N_14209);
xnor U14414 (N_14414,N_14348,N_14287);
and U14415 (N_14415,N_14343,N_14335);
nand U14416 (N_14416,N_14301,N_14375);
or U14417 (N_14417,N_14212,N_14376);
nand U14418 (N_14418,N_14372,N_14274);
nand U14419 (N_14419,N_14311,N_14323);
nand U14420 (N_14420,N_14243,N_14377);
xnor U14421 (N_14421,N_14308,N_14351);
or U14422 (N_14422,N_14225,N_14262);
or U14423 (N_14423,N_14220,N_14364);
nor U14424 (N_14424,N_14303,N_14305);
nor U14425 (N_14425,N_14349,N_14219);
or U14426 (N_14426,N_14222,N_14369);
nand U14427 (N_14427,N_14227,N_14382);
nand U14428 (N_14428,N_14389,N_14246);
xnor U14429 (N_14429,N_14354,N_14359);
and U14430 (N_14430,N_14306,N_14259);
xnor U14431 (N_14431,N_14313,N_14358);
and U14432 (N_14432,N_14342,N_14281);
and U14433 (N_14433,N_14241,N_14254);
nand U14434 (N_14434,N_14224,N_14368);
nor U14435 (N_14435,N_14360,N_14284);
and U14436 (N_14436,N_14249,N_14266);
and U14437 (N_14437,N_14253,N_14223);
nor U14438 (N_14438,N_14257,N_14340);
and U14439 (N_14439,N_14208,N_14336);
and U14440 (N_14440,N_14363,N_14330);
xnor U14441 (N_14441,N_14322,N_14395);
xnor U14442 (N_14442,N_14393,N_14292);
nor U14443 (N_14443,N_14352,N_14271);
xnor U14444 (N_14444,N_14207,N_14236);
and U14445 (N_14445,N_14309,N_14339);
nand U14446 (N_14446,N_14317,N_14232);
or U14447 (N_14447,N_14291,N_14385);
or U14448 (N_14448,N_14251,N_14296);
nor U14449 (N_14449,N_14312,N_14367);
nand U14450 (N_14450,N_14234,N_14371);
or U14451 (N_14451,N_14247,N_14226);
and U14452 (N_14452,N_14329,N_14214);
xor U14453 (N_14453,N_14387,N_14286);
xnor U14454 (N_14454,N_14265,N_14332);
xor U14455 (N_14455,N_14334,N_14289);
nor U14456 (N_14456,N_14331,N_14386);
xor U14457 (N_14457,N_14320,N_14228);
nand U14458 (N_14458,N_14273,N_14229);
nand U14459 (N_14459,N_14379,N_14205);
and U14460 (N_14460,N_14231,N_14221);
nand U14461 (N_14461,N_14337,N_14293);
nor U14462 (N_14462,N_14258,N_14338);
nor U14463 (N_14463,N_14350,N_14390);
and U14464 (N_14464,N_14238,N_14213);
nor U14465 (N_14465,N_14277,N_14314);
or U14466 (N_14466,N_14384,N_14304);
and U14467 (N_14467,N_14300,N_14315);
and U14468 (N_14468,N_14268,N_14362);
xor U14469 (N_14469,N_14242,N_14318);
nand U14470 (N_14470,N_14211,N_14244);
and U14471 (N_14471,N_14206,N_14260);
nand U14472 (N_14472,N_14269,N_14280);
and U14473 (N_14473,N_14272,N_14325);
nor U14474 (N_14474,N_14264,N_14392);
nand U14475 (N_14475,N_14380,N_14347);
or U14476 (N_14476,N_14326,N_14399);
and U14477 (N_14477,N_14378,N_14240);
and U14478 (N_14478,N_14263,N_14233);
or U14479 (N_14479,N_14319,N_14346);
xnor U14480 (N_14480,N_14285,N_14252);
or U14481 (N_14481,N_14267,N_14279);
nand U14482 (N_14482,N_14370,N_14278);
nand U14483 (N_14483,N_14235,N_14256);
nor U14484 (N_14484,N_14237,N_14394);
or U14485 (N_14485,N_14202,N_14245);
or U14486 (N_14486,N_14381,N_14357);
xnor U14487 (N_14487,N_14288,N_14361);
or U14488 (N_14488,N_14345,N_14248);
nand U14489 (N_14489,N_14275,N_14328);
xnor U14490 (N_14490,N_14290,N_14239);
and U14491 (N_14491,N_14365,N_14201);
and U14492 (N_14492,N_14383,N_14391);
nand U14493 (N_14493,N_14373,N_14299);
nor U14494 (N_14494,N_14210,N_14261);
and U14495 (N_14495,N_14276,N_14396);
nor U14496 (N_14496,N_14255,N_14341);
nor U14497 (N_14497,N_14388,N_14353);
and U14498 (N_14498,N_14327,N_14203);
xnor U14499 (N_14499,N_14294,N_14297);
and U14500 (N_14500,N_14382,N_14252);
and U14501 (N_14501,N_14366,N_14270);
or U14502 (N_14502,N_14395,N_14294);
or U14503 (N_14503,N_14312,N_14360);
or U14504 (N_14504,N_14216,N_14354);
and U14505 (N_14505,N_14295,N_14343);
xnor U14506 (N_14506,N_14354,N_14305);
xnor U14507 (N_14507,N_14358,N_14339);
or U14508 (N_14508,N_14285,N_14396);
xnor U14509 (N_14509,N_14276,N_14382);
and U14510 (N_14510,N_14309,N_14315);
nor U14511 (N_14511,N_14287,N_14368);
nor U14512 (N_14512,N_14348,N_14376);
and U14513 (N_14513,N_14335,N_14364);
or U14514 (N_14514,N_14332,N_14252);
or U14515 (N_14515,N_14296,N_14375);
xor U14516 (N_14516,N_14243,N_14266);
xnor U14517 (N_14517,N_14371,N_14269);
nand U14518 (N_14518,N_14374,N_14282);
or U14519 (N_14519,N_14360,N_14310);
nand U14520 (N_14520,N_14334,N_14283);
nor U14521 (N_14521,N_14217,N_14398);
or U14522 (N_14522,N_14278,N_14215);
or U14523 (N_14523,N_14335,N_14250);
nor U14524 (N_14524,N_14246,N_14308);
or U14525 (N_14525,N_14336,N_14237);
and U14526 (N_14526,N_14344,N_14356);
nand U14527 (N_14527,N_14248,N_14315);
nor U14528 (N_14528,N_14218,N_14243);
and U14529 (N_14529,N_14246,N_14228);
xor U14530 (N_14530,N_14322,N_14242);
or U14531 (N_14531,N_14206,N_14262);
and U14532 (N_14532,N_14212,N_14378);
or U14533 (N_14533,N_14304,N_14292);
and U14534 (N_14534,N_14285,N_14316);
and U14535 (N_14535,N_14393,N_14216);
and U14536 (N_14536,N_14398,N_14220);
nand U14537 (N_14537,N_14314,N_14386);
or U14538 (N_14538,N_14233,N_14267);
or U14539 (N_14539,N_14360,N_14367);
and U14540 (N_14540,N_14297,N_14228);
and U14541 (N_14541,N_14277,N_14365);
xnor U14542 (N_14542,N_14321,N_14221);
or U14543 (N_14543,N_14215,N_14242);
and U14544 (N_14544,N_14329,N_14361);
xnor U14545 (N_14545,N_14200,N_14203);
or U14546 (N_14546,N_14209,N_14328);
nand U14547 (N_14547,N_14293,N_14270);
or U14548 (N_14548,N_14315,N_14261);
nor U14549 (N_14549,N_14212,N_14395);
and U14550 (N_14550,N_14275,N_14278);
xor U14551 (N_14551,N_14345,N_14336);
nor U14552 (N_14552,N_14237,N_14240);
and U14553 (N_14553,N_14319,N_14360);
nor U14554 (N_14554,N_14228,N_14391);
and U14555 (N_14555,N_14329,N_14306);
and U14556 (N_14556,N_14288,N_14203);
nand U14557 (N_14557,N_14271,N_14235);
and U14558 (N_14558,N_14384,N_14280);
or U14559 (N_14559,N_14300,N_14278);
or U14560 (N_14560,N_14253,N_14248);
and U14561 (N_14561,N_14257,N_14300);
and U14562 (N_14562,N_14380,N_14215);
nor U14563 (N_14563,N_14269,N_14389);
or U14564 (N_14564,N_14396,N_14308);
nand U14565 (N_14565,N_14248,N_14389);
xnor U14566 (N_14566,N_14267,N_14265);
and U14567 (N_14567,N_14245,N_14240);
nor U14568 (N_14568,N_14380,N_14254);
nor U14569 (N_14569,N_14273,N_14354);
and U14570 (N_14570,N_14395,N_14388);
nor U14571 (N_14571,N_14396,N_14326);
and U14572 (N_14572,N_14327,N_14392);
or U14573 (N_14573,N_14325,N_14319);
or U14574 (N_14574,N_14206,N_14291);
nor U14575 (N_14575,N_14219,N_14256);
nand U14576 (N_14576,N_14261,N_14202);
xnor U14577 (N_14577,N_14304,N_14261);
or U14578 (N_14578,N_14247,N_14380);
and U14579 (N_14579,N_14397,N_14391);
nor U14580 (N_14580,N_14311,N_14356);
or U14581 (N_14581,N_14327,N_14344);
xor U14582 (N_14582,N_14324,N_14361);
nor U14583 (N_14583,N_14240,N_14270);
nor U14584 (N_14584,N_14385,N_14248);
nand U14585 (N_14585,N_14386,N_14294);
nand U14586 (N_14586,N_14327,N_14307);
xnor U14587 (N_14587,N_14269,N_14333);
nand U14588 (N_14588,N_14261,N_14378);
or U14589 (N_14589,N_14398,N_14238);
and U14590 (N_14590,N_14365,N_14227);
nand U14591 (N_14591,N_14304,N_14246);
nand U14592 (N_14592,N_14287,N_14329);
xor U14593 (N_14593,N_14307,N_14303);
and U14594 (N_14594,N_14370,N_14324);
or U14595 (N_14595,N_14397,N_14398);
xnor U14596 (N_14596,N_14300,N_14284);
or U14597 (N_14597,N_14330,N_14211);
nand U14598 (N_14598,N_14300,N_14267);
xor U14599 (N_14599,N_14322,N_14270);
xnor U14600 (N_14600,N_14445,N_14545);
nor U14601 (N_14601,N_14546,N_14485);
xnor U14602 (N_14602,N_14450,N_14573);
and U14603 (N_14603,N_14424,N_14409);
or U14604 (N_14604,N_14444,N_14541);
xor U14605 (N_14605,N_14499,N_14598);
nand U14606 (N_14606,N_14454,N_14477);
nand U14607 (N_14607,N_14407,N_14491);
nor U14608 (N_14608,N_14456,N_14542);
xnor U14609 (N_14609,N_14516,N_14514);
and U14610 (N_14610,N_14552,N_14536);
nand U14611 (N_14611,N_14522,N_14404);
and U14612 (N_14612,N_14592,N_14558);
xor U14613 (N_14613,N_14588,N_14420);
xnor U14614 (N_14614,N_14433,N_14412);
nand U14615 (N_14615,N_14490,N_14438);
and U14616 (N_14616,N_14557,N_14482);
xor U14617 (N_14617,N_14535,N_14565);
nor U14618 (N_14618,N_14504,N_14550);
nor U14619 (N_14619,N_14524,N_14411);
nand U14620 (N_14620,N_14540,N_14478);
or U14621 (N_14621,N_14533,N_14572);
nor U14622 (N_14622,N_14589,N_14419);
and U14623 (N_14623,N_14455,N_14489);
and U14624 (N_14624,N_14422,N_14510);
and U14625 (N_14625,N_14492,N_14580);
or U14626 (N_14626,N_14447,N_14413);
nand U14627 (N_14627,N_14556,N_14562);
or U14628 (N_14628,N_14576,N_14579);
nand U14629 (N_14629,N_14534,N_14594);
nor U14630 (N_14630,N_14507,N_14437);
nor U14631 (N_14631,N_14432,N_14453);
xor U14632 (N_14632,N_14520,N_14584);
and U14633 (N_14633,N_14566,N_14476);
xnor U14634 (N_14634,N_14505,N_14560);
and U14635 (N_14635,N_14449,N_14434);
or U14636 (N_14636,N_14425,N_14486);
nand U14637 (N_14637,N_14513,N_14537);
nand U14638 (N_14638,N_14528,N_14578);
nand U14639 (N_14639,N_14583,N_14549);
nand U14640 (N_14640,N_14501,N_14443);
xor U14641 (N_14641,N_14408,N_14543);
and U14642 (N_14642,N_14400,N_14519);
nor U14643 (N_14643,N_14575,N_14568);
or U14644 (N_14644,N_14547,N_14431);
or U14645 (N_14645,N_14590,N_14571);
nand U14646 (N_14646,N_14471,N_14487);
nand U14647 (N_14647,N_14585,N_14500);
and U14648 (N_14648,N_14531,N_14591);
nand U14649 (N_14649,N_14523,N_14496);
xor U14650 (N_14650,N_14518,N_14439);
and U14651 (N_14651,N_14430,N_14581);
or U14652 (N_14652,N_14483,N_14506);
or U14653 (N_14653,N_14452,N_14423);
and U14654 (N_14654,N_14587,N_14475);
nor U14655 (N_14655,N_14498,N_14561);
nor U14656 (N_14656,N_14508,N_14529);
and U14657 (N_14657,N_14551,N_14570);
xnor U14658 (N_14658,N_14410,N_14402);
xor U14659 (N_14659,N_14401,N_14509);
and U14660 (N_14660,N_14493,N_14466);
and U14661 (N_14661,N_14427,N_14479);
and U14662 (N_14662,N_14461,N_14469);
xnor U14663 (N_14663,N_14544,N_14448);
nand U14664 (N_14664,N_14414,N_14480);
xor U14665 (N_14665,N_14586,N_14511);
nand U14666 (N_14666,N_14460,N_14468);
xor U14667 (N_14667,N_14472,N_14488);
or U14668 (N_14668,N_14563,N_14462);
and U14669 (N_14669,N_14539,N_14484);
or U14670 (N_14670,N_14418,N_14467);
and U14671 (N_14671,N_14548,N_14415);
xnor U14672 (N_14672,N_14559,N_14569);
and U14673 (N_14673,N_14503,N_14497);
or U14674 (N_14674,N_14596,N_14458);
nor U14675 (N_14675,N_14494,N_14554);
xnor U14676 (N_14676,N_14481,N_14428);
xor U14677 (N_14677,N_14463,N_14582);
and U14678 (N_14678,N_14515,N_14451);
or U14679 (N_14679,N_14421,N_14446);
nand U14680 (N_14680,N_14459,N_14574);
or U14681 (N_14681,N_14440,N_14532);
xnor U14682 (N_14682,N_14436,N_14464);
or U14683 (N_14683,N_14593,N_14435);
xor U14684 (N_14684,N_14526,N_14555);
nand U14685 (N_14685,N_14597,N_14406);
nand U14686 (N_14686,N_14599,N_14470);
xnor U14687 (N_14687,N_14429,N_14416);
nor U14688 (N_14688,N_14457,N_14426);
or U14689 (N_14689,N_14495,N_14465);
and U14690 (N_14690,N_14502,N_14577);
xnor U14691 (N_14691,N_14567,N_14473);
and U14692 (N_14692,N_14442,N_14527);
or U14693 (N_14693,N_14595,N_14530);
xnor U14694 (N_14694,N_14553,N_14403);
and U14695 (N_14695,N_14441,N_14512);
nand U14696 (N_14696,N_14474,N_14517);
nand U14697 (N_14697,N_14538,N_14564);
nand U14698 (N_14698,N_14405,N_14417);
or U14699 (N_14699,N_14525,N_14521);
or U14700 (N_14700,N_14409,N_14473);
and U14701 (N_14701,N_14511,N_14417);
nor U14702 (N_14702,N_14422,N_14501);
and U14703 (N_14703,N_14416,N_14557);
nand U14704 (N_14704,N_14508,N_14598);
nor U14705 (N_14705,N_14521,N_14553);
nand U14706 (N_14706,N_14592,N_14455);
xor U14707 (N_14707,N_14495,N_14419);
and U14708 (N_14708,N_14466,N_14558);
xor U14709 (N_14709,N_14581,N_14465);
or U14710 (N_14710,N_14581,N_14475);
nand U14711 (N_14711,N_14485,N_14468);
and U14712 (N_14712,N_14503,N_14403);
nor U14713 (N_14713,N_14564,N_14485);
nand U14714 (N_14714,N_14429,N_14474);
nand U14715 (N_14715,N_14436,N_14415);
nor U14716 (N_14716,N_14446,N_14534);
and U14717 (N_14717,N_14440,N_14507);
nand U14718 (N_14718,N_14445,N_14437);
xnor U14719 (N_14719,N_14435,N_14538);
nand U14720 (N_14720,N_14413,N_14517);
or U14721 (N_14721,N_14464,N_14428);
and U14722 (N_14722,N_14447,N_14537);
or U14723 (N_14723,N_14532,N_14447);
xor U14724 (N_14724,N_14581,N_14451);
and U14725 (N_14725,N_14562,N_14501);
and U14726 (N_14726,N_14599,N_14479);
or U14727 (N_14727,N_14452,N_14498);
and U14728 (N_14728,N_14447,N_14496);
nor U14729 (N_14729,N_14583,N_14406);
and U14730 (N_14730,N_14450,N_14583);
xor U14731 (N_14731,N_14546,N_14514);
and U14732 (N_14732,N_14576,N_14404);
and U14733 (N_14733,N_14499,N_14496);
nor U14734 (N_14734,N_14559,N_14452);
or U14735 (N_14735,N_14592,N_14422);
or U14736 (N_14736,N_14465,N_14418);
nand U14737 (N_14737,N_14464,N_14594);
nand U14738 (N_14738,N_14469,N_14406);
xnor U14739 (N_14739,N_14594,N_14434);
and U14740 (N_14740,N_14581,N_14407);
or U14741 (N_14741,N_14577,N_14583);
nand U14742 (N_14742,N_14587,N_14503);
or U14743 (N_14743,N_14497,N_14409);
nor U14744 (N_14744,N_14522,N_14432);
nor U14745 (N_14745,N_14555,N_14412);
nor U14746 (N_14746,N_14569,N_14482);
nor U14747 (N_14747,N_14494,N_14508);
xor U14748 (N_14748,N_14558,N_14524);
xor U14749 (N_14749,N_14516,N_14508);
nand U14750 (N_14750,N_14533,N_14549);
and U14751 (N_14751,N_14593,N_14584);
nand U14752 (N_14752,N_14481,N_14402);
nor U14753 (N_14753,N_14525,N_14562);
xnor U14754 (N_14754,N_14474,N_14434);
and U14755 (N_14755,N_14401,N_14488);
and U14756 (N_14756,N_14409,N_14523);
or U14757 (N_14757,N_14523,N_14504);
nor U14758 (N_14758,N_14532,N_14426);
xor U14759 (N_14759,N_14571,N_14551);
nor U14760 (N_14760,N_14422,N_14558);
nor U14761 (N_14761,N_14544,N_14584);
nor U14762 (N_14762,N_14500,N_14536);
nor U14763 (N_14763,N_14560,N_14477);
nor U14764 (N_14764,N_14575,N_14567);
and U14765 (N_14765,N_14571,N_14472);
or U14766 (N_14766,N_14434,N_14523);
nor U14767 (N_14767,N_14433,N_14420);
xor U14768 (N_14768,N_14486,N_14592);
nand U14769 (N_14769,N_14453,N_14400);
nand U14770 (N_14770,N_14422,N_14541);
and U14771 (N_14771,N_14576,N_14499);
xnor U14772 (N_14772,N_14515,N_14526);
nand U14773 (N_14773,N_14535,N_14436);
nor U14774 (N_14774,N_14547,N_14592);
nor U14775 (N_14775,N_14478,N_14492);
nor U14776 (N_14776,N_14509,N_14480);
nor U14777 (N_14777,N_14473,N_14489);
and U14778 (N_14778,N_14518,N_14480);
nor U14779 (N_14779,N_14413,N_14400);
or U14780 (N_14780,N_14567,N_14422);
xnor U14781 (N_14781,N_14549,N_14587);
nand U14782 (N_14782,N_14460,N_14501);
nor U14783 (N_14783,N_14447,N_14432);
and U14784 (N_14784,N_14539,N_14530);
xnor U14785 (N_14785,N_14436,N_14529);
or U14786 (N_14786,N_14445,N_14507);
nor U14787 (N_14787,N_14463,N_14596);
or U14788 (N_14788,N_14494,N_14556);
nand U14789 (N_14789,N_14437,N_14582);
or U14790 (N_14790,N_14526,N_14473);
nor U14791 (N_14791,N_14430,N_14418);
xor U14792 (N_14792,N_14544,N_14573);
or U14793 (N_14793,N_14571,N_14470);
nand U14794 (N_14794,N_14580,N_14562);
and U14795 (N_14795,N_14524,N_14440);
nand U14796 (N_14796,N_14472,N_14563);
and U14797 (N_14797,N_14405,N_14425);
nor U14798 (N_14798,N_14573,N_14425);
nor U14799 (N_14799,N_14478,N_14548);
nor U14800 (N_14800,N_14699,N_14661);
xnor U14801 (N_14801,N_14759,N_14748);
xnor U14802 (N_14802,N_14691,N_14666);
and U14803 (N_14803,N_14637,N_14774);
or U14804 (N_14804,N_14631,N_14690);
nand U14805 (N_14805,N_14708,N_14744);
nor U14806 (N_14806,N_14641,N_14706);
and U14807 (N_14807,N_14632,N_14634);
xnor U14808 (N_14808,N_14628,N_14607);
and U14809 (N_14809,N_14784,N_14646);
or U14810 (N_14810,N_14602,N_14705);
xor U14811 (N_14811,N_14648,N_14605);
nand U14812 (N_14812,N_14766,N_14664);
nand U14813 (N_14813,N_14787,N_14617);
and U14814 (N_14814,N_14716,N_14678);
and U14815 (N_14815,N_14712,N_14680);
and U14816 (N_14816,N_14669,N_14717);
xor U14817 (N_14817,N_14612,N_14609);
or U14818 (N_14818,N_14729,N_14613);
or U14819 (N_14819,N_14772,N_14786);
and U14820 (N_14820,N_14677,N_14737);
nor U14821 (N_14821,N_14740,N_14765);
nand U14822 (N_14822,N_14643,N_14697);
xnor U14823 (N_14823,N_14734,N_14684);
xnor U14824 (N_14824,N_14771,N_14660);
or U14825 (N_14825,N_14640,N_14624);
and U14826 (N_14826,N_14749,N_14606);
xor U14827 (N_14827,N_14788,N_14743);
xor U14828 (N_14828,N_14603,N_14656);
or U14829 (N_14829,N_14770,N_14611);
or U14830 (N_14830,N_14638,N_14618);
nand U14831 (N_14831,N_14693,N_14736);
or U14832 (N_14832,N_14604,N_14727);
xnor U14833 (N_14833,N_14630,N_14713);
xnor U14834 (N_14834,N_14614,N_14763);
nand U14835 (N_14835,N_14670,N_14703);
nand U14836 (N_14836,N_14700,N_14667);
or U14837 (N_14837,N_14783,N_14782);
and U14838 (N_14838,N_14742,N_14764);
xnor U14839 (N_14839,N_14781,N_14775);
and U14840 (N_14840,N_14710,N_14768);
xor U14841 (N_14841,N_14674,N_14636);
and U14842 (N_14842,N_14778,N_14639);
and U14843 (N_14843,N_14653,N_14719);
nand U14844 (N_14844,N_14725,N_14792);
and U14845 (N_14845,N_14791,N_14761);
nor U14846 (N_14846,N_14668,N_14696);
xor U14847 (N_14847,N_14673,N_14754);
or U14848 (N_14848,N_14789,N_14780);
xnor U14849 (N_14849,N_14659,N_14663);
nand U14850 (N_14850,N_14651,N_14658);
or U14851 (N_14851,N_14623,N_14649);
or U14852 (N_14852,N_14654,N_14635);
nor U14853 (N_14853,N_14704,N_14616);
nand U14854 (N_14854,N_14620,N_14799);
nand U14855 (N_14855,N_14753,N_14672);
and U14856 (N_14856,N_14608,N_14755);
nor U14857 (N_14857,N_14702,N_14724);
and U14858 (N_14858,N_14796,N_14715);
nor U14859 (N_14859,N_14714,N_14642);
or U14860 (N_14860,N_14720,N_14665);
nor U14861 (N_14861,N_14655,N_14644);
nand U14862 (N_14862,N_14752,N_14757);
or U14863 (N_14863,N_14730,N_14692);
xor U14864 (N_14864,N_14785,N_14647);
xor U14865 (N_14865,N_14769,N_14679);
xnor U14866 (N_14866,N_14707,N_14681);
xor U14867 (N_14867,N_14735,N_14779);
nand U14868 (N_14868,N_14621,N_14688);
and U14869 (N_14869,N_14662,N_14777);
nand U14870 (N_14870,N_14619,N_14747);
and U14871 (N_14871,N_14652,N_14610);
nor U14872 (N_14872,N_14682,N_14794);
xnor U14873 (N_14873,N_14626,N_14746);
and U14874 (N_14874,N_14683,N_14615);
nor U14875 (N_14875,N_14711,N_14728);
nand U14876 (N_14876,N_14797,N_14622);
nand U14877 (N_14877,N_14758,N_14760);
and U14878 (N_14878,N_14675,N_14698);
nor U14879 (N_14879,N_14709,N_14793);
or U14880 (N_14880,N_14625,N_14671);
xor U14881 (N_14881,N_14695,N_14726);
and U14882 (N_14882,N_14629,N_14676);
and U14883 (N_14883,N_14633,N_14718);
nor U14884 (N_14884,N_14650,N_14657);
nand U14885 (N_14885,N_14722,N_14731);
xnor U14886 (N_14886,N_14686,N_14751);
xnor U14887 (N_14887,N_14745,N_14750);
xnor U14888 (N_14888,N_14701,N_14790);
nor U14889 (N_14889,N_14600,N_14685);
or U14890 (N_14890,N_14694,N_14776);
nand U14891 (N_14891,N_14741,N_14627);
or U14892 (N_14892,N_14733,N_14756);
and U14893 (N_14893,N_14645,N_14795);
nand U14894 (N_14894,N_14767,N_14732);
and U14895 (N_14895,N_14721,N_14773);
nor U14896 (N_14896,N_14739,N_14601);
nand U14897 (N_14897,N_14762,N_14689);
nand U14898 (N_14898,N_14738,N_14723);
or U14899 (N_14899,N_14687,N_14798);
nor U14900 (N_14900,N_14702,N_14679);
xnor U14901 (N_14901,N_14734,N_14796);
nor U14902 (N_14902,N_14715,N_14663);
or U14903 (N_14903,N_14689,N_14647);
nor U14904 (N_14904,N_14648,N_14700);
xnor U14905 (N_14905,N_14729,N_14685);
or U14906 (N_14906,N_14689,N_14733);
xnor U14907 (N_14907,N_14662,N_14779);
nand U14908 (N_14908,N_14606,N_14600);
nor U14909 (N_14909,N_14691,N_14780);
and U14910 (N_14910,N_14622,N_14735);
or U14911 (N_14911,N_14783,N_14792);
xnor U14912 (N_14912,N_14603,N_14785);
and U14913 (N_14913,N_14601,N_14690);
nand U14914 (N_14914,N_14615,N_14724);
and U14915 (N_14915,N_14649,N_14610);
nor U14916 (N_14916,N_14663,N_14648);
nand U14917 (N_14917,N_14618,N_14645);
or U14918 (N_14918,N_14726,N_14769);
or U14919 (N_14919,N_14752,N_14671);
nand U14920 (N_14920,N_14799,N_14696);
and U14921 (N_14921,N_14607,N_14650);
nor U14922 (N_14922,N_14618,N_14620);
nand U14923 (N_14923,N_14725,N_14747);
and U14924 (N_14924,N_14793,N_14722);
nor U14925 (N_14925,N_14629,N_14715);
nor U14926 (N_14926,N_14719,N_14640);
or U14927 (N_14927,N_14601,N_14701);
or U14928 (N_14928,N_14798,N_14618);
nor U14929 (N_14929,N_14607,N_14776);
nor U14930 (N_14930,N_14699,N_14792);
xnor U14931 (N_14931,N_14638,N_14602);
nand U14932 (N_14932,N_14714,N_14732);
nor U14933 (N_14933,N_14626,N_14797);
nand U14934 (N_14934,N_14603,N_14602);
xor U14935 (N_14935,N_14600,N_14646);
xor U14936 (N_14936,N_14635,N_14738);
or U14937 (N_14937,N_14613,N_14686);
xor U14938 (N_14938,N_14730,N_14678);
nand U14939 (N_14939,N_14671,N_14735);
xnor U14940 (N_14940,N_14651,N_14715);
nor U14941 (N_14941,N_14681,N_14726);
or U14942 (N_14942,N_14662,N_14631);
or U14943 (N_14943,N_14662,N_14684);
or U14944 (N_14944,N_14700,N_14614);
nand U14945 (N_14945,N_14693,N_14688);
xor U14946 (N_14946,N_14726,N_14697);
and U14947 (N_14947,N_14776,N_14661);
nor U14948 (N_14948,N_14691,N_14725);
or U14949 (N_14949,N_14722,N_14778);
or U14950 (N_14950,N_14622,N_14744);
or U14951 (N_14951,N_14601,N_14716);
xnor U14952 (N_14952,N_14654,N_14727);
nand U14953 (N_14953,N_14733,N_14674);
or U14954 (N_14954,N_14611,N_14711);
xnor U14955 (N_14955,N_14735,N_14763);
xor U14956 (N_14956,N_14766,N_14718);
nor U14957 (N_14957,N_14755,N_14678);
and U14958 (N_14958,N_14775,N_14675);
xor U14959 (N_14959,N_14791,N_14730);
nor U14960 (N_14960,N_14621,N_14686);
nand U14961 (N_14961,N_14780,N_14738);
xnor U14962 (N_14962,N_14714,N_14672);
and U14963 (N_14963,N_14650,N_14706);
and U14964 (N_14964,N_14649,N_14657);
xor U14965 (N_14965,N_14774,N_14795);
and U14966 (N_14966,N_14785,N_14703);
nor U14967 (N_14967,N_14680,N_14658);
and U14968 (N_14968,N_14707,N_14742);
or U14969 (N_14969,N_14700,N_14771);
or U14970 (N_14970,N_14749,N_14793);
nor U14971 (N_14971,N_14767,N_14662);
xor U14972 (N_14972,N_14784,N_14697);
nand U14973 (N_14973,N_14714,N_14707);
nand U14974 (N_14974,N_14696,N_14767);
xor U14975 (N_14975,N_14674,N_14737);
or U14976 (N_14976,N_14663,N_14701);
and U14977 (N_14977,N_14729,N_14612);
xor U14978 (N_14978,N_14675,N_14738);
nand U14979 (N_14979,N_14625,N_14715);
nor U14980 (N_14980,N_14778,N_14714);
and U14981 (N_14981,N_14659,N_14613);
nor U14982 (N_14982,N_14617,N_14739);
nor U14983 (N_14983,N_14609,N_14721);
and U14984 (N_14984,N_14784,N_14725);
nand U14985 (N_14985,N_14635,N_14649);
xor U14986 (N_14986,N_14709,N_14689);
nand U14987 (N_14987,N_14646,N_14793);
nand U14988 (N_14988,N_14629,N_14625);
or U14989 (N_14989,N_14606,N_14753);
and U14990 (N_14990,N_14655,N_14745);
or U14991 (N_14991,N_14733,N_14764);
or U14992 (N_14992,N_14655,N_14704);
nand U14993 (N_14993,N_14661,N_14629);
nand U14994 (N_14994,N_14604,N_14706);
and U14995 (N_14995,N_14785,N_14732);
nand U14996 (N_14996,N_14737,N_14740);
nor U14997 (N_14997,N_14749,N_14618);
and U14998 (N_14998,N_14644,N_14678);
or U14999 (N_14999,N_14612,N_14696);
or U15000 (N_15000,N_14818,N_14996);
nor U15001 (N_15001,N_14868,N_14886);
and U15002 (N_15002,N_14890,N_14845);
and U15003 (N_15003,N_14903,N_14877);
xnor U15004 (N_15004,N_14949,N_14927);
or U15005 (N_15005,N_14912,N_14973);
nor U15006 (N_15006,N_14917,N_14867);
nand U15007 (N_15007,N_14839,N_14929);
and U15008 (N_15008,N_14935,N_14872);
and U15009 (N_15009,N_14966,N_14953);
nor U15010 (N_15010,N_14863,N_14820);
nand U15011 (N_15011,N_14972,N_14937);
or U15012 (N_15012,N_14978,N_14908);
nand U15013 (N_15013,N_14964,N_14984);
nand U15014 (N_15014,N_14888,N_14833);
nand U15015 (N_15015,N_14914,N_14826);
or U15016 (N_15016,N_14898,N_14962);
nand U15017 (N_15017,N_14813,N_14878);
and U15018 (N_15018,N_14836,N_14852);
nand U15019 (N_15019,N_14889,N_14842);
xor U15020 (N_15020,N_14938,N_14926);
nor U15021 (N_15021,N_14800,N_14998);
or U15022 (N_15022,N_14987,N_14940);
nor U15023 (N_15023,N_14967,N_14835);
and U15024 (N_15024,N_14932,N_14849);
nor U15025 (N_15025,N_14854,N_14944);
nand U15026 (N_15026,N_14858,N_14834);
or U15027 (N_15027,N_14915,N_14906);
nand U15028 (N_15028,N_14832,N_14986);
nor U15029 (N_15029,N_14913,N_14840);
or U15030 (N_15030,N_14943,N_14866);
and U15031 (N_15031,N_14851,N_14985);
or U15032 (N_15032,N_14933,N_14814);
and U15033 (N_15033,N_14805,N_14995);
and U15034 (N_15034,N_14844,N_14961);
or U15035 (N_15035,N_14952,N_14801);
xnor U15036 (N_15036,N_14930,N_14853);
or U15037 (N_15037,N_14883,N_14823);
nand U15038 (N_15038,N_14880,N_14936);
xnor U15039 (N_15039,N_14921,N_14956);
nand U15040 (N_15040,N_14875,N_14893);
xor U15041 (N_15041,N_14896,N_14892);
and U15042 (N_15042,N_14825,N_14855);
or U15043 (N_15043,N_14948,N_14870);
nand U15044 (N_15044,N_14955,N_14869);
nand U15045 (N_15045,N_14822,N_14860);
and U15046 (N_15046,N_14969,N_14876);
nor U15047 (N_15047,N_14811,N_14827);
and U15048 (N_15048,N_14924,N_14991);
nor U15049 (N_15049,N_14843,N_14904);
and U15050 (N_15050,N_14862,N_14957);
and U15051 (N_15051,N_14992,N_14838);
xor U15052 (N_15052,N_14997,N_14871);
and U15053 (N_15053,N_14803,N_14900);
or U15054 (N_15054,N_14928,N_14994);
xnor U15055 (N_15055,N_14816,N_14907);
nand U15056 (N_15056,N_14941,N_14828);
xnor U15057 (N_15057,N_14939,N_14905);
nor U15058 (N_15058,N_14887,N_14884);
nor U15059 (N_15059,N_14873,N_14946);
and U15060 (N_15060,N_14945,N_14918);
and U15061 (N_15061,N_14885,N_14861);
or U15062 (N_15062,N_14895,N_14989);
xor U15063 (N_15063,N_14879,N_14993);
nor U15064 (N_15064,N_14831,N_14958);
and U15065 (N_15065,N_14902,N_14807);
nor U15066 (N_15066,N_14812,N_14881);
or U15067 (N_15067,N_14865,N_14976);
nor U15068 (N_15068,N_14979,N_14824);
or U15069 (N_15069,N_14857,N_14804);
nand U15070 (N_15070,N_14981,N_14971);
nor U15071 (N_15071,N_14874,N_14977);
nand U15072 (N_15072,N_14864,N_14965);
and U15073 (N_15073,N_14809,N_14934);
and U15074 (N_15074,N_14894,N_14970);
nand U15075 (N_15075,N_14841,N_14848);
or U15076 (N_15076,N_14942,N_14974);
nor U15077 (N_15077,N_14931,N_14999);
and U15078 (N_15078,N_14963,N_14830);
nand U15079 (N_15079,N_14920,N_14982);
or U15080 (N_15080,N_14975,N_14850);
nand U15081 (N_15081,N_14859,N_14988);
xnor U15082 (N_15082,N_14910,N_14954);
or U15083 (N_15083,N_14980,N_14909);
and U15084 (N_15084,N_14911,N_14901);
xor U15085 (N_15085,N_14923,N_14847);
nand U15086 (N_15086,N_14950,N_14990);
nor U15087 (N_15087,N_14947,N_14821);
and U15088 (N_15088,N_14968,N_14960);
or U15089 (N_15089,N_14983,N_14919);
xnor U15090 (N_15090,N_14815,N_14899);
nor U15091 (N_15091,N_14959,N_14882);
nor U15092 (N_15092,N_14810,N_14916);
or U15093 (N_15093,N_14806,N_14817);
nor U15094 (N_15094,N_14829,N_14856);
and U15095 (N_15095,N_14837,N_14846);
nor U15096 (N_15096,N_14925,N_14951);
or U15097 (N_15097,N_14922,N_14802);
or U15098 (N_15098,N_14819,N_14891);
nor U15099 (N_15099,N_14808,N_14897);
xnor U15100 (N_15100,N_14918,N_14936);
and U15101 (N_15101,N_14869,N_14841);
xnor U15102 (N_15102,N_14886,N_14890);
nor U15103 (N_15103,N_14857,N_14811);
or U15104 (N_15104,N_14840,N_14851);
nor U15105 (N_15105,N_14958,N_14853);
xnor U15106 (N_15106,N_14806,N_14862);
or U15107 (N_15107,N_14899,N_14944);
and U15108 (N_15108,N_14811,N_14834);
and U15109 (N_15109,N_14900,N_14989);
xnor U15110 (N_15110,N_14840,N_14995);
nand U15111 (N_15111,N_14977,N_14880);
or U15112 (N_15112,N_14960,N_14849);
xnor U15113 (N_15113,N_14914,N_14874);
and U15114 (N_15114,N_14844,N_14891);
and U15115 (N_15115,N_14803,N_14800);
and U15116 (N_15116,N_14847,N_14962);
and U15117 (N_15117,N_14950,N_14930);
and U15118 (N_15118,N_14988,N_14946);
or U15119 (N_15119,N_14913,N_14854);
or U15120 (N_15120,N_14952,N_14887);
nor U15121 (N_15121,N_14889,N_14992);
nor U15122 (N_15122,N_14843,N_14940);
or U15123 (N_15123,N_14824,N_14839);
xor U15124 (N_15124,N_14989,N_14932);
or U15125 (N_15125,N_14909,N_14858);
nor U15126 (N_15126,N_14818,N_14870);
xor U15127 (N_15127,N_14887,N_14821);
xnor U15128 (N_15128,N_14909,N_14911);
nor U15129 (N_15129,N_14837,N_14820);
or U15130 (N_15130,N_14940,N_14859);
nor U15131 (N_15131,N_14985,N_14964);
and U15132 (N_15132,N_14850,N_14841);
and U15133 (N_15133,N_14853,N_14807);
xnor U15134 (N_15134,N_14804,N_14904);
xor U15135 (N_15135,N_14994,N_14939);
and U15136 (N_15136,N_14866,N_14845);
xor U15137 (N_15137,N_14988,N_14928);
xor U15138 (N_15138,N_14808,N_14902);
or U15139 (N_15139,N_14929,N_14886);
nand U15140 (N_15140,N_14908,N_14871);
and U15141 (N_15141,N_14986,N_14816);
nor U15142 (N_15142,N_14978,N_14951);
xnor U15143 (N_15143,N_14923,N_14832);
and U15144 (N_15144,N_14859,N_14846);
and U15145 (N_15145,N_14819,N_14995);
and U15146 (N_15146,N_14830,N_14896);
nor U15147 (N_15147,N_14830,N_14861);
or U15148 (N_15148,N_14910,N_14868);
and U15149 (N_15149,N_14962,N_14998);
nand U15150 (N_15150,N_14943,N_14971);
xor U15151 (N_15151,N_14945,N_14802);
xnor U15152 (N_15152,N_14915,N_14932);
and U15153 (N_15153,N_14946,N_14920);
or U15154 (N_15154,N_14836,N_14830);
and U15155 (N_15155,N_14999,N_14927);
and U15156 (N_15156,N_14989,N_14923);
nor U15157 (N_15157,N_14913,N_14855);
or U15158 (N_15158,N_14825,N_14998);
nor U15159 (N_15159,N_14928,N_14933);
or U15160 (N_15160,N_14917,N_14936);
xnor U15161 (N_15161,N_14872,N_14898);
or U15162 (N_15162,N_14838,N_14990);
nor U15163 (N_15163,N_14971,N_14979);
xnor U15164 (N_15164,N_14973,N_14931);
xor U15165 (N_15165,N_14863,N_14971);
and U15166 (N_15166,N_14963,N_14889);
or U15167 (N_15167,N_14946,N_14898);
xor U15168 (N_15168,N_14897,N_14849);
nor U15169 (N_15169,N_14903,N_14963);
nand U15170 (N_15170,N_14917,N_14831);
xor U15171 (N_15171,N_14979,N_14944);
and U15172 (N_15172,N_14824,N_14850);
or U15173 (N_15173,N_14939,N_14926);
xor U15174 (N_15174,N_14919,N_14994);
xor U15175 (N_15175,N_14882,N_14952);
nor U15176 (N_15176,N_14952,N_14939);
and U15177 (N_15177,N_14920,N_14803);
xnor U15178 (N_15178,N_14966,N_14859);
nor U15179 (N_15179,N_14866,N_14934);
nand U15180 (N_15180,N_14959,N_14950);
and U15181 (N_15181,N_14998,N_14841);
and U15182 (N_15182,N_14929,N_14829);
or U15183 (N_15183,N_14826,N_14867);
nand U15184 (N_15184,N_14819,N_14806);
or U15185 (N_15185,N_14932,N_14833);
nor U15186 (N_15186,N_14973,N_14954);
xor U15187 (N_15187,N_14949,N_14978);
or U15188 (N_15188,N_14862,N_14896);
and U15189 (N_15189,N_14950,N_14875);
nand U15190 (N_15190,N_14921,N_14936);
nand U15191 (N_15191,N_14968,N_14940);
or U15192 (N_15192,N_14808,N_14836);
nand U15193 (N_15193,N_14905,N_14950);
nor U15194 (N_15194,N_14976,N_14951);
and U15195 (N_15195,N_14935,N_14932);
xnor U15196 (N_15196,N_14961,N_14930);
xor U15197 (N_15197,N_14913,N_14875);
nor U15198 (N_15198,N_14914,N_14857);
or U15199 (N_15199,N_14913,N_14907);
or U15200 (N_15200,N_15042,N_15027);
and U15201 (N_15201,N_15029,N_15104);
nand U15202 (N_15202,N_15069,N_15190);
and U15203 (N_15203,N_15116,N_15121);
nor U15204 (N_15204,N_15179,N_15187);
or U15205 (N_15205,N_15053,N_15033);
nand U15206 (N_15206,N_15063,N_15158);
nor U15207 (N_15207,N_15092,N_15052);
nor U15208 (N_15208,N_15180,N_15058);
or U15209 (N_15209,N_15001,N_15041);
nor U15210 (N_15210,N_15006,N_15147);
nand U15211 (N_15211,N_15094,N_15068);
nor U15212 (N_15212,N_15136,N_15011);
xor U15213 (N_15213,N_15165,N_15049);
xor U15214 (N_15214,N_15072,N_15083);
nand U15215 (N_15215,N_15185,N_15095);
nand U15216 (N_15216,N_15122,N_15118);
or U15217 (N_15217,N_15054,N_15076);
and U15218 (N_15218,N_15101,N_15197);
and U15219 (N_15219,N_15007,N_15009);
or U15220 (N_15220,N_15157,N_15023);
and U15221 (N_15221,N_15039,N_15126);
nor U15222 (N_15222,N_15152,N_15074);
nor U15223 (N_15223,N_15169,N_15191);
nor U15224 (N_15224,N_15102,N_15008);
nand U15225 (N_15225,N_15056,N_15035);
xor U15226 (N_15226,N_15080,N_15077);
nor U15227 (N_15227,N_15161,N_15159);
or U15228 (N_15228,N_15186,N_15098);
or U15229 (N_15229,N_15110,N_15106);
or U15230 (N_15230,N_15189,N_15132);
and U15231 (N_15231,N_15034,N_15002);
nand U15232 (N_15232,N_15016,N_15019);
nand U15233 (N_15233,N_15040,N_15162);
xnor U15234 (N_15234,N_15178,N_15060);
nand U15235 (N_15235,N_15127,N_15099);
nor U15236 (N_15236,N_15140,N_15048);
or U15237 (N_15237,N_15143,N_15051);
nand U15238 (N_15238,N_15091,N_15031);
xnor U15239 (N_15239,N_15112,N_15081);
and U15240 (N_15240,N_15117,N_15199);
xor U15241 (N_15241,N_15107,N_15004);
xor U15242 (N_15242,N_15075,N_15037);
or U15243 (N_15243,N_15193,N_15082);
nand U15244 (N_15244,N_15172,N_15070);
or U15245 (N_15245,N_15105,N_15196);
nand U15246 (N_15246,N_15130,N_15057);
xor U15247 (N_15247,N_15046,N_15043);
xnor U15248 (N_15248,N_15171,N_15028);
xnor U15249 (N_15249,N_15167,N_15022);
nand U15250 (N_15250,N_15124,N_15164);
or U15251 (N_15251,N_15156,N_15088);
nor U15252 (N_15252,N_15087,N_15062);
or U15253 (N_15253,N_15050,N_15097);
nand U15254 (N_15254,N_15129,N_15145);
and U15255 (N_15255,N_15067,N_15079);
nor U15256 (N_15256,N_15181,N_15150);
or U15257 (N_15257,N_15086,N_15138);
or U15258 (N_15258,N_15141,N_15078);
xor U15259 (N_15259,N_15155,N_15175);
nand U15260 (N_15260,N_15071,N_15000);
or U15261 (N_15261,N_15036,N_15120);
or U15262 (N_15262,N_15137,N_15133);
and U15263 (N_15263,N_15030,N_15115);
or U15264 (N_15264,N_15025,N_15198);
nor U15265 (N_15265,N_15182,N_15044);
and U15266 (N_15266,N_15192,N_15184);
or U15267 (N_15267,N_15012,N_15065);
nand U15268 (N_15268,N_15123,N_15038);
and U15269 (N_15269,N_15174,N_15109);
nor U15270 (N_15270,N_15055,N_15125);
and U15271 (N_15271,N_15017,N_15170);
nand U15272 (N_15272,N_15154,N_15146);
or U15273 (N_15273,N_15177,N_15032);
nor U15274 (N_15274,N_15047,N_15149);
xnor U15275 (N_15275,N_15108,N_15173);
nand U15276 (N_15276,N_15026,N_15093);
nor U15277 (N_15277,N_15024,N_15128);
and U15278 (N_15278,N_15168,N_15166);
or U15279 (N_15279,N_15021,N_15194);
xor U15280 (N_15280,N_15015,N_15163);
nand U15281 (N_15281,N_15148,N_15066);
nor U15282 (N_15282,N_15183,N_15131);
or U15283 (N_15283,N_15176,N_15085);
and U15284 (N_15284,N_15045,N_15084);
nor U15285 (N_15285,N_15195,N_15151);
or U15286 (N_15286,N_15103,N_15073);
or U15287 (N_15287,N_15010,N_15188);
xnor U15288 (N_15288,N_15135,N_15114);
xor U15289 (N_15289,N_15113,N_15153);
xnor U15290 (N_15290,N_15020,N_15089);
nand U15291 (N_15291,N_15139,N_15059);
xor U15292 (N_15292,N_15100,N_15111);
nor U15293 (N_15293,N_15061,N_15096);
or U15294 (N_15294,N_15142,N_15119);
xor U15295 (N_15295,N_15090,N_15160);
xnor U15296 (N_15296,N_15018,N_15013);
xnor U15297 (N_15297,N_15014,N_15064);
nor U15298 (N_15298,N_15005,N_15144);
nor U15299 (N_15299,N_15003,N_15134);
nor U15300 (N_15300,N_15042,N_15182);
and U15301 (N_15301,N_15188,N_15165);
or U15302 (N_15302,N_15095,N_15093);
and U15303 (N_15303,N_15182,N_15120);
nand U15304 (N_15304,N_15097,N_15077);
nand U15305 (N_15305,N_15076,N_15027);
nand U15306 (N_15306,N_15112,N_15072);
nand U15307 (N_15307,N_15154,N_15061);
and U15308 (N_15308,N_15195,N_15053);
nand U15309 (N_15309,N_15051,N_15081);
xnor U15310 (N_15310,N_15096,N_15093);
and U15311 (N_15311,N_15090,N_15167);
or U15312 (N_15312,N_15006,N_15066);
and U15313 (N_15313,N_15084,N_15021);
and U15314 (N_15314,N_15027,N_15173);
nor U15315 (N_15315,N_15187,N_15111);
and U15316 (N_15316,N_15027,N_15095);
xor U15317 (N_15317,N_15190,N_15085);
xnor U15318 (N_15318,N_15169,N_15195);
and U15319 (N_15319,N_15172,N_15169);
nor U15320 (N_15320,N_15000,N_15141);
nor U15321 (N_15321,N_15161,N_15123);
xor U15322 (N_15322,N_15170,N_15147);
and U15323 (N_15323,N_15082,N_15067);
or U15324 (N_15324,N_15085,N_15100);
and U15325 (N_15325,N_15021,N_15022);
and U15326 (N_15326,N_15077,N_15123);
xor U15327 (N_15327,N_15058,N_15116);
nor U15328 (N_15328,N_15093,N_15047);
nor U15329 (N_15329,N_15069,N_15100);
nor U15330 (N_15330,N_15184,N_15157);
nor U15331 (N_15331,N_15127,N_15070);
or U15332 (N_15332,N_15040,N_15036);
nand U15333 (N_15333,N_15092,N_15048);
or U15334 (N_15334,N_15005,N_15060);
or U15335 (N_15335,N_15184,N_15191);
xor U15336 (N_15336,N_15048,N_15147);
or U15337 (N_15337,N_15170,N_15099);
nand U15338 (N_15338,N_15046,N_15130);
or U15339 (N_15339,N_15017,N_15131);
nand U15340 (N_15340,N_15035,N_15054);
nand U15341 (N_15341,N_15158,N_15182);
nor U15342 (N_15342,N_15124,N_15017);
or U15343 (N_15343,N_15125,N_15148);
and U15344 (N_15344,N_15131,N_15169);
nor U15345 (N_15345,N_15131,N_15046);
or U15346 (N_15346,N_15105,N_15182);
xor U15347 (N_15347,N_15133,N_15062);
and U15348 (N_15348,N_15169,N_15040);
or U15349 (N_15349,N_15156,N_15115);
or U15350 (N_15350,N_15188,N_15186);
xnor U15351 (N_15351,N_15013,N_15177);
nand U15352 (N_15352,N_15199,N_15028);
nor U15353 (N_15353,N_15141,N_15084);
nand U15354 (N_15354,N_15107,N_15028);
nor U15355 (N_15355,N_15190,N_15134);
xor U15356 (N_15356,N_15162,N_15150);
or U15357 (N_15357,N_15044,N_15057);
xor U15358 (N_15358,N_15005,N_15027);
nor U15359 (N_15359,N_15013,N_15098);
xnor U15360 (N_15360,N_15043,N_15169);
nand U15361 (N_15361,N_15064,N_15099);
nor U15362 (N_15362,N_15165,N_15053);
nand U15363 (N_15363,N_15041,N_15016);
or U15364 (N_15364,N_15091,N_15094);
nor U15365 (N_15365,N_15065,N_15061);
or U15366 (N_15366,N_15163,N_15141);
and U15367 (N_15367,N_15190,N_15162);
xnor U15368 (N_15368,N_15008,N_15078);
xnor U15369 (N_15369,N_15027,N_15044);
xnor U15370 (N_15370,N_15157,N_15009);
nand U15371 (N_15371,N_15074,N_15001);
and U15372 (N_15372,N_15046,N_15052);
nor U15373 (N_15373,N_15060,N_15013);
or U15374 (N_15374,N_15150,N_15102);
nand U15375 (N_15375,N_15109,N_15000);
nor U15376 (N_15376,N_15142,N_15189);
and U15377 (N_15377,N_15039,N_15097);
and U15378 (N_15378,N_15109,N_15175);
nor U15379 (N_15379,N_15110,N_15153);
nor U15380 (N_15380,N_15013,N_15031);
and U15381 (N_15381,N_15022,N_15110);
and U15382 (N_15382,N_15125,N_15121);
nand U15383 (N_15383,N_15048,N_15049);
nor U15384 (N_15384,N_15047,N_15071);
nor U15385 (N_15385,N_15093,N_15181);
or U15386 (N_15386,N_15053,N_15010);
nand U15387 (N_15387,N_15141,N_15104);
xor U15388 (N_15388,N_15167,N_15051);
or U15389 (N_15389,N_15149,N_15160);
nor U15390 (N_15390,N_15100,N_15182);
xor U15391 (N_15391,N_15104,N_15081);
or U15392 (N_15392,N_15095,N_15144);
and U15393 (N_15393,N_15064,N_15018);
nand U15394 (N_15394,N_15144,N_15056);
or U15395 (N_15395,N_15185,N_15001);
or U15396 (N_15396,N_15119,N_15109);
and U15397 (N_15397,N_15000,N_15099);
nor U15398 (N_15398,N_15071,N_15017);
nand U15399 (N_15399,N_15101,N_15180);
xnor U15400 (N_15400,N_15331,N_15250);
xor U15401 (N_15401,N_15273,N_15260);
or U15402 (N_15402,N_15336,N_15258);
nor U15403 (N_15403,N_15209,N_15298);
xor U15404 (N_15404,N_15243,N_15281);
xnor U15405 (N_15405,N_15374,N_15329);
xor U15406 (N_15406,N_15236,N_15399);
and U15407 (N_15407,N_15254,N_15289);
or U15408 (N_15408,N_15299,N_15391);
nor U15409 (N_15409,N_15245,N_15381);
and U15410 (N_15410,N_15338,N_15208);
xor U15411 (N_15411,N_15388,N_15327);
nor U15412 (N_15412,N_15382,N_15385);
nand U15413 (N_15413,N_15353,N_15351);
or U15414 (N_15414,N_15300,N_15350);
or U15415 (N_15415,N_15359,N_15200);
or U15416 (N_15416,N_15397,N_15277);
nand U15417 (N_15417,N_15288,N_15270);
or U15418 (N_15418,N_15274,N_15257);
or U15419 (N_15419,N_15237,N_15312);
and U15420 (N_15420,N_15223,N_15384);
xnor U15421 (N_15421,N_15287,N_15364);
nor U15422 (N_15422,N_15361,N_15335);
nand U15423 (N_15423,N_15240,N_15305);
or U15424 (N_15424,N_15217,N_15314);
nor U15425 (N_15425,N_15292,N_15318);
and U15426 (N_15426,N_15230,N_15275);
and U15427 (N_15427,N_15326,N_15249);
and U15428 (N_15428,N_15328,N_15310);
or U15429 (N_15429,N_15233,N_15222);
nand U15430 (N_15430,N_15206,N_15221);
xnor U15431 (N_15431,N_15271,N_15235);
or U15432 (N_15432,N_15358,N_15239);
xor U15433 (N_15433,N_15316,N_15301);
or U15434 (N_15434,N_15317,N_15255);
or U15435 (N_15435,N_15205,N_15283);
xnor U15436 (N_15436,N_15356,N_15296);
nor U15437 (N_15437,N_15313,N_15337);
xnor U15438 (N_15438,N_15349,N_15380);
or U15439 (N_15439,N_15308,N_15248);
nor U15440 (N_15440,N_15263,N_15398);
nand U15441 (N_15441,N_15393,N_15212);
and U15442 (N_15442,N_15238,N_15319);
xor U15443 (N_15443,N_15341,N_15268);
nor U15444 (N_15444,N_15311,N_15363);
and U15445 (N_15445,N_15383,N_15365);
nor U15446 (N_15446,N_15378,N_15355);
nand U15447 (N_15447,N_15219,N_15323);
nor U15448 (N_15448,N_15272,N_15278);
nand U15449 (N_15449,N_15247,N_15321);
nand U15450 (N_15450,N_15213,N_15322);
and U15451 (N_15451,N_15246,N_15203);
xnor U15452 (N_15452,N_15259,N_15377);
xor U15453 (N_15453,N_15231,N_15396);
nand U15454 (N_15454,N_15309,N_15252);
and U15455 (N_15455,N_15343,N_15304);
xor U15456 (N_15456,N_15261,N_15346);
and U15457 (N_15457,N_15370,N_15229);
or U15458 (N_15458,N_15285,N_15348);
nor U15459 (N_15459,N_15211,N_15303);
or U15460 (N_15460,N_15280,N_15286);
and U15461 (N_15461,N_15387,N_15215);
xnor U15462 (N_15462,N_15375,N_15357);
xor U15463 (N_15463,N_15306,N_15395);
and U15464 (N_15464,N_15244,N_15201);
nor U15465 (N_15465,N_15251,N_15389);
nand U15466 (N_15466,N_15372,N_15207);
and U15467 (N_15467,N_15315,N_15220);
and U15468 (N_15468,N_15394,N_15373);
nor U15469 (N_15469,N_15264,N_15392);
nor U15470 (N_15470,N_15291,N_15227);
xnor U15471 (N_15471,N_15262,N_15347);
and U15472 (N_15472,N_15371,N_15269);
nand U15473 (N_15473,N_15307,N_15294);
xnor U15474 (N_15474,N_15390,N_15276);
or U15475 (N_15475,N_15228,N_15225);
nor U15476 (N_15476,N_15345,N_15256);
nor U15477 (N_15477,N_15342,N_15325);
nand U15478 (N_15478,N_15210,N_15368);
xnor U15479 (N_15479,N_15352,N_15360);
xor U15480 (N_15480,N_15265,N_15330);
or U15481 (N_15481,N_15295,N_15204);
nand U15482 (N_15482,N_15297,N_15354);
xor U15483 (N_15483,N_15293,N_15216);
or U15484 (N_15484,N_15284,N_15242);
or U15485 (N_15485,N_15214,N_15320);
xnor U15486 (N_15486,N_15362,N_15279);
nand U15487 (N_15487,N_15376,N_15332);
xnor U15488 (N_15488,N_15282,N_15340);
nand U15489 (N_15489,N_15333,N_15218);
or U15490 (N_15490,N_15369,N_15344);
or U15491 (N_15491,N_15267,N_15226);
xnor U15492 (N_15492,N_15234,N_15232);
nand U15493 (N_15493,N_15339,N_15224);
and U15494 (N_15494,N_15202,N_15379);
nor U15495 (N_15495,N_15302,N_15367);
or U15496 (N_15496,N_15324,N_15241);
or U15497 (N_15497,N_15266,N_15334);
nand U15498 (N_15498,N_15366,N_15386);
and U15499 (N_15499,N_15290,N_15253);
nand U15500 (N_15500,N_15264,N_15395);
xor U15501 (N_15501,N_15250,N_15214);
nand U15502 (N_15502,N_15213,N_15247);
xor U15503 (N_15503,N_15204,N_15283);
xnor U15504 (N_15504,N_15343,N_15253);
nor U15505 (N_15505,N_15344,N_15229);
nor U15506 (N_15506,N_15386,N_15254);
or U15507 (N_15507,N_15347,N_15373);
xor U15508 (N_15508,N_15259,N_15274);
or U15509 (N_15509,N_15227,N_15326);
or U15510 (N_15510,N_15342,N_15270);
xnor U15511 (N_15511,N_15374,N_15380);
nor U15512 (N_15512,N_15396,N_15356);
nand U15513 (N_15513,N_15282,N_15240);
or U15514 (N_15514,N_15206,N_15346);
nor U15515 (N_15515,N_15351,N_15221);
and U15516 (N_15516,N_15302,N_15377);
nand U15517 (N_15517,N_15293,N_15396);
nor U15518 (N_15518,N_15365,N_15309);
and U15519 (N_15519,N_15346,N_15310);
xor U15520 (N_15520,N_15273,N_15361);
nand U15521 (N_15521,N_15283,N_15324);
xor U15522 (N_15522,N_15267,N_15330);
and U15523 (N_15523,N_15357,N_15334);
nor U15524 (N_15524,N_15359,N_15373);
xnor U15525 (N_15525,N_15362,N_15249);
nor U15526 (N_15526,N_15242,N_15373);
or U15527 (N_15527,N_15200,N_15209);
and U15528 (N_15528,N_15225,N_15290);
and U15529 (N_15529,N_15302,N_15220);
xor U15530 (N_15530,N_15210,N_15245);
or U15531 (N_15531,N_15375,N_15206);
nor U15532 (N_15532,N_15227,N_15211);
xnor U15533 (N_15533,N_15276,N_15320);
xor U15534 (N_15534,N_15257,N_15361);
nor U15535 (N_15535,N_15339,N_15265);
nand U15536 (N_15536,N_15297,N_15248);
and U15537 (N_15537,N_15229,N_15202);
and U15538 (N_15538,N_15310,N_15313);
xnor U15539 (N_15539,N_15377,N_15364);
nand U15540 (N_15540,N_15207,N_15266);
and U15541 (N_15541,N_15242,N_15388);
or U15542 (N_15542,N_15212,N_15368);
nand U15543 (N_15543,N_15312,N_15309);
nand U15544 (N_15544,N_15289,N_15247);
nand U15545 (N_15545,N_15243,N_15297);
or U15546 (N_15546,N_15356,N_15209);
nand U15547 (N_15547,N_15232,N_15366);
nor U15548 (N_15548,N_15266,N_15368);
nand U15549 (N_15549,N_15372,N_15373);
and U15550 (N_15550,N_15323,N_15319);
or U15551 (N_15551,N_15392,N_15270);
or U15552 (N_15552,N_15376,N_15238);
nand U15553 (N_15553,N_15287,N_15320);
or U15554 (N_15554,N_15252,N_15232);
nor U15555 (N_15555,N_15248,N_15342);
and U15556 (N_15556,N_15366,N_15293);
nor U15557 (N_15557,N_15362,N_15396);
nand U15558 (N_15558,N_15368,N_15268);
nand U15559 (N_15559,N_15260,N_15201);
nor U15560 (N_15560,N_15285,N_15280);
xor U15561 (N_15561,N_15394,N_15282);
and U15562 (N_15562,N_15341,N_15308);
nand U15563 (N_15563,N_15299,N_15273);
nor U15564 (N_15564,N_15317,N_15387);
or U15565 (N_15565,N_15329,N_15398);
or U15566 (N_15566,N_15386,N_15307);
and U15567 (N_15567,N_15206,N_15272);
and U15568 (N_15568,N_15275,N_15300);
nor U15569 (N_15569,N_15381,N_15259);
or U15570 (N_15570,N_15373,N_15367);
nand U15571 (N_15571,N_15227,N_15379);
nand U15572 (N_15572,N_15333,N_15383);
xnor U15573 (N_15573,N_15258,N_15293);
or U15574 (N_15574,N_15287,N_15288);
nor U15575 (N_15575,N_15228,N_15290);
nor U15576 (N_15576,N_15325,N_15298);
nand U15577 (N_15577,N_15203,N_15251);
or U15578 (N_15578,N_15255,N_15332);
or U15579 (N_15579,N_15323,N_15285);
xnor U15580 (N_15580,N_15302,N_15232);
xnor U15581 (N_15581,N_15216,N_15295);
nor U15582 (N_15582,N_15217,N_15205);
nor U15583 (N_15583,N_15266,N_15238);
and U15584 (N_15584,N_15377,N_15202);
nor U15585 (N_15585,N_15253,N_15263);
nand U15586 (N_15586,N_15301,N_15305);
nand U15587 (N_15587,N_15295,N_15217);
xor U15588 (N_15588,N_15352,N_15340);
nand U15589 (N_15589,N_15265,N_15257);
and U15590 (N_15590,N_15291,N_15336);
and U15591 (N_15591,N_15286,N_15333);
xnor U15592 (N_15592,N_15262,N_15227);
and U15593 (N_15593,N_15385,N_15396);
nor U15594 (N_15594,N_15362,N_15381);
nor U15595 (N_15595,N_15246,N_15325);
nor U15596 (N_15596,N_15345,N_15355);
or U15597 (N_15597,N_15305,N_15229);
or U15598 (N_15598,N_15364,N_15222);
nor U15599 (N_15599,N_15291,N_15387);
and U15600 (N_15600,N_15596,N_15452);
nand U15601 (N_15601,N_15581,N_15592);
nand U15602 (N_15602,N_15563,N_15540);
xnor U15603 (N_15603,N_15492,N_15516);
xnor U15604 (N_15604,N_15580,N_15593);
xor U15605 (N_15605,N_15579,N_15577);
or U15606 (N_15606,N_15423,N_15460);
or U15607 (N_15607,N_15408,N_15539);
nor U15608 (N_15608,N_15464,N_15517);
and U15609 (N_15609,N_15471,N_15424);
nor U15610 (N_15610,N_15439,N_15551);
nand U15611 (N_15611,N_15533,N_15448);
nand U15612 (N_15612,N_15590,N_15473);
and U15613 (N_15613,N_15537,N_15582);
or U15614 (N_15614,N_15422,N_15559);
xnor U15615 (N_15615,N_15466,N_15586);
or U15616 (N_15616,N_15576,N_15558);
xnor U15617 (N_15617,N_15525,N_15567);
nand U15618 (N_15618,N_15481,N_15402);
nand U15619 (N_15619,N_15434,N_15445);
and U15620 (N_15620,N_15534,N_15485);
and U15621 (N_15621,N_15440,N_15479);
nand U15622 (N_15622,N_15429,N_15511);
nor U15623 (N_15623,N_15588,N_15500);
and U15624 (N_15624,N_15411,N_15414);
nand U15625 (N_15625,N_15453,N_15510);
nor U15626 (N_15626,N_15556,N_15483);
xor U15627 (N_15627,N_15497,N_15566);
and U15628 (N_15628,N_15515,N_15431);
xnor U15629 (N_15629,N_15527,N_15589);
nor U15630 (N_15630,N_15405,N_15409);
nor U15631 (N_15631,N_15501,N_15450);
nor U15632 (N_15632,N_15412,N_15542);
xor U15633 (N_15633,N_15503,N_15532);
nor U15634 (N_15634,N_15410,N_15570);
nand U15635 (N_15635,N_15462,N_15508);
xor U15636 (N_15636,N_15461,N_15564);
or U15637 (N_15637,N_15530,N_15430);
nor U15638 (N_15638,N_15478,N_15528);
nor U15639 (N_15639,N_15421,N_15502);
nor U15640 (N_15640,N_15488,N_15513);
and U15641 (N_15641,N_15544,N_15472);
nand U15642 (N_15642,N_15569,N_15561);
nor U15643 (N_15643,N_15490,N_15543);
or U15644 (N_15644,N_15442,N_15444);
and U15645 (N_15645,N_15523,N_15529);
xor U15646 (N_15646,N_15451,N_15443);
or U15647 (N_15647,N_15499,N_15557);
or U15648 (N_15648,N_15403,N_15416);
nor U15649 (N_15649,N_15417,N_15521);
and U15650 (N_15650,N_15477,N_15489);
xnor U15651 (N_15651,N_15415,N_15420);
nand U15652 (N_15652,N_15495,N_15549);
xnor U15653 (N_15653,N_15531,N_15512);
nor U15654 (N_15654,N_15433,N_15463);
or U15655 (N_15655,N_15470,N_15419);
or U15656 (N_15656,N_15524,N_15468);
nor U15657 (N_15657,N_15587,N_15550);
xnor U15658 (N_15658,N_15484,N_15455);
xnor U15659 (N_15659,N_15400,N_15555);
nand U15660 (N_15660,N_15475,N_15506);
nand U15661 (N_15661,N_15572,N_15546);
xnor U15662 (N_15662,N_15432,N_15595);
nand U15663 (N_15663,N_15599,N_15449);
xor U15664 (N_15664,N_15426,N_15487);
nor U15665 (N_15665,N_15560,N_15552);
nor U15666 (N_15666,N_15562,N_15573);
xor U15667 (N_15667,N_15456,N_15597);
and U15668 (N_15668,N_15418,N_15526);
nand U15669 (N_15669,N_15437,N_15575);
nor U15670 (N_15670,N_15553,N_15520);
nand U15671 (N_15671,N_15585,N_15574);
nor U15672 (N_15672,N_15457,N_15482);
or U15673 (N_15673,N_15404,N_15441);
and U15674 (N_15674,N_15413,N_15438);
xor U15675 (N_15675,N_15446,N_15436);
nand U15676 (N_15676,N_15476,N_15514);
or U15677 (N_15677,N_15459,N_15493);
or U15678 (N_15678,N_15594,N_15598);
nand U15679 (N_15679,N_15498,N_15507);
or U15680 (N_15680,N_15427,N_15522);
nand U15681 (N_15681,N_15494,N_15518);
and U15682 (N_15682,N_15535,N_15474);
xnor U15683 (N_15683,N_15583,N_15565);
xnor U15684 (N_15684,N_15584,N_15545);
xor U15685 (N_15685,N_15407,N_15465);
xor U15686 (N_15686,N_15548,N_15496);
nor U15687 (N_15687,N_15547,N_15509);
nor U15688 (N_15688,N_15428,N_15541);
or U15689 (N_15689,N_15536,N_15454);
or U15690 (N_15690,N_15467,N_15406);
xor U15691 (N_15691,N_15435,N_15554);
nand U15692 (N_15692,N_15447,N_15486);
xnor U15693 (N_15693,N_15504,N_15578);
and U15694 (N_15694,N_15571,N_15519);
nand U15695 (N_15695,N_15505,N_15480);
nor U15696 (N_15696,N_15538,N_15469);
or U15697 (N_15697,N_15401,N_15491);
xor U15698 (N_15698,N_15458,N_15425);
or U15699 (N_15699,N_15568,N_15591);
or U15700 (N_15700,N_15414,N_15484);
and U15701 (N_15701,N_15487,N_15480);
nand U15702 (N_15702,N_15445,N_15522);
or U15703 (N_15703,N_15524,N_15586);
nand U15704 (N_15704,N_15461,N_15549);
nor U15705 (N_15705,N_15516,N_15544);
nor U15706 (N_15706,N_15450,N_15428);
nand U15707 (N_15707,N_15508,N_15527);
or U15708 (N_15708,N_15549,N_15575);
xor U15709 (N_15709,N_15552,N_15553);
and U15710 (N_15710,N_15535,N_15412);
xor U15711 (N_15711,N_15408,N_15416);
nand U15712 (N_15712,N_15435,N_15599);
nand U15713 (N_15713,N_15538,N_15550);
nand U15714 (N_15714,N_15437,N_15529);
and U15715 (N_15715,N_15585,N_15598);
nand U15716 (N_15716,N_15514,N_15409);
nor U15717 (N_15717,N_15540,N_15468);
and U15718 (N_15718,N_15572,N_15582);
nand U15719 (N_15719,N_15593,N_15555);
or U15720 (N_15720,N_15486,N_15591);
or U15721 (N_15721,N_15488,N_15464);
or U15722 (N_15722,N_15544,N_15596);
and U15723 (N_15723,N_15470,N_15423);
or U15724 (N_15724,N_15444,N_15465);
nand U15725 (N_15725,N_15571,N_15513);
nand U15726 (N_15726,N_15576,N_15419);
and U15727 (N_15727,N_15536,N_15461);
nor U15728 (N_15728,N_15554,N_15491);
xnor U15729 (N_15729,N_15552,N_15565);
and U15730 (N_15730,N_15537,N_15485);
xnor U15731 (N_15731,N_15554,N_15477);
and U15732 (N_15732,N_15594,N_15543);
or U15733 (N_15733,N_15448,N_15446);
nor U15734 (N_15734,N_15531,N_15548);
or U15735 (N_15735,N_15520,N_15544);
or U15736 (N_15736,N_15410,N_15583);
xor U15737 (N_15737,N_15479,N_15445);
and U15738 (N_15738,N_15435,N_15421);
nand U15739 (N_15739,N_15513,N_15521);
nor U15740 (N_15740,N_15491,N_15570);
nor U15741 (N_15741,N_15556,N_15514);
and U15742 (N_15742,N_15401,N_15518);
or U15743 (N_15743,N_15408,N_15574);
or U15744 (N_15744,N_15467,N_15577);
xor U15745 (N_15745,N_15466,N_15573);
nor U15746 (N_15746,N_15452,N_15597);
xnor U15747 (N_15747,N_15509,N_15562);
nand U15748 (N_15748,N_15462,N_15594);
nand U15749 (N_15749,N_15464,N_15436);
xor U15750 (N_15750,N_15469,N_15425);
nand U15751 (N_15751,N_15448,N_15575);
nand U15752 (N_15752,N_15415,N_15471);
nand U15753 (N_15753,N_15448,N_15478);
nor U15754 (N_15754,N_15517,N_15500);
nor U15755 (N_15755,N_15579,N_15438);
and U15756 (N_15756,N_15578,N_15529);
or U15757 (N_15757,N_15465,N_15448);
xnor U15758 (N_15758,N_15481,N_15532);
and U15759 (N_15759,N_15529,N_15420);
xnor U15760 (N_15760,N_15572,N_15541);
nand U15761 (N_15761,N_15483,N_15465);
or U15762 (N_15762,N_15493,N_15495);
nor U15763 (N_15763,N_15490,N_15584);
nor U15764 (N_15764,N_15435,N_15583);
or U15765 (N_15765,N_15541,N_15469);
xnor U15766 (N_15766,N_15453,N_15433);
nor U15767 (N_15767,N_15460,N_15421);
nor U15768 (N_15768,N_15483,N_15504);
xnor U15769 (N_15769,N_15482,N_15442);
xnor U15770 (N_15770,N_15569,N_15447);
xor U15771 (N_15771,N_15400,N_15531);
xnor U15772 (N_15772,N_15573,N_15436);
xnor U15773 (N_15773,N_15519,N_15497);
and U15774 (N_15774,N_15473,N_15401);
or U15775 (N_15775,N_15549,N_15455);
and U15776 (N_15776,N_15467,N_15487);
or U15777 (N_15777,N_15540,N_15422);
or U15778 (N_15778,N_15529,N_15570);
or U15779 (N_15779,N_15424,N_15513);
nand U15780 (N_15780,N_15474,N_15543);
nor U15781 (N_15781,N_15496,N_15578);
nand U15782 (N_15782,N_15516,N_15496);
nor U15783 (N_15783,N_15505,N_15523);
xnor U15784 (N_15784,N_15578,N_15462);
or U15785 (N_15785,N_15412,N_15476);
nor U15786 (N_15786,N_15430,N_15499);
xor U15787 (N_15787,N_15528,N_15547);
nand U15788 (N_15788,N_15534,N_15557);
nor U15789 (N_15789,N_15591,N_15411);
or U15790 (N_15790,N_15486,N_15540);
and U15791 (N_15791,N_15548,N_15475);
nand U15792 (N_15792,N_15592,N_15406);
and U15793 (N_15793,N_15558,N_15516);
nand U15794 (N_15794,N_15401,N_15535);
or U15795 (N_15795,N_15419,N_15403);
or U15796 (N_15796,N_15435,N_15430);
xor U15797 (N_15797,N_15536,N_15427);
xor U15798 (N_15798,N_15433,N_15460);
nor U15799 (N_15799,N_15472,N_15571);
or U15800 (N_15800,N_15732,N_15770);
nand U15801 (N_15801,N_15675,N_15775);
nor U15802 (N_15802,N_15793,N_15665);
xor U15803 (N_15803,N_15714,N_15625);
nor U15804 (N_15804,N_15631,N_15605);
xor U15805 (N_15805,N_15673,N_15649);
nand U15806 (N_15806,N_15730,N_15710);
nor U15807 (N_15807,N_15725,N_15738);
nor U15808 (N_15808,N_15771,N_15691);
and U15809 (N_15809,N_15777,N_15769);
and U15810 (N_15810,N_15661,N_15653);
nand U15811 (N_15811,N_15729,N_15646);
nand U15812 (N_15812,N_15623,N_15648);
nand U15813 (N_15813,N_15606,N_15633);
nand U15814 (N_15814,N_15600,N_15620);
xor U15815 (N_15815,N_15754,N_15756);
xor U15816 (N_15816,N_15604,N_15684);
and U15817 (N_15817,N_15702,N_15690);
nand U15818 (N_15818,N_15635,N_15723);
or U15819 (N_15819,N_15750,N_15626);
xor U15820 (N_15820,N_15644,N_15681);
and U15821 (N_15821,N_15790,N_15632);
and U15822 (N_15822,N_15615,N_15784);
and U15823 (N_15823,N_15656,N_15658);
nor U15824 (N_15824,N_15664,N_15694);
or U15825 (N_15825,N_15707,N_15613);
nor U15826 (N_15826,N_15634,N_15772);
nand U15827 (N_15827,N_15671,N_15679);
and U15828 (N_15828,N_15715,N_15741);
nand U15829 (N_15829,N_15652,N_15650);
nand U15830 (N_15830,N_15795,N_15787);
nand U15831 (N_15831,N_15689,N_15651);
xnor U15832 (N_15832,N_15753,N_15767);
nand U15833 (N_15833,N_15735,N_15686);
nand U15834 (N_15834,N_15642,N_15751);
nor U15835 (N_15835,N_15726,N_15603);
nor U15836 (N_15836,N_15724,N_15697);
or U15837 (N_15837,N_15641,N_15739);
nor U15838 (N_15838,N_15695,N_15657);
or U15839 (N_15839,N_15781,N_15701);
nor U15840 (N_15840,N_15668,N_15779);
xnor U15841 (N_15841,N_15737,N_15733);
xnor U15842 (N_15842,N_15610,N_15749);
and U15843 (N_15843,N_15709,N_15745);
xnor U15844 (N_15844,N_15748,N_15674);
nand U15845 (N_15845,N_15744,N_15677);
and U15846 (N_15846,N_15612,N_15663);
or U15847 (N_15847,N_15743,N_15609);
nor U15848 (N_15848,N_15616,N_15682);
nor U15849 (N_15849,N_15768,N_15788);
and U15850 (N_15850,N_15676,N_15667);
nand U15851 (N_15851,N_15624,N_15778);
nand U15852 (N_15852,N_15621,N_15706);
and U15853 (N_15853,N_15708,N_15692);
xor U15854 (N_15854,N_15766,N_15740);
and U15855 (N_15855,N_15782,N_15672);
xor U15856 (N_15856,N_15601,N_15762);
and U15857 (N_15857,N_15617,N_15742);
or U15858 (N_15858,N_15629,N_15719);
nor U15859 (N_15859,N_15713,N_15602);
and U15860 (N_15860,N_15796,N_15699);
and U15861 (N_15861,N_15680,N_15660);
or U15862 (N_15862,N_15761,N_15608);
nor U15863 (N_15863,N_15718,N_15627);
and U15864 (N_15864,N_15637,N_15786);
nor U15865 (N_15865,N_15776,N_15734);
xor U15866 (N_15866,N_15678,N_15797);
xnor U15867 (N_15867,N_15764,N_15638);
nand U15868 (N_15868,N_15711,N_15727);
or U15869 (N_15869,N_15666,N_15628);
nor U15870 (N_15870,N_15611,N_15654);
xor U15871 (N_15871,N_15789,N_15645);
or U15872 (N_15872,N_15792,N_15722);
nor U15873 (N_15873,N_15791,N_15763);
nand U15874 (N_15874,N_15655,N_15758);
nand U15875 (N_15875,N_15705,N_15636);
xor U15876 (N_15876,N_15712,N_15798);
or U15877 (N_15877,N_15752,N_15747);
or U15878 (N_15878,N_15783,N_15659);
nor U15879 (N_15879,N_15780,N_15728);
and U15880 (N_15880,N_15703,N_15696);
nor U15881 (N_15881,N_15759,N_15607);
nor U15882 (N_15882,N_15794,N_15755);
xor U15883 (N_15883,N_15746,N_15785);
or U15884 (N_15884,N_15716,N_15717);
nand U15885 (N_15885,N_15639,N_15720);
nand U15886 (N_15886,N_15700,N_15619);
nor U15887 (N_15887,N_15731,N_15662);
xor U15888 (N_15888,N_15622,N_15773);
xor U15889 (N_15889,N_15698,N_15643);
nor U15890 (N_15890,N_15799,N_15688);
nor U15891 (N_15891,N_15640,N_15760);
xnor U15892 (N_15892,N_15614,N_15670);
and U15893 (N_15893,N_15683,N_15693);
or U15894 (N_15894,N_15687,N_15721);
nor U15895 (N_15895,N_15765,N_15704);
nor U15896 (N_15896,N_15774,N_15669);
and U15897 (N_15897,N_15647,N_15736);
and U15898 (N_15898,N_15757,N_15618);
nand U15899 (N_15899,N_15685,N_15630);
nor U15900 (N_15900,N_15713,N_15651);
or U15901 (N_15901,N_15791,N_15605);
nor U15902 (N_15902,N_15787,N_15753);
xor U15903 (N_15903,N_15619,N_15741);
xor U15904 (N_15904,N_15699,N_15771);
or U15905 (N_15905,N_15753,N_15768);
and U15906 (N_15906,N_15702,N_15751);
or U15907 (N_15907,N_15753,N_15617);
or U15908 (N_15908,N_15790,N_15716);
nor U15909 (N_15909,N_15726,N_15677);
and U15910 (N_15910,N_15723,N_15640);
and U15911 (N_15911,N_15609,N_15626);
or U15912 (N_15912,N_15771,N_15714);
or U15913 (N_15913,N_15624,N_15714);
nor U15914 (N_15914,N_15658,N_15745);
nor U15915 (N_15915,N_15663,N_15614);
or U15916 (N_15916,N_15789,N_15695);
xnor U15917 (N_15917,N_15727,N_15626);
or U15918 (N_15918,N_15724,N_15757);
or U15919 (N_15919,N_15694,N_15693);
xor U15920 (N_15920,N_15796,N_15777);
and U15921 (N_15921,N_15706,N_15655);
nand U15922 (N_15922,N_15609,N_15659);
nor U15923 (N_15923,N_15731,N_15637);
and U15924 (N_15924,N_15769,N_15658);
or U15925 (N_15925,N_15677,N_15711);
and U15926 (N_15926,N_15706,N_15794);
or U15927 (N_15927,N_15687,N_15702);
xnor U15928 (N_15928,N_15768,N_15644);
nor U15929 (N_15929,N_15622,N_15626);
nor U15930 (N_15930,N_15666,N_15695);
or U15931 (N_15931,N_15705,N_15689);
xnor U15932 (N_15932,N_15705,N_15758);
xor U15933 (N_15933,N_15620,N_15659);
nand U15934 (N_15934,N_15612,N_15640);
xor U15935 (N_15935,N_15685,N_15760);
or U15936 (N_15936,N_15795,N_15659);
nor U15937 (N_15937,N_15639,N_15669);
nand U15938 (N_15938,N_15791,N_15627);
nand U15939 (N_15939,N_15656,N_15602);
or U15940 (N_15940,N_15745,N_15713);
or U15941 (N_15941,N_15766,N_15646);
or U15942 (N_15942,N_15659,N_15650);
and U15943 (N_15943,N_15612,N_15754);
nand U15944 (N_15944,N_15696,N_15659);
xnor U15945 (N_15945,N_15710,N_15654);
or U15946 (N_15946,N_15666,N_15754);
xor U15947 (N_15947,N_15679,N_15604);
nand U15948 (N_15948,N_15792,N_15704);
nand U15949 (N_15949,N_15651,N_15701);
nand U15950 (N_15950,N_15653,N_15791);
and U15951 (N_15951,N_15790,N_15643);
or U15952 (N_15952,N_15732,N_15711);
and U15953 (N_15953,N_15771,N_15748);
nor U15954 (N_15954,N_15612,N_15695);
or U15955 (N_15955,N_15771,N_15645);
nor U15956 (N_15956,N_15636,N_15713);
nand U15957 (N_15957,N_15606,N_15776);
nand U15958 (N_15958,N_15670,N_15711);
nor U15959 (N_15959,N_15691,N_15696);
xor U15960 (N_15960,N_15694,N_15732);
nand U15961 (N_15961,N_15731,N_15784);
or U15962 (N_15962,N_15784,N_15693);
and U15963 (N_15963,N_15663,N_15725);
nand U15964 (N_15964,N_15608,N_15755);
and U15965 (N_15965,N_15787,N_15633);
nand U15966 (N_15966,N_15740,N_15763);
xnor U15967 (N_15967,N_15630,N_15664);
nor U15968 (N_15968,N_15601,N_15728);
nand U15969 (N_15969,N_15763,N_15753);
nor U15970 (N_15970,N_15640,N_15604);
nand U15971 (N_15971,N_15685,N_15738);
nor U15972 (N_15972,N_15781,N_15742);
xnor U15973 (N_15973,N_15672,N_15753);
xnor U15974 (N_15974,N_15763,N_15755);
nand U15975 (N_15975,N_15762,N_15727);
nor U15976 (N_15976,N_15678,N_15691);
and U15977 (N_15977,N_15725,N_15727);
nand U15978 (N_15978,N_15605,N_15702);
xor U15979 (N_15979,N_15641,N_15686);
xnor U15980 (N_15980,N_15762,N_15625);
nor U15981 (N_15981,N_15670,N_15730);
nor U15982 (N_15982,N_15614,N_15732);
and U15983 (N_15983,N_15707,N_15667);
xnor U15984 (N_15984,N_15731,N_15763);
or U15985 (N_15985,N_15602,N_15740);
nor U15986 (N_15986,N_15601,N_15791);
or U15987 (N_15987,N_15721,N_15743);
nor U15988 (N_15988,N_15685,N_15610);
or U15989 (N_15989,N_15614,N_15665);
xnor U15990 (N_15990,N_15631,N_15792);
nand U15991 (N_15991,N_15742,N_15768);
or U15992 (N_15992,N_15678,N_15656);
and U15993 (N_15993,N_15669,N_15698);
nor U15994 (N_15994,N_15624,N_15701);
or U15995 (N_15995,N_15745,N_15762);
nand U15996 (N_15996,N_15785,N_15772);
nand U15997 (N_15997,N_15668,N_15665);
nor U15998 (N_15998,N_15663,N_15789);
and U15999 (N_15999,N_15773,N_15603);
nor U16000 (N_16000,N_15848,N_15866);
or U16001 (N_16001,N_15860,N_15819);
xnor U16002 (N_16002,N_15878,N_15982);
nand U16003 (N_16003,N_15825,N_15946);
and U16004 (N_16004,N_15869,N_15962);
xnor U16005 (N_16005,N_15986,N_15914);
xor U16006 (N_16006,N_15823,N_15961);
and U16007 (N_16007,N_15892,N_15880);
nor U16008 (N_16008,N_15885,N_15856);
nor U16009 (N_16009,N_15841,N_15971);
nand U16010 (N_16010,N_15909,N_15980);
xor U16011 (N_16011,N_15916,N_15940);
or U16012 (N_16012,N_15922,N_15822);
and U16013 (N_16013,N_15836,N_15824);
or U16014 (N_16014,N_15978,N_15872);
nand U16015 (N_16015,N_15889,N_15847);
nor U16016 (N_16016,N_15907,N_15808);
nor U16017 (N_16017,N_15925,N_15876);
and U16018 (N_16018,N_15842,N_15924);
nand U16019 (N_16019,N_15934,N_15887);
nor U16020 (N_16020,N_15930,N_15953);
xor U16021 (N_16021,N_15806,N_15871);
xor U16022 (N_16022,N_15979,N_15923);
xor U16023 (N_16023,N_15894,N_15919);
xor U16024 (N_16024,N_15843,N_15849);
and U16025 (N_16025,N_15935,N_15938);
or U16026 (N_16026,N_15800,N_15851);
nand U16027 (N_16027,N_15827,N_15968);
or U16028 (N_16028,N_15868,N_15984);
xor U16029 (N_16029,N_15820,N_15890);
nand U16030 (N_16030,N_15973,N_15951);
xor U16031 (N_16031,N_15998,N_15928);
nand U16032 (N_16032,N_15855,N_15918);
and U16033 (N_16033,N_15932,N_15807);
or U16034 (N_16034,N_15942,N_15832);
xnor U16035 (N_16035,N_15969,N_15850);
nor U16036 (N_16036,N_15844,N_15936);
nand U16037 (N_16037,N_15897,N_15939);
nor U16038 (N_16038,N_15944,N_15867);
xnor U16039 (N_16039,N_15983,N_15910);
and U16040 (N_16040,N_15816,N_15839);
nor U16041 (N_16041,N_15877,N_15835);
nor U16042 (N_16042,N_15801,N_15988);
nor U16043 (N_16043,N_15900,N_15927);
and U16044 (N_16044,N_15837,N_15846);
and U16045 (N_16045,N_15821,N_15999);
xnor U16046 (N_16046,N_15882,N_15994);
and U16047 (N_16047,N_15875,N_15828);
nor U16048 (N_16048,N_15865,N_15861);
nor U16049 (N_16049,N_15992,N_15874);
nor U16050 (N_16050,N_15845,N_15985);
nand U16051 (N_16051,N_15854,N_15915);
and U16052 (N_16052,N_15852,N_15802);
xor U16053 (N_16053,N_15960,N_15904);
and U16054 (N_16054,N_15895,N_15929);
and U16055 (N_16055,N_15859,N_15997);
nand U16056 (N_16056,N_15812,N_15931);
xnor U16057 (N_16057,N_15949,N_15972);
xor U16058 (N_16058,N_15886,N_15920);
or U16059 (N_16059,N_15906,N_15809);
nand U16060 (N_16060,N_15834,N_15956);
and U16061 (N_16061,N_15933,N_15977);
nand U16062 (N_16062,N_15950,N_15976);
xnor U16063 (N_16063,N_15975,N_15990);
and U16064 (N_16064,N_15989,N_15921);
xnor U16065 (N_16065,N_15853,N_15838);
or U16066 (N_16066,N_15888,N_15864);
xnor U16067 (N_16067,N_15829,N_15954);
nand U16068 (N_16068,N_15970,N_15857);
nand U16069 (N_16069,N_15805,N_15811);
xnor U16070 (N_16070,N_15967,N_15913);
and U16071 (N_16071,N_15899,N_15858);
and U16072 (N_16072,N_15818,N_15903);
and U16073 (N_16073,N_15898,N_15965);
nand U16074 (N_16074,N_15937,N_15905);
or U16075 (N_16075,N_15879,N_15817);
and U16076 (N_16076,N_15957,N_15948);
and U16077 (N_16077,N_15830,N_15831);
and U16078 (N_16078,N_15981,N_15902);
nand U16079 (N_16079,N_15804,N_15881);
or U16080 (N_16080,N_15952,N_15966);
nand U16081 (N_16081,N_15896,N_15893);
xor U16082 (N_16082,N_15810,N_15943);
or U16083 (N_16083,N_15959,N_15945);
or U16084 (N_16084,N_15840,N_15863);
nand U16085 (N_16085,N_15941,N_15987);
and U16086 (N_16086,N_15995,N_15815);
xor U16087 (N_16087,N_15947,N_15803);
or U16088 (N_16088,N_15991,N_15964);
nor U16089 (N_16089,N_15911,N_15814);
xnor U16090 (N_16090,N_15891,N_15884);
xnor U16091 (N_16091,N_15955,N_15908);
and U16092 (N_16092,N_15901,N_15926);
and U16093 (N_16093,N_15974,N_15813);
nand U16094 (N_16094,N_15883,N_15870);
nand U16095 (N_16095,N_15862,N_15993);
nand U16096 (N_16096,N_15912,N_15963);
or U16097 (N_16097,N_15826,N_15917);
nand U16098 (N_16098,N_15873,N_15996);
nand U16099 (N_16099,N_15833,N_15958);
xnor U16100 (N_16100,N_15881,N_15941);
or U16101 (N_16101,N_15922,N_15998);
or U16102 (N_16102,N_15942,N_15868);
xor U16103 (N_16103,N_15869,N_15854);
or U16104 (N_16104,N_15949,N_15989);
or U16105 (N_16105,N_15985,N_15818);
or U16106 (N_16106,N_15906,N_15862);
nor U16107 (N_16107,N_15909,N_15880);
and U16108 (N_16108,N_15922,N_15906);
nand U16109 (N_16109,N_15868,N_15940);
nand U16110 (N_16110,N_15907,N_15985);
nand U16111 (N_16111,N_15836,N_15865);
or U16112 (N_16112,N_15931,N_15884);
xnor U16113 (N_16113,N_15964,N_15954);
or U16114 (N_16114,N_15839,N_15988);
xnor U16115 (N_16115,N_15835,N_15984);
nor U16116 (N_16116,N_15916,N_15890);
nand U16117 (N_16117,N_15937,N_15975);
nor U16118 (N_16118,N_15954,N_15881);
xor U16119 (N_16119,N_15800,N_15812);
xor U16120 (N_16120,N_15933,N_15996);
and U16121 (N_16121,N_15879,N_15918);
nand U16122 (N_16122,N_15880,N_15856);
xnor U16123 (N_16123,N_15928,N_15913);
xor U16124 (N_16124,N_15802,N_15828);
nand U16125 (N_16125,N_15950,N_15890);
or U16126 (N_16126,N_15959,N_15861);
nor U16127 (N_16127,N_15859,N_15892);
nand U16128 (N_16128,N_15891,N_15937);
and U16129 (N_16129,N_15948,N_15958);
or U16130 (N_16130,N_15845,N_15835);
and U16131 (N_16131,N_15957,N_15903);
nand U16132 (N_16132,N_15904,N_15956);
xor U16133 (N_16133,N_15957,N_15964);
or U16134 (N_16134,N_15868,N_15902);
nor U16135 (N_16135,N_15819,N_15996);
or U16136 (N_16136,N_15946,N_15830);
or U16137 (N_16137,N_15847,N_15801);
nor U16138 (N_16138,N_15909,N_15925);
and U16139 (N_16139,N_15945,N_15894);
nor U16140 (N_16140,N_15801,N_15834);
nand U16141 (N_16141,N_15919,N_15867);
xor U16142 (N_16142,N_15898,N_15970);
nor U16143 (N_16143,N_15832,N_15967);
nor U16144 (N_16144,N_15892,N_15918);
nor U16145 (N_16145,N_15869,N_15815);
or U16146 (N_16146,N_15927,N_15801);
nand U16147 (N_16147,N_15836,N_15914);
nand U16148 (N_16148,N_15945,N_15803);
and U16149 (N_16149,N_15820,N_15910);
or U16150 (N_16150,N_15952,N_15922);
nor U16151 (N_16151,N_15883,N_15998);
nor U16152 (N_16152,N_15928,N_15880);
xnor U16153 (N_16153,N_15980,N_15900);
xor U16154 (N_16154,N_15893,N_15865);
xnor U16155 (N_16155,N_15889,N_15803);
and U16156 (N_16156,N_15887,N_15892);
or U16157 (N_16157,N_15830,N_15884);
and U16158 (N_16158,N_15896,N_15811);
or U16159 (N_16159,N_15948,N_15975);
or U16160 (N_16160,N_15810,N_15985);
nand U16161 (N_16161,N_15800,N_15862);
and U16162 (N_16162,N_15864,N_15947);
or U16163 (N_16163,N_15872,N_15932);
nor U16164 (N_16164,N_15821,N_15923);
nand U16165 (N_16165,N_15933,N_15961);
xor U16166 (N_16166,N_15875,N_15989);
nand U16167 (N_16167,N_15952,N_15948);
or U16168 (N_16168,N_15990,N_15814);
or U16169 (N_16169,N_15835,N_15954);
nand U16170 (N_16170,N_15928,N_15883);
nand U16171 (N_16171,N_15962,N_15941);
xor U16172 (N_16172,N_15939,N_15873);
nand U16173 (N_16173,N_15839,N_15834);
nor U16174 (N_16174,N_15859,N_15918);
or U16175 (N_16175,N_15920,N_15993);
and U16176 (N_16176,N_15908,N_15984);
or U16177 (N_16177,N_15884,N_15992);
nand U16178 (N_16178,N_15869,N_15856);
xnor U16179 (N_16179,N_15910,N_15915);
xor U16180 (N_16180,N_15949,N_15951);
or U16181 (N_16181,N_15908,N_15981);
xor U16182 (N_16182,N_15928,N_15985);
nor U16183 (N_16183,N_15917,N_15976);
or U16184 (N_16184,N_15891,N_15927);
nor U16185 (N_16185,N_15993,N_15984);
nor U16186 (N_16186,N_15800,N_15838);
and U16187 (N_16187,N_15950,N_15838);
and U16188 (N_16188,N_15939,N_15806);
and U16189 (N_16189,N_15831,N_15932);
nand U16190 (N_16190,N_15853,N_15987);
nand U16191 (N_16191,N_15816,N_15929);
nor U16192 (N_16192,N_15953,N_15869);
or U16193 (N_16193,N_15994,N_15976);
xnor U16194 (N_16194,N_15828,N_15994);
nand U16195 (N_16195,N_15929,N_15878);
nand U16196 (N_16196,N_15955,N_15863);
and U16197 (N_16197,N_15922,N_15831);
nand U16198 (N_16198,N_15825,N_15822);
and U16199 (N_16199,N_15876,N_15834);
xnor U16200 (N_16200,N_16031,N_16192);
or U16201 (N_16201,N_16067,N_16033);
nor U16202 (N_16202,N_16105,N_16030);
nor U16203 (N_16203,N_16189,N_16004);
nand U16204 (N_16204,N_16008,N_16195);
and U16205 (N_16205,N_16072,N_16056);
nand U16206 (N_16206,N_16048,N_16146);
or U16207 (N_16207,N_16168,N_16111);
nor U16208 (N_16208,N_16161,N_16139);
or U16209 (N_16209,N_16035,N_16135);
xor U16210 (N_16210,N_16171,N_16132);
nor U16211 (N_16211,N_16042,N_16175);
xnor U16212 (N_16212,N_16194,N_16186);
xor U16213 (N_16213,N_16063,N_16040);
nand U16214 (N_16214,N_16047,N_16143);
and U16215 (N_16215,N_16115,N_16037);
nand U16216 (N_16216,N_16122,N_16112);
or U16217 (N_16217,N_16180,N_16177);
or U16218 (N_16218,N_16019,N_16165);
nor U16219 (N_16219,N_16087,N_16016);
nand U16220 (N_16220,N_16098,N_16155);
nand U16221 (N_16221,N_16092,N_16134);
nand U16222 (N_16222,N_16064,N_16170);
nand U16223 (N_16223,N_16094,N_16066);
nor U16224 (N_16224,N_16058,N_16153);
and U16225 (N_16225,N_16156,N_16107);
xor U16226 (N_16226,N_16051,N_16078);
nand U16227 (N_16227,N_16068,N_16181);
xor U16228 (N_16228,N_16129,N_16158);
or U16229 (N_16229,N_16059,N_16147);
nor U16230 (N_16230,N_16150,N_16187);
and U16231 (N_16231,N_16009,N_16079);
nand U16232 (N_16232,N_16084,N_16069);
nor U16233 (N_16233,N_16091,N_16032);
nand U16234 (N_16234,N_16025,N_16045);
and U16235 (N_16235,N_16123,N_16061);
or U16236 (N_16236,N_16073,N_16082);
xor U16237 (N_16237,N_16071,N_16006);
and U16238 (N_16238,N_16014,N_16010);
and U16239 (N_16239,N_16164,N_16011);
xor U16240 (N_16240,N_16027,N_16160);
or U16241 (N_16241,N_16121,N_16081);
nor U16242 (N_16242,N_16172,N_16038);
nand U16243 (N_16243,N_16012,N_16050);
or U16244 (N_16244,N_16023,N_16039);
xor U16245 (N_16245,N_16093,N_16149);
nand U16246 (N_16246,N_16106,N_16000);
or U16247 (N_16247,N_16136,N_16103);
or U16248 (N_16248,N_16113,N_16024);
nor U16249 (N_16249,N_16085,N_16097);
xnor U16250 (N_16250,N_16088,N_16017);
nor U16251 (N_16251,N_16052,N_16159);
and U16252 (N_16252,N_16182,N_16196);
and U16253 (N_16253,N_16128,N_16070);
xnor U16254 (N_16254,N_16086,N_16057);
nor U16255 (N_16255,N_16183,N_16133);
or U16256 (N_16256,N_16166,N_16074);
nand U16257 (N_16257,N_16169,N_16154);
or U16258 (N_16258,N_16176,N_16167);
and U16259 (N_16259,N_16055,N_16044);
nand U16260 (N_16260,N_16108,N_16101);
and U16261 (N_16261,N_16100,N_16138);
xnor U16262 (N_16262,N_16117,N_16173);
nor U16263 (N_16263,N_16102,N_16185);
and U16264 (N_16264,N_16190,N_16157);
nor U16265 (N_16265,N_16007,N_16140);
xor U16266 (N_16266,N_16184,N_16003);
or U16267 (N_16267,N_16095,N_16026);
xor U16268 (N_16268,N_16077,N_16178);
or U16269 (N_16269,N_16193,N_16174);
or U16270 (N_16270,N_16163,N_16145);
xnor U16271 (N_16271,N_16130,N_16199);
and U16272 (N_16272,N_16198,N_16076);
nand U16273 (N_16273,N_16080,N_16148);
or U16274 (N_16274,N_16036,N_16197);
nand U16275 (N_16275,N_16131,N_16162);
nand U16276 (N_16276,N_16152,N_16075);
nand U16277 (N_16277,N_16002,N_16142);
and U16278 (N_16278,N_16043,N_16125);
and U16279 (N_16279,N_16151,N_16049);
xor U16280 (N_16280,N_16114,N_16041);
nor U16281 (N_16281,N_16096,N_16022);
nor U16282 (N_16282,N_16021,N_16099);
or U16283 (N_16283,N_16116,N_16034);
and U16284 (N_16284,N_16046,N_16065);
nor U16285 (N_16285,N_16144,N_16083);
or U16286 (N_16286,N_16028,N_16060);
nand U16287 (N_16287,N_16124,N_16179);
xor U16288 (N_16288,N_16029,N_16089);
xnor U16289 (N_16289,N_16054,N_16001);
xor U16290 (N_16290,N_16188,N_16110);
nand U16291 (N_16291,N_16018,N_16015);
or U16292 (N_16292,N_16126,N_16062);
nand U16293 (N_16293,N_16005,N_16013);
or U16294 (N_16294,N_16119,N_16118);
and U16295 (N_16295,N_16137,N_16104);
and U16296 (N_16296,N_16090,N_16053);
and U16297 (N_16297,N_16109,N_16141);
or U16298 (N_16298,N_16127,N_16020);
and U16299 (N_16299,N_16120,N_16191);
nand U16300 (N_16300,N_16016,N_16120);
nor U16301 (N_16301,N_16090,N_16138);
and U16302 (N_16302,N_16175,N_16170);
nor U16303 (N_16303,N_16149,N_16011);
xor U16304 (N_16304,N_16179,N_16090);
nand U16305 (N_16305,N_16197,N_16002);
xnor U16306 (N_16306,N_16041,N_16095);
nand U16307 (N_16307,N_16197,N_16143);
nand U16308 (N_16308,N_16102,N_16073);
or U16309 (N_16309,N_16186,N_16063);
nand U16310 (N_16310,N_16066,N_16124);
or U16311 (N_16311,N_16039,N_16110);
xor U16312 (N_16312,N_16020,N_16004);
and U16313 (N_16313,N_16075,N_16092);
nand U16314 (N_16314,N_16081,N_16190);
and U16315 (N_16315,N_16099,N_16061);
and U16316 (N_16316,N_16171,N_16147);
and U16317 (N_16317,N_16113,N_16158);
nand U16318 (N_16318,N_16030,N_16181);
or U16319 (N_16319,N_16188,N_16163);
or U16320 (N_16320,N_16110,N_16040);
xnor U16321 (N_16321,N_16083,N_16152);
xor U16322 (N_16322,N_16112,N_16116);
nor U16323 (N_16323,N_16122,N_16019);
nand U16324 (N_16324,N_16012,N_16125);
nand U16325 (N_16325,N_16072,N_16043);
or U16326 (N_16326,N_16120,N_16093);
and U16327 (N_16327,N_16190,N_16093);
nand U16328 (N_16328,N_16059,N_16005);
xnor U16329 (N_16329,N_16145,N_16054);
and U16330 (N_16330,N_16073,N_16172);
xnor U16331 (N_16331,N_16139,N_16085);
and U16332 (N_16332,N_16141,N_16180);
nand U16333 (N_16333,N_16020,N_16133);
nand U16334 (N_16334,N_16046,N_16099);
xor U16335 (N_16335,N_16090,N_16165);
and U16336 (N_16336,N_16177,N_16057);
and U16337 (N_16337,N_16056,N_16184);
and U16338 (N_16338,N_16065,N_16000);
nor U16339 (N_16339,N_16160,N_16060);
xnor U16340 (N_16340,N_16075,N_16124);
xnor U16341 (N_16341,N_16187,N_16064);
xor U16342 (N_16342,N_16181,N_16069);
nor U16343 (N_16343,N_16021,N_16127);
nor U16344 (N_16344,N_16018,N_16050);
nor U16345 (N_16345,N_16114,N_16191);
nand U16346 (N_16346,N_16081,N_16067);
and U16347 (N_16347,N_16141,N_16011);
xnor U16348 (N_16348,N_16009,N_16091);
and U16349 (N_16349,N_16060,N_16183);
and U16350 (N_16350,N_16028,N_16182);
xnor U16351 (N_16351,N_16086,N_16101);
or U16352 (N_16352,N_16129,N_16008);
nor U16353 (N_16353,N_16069,N_16037);
nand U16354 (N_16354,N_16034,N_16101);
nand U16355 (N_16355,N_16004,N_16050);
nand U16356 (N_16356,N_16048,N_16191);
nand U16357 (N_16357,N_16007,N_16019);
nand U16358 (N_16358,N_16112,N_16015);
or U16359 (N_16359,N_16038,N_16103);
and U16360 (N_16360,N_16124,N_16029);
nand U16361 (N_16361,N_16048,N_16174);
nand U16362 (N_16362,N_16116,N_16123);
nand U16363 (N_16363,N_16044,N_16106);
or U16364 (N_16364,N_16078,N_16103);
nor U16365 (N_16365,N_16050,N_16009);
and U16366 (N_16366,N_16166,N_16085);
nor U16367 (N_16367,N_16045,N_16143);
and U16368 (N_16368,N_16067,N_16095);
nand U16369 (N_16369,N_16000,N_16066);
nand U16370 (N_16370,N_16169,N_16122);
or U16371 (N_16371,N_16195,N_16194);
nand U16372 (N_16372,N_16173,N_16067);
nor U16373 (N_16373,N_16013,N_16043);
and U16374 (N_16374,N_16192,N_16179);
or U16375 (N_16375,N_16058,N_16020);
nand U16376 (N_16376,N_16117,N_16110);
and U16377 (N_16377,N_16079,N_16054);
xnor U16378 (N_16378,N_16145,N_16005);
and U16379 (N_16379,N_16154,N_16173);
xor U16380 (N_16380,N_16056,N_16179);
or U16381 (N_16381,N_16035,N_16115);
nand U16382 (N_16382,N_16061,N_16046);
nand U16383 (N_16383,N_16073,N_16020);
nor U16384 (N_16384,N_16161,N_16154);
and U16385 (N_16385,N_16196,N_16125);
and U16386 (N_16386,N_16122,N_16067);
or U16387 (N_16387,N_16054,N_16126);
nand U16388 (N_16388,N_16138,N_16035);
nor U16389 (N_16389,N_16078,N_16188);
nand U16390 (N_16390,N_16155,N_16084);
and U16391 (N_16391,N_16062,N_16049);
nand U16392 (N_16392,N_16140,N_16012);
nor U16393 (N_16393,N_16024,N_16051);
nor U16394 (N_16394,N_16043,N_16114);
nand U16395 (N_16395,N_16116,N_16188);
and U16396 (N_16396,N_16094,N_16161);
nand U16397 (N_16397,N_16007,N_16086);
and U16398 (N_16398,N_16055,N_16030);
nand U16399 (N_16399,N_16044,N_16107);
nor U16400 (N_16400,N_16272,N_16365);
xnor U16401 (N_16401,N_16275,N_16261);
xor U16402 (N_16402,N_16246,N_16293);
nand U16403 (N_16403,N_16311,N_16255);
or U16404 (N_16404,N_16273,N_16395);
nor U16405 (N_16405,N_16238,N_16288);
xnor U16406 (N_16406,N_16374,N_16203);
and U16407 (N_16407,N_16339,N_16333);
and U16408 (N_16408,N_16377,N_16223);
xnor U16409 (N_16409,N_16356,N_16259);
and U16410 (N_16410,N_16282,N_16392);
nand U16411 (N_16411,N_16300,N_16207);
nor U16412 (N_16412,N_16280,N_16228);
nor U16413 (N_16413,N_16310,N_16361);
nand U16414 (N_16414,N_16347,N_16294);
or U16415 (N_16415,N_16299,N_16321);
xnor U16416 (N_16416,N_16370,N_16235);
nor U16417 (N_16417,N_16380,N_16285);
nor U16418 (N_16418,N_16357,N_16268);
or U16419 (N_16419,N_16390,N_16263);
or U16420 (N_16420,N_16305,N_16260);
nor U16421 (N_16421,N_16215,N_16249);
nor U16422 (N_16422,N_16327,N_16338);
nor U16423 (N_16423,N_16329,N_16369);
xor U16424 (N_16424,N_16386,N_16232);
and U16425 (N_16425,N_16334,N_16391);
nand U16426 (N_16426,N_16258,N_16319);
or U16427 (N_16427,N_16332,N_16382);
nand U16428 (N_16428,N_16242,N_16267);
xnor U16429 (N_16429,N_16396,N_16230);
nand U16430 (N_16430,N_16211,N_16381);
nand U16431 (N_16431,N_16291,N_16297);
nand U16432 (N_16432,N_16353,N_16237);
nor U16433 (N_16433,N_16359,N_16313);
or U16434 (N_16434,N_16385,N_16284);
nand U16435 (N_16435,N_16204,N_16248);
xor U16436 (N_16436,N_16229,N_16378);
nor U16437 (N_16437,N_16373,N_16308);
and U16438 (N_16438,N_16241,N_16205);
or U16439 (N_16439,N_16227,N_16325);
nor U16440 (N_16440,N_16399,N_16234);
or U16441 (N_16441,N_16328,N_16340);
nor U16442 (N_16442,N_16362,N_16271);
nand U16443 (N_16443,N_16336,N_16335);
or U16444 (N_16444,N_16345,N_16371);
nand U16445 (N_16445,N_16262,N_16375);
nand U16446 (N_16446,N_16312,N_16276);
or U16447 (N_16447,N_16298,N_16253);
and U16448 (N_16448,N_16344,N_16279);
and U16449 (N_16449,N_16358,N_16309);
and U16450 (N_16450,N_16323,N_16202);
or U16451 (N_16451,N_16292,N_16214);
xor U16452 (N_16452,N_16383,N_16351);
nand U16453 (N_16453,N_16303,N_16316);
and U16454 (N_16454,N_16247,N_16252);
nand U16455 (N_16455,N_16257,N_16337);
and U16456 (N_16456,N_16317,N_16213);
nand U16457 (N_16457,N_16278,N_16239);
and U16458 (N_16458,N_16240,N_16265);
xnor U16459 (N_16459,N_16219,N_16314);
or U16460 (N_16460,N_16283,N_16307);
and U16461 (N_16461,N_16368,N_16286);
nor U16462 (N_16462,N_16210,N_16243);
or U16463 (N_16463,N_16302,N_16388);
nand U16464 (N_16464,N_16320,N_16331);
nand U16465 (N_16465,N_16231,N_16245);
xor U16466 (N_16466,N_16226,N_16206);
xor U16467 (N_16467,N_16296,N_16366);
nand U16468 (N_16468,N_16360,N_16364);
xor U16469 (N_16469,N_16346,N_16270);
nor U16470 (N_16470,N_16304,N_16269);
or U16471 (N_16471,N_16287,N_16301);
and U16472 (N_16472,N_16251,N_16306);
nor U16473 (N_16473,N_16341,N_16394);
nor U16474 (N_16474,N_16281,N_16224);
nor U16475 (N_16475,N_16256,N_16221);
nand U16476 (N_16476,N_16355,N_16350);
or U16477 (N_16477,N_16289,N_16326);
or U16478 (N_16478,N_16212,N_16384);
and U16479 (N_16479,N_16254,N_16372);
nor U16480 (N_16480,N_16387,N_16200);
xor U16481 (N_16481,N_16244,N_16222);
or U16482 (N_16482,N_16277,N_16322);
xnor U16483 (N_16483,N_16352,N_16363);
xor U16484 (N_16484,N_16290,N_16349);
nand U16485 (N_16485,N_16354,N_16330);
xor U16486 (N_16486,N_16266,N_16201);
or U16487 (N_16487,N_16318,N_16376);
nor U16488 (N_16488,N_16367,N_16393);
xor U16489 (N_16489,N_16216,N_16389);
and U16490 (N_16490,N_16225,N_16295);
or U16491 (N_16491,N_16324,N_16379);
and U16492 (N_16492,N_16233,N_16220);
or U16493 (N_16493,N_16217,N_16236);
nor U16494 (N_16494,N_16274,N_16398);
xnor U16495 (N_16495,N_16218,N_16342);
or U16496 (N_16496,N_16315,N_16264);
nand U16497 (N_16497,N_16397,N_16348);
nand U16498 (N_16498,N_16209,N_16208);
and U16499 (N_16499,N_16343,N_16250);
nand U16500 (N_16500,N_16212,N_16309);
nand U16501 (N_16501,N_16219,N_16201);
nor U16502 (N_16502,N_16354,N_16316);
and U16503 (N_16503,N_16388,N_16363);
xor U16504 (N_16504,N_16348,N_16328);
or U16505 (N_16505,N_16233,N_16367);
and U16506 (N_16506,N_16309,N_16249);
or U16507 (N_16507,N_16319,N_16266);
xor U16508 (N_16508,N_16230,N_16276);
xnor U16509 (N_16509,N_16356,N_16343);
nor U16510 (N_16510,N_16386,N_16365);
nand U16511 (N_16511,N_16210,N_16230);
xnor U16512 (N_16512,N_16310,N_16351);
and U16513 (N_16513,N_16293,N_16316);
nor U16514 (N_16514,N_16246,N_16272);
nand U16515 (N_16515,N_16224,N_16325);
nor U16516 (N_16516,N_16390,N_16386);
nor U16517 (N_16517,N_16267,N_16286);
xor U16518 (N_16518,N_16250,N_16202);
xor U16519 (N_16519,N_16356,N_16394);
and U16520 (N_16520,N_16367,N_16293);
nor U16521 (N_16521,N_16375,N_16254);
or U16522 (N_16522,N_16259,N_16217);
or U16523 (N_16523,N_16223,N_16269);
xor U16524 (N_16524,N_16300,N_16376);
xor U16525 (N_16525,N_16358,N_16245);
nor U16526 (N_16526,N_16278,N_16375);
nor U16527 (N_16527,N_16274,N_16285);
and U16528 (N_16528,N_16351,N_16278);
nand U16529 (N_16529,N_16236,N_16289);
nand U16530 (N_16530,N_16233,N_16361);
xor U16531 (N_16531,N_16222,N_16371);
and U16532 (N_16532,N_16306,N_16356);
nand U16533 (N_16533,N_16356,N_16230);
nor U16534 (N_16534,N_16378,N_16247);
and U16535 (N_16535,N_16213,N_16217);
xor U16536 (N_16536,N_16252,N_16325);
and U16537 (N_16537,N_16337,N_16393);
nand U16538 (N_16538,N_16203,N_16258);
xor U16539 (N_16539,N_16322,N_16319);
and U16540 (N_16540,N_16263,N_16331);
xor U16541 (N_16541,N_16376,N_16367);
nor U16542 (N_16542,N_16335,N_16384);
and U16543 (N_16543,N_16235,N_16277);
nor U16544 (N_16544,N_16238,N_16223);
nand U16545 (N_16545,N_16278,N_16299);
nor U16546 (N_16546,N_16322,N_16269);
and U16547 (N_16547,N_16369,N_16343);
or U16548 (N_16548,N_16314,N_16316);
xor U16549 (N_16549,N_16366,N_16343);
nand U16550 (N_16550,N_16384,N_16224);
or U16551 (N_16551,N_16200,N_16219);
and U16552 (N_16552,N_16262,N_16208);
and U16553 (N_16553,N_16264,N_16287);
or U16554 (N_16554,N_16395,N_16308);
and U16555 (N_16555,N_16274,N_16204);
nand U16556 (N_16556,N_16254,N_16227);
nand U16557 (N_16557,N_16383,N_16387);
or U16558 (N_16558,N_16358,N_16272);
xnor U16559 (N_16559,N_16378,N_16360);
or U16560 (N_16560,N_16253,N_16373);
and U16561 (N_16561,N_16357,N_16254);
nand U16562 (N_16562,N_16238,N_16259);
or U16563 (N_16563,N_16371,N_16293);
or U16564 (N_16564,N_16229,N_16283);
xnor U16565 (N_16565,N_16368,N_16390);
nor U16566 (N_16566,N_16224,N_16338);
xnor U16567 (N_16567,N_16236,N_16220);
or U16568 (N_16568,N_16248,N_16365);
nor U16569 (N_16569,N_16338,N_16331);
xnor U16570 (N_16570,N_16209,N_16379);
xnor U16571 (N_16571,N_16286,N_16273);
and U16572 (N_16572,N_16374,N_16397);
and U16573 (N_16573,N_16238,N_16284);
nand U16574 (N_16574,N_16309,N_16205);
nor U16575 (N_16575,N_16239,N_16312);
or U16576 (N_16576,N_16208,N_16244);
or U16577 (N_16577,N_16329,N_16392);
or U16578 (N_16578,N_16259,N_16351);
nor U16579 (N_16579,N_16373,N_16372);
nand U16580 (N_16580,N_16274,N_16216);
nand U16581 (N_16581,N_16357,N_16384);
and U16582 (N_16582,N_16278,N_16358);
nor U16583 (N_16583,N_16389,N_16378);
nand U16584 (N_16584,N_16356,N_16353);
nor U16585 (N_16585,N_16345,N_16361);
and U16586 (N_16586,N_16397,N_16260);
nand U16587 (N_16587,N_16385,N_16225);
nor U16588 (N_16588,N_16322,N_16214);
or U16589 (N_16589,N_16241,N_16217);
xnor U16590 (N_16590,N_16248,N_16371);
and U16591 (N_16591,N_16252,N_16306);
xor U16592 (N_16592,N_16396,N_16326);
nand U16593 (N_16593,N_16201,N_16286);
and U16594 (N_16594,N_16308,N_16362);
xnor U16595 (N_16595,N_16368,N_16277);
nand U16596 (N_16596,N_16371,N_16389);
or U16597 (N_16597,N_16358,N_16286);
xor U16598 (N_16598,N_16214,N_16371);
xor U16599 (N_16599,N_16313,N_16293);
and U16600 (N_16600,N_16591,N_16561);
and U16601 (N_16601,N_16531,N_16406);
and U16602 (N_16602,N_16400,N_16490);
nand U16603 (N_16603,N_16555,N_16527);
and U16604 (N_16604,N_16467,N_16488);
and U16605 (N_16605,N_16435,N_16510);
and U16606 (N_16606,N_16525,N_16568);
nand U16607 (N_16607,N_16486,N_16564);
and U16608 (N_16608,N_16562,N_16468);
nor U16609 (N_16609,N_16418,N_16457);
nor U16610 (N_16610,N_16407,N_16502);
or U16611 (N_16611,N_16405,N_16432);
nand U16612 (N_16612,N_16491,N_16416);
and U16613 (N_16613,N_16574,N_16483);
and U16614 (N_16614,N_16499,N_16542);
nand U16615 (N_16615,N_16466,N_16414);
nor U16616 (N_16616,N_16547,N_16598);
xnor U16617 (N_16617,N_16514,N_16540);
or U16618 (N_16618,N_16410,N_16520);
and U16619 (N_16619,N_16589,N_16427);
and U16620 (N_16620,N_16492,N_16539);
or U16621 (N_16621,N_16523,N_16597);
or U16622 (N_16622,N_16595,N_16469);
nor U16623 (N_16623,N_16573,N_16579);
nand U16624 (N_16624,N_16541,N_16534);
nor U16625 (N_16625,N_16478,N_16455);
xor U16626 (N_16626,N_16423,N_16585);
xor U16627 (N_16627,N_16484,N_16563);
and U16628 (N_16628,N_16460,N_16402);
xnor U16629 (N_16629,N_16553,N_16463);
or U16630 (N_16630,N_16425,N_16507);
and U16631 (N_16631,N_16503,N_16551);
or U16632 (N_16632,N_16528,N_16538);
or U16633 (N_16633,N_16442,N_16493);
or U16634 (N_16634,N_16560,N_16586);
and U16635 (N_16635,N_16565,N_16494);
nor U16636 (N_16636,N_16530,N_16496);
xnor U16637 (N_16637,N_16417,N_16409);
and U16638 (N_16638,N_16446,N_16479);
and U16639 (N_16639,N_16545,N_16511);
nand U16640 (N_16640,N_16576,N_16566);
xnor U16641 (N_16641,N_16512,N_16537);
nor U16642 (N_16642,N_16515,N_16567);
nor U16643 (N_16643,N_16558,N_16428);
or U16644 (N_16644,N_16495,N_16554);
and U16645 (N_16645,N_16453,N_16521);
nand U16646 (N_16646,N_16408,N_16403);
or U16647 (N_16647,N_16588,N_16487);
or U16648 (N_16648,N_16412,N_16451);
nand U16649 (N_16649,N_16519,N_16533);
nor U16650 (N_16650,N_16454,N_16536);
xor U16651 (N_16651,N_16508,N_16522);
nor U16652 (N_16652,N_16549,N_16433);
or U16653 (N_16653,N_16584,N_16535);
and U16654 (N_16654,N_16594,N_16476);
nor U16655 (N_16655,N_16420,N_16570);
and U16656 (N_16656,N_16459,N_16571);
nor U16657 (N_16657,N_16404,N_16413);
nand U16658 (N_16658,N_16415,N_16444);
xor U16659 (N_16659,N_16472,N_16548);
xnor U16660 (N_16660,N_16504,N_16532);
nor U16661 (N_16661,N_16434,N_16458);
xnor U16662 (N_16662,N_16481,N_16431);
nand U16663 (N_16663,N_16578,N_16518);
or U16664 (N_16664,N_16580,N_16572);
nand U16665 (N_16665,N_16498,N_16430);
and U16666 (N_16666,N_16582,N_16445);
nand U16667 (N_16667,N_16526,N_16475);
or U16668 (N_16668,N_16443,N_16439);
nand U16669 (N_16669,N_16456,N_16470);
or U16670 (N_16670,N_16422,N_16421);
and U16671 (N_16671,N_16517,N_16452);
nand U16672 (N_16672,N_16473,N_16401);
nand U16673 (N_16673,N_16524,N_16429);
xnor U16674 (N_16674,N_16447,N_16592);
or U16675 (N_16675,N_16449,N_16419);
or U16676 (N_16676,N_16424,N_16596);
xor U16677 (N_16677,N_16544,N_16552);
xnor U16678 (N_16678,N_16529,N_16497);
nor U16679 (N_16679,N_16437,N_16461);
nand U16680 (N_16680,N_16465,N_16546);
nand U16681 (N_16681,N_16581,N_16575);
nor U16682 (N_16682,N_16448,N_16569);
and U16683 (N_16683,N_16509,N_16505);
xor U16684 (N_16684,N_16559,N_16516);
xnor U16685 (N_16685,N_16506,N_16450);
nor U16686 (N_16686,N_16599,N_16556);
xor U16687 (N_16687,N_16590,N_16587);
xor U16688 (N_16688,N_16500,N_16550);
xor U16689 (N_16689,N_16464,N_16426);
or U16690 (N_16690,N_16482,N_16543);
nand U16691 (N_16691,N_16462,N_16577);
and U16692 (N_16692,N_16501,N_16480);
xor U16693 (N_16693,N_16440,N_16489);
xnor U16694 (N_16694,N_16485,N_16474);
and U16695 (N_16695,N_16513,N_16471);
nand U16696 (N_16696,N_16436,N_16583);
nor U16697 (N_16697,N_16557,N_16593);
xnor U16698 (N_16698,N_16441,N_16438);
xnor U16699 (N_16699,N_16411,N_16477);
nand U16700 (N_16700,N_16450,N_16548);
nand U16701 (N_16701,N_16424,N_16415);
xnor U16702 (N_16702,N_16482,N_16549);
xor U16703 (N_16703,N_16471,N_16494);
nor U16704 (N_16704,N_16509,N_16433);
nand U16705 (N_16705,N_16537,N_16477);
xor U16706 (N_16706,N_16401,N_16429);
nor U16707 (N_16707,N_16505,N_16494);
and U16708 (N_16708,N_16458,N_16550);
xnor U16709 (N_16709,N_16557,N_16439);
xnor U16710 (N_16710,N_16585,N_16402);
nand U16711 (N_16711,N_16429,N_16554);
nand U16712 (N_16712,N_16480,N_16510);
or U16713 (N_16713,N_16583,N_16509);
or U16714 (N_16714,N_16414,N_16577);
nand U16715 (N_16715,N_16468,N_16460);
or U16716 (N_16716,N_16588,N_16499);
or U16717 (N_16717,N_16486,N_16424);
or U16718 (N_16718,N_16428,N_16520);
and U16719 (N_16719,N_16458,N_16438);
or U16720 (N_16720,N_16528,N_16506);
nand U16721 (N_16721,N_16511,N_16453);
xnor U16722 (N_16722,N_16584,N_16475);
or U16723 (N_16723,N_16578,N_16415);
xnor U16724 (N_16724,N_16564,N_16547);
nor U16725 (N_16725,N_16499,N_16553);
or U16726 (N_16726,N_16439,N_16462);
or U16727 (N_16727,N_16430,N_16580);
xor U16728 (N_16728,N_16445,N_16493);
nand U16729 (N_16729,N_16590,N_16419);
nand U16730 (N_16730,N_16481,N_16434);
or U16731 (N_16731,N_16402,N_16532);
nor U16732 (N_16732,N_16511,N_16480);
and U16733 (N_16733,N_16516,N_16476);
nand U16734 (N_16734,N_16556,N_16447);
nor U16735 (N_16735,N_16493,N_16403);
nor U16736 (N_16736,N_16579,N_16591);
or U16737 (N_16737,N_16400,N_16420);
xnor U16738 (N_16738,N_16570,N_16455);
or U16739 (N_16739,N_16476,N_16437);
xnor U16740 (N_16740,N_16444,N_16486);
nand U16741 (N_16741,N_16524,N_16476);
nand U16742 (N_16742,N_16457,N_16505);
nand U16743 (N_16743,N_16504,N_16456);
xor U16744 (N_16744,N_16462,N_16551);
nor U16745 (N_16745,N_16532,N_16468);
or U16746 (N_16746,N_16586,N_16487);
or U16747 (N_16747,N_16576,N_16597);
nand U16748 (N_16748,N_16455,N_16479);
and U16749 (N_16749,N_16468,N_16432);
and U16750 (N_16750,N_16495,N_16555);
nand U16751 (N_16751,N_16454,N_16554);
nand U16752 (N_16752,N_16473,N_16443);
and U16753 (N_16753,N_16540,N_16479);
nor U16754 (N_16754,N_16585,N_16455);
and U16755 (N_16755,N_16470,N_16400);
nor U16756 (N_16756,N_16488,N_16431);
and U16757 (N_16757,N_16545,N_16401);
or U16758 (N_16758,N_16407,N_16487);
or U16759 (N_16759,N_16423,N_16411);
nor U16760 (N_16760,N_16589,N_16494);
xor U16761 (N_16761,N_16594,N_16565);
xnor U16762 (N_16762,N_16540,N_16557);
xor U16763 (N_16763,N_16468,N_16583);
or U16764 (N_16764,N_16482,N_16535);
xor U16765 (N_16765,N_16420,N_16481);
xnor U16766 (N_16766,N_16427,N_16478);
xnor U16767 (N_16767,N_16449,N_16536);
xor U16768 (N_16768,N_16504,N_16403);
xnor U16769 (N_16769,N_16561,N_16510);
nand U16770 (N_16770,N_16561,N_16592);
nor U16771 (N_16771,N_16488,N_16425);
xnor U16772 (N_16772,N_16596,N_16487);
xnor U16773 (N_16773,N_16541,N_16494);
nand U16774 (N_16774,N_16493,N_16499);
or U16775 (N_16775,N_16585,N_16557);
and U16776 (N_16776,N_16439,N_16470);
nand U16777 (N_16777,N_16564,N_16452);
nand U16778 (N_16778,N_16562,N_16436);
nor U16779 (N_16779,N_16547,N_16572);
and U16780 (N_16780,N_16436,N_16428);
and U16781 (N_16781,N_16460,N_16470);
xnor U16782 (N_16782,N_16421,N_16576);
and U16783 (N_16783,N_16519,N_16472);
nor U16784 (N_16784,N_16402,N_16544);
and U16785 (N_16785,N_16540,N_16545);
nor U16786 (N_16786,N_16439,N_16568);
and U16787 (N_16787,N_16539,N_16574);
nor U16788 (N_16788,N_16554,N_16581);
nand U16789 (N_16789,N_16474,N_16520);
nand U16790 (N_16790,N_16514,N_16577);
and U16791 (N_16791,N_16478,N_16460);
xnor U16792 (N_16792,N_16574,N_16564);
xor U16793 (N_16793,N_16404,N_16582);
or U16794 (N_16794,N_16580,N_16565);
nor U16795 (N_16795,N_16547,N_16494);
nand U16796 (N_16796,N_16590,N_16428);
xnor U16797 (N_16797,N_16589,N_16569);
or U16798 (N_16798,N_16548,N_16527);
xnor U16799 (N_16799,N_16444,N_16485);
xnor U16800 (N_16800,N_16741,N_16708);
and U16801 (N_16801,N_16793,N_16619);
or U16802 (N_16802,N_16611,N_16655);
nor U16803 (N_16803,N_16640,N_16624);
xor U16804 (N_16804,N_16766,N_16769);
nand U16805 (N_16805,N_16789,N_16767);
nand U16806 (N_16806,N_16790,N_16719);
nand U16807 (N_16807,N_16696,N_16758);
nor U16808 (N_16808,N_16765,N_16697);
nor U16809 (N_16809,N_16603,N_16623);
nand U16810 (N_16810,N_16717,N_16667);
and U16811 (N_16811,N_16636,N_16706);
and U16812 (N_16812,N_16771,N_16651);
xnor U16813 (N_16813,N_16720,N_16698);
nor U16814 (N_16814,N_16723,N_16763);
or U16815 (N_16815,N_16747,N_16736);
and U16816 (N_16816,N_16710,N_16722);
and U16817 (N_16817,N_16703,N_16709);
xor U16818 (N_16818,N_16671,N_16725);
or U16819 (N_16819,N_16783,N_16733);
xnor U16820 (N_16820,N_16724,N_16660);
or U16821 (N_16821,N_16687,N_16744);
and U16822 (N_16822,N_16694,N_16662);
and U16823 (N_16823,N_16704,N_16738);
xnor U16824 (N_16824,N_16643,N_16677);
xnor U16825 (N_16825,N_16727,N_16641);
xnor U16826 (N_16826,N_16761,N_16752);
nand U16827 (N_16827,N_16701,N_16787);
nand U16828 (N_16828,N_16755,N_16748);
and U16829 (N_16829,N_16777,N_16718);
and U16830 (N_16830,N_16616,N_16735);
nor U16831 (N_16831,N_16740,N_16684);
or U16832 (N_16832,N_16670,N_16776);
or U16833 (N_16833,N_16689,N_16672);
nor U16834 (N_16834,N_16786,N_16605);
or U16835 (N_16835,N_16768,N_16764);
or U16836 (N_16836,N_16679,N_16760);
or U16837 (N_16837,N_16652,N_16642);
nor U16838 (N_16838,N_16699,N_16618);
or U16839 (N_16839,N_16762,N_16692);
or U16840 (N_16840,N_16609,N_16665);
xnor U16841 (N_16841,N_16678,N_16686);
nor U16842 (N_16842,N_16732,N_16756);
and U16843 (N_16843,N_16743,N_16635);
or U16844 (N_16844,N_16674,N_16680);
or U16845 (N_16845,N_16625,N_16796);
or U16846 (N_16846,N_16614,N_16633);
nand U16847 (N_16847,N_16770,N_16647);
nor U16848 (N_16848,N_16649,N_16601);
nand U16849 (N_16849,N_16658,N_16773);
nand U16850 (N_16850,N_16673,N_16745);
xor U16851 (N_16851,N_16757,N_16685);
or U16852 (N_16852,N_16659,N_16690);
nand U16853 (N_16853,N_16664,N_16617);
nor U16854 (N_16854,N_16737,N_16791);
or U16855 (N_16855,N_16713,N_16782);
nand U16856 (N_16856,N_16646,N_16666);
xor U16857 (N_16857,N_16688,N_16648);
nor U16858 (N_16858,N_16612,N_16691);
xnor U16859 (N_16859,N_16602,N_16778);
nand U16860 (N_16860,N_16600,N_16731);
and U16861 (N_16861,N_16775,N_16693);
xnor U16862 (N_16862,N_16661,N_16622);
and U16863 (N_16863,N_16606,N_16610);
or U16864 (N_16864,N_16750,N_16754);
xnor U16865 (N_16865,N_16668,N_16656);
or U16866 (N_16866,N_16607,N_16639);
xor U16867 (N_16867,N_16749,N_16638);
nand U16868 (N_16868,N_16779,N_16608);
or U16869 (N_16869,N_16728,N_16739);
or U16870 (N_16870,N_16729,N_16785);
and U16871 (N_16871,N_16734,N_16798);
or U16872 (N_16872,N_16781,N_16797);
nand U16873 (N_16873,N_16645,N_16628);
or U16874 (N_16874,N_16682,N_16759);
or U16875 (N_16875,N_16746,N_16712);
nor U16876 (N_16876,N_16695,N_16751);
and U16877 (N_16877,N_16784,N_16632);
and U16878 (N_16878,N_16621,N_16615);
nand U16879 (N_16879,N_16650,N_16788);
nor U16880 (N_16880,N_16794,N_16604);
nor U16881 (N_16881,N_16700,N_16795);
xor U16882 (N_16882,N_16711,N_16753);
nand U16883 (N_16883,N_16629,N_16705);
and U16884 (N_16884,N_16730,N_16721);
or U16885 (N_16885,N_16644,N_16627);
nor U16886 (N_16886,N_16669,N_16681);
or U16887 (N_16887,N_16702,N_16707);
nand U16888 (N_16888,N_16613,N_16716);
nor U16889 (N_16889,N_16792,N_16620);
or U16890 (N_16890,N_16714,N_16715);
or U16891 (N_16891,N_16742,N_16676);
nand U16892 (N_16892,N_16675,N_16653);
and U16893 (N_16893,N_16683,N_16634);
or U16894 (N_16894,N_16774,N_16663);
and U16895 (N_16895,N_16657,N_16637);
xor U16896 (N_16896,N_16654,N_16726);
xor U16897 (N_16897,N_16631,N_16626);
nor U16898 (N_16898,N_16799,N_16780);
xor U16899 (N_16899,N_16630,N_16772);
nand U16900 (N_16900,N_16609,N_16796);
or U16901 (N_16901,N_16705,N_16647);
xor U16902 (N_16902,N_16657,N_16603);
and U16903 (N_16903,N_16765,N_16761);
and U16904 (N_16904,N_16679,N_16701);
nand U16905 (N_16905,N_16729,N_16710);
nor U16906 (N_16906,N_16776,N_16647);
or U16907 (N_16907,N_16692,N_16635);
xor U16908 (N_16908,N_16638,N_16702);
nand U16909 (N_16909,N_16749,N_16640);
and U16910 (N_16910,N_16636,N_16612);
nand U16911 (N_16911,N_16696,N_16609);
xor U16912 (N_16912,N_16614,N_16664);
nor U16913 (N_16913,N_16735,N_16729);
nand U16914 (N_16914,N_16732,N_16759);
nand U16915 (N_16915,N_16746,N_16681);
xor U16916 (N_16916,N_16661,N_16680);
xor U16917 (N_16917,N_16717,N_16629);
nand U16918 (N_16918,N_16661,N_16700);
xnor U16919 (N_16919,N_16626,N_16630);
nand U16920 (N_16920,N_16790,N_16672);
and U16921 (N_16921,N_16780,N_16602);
xor U16922 (N_16922,N_16786,N_16612);
and U16923 (N_16923,N_16670,N_16714);
or U16924 (N_16924,N_16601,N_16728);
and U16925 (N_16925,N_16775,N_16711);
and U16926 (N_16926,N_16742,N_16602);
and U16927 (N_16927,N_16677,N_16610);
xor U16928 (N_16928,N_16765,N_16755);
nor U16929 (N_16929,N_16782,N_16626);
nand U16930 (N_16930,N_16791,N_16620);
xnor U16931 (N_16931,N_16767,N_16742);
or U16932 (N_16932,N_16701,N_16691);
or U16933 (N_16933,N_16697,N_16664);
xnor U16934 (N_16934,N_16624,N_16715);
nor U16935 (N_16935,N_16636,N_16758);
nor U16936 (N_16936,N_16712,N_16623);
or U16937 (N_16937,N_16737,N_16771);
nand U16938 (N_16938,N_16683,N_16670);
or U16939 (N_16939,N_16618,N_16660);
and U16940 (N_16940,N_16757,N_16652);
and U16941 (N_16941,N_16640,N_16634);
xor U16942 (N_16942,N_16609,N_16625);
and U16943 (N_16943,N_16787,N_16799);
and U16944 (N_16944,N_16715,N_16600);
and U16945 (N_16945,N_16668,N_16788);
or U16946 (N_16946,N_16748,N_16666);
nor U16947 (N_16947,N_16761,N_16674);
xor U16948 (N_16948,N_16690,N_16650);
nor U16949 (N_16949,N_16604,N_16753);
nor U16950 (N_16950,N_16771,N_16722);
nand U16951 (N_16951,N_16788,N_16696);
and U16952 (N_16952,N_16633,N_16670);
nor U16953 (N_16953,N_16787,N_16792);
xnor U16954 (N_16954,N_16766,N_16785);
and U16955 (N_16955,N_16742,N_16704);
nor U16956 (N_16956,N_16617,N_16686);
nor U16957 (N_16957,N_16660,N_16791);
xor U16958 (N_16958,N_16675,N_16664);
xnor U16959 (N_16959,N_16670,N_16663);
and U16960 (N_16960,N_16762,N_16678);
or U16961 (N_16961,N_16630,N_16790);
or U16962 (N_16962,N_16731,N_16784);
or U16963 (N_16963,N_16645,N_16644);
nand U16964 (N_16964,N_16613,N_16610);
and U16965 (N_16965,N_16767,N_16711);
or U16966 (N_16966,N_16712,N_16702);
nand U16967 (N_16967,N_16793,N_16695);
nor U16968 (N_16968,N_16764,N_16607);
nor U16969 (N_16969,N_16753,N_16747);
and U16970 (N_16970,N_16664,N_16677);
xnor U16971 (N_16971,N_16701,N_16639);
xnor U16972 (N_16972,N_16787,N_16679);
xor U16973 (N_16973,N_16748,N_16627);
or U16974 (N_16974,N_16647,N_16755);
nor U16975 (N_16975,N_16768,N_16644);
and U16976 (N_16976,N_16713,N_16753);
xor U16977 (N_16977,N_16645,N_16685);
or U16978 (N_16978,N_16624,N_16770);
and U16979 (N_16979,N_16663,N_16720);
and U16980 (N_16980,N_16711,N_16714);
nand U16981 (N_16981,N_16631,N_16669);
or U16982 (N_16982,N_16665,N_16653);
xnor U16983 (N_16983,N_16629,N_16700);
nand U16984 (N_16984,N_16794,N_16737);
xnor U16985 (N_16985,N_16791,N_16664);
nor U16986 (N_16986,N_16690,N_16694);
xnor U16987 (N_16987,N_16725,N_16720);
nand U16988 (N_16988,N_16737,N_16690);
nor U16989 (N_16989,N_16712,N_16700);
nand U16990 (N_16990,N_16682,N_16773);
nor U16991 (N_16991,N_16768,N_16657);
xnor U16992 (N_16992,N_16606,N_16739);
nand U16993 (N_16993,N_16767,N_16631);
nor U16994 (N_16994,N_16644,N_16770);
or U16995 (N_16995,N_16682,N_16649);
nor U16996 (N_16996,N_16777,N_16798);
nand U16997 (N_16997,N_16774,N_16743);
nand U16998 (N_16998,N_16618,N_16746);
and U16999 (N_16999,N_16786,N_16607);
nor U17000 (N_17000,N_16801,N_16915);
nor U17001 (N_17001,N_16832,N_16932);
nand U17002 (N_17002,N_16982,N_16959);
and U17003 (N_17003,N_16993,N_16933);
nor U17004 (N_17004,N_16828,N_16950);
and U17005 (N_17005,N_16805,N_16877);
nand U17006 (N_17006,N_16968,N_16897);
nor U17007 (N_17007,N_16906,N_16857);
or U17008 (N_17008,N_16967,N_16984);
xor U17009 (N_17009,N_16973,N_16889);
and U17010 (N_17010,N_16917,N_16859);
and U17011 (N_17011,N_16909,N_16987);
nand U17012 (N_17012,N_16800,N_16818);
nand U17013 (N_17013,N_16895,N_16998);
and U17014 (N_17014,N_16927,N_16823);
xor U17015 (N_17015,N_16937,N_16876);
nor U17016 (N_17016,N_16843,N_16885);
or U17017 (N_17017,N_16899,N_16854);
or U17018 (N_17018,N_16913,N_16955);
nand U17019 (N_17019,N_16958,N_16803);
or U17020 (N_17020,N_16979,N_16995);
and U17021 (N_17021,N_16947,N_16893);
and U17022 (N_17022,N_16983,N_16848);
xnor U17023 (N_17023,N_16837,N_16992);
nand U17024 (N_17024,N_16864,N_16817);
xor U17025 (N_17025,N_16901,N_16902);
nand U17026 (N_17026,N_16989,N_16980);
or U17027 (N_17027,N_16939,N_16841);
nor U17028 (N_17028,N_16840,N_16863);
or U17029 (N_17029,N_16809,N_16961);
xnor U17030 (N_17030,N_16861,N_16886);
and U17031 (N_17031,N_16804,N_16948);
xor U17032 (N_17032,N_16997,N_16810);
xor U17033 (N_17033,N_16911,N_16918);
or U17034 (N_17034,N_16966,N_16925);
and U17035 (N_17035,N_16962,N_16881);
nand U17036 (N_17036,N_16905,N_16985);
nor U17037 (N_17037,N_16926,N_16855);
or U17038 (N_17038,N_16976,N_16875);
nand U17039 (N_17039,N_16922,N_16816);
nand U17040 (N_17040,N_16956,N_16891);
xnor U17041 (N_17041,N_16806,N_16953);
or U17042 (N_17042,N_16991,N_16934);
xor U17043 (N_17043,N_16943,N_16900);
and U17044 (N_17044,N_16825,N_16888);
or U17045 (N_17045,N_16957,N_16868);
or U17046 (N_17046,N_16839,N_16972);
xnor U17047 (N_17047,N_16894,N_16879);
nand U17048 (N_17048,N_16990,N_16834);
nand U17049 (N_17049,N_16963,N_16988);
nor U17050 (N_17050,N_16812,N_16960);
and U17051 (N_17051,N_16846,N_16996);
or U17052 (N_17052,N_16929,N_16849);
or U17053 (N_17053,N_16870,N_16999);
xor U17054 (N_17054,N_16836,N_16852);
nand U17055 (N_17055,N_16814,N_16907);
xor U17056 (N_17056,N_16819,N_16952);
nand U17057 (N_17057,N_16903,N_16887);
nor U17058 (N_17058,N_16942,N_16978);
nand U17059 (N_17059,N_16935,N_16826);
xnor U17060 (N_17060,N_16871,N_16945);
or U17061 (N_17061,N_16930,N_16873);
nand U17062 (N_17062,N_16986,N_16884);
nor U17063 (N_17063,N_16892,N_16851);
nand U17064 (N_17064,N_16890,N_16970);
or U17065 (N_17065,N_16811,N_16951);
xor U17066 (N_17066,N_16833,N_16938);
xnor U17067 (N_17067,N_16920,N_16872);
xor U17068 (N_17068,N_16827,N_16842);
nand U17069 (N_17069,N_16866,N_16975);
or U17070 (N_17070,N_16844,N_16820);
nor U17071 (N_17071,N_16944,N_16824);
nand U17072 (N_17072,N_16822,N_16882);
xor U17073 (N_17073,N_16896,N_16821);
nor U17074 (N_17074,N_16874,N_16981);
nand U17075 (N_17075,N_16831,N_16928);
and U17076 (N_17076,N_16914,N_16847);
or U17077 (N_17077,N_16862,N_16835);
nor U17078 (N_17078,N_16964,N_16880);
nor U17079 (N_17079,N_16908,N_16838);
nor U17080 (N_17080,N_16904,N_16853);
xor U17081 (N_17081,N_16829,N_16865);
and U17082 (N_17082,N_16910,N_16808);
nor U17083 (N_17083,N_16916,N_16878);
or U17084 (N_17084,N_16813,N_16969);
and U17085 (N_17085,N_16860,N_16940);
nand U17086 (N_17086,N_16965,N_16921);
nand U17087 (N_17087,N_16858,N_16946);
nor U17088 (N_17088,N_16912,N_16898);
and U17089 (N_17089,N_16954,N_16941);
or U17090 (N_17090,N_16974,N_16919);
and U17091 (N_17091,N_16815,N_16924);
and U17092 (N_17092,N_16867,N_16923);
nand U17093 (N_17093,N_16850,N_16931);
nor U17094 (N_17094,N_16869,N_16977);
xnor U17095 (N_17095,N_16936,N_16856);
xnor U17096 (N_17096,N_16830,N_16802);
nand U17097 (N_17097,N_16949,N_16994);
nand U17098 (N_17098,N_16971,N_16883);
nor U17099 (N_17099,N_16845,N_16807);
nand U17100 (N_17100,N_16964,N_16892);
nand U17101 (N_17101,N_16972,N_16892);
nand U17102 (N_17102,N_16888,N_16827);
and U17103 (N_17103,N_16851,N_16883);
nand U17104 (N_17104,N_16807,N_16947);
nor U17105 (N_17105,N_16962,N_16822);
nand U17106 (N_17106,N_16871,N_16971);
xnor U17107 (N_17107,N_16849,N_16819);
xnor U17108 (N_17108,N_16800,N_16946);
and U17109 (N_17109,N_16983,N_16868);
xor U17110 (N_17110,N_16964,N_16928);
nor U17111 (N_17111,N_16969,N_16889);
xnor U17112 (N_17112,N_16816,N_16851);
or U17113 (N_17113,N_16876,N_16975);
or U17114 (N_17114,N_16826,N_16941);
and U17115 (N_17115,N_16991,N_16931);
and U17116 (N_17116,N_16912,N_16991);
nor U17117 (N_17117,N_16815,N_16913);
or U17118 (N_17118,N_16967,N_16874);
nand U17119 (N_17119,N_16956,N_16982);
and U17120 (N_17120,N_16837,N_16829);
nand U17121 (N_17121,N_16886,N_16924);
or U17122 (N_17122,N_16885,N_16973);
xor U17123 (N_17123,N_16962,N_16985);
nand U17124 (N_17124,N_16906,N_16967);
nand U17125 (N_17125,N_16885,N_16851);
and U17126 (N_17126,N_16920,N_16939);
and U17127 (N_17127,N_16937,N_16971);
and U17128 (N_17128,N_16914,N_16866);
nor U17129 (N_17129,N_16944,N_16985);
nand U17130 (N_17130,N_16926,N_16904);
nand U17131 (N_17131,N_16802,N_16891);
and U17132 (N_17132,N_16945,N_16830);
xor U17133 (N_17133,N_16902,N_16889);
nor U17134 (N_17134,N_16907,N_16988);
and U17135 (N_17135,N_16809,N_16905);
and U17136 (N_17136,N_16910,N_16989);
and U17137 (N_17137,N_16821,N_16883);
nor U17138 (N_17138,N_16858,N_16893);
nor U17139 (N_17139,N_16903,N_16831);
nand U17140 (N_17140,N_16859,N_16944);
and U17141 (N_17141,N_16877,N_16913);
xor U17142 (N_17142,N_16869,N_16909);
nor U17143 (N_17143,N_16991,N_16894);
or U17144 (N_17144,N_16929,N_16847);
or U17145 (N_17145,N_16822,N_16971);
xor U17146 (N_17146,N_16873,N_16935);
or U17147 (N_17147,N_16919,N_16965);
and U17148 (N_17148,N_16889,N_16942);
nand U17149 (N_17149,N_16864,N_16984);
xnor U17150 (N_17150,N_16809,N_16980);
nand U17151 (N_17151,N_16842,N_16838);
nor U17152 (N_17152,N_16992,N_16870);
xnor U17153 (N_17153,N_16829,N_16838);
nand U17154 (N_17154,N_16893,N_16984);
and U17155 (N_17155,N_16989,N_16997);
nand U17156 (N_17156,N_16894,N_16928);
and U17157 (N_17157,N_16888,N_16867);
xor U17158 (N_17158,N_16950,N_16989);
or U17159 (N_17159,N_16843,N_16815);
and U17160 (N_17160,N_16864,N_16976);
xnor U17161 (N_17161,N_16933,N_16876);
and U17162 (N_17162,N_16967,N_16805);
or U17163 (N_17163,N_16803,N_16911);
or U17164 (N_17164,N_16954,N_16979);
nand U17165 (N_17165,N_16923,N_16991);
nand U17166 (N_17166,N_16817,N_16843);
nand U17167 (N_17167,N_16820,N_16922);
nor U17168 (N_17168,N_16811,N_16954);
nand U17169 (N_17169,N_16826,N_16987);
nand U17170 (N_17170,N_16993,N_16991);
nor U17171 (N_17171,N_16865,N_16819);
nand U17172 (N_17172,N_16908,N_16939);
nor U17173 (N_17173,N_16826,N_16816);
nor U17174 (N_17174,N_16998,N_16924);
nand U17175 (N_17175,N_16990,N_16853);
xnor U17176 (N_17176,N_16977,N_16938);
xor U17177 (N_17177,N_16864,N_16909);
or U17178 (N_17178,N_16820,N_16982);
and U17179 (N_17179,N_16931,N_16812);
or U17180 (N_17180,N_16823,N_16880);
nor U17181 (N_17181,N_16967,N_16916);
xor U17182 (N_17182,N_16948,N_16809);
nand U17183 (N_17183,N_16927,N_16898);
nor U17184 (N_17184,N_16800,N_16826);
nand U17185 (N_17185,N_16918,N_16966);
and U17186 (N_17186,N_16858,N_16867);
nor U17187 (N_17187,N_16863,N_16857);
nand U17188 (N_17188,N_16831,N_16857);
or U17189 (N_17189,N_16875,N_16879);
nor U17190 (N_17190,N_16809,N_16956);
xor U17191 (N_17191,N_16872,N_16891);
or U17192 (N_17192,N_16867,N_16936);
nand U17193 (N_17193,N_16921,N_16907);
xor U17194 (N_17194,N_16892,N_16959);
and U17195 (N_17195,N_16928,N_16957);
or U17196 (N_17196,N_16993,N_16866);
nor U17197 (N_17197,N_16811,N_16827);
or U17198 (N_17198,N_16989,N_16995);
nand U17199 (N_17199,N_16924,N_16807);
or U17200 (N_17200,N_17066,N_17100);
or U17201 (N_17201,N_17162,N_17133);
or U17202 (N_17202,N_17134,N_17157);
nand U17203 (N_17203,N_17171,N_17011);
or U17204 (N_17204,N_17160,N_17057);
and U17205 (N_17205,N_17056,N_17074);
nand U17206 (N_17206,N_17181,N_17075);
nor U17207 (N_17207,N_17091,N_17029);
nor U17208 (N_17208,N_17048,N_17019);
nand U17209 (N_17209,N_17197,N_17046);
or U17210 (N_17210,N_17071,N_17077);
nor U17211 (N_17211,N_17065,N_17002);
and U17212 (N_17212,N_17190,N_17185);
xor U17213 (N_17213,N_17158,N_17062);
nand U17214 (N_17214,N_17047,N_17052);
nand U17215 (N_17215,N_17196,N_17055);
or U17216 (N_17216,N_17189,N_17131);
and U17217 (N_17217,N_17126,N_17170);
or U17218 (N_17218,N_17164,N_17166);
and U17219 (N_17219,N_17043,N_17012);
xor U17220 (N_17220,N_17022,N_17099);
or U17221 (N_17221,N_17060,N_17027);
nand U17222 (N_17222,N_17064,N_17005);
nor U17223 (N_17223,N_17081,N_17184);
nand U17224 (N_17224,N_17146,N_17032);
and U17225 (N_17225,N_17087,N_17169);
nand U17226 (N_17226,N_17036,N_17021);
or U17227 (N_17227,N_17173,N_17085);
or U17228 (N_17228,N_17199,N_17030);
nand U17229 (N_17229,N_17063,N_17093);
xor U17230 (N_17230,N_17183,N_17023);
xnor U17231 (N_17231,N_17038,N_17165);
nand U17232 (N_17232,N_17139,N_17026);
xor U17233 (N_17233,N_17051,N_17000);
nand U17234 (N_17234,N_17084,N_17006);
and U17235 (N_17235,N_17128,N_17145);
xor U17236 (N_17236,N_17059,N_17167);
nand U17237 (N_17237,N_17110,N_17122);
xor U17238 (N_17238,N_17001,N_17086);
or U17239 (N_17239,N_17016,N_17194);
or U17240 (N_17240,N_17013,N_17130);
xnor U17241 (N_17241,N_17049,N_17034);
xor U17242 (N_17242,N_17187,N_17193);
and U17243 (N_17243,N_17125,N_17121);
xor U17244 (N_17244,N_17061,N_17109);
and U17245 (N_17245,N_17092,N_17089);
or U17246 (N_17246,N_17140,N_17035);
xnor U17247 (N_17247,N_17094,N_17191);
nor U17248 (N_17248,N_17152,N_17142);
and U17249 (N_17249,N_17143,N_17117);
nor U17250 (N_17250,N_17174,N_17147);
xor U17251 (N_17251,N_17179,N_17040);
xor U17252 (N_17252,N_17186,N_17020);
nor U17253 (N_17253,N_17105,N_17192);
and U17254 (N_17254,N_17028,N_17102);
nor U17255 (N_17255,N_17096,N_17163);
xor U17256 (N_17256,N_17082,N_17113);
xor U17257 (N_17257,N_17076,N_17120);
or U17258 (N_17258,N_17115,N_17106);
nand U17259 (N_17259,N_17114,N_17041);
xor U17260 (N_17260,N_17018,N_17175);
and U17261 (N_17261,N_17031,N_17172);
nand U17262 (N_17262,N_17072,N_17009);
and U17263 (N_17263,N_17010,N_17083);
nand U17264 (N_17264,N_17111,N_17182);
nor U17265 (N_17265,N_17042,N_17150);
xnor U17266 (N_17266,N_17015,N_17195);
nor U17267 (N_17267,N_17073,N_17141);
or U17268 (N_17268,N_17149,N_17078);
nor U17269 (N_17269,N_17025,N_17119);
nand U17270 (N_17270,N_17104,N_17098);
nor U17271 (N_17271,N_17129,N_17124);
nand U17272 (N_17272,N_17156,N_17135);
nor U17273 (N_17273,N_17050,N_17178);
xnor U17274 (N_17274,N_17008,N_17123);
nor U17275 (N_17275,N_17198,N_17067);
nand U17276 (N_17276,N_17037,N_17103);
nand U17277 (N_17277,N_17017,N_17097);
or U17278 (N_17278,N_17161,N_17044);
or U17279 (N_17279,N_17132,N_17180);
or U17280 (N_17280,N_17159,N_17058);
or U17281 (N_17281,N_17024,N_17053);
xor U17282 (N_17282,N_17004,N_17088);
or U17283 (N_17283,N_17188,N_17153);
xnor U17284 (N_17284,N_17045,N_17069);
nand U17285 (N_17285,N_17148,N_17079);
xor U17286 (N_17286,N_17014,N_17138);
or U17287 (N_17287,N_17039,N_17068);
nand U17288 (N_17288,N_17090,N_17007);
and U17289 (N_17289,N_17168,N_17176);
xor U17290 (N_17290,N_17154,N_17137);
and U17291 (N_17291,N_17095,N_17112);
nor U17292 (N_17292,N_17033,N_17107);
xor U17293 (N_17293,N_17080,N_17136);
and U17294 (N_17294,N_17127,N_17155);
or U17295 (N_17295,N_17070,N_17116);
and U17296 (N_17296,N_17177,N_17151);
nand U17297 (N_17297,N_17144,N_17118);
xnor U17298 (N_17298,N_17108,N_17054);
and U17299 (N_17299,N_17101,N_17003);
and U17300 (N_17300,N_17099,N_17111);
xor U17301 (N_17301,N_17185,N_17140);
or U17302 (N_17302,N_17012,N_17013);
and U17303 (N_17303,N_17164,N_17030);
and U17304 (N_17304,N_17190,N_17021);
xnor U17305 (N_17305,N_17125,N_17187);
nand U17306 (N_17306,N_17047,N_17048);
and U17307 (N_17307,N_17089,N_17039);
nand U17308 (N_17308,N_17093,N_17135);
nor U17309 (N_17309,N_17057,N_17195);
and U17310 (N_17310,N_17082,N_17067);
nand U17311 (N_17311,N_17119,N_17160);
nand U17312 (N_17312,N_17010,N_17154);
and U17313 (N_17313,N_17048,N_17096);
or U17314 (N_17314,N_17063,N_17173);
and U17315 (N_17315,N_17148,N_17197);
or U17316 (N_17316,N_17146,N_17087);
nor U17317 (N_17317,N_17154,N_17045);
and U17318 (N_17318,N_17091,N_17062);
or U17319 (N_17319,N_17184,N_17040);
xor U17320 (N_17320,N_17195,N_17096);
nor U17321 (N_17321,N_17167,N_17163);
nand U17322 (N_17322,N_17193,N_17171);
or U17323 (N_17323,N_17084,N_17107);
nand U17324 (N_17324,N_17132,N_17192);
and U17325 (N_17325,N_17191,N_17185);
xor U17326 (N_17326,N_17125,N_17111);
and U17327 (N_17327,N_17060,N_17014);
nor U17328 (N_17328,N_17197,N_17156);
nand U17329 (N_17329,N_17015,N_17037);
and U17330 (N_17330,N_17077,N_17045);
nand U17331 (N_17331,N_17111,N_17102);
nor U17332 (N_17332,N_17144,N_17019);
nand U17333 (N_17333,N_17142,N_17073);
nor U17334 (N_17334,N_17013,N_17192);
and U17335 (N_17335,N_17068,N_17145);
nand U17336 (N_17336,N_17198,N_17066);
or U17337 (N_17337,N_17063,N_17088);
and U17338 (N_17338,N_17086,N_17056);
and U17339 (N_17339,N_17131,N_17194);
and U17340 (N_17340,N_17127,N_17102);
or U17341 (N_17341,N_17084,N_17162);
nand U17342 (N_17342,N_17092,N_17122);
or U17343 (N_17343,N_17054,N_17030);
nor U17344 (N_17344,N_17084,N_17148);
xnor U17345 (N_17345,N_17058,N_17064);
nand U17346 (N_17346,N_17152,N_17055);
nor U17347 (N_17347,N_17010,N_17136);
nand U17348 (N_17348,N_17116,N_17194);
nand U17349 (N_17349,N_17174,N_17139);
and U17350 (N_17350,N_17186,N_17074);
nand U17351 (N_17351,N_17081,N_17058);
and U17352 (N_17352,N_17081,N_17040);
xor U17353 (N_17353,N_17057,N_17089);
nor U17354 (N_17354,N_17186,N_17083);
nand U17355 (N_17355,N_17198,N_17116);
xor U17356 (N_17356,N_17036,N_17054);
or U17357 (N_17357,N_17061,N_17042);
nand U17358 (N_17358,N_17099,N_17100);
nor U17359 (N_17359,N_17090,N_17047);
or U17360 (N_17360,N_17154,N_17152);
xnor U17361 (N_17361,N_17140,N_17169);
or U17362 (N_17362,N_17025,N_17087);
or U17363 (N_17363,N_17078,N_17145);
or U17364 (N_17364,N_17140,N_17014);
and U17365 (N_17365,N_17175,N_17122);
nor U17366 (N_17366,N_17163,N_17093);
nor U17367 (N_17367,N_17041,N_17022);
xor U17368 (N_17368,N_17197,N_17102);
or U17369 (N_17369,N_17003,N_17134);
nor U17370 (N_17370,N_17077,N_17055);
and U17371 (N_17371,N_17154,N_17044);
nor U17372 (N_17372,N_17020,N_17051);
nand U17373 (N_17373,N_17188,N_17050);
xor U17374 (N_17374,N_17082,N_17050);
and U17375 (N_17375,N_17181,N_17097);
nand U17376 (N_17376,N_17132,N_17155);
nor U17377 (N_17377,N_17160,N_17084);
or U17378 (N_17378,N_17043,N_17054);
xor U17379 (N_17379,N_17048,N_17085);
and U17380 (N_17380,N_17060,N_17159);
nor U17381 (N_17381,N_17186,N_17034);
or U17382 (N_17382,N_17178,N_17109);
nand U17383 (N_17383,N_17031,N_17099);
and U17384 (N_17384,N_17124,N_17123);
xnor U17385 (N_17385,N_17147,N_17021);
and U17386 (N_17386,N_17187,N_17109);
or U17387 (N_17387,N_17114,N_17144);
nor U17388 (N_17388,N_17173,N_17080);
nand U17389 (N_17389,N_17021,N_17143);
and U17390 (N_17390,N_17176,N_17074);
xor U17391 (N_17391,N_17137,N_17063);
nand U17392 (N_17392,N_17183,N_17006);
nand U17393 (N_17393,N_17008,N_17035);
or U17394 (N_17394,N_17055,N_17048);
and U17395 (N_17395,N_17130,N_17169);
and U17396 (N_17396,N_17013,N_17001);
xnor U17397 (N_17397,N_17003,N_17178);
or U17398 (N_17398,N_17094,N_17074);
or U17399 (N_17399,N_17014,N_17065);
nor U17400 (N_17400,N_17341,N_17209);
nor U17401 (N_17401,N_17231,N_17354);
xor U17402 (N_17402,N_17309,N_17291);
nand U17403 (N_17403,N_17284,N_17299);
xnor U17404 (N_17404,N_17232,N_17392);
nor U17405 (N_17405,N_17337,N_17347);
or U17406 (N_17406,N_17246,N_17338);
and U17407 (N_17407,N_17286,N_17377);
nand U17408 (N_17408,N_17273,N_17224);
xnor U17409 (N_17409,N_17390,N_17313);
nand U17410 (N_17410,N_17201,N_17305);
and U17411 (N_17411,N_17387,N_17397);
or U17412 (N_17412,N_17367,N_17346);
nor U17413 (N_17413,N_17202,N_17311);
nand U17414 (N_17414,N_17215,N_17205);
nor U17415 (N_17415,N_17266,N_17385);
nand U17416 (N_17416,N_17372,N_17348);
nand U17417 (N_17417,N_17344,N_17303);
or U17418 (N_17418,N_17359,N_17378);
or U17419 (N_17419,N_17331,N_17362);
xnor U17420 (N_17420,N_17389,N_17342);
and U17421 (N_17421,N_17376,N_17307);
xnor U17422 (N_17422,N_17319,N_17276);
or U17423 (N_17423,N_17265,N_17287);
nand U17424 (N_17424,N_17290,N_17351);
nor U17425 (N_17425,N_17203,N_17261);
xor U17426 (N_17426,N_17358,N_17398);
nor U17427 (N_17427,N_17332,N_17235);
xor U17428 (N_17428,N_17393,N_17256);
nor U17429 (N_17429,N_17335,N_17289);
nor U17430 (N_17430,N_17249,N_17345);
xnor U17431 (N_17431,N_17292,N_17223);
nand U17432 (N_17432,N_17322,N_17254);
xor U17433 (N_17433,N_17356,N_17381);
xnor U17434 (N_17434,N_17352,N_17315);
nor U17435 (N_17435,N_17300,N_17302);
and U17436 (N_17436,N_17366,N_17257);
or U17437 (N_17437,N_17304,N_17214);
nor U17438 (N_17438,N_17251,N_17281);
xor U17439 (N_17439,N_17317,N_17274);
nand U17440 (N_17440,N_17343,N_17386);
nor U17441 (N_17441,N_17239,N_17270);
nand U17442 (N_17442,N_17253,N_17295);
nor U17443 (N_17443,N_17207,N_17321);
xnor U17444 (N_17444,N_17339,N_17260);
or U17445 (N_17445,N_17259,N_17395);
xor U17446 (N_17446,N_17320,N_17382);
nor U17447 (N_17447,N_17380,N_17245);
nor U17448 (N_17448,N_17237,N_17255);
nand U17449 (N_17449,N_17241,N_17220);
nor U17450 (N_17450,N_17364,N_17388);
or U17451 (N_17451,N_17250,N_17244);
nor U17452 (N_17452,N_17350,N_17211);
or U17453 (N_17453,N_17399,N_17233);
nor U17454 (N_17454,N_17204,N_17258);
nand U17455 (N_17455,N_17323,N_17324);
or U17456 (N_17456,N_17328,N_17293);
nand U17457 (N_17457,N_17333,N_17221);
xor U17458 (N_17458,N_17275,N_17310);
xor U17459 (N_17459,N_17210,N_17368);
nor U17460 (N_17460,N_17247,N_17282);
xor U17461 (N_17461,N_17361,N_17213);
or U17462 (N_17462,N_17327,N_17252);
xnor U17463 (N_17463,N_17242,N_17271);
and U17464 (N_17464,N_17312,N_17285);
nand U17465 (N_17465,N_17228,N_17325);
and U17466 (N_17466,N_17314,N_17301);
and U17467 (N_17467,N_17208,N_17225);
xnor U17468 (N_17468,N_17283,N_17272);
nor U17469 (N_17469,N_17217,N_17297);
nand U17470 (N_17470,N_17206,N_17316);
nand U17471 (N_17471,N_17218,N_17234);
nor U17472 (N_17472,N_17216,N_17391);
xor U17473 (N_17473,N_17353,N_17280);
or U17474 (N_17474,N_17371,N_17263);
xor U17475 (N_17475,N_17298,N_17326);
or U17476 (N_17476,N_17396,N_17240);
or U17477 (N_17477,N_17383,N_17369);
and U17478 (N_17478,N_17264,N_17212);
or U17479 (N_17479,N_17355,N_17288);
nor U17480 (N_17480,N_17278,N_17394);
and U17481 (N_17481,N_17330,N_17230);
or U17482 (N_17482,N_17226,N_17349);
nand U17483 (N_17483,N_17267,N_17363);
xnor U17484 (N_17484,N_17296,N_17357);
xor U17485 (N_17485,N_17200,N_17334);
nor U17486 (N_17486,N_17370,N_17279);
nand U17487 (N_17487,N_17375,N_17238);
xor U17488 (N_17488,N_17219,N_17248);
or U17489 (N_17489,N_17269,N_17308);
or U17490 (N_17490,N_17318,N_17340);
nor U17491 (N_17491,N_17329,N_17236);
nand U17492 (N_17492,N_17379,N_17373);
nand U17493 (N_17493,N_17374,N_17229);
nor U17494 (N_17494,N_17360,N_17277);
nand U17495 (N_17495,N_17306,N_17227);
xnor U17496 (N_17496,N_17262,N_17268);
or U17497 (N_17497,N_17336,N_17384);
or U17498 (N_17498,N_17222,N_17365);
xor U17499 (N_17499,N_17243,N_17294);
nand U17500 (N_17500,N_17209,N_17275);
or U17501 (N_17501,N_17333,N_17349);
nand U17502 (N_17502,N_17215,N_17354);
and U17503 (N_17503,N_17235,N_17352);
nand U17504 (N_17504,N_17266,N_17201);
and U17505 (N_17505,N_17352,N_17245);
nor U17506 (N_17506,N_17215,N_17282);
or U17507 (N_17507,N_17215,N_17387);
nand U17508 (N_17508,N_17288,N_17245);
or U17509 (N_17509,N_17212,N_17365);
xnor U17510 (N_17510,N_17318,N_17392);
or U17511 (N_17511,N_17297,N_17388);
and U17512 (N_17512,N_17261,N_17322);
and U17513 (N_17513,N_17379,N_17222);
nand U17514 (N_17514,N_17335,N_17240);
nor U17515 (N_17515,N_17392,N_17279);
and U17516 (N_17516,N_17350,N_17272);
or U17517 (N_17517,N_17316,N_17310);
or U17518 (N_17518,N_17364,N_17289);
nand U17519 (N_17519,N_17203,N_17304);
nor U17520 (N_17520,N_17348,N_17345);
nand U17521 (N_17521,N_17239,N_17283);
and U17522 (N_17522,N_17260,N_17364);
nor U17523 (N_17523,N_17266,N_17239);
nor U17524 (N_17524,N_17231,N_17374);
xnor U17525 (N_17525,N_17281,N_17302);
or U17526 (N_17526,N_17332,N_17311);
and U17527 (N_17527,N_17216,N_17266);
xor U17528 (N_17528,N_17201,N_17323);
and U17529 (N_17529,N_17367,N_17229);
nand U17530 (N_17530,N_17323,N_17213);
nand U17531 (N_17531,N_17253,N_17336);
or U17532 (N_17532,N_17285,N_17337);
and U17533 (N_17533,N_17210,N_17393);
nor U17534 (N_17534,N_17308,N_17310);
nor U17535 (N_17535,N_17213,N_17262);
xor U17536 (N_17536,N_17391,N_17290);
and U17537 (N_17537,N_17233,N_17281);
nor U17538 (N_17538,N_17282,N_17297);
or U17539 (N_17539,N_17326,N_17379);
and U17540 (N_17540,N_17399,N_17338);
or U17541 (N_17541,N_17325,N_17363);
xor U17542 (N_17542,N_17210,N_17342);
or U17543 (N_17543,N_17206,N_17268);
nor U17544 (N_17544,N_17229,N_17293);
or U17545 (N_17545,N_17222,N_17316);
nand U17546 (N_17546,N_17325,N_17289);
or U17547 (N_17547,N_17367,N_17368);
and U17548 (N_17548,N_17254,N_17307);
and U17549 (N_17549,N_17334,N_17382);
nand U17550 (N_17550,N_17361,N_17316);
or U17551 (N_17551,N_17326,N_17391);
xnor U17552 (N_17552,N_17319,N_17300);
nor U17553 (N_17553,N_17333,N_17297);
or U17554 (N_17554,N_17231,N_17397);
xnor U17555 (N_17555,N_17341,N_17304);
or U17556 (N_17556,N_17267,N_17300);
or U17557 (N_17557,N_17370,N_17246);
or U17558 (N_17558,N_17256,N_17328);
and U17559 (N_17559,N_17301,N_17267);
and U17560 (N_17560,N_17399,N_17223);
and U17561 (N_17561,N_17312,N_17211);
or U17562 (N_17562,N_17290,N_17320);
xor U17563 (N_17563,N_17389,N_17204);
or U17564 (N_17564,N_17389,N_17287);
xnor U17565 (N_17565,N_17399,N_17230);
and U17566 (N_17566,N_17302,N_17295);
or U17567 (N_17567,N_17324,N_17207);
xnor U17568 (N_17568,N_17268,N_17315);
nand U17569 (N_17569,N_17286,N_17371);
xor U17570 (N_17570,N_17370,N_17248);
xnor U17571 (N_17571,N_17200,N_17301);
xnor U17572 (N_17572,N_17399,N_17322);
or U17573 (N_17573,N_17275,N_17365);
or U17574 (N_17574,N_17287,N_17288);
or U17575 (N_17575,N_17319,N_17225);
or U17576 (N_17576,N_17387,N_17231);
and U17577 (N_17577,N_17371,N_17363);
xor U17578 (N_17578,N_17214,N_17322);
xor U17579 (N_17579,N_17216,N_17287);
or U17580 (N_17580,N_17366,N_17335);
xor U17581 (N_17581,N_17285,N_17384);
or U17582 (N_17582,N_17359,N_17390);
nor U17583 (N_17583,N_17219,N_17285);
xor U17584 (N_17584,N_17313,N_17239);
nand U17585 (N_17585,N_17254,N_17200);
and U17586 (N_17586,N_17319,N_17268);
or U17587 (N_17587,N_17307,N_17220);
xnor U17588 (N_17588,N_17282,N_17335);
nor U17589 (N_17589,N_17396,N_17306);
nor U17590 (N_17590,N_17245,N_17238);
nand U17591 (N_17591,N_17216,N_17304);
nand U17592 (N_17592,N_17283,N_17360);
or U17593 (N_17593,N_17354,N_17208);
xor U17594 (N_17594,N_17252,N_17213);
nand U17595 (N_17595,N_17373,N_17358);
nand U17596 (N_17596,N_17214,N_17303);
or U17597 (N_17597,N_17219,N_17282);
nor U17598 (N_17598,N_17367,N_17399);
and U17599 (N_17599,N_17398,N_17285);
xor U17600 (N_17600,N_17428,N_17483);
and U17601 (N_17601,N_17429,N_17595);
nand U17602 (N_17602,N_17476,N_17516);
xor U17603 (N_17603,N_17419,N_17569);
and U17604 (N_17604,N_17471,N_17507);
or U17605 (N_17605,N_17518,N_17548);
and U17606 (N_17606,N_17404,N_17413);
nand U17607 (N_17607,N_17453,N_17547);
nand U17608 (N_17608,N_17524,N_17436);
and U17609 (N_17609,N_17564,N_17540);
nor U17610 (N_17610,N_17552,N_17583);
and U17611 (N_17611,N_17504,N_17514);
and U17612 (N_17612,N_17489,N_17472);
or U17613 (N_17613,N_17508,N_17458);
nor U17614 (N_17614,N_17588,N_17491);
and U17615 (N_17615,N_17573,N_17561);
nor U17616 (N_17616,N_17537,N_17584);
and U17617 (N_17617,N_17481,N_17401);
nand U17618 (N_17618,N_17410,N_17593);
and U17619 (N_17619,N_17551,N_17509);
or U17620 (N_17620,N_17434,N_17598);
and U17621 (N_17621,N_17443,N_17579);
or U17622 (N_17622,N_17446,N_17455);
or U17623 (N_17623,N_17546,N_17486);
and U17624 (N_17624,N_17535,N_17506);
nand U17625 (N_17625,N_17441,N_17529);
xor U17626 (N_17626,N_17580,N_17502);
nand U17627 (N_17627,N_17469,N_17526);
or U17628 (N_17628,N_17478,N_17543);
nand U17629 (N_17629,N_17575,N_17542);
and U17630 (N_17630,N_17566,N_17406);
and U17631 (N_17631,N_17534,N_17517);
nand U17632 (N_17632,N_17556,N_17470);
xnor U17633 (N_17633,N_17400,N_17444);
nand U17634 (N_17634,N_17468,N_17586);
and U17635 (N_17635,N_17565,N_17467);
xor U17636 (N_17636,N_17431,N_17505);
and U17637 (N_17637,N_17432,N_17480);
xnor U17638 (N_17638,N_17488,N_17430);
nand U17639 (N_17639,N_17555,N_17525);
xnor U17640 (N_17640,N_17578,N_17545);
and U17641 (N_17641,N_17426,N_17485);
xnor U17642 (N_17642,N_17450,N_17590);
nand U17643 (N_17643,N_17459,N_17597);
or U17644 (N_17644,N_17541,N_17527);
and U17645 (N_17645,N_17574,N_17511);
and U17646 (N_17646,N_17528,N_17570);
and U17647 (N_17647,N_17493,N_17412);
nor U17648 (N_17648,N_17563,N_17449);
xor U17649 (N_17649,N_17587,N_17568);
xnor U17650 (N_17650,N_17463,N_17560);
nor U17651 (N_17651,N_17479,N_17451);
and U17652 (N_17652,N_17503,N_17460);
or U17653 (N_17653,N_17531,N_17420);
nand U17654 (N_17654,N_17482,N_17425);
xnor U17655 (N_17655,N_17553,N_17512);
nor U17656 (N_17656,N_17572,N_17409);
nand U17657 (N_17657,N_17440,N_17496);
xnor U17658 (N_17658,N_17501,N_17442);
or U17659 (N_17659,N_17473,N_17427);
nor U17660 (N_17660,N_17510,N_17464);
nor U17661 (N_17661,N_17549,N_17550);
and U17662 (N_17662,N_17592,N_17474);
nand U17663 (N_17663,N_17424,N_17421);
xnor U17664 (N_17664,N_17402,N_17437);
nor U17665 (N_17665,N_17554,N_17417);
xnor U17666 (N_17666,N_17523,N_17414);
xor U17667 (N_17667,N_17591,N_17559);
xnor U17668 (N_17668,N_17533,N_17416);
xor U17669 (N_17669,N_17596,N_17405);
nor U17670 (N_17670,N_17521,N_17466);
and U17671 (N_17671,N_17484,N_17562);
nand U17672 (N_17672,N_17495,N_17519);
and U17673 (N_17673,N_17522,N_17577);
xnor U17674 (N_17674,N_17515,N_17492);
or U17675 (N_17675,N_17544,N_17490);
nand U17676 (N_17676,N_17438,N_17445);
xnor U17677 (N_17677,N_17456,N_17448);
nand U17678 (N_17678,N_17403,N_17520);
and U17679 (N_17679,N_17477,N_17494);
and U17680 (N_17680,N_17557,N_17408);
or U17681 (N_17681,N_17576,N_17599);
xor U17682 (N_17682,N_17418,N_17558);
or U17683 (N_17683,N_17447,N_17589);
or U17684 (N_17684,N_17513,N_17500);
nand U17685 (N_17685,N_17435,N_17567);
or U17686 (N_17686,N_17487,N_17433);
nand U17687 (N_17687,N_17461,N_17465);
or U17688 (N_17688,N_17407,N_17538);
nor U17689 (N_17689,N_17539,N_17498);
or U17690 (N_17690,N_17497,N_17582);
xor U17691 (N_17691,N_17594,N_17439);
or U17692 (N_17692,N_17475,N_17462);
xnor U17693 (N_17693,N_17530,N_17532);
or U17694 (N_17694,N_17457,N_17581);
nand U17695 (N_17695,N_17499,N_17423);
xnor U17696 (N_17696,N_17585,N_17571);
nand U17697 (N_17697,N_17536,N_17452);
nor U17698 (N_17698,N_17411,N_17454);
nor U17699 (N_17699,N_17422,N_17415);
xor U17700 (N_17700,N_17456,N_17533);
xor U17701 (N_17701,N_17586,N_17532);
nand U17702 (N_17702,N_17577,N_17493);
xor U17703 (N_17703,N_17587,N_17454);
xnor U17704 (N_17704,N_17514,N_17585);
xor U17705 (N_17705,N_17529,N_17520);
nand U17706 (N_17706,N_17471,N_17524);
xnor U17707 (N_17707,N_17422,N_17523);
and U17708 (N_17708,N_17477,N_17457);
or U17709 (N_17709,N_17509,N_17569);
or U17710 (N_17710,N_17522,N_17438);
nand U17711 (N_17711,N_17577,N_17435);
nor U17712 (N_17712,N_17512,N_17563);
or U17713 (N_17713,N_17534,N_17402);
xor U17714 (N_17714,N_17450,N_17521);
or U17715 (N_17715,N_17449,N_17530);
or U17716 (N_17716,N_17483,N_17404);
or U17717 (N_17717,N_17485,N_17421);
and U17718 (N_17718,N_17533,N_17491);
nand U17719 (N_17719,N_17437,N_17466);
nand U17720 (N_17720,N_17441,N_17463);
and U17721 (N_17721,N_17518,N_17532);
nor U17722 (N_17722,N_17548,N_17459);
nor U17723 (N_17723,N_17511,N_17552);
and U17724 (N_17724,N_17490,N_17434);
nor U17725 (N_17725,N_17508,N_17522);
or U17726 (N_17726,N_17556,N_17526);
nand U17727 (N_17727,N_17458,N_17412);
xnor U17728 (N_17728,N_17578,N_17434);
or U17729 (N_17729,N_17427,N_17591);
nand U17730 (N_17730,N_17450,N_17445);
and U17731 (N_17731,N_17478,N_17482);
or U17732 (N_17732,N_17556,N_17435);
nand U17733 (N_17733,N_17517,N_17555);
and U17734 (N_17734,N_17532,N_17564);
and U17735 (N_17735,N_17558,N_17555);
xnor U17736 (N_17736,N_17464,N_17537);
xnor U17737 (N_17737,N_17570,N_17581);
nand U17738 (N_17738,N_17485,N_17585);
nand U17739 (N_17739,N_17529,N_17424);
or U17740 (N_17740,N_17496,N_17564);
xnor U17741 (N_17741,N_17436,N_17533);
nor U17742 (N_17742,N_17584,N_17525);
nand U17743 (N_17743,N_17445,N_17517);
and U17744 (N_17744,N_17420,N_17403);
or U17745 (N_17745,N_17419,N_17468);
and U17746 (N_17746,N_17433,N_17510);
or U17747 (N_17747,N_17562,N_17561);
or U17748 (N_17748,N_17582,N_17474);
and U17749 (N_17749,N_17412,N_17520);
or U17750 (N_17750,N_17538,N_17520);
nand U17751 (N_17751,N_17422,N_17451);
nor U17752 (N_17752,N_17498,N_17528);
and U17753 (N_17753,N_17520,N_17548);
nand U17754 (N_17754,N_17516,N_17523);
nor U17755 (N_17755,N_17451,N_17431);
nand U17756 (N_17756,N_17458,N_17465);
or U17757 (N_17757,N_17517,N_17459);
xor U17758 (N_17758,N_17571,N_17509);
or U17759 (N_17759,N_17420,N_17418);
xnor U17760 (N_17760,N_17568,N_17478);
nand U17761 (N_17761,N_17458,N_17542);
xnor U17762 (N_17762,N_17410,N_17434);
and U17763 (N_17763,N_17545,N_17583);
nand U17764 (N_17764,N_17402,N_17509);
nand U17765 (N_17765,N_17596,N_17510);
nor U17766 (N_17766,N_17518,N_17574);
and U17767 (N_17767,N_17497,N_17530);
nor U17768 (N_17768,N_17483,N_17429);
nand U17769 (N_17769,N_17400,N_17565);
xor U17770 (N_17770,N_17409,N_17525);
nor U17771 (N_17771,N_17432,N_17552);
and U17772 (N_17772,N_17528,N_17468);
nand U17773 (N_17773,N_17516,N_17515);
xor U17774 (N_17774,N_17488,N_17420);
nand U17775 (N_17775,N_17551,N_17512);
and U17776 (N_17776,N_17407,N_17430);
or U17777 (N_17777,N_17409,N_17510);
xor U17778 (N_17778,N_17456,N_17566);
or U17779 (N_17779,N_17516,N_17594);
xnor U17780 (N_17780,N_17485,N_17559);
xor U17781 (N_17781,N_17458,N_17484);
nor U17782 (N_17782,N_17438,N_17449);
and U17783 (N_17783,N_17421,N_17540);
or U17784 (N_17784,N_17595,N_17586);
or U17785 (N_17785,N_17524,N_17559);
nand U17786 (N_17786,N_17464,N_17482);
and U17787 (N_17787,N_17498,N_17554);
or U17788 (N_17788,N_17443,N_17442);
or U17789 (N_17789,N_17420,N_17452);
xnor U17790 (N_17790,N_17563,N_17410);
or U17791 (N_17791,N_17512,N_17437);
nor U17792 (N_17792,N_17521,N_17419);
and U17793 (N_17793,N_17496,N_17426);
nand U17794 (N_17794,N_17528,N_17533);
nor U17795 (N_17795,N_17533,N_17598);
nand U17796 (N_17796,N_17447,N_17517);
nand U17797 (N_17797,N_17400,N_17408);
nand U17798 (N_17798,N_17516,N_17409);
xor U17799 (N_17799,N_17576,N_17529);
or U17800 (N_17800,N_17651,N_17637);
and U17801 (N_17801,N_17666,N_17609);
nand U17802 (N_17802,N_17636,N_17735);
nand U17803 (N_17803,N_17685,N_17712);
nor U17804 (N_17804,N_17639,N_17648);
or U17805 (N_17805,N_17616,N_17659);
nand U17806 (N_17806,N_17718,N_17691);
and U17807 (N_17807,N_17775,N_17771);
or U17808 (N_17808,N_17799,N_17698);
and U17809 (N_17809,N_17761,N_17758);
xor U17810 (N_17810,N_17617,N_17769);
and U17811 (N_17811,N_17791,N_17649);
nand U17812 (N_17812,N_17628,N_17716);
nand U17813 (N_17813,N_17725,N_17796);
xnor U17814 (N_17814,N_17690,N_17654);
and U17815 (N_17815,N_17773,N_17701);
nor U17816 (N_17816,N_17734,N_17715);
or U17817 (N_17817,N_17693,N_17729);
nand U17818 (N_17818,N_17658,N_17663);
or U17819 (N_17819,N_17795,N_17619);
and U17820 (N_17820,N_17696,N_17749);
nor U17821 (N_17821,N_17705,N_17724);
and U17822 (N_17822,N_17754,N_17655);
nor U17823 (N_17823,N_17731,N_17764);
xnor U17824 (N_17824,N_17687,N_17660);
nor U17825 (N_17825,N_17607,N_17717);
and U17826 (N_17826,N_17602,N_17732);
nor U17827 (N_17827,N_17667,N_17642);
and U17828 (N_17828,N_17664,N_17633);
xnor U17829 (N_17829,N_17620,N_17683);
nor U17830 (N_17830,N_17623,N_17618);
nand U17831 (N_17831,N_17782,N_17702);
nor U17832 (N_17832,N_17781,N_17680);
and U17833 (N_17833,N_17772,N_17677);
nor U17834 (N_17834,N_17656,N_17638);
nor U17835 (N_17835,N_17706,N_17747);
and U17836 (N_17836,N_17780,N_17776);
nor U17837 (N_17837,N_17610,N_17710);
nand U17838 (N_17838,N_17682,N_17721);
and U17839 (N_17839,N_17622,N_17675);
nand U17840 (N_17840,N_17614,N_17601);
nand U17841 (N_17841,N_17763,N_17703);
nand U17842 (N_17842,N_17689,N_17736);
nand U17843 (N_17843,N_17699,N_17624);
and U17844 (N_17844,N_17738,N_17668);
or U17845 (N_17845,N_17625,N_17751);
or U17846 (N_17846,N_17665,N_17788);
nand U17847 (N_17847,N_17766,N_17644);
nor U17848 (N_17848,N_17783,N_17704);
nor U17849 (N_17849,N_17730,N_17760);
xnor U17850 (N_17850,N_17708,N_17774);
xor U17851 (N_17851,N_17671,N_17645);
or U17852 (N_17852,N_17632,N_17603);
nand U17853 (N_17853,N_17640,N_17793);
nor U17854 (N_17854,N_17798,N_17700);
and U17855 (N_17855,N_17786,N_17631);
xor U17856 (N_17856,N_17646,N_17726);
nand U17857 (N_17857,N_17742,N_17684);
and U17858 (N_17858,N_17626,N_17744);
or U17859 (N_17859,N_17695,N_17741);
or U17860 (N_17860,N_17676,N_17719);
and U17861 (N_17861,N_17714,N_17688);
nor U17862 (N_17862,N_17739,N_17711);
nand U17863 (N_17863,N_17612,N_17756);
xnor U17864 (N_17864,N_17737,N_17777);
and U17865 (N_17865,N_17600,N_17604);
and U17866 (N_17866,N_17650,N_17797);
and U17867 (N_17867,N_17652,N_17755);
and U17868 (N_17868,N_17743,N_17672);
or U17869 (N_17869,N_17621,N_17681);
and U17870 (N_17870,N_17709,N_17673);
or U17871 (N_17871,N_17790,N_17794);
nor U17872 (N_17872,N_17678,N_17720);
or U17873 (N_17873,N_17767,N_17779);
or U17874 (N_17874,N_17707,N_17727);
nor U17875 (N_17875,N_17605,N_17643);
nand U17876 (N_17876,N_17635,N_17641);
nand U17877 (N_17877,N_17674,N_17757);
and U17878 (N_17878,N_17770,N_17657);
nand U17879 (N_17879,N_17740,N_17785);
nand U17880 (N_17880,N_17750,N_17765);
nor U17881 (N_17881,N_17661,N_17634);
xor U17882 (N_17882,N_17713,N_17753);
or U17883 (N_17883,N_17694,N_17647);
or U17884 (N_17884,N_17746,N_17686);
and U17885 (N_17885,N_17662,N_17611);
and U17886 (N_17886,N_17722,N_17613);
and U17887 (N_17887,N_17627,N_17692);
nand U17888 (N_17888,N_17630,N_17629);
nor U17889 (N_17889,N_17728,N_17789);
xor U17890 (N_17890,N_17733,N_17615);
and U17891 (N_17891,N_17723,N_17679);
and U17892 (N_17892,N_17606,N_17787);
xor U17893 (N_17893,N_17792,N_17768);
or U17894 (N_17894,N_17653,N_17784);
and U17895 (N_17895,N_17697,N_17762);
nand U17896 (N_17896,N_17670,N_17745);
and U17897 (N_17897,N_17759,N_17778);
and U17898 (N_17898,N_17669,N_17748);
or U17899 (N_17899,N_17608,N_17752);
nand U17900 (N_17900,N_17613,N_17696);
or U17901 (N_17901,N_17697,N_17738);
nand U17902 (N_17902,N_17681,N_17784);
or U17903 (N_17903,N_17662,N_17687);
or U17904 (N_17904,N_17713,N_17744);
nor U17905 (N_17905,N_17782,N_17673);
nor U17906 (N_17906,N_17661,N_17767);
nand U17907 (N_17907,N_17688,N_17658);
xnor U17908 (N_17908,N_17752,N_17792);
or U17909 (N_17909,N_17606,N_17669);
nor U17910 (N_17910,N_17606,N_17734);
xor U17911 (N_17911,N_17721,N_17629);
or U17912 (N_17912,N_17757,N_17675);
xnor U17913 (N_17913,N_17748,N_17612);
nand U17914 (N_17914,N_17654,N_17733);
and U17915 (N_17915,N_17702,N_17732);
or U17916 (N_17916,N_17618,N_17693);
nand U17917 (N_17917,N_17621,N_17691);
nor U17918 (N_17918,N_17787,N_17717);
xnor U17919 (N_17919,N_17728,N_17641);
nor U17920 (N_17920,N_17673,N_17755);
nor U17921 (N_17921,N_17786,N_17662);
xor U17922 (N_17922,N_17793,N_17683);
and U17923 (N_17923,N_17754,N_17625);
and U17924 (N_17924,N_17791,N_17612);
nor U17925 (N_17925,N_17798,N_17787);
xnor U17926 (N_17926,N_17624,N_17765);
and U17927 (N_17927,N_17709,N_17700);
nand U17928 (N_17928,N_17647,N_17705);
nor U17929 (N_17929,N_17628,N_17693);
xor U17930 (N_17930,N_17636,N_17757);
nand U17931 (N_17931,N_17790,N_17634);
or U17932 (N_17932,N_17709,N_17602);
nand U17933 (N_17933,N_17757,N_17788);
nand U17934 (N_17934,N_17738,N_17793);
xnor U17935 (N_17935,N_17659,N_17727);
and U17936 (N_17936,N_17657,N_17792);
xor U17937 (N_17937,N_17628,N_17733);
nand U17938 (N_17938,N_17721,N_17683);
nand U17939 (N_17939,N_17635,N_17704);
xor U17940 (N_17940,N_17665,N_17752);
or U17941 (N_17941,N_17649,N_17716);
and U17942 (N_17942,N_17735,N_17674);
or U17943 (N_17943,N_17779,N_17640);
nand U17944 (N_17944,N_17618,N_17737);
nor U17945 (N_17945,N_17659,N_17677);
xor U17946 (N_17946,N_17686,N_17724);
and U17947 (N_17947,N_17770,N_17606);
nand U17948 (N_17948,N_17734,N_17774);
nand U17949 (N_17949,N_17623,N_17703);
or U17950 (N_17950,N_17681,N_17742);
xor U17951 (N_17951,N_17772,N_17720);
nor U17952 (N_17952,N_17740,N_17646);
or U17953 (N_17953,N_17751,N_17649);
xor U17954 (N_17954,N_17627,N_17608);
xnor U17955 (N_17955,N_17681,N_17787);
xor U17956 (N_17956,N_17674,N_17782);
or U17957 (N_17957,N_17666,N_17619);
xnor U17958 (N_17958,N_17698,N_17687);
and U17959 (N_17959,N_17620,N_17722);
or U17960 (N_17960,N_17709,N_17629);
and U17961 (N_17961,N_17747,N_17637);
nand U17962 (N_17962,N_17673,N_17776);
xnor U17963 (N_17963,N_17726,N_17693);
nand U17964 (N_17964,N_17706,N_17667);
nand U17965 (N_17965,N_17780,N_17702);
nand U17966 (N_17966,N_17778,N_17751);
and U17967 (N_17967,N_17669,N_17677);
nand U17968 (N_17968,N_17665,N_17775);
nand U17969 (N_17969,N_17656,N_17652);
nand U17970 (N_17970,N_17730,N_17757);
xor U17971 (N_17971,N_17711,N_17760);
nor U17972 (N_17972,N_17768,N_17657);
and U17973 (N_17973,N_17623,N_17747);
nor U17974 (N_17974,N_17727,N_17648);
and U17975 (N_17975,N_17609,N_17758);
and U17976 (N_17976,N_17774,N_17613);
nor U17977 (N_17977,N_17621,N_17640);
nor U17978 (N_17978,N_17715,N_17718);
xnor U17979 (N_17979,N_17730,N_17652);
and U17980 (N_17980,N_17706,N_17715);
nand U17981 (N_17981,N_17697,N_17657);
and U17982 (N_17982,N_17635,N_17727);
and U17983 (N_17983,N_17615,N_17607);
nand U17984 (N_17984,N_17704,N_17700);
nor U17985 (N_17985,N_17708,N_17704);
nand U17986 (N_17986,N_17702,N_17604);
xnor U17987 (N_17987,N_17727,N_17775);
nor U17988 (N_17988,N_17705,N_17650);
and U17989 (N_17989,N_17765,N_17724);
xor U17990 (N_17990,N_17632,N_17707);
or U17991 (N_17991,N_17657,N_17667);
or U17992 (N_17992,N_17658,N_17620);
xnor U17993 (N_17993,N_17619,N_17617);
and U17994 (N_17994,N_17711,N_17702);
nand U17995 (N_17995,N_17753,N_17671);
xor U17996 (N_17996,N_17769,N_17758);
xnor U17997 (N_17997,N_17792,N_17632);
nand U17998 (N_17998,N_17797,N_17678);
nor U17999 (N_17999,N_17772,N_17743);
nor U18000 (N_18000,N_17836,N_17823);
xor U18001 (N_18001,N_17989,N_17856);
xnor U18002 (N_18002,N_17961,N_17949);
or U18003 (N_18003,N_17992,N_17822);
nand U18004 (N_18004,N_17944,N_17951);
nand U18005 (N_18005,N_17978,N_17834);
and U18006 (N_18006,N_17991,N_17930);
nand U18007 (N_18007,N_17833,N_17953);
nor U18008 (N_18008,N_17863,N_17804);
nor U18009 (N_18009,N_17920,N_17879);
xor U18010 (N_18010,N_17999,N_17966);
nand U18011 (N_18011,N_17911,N_17973);
nor U18012 (N_18012,N_17807,N_17891);
xnor U18013 (N_18013,N_17875,N_17810);
nor U18014 (N_18014,N_17809,N_17881);
and U18015 (N_18015,N_17840,N_17876);
nand U18016 (N_18016,N_17910,N_17977);
nand U18017 (N_18017,N_17902,N_17904);
xnor U18018 (N_18018,N_17865,N_17955);
or U18019 (N_18019,N_17812,N_17888);
nand U18020 (N_18020,N_17867,N_17899);
and U18021 (N_18021,N_17984,N_17996);
and U18022 (N_18022,N_17858,N_17907);
nand U18023 (N_18023,N_17974,N_17998);
nor U18024 (N_18024,N_17970,N_17898);
nand U18025 (N_18025,N_17969,N_17918);
and U18026 (N_18026,N_17962,N_17854);
or U18027 (N_18027,N_17883,N_17926);
xnor U18028 (N_18028,N_17908,N_17941);
or U18029 (N_18029,N_17895,N_17857);
nand U18030 (N_18030,N_17919,N_17968);
xor U18031 (N_18031,N_17873,N_17817);
nor U18032 (N_18032,N_17853,N_17831);
and U18033 (N_18033,N_17985,N_17972);
xor U18034 (N_18034,N_17887,N_17839);
and U18035 (N_18035,N_17936,N_17921);
and U18036 (N_18036,N_17847,N_17869);
xor U18037 (N_18037,N_17868,N_17925);
or U18038 (N_18038,N_17886,N_17923);
nand U18039 (N_18039,N_17821,N_17877);
and U18040 (N_18040,N_17960,N_17945);
or U18041 (N_18041,N_17878,N_17845);
xor U18042 (N_18042,N_17893,N_17980);
nor U18043 (N_18043,N_17874,N_17975);
nor U18044 (N_18044,N_17852,N_17880);
or U18045 (N_18045,N_17957,N_17901);
nor U18046 (N_18046,N_17849,N_17860);
xor U18047 (N_18047,N_17835,N_17859);
nand U18048 (N_18048,N_17982,N_17870);
and U18049 (N_18049,N_17929,N_17946);
nand U18050 (N_18050,N_17933,N_17844);
or U18051 (N_18051,N_17914,N_17965);
xnor U18052 (N_18052,N_17872,N_17829);
and U18053 (N_18053,N_17894,N_17912);
or U18054 (N_18054,N_17913,N_17993);
and U18055 (N_18055,N_17813,N_17900);
or U18056 (N_18056,N_17964,N_17841);
nand U18057 (N_18057,N_17842,N_17954);
or U18058 (N_18058,N_17806,N_17938);
or U18059 (N_18059,N_17937,N_17958);
xor U18060 (N_18060,N_17942,N_17802);
nor U18061 (N_18061,N_17915,N_17890);
and U18062 (N_18062,N_17861,N_17826);
and U18063 (N_18063,N_17862,N_17917);
xnor U18064 (N_18064,N_17825,N_17820);
or U18065 (N_18065,N_17882,N_17818);
nand U18066 (N_18066,N_17892,N_17801);
or U18067 (N_18067,N_17846,N_17967);
or U18068 (N_18068,N_17808,N_17885);
or U18069 (N_18069,N_17843,N_17931);
xor U18070 (N_18070,N_17924,N_17803);
and U18071 (N_18071,N_17855,N_17815);
and U18072 (N_18072,N_17995,N_17864);
xnor U18073 (N_18073,N_17922,N_17916);
nand U18074 (N_18074,N_17827,N_17959);
or U18075 (N_18075,N_17837,N_17994);
xor U18076 (N_18076,N_17934,N_17871);
and U18077 (N_18077,N_17814,N_17997);
nand U18078 (N_18078,N_17928,N_17906);
nand U18079 (N_18079,N_17987,N_17838);
nand U18080 (N_18080,N_17828,N_17830);
xor U18081 (N_18081,N_17832,N_17824);
xnor U18082 (N_18082,N_17889,N_17932);
and U18083 (N_18083,N_17811,N_17983);
and U18084 (N_18084,N_17848,N_17963);
nand U18085 (N_18085,N_17927,N_17819);
and U18086 (N_18086,N_17990,N_17981);
nor U18087 (N_18087,N_17947,N_17988);
and U18088 (N_18088,N_17979,N_17905);
xor U18089 (N_18089,N_17940,N_17896);
nor U18090 (N_18090,N_17939,N_17950);
or U18091 (N_18091,N_17884,N_17952);
nor U18092 (N_18092,N_17897,N_17816);
nor U18093 (N_18093,N_17935,N_17850);
and U18094 (N_18094,N_17976,N_17909);
nor U18095 (N_18095,N_17956,N_17943);
or U18096 (N_18096,N_17851,N_17800);
nor U18097 (N_18097,N_17866,N_17903);
nor U18098 (N_18098,N_17948,N_17971);
xor U18099 (N_18099,N_17805,N_17986);
and U18100 (N_18100,N_17847,N_17858);
nor U18101 (N_18101,N_17838,N_17986);
nand U18102 (N_18102,N_17899,N_17831);
or U18103 (N_18103,N_17954,N_17920);
and U18104 (N_18104,N_17820,N_17949);
xnor U18105 (N_18105,N_17880,N_17981);
or U18106 (N_18106,N_17991,N_17897);
or U18107 (N_18107,N_17923,N_17856);
nor U18108 (N_18108,N_17972,N_17844);
nor U18109 (N_18109,N_17899,N_17872);
xor U18110 (N_18110,N_17942,N_17993);
or U18111 (N_18111,N_17826,N_17917);
nor U18112 (N_18112,N_17828,N_17942);
nand U18113 (N_18113,N_17974,N_17905);
nand U18114 (N_18114,N_17860,N_17921);
or U18115 (N_18115,N_17968,N_17888);
xor U18116 (N_18116,N_17867,N_17890);
or U18117 (N_18117,N_17990,N_17978);
nor U18118 (N_18118,N_17928,N_17951);
nand U18119 (N_18119,N_17914,N_17917);
or U18120 (N_18120,N_17886,N_17988);
nor U18121 (N_18121,N_17877,N_17945);
or U18122 (N_18122,N_17892,N_17906);
xnor U18123 (N_18123,N_17956,N_17960);
nand U18124 (N_18124,N_17986,N_17864);
and U18125 (N_18125,N_17959,N_17898);
nor U18126 (N_18126,N_17947,N_17869);
nand U18127 (N_18127,N_17942,N_17863);
xnor U18128 (N_18128,N_17920,N_17847);
nor U18129 (N_18129,N_17860,N_17841);
nand U18130 (N_18130,N_17977,N_17876);
and U18131 (N_18131,N_17940,N_17837);
xor U18132 (N_18132,N_17863,N_17953);
xnor U18133 (N_18133,N_17934,N_17858);
nor U18134 (N_18134,N_17959,N_17923);
nor U18135 (N_18135,N_17845,N_17978);
or U18136 (N_18136,N_17854,N_17965);
xor U18137 (N_18137,N_17932,N_17861);
xnor U18138 (N_18138,N_17956,N_17930);
or U18139 (N_18139,N_17923,N_17863);
or U18140 (N_18140,N_17933,N_17806);
nand U18141 (N_18141,N_17906,N_17917);
and U18142 (N_18142,N_17850,N_17848);
nand U18143 (N_18143,N_17966,N_17856);
nand U18144 (N_18144,N_17968,N_17965);
nand U18145 (N_18145,N_17802,N_17843);
and U18146 (N_18146,N_17932,N_17906);
nor U18147 (N_18147,N_17946,N_17867);
xnor U18148 (N_18148,N_17889,N_17887);
and U18149 (N_18149,N_17991,N_17961);
or U18150 (N_18150,N_17885,N_17807);
or U18151 (N_18151,N_17814,N_17805);
xnor U18152 (N_18152,N_17878,N_17849);
and U18153 (N_18153,N_17893,N_17904);
or U18154 (N_18154,N_17830,N_17930);
or U18155 (N_18155,N_17884,N_17999);
nand U18156 (N_18156,N_17874,N_17825);
and U18157 (N_18157,N_17960,N_17978);
or U18158 (N_18158,N_17881,N_17852);
and U18159 (N_18159,N_17876,N_17885);
or U18160 (N_18160,N_17888,N_17814);
xnor U18161 (N_18161,N_17902,N_17996);
nor U18162 (N_18162,N_17964,N_17876);
or U18163 (N_18163,N_17970,N_17884);
and U18164 (N_18164,N_17993,N_17960);
or U18165 (N_18165,N_17857,N_17841);
xor U18166 (N_18166,N_17970,N_17842);
xor U18167 (N_18167,N_17811,N_17934);
and U18168 (N_18168,N_17897,N_17920);
nand U18169 (N_18169,N_17808,N_17890);
nand U18170 (N_18170,N_17836,N_17879);
or U18171 (N_18171,N_17886,N_17818);
and U18172 (N_18172,N_17915,N_17857);
or U18173 (N_18173,N_17856,N_17944);
xnor U18174 (N_18174,N_17956,N_17991);
or U18175 (N_18175,N_17907,N_17834);
xor U18176 (N_18176,N_17998,N_17824);
nor U18177 (N_18177,N_17808,N_17918);
and U18178 (N_18178,N_17853,N_17939);
nand U18179 (N_18179,N_17861,N_17997);
xor U18180 (N_18180,N_17954,N_17896);
xor U18181 (N_18181,N_17800,N_17944);
nor U18182 (N_18182,N_17897,N_17893);
or U18183 (N_18183,N_17814,N_17987);
nand U18184 (N_18184,N_17973,N_17929);
nand U18185 (N_18185,N_17806,N_17975);
nand U18186 (N_18186,N_17808,N_17889);
or U18187 (N_18187,N_17873,N_17845);
nor U18188 (N_18188,N_17927,N_17987);
or U18189 (N_18189,N_17902,N_17989);
and U18190 (N_18190,N_17859,N_17808);
or U18191 (N_18191,N_17812,N_17801);
xnor U18192 (N_18192,N_17815,N_17933);
nand U18193 (N_18193,N_17828,N_17811);
nor U18194 (N_18194,N_17939,N_17852);
nor U18195 (N_18195,N_17980,N_17922);
or U18196 (N_18196,N_17953,N_17962);
nor U18197 (N_18197,N_17853,N_17827);
nand U18198 (N_18198,N_17932,N_17846);
nand U18199 (N_18199,N_17875,N_17967);
and U18200 (N_18200,N_18000,N_18085);
or U18201 (N_18201,N_18168,N_18018);
or U18202 (N_18202,N_18147,N_18097);
nor U18203 (N_18203,N_18112,N_18101);
or U18204 (N_18204,N_18192,N_18020);
xor U18205 (N_18205,N_18056,N_18071);
or U18206 (N_18206,N_18121,N_18012);
nor U18207 (N_18207,N_18175,N_18036);
and U18208 (N_18208,N_18050,N_18140);
xor U18209 (N_18209,N_18084,N_18027);
and U18210 (N_18210,N_18125,N_18098);
nand U18211 (N_18211,N_18040,N_18086);
nor U18212 (N_18212,N_18134,N_18185);
xor U18213 (N_18213,N_18061,N_18102);
and U18214 (N_18214,N_18156,N_18001);
and U18215 (N_18215,N_18108,N_18117);
nor U18216 (N_18216,N_18015,N_18014);
nand U18217 (N_18217,N_18114,N_18022);
nand U18218 (N_18218,N_18008,N_18116);
nand U18219 (N_18219,N_18195,N_18166);
nor U18220 (N_18220,N_18094,N_18180);
or U18221 (N_18221,N_18044,N_18011);
or U18222 (N_18222,N_18127,N_18088);
xnor U18223 (N_18223,N_18129,N_18041);
or U18224 (N_18224,N_18138,N_18187);
and U18225 (N_18225,N_18106,N_18074);
nand U18226 (N_18226,N_18169,N_18188);
and U18227 (N_18227,N_18142,N_18146);
nand U18228 (N_18228,N_18190,N_18165);
nand U18229 (N_18229,N_18105,N_18184);
nand U18230 (N_18230,N_18029,N_18089);
nor U18231 (N_18231,N_18066,N_18073);
nand U18232 (N_18232,N_18103,N_18181);
nand U18233 (N_18233,N_18057,N_18064);
nand U18234 (N_18234,N_18182,N_18046);
and U18235 (N_18235,N_18058,N_18162);
nor U18236 (N_18236,N_18070,N_18055);
xor U18237 (N_18237,N_18004,N_18171);
nand U18238 (N_18238,N_18130,N_18002);
nor U18239 (N_18239,N_18150,N_18136);
nand U18240 (N_18240,N_18178,N_18090);
nor U18241 (N_18241,N_18115,N_18021);
and U18242 (N_18242,N_18191,N_18143);
nor U18243 (N_18243,N_18151,N_18049);
xnor U18244 (N_18244,N_18124,N_18081);
nor U18245 (N_18245,N_18155,N_18135);
xnor U18246 (N_18246,N_18164,N_18045);
or U18247 (N_18247,N_18170,N_18009);
or U18248 (N_18248,N_18199,N_18107);
and U18249 (N_18249,N_18119,N_18052);
xor U18250 (N_18250,N_18128,N_18054);
nand U18251 (N_18251,N_18038,N_18026);
nand U18252 (N_18252,N_18154,N_18051);
nand U18253 (N_18253,N_18031,N_18152);
nand U18254 (N_18254,N_18013,N_18059);
and U18255 (N_18255,N_18194,N_18062);
nand U18256 (N_18256,N_18024,N_18019);
nor U18257 (N_18257,N_18139,N_18030);
and U18258 (N_18258,N_18126,N_18096);
nor U18259 (N_18259,N_18072,N_18039);
nor U18260 (N_18260,N_18122,N_18197);
nor U18261 (N_18261,N_18063,N_18042);
or U18262 (N_18262,N_18033,N_18093);
and U18263 (N_18263,N_18159,N_18076);
xor U18264 (N_18264,N_18163,N_18153);
and U18265 (N_18265,N_18174,N_18035);
and U18266 (N_18266,N_18028,N_18144);
xnor U18267 (N_18267,N_18172,N_18082);
nor U18268 (N_18268,N_18083,N_18095);
xnor U18269 (N_18269,N_18186,N_18003);
nor U18270 (N_18270,N_18157,N_18141);
nor U18271 (N_18271,N_18065,N_18198);
and U18272 (N_18272,N_18167,N_18145);
xor U18273 (N_18273,N_18069,N_18079);
nor U18274 (N_18274,N_18047,N_18160);
xnor U18275 (N_18275,N_18173,N_18092);
nor U18276 (N_18276,N_18053,N_18016);
nand U18277 (N_18277,N_18023,N_18080);
and U18278 (N_18278,N_18110,N_18099);
or U18279 (N_18279,N_18091,N_18060);
and U18280 (N_18280,N_18006,N_18148);
and U18281 (N_18281,N_18100,N_18104);
xor U18282 (N_18282,N_18032,N_18078);
nor U18283 (N_18283,N_18037,N_18193);
and U18284 (N_18284,N_18067,N_18109);
xnor U18285 (N_18285,N_18133,N_18123);
nor U18286 (N_18286,N_18010,N_18005);
nand U18287 (N_18287,N_18017,N_18048);
nor U18288 (N_18288,N_18132,N_18111);
or U18289 (N_18289,N_18137,N_18177);
nand U18290 (N_18290,N_18087,N_18179);
nand U18291 (N_18291,N_18075,N_18196);
nor U18292 (N_18292,N_18113,N_18120);
xor U18293 (N_18293,N_18189,N_18183);
nand U18294 (N_18294,N_18007,N_18149);
and U18295 (N_18295,N_18176,N_18043);
and U18296 (N_18296,N_18068,N_18034);
xnor U18297 (N_18297,N_18118,N_18158);
xor U18298 (N_18298,N_18161,N_18077);
or U18299 (N_18299,N_18131,N_18025);
xor U18300 (N_18300,N_18058,N_18010);
and U18301 (N_18301,N_18082,N_18183);
nand U18302 (N_18302,N_18101,N_18119);
or U18303 (N_18303,N_18142,N_18121);
xnor U18304 (N_18304,N_18133,N_18124);
nor U18305 (N_18305,N_18104,N_18066);
and U18306 (N_18306,N_18079,N_18001);
or U18307 (N_18307,N_18038,N_18099);
xnor U18308 (N_18308,N_18117,N_18068);
and U18309 (N_18309,N_18135,N_18104);
xor U18310 (N_18310,N_18096,N_18102);
and U18311 (N_18311,N_18149,N_18053);
or U18312 (N_18312,N_18175,N_18095);
nor U18313 (N_18313,N_18127,N_18069);
or U18314 (N_18314,N_18193,N_18124);
xor U18315 (N_18315,N_18091,N_18164);
and U18316 (N_18316,N_18058,N_18047);
and U18317 (N_18317,N_18159,N_18055);
xor U18318 (N_18318,N_18000,N_18037);
nor U18319 (N_18319,N_18109,N_18139);
or U18320 (N_18320,N_18043,N_18053);
xor U18321 (N_18321,N_18006,N_18185);
and U18322 (N_18322,N_18056,N_18023);
and U18323 (N_18323,N_18180,N_18152);
xnor U18324 (N_18324,N_18100,N_18054);
nand U18325 (N_18325,N_18002,N_18057);
xor U18326 (N_18326,N_18111,N_18112);
or U18327 (N_18327,N_18178,N_18153);
xnor U18328 (N_18328,N_18027,N_18138);
and U18329 (N_18329,N_18142,N_18129);
nor U18330 (N_18330,N_18122,N_18005);
xnor U18331 (N_18331,N_18100,N_18053);
and U18332 (N_18332,N_18169,N_18092);
or U18333 (N_18333,N_18025,N_18143);
nor U18334 (N_18334,N_18050,N_18100);
or U18335 (N_18335,N_18134,N_18111);
or U18336 (N_18336,N_18030,N_18044);
nand U18337 (N_18337,N_18034,N_18078);
xnor U18338 (N_18338,N_18123,N_18196);
or U18339 (N_18339,N_18133,N_18063);
xor U18340 (N_18340,N_18037,N_18180);
xnor U18341 (N_18341,N_18018,N_18176);
and U18342 (N_18342,N_18001,N_18080);
and U18343 (N_18343,N_18047,N_18035);
and U18344 (N_18344,N_18140,N_18020);
and U18345 (N_18345,N_18017,N_18005);
and U18346 (N_18346,N_18154,N_18031);
and U18347 (N_18347,N_18110,N_18192);
xor U18348 (N_18348,N_18074,N_18098);
and U18349 (N_18349,N_18021,N_18049);
xnor U18350 (N_18350,N_18011,N_18139);
and U18351 (N_18351,N_18130,N_18016);
nand U18352 (N_18352,N_18037,N_18104);
nor U18353 (N_18353,N_18120,N_18167);
nor U18354 (N_18354,N_18017,N_18084);
nand U18355 (N_18355,N_18050,N_18017);
nand U18356 (N_18356,N_18098,N_18153);
xor U18357 (N_18357,N_18087,N_18016);
xor U18358 (N_18358,N_18132,N_18005);
and U18359 (N_18359,N_18044,N_18097);
xor U18360 (N_18360,N_18057,N_18105);
and U18361 (N_18361,N_18185,N_18184);
xor U18362 (N_18362,N_18030,N_18033);
xor U18363 (N_18363,N_18013,N_18132);
xnor U18364 (N_18364,N_18181,N_18049);
nand U18365 (N_18365,N_18166,N_18050);
and U18366 (N_18366,N_18053,N_18099);
nor U18367 (N_18367,N_18169,N_18159);
and U18368 (N_18368,N_18141,N_18129);
nor U18369 (N_18369,N_18066,N_18067);
nand U18370 (N_18370,N_18019,N_18184);
nor U18371 (N_18371,N_18157,N_18182);
xnor U18372 (N_18372,N_18193,N_18145);
and U18373 (N_18373,N_18106,N_18044);
or U18374 (N_18374,N_18111,N_18044);
xor U18375 (N_18375,N_18017,N_18076);
nor U18376 (N_18376,N_18079,N_18199);
or U18377 (N_18377,N_18051,N_18072);
xor U18378 (N_18378,N_18107,N_18144);
or U18379 (N_18379,N_18175,N_18091);
or U18380 (N_18380,N_18077,N_18096);
nand U18381 (N_18381,N_18035,N_18059);
or U18382 (N_18382,N_18022,N_18065);
nand U18383 (N_18383,N_18196,N_18132);
or U18384 (N_18384,N_18125,N_18034);
nor U18385 (N_18385,N_18117,N_18146);
nand U18386 (N_18386,N_18175,N_18172);
nor U18387 (N_18387,N_18158,N_18147);
or U18388 (N_18388,N_18119,N_18105);
or U18389 (N_18389,N_18021,N_18119);
nand U18390 (N_18390,N_18084,N_18142);
nand U18391 (N_18391,N_18001,N_18019);
or U18392 (N_18392,N_18032,N_18103);
or U18393 (N_18393,N_18187,N_18111);
nor U18394 (N_18394,N_18011,N_18188);
or U18395 (N_18395,N_18198,N_18111);
or U18396 (N_18396,N_18146,N_18175);
or U18397 (N_18397,N_18104,N_18060);
and U18398 (N_18398,N_18179,N_18057);
xor U18399 (N_18399,N_18100,N_18067);
nand U18400 (N_18400,N_18220,N_18251);
nor U18401 (N_18401,N_18200,N_18386);
xor U18402 (N_18402,N_18261,N_18375);
nor U18403 (N_18403,N_18284,N_18316);
nand U18404 (N_18404,N_18358,N_18339);
or U18405 (N_18405,N_18393,N_18288);
and U18406 (N_18406,N_18275,N_18348);
nand U18407 (N_18407,N_18268,N_18292);
nor U18408 (N_18408,N_18346,N_18303);
and U18409 (N_18409,N_18307,N_18293);
xnor U18410 (N_18410,N_18267,N_18235);
nand U18411 (N_18411,N_18330,N_18334);
nand U18412 (N_18412,N_18229,N_18382);
and U18413 (N_18413,N_18387,N_18398);
nand U18414 (N_18414,N_18390,N_18364);
or U18415 (N_18415,N_18389,N_18244);
nand U18416 (N_18416,N_18299,N_18266);
xor U18417 (N_18417,N_18372,N_18278);
nor U18418 (N_18418,N_18373,N_18304);
and U18419 (N_18419,N_18357,N_18306);
nor U18420 (N_18420,N_18343,N_18240);
nand U18421 (N_18421,N_18344,N_18248);
or U18422 (N_18422,N_18279,N_18350);
xnor U18423 (N_18423,N_18301,N_18361);
nor U18424 (N_18424,N_18219,N_18383);
xor U18425 (N_18425,N_18399,N_18381);
xnor U18426 (N_18426,N_18236,N_18388);
xnor U18427 (N_18427,N_18242,N_18216);
nor U18428 (N_18428,N_18222,N_18298);
xnor U18429 (N_18429,N_18239,N_18221);
or U18430 (N_18430,N_18243,N_18341);
and U18431 (N_18431,N_18327,N_18258);
nor U18432 (N_18432,N_18379,N_18207);
xor U18433 (N_18433,N_18213,N_18203);
or U18434 (N_18434,N_18300,N_18217);
xnor U18435 (N_18435,N_18319,N_18255);
nand U18436 (N_18436,N_18362,N_18246);
nand U18437 (N_18437,N_18332,N_18384);
xnor U18438 (N_18438,N_18295,N_18276);
nor U18439 (N_18439,N_18366,N_18228);
or U18440 (N_18440,N_18356,N_18272);
xor U18441 (N_18441,N_18367,N_18215);
and U18442 (N_18442,N_18237,N_18297);
nand U18443 (N_18443,N_18359,N_18337);
nor U18444 (N_18444,N_18308,N_18397);
nand U18445 (N_18445,N_18290,N_18391);
nor U18446 (N_18446,N_18321,N_18206);
xor U18447 (N_18447,N_18286,N_18269);
or U18448 (N_18448,N_18260,N_18225);
xor U18449 (N_18449,N_18287,N_18296);
nor U18450 (N_18450,N_18318,N_18281);
xnor U18451 (N_18451,N_18324,N_18325);
and U18452 (N_18452,N_18340,N_18342);
nor U18453 (N_18453,N_18309,N_18257);
nor U18454 (N_18454,N_18352,N_18310);
or U18455 (N_18455,N_18265,N_18283);
and U18456 (N_18456,N_18355,N_18320);
and U18457 (N_18457,N_18205,N_18253);
nand U18458 (N_18458,N_18333,N_18368);
nor U18459 (N_18459,N_18227,N_18302);
nand U18460 (N_18460,N_18263,N_18365);
and U18461 (N_18461,N_18395,N_18289);
nand U18462 (N_18462,N_18204,N_18282);
nand U18463 (N_18463,N_18347,N_18226);
nand U18464 (N_18464,N_18285,N_18241);
xnor U18465 (N_18465,N_18234,N_18315);
nand U18466 (N_18466,N_18233,N_18210);
or U18467 (N_18467,N_18280,N_18311);
nor U18468 (N_18468,N_18392,N_18378);
or U18469 (N_18469,N_18294,N_18328);
nand U18470 (N_18470,N_18247,N_18312);
or U18471 (N_18471,N_18376,N_18323);
and U18472 (N_18472,N_18259,N_18252);
xor U18473 (N_18473,N_18370,N_18394);
nor U18474 (N_18474,N_18224,N_18369);
nand U18475 (N_18475,N_18250,N_18322);
or U18476 (N_18476,N_18231,N_18273);
nor U18477 (N_18477,N_18291,N_18238);
nand U18478 (N_18478,N_18305,N_18201);
nor U18479 (N_18479,N_18274,N_18218);
and U18480 (N_18480,N_18214,N_18249);
and U18481 (N_18481,N_18254,N_18329);
nor U18482 (N_18482,N_18360,N_18377);
and U18483 (N_18483,N_18232,N_18336);
xnor U18484 (N_18484,N_18230,N_18211);
or U18485 (N_18485,N_18345,N_18374);
xnor U18486 (N_18486,N_18313,N_18245);
xnor U18487 (N_18487,N_18317,N_18208);
nor U18488 (N_18488,N_18371,N_18338);
xnor U18489 (N_18489,N_18209,N_18385);
xnor U18490 (N_18490,N_18396,N_18264);
nor U18491 (N_18491,N_18223,N_18380);
or U18492 (N_18492,N_18351,N_18212);
nor U18493 (N_18493,N_18335,N_18277);
or U18494 (N_18494,N_18363,N_18262);
nand U18495 (N_18495,N_18326,N_18353);
nor U18496 (N_18496,N_18314,N_18331);
and U18497 (N_18497,N_18256,N_18354);
nand U18498 (N_18498,N_18271,N_18349);
nor U18499 (N_18499,N_18202,N_18270);
or U18500 (N_18500,N_18213,N_18319);
xnor U18501 (N_18501,N_18366,N_18343);
and U18502 (N_18502,N_18348,N_18223);
nor U18503 (N_18503,N_18323,N_18245);
nor U18504 (N_18504,N_18230,N_18256);
and U18505 (N_18505,N_18332,N_18278);
nand U18506 (N_18506,N_18266,N_18355);
or U18507 (N_18507,N_18284,N_18204);
nor U18508 (N_18508,N_18293,N_18390);
nor U18509 (N_18509,N_18241,N_18226);
nand U18510 (N_18510,N_18315,N_18336);
nand U18511 (N_18511,N_18204,N_18248);
and U18512 (N_18512,N_18280,N_18266);
nor U18513 (N_18513,N_18261,N_18240);
nor U18514 (N_18514,N_18312,N_18342);
nand U18515 (N_18515,N_18376,N_18395);
xnor U18516 (N_18516,N_18252,N_18360);
nor U18517 (N_18517,N_18355,N_18328);
nor U18518 (N_18518,N_18239,N_18295);
and U18519 (N_18519,N_18317,N_18351);
xor U18520 (N_18520,N_18245,N_18339);
xor U18521 (N_18521,N_18279,N_18245);
nor U18522 (N_18522,N_18219,N_18213);
xnor U18523 (N_18523,N_18269,N_18355);
and U18524 (N_18524,N_18279,N_18356);
and U18525 (N_18525,N_18284,N_18261);
xnor U18526 (N_18526,N_18353,N_18200);
nor U18527 (N_18527,N_18326,N_18384);
nor U18528 (N_18528,N_18373,N_18305);
and U18529 (N_18529,N_18358,N_18224);
nand U18530 (N_18530,N_18200,N_18366);
xnor U18531 (N_18531,N_18240,N_18243);
nand U18532 (N_18532,N_18338,N_18240);
xnor U18533 (N_18533,N_18250,N_18260);
nand U18534 (N_18534,N_18330,N_18343);
and U18535 (N_18535,N_18378,N_18282);
xor U18536 (N_18536,N_18248,N_18363);
xnor U18537 (N_18537,N_18315,N_18389);
xor U18538 (N_18538,N_18309,N_18208);
xnor U18539 (N_18539,N_18347,N_18286);
or U18540 (N_18540,N_18276,N_18307);
nand U18541 (N_18541,N_18268,N_18365);
and U18542 (N_18542,N_18255,N_18252);
nand U18543 (N_18543,N_18391,N_18355);
or U18544 (N_18544,N_18326,N_18210);
xnor U18545 (N_18545,N_18340,N_18274);
xor U18546 (N_18546,N_18390,N_18288);
or U18547 (N_18547,N_18225,N_18256);
nand U18548 (N_18548,N_18242,N_18280);
nor U18549 (N_18549,N_18384,N_18287);
xnor U18550 (N_18550,N_18223,N_18228);
and U18551 (N_18551,N_18371,N_18318);
xor U18552 (N_18552,N_18372,N_18279);
nand U18553 (N_18553,N_18254,N_18206);
nor U18554 (N_18554,N_18267,N_18218);
and U18555 (N_18555,N_18348,N_18387);
nand U18556 (N_18556,N_18237,N_18274);
or U18557 (N_18557,N_18202,N_18219);
or U18558 (N_18558,N_18301,N_18310);
nand U18559 (N_18559,N_18341,N_18212);
and U18560 (N_18560,N_18229,N_18341);
xnor U18561 (N_18561,N_18333,N_18331);
or U18562 (N_18562,N_18208,N_18257);
or U18563 (N_18563,N_18303,N_18290);
xnor U18564 (N_18564,N_18388,N_18381);
nand U18565 (N_18565,N_18250,N_18320);
nor U18566 (N_18566,N_18350,N_18287);
or U18567 (N_18567,N_18376,N_18260);
nand U18568 (N_18568,N_18380,N_18212);
and U18569 (N_18569,N_18313,N_18272);
and U18570 (N_18570,N_18214,N_18206);
nand U18571 (N_18571,N_18222,N_18218);
xnor U18572 (N_18572,N_18251,N_18201);
xor U18573 (N_18573,N_18285,N_18253);
nand U18574 (N_18574,N_18398,N_18336);
nor U18575 (N_18575,N_18221,N_18373);
or U18576 (N_18576,N_18269,N_18291);
or U18577 (N_18577,N_18247,N_18250);
or U18578 (N_18578,N_18201,N_18291);
nor U18579 (N_18579,N_18379,N_18247);
nand U18580 (N_18580,N_18254,N_18229);
nand U18581 (N_18581,N_18353,N_18231);
xnor U18582 (N_18582,N_18286,N_18365);
nor U18583 (N_18583,N_18273,N_18397);
nand U18584 (N_18584,N_18204,N_18398);
or U18585 (N_18585,N_18285,N_18209);
and U18586 (N_18586,N_18394,N_18227);
and U18587 (N_18587,N_18333,N_18326);
nand U18588 (N_18588,N_18247,N_18324);
nand U18589 (N_18589,N_18380,N_18202);
nor U18590 (N_18590,N_18271,N_18353);
xor U18591 (N_18591,N_18378,N_18308);
or U18592 (N_18592,N_18371,N_18246);
nand U18593 (N_18593,N_18239,N_18348);
nand U18594 (N_18594,N_18282,N_18348);
nand U18595 (N_18595,N_18332,N_18299);
or U18596 (N_18596,N_18378,N_18344);
nor U18597 (N_18597,N_18257,N_18363);
and U18598 (N_18598,N_18216,N_18398);
and U18599 (N_18599,N_18255,N_18361);
nand U18600 (N_18600,N_18533,N_18418);
nor U18601 (N_18601,N_18413,N_18446);
xor U18602 (N_18602,N_18549,N_18469);
nand U18603 (N_18603,N_18504,N_18441);
xor U18604 (N_18604,N_18415,N_18589);
or U18605 (N_18605,N_18405,N_18482);
nand U18606 (N_18606,N_18567,N_18524);
or U18607 (N_18607,N_18519,N_18512);
nor U18608 (N_18608,N_18464,N_18546);
and U18609 (N_18609,N_18596,N_18428);
or U18610 (N_18610,N_18516,N_18445);
and U18611 (N_18611,N_18494,N_18444);
nor U18612 (N_18612,N_18500,N_18556);
or U18613 (N_18613,N_18401,N_18518);
or U18614 (N_18614,N_18417,N_18575);
nand U18615 (N_18615,N_18410,N_18552);
xor U18616 (N_18616,N_18560,N_18566);
nand U18617 (N_18617,N_18424,N_18574);
nor U18618 (N_18618,N_18577,N_18407);
nand U18619 (N_18619,N_18585,N_18453);
and U18620 (N_18620,N_18576,N_18511);
nand U18621 (N_18621,N_18471,N_18578);
or U18622 (N_18622,N_18543,N_18558);
and U18623 (N_18623,N_18528,N_18565);
and U18624 (N_18624,N_18535,N_18579);
or U18625 (N_18625,N_18509,N_18573);
and U18626 (N_18626,N_18544,N_18443);
nand U18627 (N_18627,N_18473,N_18406);
and U18628 (N_18628,N_18484,N_18536);
or U18629 (N_18629,N_18427,N_18548);
or U18630 (N_18630,N_18540,N_18476);
nand U18631 (N_18631,N_18423,N_18409);
and U18632 (N_18632,N_18495,N_18571);
or U18633 (N_18633,N_18483,N_18437);
nand U18634 (N_18634,N_18547,N_18563);
nand U18635 (N_18635,N_18463,N_18442);
and U18636 (N_18636,N_18582,N_18523);
xor U18637 (N_18637,N_18590,N_18431);
or U18638 (N_18638,N_18595,N_18538);
and U18639 (N_18639,N_18522,N_18513);
nor U18640 (N_18640,N_18599,N_18485);
nand U18641 (N_18641,N_18532,N_18489);
or U18642 (N_18642,N_18474,N_18490);
or U18643 (N_18643,N_18587,N_18527);
nand U18644 (N_18644,N_18435,N_18457);
nand U18645 (N_18645,N_18488,N_18531);
xnor U18646 (N_18646,N_18467,N_18480);
or U18647 (N_18647,N_18411,N_18597);
xnor U18648 (N_18648,N_18404,N_18561);
and U18649 (N_18649,N_18551,N_18506);
nor U18650 (N_18650,N_18429,N_18412);
nand U18651 (N_18651,N_18588,N_18439);
nand U18652 (N_18652,N_18541,N_18502);
and U18653 (N_18653,N_18434,N_18419);
nand U18654 (N_18654,N_18496,N_18452);
nand U18655 (N_18655,N_18529,N_18477);
or U18656 (N_18656,N_18553,N_18537);
nor U18657 (N_18657,N_18472,N_18598);
or U18658 (N_18658,N_18498,N_18534);
or U18659 (N_18659,N_18525,N_18581);
or U18660 (N_18660,N_18583,N_18436);
and U18661 (N_18661,N_18479,N_18440);
and U18662 (N_18662,N_18569,N_18550);
and U18663 (N_18663,N_18449,N_18475);
and U18664 (N_18664,N_18478,N_18491);
or U18665 (N_18665,N_18572,N_18564);
nand U18666 (N_18666,N_18508,N_18584);
nor U18667 (N_18667,N_18425,N_18466);
and U18668 (N_18668,N_18492,N_18433);
xnor U18669 (N_18669,N_18454,N_18594);
nor U18670 (N_18670,N_18420,N_18517);
xnor U18671 (N_18671,N_18493,N_18507);
xnor U18672 (N_18672,N_18545,N_18487);
xnor U18673 (N_18673,N_18530,N_18421);
or U18674 (N_18674,N_18539,N_18592);
xnor U18675 (N_18675,N_18562,N_18447);
nand U18676 (N_18676,N_18461,N_18400);
or U18677 (N_18677,N_18497,N_18542);
nand U18678 (N_18678,N_18591,N_18505);
nor U18679 (N_18679,N_18468,N_18510);
xor U18680 (N_18680,N_18459,N_18514);
xor U18681 (N_18681,N_18521,N_18450);
nor U18682 (N_18682,N_18462,N_18458);
xnor U18683 (N_18683,N_18460,N_18580);
or U18684 (N_18684,N_18430,N_18554);
nor U18685 (N_18685,N_18568,N_18455);
nand U18686 (N_18686,N_18526,N_18470);
nor U18687 (N_18687,N_18456,N_18499);
nand U18688 (N_18688,N_18486,N_18503);
xor U18689 (N_18689,N_18432,N_18422);
and U18690 (N_18690,N_18403,N_18448);
or U18691 (N_18691,N_18555,N_18414);
nor U18692 (N_18692,N_18481,N_18402);
nand U18693 (N_18693,N_18438,N_18426);
or U18694 (N_18694,N_18520,N_18557);
xor U18695 (N_18695,N_18593,N_18451);
and U18696 (N_18696,N_18408,N_18465);
nand U18697 (N_18697,N_18501,N_18586);
xnor U18698 (N_18698,N_18570,N_18559);
nor U18699 (N_18699,N_18416,N_18515);
nor U18700 (N_18700,N_18595,N_18491);
or U18701 (N_18701,N_18568,N_18566);
xnor U18702 (N_18702,N_18596,N_18504);
xnor U18703 (N_18703,N_18470,N_18506);
nor U18704 (N_18704,N_18550,N_18537);
nor U18705 (N_18705,N_18513,N_18599);
or U18706 (N_18706,N_18439,N_18495);
nand U18707 (N_18707,N_18437,N_18553);
xor U18708 (N_18708,N_18536,N_18533);
xor U18709 (N_18709,N_18556,N_18512);
and U18710 (N_18710,N_18570,N_18517);
nand U18711 (N_18711,N_18585,N_18450);
nor U18712 (N_18712,N_18595,N_18439);
xnor U18713 (N_18713,N_18484,N_18546);
nand U18714 (N_18714,N_18555,N_18519);
or U18715 (N_18715,N_18458,N_18575);
and U18716 (N_18716,N_18584,N_18497);
nor U18717 (N_18717,N_18439,N_18475);
nand U18718 (N_18718,N_18433,N_18400);
xnor U18719 (N_18719,N_18449,N_18466);
nand U18720 (N_18720,N_18505,N_18483);
xnor U18721 (N_18721,N_18479,N_18569);
or U18722 (N_18722,N_18468,N_18408);
or U18723 (N_18723,N_18485,N_18401);
or U18724 (N_18724,N_18510,N_18473);
or U18725 (N_18725,N_18522,N_18449);
or U18726 (N_18726,N_18475,N_18534);
and U18727 (N_18727,N_18444,N_18523);
nand U18728 (N_18728,N_18536,N_18436);
xnor U18729 (N_18729,N_18592,N_18521);
nand U18730 (N_18730,N_18473,N_18491);
and U18731 (N_18731,N_18442,N_18546);
xor U18732 (N_18732,N_18550,N_18529);
nor U18733 (N_18733,N_18427,N_18445);
nor U18734 (N_18734,N_18592,N_18517);
nor U18735 (N_18735,N_18407,N_18500);
nand U18736 (N_18736,N_18578,N_18474);
nand U18737 (N_18737,N_18526,N_18518);
nor U18738 (N_18738,N_18597,N_18430);
xnor U18739 (N_18739,N_18543,N_18418);
or U18740 (N_18740,N_18425,N_18405);
or U18741 (N_18741,N_18427,N_18574);
xnor U18742 (N_18742,N_18442,N_18585);
nor U18743 (N_18743,N_18560,N_18569);
nor U18744 (N_18744,N_18499,N_18579);
xor U18745 (N_18745,N_18494,N_18513);
nand U18746 (N_18746,N_18414,N_18561);
and U18747 (N_18747,N_18532,N_18577);
and U18748 (N_18748,N_18458,N_18523);
or U18749 (N_18749,N_18505,N_18419);
nand U18750 (N_18750,N_18558,N_18468);
nand U18751 (N_18751,N_18404,N_18528);
or U18752 (N_18752,N_18591,N_18451);
or U18753 (N_18753,N_18597,N_18433);
or U18754 (N_18754,N_18551,N_18410);
or U18755 (N_18755,N_18406,N_18530);
nand U18756 (N_18756,N_18574,N_18484);
xor U18757 (N_18757,N_18553,N_18597);
xnor U18758 (N_18758,N_18469,N_18553);
and U18759 (N_18759,N_18516,N_18469);
nand U18760 (N_18760,N_18530,N_18523);
nand U18761 (N_18761,N_18517,N_18549);
xor U18762 (N_18762,N_18492,N_18560);
nand U18763 (N_18763,N_18551,N_18404);
nor U18764 (N_18764,N_18429,N_18538);
nand U18765 (N_18765,N_18465,N_18585);
nor U18766 (N_18766,N_18553,N_18434);
nor U18767 (N_18767,N_18439,N_18582);
nand U18768 (N_18768,N_18560,N_18495);
nor U18769 (N_18769,N_18519,N_18533);
nand U18770 (N_18770,N_18466,N_18516);
nor U18771 (N_18771,N_18489,N_18460);
and U18772 (N_18772,N_18463,N_18512);
nor U18773 (N_18773,N_18449,N_18477);
and U18774 (N_18774,N_18414,N_18460);
nor U18775 (N_18775,N_18552,N_18534);
xor U18776 (N_18776,N_18474,N_18471);
nand U18777 (N_18777,N_18591,N_18458);
nand U18778 (N_18778,N_18599,N_18528);
nor U18779 (N_18779,N_18490,N_18559);
xnor U18780 (N_18780,N_18587,N_18499);
nor U18781 (N_18781,N_18591,N_18542);
nand U18782 (N_18782,N_18589,N_18455);
or U18783 (N_18783,N_18533,N_18495);
nand U18784 (N_18784,N_18560,N_18465);
nor U18785 (N_18785,N_18469,N_18594);
nor U18786 (N_18786,N_18401,N_18443);
nand U18787 (N_18787,N_18597,N_18464);
or U18788 (N_18788,N_18545,N_18562);
nor U18789 (N_18789,N_18579,N_18575);
nor U18790 (N_18790,N_18591,N_18520);
nor U18791 (N_18791,N_18434,N_18411);
and U18792 (N_18792,N_18436,N_18442);
xor U18793 (N_18793,N_18415,N_18528);
xnor U18794 (N_18794,N_18402,N_18520);
and U18795 (N_18795,N_18459,N_18572);
nand U18796 (N_18796,N_18545,N_18577);
nor U18797 (N_18797,N_18577,N_18590);
or U18798 (N_18798,N_18555,N_18597);
xnor U18799 (N_18799,N_18442,N_18479);
or U18800 (N_18800,N_18731,N_18647);
nand U18801 (N_18801,N_18630,N_18669);
nand U18802 (N_18802,N_18651,N_18737);
xnor U18803 (N_18803,N_18629,N_18762);
nand U18804 (N_18804,N_18634,N_18710);
and U18805 (N_18805,N_18705,N_18702);
or U18806 (N_18806,N_18645,N_18641);
nor U18807 (N_18807,N_18712,N_18604);
nor U18808 (N_18808,N_18750,N_18779);
or U18809 (N_18809,N_18755,N_18660);
or U18810 (N_18810,N_18619,N_18766);
and U18811 (N_18811,N_18740,N_18663);
nand U18812 (N_18812,N_18717,N_18721);
or U18813 (N_18813,N_18610,N_18690);
or U18814 (N_18814,N_18677,N_18681);
xnor U18815 (N_18815,N_18603,N_18780);
or U18816 (N_18816,N_18646,N_18682);
nand U18817 (N_18817,N_18614,N_18632);
nand U18818 (N_18818,N_18738,N_18767);
and U18819 (N_18819,N_18623,N_18709);
or U18820 (N_18820,N_18640,N_18667);
xor U18821 (N_18821,N_18622,N_18714);
or U18822 (N_18822,N_18633,N_18616);
xnor U18823 (N_18823,N_18782,N_18786);
nor U18824 (N_18824,N_18668,N_18763);
and U18825 (N_18825,N_18795,N_18676);
and U18826 (N_18826,N_18765,N_18708);
and U18827 (N_18827,N_18788,N_18725);
xor U18828 (N_18828,N_18678,N_18688);
nor U18829 (N_18829,N_18699,N_18711);
nor U18830 (N_18830,N_18716,N_18670);
xor U18831 (N_18831,N_18635,N_18696);
or U18832 (N_18832,N_18754,N_18791);
xor U18833 (N_18833,N_18602,N_18661);
or U18834 (N_18834,N_18726,N_18697);
or U18835 (N_18835,N_18664,N_18722);
xnor U18836 (N_18836,N_18793,N_18608);
xor U18837 (N_18837,N_18680,N_18774);
xnor U18838 (N_18838,N_18691,N_18797);
and U18839 (N_18839,N_18659,N_18666);
and U18840 (N_18840,N_18729,N_18761);
nor U18841 (N_18841,N_18615,N_18747);
and U18842 (N_18842,N_18784,N_18776);
xor U18843 (N_18843,N_18799,N_18768);
nor U18844 (N_18844,N_18777,N_18673);
nand U18845 (N_18845,N_18639,N_18636);
xor U18846 (N_18846,N_18662,N_18798);
nand U18847 (N_18847,N_18706,N_18787);
nor U18848 (N_18848,N_18649,N_18644);
nor U18849 (N_18849,N_18744,N_18684);
nand U18850 (N_18850,N_18718,N_18772);
nor U18851 (N_18851,N_18600,N_18758);
nand U18852 (N_18852,N_18781,N_18730);
nor U18853 (N_18853,N_18685,N_18759);
nand U18854 (N_18854,N_18692,N_18693);
nor U18855 (N_18855,N_18679,N_18741);
nor U18856 (N_18856,N_18720,N_18665);
xnor U18857 (N_18857,N_18689,N_18612);
nand U18858 (N_18858,N_18631,N_18783);
nand U18859 (N_18859,N_18732,N_18655);
or U18860 (N_18860,N_18743,N_18753);
xnor U18861 (N_18861,N_18642,N_18728);
and U18862 (N_18862,N_18727,N_18626);
nand U18863 (N_18863,N_18792,N_18757);
xor U18864 (N_18864,N_18736,N_18724);
or U18865 (N_18865,N_18742,N_18707);
xor U18866 (N_18866,N_18658,N_18746);
nand U18867 (N_18867,N_18609,N_18628);
nor U18868 (N_18868,N_18789,N_18613);
or U18869 (N_18869,N_18625,N_18713);
xnor U18870 (N_18870,N_18771,N_18701);
xnor U18871 (N_18871,N_18764,N_18627);
nor U18872 (N_18872,N_18611,N_18773);
or U18873 (N_18873,N_18617,N_18739);
xnor U18874 (N_18874,N_18671,N_18653);
xor U18875 (N_18875,N_18686,N_18675);
and U18876 (N_18876,N_18785,N_18745);
nand U18877 (N_18877,N_18621,N_18674);
xnor U18878 (N_18878,N_18624,N_18698);
and U18879 (N_18879,N_18719,N_18643);
or U18880 (N_18880,N_18620,N_18683);
and U18881 (N_18881,N_18601,N_18700);
and U18882 (N_18882,N_18652,N_18607);
or U18883 (N_18883,N_18715,N_18734);
nand U18884 (N_18884,N_18748,N_18648);
xor U18885 (N_18885,N_18638,N_18794);
xor U18886 (N_18886,N_18775,N_18796);
xor U18887 (N_18887,N_18637,N_18695);
xnor U18888 (N_18888,N_18769,N_18618);
nor U18889 (N_18889,N_18656,N_18723);
or U18890 (N_18890,N_18672,N_18687);
or U18891 (N_18891,N_18749,N_18733);
or U18892 (N_18892,N_18657,N_18778);
nor U18893 (N_18893,N_18650,N_18694);
nand U18894 (N_18894,N_18606,N_18790);
xnor U18895 (N_18895,N_18704,N_18703);
or U18896 (N_18896,N_18735,N_18760);
and U18897 (N_18897,N_18654,N_18770);
nor U18898 (N_18898,N_18752,N_18751);
and U18899 (N_18899,N_18756,N_18605);
nand U18900 (N_18900,N_18762,N_18759);
or U18901 (N_18901,N_18719,N_18689);
or U18902 (N_18902,N_18630,N_18670);
or U18903 (N_18903,N_18657,N_18787);
xor U18904 (N_18904,N_18659,N_18611);
nor U18905 (N_18905,N_18632,N_18766);
or U18906 (N_18906,N_18779,N_18718);
nand U18907 (N_18907,N_18699,N_18702);
and U18908 (N_18908,N_18674,N_18753);
and U18909 (N_18909,N_18646,N_18681);
nand U18910 (N_18910,N_18698,N_18658);
and U18911 (N_18911,N_18648,N_18684);
nor U18912 (N_18912,N_18771,N_18678);
nand U18913 (N_18913,N_18687,N_18769);
and U18914 (N_18914,N_18649,N_18622);
or U18915 (N_18915,N_18769,N_18619);
xor U18916 (N_18916,N_18646,N_18736);
xor U18917 (N_18917,N_18629,N_18690);
and U18918 (N_18918,N_18694,N_18652);
or U18919 (N_18919,N_18730,N_18633);
and U18920 (N_18920,N_18600,N_18742);
or U18921 (N_18921,N_18671,N_18642);
nor U18922 (N_18922,N_18772,N_18762);
and U18923 (N_18923,N_18601,N_18791);
nand U18924 (N_18924,N_18651,N_18741);
xnor U18925 (N_18925,N_18603,N_18758);
and U18926 (N_18926,N_18680,N_18741);
nand U18927 (N_18927,N_18781,N_18636);
or U18928 (N_18928,N_18669,N_18625);
xor U18929 (N_18929,N_18715,N_18620);
or U18930 (N_18930,N_18701,N_18676);
and U18931 (N_18931,N_18657,N_18683);
nand U18932 (N_18932,N_18734,N_18615);
nor U18933 (N_18933,N_18717,N_18754);
xor U18934 (N_18934,N_18759,N_18605);
or U18935 (N_18935,N_18653,N_18739);
and U18936 (N_18936,N_18746,N_18756);
and U18937 (N_18937,N_18643,N_18738);
or U18938 (N_18938,N_18600,N_18608);
nor U18939 (N_18939,N_18755,N_18763);
xor U18940 (N_18940,N_18780,N_18724);
nor U18941 (N_18941,N_18735,N_18632);
nand U18942 (N_18942,N_18764,N_18728);
xnor U18943 (N_18943,N_18639,N_18760);
or U18944 (N_18944,N_18796,N_18658);
nor U18945 (N_18945,N_18752,N_18641);
xnor U18946 (N_18946,N_18719,N_18635);
or U18947 (N_18947,N_18674,N_18622);
and U18948 (N_18948,N_18705,N_18627);
nor U18949 (N_18949,N_18780,N_18799);
xor U18950 (N_18950,N_18772,N_18780);
xnor U18951 (N_18951,N_18755,N_18613);
xnor U18952 (N_18952,N_18764,N_18762);
nor U18953 (N_18953,N_18636,N_18766);
nor U18954 (N_18954,N_18765,N_18717);
or U18955 (N_18955,N_18737,N_18749);
nor U18956 (N_18956,N_18670,N_18679);
or U18957 (N_18957,N_18673,N_18761);
xnor U18958 (N_18958,N_18775,N_18773);
nand U18959 (N_18959,N_18786,N_18791);
or U18960 (N_18960,N_18635,N_18602);
or U18961 (N_18961,N_18702,N_18610);
and U18962 (N_18962,N_18619,N_18716);
and U18963 (N_18963,N_18637,N_18765);
nor U18964 (N_18964,N_18768,N_18724);
xnor U18965 (N_18965,N_18741,N_18772);
nor U18966 (N_18966,N_18637,N_18716);
and U18967 (N_18967,N_18677,N_18685);
and U18968 (N_18968,N_18677,N_18741);
xor U18969 (N_18969,N_18603,N_18785);
nand U18970 (N_18970,N_18684,N_18745);
and U18971 (N_18971,N_18632,N_18654);
or U18972 (N_18972,N_18603,N_18645);
or U18973 (N_18973,N_18706,N_18618);
xor U18974 (N_18974,N_18704,N_18775);
xor U18975 (N_18975,N_18680,N_18751);
nor U18976 (N_18976,N_18681,N_18628);
or U18977 (N_18977,N_18656,N_18644);
and U18978 (N_18978,N_18786,N_18637);
nor U18979 (N_18979,N_18629,N_18662);
or U18980 (N_18980,N_18754,N_18600);
or U18981 (N_18981,N_18748,N_18766);
xor U18982 (N_18982,N_18639,N_18622);
nor U18983 (N_18983,N_18749,N_18663);
and U18984 (N_18984,N_18799,N_18643);
or U18985 (N_18985,N_18683,N_18696);
or U18986 (N_18986,N_18711,N_18782);
or U18987 (N_18987,N_18627,N_18735);
nor U18988 (N_18988,N_18668,N_18657);
and U18989 (N_18989,N_18732,N_18636);
nor U18990 (N_18990,N_18794,N_18690);
nand U18991 (N_18991,N_18731,N_18772);
and U18992 (N_18992,N_18619,N_18652);
and U18993 (N_18993,N_18768,N_18642);
xor U18994 (N_18994,N_18659,N_18722);
or U18995 (N_18995,N_18718,N_18656);
nor U18996 (N_18996,N_18649,N_18795);
nor U18997 (N_18997,N_18621,N_18786);
nand U18998 (N_18998,N_18683,N_18734);
or U18999 (N_18999,N_18630,N_18757);
xnor U19000 (N_19000,N_18917,N_18975);
xor U19001 (N_19001,N_18951,N_18990);
nand U19002 (N_19002,N_18882,N_18803);
or U19003 (N_19003,N_18855,N_18937);
xor U19004 (N_19004,N_18897,N_18867);
xnor U19005 (N_19005,N_18864,N_18842);
or U19006 (N_19006,N_18869,N_18874);
or U19007 (N_19007,N_18868,N_18865);
xnor U19008 (N_19008,N_18941,N_18978);
xnor U19009 (N_19009,N_18844,N_18888);
nand U19010 (N_19010,N_18817,N_18801);
nor U19011 (N_19011,N_18822,N_18945);
xor U19012 (N_19012,N_18965,N_18830);
xnor U19013 (N_19013,N_18833,N_18805);
or U19014 (N_19014,N_18906,N_18922);
xnor U19015 (N_19015,N_18918,N_18889);
nor U19016 (N_19016,N_18826,N_18960);
nor U19017 (N_19017,N_18985,N_18993);
and U19018 (N_19018,N_18849,N_18954);
or U19019 (N_19019,N_18992,N_18900);
nor U19020 (N_19020,N_18902,N_18995);
or U19021 (N_19021,N_18914,N_18967);
and U19022 (N_19022,N_18972,N_18934);
or U19023 (N_19023,N_18832,N_18932);
nor U19024 (N_19024,N_18870,N_18921);
xor U19025 (N_19025,N_18959,N_18892);
xnor U19026 (N_19026,N_18950,N_18858);
xor U19027 (N_19027,N_18880,N_18829);
and U19028 (N_19028,N_18938,N_18852);
xnor U19029 (N_19029,N_18894,N_18881);
nand U19030 (N_19030,N_18983,N_18839);
and U19031 (N_19031,N_18991,N_18891);
nor U19032 (N_19032,N_18814,N_18856);
nand U19033 (N_19033,N_18903,N_18929);
nand U19034 (N_19034,N_18928,N_18925);
nand U19035 (N_19035,N_18943,N_18847);
or U19036 (N_19036,N_18893,N_18963);
nand U19037 (N_19037,N_18875,N_18936);
or U19038 (N_19038,N_18848,N_18804);
and U19039 (N_19039,N_18911,N_18896);
and U19040 (N_19040,N_18904,N_18820);
or U19041 (N_19041,N_18890,N_18910);
and U19042 (N_19042,N_18876,N_18976);
or U19043 (N_19043,N_18974,N_18912);
xnor U19044 (N_19044,N_18857,N_18802);
or U19045 (N_19045,N_18988,N_18905);
nand U19046 (N_19046,N_18818,N_18871);
xnor U19047 (N_19047,N_18935,N_18987);
or U19048 (N_19048,N_18859,N_18939);
and U19049 (N_19049,N_18836,N_18961);
or U19050 (N_19050,N_18809,N_18873);
and U19051 (N_19051,N_18980,N_18860);
nor U19052 (N_19052,N_18846,N_18982);
nand U19053 (N_19053,N_18800,N_18821);
and U19054 (N_19054,N_18919,N_18947);
xor U19055 (N_19055,N_18907,N_18825);
and U19056 (N_19056,N_18927,N_18930);
nor U19057 (N_19057,N_18962,N_18949);
and U19058 (N_19058,N_18887,N_18970);
or U19059 (N_19059,N_18901,N_18964);
nand U19060 (N_19060,N_18920,N_18834);
and U19061 (N_19061,N_18916,N_18812);
nor U19062 (N_19062,N_18863,N_18956);
nand U19063 (N_19063,N_18926,N_18866);
xor U19064 (N_19064,N_18898,N_18885);
nor U19065 (N_19065,N_18966,N_18824);
nand U19066 (N_19066,N_18831,N_18823);
or U19067 (N_19067,N_18883,N_18808);
or U19068 (N_19068,N_18994,N_18806);
xnor U19069 (N_19069,N_18828,N_18986);
nor U19070 (N_19070,N_18933,N_18989);
nor U19071 (N_19071,N_18958,N_18843);
xor U19072 (N_19072,N_18815,N_18979);
xor U19073 (N_19073,N_18884,N_18886);
nand U19074 (N_19074,N_18879,N_18942);
nand U19075 (N_19075,N_18877,N_18969);
and U19076 (N_19076,N_18813,N_18816);
and U19077 (N_19077,N_18853,N_18981);
nand U19078 (N_19078,N_18835,N_18895);
or U19079 (N_19079,N_18811,N_18913);
or U19080 (N_19080,N_18953,N_18955);
nor U19081 (N_19081,N_18841,N_18999);
and U19082 (N_19082,N_18996,N_18957);
nor U19083 (N_19083,N_18952,N_18915);
nor U19084 (N_19084,N_18861,N_18924);
or U19085 (N_19085,N_18971,N_18837);
or U19086 (N_19086,N_18968,N_18940);
nand U19087 (N_19087,N_18845,N_18899);
xnor U19088 (N_19088,N_18944,N_18851);
xnor U19089 (N_19089,N_18998,N_18977);
xnor U19090 (N_19090,N_18878,N_18908);
xor U19091 (N_19091,N_18827,N_18810);
and U19092 (N_19092,N_18931,N_18973);
and U19093 (N_19093,N_18948,N_18946);
nand U19094 (N_19094,N_18854,N_18840);
and U19095 (N_19095,N_18807,N_18872);
or U19096 (N_19096,N_18850,N_18819);
nor U19097 (N_19097,N_18984,N_18923);
xnor U19098 (N_19098,N_18838,N_18997);
xnor U19099 (N_19099,N_18862,N_18909);
nand U19100 (N_19100,N_18890,N_18985);
or U19101 (N_19101,N_18939,N_18825);
xnor U19102 (N_19102,N_18846,N_18814);
nor U19103 (N_19103,N_18930,N_18811);
nor U19104 (N_19104,N_18890,N_18832);
and U19105 (N_19105,N_18888,N_18858);
xor U19106 (N_19106,N_18962,N_18953);
nand U19107 (N_19107,N_18862,N_18851);
nand U19108 (N_19108,N_18916,N_18805);
or U19109 (N_19109,N_18857,N_18910);
or U19110 (N_19110,N_18983,N_18909);
nand U19111 (N_19111,N_18985,N_18814);
xnor U19112 (N_19112,N_18972,N_18847);
and U19113 (N_19113,N_18836,N_18908);
or U19114 (N_19114,N_18933,N_18878);
nor U19115 (N_19115,N_18867,N_18999);
nand U19116 (N_19116,N_18977,N_18814);
or U19117 (N_19117,N_18988,N_18933);
xnor U19118 (N_19118,N_18964,N_18897);
nand U19119 (N_19119,N_18808,N_18870);
and U19120 (N_19120,N_18948,N_18887);
nand U19121 (N_19121,N_18940,N_18819);
nor U19122 (N_19122,N_18877,N_18874);
nor U19123 (N_19123,N_18820,N_18907);
nor U19124 (N_19124,N_18826,N_18871);
nor U19125 (N_19125,N_18984,N_18832);
and U19126 (N_19126,N_18920,N_18978);
nor U19127 (N_19127,N_18826,N_18838);
or U19128 (N_19128,N_18899,N_18872);
xnor U19129 (N_19129,N_18983,N_18966);
or U19130 (N_19130,N_18971,N_18867);
and U19131 (N_19131,N_18822,N_18987);
nand U19132 (N_19132,N_18828,N_18901);
xnor U19133 (N_19133,N_18902,N_18982);
xnor U19134 (N_19134,N_18906,N_18964);
nand U19135 (N_19135,N_18962,N_18896);
and U19136 (N_19136,N_18881,N_18994);
xor U19137 (N_19137,N_18840,N_18820);
nand U19138 (N_19138,N_18973,N_18876);
xor U19139 (N_19139,N_18903,N_18880);
xor U19140 (N_19140,N_18945,N_18889);
nand U19141 (N_19141,N_18959,N_18863);
xnor U19142 (N_19142,N_18852,N_18871);
nor U19143 (N_19143,N_18874,N_18949);
xor U19144 (N_19144,N_18965,N_18931);
xnor U19145 (N_19145,N_18930,N_18850);
nor U19146 (N_19146,N_18839,N_18855);
nand U19147 (N_19147,N_18902,N_18989);
or U19148 (N_19148,N_18874,N_18970);
xnor U19149 (N_19149,N_18994,N_18890);
and U19150 (N_19150,N_18930,N_18880);
xnor U19151 (N_19151,N_18969,N_18812);
xnor U19152 (N_19152,N_18923,N_18863);
xnor U19153 (N_19153,N_18898,N_18916);
nand U19154 (N_19154,N_18872,N_18841);
or U19155 (N_19155,N_18866,N_18872);
nand U19156 (N_19156,N_18958,N_18886);
xnor U19157 (N_19157,N_18871,N_18919);
nor U19158 (N_19158,N_18899,N_18831);
and U19159 (N_19159,N_18868,N_18927);
and U19160 (N_19160,N_18922,N_18817);
and U19161 (N_19161,N_18877,N_18814);
or U19162 (N_19162,N_18982,N_18886);
xor U19163 (N_19163,N_18841,N_18876);
or U19164 (N_19164,N_18892,N_18890);
nor U19165 (N_19165,N_18983,N_18926);
nor U19166 (N_19166,N_18913,N_18918);
xor U19167 (N_19167,N_18933,N_18869);
nand U19168 (N_19168,N_18878,N_18920);
xnor U19169 (N_19169,N_18884,N_18883);
or U19170 (N_19170,N_18911,N_18988);
nand U19171 (N_19171,N_18917,N_18867);
and U19172 (N_19172,N_18946,N_18963);
and U19173 (N_19173,N_18874,N_18821);
or U19174 (N_19174,N_18883,N_18868);
xor U19175 (N_19175,N_18947,N_18959);
and U19176 (N_19176,N_18896,N_18830);
nor U19177 (N_19177,N_18884,N_18997);
nor U19178 (N_19178,N_18997,N_18910);
nand U19179 (N_19179,N_18871,N_18914);
and U19180 (N_19180,N_18990,N_18820);
nor U19181 (N_19181,N_18846,N_18968);
and U19182 (N_19182,N_18831,N_18840);
nand U19183 (N_19183,N_18991,N_18984);
or U19184 (N_19184,N_18956,N_18960);
xor U19185 (N_19185,N_18949,N_18868);
xor U19186 (N_19186,N_18918,N_18956);
and U19187 (N_19187,N_18895,N_18931);
or U19188 (N_19188,N_18895,N_18972);
or U19189 (N_19189,N_18850,N_18853);
xnor U19190 (N_19190,N_18981,N_18898);
nor U19191 (N_19191,N_18842,N_18933);
and U19192 (N_19192,N_18946,N_18827);
nor U19193 (N_19193,N_18947,N_18816);
and U19194 (N_19194,N_18889,N_18950);
nand U19195 (N_19195,N_18914,N_18844);
or U19196 (N_19196,N_18903,N_18935);
and U19197 (N_19197,N_18952,N_18956);
or U19198 (N_19198,N_18947,N_18849);
nand U19199 (N_19199,N_18898,N_18920);
nand U19200 (N_19200,N_19116,N_19049);
nand U19201 (N_19201,N_19059,N_19144);
nand U19202 (N_19202,N_19052,N_19147);
or U19203 (N_19203,N_19021,N_19075);
and U19204 (N_19204,N_19025,N_19104);
and U19205 (N_19205,N_19089,N_19031);
nor U19206 (N_19206,N_19030,N_19132);
nand U19207 (N_19207,N_19152,N_19118);
xnor U19208 (N_19208,N_19085,N_19166);
nand U19209 (N_19209,N_19157,N_19057);
xnor U19210 (N_19210,N_19051,N_19163);
nor U19211 (N_19211,N_19113,N_19047);
xnor U19212 (N_19212,N_19172,N_19107);
nor U19213 (N_19213,N_19150,N_19036);
or U19214 (N_19214,N_19156,N_19151);
xnor U19215 (N_19215,N_19190,N_19082);
and U19216 (N_19216,N_19187,N_19041);
xnor U19217 (N_19217,N_19142,N_19176);
and U19218 (N_19218,N_19022,N_19197);
and U19219 (N_19219,N_19159,N_19092);
nand U19220 (N_19220,N_19103,N_19110);
nand U19221 (N_19221,N_19066,N_19135);
xor U19222 (N_19222,N_19140,N_19122);
and U19223 (N_19223,N_19019,N_19018);
or U19224 (N_19224,N_19029,N_19027);
nand U19225 (N_19225,N_19042,N_19155);
nor U19226 (N_19226,N_19100,N_19112);
and U19227 (N_19227,N_19003,N_19183);
nor U19228 (N_19228,N_19148,N_19131);
xor U19229 (N_19229,N_19055,N_19121);
nand U19230 (N_19230,N_19081,N_19141);
or U19231 (N_19231,N_19069,N_19032);
and U19232 (N_19232,N_19138,N_19180);
nor U19233 (N_19233,N_19119,N_19145);
xor U19234 (N_19234,N_19050,N_19153);
and U19235 (N_19235,N_19053,N_19184);
nand U19236 (N_19236,N_19111,N_19181);
and U19237 (N_19237,N_19175,N_19012);
nand U19238 (N_19238,N_19136,N_19098);
xnor U19239 (N_19239,N_19005,N_19129);
nor U19240 (N_19240,N_19128,N_19164);
or U19241 (N_19241,N_19016,N_19035);
and U19242 (N_19242,N_19170,N_19126);
xor U19243 (N_19243,N_19045,N_19090);
xor U19244 (N_19244,N_19024,N_19039);
nand U19245 (N_19245,N_19173,N_19114);
nand U19246 (N_19246,N_19109,N_19010);
xor U19247 (N_19247,N_19179,N_19061);
nand U19248 (N_19248,N_19058,N_19014);
and U19249 (N_19249,N_19178,N_19023);
and U19250 (N_19250,N_19198,N_19068);
xnor U19251 (N_19251,N_19102,N_19185);
nor U19252 (N_19252,N_19087,N_19076);
nand U19253 (N_19253,N_19034,N_19088);
or U19254 (N_19254,N_19037,N_19086);
xor U19255 (N_19255,N_19004,N_19074);
nand U19256 (N_19256,N_19067,N_19007);
xor U19257 (N_19257,N_19192,N_19028);
xnor U19258 (N_19258,N_19070,N_19124);
or U19259 (N_19259,N_19149,N_19063);
or U19260 (N_19260,N_19191,N_19120);
or U19261 (N_19261,N_19026,N_19078);
and U19262 (N_19262,N_19096,N_19117);
xor U19263 (N_19263,N_19174,N_19084);
nor U19264 (N_19264,N_19002,N_19046);
or U19265 (N_19265,N_19013,N_19020);
nand U19266 (N_19266,N_19139,N_19099);
or U19267 (N_19267,N_19137,N_19162);
nand U19268 (N_19268,N_19094,N_19033);
and U19269 (N_19269,N_19091,N_19160);
nand U19270 (N_19270,N_19182,N_19154);
nor U19271 (N_19271,N_19009,N_19054);
nor U19272 (N_19272,N_19095,N_19134);
nor U19273 (N_19273,N_19189,N_19000);
and U19274 (N_19274,N_19186,N_19130);
xor U19275 (N_19275,N_19006,N_19056);
xnor U19276 (N_19276,N_19064,N_19093);
and U19277 (N_19277,N_19108,N_19177);
and U19278 (N_19278,N_19097,N_19017);
xnor U19279 (N_19279,N_19167,N_19196);
or U19280 (N_19280,N_19072,N_19188);
or U19281 (N_19281,N_19165,N_19195);
xnor U19282 (N_19282,N_19101,N_19062);
nor U19283 (N_19283,N_19143,N_19123);
and U19284 (N_19284,N_19106,N_19038);
nand U19285 (N_19285,N_19127,N_19105);
nor U19286 (N_19286,N_19125,N_19171);
nand U19287 (N_19287,N_19168,N_19133);
nor U19288 (N_19288,N_19077,N_19048);
nand U19289 (N_19289,N_19071,N_19080);
or U19290 (N_19290,N_19060,N_19043);
nand U19291 (N_19291,N_19040,N_19073);
and U19292 (N_19292,N_19044,N_19161);
or U19293 (N_19293,N_19199,N_19001);
xnor U19294 (N_19294,N_19146,N_19008);
xor U19295 (N_19295,N_19169,N_19115);
nor U19296 (N_19296,N_19065,N_19193);
xnor U19297 (N_19297,N_19158,N_19194);
nand U19298 (N_19298,N_19079,N_19015);
and U19299 (N_19299,N_19083,N_19011);
and U19300 (N_19300,N_19196,N_19040);
and U19301 (N_19301,N_19032,N_19074);
nand U19302 (N_19302,N_19160,N_19175);
and U19303 (N_19303,N_19030,N_19054);
xor U19304 (N_19304,N_19196,N_19023);
and U19305 (N_19305,N_19157,N_19099);
nand U19306 (N_19306,N_19046,N_19064);
nand U19307 (N_19307,N_19125,N_19015);
nand U19308 (N_19308,N_19140,N_19093);
and U19309 (N_19309,N_19034,N_19092);
nand U19310 (N_19310,N_19186,N_19085);
nand U19311 (N_19311,N_19077,N_19151);
or U19312 (N_19312,N_19174,N_19104);
and U19313 (N_19313,N_19120,N_19103);
xor U19314 (N_19314,N_19045,N_19096);
and U19315 (N_19315,N_19065,N_19194);
xor U19316 (N_19316,N_19042,N_19148);
nand U19317 (N_19317,N_19135,N_19091);
xnor U19318 (N_19318,N_19136,N_19092);
and U19319 (N_19319,N_19092,N_19066);
nand U19320 (N_19320,N_19193,N_19181);
or U19321 (N_19321,N_19092,N_19194);
and U19322 (N_19322,N_19111,N_19116);
xnor U19323 (N_19323,N_19041,N_19063);
or U19324 (N_19324,N_19052,N_19065);
nand U19325 (N_19325,N_19063,N_19078);
nor U19326 (N_19326,N_19078,N_19093);
or U19327 (N_19327,N_19180,N_19120);
or U19328 (N_19328,N_19177,N_19023);
nor U19329 (N_19329,N_19076,N_19106);
and U19330 (N_19330,N_19019,N_19020);
nand U19331 (N_19331,N_19068,N_19195);
and U19332 (N_19332,N_19159,N_19108);
xor U19333 (N_19333,N_19183,N_19133);
or U19334 (N_19334,N_19071,N_19103);
xnor U19335 (N_19335,N_19009,N_19138);
xor U19336 (N_19336,N_19018,N_19095);
or U19337 (N_19337,N_19124,N_19087);
nor U19338 (N_19338,N_19116,N_19165);
xor U19339 (N_19339,N_19142,N_19088);
nor U19340 (N_19340,N_19137,N_19009);
nor U19341 (N_19341,N_19126,N_19039);
and U19342 (N_19342,N_19024,N_19174);
and U19343 (N_19343,N_19115,N_19079);
or U19344 (N_19344,N_19029,N_19095);
and U19345 (N_19345,N_19175,N_19098);
nor U19346 (N_19346,N_19137,N_19026);
nand U19347 (N_19347,N_19015,N_19077);
nor U19348 (N_19348,N_19189,N_19029);
nor U19349 (N_19349,N_19070,N_19173);
or U19350 (N_19350,N_19191,N_19092);
or U19351 (N_19351,N_19159,N_19127);
xor U19352 (N_19352,N_19028,N_19144);
nand U19353 (N_19353,N_19008,N_19170);
nand U19354 (N_19354,N_19041,N_19093);
and U19355 (N_19355,N_19051,N_19154);
xor U19356 (N_19356,N_19097,N_19061);
and U19357 (N_19357,N_19121,N_19098);
nand U19358 (N_19358,N_19072,N_19191);
and U19359 (N_19359,N_19184,N_19024);
or U19360 (N_19360,N_19082,N_19067);
and U19361 (N_19361,N_19052,N_19149);
or U19362 (N_19362,N_19143,N_19170);
and U19363 (N_19363,N_19022,N_19119);
nor U19364 (N_19364,N_19160,N_19056);
xnor U19365 (N_19365,N_19165,N_19159);
and U19366 (N_19366,N_19143,N_19130);
nor U19367 (N_19367,N_19020,N_19191);
nor U19368 (N_19368,N_19031,N_19118);
nand U19369 (N_19369,N_19054,N_19011);
xor U19370 (N_19370,N_19152,N_19089);
or U19371 (N_19371,N_19179,N_19163);
or U19372 (N_19372,N_19043,N_19126);
and U19373 (N_19373,N_19154,N_19190);
or U19374 (N_19374,N_19113,N_19131);
or U19375 (N_19375,N_19134,N_19125);
xnor U19376 (N_19376,N_19047,N_19067);
or U19377 (N_19377,N_19177,N_19011);
xor U19378 (N_19378,N_19148,N_19094);
xnor U19379 (N_19379,N_19129,N_19069);
and U19380 (N_19380,N_19077,N_19026);
and U19381 (N_19381,N_19076,N_19042);
and U19382 (N_19382,N_19042,N_19074);
nor U19383 (N_19383,N_19165,N_19061);
nor U19384 (N_19384,N_19090,N_19175);
and U19385 (N_19385,N_19186,N_19074);
nor U19386 (N_19386,N_19184,N_19110);
xor U19387 (N_19387,N_19117,N_19186);
xnor U19388 (N_19388,N_19046,N_19061);
nor U19389 (N_19389,N_19038,N_19107);
xnor U19390 (N_19390,N_19022,N_19006);
and U19391 (N_19391,N_19176,N_19014);
or U19392 (N_19392,N_19073,N_19079);
or U19393 (N_19393,N_19095,N_19039);
nand U19394 (N_19394,N_19062,N_19087);
nor U19395 (N_19395,N_19000,N_19026);
and U19396 (N_19396,N_19141,N_19182);
and U19397 (N_19397,N_19081,N_19042);
nand U19398 (N_19398,N_19038,N_19132);
nand U19399 (N_19399,N_19166,N_19191);
nand U19400 (N_19400,N_19268,N_19358);
nor U19401 (N_19401,N_19350,N_19399);
nor U19402 (N_19402,N_19351,N_19306);
nand U19403 (N_19403,N_19390,N_19389);
and U19404 (N_19404,N_19342,N_19295);
xnor U19405 (N_19405,N_19285,N_19201);
and U19406 (N_19406,N_19259,N_19303);
nor U19407 (N_19407,N_19229,N_19353);
or U19408 (N_19408,N_19234,N_19383);
and U19409 (N_19409,N_19377,N_19224);
or U19410 (N_19410,N_19283,N_19324);
xnor U19411 (N_19411,N_19352,N_19311);
xnor U19412 (N_19412,N_19271,N_19305);
nand U19413 (N_19413,N_19322,N_19273);
xnor U19414 (N_19414,N_19378,N_19215);
or U19415 (N_19415,N_19262,N_19252);
nor U19416 (N_19416,N_19313,N_19277);
nand U19417 (N_19417,N_19255,N_19242);
nor U19418 (N_19418,N_19336,N_19343);
or U19419 (N_19419,N_19294,N_19357);
nor U19420 (N_19420,N_19220,N_19231);
or U19421 (N_19421,N_19361,N_19327);
nand U19422 (N_19422,N_19219,N_19301);
nand U19423 (N_19423,N_19335,N_19359);
or U19424 (N_19424,N_19360,N_19387);
nand U19425 (N_19425,N_19304,N_19310);
nand U19426 (N_19426,N_19369,N_19368);
nand U19427 (N_19427,N_19243,N_19302);
nand U19428 (N_19428,N_19209,N_19202);
nand U19429 (N_19429,N_19349,N_19372);
or U19430 (N_19430,N_19249,N_19348);
and U19431 (N_19431,N_19370,N_19320);
and U19432 (N_19432,N_19307,N_19221);
nor U19433 (N_19433,N_19275,N_19382);
nor U19434 (N_19434,N_19274,N_19269);
xnor U19435 (N_19435,N_19398,N_19338);
nor U19436 (N_19436,N_19256,N_19319);
nand U19437 (N_19437,N_19346,N_19250);
nand U19438 (N_19438,N_19270,N_19325);
xnor U19439 (N_19439,N_19254,N_19245);
xor U19440 (N_19440,N_19247,N_19300);
or U19441 (N_19441,N_19363,N_19225);
or U19442 (N_19442,N_19292,N_19396);
and U19443 (N_19443,N_19291,N_19272);
or U19444 (N_19444,N_19341,N_19241);
and U19445 (N_19445,N_19296,N_19276);
nor U19446 (N_19446,N_19263,N_19395);
xor U19447 (N_19447,N_19280,N_19200);
nand U19448 (N_19448,N_19355,N_19207);
or U19449 (N_19449,N_19235,N_19246);
nand U19450 (N_19450,N_19397,N_19212);
or U19451 (N_19451,N_19266,N_19205);
nand U19452 (N_19452,N_19384,N_19308);
or U19453 (N_19453,N_19344,N_19339);
xor U19454 (N_19454,N_19244,N_19366);
nor U19455 (N_19455,N_19340,N_19354);
nand U19456 (N_19456,N_19286,N_19380);
or U19457 (N_19457,N_19238,N_19248);
nand U19458 (N_19458,N_19203,N_19337);
nand U19459 (N_19459,N_19333,N_19282);
xor U19460 (N_19460,N_19317,N_19391);
and U19461 (N_19461,N_19253,N_19284);
nand U19462 (N_19462,N_19323,N_19293);
and U19463 (N_19463,N_19379,N_19251);
nand U19464 (N_19464,N_19329,N_19386);
and U19465 (N_19465,N_19206,N_19332);
and U19466 (N_19466,N_19297,N_19321);
and U19467 (N_19467,N_19385,N_19381);
nand U19468 (N_19468,N_19347,N_19218);
nor U19469 (N_19469,N_19394,N_19388);
nand U19470 (N_19470,N_19287,N_19240);
nor U19471 (N_19471,N_19289,N_19373);
xnor U19472 (N_19472,N_19376,N_19392);
xnor U19473 (N_19473,N_19318,N_19233);
or U19474 (N_19474,N_19261,N_19316);
nand U19475 (N_19475,N_19239,N_19211);
nor U19476 (N_19476,N_19264,N_19260);
xnor U19477 (N_19477,N_19393,N_19278);
xor U19478 (N_19478,N_19362,N_19237);
xnor U19479 (N_19479,N_19371,N_19279);
and U19480 (N_19480,N_19331,N_19204);
nand U19481 (N_19481,N_19257,N_19288);
or U19482 (N_19482,N_19281,N_19375);
xnor U19483 (N_19483,N_19265,N_19367);
nor U19484 (N_19484,N_19312,N_19345);
or U19485 (N_19485,N_19228,N_19365);
xnor U19486 (N_19486,N_19328,N_19227);
nor U19487 (N_19487,N_19216,N_19326);
or U19488 (N_19488,N_19222,N_19364);
nor U19489 (N_19489,N_19374,N_19290);
nand U19490 (N_19490,N_19314,N_19230);
nand U19491 (N_19491,N_19334,N_19213);
and U19492 (N_19492,N_19330,N_19298);
nor U19493 (N_19493,N_19299,N_19217);
xor U19494 (N_19494,N_19267,N_19315);
nand U19495 (N_19495,N_19236,N_19258);
or U19496 (N_19496,N_19223,N_19232);
xnor U19497 (N_19497,N_19226,N_19356);
nand U19498 (N_19498,N_19208,N_19210);
and U19499 (N_19499,N_19309,N_19214);
nand U19500 (N_19500,N_19259,N_19313);
nor U19501 (N_19501,N_19340,N_19201);
nor U19502 (N_19502,N_19293,N_19248);
xor U19503 (N_19503,N_19250,N_19344);
nand U19504 (N_19504,N_19350,N_19248);
and U19505 (N_19505,N_19391,N_19234);
xnor U19506 (N_19506,N_19238,N_19242);
xor U19507 (N_19507,N_19374,N_19202);
or U19508 (N_19508,N_19216,N_19307);
nand U19509 (N_19509,N_19373,N_19290);
nand U19510 (N_19510,N_19316,N_19315);
or U19511 (N_19511,N_19201,N_19388);
and U19512 (N_19512,N_19360,N_19331);
or U19513 (N_19513,N_19240,N_19371);
xnor U19514 (N_19514,N_19305,N_19257);
or U19515 (N_19515,N_19297,N_19349);
nor U19516 (N_19516,N_19367,N_19386);
or U19517 (N_19517,N_19207,N_19285);
nand U19518 (N_19518,N_19333,N_19252);
xor U19519 (N_19519,N_19205,N_19269);
xor U19520 (N_19520,N_19398,N_19211);
nand U19521 (N_19521,N_19296,N_19239);
nor U19522 (N_19522,N_19391,N_19314);
nor U19523 (N_19523,N_19281,N_19290);
and U19524 (N_19524,N_19301,N_19224);
and U19525 (N_19525,N_19293,N_19214);
and U19526 (N_19526,N_19252,N_19259);
nor U19527 (N_19527,N_19396,N_19210);
nor U19528 (N_19528,N_19368,N_19215);
and U19529 (N_19529,N_19357,N_19235);
nand U19530 (N_19530,N_19344,N_19357);
and U19531 (N_19531,N_19355,N_19301);
and U19532 (N_19532,N_19368,N_19248);
xnor U19533 (N_19533,N_19218,N_19328);
nand U19534 (N_19534,N_19356,N_19251);
xor U19535 (N_19535,N_19277,N_19398);
and U19536 (N_19536,N_19380,N_19295);
nor U19537 (N_19537,N_19308,N_19259);
and U19538 (N_19538,N_19385,N_19240);
or U19539 (N_19539,N_19234,N_19315);
nor U19540 (N_19540,N_19222,N_19200);
xnor U19541 (N_19541,N_19319,N_19276);
or U19542 (N_19542,N_19272,N_19313);
nand U19543 (N_19543,N_19208,N_19312);
or U19544 (N_19544,N_19387,N_19241);
or U19545 (N_19545,N_19225,N_19365);
xor U19546 (N_19546,N_19340,N_19261);
nand U19547 (N_19547,N_19206,N_19252);
and U19548 (N_19548,N_19320,N_19358);
nor U19549 (N_19549,N_19351,N_19325);
nand U19550 (N_19550,N_19282,N_19368);
xor U19551 (N_19551,N_19353,N_19286);
xnor U19552 (N_19552,N_19265,N_19307);
xnor U19553 (N_19553,N_19307,N_19294);
nor U19554 (N_19554,N_19342,N_19378);
xnor U19555 (N_19555,N_19290,N_19366);
nand U19556 (N_19556,N_19213,N_19388);
nor U19557 (N_19557,N_19214,N_19323);
xnor U19558 (N_19558,N_19219,N_19229);
and U19559 (N_19559,N_19285,N_19200);
and U19560 (N_19560,N_19362,N_19391);
and U19561 (N_19561,N_19229,N_19249);
nand U19562 (N_19562,N_19292,N_19281);
or U19563 (N_19563,N_19397,N_19396);
nand U19564 (N_19564,N_19399,N_19237);
nand U19565 (N_19565,N_19235,N_19275);
or U19566 (N_19566,N_19321,N_19225);
nor U19567 (N_19567,N_19369,N_19228);
and U19568 (N_19568,N_19240,N_19320);
nand U19569 (N_19569,N_19323,N_19381);
and U19570 (N_19570,N_19231,N_19225);
and U19571 (N_19571,N_19234,N_19322);
xnor U19572 (N_19572,N_19312,N_19250);
or U19573 (N_19573,N_19243,N_19275);
or U19574 (N_19574,N_19280,N_19250);
and U19575 (N_19575,N_19233,N_19341);
or U19576 (N_19576,N_19214,N_19269);
nor U19577 (N_19577,N_19293,N_19393);
nand U19578 (N_19578,N_19206,N_19339);
nand U19579 (N_19579,N_19366,N_19315);
or U19580 (N_19580,N_19268,N_19246);
nand U19581 (N_19581,N_19274,N_19285);
nor U19582 (N_19582,N_19365,N_19377);
or U19583 (N_19583,N_19368,N_19271);
nand U19584 (N_19584,N_19387,N_19254);
nand U19585 (N_19585,N_19249,N_19351);
nand U19586 (N_19586,N_19201,N_19301);
and U19587 (N_19587,N_19331,N_19292);
nor U19588 (N_19588,N_19358,N_19363);
xnor U19589 (N_19589,N_19374,N_19256);
nor U19590 (N_19590,N_19387,N_19261);
nor U19591 (N_19591,N_19385,N_19293);
xnor U19592 (N_19592,N_19245,N_19283);
nor U19593 (N_19593,N_19255,N_19288);
nand U19594 (N_19594,N_19311,N_19212);
xor U19595 (N_19595,N_19244,N_19316);
and U19596 (N_19596,N_19285,N_19322);
xor U19597 (N_19597,N_19286,N_19272);
xnor U19598 (N_19598,N_19211,N_19219);
nand U19599 (N_19599,N_19341,N_19276);
and U19600 (N_19600,N_19504,N_19586);
nor U19601 (N_19601,N_19513,N_19429);
nand U19602 (N_19602,N_19467,N_19556);
nand U19603 (N_19603,N_19541,N_19531);
nand U19604 (N_19604,N_19445,N_19580);
nor U19605 (N_19605,N_19506,N_19590);
nor U19606 (N_19606,N_19588,N_19446);
or U19607 (N_19607,N_19501,N_19426);
nand U19608 (N_19608,N_19497,N_19487);
xor U19609 (N_19609,N_19542,N_19557);
and U19610 (N_19610,N_19453,N_19536);
nor U19611 (N_19611,N_19544,N_19539);
and U19612 (N_19612,N_19428,N_19595);
or U19613 (N_19613,N_19495,N_19510);
or U19614 (N_19614,N_19416,N_19566);
nor U19615 (N_19615,N_19507,N_19465);
nand U19616 (N_19616,N_19441,N_19559);
xor U19617 (N_19617,N_19411,N_19458);
or U19618 (N_19618,N_19442,N_19420);
nor U19619 (N_19619,N_19524,N_19555);
and U19620 (N_19620,N_19597,N_19449);
nand U19621 (N_19621,N_19410,N_19460);
and U19622 (N_19622,N_19401,N_19422);
and U19623 (N_19623,N_19480,N_19424);
and U19624 (N_19624,N_19454,N_19552);
nand U19625 (N_19625,N_19477,N_19434);
nor U19626 (N_19626,N_19484,N_19514);
nor U19627 (N_19627,N_19415,N_19563);
and U19628 (N_19628,N_19550,N_19570);
xor U19629 (N_19629,N_19430,N_19599);
xor U19630 (N_19630,N_19578,N_19475);
nand U19631 (N_19631,N_19587,N_19526);
xnor U19632 (N_19632,N_19508,N_19469);
and U19633 (N_19633,N_19522,N_19400);
nand U19634 (N_19634,N_19538,N_19466);
nor U19635 (N_19635,N_19502,N_19461);
or U19636 (N_19636,N_19443,N_19521);
xor U19637 (N_19637,N_19523,N_19574);
nand U19638 (N_19638,N_19528,N_19565);
and U19639 (N_19639,N_19537,N_19432);
xor U19640 (N_19640,N_19575,N_19489);
nor U19641 (N_19641,N_19511,N_19455);
or U19642 (N_19642,N_19450,N_19562);
nor U19643 (N_19643,N_19463,N_19409);
nor U19644 (N_19644,N_19509,N_19560);
or U19645 (N_19645,N_19407,N_19515);
and U19646 (N_19646,N_19412,N_19518);
xor U19647 (N_19647,N_19483,N_19505);
nand U19648 (N_19648,N_19468,N_19421);
or U19649 (N_19649,N_19564,N_19473);
and U19650 (N_19650,N_19431,N_19533);
or U19651 (N_19651,N_19459,N_19568);
and U19652 (N_19652,N_19496,N_19553);
and U19653 (N_19653,N_19512,N_19543);
or U19654 (N_19654,N_19520,N_19457);
xor U19655 (N_19655,N_19589,N_19535);
and U19656 (N_19656,N_19585,N_19406);
and U19657 (N_19657,N_19579,N_19548);
nand U19658 (N_19658,N_19402,N_19593);
nand U19659 (N_19659,N_19481,N_19567);
nand U19660 (N_19660,N_19404,N_19494);
or U19661 (N_19661,N_19464,N_19525);
xor U19662 (N_19662,N_19476,N_19470);
xor U19663 (N_19663,N_19423,N_19478);
or U19664 (N_19664,N_19403,N_19427);
xor U19665 (N_19665,N_19516,N_19408);
xnor U19666 (N_19666,N_19500,N_19573);
nor U19667 (N_19667,N_19577,N_19547);
and U19668 (N_19668,N_19486,N_19435);
or U19669 (N_19669,N_19488,N_19554);
nand U19670 (N_19670,N_19456,N_19474);
nand U19671 (N_19671,N_19582,N_19437);
nand U19672 (N_19672,N_19546,N_19425);
and U19673 (N_19673,N_19485,N_19551);
nor U19674 (N_19674,N_19451,N_19482);
xnor U19675 (N_19675,N_19472,N_19592);
xor U19676 (N_19676,N_19436,N_19576);
xnor U19677 (N_19677,N_19444,N_19413);
or U19678 (N_19678,N_19492,N_19405);
nor U19679 (N_19679,N_19591,N_19545);
xor U19680 (N_19680,N_19558,N_19491);
xor U19681 (N_19681,N_19471,N_19503);
or U19682 (N_19682,N_19534,N_19572);
xor U19683 (N_19683,N_19414,N_19440);
and U19684 (N_19684,N_19571,N_19561);
and U19685 (N_19685,N_19493,N_19594);
nand U19686 (N_19686,N_19540,N_19530);
and U19687 (N_19687,N_19569,N_19462);
or U19688 (N_19688,N_19418,N_19419);
nor U19689 (N_19689,N_19452,N_19598);
nor U19690 (N_19690,N_19479,N_19583);
nor U19691 (N_19691,N_19581,N_19448);
nor U19692 (N_19692,N_19499,N_19517);
nor U19693 (N_19693,N_19519,N_19532);
nand U19694 (N_19694,N_19527,N_19433);
xor U19695 (N_19695,N_19498,N_19596);
nor U19696 (N_19696,N_19439,N_19584);
nor U19697 (N_19697,N_19417,N_19529);
nor U19698 (N_19698,N_19447,N_19549);
nor U19699 (N_19699,N_19490,N_19438);
or U19700 (N_19700,N_19503,N_19467);
nand U19701 (N_19701,N_19579,N_19404);
nand U19702 (N_19702,N_19572,N_19562);
or U19703 (N_19703,N_19422,N_19589);
and U19704 (N_19704,N_19590,N_19408);
or U19705 (N_19705,N_19403,N_19413);
nand U19706 (N_19706,N_19435,N_19578);
xor U19707 (N_19707,N_19478,N_19582);
and U19708 (N_19708,N_19539,N_19431);
nor U19709 (N_19709,N_19543,N_19565);
or U19710 (N_19710,N_19466,N_19432);
nor U19711 (N_19711,N_19468,N_19413);
nand U19712 (N_19712,N_19461,N_19554);
and U19713 (N_19713,N_19401,N_19508);
and U19714 (N_19714,N_19572,N_19513);
or U19715 (N_19715,N_19591,N_19493);
and U19716 (N_19716,N_19479,N_19554);
and U19717 (N_19717,N_19468,N_19488);
nor U19718 (N_19718,N_19475,N_19492);
and U19719 (N_19719,N_19519,N_19514);
or U19720 (N_19720,N_19595,N_19578);
nand U19721 (N_19721,N_19419,N_19516);
or U19722 (N_19722,N_19417,N_19572);
xor U19723 (N_19723,N_19418,N_19574);
and U19724 (N_19724,N_19490,N_19432);
nor U19725 (N_19725,N_19445,N_19402);
nand U19726 (N_19726,N_19584,N_19585);
or U19727 (N_19727,N_19451,N_19496);
or U19728 (N_19728,N_19470,N_19593);
and U19729 (N_19729,N_19516,N_19495);
or U19730 (N_19730,N_19538,N_19571);
nand U19731 (N_19731,N_19489,N_19551);
nor U19732 (N_19732,N_19504,N_19593);
or U19733 (N_19733,N_19525,N_19548);
xor U19734 (N_19734,N_19576,N_19538);
nor U19735 (N_19735,N_19559,N_19556);
nor U19736 (N_19736,N_19521,N_19440);
xor U19737 (N_19737,N_19593,N_19574);
nand U19738 (N_19738,N_19585,N_19421);
nor U19739 (N_19739,N_19426,N_19402);
nand U19740 (N_19740,N_19595,N_19447);
or U19741 (N_19741,N_19498,N_19597);
nand U19742 (N_19742,N_19500,N_19471);
xnor U19743 (N_19743,N_19457,N_19515);
and U19744 (N_19744,N_19542,N_19514);
nand U19745 (N_19745,N_19510,N_19541);
nand U19746 (N_19746,N_19501,N_19439);
or U19747 (N_19747,N_19492,N_19484);
xnor U19748 (N_19748,N_19434,N_19454);
xor U19749 (N_19749,N_19423,N_19411);
nor U19750 (N_19750,N_19445,N_19508);
and U19751 (N_19751,N_19493,N_19408);
nand U19752 (N_19752,N_19597,N_19477);
xor U19753 (N_19753,N_19457,N_19578);
xor U19754 (N_19754,N_19541,N_19496);
or U19755 (N_19755,N_19406,N_19562);
xnor U19756 (N_19756,N_19546,N_19544);
and U19757 (N_19757,N_19464,N_19491);
and U19758 (N_19758,N_19466,N_19409);
nor U19759 (N_19759,N_19491,N_19436);
xor U19760 (N_19760,N_19493,N_19446);
xnor U19761 (N_19761,N_19513,N_19435);
nand U19762 (N_19762,N_19406,N_19450);
nor U19763 (N_19763,N_19593,N_19449);
xor U19764 (N_19764,N_19584,N_19418);
xnor U19765 (N_19765,N_19415,N_19483);
or U19766 (N_19766,N_19595,N_19479);
and U19767 (N_19767,N_19494,N_19528);
nor U19768 (N_19768,N_19477,N_19469);
and U19769 (N_19769,N_19552,N_19472);
or U19770 (N_19770,N_19444,N_19488);
nand U19771 (N_19771,N_19531,N_19534);
and U19772 (N_19772,N_19472,N_19590);
and U19773 (N_19773,N_19529,N_19508);
or U19774 (N_19774,N_19557,N_19556);
xnor U19775 (N_19775,N_19598,N_19579);
nand U19776 (N_19776,N_19569,N_19466);
or U19777 (N_19777,N_19527,N_19487);
xor U19778 (N_19778,N_19477,N_19443);
nor U19779 (N_19779,N_19546,N_19423);
nand U19780 (N_19780,N_19532,N_19400);
nor U19781 (N_19781,N_19583,N_19411);
or U19782 (N_19782,N_19549,N_19414);
xnor U19783 (N_19783,N_19569,N_19512);
or U19784 (N_19784,N_19581,N_19463);
xnor U19785 (N_19785,N_19458,N_19599);
nor U19786 (N_19786,N_19573,N_19416);
and U19787 (N_19787,N_19460,N_19588);
nand U19788 (N_19788,N_19546,N_19443);
and U19789 (N_19789,N_19448,N_19546);
and U19790 (N_19790,N_19567,N_19409);
xor U19791 (N_19791,N_19584,N_19548);
nand U19792 (N_19792,N_19500,N_19555);
xnor U19793 (N_19793,N_19536,N_19589);
nor U19794 (N_19794,N_19519,N_19425);
or U19795 (N_19795,N_19488,N_19427);
nor U19796 (N_19796,N_19544,N_19585);
xnor U19797 (N_19797,N_19570,N_19546);
xnor U19798 (N_19798,N_19430,N_19511);
nand U19799 (N_19799,N_19598,N_19541);
xor U19800 (N_19800,N_19612,N_19787);
or U19801 (N_19801,N_19722,N_19622);
or U19802 (N_19802,N_19662,N_19777);
xnor U19803 (N_19803,N_19758,N_19682);
nor U19804 (N_19804,N_19626,N_19608);
xor U19805 (N_19805,N_19679,N_19779);
nand U19806 (N_19806,N_19708,N_19646);
xor U19807 (N_19807,N_19645,N_19761);
nand U19808 (N_19808,N_19638,N_19664);
nand U19809 (N_19809,N_19794,N_19668);
nand U19810 (N_19810,N_19629,N_19716);
xor U19811 (N_19811,N_19654,N_19760);
or U19812 (N_19812,N_19737,N_19661);
nor U19813 (N_19813,N_19653,N_19755);
and U19814 (N_19814,N_19730,N_19764);
and U19815 (N_19815,N_19727,N_19799);
or U19816 (N_19816,N_19718,N_19632);
xnor U19817 (N_19817,N_19619,N_19655);
or U19818 (N_19818,N_19667,N_19610);
or U19819 (N_19819,N_19620,N_19773);
nand U19820 (N_19820,N_19607,N_19770);
xnor U19821 (N_19821,N_19688,N_19691);
nand U19822 (N_19822,N_19651,N_19757);
nand U19823 (N_19823,N_19750,N_19658);
or U19824 (N_19824,N_19639,N_19657);
nand U19825 (N_19825,N_19603,N_19636);
or U19826 (N_19826,N_19643,N_19644);
xnor U19827 (N_19827,N_19614,N_19685);
nor U19828 (N_19828,N_19736,N_19713);
nor U19829 (N_19829,N_19683,N_19623);
xnor U19830 (N_19830,N_19738,N_19707);
and U19831 (N_19831,N_19774,N_19746);
nand U19832 (N_19832,N_19648,N_19768);
nor U19833 (N_19833,N_19676,N_19624);
nand U19834 (N_19834,N_19717,N_19641);
xnor U19835 (N_19835,N_19635,N_19696);
and U19836 (N_19836,N_19631,N_19686);
xnor U19837 (N_19837,N_19634,N_19744);
or U19838 (N_19838,N_19725,N_19652);
or U19839 (N_19839,N_19678,N_19756);
nand U19840 (N_19840,N_19618,N_19649);
nand U19841 (N_19841,N_19609,N_19659);
nand U19842 (N_19842,N_19621,N_19711);
xnor U19843 (N_19843,N_19765,N_19743);
xnor U19844 (N_19844,N_19791,N_19766);
nand U19845 (N_19845,N_19798,N_19702);
xor U19846 (N_19846,N_19642,N_19606);
or U19847 (N_19847,N_19630,N_19703);
nor U19848 (N_19848,N_19650,N_19778);
nand U19849 (N_19849,N_19769,N_19796);
xnor U19850 (N_19850,N_19749,N_19693);
xnor U19851 (N_19851,N_19613,N_19782);
and U19852 (N_19852,N_19669,N_19742);
nand U19853 (N_19853,N_19786,N_19660);
xor U19854 (N_19854,N_19759,N_19771);
xnor U19855 (N_19855,N_19724,N_19627);
nand U19856 (N_19856,N_19602,N_19780);
nand U19857 (N_19857,N_19704,N_19692);
or U19858 (N_19858,N_19748,N_19640);
or U19859 (N_19859,N_19617,N_19677);
xnor U19860 (N_19860,N_19767,N_19754);
and U19861 (N_19861,N_19785,N_19605);
and U19862 (N_19862,N_19735,N_19732);
nand U19863 (N_19863,N_19751,N_19734);
nor U19864 (N_19864,N_19781,N_19752);
xnor U19865 (N_19865,N_19675,N_19611);
and U19866 (N_19866,N_19710,N_19689);
nor U19867 (N_19867,N_19628,N_19687);
or U19868 (N_19868,N_19731,N_19753);
nor U19869 (N_19869,N_19666,N_19728);
or U19870 (N_19870,N_19705,N_19776);
nand U19871 (N_19871,N_19699,N_19615);
nand U19872 (N_19872,N_19795,N_19747);
nor U19873 (N_19873,N_19763,N_19772);
nand U19874 (N_19874,N_19709,N_19633);
nor U19875 (N_19875,N_19694,N_19793);
xnor U19876 (N_19876,N_19745,N_19601);
xnor U19877 (N_19877,N_19670,N_19604);
and U19878 (N_19878,N_19726,N_19625);
and U19879 (N_19879,N_19647,N_19680);
xnor U19880 (N_19880,N_19600,N_19719);
xnor U19881 (N_19881,N_19681,N_19706);
nor U19882 (N_19882,N_19695,N_19733);
nor U19883 (N_19883,N_19762,N_19690);
xor U19884 (N_19884,N_19783,N_19698);
xor U19885 (N_19885,N_19797,N_19721);
and U19886 (N_19886,N_19663,N_19701);
nand U19887 (N_19887,N_19720,N_19739);
or U19888 (N_19888,N_19697,N_19789);
or U19889 (N_19889,N_19784,N_19616);
xnor U19890 (N_19890,N_19790,N_19741);
and U19891 (N_19891,N_19637,N_19792);
or U19892 (N_19892,N_19671,N_19674);
or U19893 (N_19893,N_19700,N_19656);
nor U19894 (N_19894,N_19788,N_19672);
nand U19895 (N_19895,N_19665,N_19729);
and U19896 (N_19896,N_19712,N_19684);
and U19897 (N_19897,N_19775,N_19723);
nor U19898 (N_19898,N_19740,N_19714);
and U19899 (N_19899,N_19715,N_19673);
and U19900 (N_19900,N_19678,N_19657);
xor U19901 (N_19901,N_19735,N_19680);
nor U19902 (N_19902,N_19680,N_19618);
nand U19903 (N_19903,N_19605,N_19773);
nand U19904 (N_19904,N_19623,N_19744);
and U19905 (N_19905,N_19648,N_19795);
nor U19906 (N_19906,N_19650,N_19644);
or U19907 (N_19907,N_19729,N_19636);
or U19908 (N_19908,N_19754,N_19641);
or U19909 (N_19909,N_19702,N_19621);
and U19910 (N_19910,N_19711,N_19678);
and U19911 (N_19911,N_19659,N_19744);
nand U19912 (N_19912,N_19664,N_19781);
xnor U19913 (N_19913,N_19716,N_19740);
xnor U19914 (N_19914,N_19744,N_19714);
and U19915 (N_19915,N_19640,N_19698);
nand U19916 (N_19916,N_19756,N_19690);
nand U19917 (N_19917,N_19700,N_19635);
xor U19918 (N_19918,N_19765,N_19654);
and U19919 (N_19919,N_19723,N_19799);
or U19920 (N_19920,N_19735,N_19624);
or U19921 (N_19921,N_19734,N_19672);
nor U19922 (N_19922,N_19601,N_19656);
or U19923 (N_19923,N_19656,N_19755);
nand U19924 (N_19924,N_19775,N_19603);
nor U19925 (N_19925,N_19727,N_19718);
nor U19926 (N_19926,N_19665,N_19792);
xnor U19927 (N_19927,N_19610,N_19769);
nor U19928 (N_19928,N_19789,N_19675);
and U19929 (N_19929,N_19724,N_19707);
nor U19930 (N_19930,N_19649,N_19653);
nor U19931 (N_19931,N_19773,N_19779);
or U19932 (N_19932,N_19750,N_19718);
nor U19933 (N_19933,N_19780,N_19656);
xnor U19934 (N_19934,N_19798,N_19634);
and U19935 (N_19935,N_19651,N_19767);
and U19936 (N_19936,N_19766,N_19602);
xor U19937 (N_19937,N_19791,N_19705);
xor U19938 (N_19938,N_19626,N_19768);
nor U19939 (N_19939,N_19608,N_19714);
xor U19940 (N_19940,N_19625,N_19706);
nand U19941 (N_19941,N_19702,N_19772);
nor U19942 (N_19942,N_19721,N_19704);
and U19943 (N_19943,N_19749,N_19793);
or U19944 (N_19944,N_19688,N_19729);
nor U19945 (N_19945,N_19634,N_19648);
xnor U19946 (N_19946,N_19685,N_19625);
xor U19947 (N_19947,N_19677,N_19628);
nor U19948 (N_19948,N_19746,N_19769);
and U19949 (N_19949,N_19792,N_19745);
and U19950 (N_19950,N_19694,N_19607);
and U19951 (N_19951,N_19736,N_19775);
nor U19952 (N_19952,N_19611,N_19764);
nand U19953 (N_19953,N_19770,N_19746);
nor U19954 (N_19954,N_19633,N_19753);
or U19955 (N_19955,N_19749,N_19796);
nor U19956 (N_19956,N_19740,N_19610);
and U19957 (N_19957,N_19642,N_19728);
nor U19958 (N_19958,N_19647,N_19628);
or U19959 (N_19959,N_19769,N_19786);
nor U19960 (N_19960,N_19796,N_19685);
and U19961 (N_19961,N_19611,N_19610);
or U19962 (N_19962,N_19706,N_19739);
nand U19963 (N_19963,N_19755,N_19686);
nand U19964 (N_19964,N_19625,N_19797);
and U19965 (N_19965,N_19726,N_19795);
xnor U19966 (N_19966,N_19608,N_19761);
nor U19967 (N_19967,N_19788,N_19775);
and U19968 (N_19968,N_19637,N_19706);
xor U19969 (N_19969,N_19750,N_19683);
nand U19970 (N_19970,N_19624,N_19673);
and U19971 (N_19971,N_19793,N_19665);
nor U19972 (N_19972,N_19654,N_19706);
or U19973 (N_19973,N_19775,N_19792);
and U19974 (N_19974,N_19665,N_19682);
and U19975 (N_19975,N_19702,N_19759);
nand U19976 (N_19976,N_19610,N_19796);
nor U19977 (N_19977,N_19630,N_19739);
and U19978 (N_19978,N_19720,N_19767);
nand U19979 (N_19979,N_19768,N_19657);
or U19980 (N_19980,N_19655,N_19682);
xnor U19981 (N_19981,N_19733,N_19776);
or U19982 (N_19982,N_19605,N_19778);
nand U19983 (N_19983,N_19758,N_19694);
and U19984 (N_19984,N_19734,N_19695);
or U19985 (N_19985,N_19743,N_19636);
nand U19986 (N_19986,N_19610,N_19757);
and U19987 (N_19987,N_19761,N_19714);
or U19988 (N_19988,N_19690,N_19712);
and U19989 (N_19989,N_19690,N_19735);
or U19990 (N_19990,N_19794,N_19648);
and U19991 (N_19991,N_19624,N_19783);
or U19992 (N_19992,N_19636,N_19721);
or U19993 (N_19993,N_19744,N_19756);
nor U19994 (N_19994,N_19771,N_19749);
or U19995 (N_19995,N_19657,N_19777);
and U19996 (N_19996,N_19636,N_19780);
or U19997 (N_19997,N_19692,N_19708);
nand U19998 (N_19998,N_19611,N_19617);
nand U19999 (N_19999,N_19696,N_19748);
or UO_0 (O_0,N_19864,N_19939);
nor UO_1 (O_1,N_19933,N_19840);
xnor UO_2 (O_2,N_19859,N_19959);
nand UO_3 (O_3,N_19874,N_19922);
xnor UO_4 (O_4,N_19876,N_19888);
and UO_5 (O_5,N_19813,N_19992);
nor UO_6 (O_6,N_19845,N_19896);
and UO_7 (O_7,N_19911,N_19898);
and UO_8 (O_8,N_19804,N_19946);
nand UO_9 (O_9,N_19853,N_19997);
or UO_10 (O_10,N_19908,N_19953);
nor UO_11 (O_11,N_19826,N_19971);
or UO_12 (O_12,N_19818,N_19968);
nand UO_13 (O_13,N_19963,N_19871);
and UO_14 (O_14,N_19920,N_19865);
or UO_15 (O_15,N_19944,N_19935);
nand UO_16 (O_16,N_19949,N_19857);
xor UO_17 (O_17,N_19975,N_19952);
nand UO_18 (O_18,N_19879,N_19885);
and UO_19 (O_19,N_19916,N_19881);
nand UO_20 (O_20,N_19834,N_19926);
nor UO_21 (O_21,N_19937,N_19900);
nor UO_22 (O_22,N_19895,N_19979);
xor UO_23 (O_23,N_19855,N_19832);
or UO_24 (O_24,N_19928,N_19849);
xnor UO_25 (O_25,N_19987,N_19852);
or UO_26 (O_26,N_19886,N_19915);
nand UO_27 (O_27,N_19810,N_19800);
xnor UO_28 (O_28,N_19829,N_19812);
nor UO_29 (O_29,N_19956,N_19996);
xor UO_30 (O_30,N_19972,N_19977);
or UO_31 (O_31,N_19938,N_19904);
or UO_32 (O_32,N_19878,N_19986);
nand UO_33 (O_33,N_19927,N_19883);
or UO_34 (O_34,N_19846,N_19993);
nor UO_35 (O_35,N_19868,N_19901);
nand UO_36 (O_36,N_19894,N_19912);
or UO_37 (O_37,N_19947,N_19801);
xor UO_38 (O_38,N_19899,N_19941);
and UO_39 (O_39,N_19906,N_19966);
or UO_40 (O_40,N_19842,N_19998);
nand UO_41 (O_41,N_19995,N_19930);
xnor UO_42 (O_42,N_19823,N_19847);
and UO_43 (O_43,N_19817,N_19809);
xnor UO_44 (O_44,N_19831,N_19989);
xnor UO_45 (O_45,N_19839,N_19820);
nand UO_46 (O_46,N_19918,N_19863);
nand UO_47 (O_47,N_19982,N_19821);
nor UO_48 (O_48,N_19836,N_19976);
nor UO_49 (O_49,N_19882,N_19805);
or UO_50 (O_50,N_19970,N_19962);
nor UO_51 (O_51,N_19932,N_19880);
xnor UO_52 (O_52,N_19897,N_19929);
nand UO_53 (O_53,N_19910,N_19940);
or UO_54 (O_54,N_19965,N_19887);
or UO_55 (O_55,N_19811,N_19819);
xnor UO_56 (O_56,N_19942,N_19914);
nand UO_57 (O_57,N_19978,N_19858);
xor UO_58 (O_58,N_19923,N_19990);
and UO_59 (O_59,N_19999,N_19815);
and UO_60 (O_60,N_19960,N_19984);
and UO_61 (O_61,N_19974,N_19850);
and UO_62 (O_62,N_19967,N_19893);
xnor UO_63 (O_63,N_19891,N_19827);
and UO_64 (O_64,N_19951,N_19843);
and UO_65 (O_65,N_19903,N_19985);
nand UO_66 (O_66,N_19860,N_19892);
nor UO_67 (O_67,N_19835,N_19861);
or UO_68 (O_68,N_19943,N_19919);
xnor UO_69 (O_69,N_19803,N_19924);
xnor UO_70 (O_70,N_19913,N_19866);
nand UO_71 (O_71,N_19807,N_19961);
and UO_72 (O_72,N_19950,N_19925);
or UO_73 (O_73,N_19981,N_19958);
xnor UO_74 (O_74,N_19802,N_19830);
and UO_75 (O_75,N_19889,N_19964);
xnor UO_76 (O_76,N_19867,N_19917);
or UO_77 (O_77,N_19870,N_19856);
nor UO_78 (O_78,N_19921,N_19988);
or UO_79 (O_79,N_19851,N_19907);
or UO_80 (O_80,N_19983,N_19973);
and UO_81 (O_81,N_19877,N_19862);
and UO_82 (O_82,N_19806,N_19844);
nor UO_83 (O_83,N_19824,N_19890);
or UO_84 (O_84,N_19948,N_19934);
xor UO_85 (O_85,N_19825,N_19969);
nor UO_86 (O_86,N_19854,N_19902);
nand UO_87 (O_87,N_19822,N_19872);
nor UO_88 (O_88,N_19875,N_19869);
nand UO_89 (O_89,N_19884,N_19837);
and UO_90 (O_90,N_19955,N_19994);
nor UO_91 (O_91,N_19954,N_19931);
nor UO_92 (O_92,N_19945,N_19873);
nor UO_93 (O_93,N_19828,N_19936);
or UO_94 (O_94,N_19838,N_19909);
nor UO_95 (O_95,N_19833,N_19991);
and UO_96 (O_96,N_19816,N_19980);
and UO_97 (O_97,N_19808,N_19841);
xnor UO_98 (O_98,N_19848,N_19957);
nor UO_99 (O_99,N_19814,N_19905);
or UO_100 (O_100,N_19807,N_19919);
nor UO_101 (O_101,N_19954,N_19899);
nor UO_102 (O_102,N_19951,N_19925);
or UO_103 (O_103,N_19913,N_19954);
xor UO_104 (O_104,N_19960,N_19815);
xnor UO_105 (O_105,N_19830,N_19890);
and UO_106 (O_106,N_19973,N_19956);
or UO_107 (O_107,N_19980,N_19800);
xnor UO_108 (O_108,N_19890,N_19884);
nand UO_109 (O_109,N_19995,N_19968);
and UO_110 (O_110,N_19811,N_19962);
nor UO_111 (O_111,N_19814,N_19823);
nand UO_112 (O_112,N_19972,N_19981);
and UO_113 (O_113,N_19897,N_19828);
or UO_114 (O_114,N_19983,N_19807);
or UO_115 (O_115,N_19883,N_19803);
nor UO_116 (O_116,N_19964,N_19941);
or UO_117 (O_117,N_19879,N_19828);
or UO_118 (O_118,N_19932,N_19824);
nor UO_119 (O_119,N_19898,N_19972);
xnor UO_120 (O_120,N_19858,N_19996);
or UO_121 (O_121,N_19927,N_19967);
or UO_122 (O_122,N_19930,N_19861);
and UO_123 (O_123,N_19870,N_19815);
and UO_124 (O_124,N_19820,N_19933);
nor UO_125 (O_125,N_19815,N_19965);
xor UO_126 (O_126,N_19803,N_19997);
or UO_127 (O_127,N_19935,N_19877);
and UO_128 (O_128,N_19998,N_19872);
xnor UO_129 (O_129,N_19897,N_19935);
nand UO_130 (O_130,N_19894,N_19818);
or UO_131 (O_131,N_19988,N_19813);
xnor UO_132 (O_132,N_19885,N_19842);
and UO_133 (O_133,N_19852,N_19983);
or UO_134 (O_134,N_19886,N_19817);
or UO_135 (O_135,N_19806,N_19870);
nor UO_136 (O_136,N_19943,N_19986);
and UO_137 (O_137,N_19915,N_19951);
nor UO_138 (O_138,N_19841,N_19992);
xor UO_139 (O_139,N_19984,N_19941);
nor UO_140 (O_140,N_19855,N_19953);
or UO_141 (O_141,N_19983,N_19800);
xnor UO_142 (O_142,N_19881,N_19891);
nand UO_143 (O_143,N_19862,N_19826);
nor UO_144 (O_144,N_19950,N_19835);
and UO_145 (O_145,N_19955,N_19924);
nor UO_146 (O_146,N_19884,N_19882);
nor UO_147 (O_147,N_19936,N_19942);
and UO_148 (O_148,N_19955,N_19995);
nor UO_149 (O_149,N_19828,N_19964);
nor UO_150 (O_150,N_19832,N_19882);
or UO_151 (O_151,N_19819,N_19930);
xor UO_152 (O_152,N_19955,N_19867);
nor UO_153 (O_153,N_19960,N_19945);
or UO_154 (O_154,N_19960,N_19840);
nor UO_155 (O_155,N_19907,N_19953);
nor UO_156 (O_156,N_19923,N_19940);
nor UO_157 (O_157,N_19984,N_19904);
xnor UO_158 (O_158,N_19840,N_19805);
xnor UO_159 (O_159,N_19830,N_19955);
xnor UO_160 (O_160,N_19988,N_19875);
and UO_161 (O_161,N_19860,N_19959);
nand UO_162 (O_162,N_19878,N_19966);
nand UO_163 (O_163,N_19808,N_19993);
nor UO_164 (O_164,N_19804,N_19816);
nand UO_165 (O_165,N_19830,N_19900);
xor UO_166 (O_166,N_19914,N_19997);
nor UO_167 (O_167,N_19803,N_19834);
nand UO_168 (O_168,N_19855,N_19811);
nand UO_169 (O_169,N_19833,N_19899);
nand UO_170 (O_170,N_19914,N_19929);
xor UO_171 (O_171,N_19851,N_19835);
and UO_172 (O_172,N_19841,N_19856);
nand UO_173 (O_173,N_19951,N_19965);
nor UO_174 (O_174,N_19842,N_19810);
nand UO_175 (O_175,N_19805,N_19812);
nor UO_176 (O_176,N_19960,N_19846);
nand UO_177 (O_177,N_19999,N_19857);
xnor UO_178 (O_178,N_19900,N_19912);
xor UO_179 (O_179,N_19879,N_19975);
xnor UO_180 (O_180,N_19979,N_19811);
or UO_181 (O_181,N_19973,N_19977);
nor UO_182 (O_182,N_19902,N_19940);
or UO_183 (O_183,N_19873,N_19991);
or UO_184 (O_184,N_19960,N_19905);
or UO_185 (O_185,N_19893,N_19952);
nor UO_186 (O_186,N_19927,N_19900);
xnor UO_187 (O_187,N_19990,N_19905);
and UO_188 (O_188,N_19837,N_19840);
or UO_189 (O_189,N_19999,N_19912);
nand UO_190 (O_190,N_19977,N_19824);
and UO_191 (O_191,N_19937,N_19973);
nand UO_192 (O_192,N_19936,N_19967);
xnor UO_193 (O_193,N_19941,N_19895);
nor UO_194 (O_194,N_19879,N_19821);
and UO_195 (O_195,N_19869,N_19977);
or UO_196 (O_196,N_19813,N_19868);
nor UO_197 (O_197,N_19843,N_19912);
and UO_198 (O_198,N_19923,N_19902);
or UO_199 (O_199,N_19878,N_19928);
and UO_200 (O_200,N_19810,N_19957);
xnor UO_201 (O_201,N_19991,N_19852);
xnor UO_202 (O_202,N_19806,N_19887);
xor UO_203 (O_203,N_19918,N_19957);
or UO_204 (O_204,N_19962,N_19940);
or UO_205 (O_205,N_19996,N_19988);
nand UO_206 (O_206,N_19860,N_19943);
or UO_207 (O_207,N_19969,N_19851);
nor UO_208 (O_208,N_19976,N_19919);
nand UO_209 (O_209,N_19958,N_19950);
xor UO_210 (O_210,N_19915,N_19972);
xnor UO_211 (O_211,N_19817,N_19959);
xnor UO_212 (O_212,N_19945,N_19919);
nor UO_213 (O_213,N_19902,N_19979);
nand UO_214 (O_214,N_19860,N_19837);
nand UO_215 (O_215,N_19911,N_19875);
and UO_216 (O_216,N_19971,N_19872);
xor UO_217 (O_217,N_19905,N_19897);
or UO_218 (O_218,N_19855,N_19914);
and UO_219 (O_219,N_19908,N_19993);
nor UO_220 (O_220,N_19879,N_19924);
xor UO_221 (O_221,N_19964,N_19980);
or UO_222 (O_222,N_19949,N_19969);
and UO_223 (O_223,N_19988,N_19824);
or UO_224 (O_224,N_19832,N_19950);
or UO_225 (O_225,N_19817,N_19824);
xnor UO_226 (O_226,N_19851,N_19818);
and UO_227 (O_227,N_19872,N_19973);
and UO_228 (O_228,N_19842,N_19928);
and UO_229 (O_229,N_19841,N_19955);
nor UO_230 (O_230,N_19812,N_19959);
nor UO_231 (O_231,N_19867,N_19810);
nand UO_232 (O_232,N_19998,N_19992);
xor UO_233 (O_233,N_19895,N_19828);
nor UO_234 (O_234,N_19988,N_19897);
or UO_235 (O_235,N_19825,N_19810);
and UO_236 (O_236,N_19892,N_19836);
and UO_237 (O_237,N_19967,N_19926);
nor UO_238 (O_238,N_19800,N_19894);
or UO_239 (O_239,N_19866,N_19993);
nand UO_240 (O_240,N_19815,N_19861);
nor UO_241 (O_241,N_19917,N_19814);
or UO_242 (O_242,N_19926,N_19913);
or UO_243 (O_243,N_19989,N_19907);
nor UO_244 (O_244,N_19975,N_19996);
nor UO_245 (O_245,N_19892,N_19980);
nand UO_246 (O_246,N_19840,N_19866);
nand UO_247 (O_247,N_19969,N_19958);
xor UO_248 (O_248,N_19843,N_19933);
xor UO_249 (O_249,N_19854,N_19992);
xnor UO_250 (O_250,N_19901,N_19946);
and UO_251 (O_251,N_19820,N_19934);
xnor UO_252 (O_252,N_19922,N_19904);
nor UO_253 (O_253,N_19834,N_19854);
and UO_254 (O_254,N_19896,N_19956);
or UO_255 (O_255,N_19870,N_19958);
xor UO_256 (O_256,N_19952,N_19946);
or UO_257 (O_257,N_19930,N_19896);
or UO_258 (O_258,N_19881,N_19850);
nor UO_259 (O_259,N_19859,N_19979);
and UO_260 (O_260,N_19957,N_19873);
nand UO_261 (O_261,N_19985,N_19840);
or UO_262 (O_262,N_19978,N_19852);
and UO_263 (O_263,N_19882,N_19967);
or UO_264 (O_264,N_19904,N_19867);
nor UO_265 (O_265,N_19858,N_19869);
xnor UO_266 (O_266,N_19919,N_19868);
nor UO_267 (O_267,N_19957,N_19983);
or UO_268 (O_268,N_19848,N_19994);
nand UO_269 (O_269,N_19900,N_19908);
nor UO_270 (O_270,N_19917,N_19992);
and UO_271 (O_271,N_19879,N_19808);
nor UO_272 (O_272,N_19867,N_19911);
and UO_273 (O_273,N_19841,N_19908);
nand UO_274 (O_274,N_19848,N_19914);
nand UO_275 (O_275,N_19815,N_19977);
and UO_276 (O_276,N_19920,N_19982);
xnor UO_277 (O_277,N_19950,N_19888);
and UO_278 (O_278,N_19851,N_19857);
xor UO_279 (O_279,N_19898,N_19851);
nand UO_280 (O_280,N_19970,N_19801);
nand UO_281 (O_281,N_19870,N_19888);
nor UO_282 (O_282,N_19954,N_19879);
xnor UO_283 (O_283,N_19983,N_19804);
xor UO_284 (O_284,N_19945,N_19822);
nand UO_285 (O_285,N_19819,N_19972);
xnor UO_286 (O_286,N_19892,N_19948);
or UO_287 (O_287,N_19941,N_19934);
xor UO_288 (O_288,N_19842,N_19804);
or UO_289 (O_289,N_19980,N_19969);
nor UO_290 (O_290,N_19904,N_19806);
nand UO_291 (O_291,N_19880,N_19930);
xnor UO_292 (O_292,N_19844,N_19883);
or UO_293 (O_293,N_19924,N_19940);
nand UO_294 (O_294,N_19973,N_19954);
nor UO_295 (O_295,N_19972,N_19946);
xor UO_296 (O_296,N_19871,N_19899);
nand UO_297 (O_297,N_19928,N_19803);
nand UO_298 (O_298,N_19896,N_19939);
or UO_299 (O_299,N_19879,N_19930);
or UO_300 (O_300,N_19881,N_19867);
nand UO_301 (O_301,N_19834,N_19832);
nand UO_302 (O_302,N_19945,N_19900);
and UO_303 (O_303,N_19938,N_19917);
nand UO_304 (O_304,N_19864,N_19964);
nand UO_305 (O_305,N_19821,N_19838);
and UO_306 (O_306,N_19996,N_19902);
nand UO_307 (O_307,N_19844,N_19846);
xnor UO_308 (O_308,N_19921,N_19925);
nor UO_309 (O_309,N_19840,N_19957);
xnor UO_310 (O_310,N_19925,N_19869);
nand UO_311 (O_311,N_19833,N_19917);
xor UO_312 (O_312,N_19998,N_19950);
nor UO_313 (O_313,N_19818,N_19829);
and UO_314 (O_314,N_19849,N_19976);
xnor UO_315 (O_315,N_19870,N_19912);
nand UO_316 (O_316,N_19954,N_19853);
nand UO_317 (O_317,N_19933,N_19826);
or UO_318 (O_318,N_19930,N_19801);
nor UO_319 (O_319,N_19876,N_19906);
nor UO_320 (O_320,N_19858,N_19900);
nand UO_321 (O_321,N_19974,N_19983);
and UO_322 (O_322,N_19977,N_19807);
and UO_323 (O_323,N_19871,N_19969);
nand UO_324 (O_324,N_19937,N_19827);
xnor UO_325 (O_325,N_19895,N_19860);
nor UO_326 (O_326,N_19882,N_19958);
nor UO_327 (O_327,N_19966,N_19978);
xor UO_328 (O_328,N_19828,N_19818);
xnor UO_329 (O_329,N_19897,N_19823);
or UO_330 (O_330,N_19804,N_19936);
and UO_331 (O_331,N_19871,N_19931);
nor UO_332 (O_332,N_19811,N_19848);
nand UO_333 (O_333,N_19916,N_19817);
xnor UO_334 (O_334,N_19850,N_19874);
or UO_335 (O_335,N_19820,N_19971);
xor UO_336 (O_336,N_19965,N_19820);
nor UO_337 (O_337,N_19839,N_19898);
nor UO_338 (O_338,N_19828,N_19991);
nand UO_339 (O_339,N_19924,N_19829);
nand UO_340 (O_340,N_19895,N_19959);
nor UO_341 (O_341,N_19873,N_19889);
nand UO_342 (O_342,N_19897,N_19923);
nor UO_343 (O_343,N_19870,N_19950);
xnor UO_344 (O_344,N_19971,N_19990);
nor UO_345 (O_345,N_19990,N_19873);
xnor UO_346 (O_346,N_19955,N_19917);
and UO_347 (O_347,N_19971,N_19807);
or UO_348 (O_348,N_19832,N_19883);
nand UO_349 (O_349,N_19932,N_19910);
nor UO_350 (O_350,N_19929,N_19848);
nor UO_351 (O_351,N_19809,N_19871);
nand UO_352 (O_352,N_19818,N_19941);
nand UO_353 (O_353,N_19866,N_19805);
and UO_354 (O_354,N_19954,N_19941);
and UO_355 (O_355,N_19915,N_19944);
xnor UO_356 (O_356,N_19883,N_19949);
or UO_357 (O_357,N_19815,N_19925);
and UO_358 (O_358,N_19856,N_19848);
xnor UO_359 (O_359,N_19820,N_19915);
xor UO_360 (O_360,N_19813,N_19878);
nor UO_361 (O_361,N_19924,N_19994);
nand UO_362 (O_362,N_19803,N_19967);
xnor UO_363 (O_363,N_19959,N_19998);
xnor UO_364 (O_364,N_19994,N_19812);
xor UO_365 (O_365,N_19961,N_19971);
nand UO_366 (O_366,N_19821,N_19817);
and UO_367 (O_367,N_19910,N_19846);
xor UO_368 (O_368,N_19938,N_19895);
and UO_369 (O_369,N_19883,N_19919);
or UO_370 (O_370,N_19847,N_19886);
and UO_371 (O_371,N_19877,N_19967);
nand UO_372 (O_372,N_19977,N_19842);
or UO_373 (O_373,N_19996,N_19946);
and UO_374 (O_374,N_19819,N_19956);
xor UO_375 (O_375,N_19813,N_19917);
nand UO_376 (O_376,N_19908,N_19976);
nand UO_377 (O_377,N_19993,N_19891);
nand UO_378 (O_378,N_19813,N_19872);
xnor UO_379 (O_379,N_19845,N_19890);
nand UO_380 (O_380,N_19846,N_19835);
or UO_381 (O_381,N_19961,N_19914);
xnor UO_382 (O_382,N_19829,N_19844);
nor UO_383 (O_383,N_19953,N_19867);
nand UO_384 (O_384,N_19811,N_19964);
nand UO_385 (O_385,N_19987,N_19898);
nand UO_386 (O_386,N_19812,N_19837);
nor UO_387 (O_387,N_19991,N_19844);
and UO_388 (O_388,N_19896,N_19849);
or UO_389 (O_389,N_19931,N_19947);
or UO_390 (O_390,N_19957,N_19994);
and UO_391 (O_391,N_19898,N_19831);
xor UO_392 (O_392,N_19925,N_19953);
xnor UO_393 (O_393,N_19955,N_19876);
xnor UO_394 (O_394,N_19963,N_19916);
nor UO_395 (O_395,N_19902,N_19990);
and UO_396 (O_396,N_19891,N_19802);
and UO_397 (O_397,N_19923,N_19961);
and UO_398 (O_398,N_19980,N_19870);
nand UO_399 (O_399,N_19909,N_19841);
nand UO_400 (O_400,N_19850,N_19911);
or UO_401 (O_401,N_19847,N_19955);
nor UO_402 (O_402,N_19970,N_19893);
or UO_403 (O_403,N_19893,N_19996);
or UO_404 (O_404,N_19924,N_19895);
and UO_405 (O_405,N_19835,N_19917);
xor UO_406 (O_406,N_19863,N_19933);
and UO_407 (O_407,N_19958,N_19817);
or UO_408 (O_408,N_19800,N_19883);
xnor UO_409 (O_409,N_19940,N_19948);
or UO_410 (O_410,N_19815,N_19955);
or UO_411 (O_411,N_19884,N_19864);
and UO_412 (O_412,N_19911,N_19869);
and UO_413 (O_413,N_19961,N_19954);
or UO_414 (O_414,N_19908,N_19940);
and UO_415 (O_415,N_19899,N_19801);
nor UO_416 (O_416,N_19922,N_19897);
nor UO_417 (O_417,N_19906,N_19904);
nand UO_418 (O_418,N_19949,N_19879);
nor UO_419 (O_419,N_19909,N_19980);
and UO_420 (O_420,N_19804,N_19801);
nand UO_421 (O_421,N_19828,N_19871);
xnor UO_422 (O_422,N_19937,N_19832);
xor UO_423 (O_423,N_19859,N_19968);
xor UO_424 (O_424,N_19925,N_19899);
xor UO_425 (O_425,N_19805,N_19913);
nor UO_426 (O_426,N_19926,N_19835);
nor UO_427 (O_427,N_19802,N_19953);
xnor UO_428 (O_428,N_19938,N_19805);
and UO_429 (O_429,N_19875,N_19824);
nor UO_430 (O_430,N_19880,N_19984);
xor UO_431 (O_431,N_19919,N_19842);
or UO_432 (O_432,N_19901,N_19932);
nand UO_433 (O_433,N_19953,N_19936);
nand UO_434 (O_434,N_19803,N_19914);
nor UO_435 (O_435,N_19983,N_19822);
nand UO_436 (O_436,N_19812,N_19811);
and UO_437 (O_437,N_19994,N_19891);
and UO_438 (O_438,N_19945,N_19812);
and UO_439 (O_439,N_19905,N_19912);
and UO_440 (O_440,N_19944,N_19882);
or UO_441 (O_441,N_19888,N_19970);
nand UO_442 (O_442,N_19891,N_19921);
or UO_443 (O_443,N_19892,N_19915);
nor UO_444 (O_444,N_19829,N_19839);
and UO_445 (O_445,N_19812,N_19897);
xor UO_446 (O_446,N_19945,N_19831);
nand UO_447 (O_447,N_19913,N_19947);
xnor UO_448 (O_448,N_19918,N_19969);
xor UO_449 (O_449,N_19928,N_19892);
nor UO_450 (O_450,N_19879,N_19957);
or UO_451 (O_451,N_19909,N_19877);
nand UO_452 (O_452,N_19843,N_19910);
and UO_453 (O_453,N_19809,N_19859);
or UO_454 (O_454,N_19964,N_19842);
or UO_455 (O_455,N_19817,N_19873);
or UO_456 (O_456,N_19951,N_19888);
nor UO_457 (O_457,N_19948,N_19838);
nand UO_458 (O_458,N_19961,N_19934);
or UO_459 (O_459,N_19839,N_19995);
nand UO_460 (O_460,N_19962,N_19835);
xor UO_461 (O_461,N_19926,N_19877);
nand UO_462 (O_462,N_19953,N_19906);
or UO_463 (O_463,N_19867,N_19981);
nor UO_464 (O_464,N_19825,N_19855);
nor UO_465 (O_465,N_19935,N_19829);
nor UO_466 (O_466,N_19920,N_19870);
and UO_467 (O_467,N_19969,N_19935);
xnor UO_468 (O_468,N_19975,N_19900);
nand UO_469 (O_469,N_19991,N_19982);
and UO_470 (O_470,N_19912,N_19829);
nand UO_471 (O_471,N_19800,N_19801);
or UO_472 (O_472,N_19958,N_19865);
or UO_473 (O_473,N_19991,N_19848);
nor UO_474 (O_474,N_19995,N_19940);
nand UO_475 (O_475,N_19843,N_19814);
nand UO_476 (O_476,N_19852,N_19898);
xnor UO_477 (O_477,N_19997,N_19974);
nor UO_478 (O_478,N_19870,N_19992);
nand UO_479 (O_479,N_19912,N_19956);
nand UO_480 (O_480,N_19881,N_19813);
and UO_481 (O_481,N_19909,N_19824);
or UO_482 (O_482,N_19956,N_19967);
nor UO_483 (O_483,N_19884,N_19989);
xor UO_484 (O_484,N_19829,N_19903);
and UO_485 (O_485,N_19999,N_19896);
or UO_486 (O_486,N_19960,N_19860);
or UO_487 (O_487,N_19996,N_19911);
xor UO_488 (O_488,N_19828,N_19996);
xor UO_489 (O_489,N_19910,N_19835);
nand UO_490 (O_490,N_19976,N_19921);
nand UO_491 (O_491,N_19806,N_19998);
nand UO_492 (O_492,N_19810,N_19996);
and UO_493 (O_493,N_19989,N_19800);
xor UO_494 (O_494,N_19927,N_19972);
nor UO_495 (O_495,N_19884,N_19994);
nand UO_496 (O_496,N_19908,N_19825);
nand UO_497 (O_497,N_19853,N_19944);
nor UO_498 (O_498,N_19898,N_19836);
nand UO_499 (O_499,N_19995,N_19965);
or UO_500 (O_500,N_19807,N_19932);
xnor UO_501 (O_501,N_19987,N_19924);
nand UO_502 (O_502,N_19811,N_19997);
or UO_503 (O_503,N_19979,N_19936);
xnor UO_504 (O_504,N_19981,N_19937);
xor UO_505 (O_505,N_19865,N_19927);
nor UO_506 (O_506,N_19988,N_19931);
and UO_507 (O_507,N_19956,N_19865);
nand UO_508 (O_508,N_19876,N_19961);
and UO_509 (O_509,N_19800,N_19915);
and UO_510 (O_510,N_19895,N_19806);
xnor UO_511 (O_511,N_19897,N_19951);
nor UO_512 (O_512,N_19916,N_19845);
xor UO_513 (O_513,N_19878,N_19863);
or UO_514 (O_514,N_19837,N_19997);
nor UO_515 (O_515,N_19977,N_19863);
xnor UO_516 (O_516,N_19885,N_19874);
or UO_517 (O_517,N_19925,N_19915);
nor UO_518 (O_518,N_19861,N_19841);
and UO_519 (O_519,N_19988,N_19930);
nand UO_520 (O_520,N_19821,N_19858);
xor UO_521 (O_521,N_19818,N_19921);
and UO_522 (O_522,N_19886,N_19830);
nor UO_523 (O_523,N_19958,N_19973);
xnor UO_524 (O_524,N_19830,N_19889);
nand UO_525 (O_525,N_19944,N_19845);
nor UO_526 (O_526,N_19824,N_19842);
xor UO_527 (O_527,N_19960,N_19855);
and UO_528 (O_528,N_19820,N_19938);
nand UO_529 (O_529,N_19850,N_19841);
or UO_530 (O_530,N_19937,N_19919);
and UO_531 (O_531,N_19981,N_19881);
xor UO_532 (O_532,N_19839,N_19948);
or UO_533 (O_533,N_19892,N_19865);
nor UO_534 (O_534,N_19864,N_19819);
and UO_535 (O_535,N_19951,N_19878);
xnor UO_536 (O_536,N_19987,N_19912);
xor UO_537 (O_537,N_19869,N_19946);
or UO_538 (O_538,N_19892,N_19995);
or UO_539 (O_539,N_19994,N_19853);
nand UO_540 (O_540,N_19971,N_19871);
or UO_541 (O_541,N_19867,N_19834);
nor UO_542 (O_542,N_19928,N_19994);
nand UO_543 (O_543,N_19847,N_19986);
or UO_544 (O_544,N_19824,N_19897);
or UO_545 (O_545,N_19832,N_19946);
and UO_546 (O_546,N_19801,N_19937);
nor UO_547 (O_547,N_19841,N_19991);
or UO_548 (O_548,N_19833,N_19983);
or UO_549 (O_549,N_19962,N_19985);
and UO_550 (O_550,N_19967,N_19891);
nand UO_551 (O_551,N_19937,N_19800);
nand UO_552 (O_552,N_19955,N_19973);
and UO_553 (O_553,N_19806,N_19948);
and UO_554 (O_554,N_19849,N_19915);
or UO_555 (O_555,N_19874,N_19800);
nor UO_556 (O_556,N_19917,N_19810);
nor UO_557 (O_557,N_19978,N_19953);
or UO_558 (O_558,N_19975,N_19974);
nand UO_559 (O_559,N_19992,N_19979);
nor UO_560 (O_560,N_19925,N_19859);
nor UO_561 (O_561,N_19818,N_19885);
nand UO_562 (O_562,N_19911,N_19975);
nand UO_563 (O_563,N_19847,N_19949);
and UO_564 (O_564,N_19901,N_19867);
nor UO_565 (O_565,N_19803,N_19876);
nand UO_566 (O_566,N_19823,N_19989);
nand UO_567 (O_567,N_19934,N_19824);
and UO_568 (O_568,N_19817,N_19806);
nor UO_569 (O_569,N_19864,N_19856);
xnor UO_570 (O_570,N_19913,N_19808);
nand UO_571 (O_571,N_19961,N_19984);
and UO_572 (O_572,N_19815,N_19973);
or UO_573 (O_573,N_19976,N_19909);
nor UO_574 (O_574,N_19963,N_19996);
xnor UO_575 (O_575,N_19944,N_19896);
and UO_576 (O_576,N_19886,N_19991);
nand UO_577 (O_577,N_19876,N_19918);
xnor UO_578 (O_578,N_19844,N_19863);
nor UO_579 (O_579,N_19874,N_19820);
xor UO_580 (O_580,N_19898,N_19946);
xor UO_581 (O_581,N_19933,N_19977);
or UO_582 (O_582,N_19965,N_19930);
or UO_583 (O_583,N_19820,N_19950);
and UO_584 (O_584,N_19945,N_19881);
nor UO_585 (O_585,N_19933,N_19898);
nand UO_586 (O_586,N_19800,N_19843);
or UO_587 (O_587,N_19991,N_19806);
or UO_588 (O_588,N_19852,N_19994);
nor UO_589 (O_589,N_19961,N_19999);
nor UO_590 (O_590,N_19873,N_19993);
and UO_591 (O_591,N_19846,N_19925);
and UO_592 (O_592,N_19855,N_19845);
or UO_593 (O_593,N_19823,N_19967);
or UO_594 (O_594,N_19849,N_19834);
or UO_595 (O_595,N_19933,N_19908);
or UO_596 (O_596,N_19869,N_19902);
and UO_597 (O_597,N_19875,N_19828);
nand UO_598 (O_598,N_19831,N_19981);
or UO_599 (O_599,N_19880,N_19949);
and UO_600 (O_600,N_19976,N_19935);
nand UO_601 (O_601,N_19994,N_19834);
xnor UO_602 (O_602,N_19971,N_19914);
nor UO_603 (O_603,N_19915,N_19983);
or UO_604 (O_604,N_19811,N_19851);
or UO_605 (O_605,N_19970,N_19819);
nor UO_606 (O_606,N_19908,N_19844);
or UO_607 (O_607,N_19921,N_19860);
and UO_608 (O_608,N_19822,N_19832);
nor UO_609 (O_609,N_19989,N_19987);
xnor UO_610 (O_610,N_19953,N_19963);
nand UO_611 (O_611,N_19970,N_19802);
nor UO_612 (O_612,N_19946,N_19954);
xnor UO_613 (O_613,N_19984,N_19927);
xor UO_614 (O_614,N_19955,N_19809);
or UO_615 (O_615,N_19817,N_19978);
xnor UO_616 (O_616,N_19955,N_19808);
xnor UO_617 (O_617,N_19939,N_19898);
nor UO_618 (O_618,N_19993,N_19801);
or UO_619 (O_619,N_19820,N_19825);
or UO_620 (O_620,N_19882,N_19835);
xor UO_621 (O_621,N_19862,N_19871);
nor UO_622 (O_622,N_19816,N_19809);
xor UO_623 (O_623,N_19827,N_19855);
xor UO_624 (O_624,N_19931,N_19803);
or UO_625 (O_625,N_19948,N_19885);
xnor UO_626 (O_626,N_19830,N_19845);
or UO_627 (O_627,N_19872,N_19883);
xnor UO_628 (O_628,N_19943,N_19893);
or UO_629 (O_629,N_19827,N_19809);
nand UO_630 (O_630,N_19870,N_19873);
and UO_631 (O_631,N_19807,N_19809);
xor UO_632 (O_632,N_19976,N_19925);
nand UO_633 (O_633,N_19939,N_19908);
or UO_634 (O_634,N_19859,N_19849);
nand UO_635 (O_635,N_19867,N_19932);
nand UO_636 (O_636,N_19965,N_19816);
nor UO_637 (O_637,N_19979,N_19978);
or UO_638 (O_638,N_19964,N_19903);
nor UO_639 (O_639,N_19921,N_19808);
and UO_640 (O_640,N_19906,N_19836);
or UO_641 (O_641,N_19983,N_19969);
xnor UO_642 (O_642,N_19804,N_19970);
nand UO_643 (O_643,N_19899,N_19857);
and UO_644 (O_644,N_19902,N_19946);
xor UO_645 (O_645,N_19913,N_19868);
nand UO_646 (O_646,N_19920,N_19964);
or UO_647 (O_647,N_19896,N_19920);
and UO_648 (O_648,N_19898,N_19955);
xor UO_649 (O_649,N_19820,N_19836);
nor UO_650 (O_650,N_19854,N_19924);
nor UO_651 (O_651,N_19884,N_19939);
nor UO_652 (O_652,N_19971,N_19815);
and UO_653 (O_653,N_19954,N_19808);
and UO_654 (O_654,N_19979,N_19800);
xnor UO_655 (O_655,N_19948,N_19836);
nor UO_656 (O_656,N_19837,N_19805);
xor UO_657 (O_657,N_19962,N_19996);
nand UO_658 (O_658,N_19983,N_19920);
xor UO_659 (O_659,N_19886,N_19855);
nor UO_660 (O_660,N_19878,N_19915);
and UO_661 (O_661,N_19990,N_19840);
or UO_662 (O_662,N_19808,N_19857);
nor UO_663 (O_663,N_19977,N_19854);
or UO_664 (O_664,N_19866,N_19986);
xor UO_665 (O_665,N_19828,N_19950);
or UO_666 (O_666,N_19875,N_19976);
or UO_667 (O_667,N_19977,N_19960);
nor UO_668 (O_668,N_19914,N_19927);
or UO_669 (O_669,N_19867,N_19830);
nand UO_670 (O_670,N_19903,N_19885);
or UO_671 (O_671,N_19939,N_19849);
nor UO_672 (O_672,N_19912,N_19951);
xnor UO_673 (O_673,N_19908,N_19823);
and UO_674 (O_674,N_19911,N_19844);
xnor UO_675 (O_675,N_19895,N_19980);
xnor UO_676 (O_676,N_19835,N_19905);
nand UO_677 (O_677,N_19804,N_19867);
nand UO_678 (O_678,N_19883,N_19909);
or UO_679 (O_679,N_19879,N_19883);
or UO_680 (O_680,N_19815,N_19826);
nand UO_681 (O_681,N_19825,N_19878);
or UO_682 (O_682,N_19905,N_19847);
and UO_683 (O_683,N_19847,N_19861);
or UO_684 (O_684,N_19866,N_19987);
or UO_685 (O_685,N_19898,N_19899);
xnor UO_686 (O_686,N_19921,N_19901);
nand UO_687 (O_687,N_19818,N_19989);
nor UO_688 (O_688,N_19812,N_19943);
or UO_689 (O_689,N_19829,N_19870);
nand UO_690 (O_690,N_19941,N_19885);
or UO_691 (O_691,N_19868,N_19871);
nor UO_692 (O_692,N_19852,N_19851);
nor UO_693 (O_693,N_19932,N_19895);
and UO_694 (O_694,N_19833,N_19846);
nand UO_695 (O_695,N_19894,N_19816);
nor UO_696 (O_696,N_19833,N_19925);
nand UO_697 (O_697,N_19920,N_19926);
or UO_698 (O_698,N_19812,N_19976);
nand UO_699 (O_699,N_19843,N_19949);
and UO_700 (O_700,N_19869,N_19992);
or UO_701 (O_701,N_19894,N_19844);
nor UO_702 (O_702,N_19866,N_19968);
or UO_703 (O_703,N_19837,N_19830);
and UO_704 (O_704,N_19834,N_19899);
xnor UO_705 (O_705,N_19887,N_19901);
xnor UO_706 (O_706,N_19823,N_19862);
and UO_707 (O_707,N_19972,N_19926);
nand UO_708 (O_708,N_19964,N_19813);
nand UO_709 (O_709,N_19893,N_19962);
nor UO_710 (O_710,N_19826,N_19915);
nor UO_711 (O_711,N_19967,N_19819);
nor UO_712 (O_712,N_19809,N_19962);
or UO_713 (O_713,N_19995,N_19994);
nor UO_714 (O_714,N_19835,N_19928);
nand UO_715 (O_715,N_19926,N_19940);
nand UO_716 (O_716,N_19939,N_19874);
nand UO_717 (O_717,N_19929,N_19865);
nor UO_718 (O_718,N_19990,N_19833);
or UO_719 (O_719,N_19896,N_19873);
or UO_720 (O_720,N_19828,N_19968);
nand UO_721 (O_721,N_19843,N_19942);
nand UO_722 (O_722,N_19856,N_19873);
and UO_723 (O_723,N_19849,N_19935);
xor UO_724 (O_724,N_19974,N_19939);
and UO_725 (O_725,N_19816,N_19978);
nor UO_726 (O_726,N_19801,N_19885);
xor UO_727 (O_727,N_19866,N_19906);
and UO_728 (O_728,N_19831,N_19811);
or UO_729 (O_729,N_19950,N_19887);
nor UO_730 (O_730,N_19880,N_19944);
and UO_731 (O_731,N_19937,N_19829);
and UO_732 (O_732,N_19862,N_19817);
nor UO_733 (O_733,N_19899,N_19988);
nor UO_734 (O_734,N_19836,N_19959);
xor UO_735 (O_735,N_19961,N_19943);
nor UO_736 (O_736,N_19922,N_19980);
xor UO_737 (O_737,N_19823,N_19832);
or UO_738 (O_738,N_19915,N_19985);
and UO_739 (O_739,N_19913,N_19943);
and UO_740 (O_740,N_19844,N_19867);
or UO_741 (O_741,N_19935,N_19864);
or UO_742 (O_742,N_19870,N_19860);
and UO_743 (O_743,N_19911,N_19838);
and UO_744 (O_744,N_19991,N_19910);
nand UO_745 (O_745,N_19970,N_19965);
or UO_746 (O_746,N_19862,N_19854);
nor UO_747 (O_747,N_19919,N_19980);
nor UO_748 (O_748,N_19896,N_19905);
nand UO_749 (O_749,N_19833,N_19886);
or UO_750 (O_750,N_19837,N_19989);
and UO_751 (O_751,N_19864,N_19835);
or UO_752 (O_752,N_19928,N_19832);
and UO_753 (O_753,N_19988,N_19963);
nor UO_754 (O_754,N_19876,N_19902);
nand UO_755 (O_755,N_19994,N_19813);
or UO_756 (O_756,N_19969,N_19818);
xnor UO_757 (O_757,N_19944,N_19819);
or UO_758 (O_758,N_19810,N_19952);
and UO_759 (O_759,N_19806,N_19860);
nand UO_760 (O_760,N_19978,N_19950);
nor UO_761 (O_761,N_19842,N_19859);
or UO_762 (O_762,N_19911,N_19904);
nor UO_763 (O_763,N_19808,N_19990);
nor UO_764 (O_764,N_19917,N_19941);
xnor UO_765 (O_765,N_19882,N_19870);
and UO_766 (O_766,N_19892,N_19874);
nor UO_767 (O_767,N_19910,N_19938);
and UO_768 (O_768,N_19947,N_19892);
nor UO_769 (O_769,N_19849,N_19816);
and UO_770 (O_770,N_19864,N_19803);
xnor UO_771 (O_771,N_19937,N_19866);
or UO_772 (O_772,N_19821,N_19944);
and UO_773 (O_773,N_19821,N_19853);
or UO_774 (O_774,N_19859,N_19818);
nand UO_775 (O_775,N_19962,N_19969);
and UO_776 (O_776,N_19886,N_19884);
xnor UO_777 (O_777,N_19832,N_19997);
nor UO_778 (O_778,N_19990,N_19972);
or UO_779 (O_779,N_19810,N_19870);
nand UO_780 (O_780,N_19925,N_19816);
or UO_781 (O_781,N_19947,N_19948);
and UO_782 (O_782,N_19814,N_19809);
and UO_783 (O_783,N_19842,N_19921);
or UO_784 (O_784,N_19997,N_19856);
nor UO_785 (O_785,N_19875,N_19964);
nor UO_786 (O_786,N_19908,N_19857);
xor UO_787 (O_787,N_19846,N_19861);
or UO_788 (O_788,N_19893,N_19927);
nor UO_789 (O_789,N_19910,N_19806);
xnor UO_790 (O_790,N_19903,N_19912);
nor UO_791 (O_791,N_19813,N_19943);
or UO_792 (O_792,N_19987,N_19993);
and UO_793 (O_793,N_19828,N_19870);
and UO_794 (O_794,N_19990,N_19804);
xor UO_795 (O_795,N_19969,N_19992);
nor UO_796 (O_796,N_19892,N_19927);
and UO_797 (O_797,N_19958,N_19922);
xor UO_798 (O_798,N_19958,N_19901);
or UO_799 (O_799,N_19927,N_19806);
or UO_800 (O_800,N_19925,N_19897);
nand UO_801 (O_801,N_19974,N_19968);
or UO_802 (O_802,N_19969,N_19916);
xnor UO_803 (O_803,N_19928,N_19807);
nand UO_804 (O_804,N_19903,N_19808);
or UO_805 (O_805,N_19867,N_19897);
or UO_806 (O_806,N_19930,N_19949);
xnor UO_807 (O_807,N_19844,N_19935);
or UO_808 (O_808,N_19862,N_19913);
and UO_809 (O_809,N_19823,N_19973);
and UO_810 (O_810,N_19966,N_19887);
nand UO_811 (O_811,N_19972,N_19879);
nand UO_812 (O_812,N_19946,N_19965);
nor UO_813 (O_813,N_19875,N_19971);
or UO_814 (O_814,N_19824,N_19954);
nor UO_815 (O_815,N_19998,N_19818);
xnor UO_816 (O_816,N_19823,N_19860);
and UO_817 (O_817,N_19972,N_19810);
xor UO_818 (O_818,N_19808,N_19825);
nor UO_819 (O_819,N_19988,N_19976);
xor UO_820 (O_820,N_19993,N_19880);
nor UO_821 (O_821,N_19928,N_19979);
nor UO_822 (O_822,N_19831,N_19853);
nor UO_823 (O_823,N_19914,N_19949);
or UO_824 (O_824,N_19897,N_19873);
nand UO_825 (O_825,N_19918,N_19994);
nand UO_826 (O_826,N_19871,N_19944);
and UO_827 (O_827,N_19931,N_19884);
nor UO_828 (O_828,N_19890,N_19834);
and UO_829 (O_829,N_19963,N_19815);
nand UO_830 (O_830,N_19867,N_19997);
nor UO_831 (O_831,N_19822,N_19909);
nor UO_832 (O_832,N_19895,N_19881);
or UO_833 (O_833,N_19814,N_19857);
xor UO_834 (O_834,N_19942,N_19869);
or UO_835 (O_835,N_19961,N_19847);
nor UO_836 (O_836,N_19994,N_19946);
nor UO_837 (O_837,N_19849,N_19965);
nand UO_838 (O_838,N_19808,N_19959);
nand UO_839 (O_839,N_19963,N_19884);
and UO_840 (O_840,N_19825,N_19814);
and UO_841 (O_841,N_19952,N_19894);
or UO_842 (O_842,N_19846,N_19831);
or UO_843 (O_843,N_19854,N_19926);
xnor UO_844 (O_844,N_19901,N_19825);
or UO_845 (O_845,N_19900,N_19976);
nand UO_846 (O_846,N_19996,N_19991);
nand UO_847 (O_847,N_19819,N_19854);
or UO_848 (O_848,N_19843,N_19811);
or UO_849 (O_849,N_19939,N_19890);
nand UO_850 (O_850,N_19831,N_19895);
nand UO_851 (O_851,N_19879,N_19804);
nand UO_852 (O_852,N_19905,N_19966);
and UO_853 (O_853,N_19980,N_19885);
xnor UO_854 (O_854,N_19983,N_19996);
or UO_855 (O_855,N_19990,N_19987);
and UO_856 (O_856,N_19829,N_19896);
or UO_857 (O_857,N_19809,N_19895);
or UO_858 (O_858,N_19851,N_19936);
or UO_859 (O_859,N_19919,N_19831);
and UO_860 (O_860,N_19836,N_19946);
nand UO_861 (O_861,N_19843,N_19804);
xnor UO_862 (O_862,N_19890,N_19871);
nand UO_863 (O_863,N_19929,N_19903);
nand UO_864 (O_864,N_19915,N_19855);
nor UO_865 (O_865,N_19929,N_19888);
and UO_866 (O_866,N_19908,N_19996);
or UO_867 (O_867,N_19975,N_19831);
and UO_868 (O_868,N_19958,N_19941);
nor UO_869 (O_869,N_19984,N_19899);
or UO_870 (O_870,N_19813,N_19871);
nor UO_871 (O_871,N_19832,N_19923);
or UO_872 (O_872,N_19947,N_19925);
or UO_873 (O_873,N_19872,N_19878);
xnor UO_874 (O_874,N_19810,N_19884);
and UO_875 (O_875,N_19828,N_19842);
or UO_876 (O_876,N_19922,N_19880);
or UO_877 (O_877,N_19808,N_19838);
nand UO_878 (O_878,N_19942,N_19922);
and UO_879 (O_879,N_19831,N_19807);
xnor UO_880 (O_880,N_19822,N_19985);
or UO_881 (O_881,N_19892,N_19838);
nand UO_882 (O_882,N_19975,N_19986);
or UO_883 (O_883,N_19890,N_19977);
xnor UO_884 (O_884,N_19974,N_19857);
or UO_885 (O_885,N_19825,N_19919);
or UO_886 (O_886,N_19851,N_19814);
xnor UO_887 (O_887,N_19853,N_19981);
xnor UO_888 (O_888,N_19911,N_19895);
or UO_889 (O_889,N_19899,N_19917);
and UO_890 (O_890,N_19843,N_19947);
nand UO_891 (O_891,N_19887,N_19995);
nor UO_892 (O_892,N_19855,N_19956);
and UO_893 (O_893,N_19950,N_19953);
and UO_894 (O_894,N_19949,N_19986);
nand UO_895 (O_895,N_19824,N_19961);
and UO_896 (O_896,N_19843,N_19945);
nor UO_897 (O_897,N_19886,N_19966);
and UO_898 (O_898,N_19925,N_19920);
xnor UO_899 (O_899,N_19963,N_19919);
xnor UO_900 (O_900,N_19884,N_19986);
xnor UO_901 (O_901,N_19817,N_19999);
and UO_902 (O_902,N_19915,N_19805);
and UO_903 (O_903,N_19917,N_19986);
nand UO_904 (O_904,N_19960,N_19850);
and UO_905 (O_905,N_19860,N_19972);
nand UO_906 (O_906,N_19898,N_19947);
xnor UO_907 (O_907,N_19812,N_19919);
xnor UO_908 (O_908,N_19988,N_19957);
and UO_909 (O_909,N_19966,N_19930);
and UO_910 (O_910,N_19817,N_19872);
nor UO_911 (O_911,N_19824,N_19927);
or UO_912 (O_912,N_19902,N_19998);
or UO_913 (O_913,N_19823,N_19898);
nor UO_914 (O_914,N_19893,N_19928);
nor UO_915 (O_915,N_19936,N_19957);
or UO_916 (O_916,N_19895,N_19835);
xnor UO_917 (O_917,N_19899,N_19916);
nor UO_918 (O_918,N_19928,N_19942);
xor UO_919 (O_919,N_19991,N_19908);
and UO_920 (O_920,N_19815,N_19929);
and UO_921 (O_921,N_19867,N_19903);
or UO_922 (O_922,N_19983,N_19968);
or UO_923 (O_923,N_19929,N_19891);
xnor UO_924 (O_924,N_19877,N_19939);
nand UO_925 (O_925,N_19803,N_19949);
and UO_926 (O_926,N_19960,N_19805);
or UO_927 (O_927,N_19843,N_19901);
nor UO_928 (O_928,N_19866,N_19871);
nand UO_929 (O_929,N_19918,N_19996);
or UO_930 (O_930,N_19957,N_19809);
xnor UO_931 (O_931,N_19883,N_19822);
or UO_932 (O_932,N_19929,N_19846);
xnor UO_933 (O_933,N_19837,N_19834);
nor UO_934 (O_934,N_19850,N_19871);
and UO_935 (O_935,N_19882,N_19815);
nand UO_936 (O_936,N_19816,N_19984);
nand UO_937 (O_937,N_19969,N_19946);
or UO_938 (O_938,N_19977,N_19875);
or UO_939 (O_939,N_19972,N_19994);
nor UO_940 (O_940,N_19818,N_19919);
xnor UO_941 (O_941,N_19844,N_19927);
nand UO_942 (O_942,N_19892,N_19800);
xnor UO_943 (O_943,N_19827,N_19861);
nand UO_944 (O_944,N_19835,N_19898);
or UO_945 (O_945,N_19956,N_19906);
or UO_946 (O_946,N_19985,N_19911);
xnor UO_947 (O_947,N_19828,N_19957);
nor UO_948 (O_948,N_19996,N_19825);
nand UO_949 (O_949,N_19905,N_19981);
xor UO_950 (O_950,N_19999,N_19979);
nor UO_951 (O_951,N_19851,N_19847);
or UO_952 (O_952,N_19901,N_19842);
nand UO_953 (O_953,N_19905,N_19926);
xnor UO_954 (O_954,N_19976,N_19814);
nand UO_955 (O_955,N_19920,N_19820);
or UO_956 (O_956,N_19808,N_19818);
nand UO_957 (O_957,N_19897,N_19958);
or UO_958 (O_958,N_19919,N_19895);
or UO_959 (O_959,N_19875,N_19913);
or UO_960 (O_960,N_19895,N_19820);
and UO_961 (O_961,N_19961,N_19926);
xor UO_962 (O_962,N_19998,N_19939);
or UO_963 (O_963,N_19856,N_19850);
xor UO_964 (O_964,N_19834,N_19883);
and UO_965 (O_965,N_19844,N_19821);
nor UO_966 (O_966,N_19968,N_19975);
and UO_967 (O_967,N_19943,N_19945);
nor UO_968 (O_968,N_19905,N_19942);
and UO_969 (O_969,N_19832,N_19842);
nand UO_970 (O_970,N_19926,N_19842);
xor UO_971 (O_971,N_19870,N_19872);
or UO_972 (O_972,N_19843,N_19990);
and UO_973 (O_973,N_19947,N_19975);
nand UO_974 (O_974,N_19882,N_19863);
nand UO_975 (O_975,N_19862,N_19908);
nor UO_976 (O_976,N_19963,N_19973);
xor UO_977 (O_977,N_19955,N_19831);
or UO_978 (O_978,N_19905,N_19859);
nor UO_979 (O_979,N_19863,N_19991);
or UO_980 (O_980,N_19889,N_19967);
and UO_981 (O_981,N_19943,N_19840);
xor UO_982 (O_982,N_19917,N_19820);
xnor UO_983 (O_983,N_19857,N_19835);
and UO_984 (O_984,N_19911,N_19857);
nand UO_985 (O_985,N_19966,N_19961);
or UO_986 (O_986,N_19924,N_19866);
nand UO_987 (O_987,N_19812,N_19833);
nand UO_988 (O_988,N_19898,N_19807);
nor UO_989 (O_989,N_19802,N_19807);
nor UO_990 (O_990,N_19929,N_19875);
nor UO_991 (O_991,N_19906,N_19929);
nand UO_992 (O_992,N_19905,N_19886);
xor UO_993 (O_993,N_19916,N_19898);
or UO_994 (O_994,N_19961,N_19937);
nor UO_995 (O_995,N_19965,N_19812);
or UO_996 (O_996,N_19880,N_19894);
xor UO_997 (O_997,N_19826,N_19979);
and UO_998 (O_998,N_19986,N_19800);
xor UO_999 (O_999,N_19803,N_19892);
nor UO_1000 (O_1000,N_19832,N_19987);
and UO_1001 (O_1001,N_19821,N_19834);
nand UO_1002 (O_1002,N_19950,N_19992);
nor UO_1003 (O_1003,N_19973,N_19836);
or UO_1004 (O_1004,N_19821,N_19971);
nor UO_1005 (O_1005,N_19891,N_19915);
and UO_1006 (O_1006,N_19863,N_19907);
or UO_1007 (O_1007,N_19840,N_19979);
nor UO_1008 (O_1008,N_19890,N_19840);
or UO_1009 (O_1009,N_19841,N_19806);
and UO_1010 (O_1010,N_19987,N_19983);
and UO_1011 (O_1011,N_19926,N_19860);
or UO_1012 (O_1012,N_19869,N_19987);
and UO_1013 (O_1013,N_19800,N_19850);
or UO_1014 (O_1014,N_19986,N_19913);
and UO_1015 (O_1015,N_19916,N_19860);
or UO_1016 (O_1016,N_19917,N_19905);
nand UO_1017 (O_1017,N_19881,N_19913);
xnor UO_1018 (O_1018,N_19931,N_19976);
xor UO_1019 (O_1019,N_19986,N_19902);
or UO_1020 (O_1020,N_19928,N_19817);
xor UO_1021 (O_1021,N_19919,N_19972);
and UO_1022 (O_1022,N_19813,N_19902);
and UO_1023 (O_1023,N_19970,N_19839);
nor UO_1024 (O_1024,N_19873,N_19976);
xor UO_1025 (O_1025,N_19957,N_19827);
nand UO_1026 (O_1026,N_19840,N_19978);
or UO_1027 (O_1027,N_19876,N_19879);
nor UO_1028 (O_1028,N_19895,N_19888);
or UO_1029 (O_1029,N_19963,N_19915);
nor UO_1030 (O_1030,N_19937,N_19810);
nand UO_1031 (O_1031,N_19858,N_19968);
xor UO_1032 (O_1032,N_19883,N_19860);
nor UO_1033 (O_1033,N_19982,N_19986);
or UO_1034 (O_1034,N_19854,N_19944);
or UO_1035 (O_1035,N_19939,N_19962);
nand UO_1036 (O_1036,N_19937,N_19859);
and UO_1037 (O_1037,N_19863,N_19920);
or UO_1038 (O_1038,N_19803,N_19826);
and UO_1039 (O_1039,N_19955,N_19806);
and UO_1040 (O_1040,N_19834,N_19810);
and UO_1041 (O_1041,N_19849,N_19867);
nor UO_1042 (O_1042,N_19852,N_19806);
and UO_1043 (O_1043,N_19990,N_19911);
nand UO_1044 (O_1044,N_19800,N_19844);
or UO_1045 (O_1045,N_19872,N_19881);
xor UO_1046 (O_1046,N_19959,N_19923);
xnor UO_1047 (O_1047,N_19877,N_19895);
and UO_1048 (O_1048,N_19984,N_19805);
nand UO_1049 (O_1049,N_19838,N_19846);
or UO_1050 (O_1050,N_19947,N_19891);
xor UO_1051 (O_1051,N_19949,N_19882);
xor UO_1052 (O_1052,N_19844,N_19836);
nand UO_1053 (O_1053,N_19820,N_19897);
and UO_1054 (O_1054,N_19856,N_19902);
nand UO_1055 (O_1055,N_19927,N_19876);
nor UO_1056 (O_1056,N_19993,N_19821);
nor UO_1057 (O_1057,N_19887,N_19826);
or UO_1058 (O_1058,N_19870,N_19905);
or UO_1059 (O_1059,N_19978,N_19890);
and UO_1060 (O_1060,N_19921,N_19950);
or UO_1061 (O_1061,N_19878,N_19918);
and UO_1062 (O_1062,N_19965,N_19884);
or UO_1063 (O_1063,N_19905,N_19962);
xnor UO_1064 (O_1064,N_19916,N_19942);
or UO_1065 (O_1065,N_19885,N_19907);
nand UO_1066 (O_1066,N_19914,N_19838);
or UO_1067 (O_1067,N_19836,N_19808);
nand UO_1068 (O_1068,N_19966,N_19898);
nor UO_1069 (O_1069,N_19845,N_19978);
xor UO_1070 (O_1070,N_19843,N_19914);
xor UO_1071 (O_1071,N_19925,N_19992);
and UO_1072 (O_1072,N_19838,N_19852);
or UO_1073 (O_1073,N_19829,N_19864);
xnor UO_1074 (O_1074,N_19965,N_19862);
or UO_1075 (O_1075,N_19926,N_19947);
and UO_1076 (O_1076,N_19829,N_19834);
xnor UO_1077 (O_1077,N_19847,N_19808);
and UO_1078 (O_1078,N_19983,N_19850);
xor UO_1079 (O_1079,N_19845,N_19985);
and UO_1080 (O_1080,N_19955,N_19929);
nand UO_1081 (O_1081,N_19981,N_19852);
or UO_1082 (O_1082,N_19954,N_19821);
xnor UO_1083 (O_1083,N_19964,N_19855);
or UO_1084 (O_1084,N_19997,N_19964);
nand UO_1085 (O_1085,N_19805,N_19961);
and UO_1086 (O_1086,N_19901,N_19968);
nand UO_1087 (O_1087,N_19969,N_19975);
nand UO_1088 (O_1088,N_19850,N_19843);
and UO_1089 (O_1089,N_19804,N_19980);
xnor UO_1090 (O_1090,N_19938,N_19963);
or UO_1091 (O_1091,N_19859,N_19802);
nor UO_1092 (O_1092,N_19884,N_19845);
nor UO_1093 (O_1093,N_19802,N_19914);
nand UO_1094 (O_1094,N_19811,N_19856);
xor UO_1095 (O_1095,N_19926,N_19853);
xor UO_1096 (O_1096,N_19935,N_19961);
or UO_1097 (O_1097,N_19966,N_19841);
nand UO_1098 (O_1098,N_19804,N_19826);
and UO_1099 (O_1099,N_19873,N_19923);
nand UO_1100 (O_1100,N_19986,N_19904);
xor UO_1101 (O_1101,N_19984,N_19905);
nor UO_1102 (O_1102,N_19859,N_19836);
xnor UO_1103 (O_1103,N_19951,N_19940);
xnor UO_1104 (O_1104,N_19823,N_19900);
or UO_1105 (O_1105,N_19883,N_19833);
nand UO_1106 (O_1106,N_19866,N_19976);
or UO_1107 (O_1107,N_19914,N_19948);
and UO_1108 (O_1108,N_19924,N_19887);
nor UO_1109 (O_1109,N_19964,N_19833);
xnor UO_1110 (O_1110,N_19897,N_19972);
and UO_1111 (O_1111,N_19869,N_19829);
and UO_1112 (O_1112,N_19873,N_19894);
nor UO_1113 (O_1113,N_19914,N_19876);
nand UO_1114 (O_1114,N_19880,N_19815);
or UO_1115 (O_1115,N_19974,N_19828);
nand UO_1116 (O_1116,N_19891,N_19923);
nor UO_1117 (O_1117,N_19978,N_19894);
nand UO_1118 (O_1118,N_19814,N_19883);
nor UO_1119 (O_1119,N_19865,N_19812);
or UO_1120 (O_1120,N_19934,N_19963);
and UO_1121 (O_1121,N_19939,N_19876);
xor UO_1122 (O_1122,N_19992,N_19895);
nand UO_1123 (O_1123,N_19981,N_19971);
xnor UO_1124 (O_1124,N_19998,N_19940);
or UO_1125 (O_1125,N_19870,N_19892);
nand UO_1126 (O_1126,N_19811,N_19917);
xnor UO_1127 (O_1127,N_19961,N_19950);
and UO_1128 (O_1128,N_19967,N_19860);
nand UO_1129 (O_1129,N_19916,N_19863);
nor UO_1130 (O_1130,N_19966,N_19987);
or UO_1131 (O_1131,N_19936,N_19980);
and UO_1132 (O_1132,N_19983,N_19836);
and UO_1133 (O_1133,N_19913,N_19825);
xor UO_1134 (O_1134,N_19959,N_19893);
nor UO_1135 (O_1135,N_19935,N_19882);
xnor UO_1136 (O_1136,N_19845,N_19876);
nand UO_1137 (O_1137,N_19939,N_19838);
xor UO_1138 (O_1138,N_19817,N_19893);
xnor UO_1139 (O_1139,N_19981,N_19976);
or UO_1140 (O_1140,N_19888,N_19956);
and UO_1141 (O_1141,N_19914,N_19883);
and UO_1142 (O_1142,N_19992,N_19858);
nor UO_1143 (O_1143,N_19971,N_19870);
nor UO_1144 (O_1144,N_19841,N_19967);
or UO_1145 (O_1145,N_19830,N_19832);
and UO_1146 (O_1146,N_19954,N_19815);
xnor UO_1147 (O_1147,N_19917,N_19964);
nor UO_1148 (O_1148,N_19853,N_19982);
nand UO_1149 (O_1149,N_19856,N_19828);
and UO_1150 (O_1150,N_19962,N_19992);
or UO_1151 (O_1151,N_19805,N_19872);
xnor UO_1152 (O_1152,N_19802,N_19896);
xor UO_1153 (O_1153,N_19806,N_19818);
or UO_1154 (O_1154,N_19970,N_19896);
xnor UO_1155 (O_1155,N_19944,N_19928);
or UO_1156 (O_1156,N_19927,N_19804);
nor UO_1157 (O_1157,N_19980,N_19933);
xnor UO_1158 (O_1158,N_19820,N_19903);
xor UO_1159 (O_1159,N_19965,N_19912);
nor UO_1160 (O_1160,N_19860,N_19974);
nand UO_1161 (O_1161,N_19872,N_19818);
xor UO_1162 (O_1162,N_19971,N_19952);
and UO_1163 (O_1163,N_19974,N_19812);
and UO_1164 (O_1164,N_19815,N_19917);
and UO_1165 (O_1165,N_19857,N_19937);
and UO_1166 (O_1166,N_19870,N_19899);
or UO_1167 (O_1167,N_19876,N_19907);
nand UO_1168 (O_1168,N_19941,N_19999);
or UO_1169 (O_1169,N_19888,N_19812);
nand UO_1170 (O_1170,N_19820,N_19884);
nor UO_1171 (O_1171,N_19993,N_19953);
or UO_1172 (O_1172,N_19840,N_19852);
or UO_1173 (O_1173,N_19909,N_19912);
nand UO_1174 (O_1174,N_19953,N_19929);
nor UO_1175 (O_1175,N_19852,N_19818);
nor UO_1176 (O_1176,N_19801,N_19841);
and UO_1177 (O_1177,N_19989,N_19955);
nand UO_1178 (O_1178,N_19833,N_19996);
xnor UO_1179 (O_1179,N_19928,N_19902);
xnor UO_1180 (O_1180,N_19975,N_19922);
nand UO_1181 (O_1181,N_19842,N_19853);
xnor UO_1182 (O_1182,N_19907,N_19911);
or UO_1183 (O_1183,N_19985,N_19850);
nor UO_1184 (O_1184,N_19972,N_19883);
nand UO_1185 (O_1185,N_19806,N_19984);
and UO_1186 (O_1186,N_19900,N_19958);
xnor UO_1187 (O_1187,N_19965,N_19960);
or UO_1188 (O_1188,N_19863,N_19813);
nand UO_1189 (O_1189,N_19816,N_19872);
nand UO_1190 (O_1190,N_19858,N_19912);
nor UO_1191 (O_1191,N_19979,N_19962);
and UO_1192 (O_1192,N_19803,N_19944);
or UO_1193 (O_1193,N_19979,N_19907);
xor UO_1194 (O_1194,N_19944,N_19926);
nand UO_1195 (O_1195,N_19830,N_19942);
and UO_1196 (O_1196,N_19894,N_19857);
or UO_1197 (O_1197,N_19862,N_19933);
xor UO_1198 (O_1198,N_19885,N_19949);
nor UO_1199 (O_1199,N_19820,N_19935);
xor UO_1200 (O_1200,N_19911,N_19921);
or UO_1201 (O_1201,N_19834,N_19969);
nor UO_1202 (O_1202,N_19956,N_19911);
xor UO_1203 (O_1203,N_19922,N_19969);
nor UO_1204 (O_1204,N_19947,N_19903);
and UO_1205 (O_1205,N_19914,N_19892);
nor UO_1206 (O_1206,N_19998,N_19888);
and UO_1207 (O_1207,N_19993,N_19877);
nor UO_1208 (O_1208,N_19992,N_19920);
nand UO_1209 (O_1209,N_19806,N_19885);
and UO_1210 (O_1210,N_19943,N_19853);
xor UO_1211 (O_1211,N_19977,N_19886);
nor UO_1212 (O_1212,N_19809,N_19999);
nor UO_1213 (O_1213,N_19935,N_19977);
and UO_1214 (O_1214,N_19867,N_19819);
nor UO_1215 (O_1215,N_19998,N_19835);
and UO_1216 (O_1216,N_19996,N_19997);
xnor UO_1217 (O_1217,N_19881,N_19883);
nand UO_1218 (O_1218,N_19878,N_19849);
nor UO_1219 (O_1219,N_19966,N_19927);
and UO_1220 (O_1220,N_19844,N_19827);
and UO_1221 (O_1221,N_19816,N_19964);
xnor UO_1222 (O_1222,N_19987,N_19868);
nand UO_1223 (O_1223,N_19852,N_19979);
nor UO_1224 (O_1224,N_19976,N_19859);
nand UO_1225 (O_1225,N_19814,N_19880);
or UO_1226 (O_1226,N_19825,N_19990);
xnor UO_1227 (O_1227,N_19958,N_19968);
nand UO_1228 (O_1228,N_19869,N_19949);
nand UO_1229 (O_1229,N_19982,N_19834);
nor UO_1230 (O_1230,N_19909,N_19858);
or UO_1231 (O_1231,N_19914,N_19806);
and UO_1232 (O_1232,N_19968,N_19879);
and UO_1233 (O_1233,N_19972,N_19868);
xor UO_1234 (O_1234,N_19984,N_19870);
xnor UO_1235 (O_1235,N_19978,N_19813);
nand UO_1236 (O_1236,N_19957,N_19917);
or UO_1237 (O_1237,N_19901,N_19964);
or UO_1238 (O_1238,N_19866,N_19843);
or UO_1239 (O_1239,N_19980,N_19961);
nor UO_1240 (O_1240,N_19828,N_19890);
or UO_1241 (O_1241,N_19804,N_19875);
or UO_1242 (O_1242,N_19800,N_19831);
nor UO_1243 (O_1243,N_19935,N_19985);
or UO_1244 (O_1244,N_19821,N_19987);
and UO_1245 (O_1245,N_19921,N_19917);
or UO_1246 (O_1246,N_19997,N_19850);
and UO_1247 (O_1247,N_19984,N_19802);
nand UO_1248 (O_1248,N_19874,N_19805);
and UO_1249 (O_1249,N_19802,N_19938);
nor UO_1250 (O_1250,N_19943,N_19873);
or UO_1251 (O_1251,N_19821,N_19812);
nor UO_1252 (O_1252,N_19963,N_19908);
or UO_1253 (O_1253,N_19963,N_19950);
nor UO_1254 (O_1254,N_19907,N_19811);
and UO_1255 (O_1255,N_19919,N_19925);
nand UO_1256 (O_1256,N_19999,N_19836);
nor UO_1257 (O_1257,N_19842,N_19814);
nor UO_1258 (O_1258,N_19923,N_19993);
or UO_1259 (O_1259,N_19958,N_19848);
or UO_1260 (O_1260,N_19995,N_19808);
or UO_1261 (O_1261,N_19800,N_19963);
or UO_1262 (O_1262,N_19873,N_19800);
and UO_1263 (O_1263,N_19841,N_19929);
nand UO_1264 (O_1264,N_19890,N_19865);
or UO_1265 (O_1265,N_19860,N_19920);
and UO_1266 (O_1266,N_19850,N_19807);
or UO_1267 (O_1267,N_19839,N_19897);
xnor UO_1268 (O_1268,N_19800,N_19910);
nor UO_1269 (O_1269,N_19829,N_19850);
and UO_1270 (O_1270,N_19801,N_19932);
or UO_1271 (O_1271,N_19876,N_19912);
or UO_1272 (O_1272,N_19934,N_19990);
and UO_1273 (O_1273,N_19816,N_19974);
nand UO_1274 (O_1274,N_19871,N_19851);
nand UO_1275 (O_1275,N_19964,N_19819);
xor UO_1276 (O_1276,N_19809,N_19948);
and UO_1277 (O_1277,N_19882,N_19984);
or UO_1278 (O_1278,N_19825,N_19980);
nor UO_1279 (O_1279,N_19886,N_19982);
or UO_1280 (O_1280,N_19897,N_19968);
xor UO_1281 (O_1281,N_19942,N_19972);
xor UO_1282 (O_1282,N_19870,N_19954);
nand UO_1283 (O_1283,N_19944,N_19889);
or UO_1284 (O_1284,N_19995,N_19862);
nand UO_1285 (O_1285,N_19805,N_19836);
or UO_1286 (O_1286,N_19804,N_19898);
and UO_1287 (O_1287,N_19803,N_19906);
nand UO_1288 (O_1288,N_19950,N_19946);
nand UO_1289 (O_1289,N_19982,N_19895);
nor UO_1290 (O_1290,N_19949,N_19878);
xnor UO_1291 (O_1291,N_19953,N_19948);
xor UO_1292 (O_1292,N_19934,N_19883);
xnor UO_1293 (O_1293,N_19826,N_19975);
and UO_1294 (O_1294,N_19971,N_19829);
nor UO_1295 (O_1295,N_19834,N_19875);
nand UO_1296 (O_1296,N_19913,N_19923);
xnor UO_1297 (O_1297,N_19903,N_19824);
nand UO_1298 (O_1298,N_19848,N_19829);
or UO_1299 (O_1299,N_19825,N_19949);
xnor UO_1300 (O_1300,N_19826,N_19844);
nor UO_1301 (O_1301,N_19883,N_19880);
xnor UO_1302 (O_1302,N_19897,N_19971);
nand UO_1303 (O_1303,N_19845,N_19806);
xor UO_1304 (O_1304,N_19847,N_19948);
nand UO_1305 (O_1305,N_19891,N_19982);
or UO_1306 (O_1306,N_19837,N_19875);
xor UO_1307 (O_1307,N_19991,N_19820);
or UO_1308 (O_1308,N_19967,N_19878);
xor UO_1309 (O_1309,N_19875,N_19960);
xnor UO_1310 (O_1310,N_19932,N_19850);
or UO_1311 (O_1311,N_19936,N_19928);
and UO_1312 (O_1312,N_19966,N_19925);
xnor UO_1313 (O_1313,N_19952,N_19889);
or UO_1314 (O_1314,N_19913,N_19874);
or UO_1315 (O_1315,N_19980,N_19902);
nor UO_1316 (O_1316,N_19948,N_19884);
or UO_1317 (O_1317,N_19984,N_19943);
or UO_1318 (O_1318,N_19811,N_19989);
nor UO_1319 (O_1319,N_19890,N_19807);
nand UO_1320 (O_1320,N_19976,N_19855);
xnor UO_1321 (O_1321,N_19814,N_19824);
nand UO_1322 (O_1322,N_19984,N_19866);
and UO_1323 (O_1323,N_19823,N_19820);
or UO_1324 (O_1324,N_19897,N_19967);
or UO_1325 (O_1325,N_19968,N_19821);
xnor UO_1326 (O_1326,N_19874,N_19980);
xor UO_1327 (O_1327,N_19886,N_19962);
xor UO_1328 (O_1328,N_19863,N_19945);
or UO_1329 (O_1329,N_19918,N_19954);
nor UO_1330 (O_1330,N_19861,N_19947);
nor UO_1331 (O_1331,N_19956,N_19991);
xnor UO_1332 (O_1332,N_19880,N_19988);
nand UO_1333 (O_1333,N_19902,N_19842);
xor UO_1334 (O_1334,N_19898,N_19919);
xor UO_1335 (O_1335,N_19832,N_19913);
xnor UO_1336 (O_1336,N_19850,N_19987);
and UO_1337 (O_1337,N_19926,N_19840);
nor UO_1338 (O_1338,N_19813,N_19987);
nor UO_1339 (O_1339,N_19881,N_19886);
xor UO_1340 (O_1340,N_19965,N_19876);
or UO_1341 (O_1341,N_19880,N_19879);
nand UO_1342 (O_1342,N_19901,N_19803);
nand UO_1343 (O_1343,N_19952,N_19879);
and UO_1344 (O_1344,N_19881,N_19985);
and UO_1345 (O_1345,N_19883,N_19967);
nand UO_1346 (O_1346,N_19874,N_19801);
nor UO_1347 (O_1347,N_19843,N_19879);
and UO_1348 (O_1348,N_19942,N_19802);
xnor UO_1349 (O_1349,N_19904,N_19825);
xor UO_1350 (O_1350,N_19982,N_19879);
or UO_1351 (O_1351,N_19801,N_19822);
or UO_1352 (O_1352,N_19996,N_19949);
nand UO_1353 (O_1353,N_19877,N_19850);
nor UO_1354 (O_1354,N_19993,N_19948);
xnor UO_1355 (O_1355,N_19848,N_19851);
xor UO_1356 (O_1356,N_19848,N_19838);
or UO_1357 (O_1357,N_19830,N_19914);
nand UO_1358 (O_1358,N_19851,N_19925);
or UO_1359 (O_1359,N_19985,N_19934);
or UO_1360 (O_1360,N_19818,N_19979);
xor UO_1361 (O_1361,N_19904,N_19883);
and UO_1362 (O_1362,N_19970,N_19870);
nor UO_1363 (O_1363,N_19804,N_19899);
or UO_1364 (O_1364,N_19855,N_19961);
and UO_1365 (O_1365,N_19965,N_19878);
nand UO_1366 (O_1366,N_19868,N_19974);
nor UO_1367 (O_1367,N_19971,N_19972);
xnor UO_1368 (O_1368,N_19804,N_19825);
xor UO_1369 (O_1369,N_19905,N_19907);
nand UO_1370 (O_1370,N_19886,N_19933);
nor UO_1371 (O_1371,N_19917,N_19996);
xnor UO_1372 (O_1372,N_19965,N_19905);
nor UO_1373 (O_1373,N_19871,N_19802);
nand UO_1374 (O_1374,N_19954,N_19999);
and UO_1375 (O_1375,N_19879,N_19865);
nand UO_1376 (O_1376,N_19971,N_19865);
nor UO_1377 (O_1377,N_19824,N_19826);
and UO_1378 (O_1378,N_19879,N_19814);
xnor UO_1379 (O_1379,N_19979,N_19801);
nand UO_1380 (O_1380,N_19881,N_19890);
and UO_1381 (O_1381,N_19862,N_19943);
or UO_1382 (O_1382,N_19809,N_19960);
nor UO_1383 (O_1383,N_19929,N_19864);
nand UO_1384 (O_1384,N_19809,N_19935);
nand UO_1385 (O_1385,N_19994,N_19992);
and UO_1386 (O_1386,N_19983,N_19890);
nor UO_1387 (O_1387,N_19895,N_19885);
or UO_1388 (O_1388,N_19892,N_19942);
nor UO_1389 (O_1389,N_19900,N_19853);
nand UO_1390 (O_1390,N_19803,N_19915);
nand UO_1391 (O_1391,N_19895,N_19904);
or UO_1392 (O_1392,N_19822,N_19814);
xor UO_1393 (O_1393,N_19850,N_19965);
or UO_1394 (O_1394,N_19838,N_19977);
nand UO_1395 (O_1395,N_19903,N_19946);
and UO_1396 (O_1396,N_19968,N_19946);
and UO_1397 (O_1397,N_19961,N_19815);
or UO_1398 (O_1398,N_19944,N_19931);
nor UO_1399 (O_1399,N_19971,N_19964);
and UO_1400 (O_1400,N_19877,N_19857);
or UO_1401 (O_1401,N_19994,N_19899);
xor UO_1402 (O_1402,N_19871,N_19829);
xor UO_1403 (O_1403,N_19964,N_19844);
or UO_1404 (O_1404,N_19886,N_19811);
or UO_1405 (O_1405,N_19959,N_19982);
nand UO_1406 (O_1406,N_19863,N_19861);
and UO_1407 (O_1407,N_19874,N_19839);
or UO_1408 (O_1408,N_19986,N_19909);
or UO_1409 (O_1409,N_19855,N_19859);
nor UO_1410 (O_1410,N_19858,N_19877);
and UO_1411 (O_1411,N_19805,N_19815);
nor UO_1412 (O_1412,N_19916,N_19935);
or UO_1413 (O_1413,N_19984,N_19974);
nand UO_1414 (O_1414,N_19997,N_19985);
xor UO_1415 (O_1415,N_19933,N_19928);
and UO_1416 (O_1416,N_19978,N_19801);
or UO_1417 (O_1417,N_19954,N_19939);
nand UO_1418 (O_1418,N_19846,N_19862);
and UO_1419 (O_1419,N_19959,N_19844);
and UO_1420 (O_1420,N_19923,N_19867);
nor UO_1421 (O_1421,N_19950,N_19867);
xnor UO_1422 (O_1422,N_19822,N_19910);
and UO_1423 (O_1423,N_19991,N_19916);
xor UO_1424 (O_1424,N_19845,N_19952);
xor UO_1425 (O_1425,N_19905,N_19940);
or UO_1426 (O_1426,N_19800,N_19806);
or UO_1427 (O_1427,N_19919,N_19969);
and UO_1428 (O_1428,N_19997,N_19986);
and UO_1429 (O_1429,N_19983,N_19821);
xnor UO_1430 (O_1430,N_19969,N_19813);
nor UO_1431 (O_1431,N_19914,N_19908);
or UO_1432 (O_1432,N_19879,N_19917);
nand UO_1433 (O_1433,N_19891,N_19811);
nor UO_1434 (O_1434,N_19909,N_19900);
nor UO_1435 (O_1435,N_19822,N_19968);
nor UO_1436 (O_1436,N_19889,N_19993);
and UO_1437 (O_1437,N_19973,N_19951);
and UO_1438 (O_1438,N_19827,N_19822);
nor UO_1439 (O_1439,N_19887,N_19977);
or UO_1440 (O_1440,N_19879,N_19838);
nor UO_1441 (O_1441,N_19830,N_19959);
or UO_1442 (O_1442,N_19965,N_19828);
nand UO_1443 (O_1443,N_19865,N_19839);
nor UO_1444 (O_1444,N_19922,N_19861);
xor UO_1445 (O_1445,N_19933,N_19929);
nand UO_1446 (O_1446,N_19813,N_19800);
xnor UO_1447 (O_1447,N_19900,N_19841);
nor UO_1448 (O_1448,N_19933,N_19828);
nor UO_1449 (O_1449,N_19846,N_19950);
xor UO_1450 (O_1450,N_19856,N_19956);
nand UO_1451 (O_1451,N_19822,N_19911);
xnor UO_1452 (O_1452,N_19920,N_19922);
nand UO_1453 (O_1453,N_19947,N_19814);
nor UO_1454 (O_1454,N_19932,N_19904);
nand UO_1455 (O_1455,N_19825,N_19862);
nor UO_1456 (O_1456,N_19912,N_19955);
and UO_1457 (O_1457,N_19968,N_19990);
or UO_1458 (O_1458,N_19834,N_19852);
nand UO_1459 (O_1459,N_19929,N_19884);
nand UO_1460 (O_1460,N_19984,N_19801);
nand UO_1461 (O_1461,N_19870,N_19854);
nor UO_1462 (O_1462,N_19844,N_19835);
and UO_1463 (O_1463,N_19991,N_19952);
or UO_1464 (O_1464,N_19938,N_19931);
nand UO_1465 (O_1465,N_19961,N_19859);
and UO_1466 (O_1466,N_19988,N_19942);
nor UO_1467 (O_1467,N_19833,N_19820);
xnor UO_1468 (O_1468,N_19932,N_19896);
nand UO_1469 (O_1469,N_19821,N_19913);
nor UO_1470 (O_1470,N_19892,N_19885);
xnor UO_1471 (O_1471,N_19973,N_19897);
nand UO_1472 (O_1472,N_19936,N_19808);
nor UO_1473 (O_1473,N_19846,N_19915);
xnor UO_1474 (O_1474,N_19971,N_19809);
or UO_1475 (O_1475,N_19830,N_19968);
and UO_1476 (O_1476,N_19823,N_19815);
and UO_1477 (O_1477,N_19901,N_19845);
nand UO_1478 (O_1478,N_19895,N_19951);
or UO_1479 (O_1479,N_19936,N_19805);
and UO_1480 (O_1480,N_19994,N_19880);
nand UO_1481 (O_1481,N_19926,N_19870);
xnor UO_1482 (O_1482,N_19812,N_19993);
nand UO_1483 (O_1483,N_19863,N_19897);
xor UO_1484 (O_1484,N_19830,N_19969);
and UO_1485 (O_1485,N_19932,N_19855);
nor UO_1486 (O_1486,N_19812,N_19955);
xor UO_1487 (O_1487,N_19894,N_19823);
or UO_1488 (O_1488,N_19819,N_19856);
and UO_1489 (O_1489,N_19936,N_19871);
nor UO_1490 (O_1490,N_19800,N_19862);
nor UO_1491 (O_1491,N_19946,N_19853);
xnor UO_1492 (O_1492,N_19821,N_19950);
nor UO_1493 (O_1493,N_19953,N_19996);
and UO_1494 (O_1494,N_19940,N_19813);
and UO_1495 (O_1495,N_19853,N_19938);
or UO_1496 (O_1496,N_19895,N_19903);
xnor UO_1497 (O_1497,N_19914,N_19857);
nor UO_1498 (O_1498,N_19805,N_19954);
and UO_1499 (O_1499,N_19840,N_19945);
and UO_1500 (O_1500,N_19825,N_19989);
and UO_1501 (O_1501,N_19947,N_19878);
nand UO_1502 (O_1502,N_19817,N_19975);
xnor UO_1503 (O_1503,N_19875,N_19943);
and UO_1504 (O_1504,N_19812,N_19951);
xor UO_1505 (O_1505,N_19862,N_19992);
and UO_1506 (O_1506,N_19929,N_19821);
nand UO_1507 (O_1507,N_19834,N_19919);
nor UO_1508 (O_1508,N_19977,N_19819);
xnor UO_1509 (O_1509,N_19882,N_19822);
and UO_1510 (O_1510,N_19910,N_19987);
nand UO_1511 (O_1511,N_19833,N_19853);
and UO_1512 (O_1512,N_19950,N_19941);
or UO_1513 (O_1513,N_19880,N_19948);
xor UO_1514 (O_1514,N_19875,N_19920);
nand UO_1515 (O_1515,N_19985,N_19949);
or UO_1516 (O_1516,N_19970,N_19875);
xor UO_1517 (O_1517,N_19931,N_19863);
nand UO_1518 (O_1518,N_19831,N_19960);
xnor UO_1519 (O_1519,N_19944,N_19919);
nand UO_1520 (O_1520,N_19800,N_19857);
nand UO_1521 (O_1521,N_19994,N_19921);
nand UO_1522 (O_1522,N_19988,N_19822);
xor UO_1523 (O_1523,N_19812,N_19963);
nand UO_1524 (O_1524,N_19958,N_19827);
and UO_1525 (O_1525,N_19966,N_19984);
or UO_1526 (O_1526,N_19936,N_19916);
xor UO_1527 (O_1527,N_19828,N_19804);
or UO_1528 (O_1528,N_19927,N_19819);
or UO_1529 (O_1529,N_19970,N_19806);
nor UO_1530 (O_1530,N_19900,N_19833);
nor UO_1531 (O_1531,N_19806,N_19824);
xnor UO_1532 (O_1532,N_19963,N_19913);
nor UO_1533 (O_1533,N_19892,N_19810);
and UO_1534 (O_1534,N_19988,N_19868);
or UO_1535 (O_1535,N_19973,N_19860);
and UO_1536 (O_1536,N_19930,N_19932);
and UO_1537 (O_1537,N_19993,N_19864);
nor UO_1538 (O_1538,N_19960,N_19895);
or UO_1539 (O_1539,N_19867,N_19933);
and UO_1540 (O_1540,N_19841,N_19973);
nor UO_1541 (O_1541,N_19841,N_19896);
nand UO_1542 (O_1542,N_19986,N_19839);
nand UO_1543 (O_1543,N_19899,N_19828);
or UO_1544 (O_1544,N_19930,N_19812);
nor UO_1545 (O_1545,N_19900,N_19991);
and UO_1546 (O_1546,N_19802,N_19928);
nor UO_1547 (O_1547,N_19961,N_19917);
nor UO_1548 (O_1548,N_19827,N_19828);
or UO_1549 (O_1549,N_19970,N_19882);
nor UO_1550 (O_1550,N_19895,N_19808);
xnor UO_1551 (O_1551,N_19824,N_19991);
and UO_1552 (O_1552,N_19891,N_19867);
xnor UO_1553 (O_1553,N_19857,N_19953);
and UO_1554 (O_1554,N_19891,N_19807);
or UO_1555 (O_1555,N_19952,N_19828);
or UO_1556 (O_1556,N_19964,N_19831);
nand UO_1557 (O_1557,N_19833,N_19903);
nand UO_1558 (O_1558,N_19878,N_19968);
and UO_1559 (O_1559,N_19895,N_19841);
or UO_1560 (O_1560,N_19955,N_19938);
xnor UO_1561 (O_1561,N_19839,N_19812);
or UO_1562 (O_1562,N_19970,N_19927);
nor UO_1563 (O_1563,N_19899,N_19934);
nor UO_1564 (O_1564,N_19975,N_19894);
nand UO_1565 (O_1565,N_19943,N_19864);
xnor UO_1566 (O_1566,N_19836,N_19807);
and UO_1567 (O_1567,N_19853,N_19914);
nor UO_1568 (O_1568,N_19860,N_19922);
and UO_1569 (O_1569,N_19949,N_19822);
xor UO_1570 (O_1570,N_19868,N_19969);
or UO_1571 (O_1571,N_19944,N_19836);
xor UO_1572 (O_1572,N_19963,N_19939);
nor UO_1573 (O_1573,N_19814,N_19885);
or UO_1574 (O_1574,N_19875,N_19807);
and UO_1575 (O_1575,N_19920,N_19956);
and UO_1576 (O_1576,N_19899,N_19946);
xor UO_1577 (O_1577,N_19951,N_19916);
or UO_1578 (O_1578,N_19975,N_19858);
or UO_1579 (O_1579,N_19888,N_19935);
xor UO_1580 (O_1580,N_19889,N_19860);
xnor UO_1581 (O_1581,N_19943,N_19925);
xnor UO_1582 (O_1582,N_19810,N_19844);
and UO_1583 (O_1583,N_19809,N_19834);
and UO_1584 (O_1584,N_19993,N_19837);
or UO_1585 (O_1585,N_19852,N_19989);
nand UO_1586 (O_1586,N_19893,N_19855);
nand UO_1587 (O_1587,N_19928,N_19958);
nor UO_1588 (O_1588,N_19978,N_19988);
and UO_1589 (O_1589,N_19935,N_19800);
or UO_1590 (O_1590,N_19808,N_19866);
xor UO_1591 (O_1591,N_19859,N_19819);
xor UO_1592 (O_1592,N_19854,N_19981);
or UO_1593 (O_1593,N_19828,N_19863);
and UO_1594 (O_1594,N_19835,N_19985);
nor UO_1595 (O_1595,N_19923,N_19998);
nand UO_1596 (O_1596,N_19837,N_19944);
nor UO_1597 (O_1597,N_19938,N_19929);
or UO_1598 (O_1598,N_19822,N_19826);
and UO_1599 (O_1599,N_19866,N_19952);
nand UO_1600 (O_1600,N_19808,N_19824);
and UO_1601 (O_1601,N_19924,N_19882);
or UO_1602 (O_1602,N_19961,N_19975);
or UO_1603 (O_1603,N_19893,N_19801);
and UO_1604 (O_1604,N_19968,N_19871);
nand UO_1605 (O_1605,N_19829,N_19835);
nor UO_1606 (O_1606,N_19963,N_19978);
xor UO_1607 (O_1607,N_19942,N_19962);
and UO_1608 (O_1608,N_19988,N_19909);
nand UO_1609 (O_1609,N_19907,N_19838);
and UO_1610 (O_1610,N_19833,N_19942);
nand UO_1611 (O_1611,N_19806,N_19920);
xor UO_1612 (O_1612,N_19823,N_19822);
nor UO_1613 (O_1613,N_19888,N_19932);
and UO_1614 (O_1614,N_19925,N_19889);
xnor UO_1615 (O_1615,N_19993,N_19939);
nand UO_1616 (O_1616,N_19958,N_19934);
nor UO_1617 (O_1617,N_19812,N_19909);
xor UO_1618 (O_1618,N_19817,N_19926);
nor UO_1619 (O_1619,N_19860,N_19844);
or UO_1620 (O_1620,N_19945,N_19967);
xnor UO_1621 (O_1621,N_19869,N_19843);
and UO_1622 (O_1622,N_19983,N_19923);
nor UO_1623 (O_1623,N_19843,N_19864);
and UO_1624 (O_1624,N_19922,N_19944);
nand UO_1625 (O_1625,N_19981,N_19828);
nand UO_1626 (O_1626,N_19956,N_19902);
and UO_1627 (O_1627,N_19951,N_19931);
or UO_1628 (O_1628,N_19880,N_19812);
or UO_1629 (O_1629,N_19993,N_19827);
xor UO_1630 (O_1630,N_19994,N_19958);
or UO_1631 (O_1631,N_19995,N_19997);
nand UO_1632 (O_1632,N_19859,N_19964);
nand UO_1633 (O_1633,N_19876,N_19880);
xnor UO_1634 (O_1634,N_19874,N_19899);
and UO_1635 (O_1635,N_19946,N_19849);
nor UO_1636 (O_1636,N_19985,N_19924);
or UO_1637 (O_1637,N_19911,N_19919);
xor UO_1638 (O_1638,N_19961,N_19827);
nand UO_1639 (O_1639,N_19950,N_19818);
or UO_1640 (O_1640,N_19819,N_19924);
or UO_1641 (O_1641,N_19967,N_19810);
nor UO_1642 (O_1642,N_19937,N_19904);
nand UO_1643 (O_1643,N_19834,N_19909);
or UO_1644 (O_1644,N_19807,N_19863);
or UO_1645 (O_1645,N_19975,N_19888);
and UO_1646 (O_1646,N_19828,N_19850);
and UO_1647 (O_1647,N_19945,N_19974);
nand UO_1648 (O_1648,N_19842,N_19929);
xor UO_1649 (O_1649,N_19871,N_19817);
xor UO_1650 (O_1650,N_19820,N_19829);
or UO_1651 (O_1651,N_19886,N_19853);
xor UO_1652 (O_1652,N_19871,N_19811);
and UO_1653 (O_1653,N_19986,N_19858);
nand UO_1654 (O_1654,N_19943,N_19996);
nand UO_1655 (O_1655,N_19998,N_19949);
nand UO_1656 (O_1656,N_19964,N_19962);
nand UO_1657 (O_1657,N_19897,N_19831);
and UO_1658 (O_1658,N_19992,N_19960);
and UO_1659 (O_1659,N_19909,N_19881);
nand UO_1660 (O_1660,N_19891,N_19972);
nor UO_1661 (O_1661,N_19856,N_19887);
or UO_1662 (O_1662,N_19893,N_19823);
nor UO_1663 (O_1663,N_19811,N_19968);
nor UO_1664 (O_1664,N_19988,N_19863);
nand UO_1665 (O_1665,N_19991,N_19851);
nand UO_1666 (O_1666,N_19835,N_19897);
nand UO_1667 (O_1667,N_19920,N_19955);
nand UO_1668 (O_1668,N_19978,N_19947);
or UO_1669 (O_1669,N_19870,N_19965);
nor UO_1670 (O_1670,N_19870,N_19995);
and UO_1671 (O_1671,N_19922,N_19908);
nand UO_1672 (O_1672,N_19891,N_19826);
or UO_1673 (O_1673,N_19940,N_19890);
or UO_1674 (O_1674,N_19891,N_19904);
xor UO_1675 (O_1675,N_19984,N_19800);
xnor UO_1676 (O_1676,N_19965,N_19874);
and UO_1677 (O_1677,N_19979,N_19989);
nor UO_1678 (O_1678,N_19922,N_19833);
nor UO_1679 (O_1679,N_19808,N_19982);
nand UO_1680 (O_1680,N_19961,N_19929);
and UO_1681 (O_1681,N_19921,N_19963);
nand UO_1682 (O_1682,N_19843,N_19841);
nor UO_1683 (O_1683,N_19915,N_19806);
or UO_1684 (O_1684,N_19977,N_19965);
nor UO_1685 (O_1685,N_19984,N_19935);
or UO_1686 (O_1686,N_19980,N_19965);
nor UO_1687 (O_1687,N_19901,N_19920);
xnor UO_1688 (O_1688,N_19850,N_19820);
nor UO_1689 (O_1689,N_19907,N_19839);
nor UO_1690 (O_1690,N_19929,N_19890);
nor UO_1691 (O_1691,N_19881,N_19800);
and UO_1692 (O_1692,N_19945,N_19832);
and UO_1693 (O_1693,N_19894,N_19811);
nand UO_1694 (O_1694,N_19916,N_19855);
xor UO_1695 (O_1695,N_19843,N_19904);
nor UO_1696 (O_1696,N_19810,N_19858);
nor UO_1697 (O_1697,N_19816,N_19903);
nor UO_1698 (O_1698,N_19814,N_19942);
and UO_1699 (O_1699,N_19998,N_19913);
nand UO_1700 (O_1700,N_19835,N_19870);
and UO_1701 (O_1701,N_19946,N_19814);
xnor UO_1702 (O_1702,N_19831,N_19946);
and UO_1703 (O_1703,N_19929,N_19981);
nor UO_1704 (O_1704,N_19816,N_19828);
nand UO_1705 (O_1705,N_19980,N_19962);
or UO_1706 (O_1706,N_19921,N_19964);
nor UO_1707 (O_1707,N_19825,N_19935);
nand UO_1708 (O_1708,N_19944,N_19847);
nor UO_1709 (O_1709,N_19974,N_19824);
nand UO_1710 (O_1710,N_19873,N_19825);
nor UO_1711 (O_1711,N_19854,N_19928);
or UO_1712 (O_1712,N_19842,N_19890);
xnor UO_1713 (O_1713,N_19881,N_19896);
nand UO_1714 (O_1714,N_19881,N_19940);
nor UO_1715 (O_1715,N_19854,N_19800);
nor UO_1716 (O_1716,N_19945,N_19934);
nor UO_1717 (O_1717,N_19988,N_19977);
nand UO_1718 (O_1718,N_19929,N_19982);
and UO_1719 (O_1719,N_19885,N_19906);
nor UO_1720 (O_1720,N_19970,N_19921);
nand UO_1721 (O_1721,N_19973,N_19919);
and UO_1722 (O_1722,N_19997,N_19929);
or UO_1723 (O_1723,N_19973,N_19949);
nor UO_1724 (O_1724,N_19936,N_19933);
nor UO_1725 (O_1725,N_19845,N_19879);
or UO_1726 (O_1726,N_19849,N_19887);
xor UO_1727 (O_1727,N_19911,N_19892);
and UO_1728 (O_1728,N_19831,N_19924);
and UO_1729 (O_1729,N_19802,N_19998);
or UO_1730 (O_1730,N_19872,N_19963);
and UO_1731 (O_1731,N_19849,N_19938);
and UO_1732 (O_1732,N_19898,N_19935);
xor UO_1733 (O_1733,N_19952,N_19943);
nand UO_1734 (O_1734,N_19953,N_19882);
xor UO_1735 (O_1735,N_19860,N_19874);
nor UO_1736 (O_1736,N_19916,N_19802);
or UO_1737 (O_1737,N_19923,N_19874);
nand UO_1738 (O_1738,N_19889,N_19859);
xnor UO_1739 (O_1739,N_19925,N_19922);
nand UO_1740 (O_1740,N_19983,N_19984);
or UO_1741 (O_1741,N_19847,N_19904);
or UO_1742 (O_1742,N_19885,N_19813);
and UO_1743 (O_1743,N_19919,N_19932);
nand UO_1744 (O_1744,N_19996,N_19847);
nor UO_1745 (O_1745,N_19857,N_19871);
xnor UO_1746 (O_1746,N_19824,N_19952);
nand UO_1747 (O_1747,N_19932,N_19893);
nor UO_1748 (O_1748,N_19909,N_19815);
or UO_1749 (O_1749,N_19941,N_19998);
nand UO_1750 (O_1750,N_19864,N_19998);
and UO_1751 (O_1751,N_19990,N_19870);
nor UO_1752 (O_1752,N_19877,N_19946);
xor UO_1753 (O_1753,N_19954,N_19847);
or UO_1754 (O_1754,N_19818,N_19958);
xnor UO_1755 (O_1755,N_19836,N_19953);
and UO_1756 (O_1756,N_19968,N_19911);
xnor UO_1757 (O_1757,N_19915,N_19845);
or UO_1758 (O_1758,N_19856,N_19805);
or UO_1759 (O_1759,N_19907,N_19991);
nor UO_1760 (O_1760,N_19955,N_19829);
xor UO_1761 (O_1761,N_19864,N_19895);
nor UO_1762 (O_1762,N_19890,N_19835);
or UO_1763 (O_1763,N_19929,N_19988);
nor UO_1764 (O_1764,N_19926,N_19973);
xor UO_1765 (O_1765,N_19848,N_19892);
and UO_1766 (O_1766,N_19885,N_19986);
nor UO_1767 (O_1767,N_19886,N_19993);
nor UO_1768 (O_1768,N_19814,N_19876);
nor UO_1769 (O_1769,N_19923,N_19975);
xor UO_1770 (O_1770,N_19892,N_19814);
and UO_1771 (O_1771,N_19816,N_19810);
or UO_1772 (O_1772,N_19894,N_19997);
nor UO_1773 (O_1773,N_19953,N_19987);
nor UO_1774 (O_1774,N_19878,N_19884);
and UO_1775 (O_1775,N_19920,N_19836);
nand UO_1776 (O_1776,N_19965,N_19800);
or UO_1777 (O_1777,N_19829,N_19996);
or UO_1778 (O_1778,N_19924,N_19935);
and UO_1779 (O_1779,N_19999,N_19890);
xnor UO_1780 (O_1780,N_19805,N_19988);
and UO_1781 (O_1781,N_19918,N_19962);
xor UO_1782 (O_1782,N_19981,N_19915);
nor UO_1783 (O_1783,N_19807,N_19993);
nand UO_1784 (O_1784,N_19983,N_19924);
and UO_1785 (O_1785,N_19914,N_19941);
or UO_1786 (O_1786,N_19878,N_19885);
and UO_1787 (O_1787,N_19817,N_19934);
nor UO_1788 (O_1788,N_19887,N_19978);
nor UO_1789 (O_1789,N_19949,N_19907);
or UO_1790 (O_1790,N_19906,N_19843);
nor UO_1791 (O_1791,N_19943,N_19931);
and UO_1792 (O_1792,N_19845,N_19846);
xor UO_1793 (O_1793,N_19864,N_19968);
or UO_1794 (O_1794,N_19995,N_19863);
and UO_1795 (O_1795,N_19866,N_19889);
or UO_1796 (O_1796,N_19860,N_19836);
or UO_1797 (O_1797,N_19994,N_19851);
or UO_1798 (O_1798,N_19956,N_19953);
or UO_1799 (O_1799,N_19850,N_19925);
nand UO_1800 (O_1800,N_19890,N_19912);
and UO_1801 (O_1801,N_19987,N_19901);
and UO_1802 (O_1802,N_19809,N_19945);
nand UO_1803 (O_1803,N_19820,N_19913);
nand UO_1804 (O_1804,N_19952,N_19987);
nor UO_1805 (O_1805,N_19931,N_19889);
and UO_1806 (O_1806,N_19932,N_19942);
xor UO_1807 (O_1807,N_19887,N_19873);
and UO_1808 (O_1808,N_19877,N_19933);
xor UO_1809 (O_1809,N_19927,N_19934);
or UO_1810 (O_1810,N_19850,N_19926);
nand UO_1811 (O_1811,N_19847,N_19870);
nor UO_1812 (O_1812,N_19958,N_19854);
and UO_1813 (O_1813,N_19883,N_19870);
nor UO_1814 (O_1814,N_19934,N_19839);
and UO_1815 (O_1815,N_19909,N_19873);
nand UO_1816 (O_1816,N_19952,N_19973);
or UO_1817 (O_1817,N_19861,N_19940);
xor UO_1818 (O_1818,N_19929,N_19986);
or UO_1819 (O_1819,N_19844,N_19820);
nor UO_1820 (O_1820,N_19917,N_19803);
and UO_1821 (O_1821,N_19857,N_19876);
nand UO_1822 (O_1822,N_19844,N_19954);
or UO_1823 (O_1823,N_19915,N_19888);
nor UO_1824 (O_1824,N_19830,N_19937);
nor UO_1825 (O_1825,N_19962,N_19834);
or UO_1826 (O_1826,N_19937,N_19806);
or UO_1827 (O_1827,N_19917,N_19880);
nor UO_1828 (O_1828,N_19971,N_19978);
nand UO_1829 (O_1829,N_19976,N_19831);
and UO_1830 (O_1830,N_19912,N_19982);
and UO_1831 (O_1831,N_19979,N_19920);
or UO_1832 (O_1832,N_19932,N_19950);
nor UO_1833 (O_1833,N_19882,N_19834);
and UO_1834 (O_1834,N_19919,N_19899);
or UO_1835 (O_1835,N_19839,N_19952);
nand UO_1836 (O_1836,N_19884,N_19817);
or UO_1837 (O_1837,N_19943,N_19921);
nand UO_1838 (O_1838,N_19809,N_19941);
or UO_1839 (O_1839,N_19862,N_19849);
and UO_1840 (O_1840,N_19883,N_19947);
and UO_1841 (O_1841,N_19867,N_19856);
or UO_1842 (O_1842,N_19828,N_19836);
nand UO_1843 (O_1843,N_19870,N_19813);
xnor UO_1844 (O_1844,N_19822,N_19893);
and UO_1845 (O_1845,N_19876,N_19837);
or UO_1846 (O_1846,N_19944,N_19924);
or UO_1847 (O_1847,N_19888,N_19811);
xor UO_1848 (O_1848,N_19863,N_19914);
xnor UO_1849 (O_1849,N_19944,N_19820);
xnor UO_1850 (O_1850,N_19908,N_19872);
nand UO_1851 (O_1851,N_19991,N_19854);
nor UO_1852 (O_1852,N_19862,N_19915);
or UO_1853 (O_1853,N_19991,N_19880);
or UO_1854 (O_1854,N_19959,N_19848);
nand UO_1855 (O_1855,N_19950,N_19857);
nor UO_1856 (O_1856,N_19909,N_19972);
xnor UO_1857 (O_1857,N_19829,N_19984);
or UO_1858 (O_1858,N_19907,N_19893);
nand UO_1859 (O_1859,N_19983,N_19982);
and UO_1860 (O_1860,N_19927,N_19842);
or UO_1861 (O_1861,N_19937,N_19843);
nor UO_1862 (O_1862,N_19879,N_19856);
xnor UO_1863 (O_1863,N_19983,N_19812);
nand UO_1864 (O_1864,N_19805,N_19981);
and UO_1865 (O_1865,N_19929,N_19822);
or UO_1866 (O_1866,N_19901,N_19878);
nor UO_1867 (O_1867,N_19989,N_19933);
nor UO_1868 (O_1868,N_19936,N_19964);
or UO_1869 (O_1869,N_19862,N_19859);
or UO_1870 (O_1870,N_19937,N_19930);
nand UO_1871 (O_1871,N_19949,N_19994);
nor UO_1872 (O_1872,N_19862,N_19964);
and UO_1873 (O_1873,N_19924,N_19871);
and UO_1874 (O_1874,N_19863,N_19808);
xor UO_1875 (O_1875,N_19920,N_19855);
or UO_1876 (O_1876,N_19818,N_19856);
and UO_1877 (O_1877,N_19898,N_19876);
or UO_1878 (O_1878,N_19899,N_19869);
and UO_1879 (O_1879,N_19987,N_19835);
nor UO_1880 (O_1880,N_19997,N_19842);
nor UO_1881 (O_1881,N_19877,N_19887);
xnor UO_1882 (O_1882,N_19935,N_19972);
nand UO_1883 (O_1883,N_19919,N_19822);
xnor UO_1884 (O_1884,N_19948,N_19944);
and UO_1885 (O_1885,N_19987,N_19935);
nor UO_1886 (O_1886,N_19901,N_19906);
and UO_1887 (O_1887,N_19918,N_19984);
nand UO_1888 (O_1888,N_19816,N_19989);
or UO_1889 (O_1889,N_19996,N_19852);
xnor UO_1890 (O_1890,N_19934,N_19922);
nand UO_1891 (O_1891,N_19866,N_19919);
xnor UO_1892 (O_1892,N_19967,N_19915);
and UO_1893 (O_1893,N_19892,N_19974);
xor UO_1894 (O_1894,N_19939,N_19941);
nor UO_1895 (O_1895,N_19923,N_19953);
and UO_1896 (O_1896,N_19879,N_19906);
and UO_1897 (O_1897,N_19945,N_19926);
nand UO_1898 (O_1898,N_19879,N_19862);
nand UO_1899 (O_1899,N_19825,N_19830);
xor UO_1900 (O_1900,N_19925,N_19932);
nand UO_1901 (O_1901,N_19808,N_19941);
or UO_1902 (O_1902,N_19964,N_19982);
nor UO_1903 (O_1903,N_19927,N_19894);
xor UO_1904 (O_1904,N_19858,N_19933);
or UO_1905 (O_1905,N_19993,N_19954);
nand UO_1906 (O_1906,N_19962,N_19803);
xor UO_1907 (O_1907,N_19937,N_19975);
nand UO_1908 (O_1908,N_19868,N_19965);
xnor UO_1909 (O_1909,N_19872,N_19832);
nand UO_1910 (O_1910,N_19842,N_19861);
nor UO_1911 (O_1911,N_19973,N_19989);
or UO_1912 (O_1912,N_19895,N_19949);
or UO_1913 (O_1913,N_19806,N_19839);
and UO_1914 (O_1914,N_19930,N_19973);
or UO_1915 (O_1915,N_19886,N_19906);
and UO_1916 (O_1916,N_19898,N_19891);
xor UO_1917 (O_1917,N_19979,N_19919);
and UO_1918 (O_1918,N_19802,N_19834);
and UO_1919 (O_1919,N_19831,N_19974);
xor UO_1920 (O_1920,N_19939,N_19829);
xor UO_1921 (O_1921,N_19922,N_19910);
nand UO_1922 (O_1922,N_19985,N_19922);
or UO_1923 (O_1923,N_19855,N_19997);
nand UO_1924 (O_1924,N_19809,N_19892);
xor UO_1925 (O_1925,N_19888,N_19918);
or UO_1926 (O_1926,N_19801,N_19927);
nand UO_1927 (O_1927,N_19872,N_19920);
xnor UO_1928 (O_1928,N_19886,N_19927);
nand UO_1929 (O_1929,N_19931,N_19917);
xnor UO_1930 (O_1930,N_19820,N_19880);
nor UO_1931 (O_1931,N_19917,N_19889);
xnor UO_1932 (O_1932,N_19943,N_19918);
xnor UO_1933 (O_1933,N_19848,N_19980);
nor UO_1934 (O_1934,N_19974,N_19807);
or UO_1935 (O_1935,N_19893,N_19995);
and UO_1936 (O_1936,N_19972,N_19983);
xnor UO_1937 (O_1937,N_19873,N_19905);
nor UO_1938 (O_1938,N_19825,N_19986);
and UO_1939 (O_1939,N_19999,N_19922);
or UO_1940 (O_1940,N_19864,N_19802);
and UO_1941 (O_1941,N_19983,N_19863);
nand UO_1942 (O_1942,N_19867,N_19967);
nand UO_1943 (O_1943,N_19883,N_19807);
nand UO_1944 (O_1944,N_19878,N_19909);
nor UO_1945 (O_1945,N_19920,N_19928);
and UO_1946 (O_1946,N_19995,N_19924);
nor UO_1947 (O_1947,N_19997,N_19957);
nand UO_1948 (O_1948,N_19977,N_19903);
xnor UO_1949 (O_1949,N_19952,N_19999);
nand UO_1950 (O_1950,N_19846,N_19811);
xnor UO_1951 (O_1951,N_19985,N_19978);
nor UO_1952 (O_1952,N_19959,N_19825);
nand UO_1953 (O_1953,N_19858,N_19917);
nand UO_1954 (O_1954,N_19844,N_19949);
and UO_1955 (O_1955,N_19875,N_19883);
nand UO_1956 (O_1956,N_19938,N_19909);
xnor UO_1957 (O_1957,N_19908,N_19913);
or UO_1958 (O_1958,N_19964,N_19832);
xnor UO_1959 (O_1959,N_19894,N_19916);
nand UO_1960 (O_1960,N_19860,N_19848);
xnor UO_1961 (O_1961,N_19923,N_19904);
xor UO_1962 (O_1962,N_19924,N_19962);
and UO_1963 (O_1963,N_19998,N_19826);
nand UO_1964 (O_1964,N_19878,N_19853);
nand UO_1965 (O_1965,N_19979,N_19850);
or UO_1966 (O_1966,N_19904,N_19878);
and UO_1967 (O_1967,N_19877,N_19995);
or UO_1968 (O_1968,N_19979,N_19823);
and UO_1969 (O_1969,N_19833,N_19836);
xor UO_1970 (O_1970,N_19910,N_19889);
nor UO_1971 (O_1971,N_19906,N_19838);
xnor UO_1972 (O_1972,N_19851,N_19903);
or UO_1973 (O_1973,N_19858,N_19940);
or UO_1974 (O_1974,N_19808,N_19966);
and UO_1975 (O_1975,N_19865,N_19972);
and UO_1976 (O_1976,N_19971,N_19967);
xor UO_1977 (O_1977,N_19800,N_19845);
nand UO_1978 (O_1978,N_19883,N_19876);
nand UO_1979 (O_1979,N_19838,N_19891);
nor UO_1980 (O_1980,N_19997,N_19944);
or UO_1981 (O_1981,N_19983,N_19877);
nor UO_1982 (O_1982,N_19881,N_19864);
and UO_1983 (O_1983,N_19949,N_19905);
or UO_1984 (O_1984,N_19911,N_19920);
nand UO_1985 (O_1985,N_19951,N_19926);
and UO_1986 (O_1986,N_19847,N_19976);
or UO_1987 (O_1987,N_19985,N_19824);
and UO_1988 (O_1988,N_19924,N_19943);
nor UO_1989 (O_1989,N_19870,N_19845);
nand UO_1990 (O_1990,N_19804,N_19887);
nor UO_1991 (O_1991,N_19806,N_19856);
and UO_1992 (O_1992,N_19844,N_19942);
xnor UO_1993 (O_1993,N_19895,N_19975);
nand UO_1994 (O_1994,N_19998,N_19968);
and UO_1995 (O_1995,N_19829,N_19974);
nor UO_1996 (O_1996,N_19923,N_19956);
and UO_1997 (O_1997,N_19916,N_19962);
nor UO_1998 (O_1998,N_19978,N_19955);
and UO_1999 (O_1999,N_19961,N_19939);
and UO_2000 (O_2000,N_19921,N_19939);
nand UO_2001 (O_2001,N_19960,N_19834);
or UO_2002 (O_2002,N_19821,N_19963);
and UO_2003 (O_2003,N_19872,N_19874);
nor UO_2004 (O_2004,N_19879,N_19895);
and UO_2005 (O_2005,N_19986,N_19821);
nor UO_2006 (O_2006,N_19856,N_19829);
nor UO_2007 (O_2007,N_19947,N_19816);
nor UO_2008 (O_2008,N_19865,N_19854);
and UO_2009 (O_2009,N_19816,N_19891);
xor UO_2010 (O_2010,N_19838,N_19883);
nand UO_2011 (O_2011,N_19998,N_19895);
and UO_2012 (O_2012,N_19865,N_19968);
xor UO_2013 (O_2013,N_19873,N_19867);
nor UO_2014 (O_2014,N_19867,N_19815);
nor UO_2015 (O_2015,N_19871,N_19867);
xor UO_2016 (O_2016,N_19856,N_19988);
or UO_2017 (O_2017,N_19814,N_19900);
xnor UO_2018 (O_2018,N_19931,N_19883);
nor UO_2019 (O_2019,N_19948,N_19860);
and UO_2020 (O_2020,N_19933,N_19966);
nand UO_2021 (O_2021,N_19968,N_19933);
nor UO_2022 (O_2022,N_19857,N_19840);
nor UO_2023 (O_2023,N_19801,N_19933);
and UO_2024 (O_2024,N_19889,N_19854);
nor UO_2025 (O_2025,N_19837,N_19921);
nand UO_2026 (O_2026,N_19937,N_19934);
and UO_2027 (O_2027,N_19985,N_19880);
or UO_2028 (O_2028,N_19934,N_19991);
nor UO_2029 (O_2029,N_19907,N_19869);
nand UO_2030 (O_2030,N_19990,N_19879);
nor UO_2031 (O_2031,N_19985,N_19817);
nor UO_2032 (O_2032,N_19840,N_19940);
xor UO_2033 (O_2033,N_19841,N_19983);
or UO_2034 (O_2034,N_19971,N_19949);
nor UO_2035 (O_2035,N_19890,N_19858);
nand UO_2036 (O_2036,N_19930,N_19860);
and UO_2037 (O_2037,N_19850,N_19813);
nor UO_2038 (O_2038,N_19991,N_19849);
and UO_2039 (O_2039,N_19804,N_19885);
or UO_2040 (O_2040,N_19895,N_19947);
or UO_2041 (O_2041,N_19913,N_19852);
xnor UO_2042 (O_2042,N_19899,N_19896);
nor UO_2043 (O_2043,N_19916,N_19805);
nand UO_2044 (O_2044,N_19817,N_19962);
or UO_2045 (O_2045,N_19997,N_19921);
and UO_2046 (O_2046,N_19889,N_19862);
nand UO_2047 (O_2047,N_19926,N_19949);
or UO_2048 (O_2048,N_19807,N_19995);
and UO_2049 (O_2049,N_19975,N_19867);
or UO_2050 (O_2050,N_19804,N_19998);
nand UO_2051 (O_2051,N_19957,N_19847);
nor UO_2052 (O_2052,N_19987,N_19848);
nand UO_2053 (O_2053,N_19844,N_19983);
and UO_2054 (O_2054,N_19967,N_19988);
or UO_2055 (O_2055,N_19832,N_19829);
nor UO_2056 (O_2056,N_19855,N_19955);
nand UO_2057 (O_2057,N_19933,N_19854);
nand UO_2058 (O_2058,N_19968,N_19977);
xor UO_2059 (O_2059,N_19969,N_19937);
nand UO_2060 (O_2060,N_19931,N_19941);
and UO_2061 (O_2061,N_19930,N_19890);
nor UO_2062 (O_2062,N_19962,N_19890);
nand UO_2063 (O_2063,N_19988,N_19951);
or UO_2064 (O_2064,N_19967,N_19973);
or UO_2065 (O_2065,N_19827,N_19813);
nand UO_2066 (O_2066,N_19991,N_19845);
nor UO_2067 (O_2067,N_19996,N_19800);
xnor UO_2068 (O_2068,N_19936,N_19912);
nand UO_2069 (O_2069,N_19871,N_19921);
nor UO_2070 (O_2070,N_19892,N_19964);
xnor UO_2071 (O_2071,N_19944,N_19834);
nand UO_2072 (O_2072,N_19846,N_19984);
and UO_2073 (O_2073,N_19921,N_19852);
or UO_2074 (O_2074,N_19916,N_19975);
nand UO_2075 (O_2075,N_19850,N_19906);
xnor UO_2076 (O_2076,N_19814,N_19844);
nor UO_2077 (O_2077,N_19918,N_19802);
and UO_2078 (O_2078,N_19966,N_19928);
and UO_2079 (O_2079,N_19870,N_19972);
xor UO_2080 (O_2080,N_19870,N_19874);
nand UO_2081 (O_2081,N_19859,N_19843);
or UO_2082 (O_2082,N_19949,N_19956);
and UO_2083 (O_2083,N_19908,N_19883);
nand UO_2084 (O_2084,N_19916,N_19943);
nand UO_2085 (O_2085,N_19909,N_19907);
or UO_2086 (O_2086,N_19912,N_19862);
or UO_2087 (O_2087,N_19992,N_19880);
or UO_2088 (O_2088,N_19831,N_19813);
nand UO_2089 (O_2089,N_19811,N_19991);
nand UO_2090 (O_2090,N_19871,N_19955);
nand UO_2091 (O_2091,N_19840,N_19855);
xor UO_2092 (O_2092,N_19940,N_19970);
nor UO_2093 (O_2093,N_19834,N_19923);
nand UO_2094 (O_2094,N_19926,N_19898);
xor UO_2095 (O_2095,N_19837,N_19938);
xor UO_2096 (O_2096,N_19881,N_19906);
or UO_2097 (O_2097,N_19987,N_19845);
xor UO_2098 (O_2098,N_19876,N_19862);
or UO_2099 (O_2099,N_19899,N_19851);
xor UO_2100 (O_2100,N_19911,N_19816);
nand UO_2101 (O_2101,N_19806,N_19938);
nand UO_2102 (O_2102,N_19818,N_19857);
nor UO_2103 (O_2103,N_19908,N_19987);
xnor UO_2104 (O_2104,N_19862,N_19969);
xor UO_2105 (O_2105,N_19875,N_19941);
xor UO_2106 (O_2106,N_19973,N_19981);
or UO_2107 (O_2107,N_19801,N_19940);
xor UO_2108 (O_2108,N_19857,N_19813);
and UO_2109 (O_2109,N_19867,N_19839);
nor UO_2110 (O_2110,N_19843,N_19860);
or UO_2111 (O_2111,N_19876,N_19892);
and UO_2112 (O_2112,N_19986,N_19826);
and UO_2113 (O_2113,N_19986,N_19855);
or UO_2114 (O_2114,N_19994,N_19833);
nor UO_2115 (O_2115,N_19823,N_19965);
and UO_2116 (O_2116,N_19946,N_19892);
nand UO_2117 (O_2117,N_19865,N_19939);
nand UO_2118 (O_2118,N_19981,N_19956);
or UO_2119 (O_2119,N_19992,N_19859);
xnor UO_2120 (O_2120,N_19950,N_19959);
xor UO_2121 (O_2121,N_19995,N_19942);
or UO_2122 (O_2122,N_19974,N_19931);
nand UO_2123 (O_2123,N_19823,N_19807);
or UO_2124 (O_2124,N_19849,N_19963);
or UO_2125 (O_2125,N_19983,N_19988);
and UO_2126 (O_2126,N_19866,N_19802);
xor UO_2127 (O_2127,N_19845,N_19814);
nor UO_2128 (O_2128,N_19886,N_19970);
nor UO_2129 (O_2129,N_19990,N_19965);
nor UO_2130 (O_2130,N_19821,N_19859);
nand UO_2131 (O_2131,N_19981,N_19989);
or UO_2132 (O_2132,N_19948,N_19859);
xnor UO_2133 (O_2133,N_19986,N_19934);
nand UO_2134 (O_2134,N_19873,N_19872);
nand UO_2135 (O_2135,N_19868,N_19883);
nand UO_2136 (O_2136,N_19857,N_19941);
nor UO_2137 (O_2137,N_19883,N_19864);
xor UO_2138 (O_2138,N_19866,N_19934);
nand UO_2139 (O_2139,N_19926,N_19995);
nand UO_2140 (O_2140,N_19985,N_19819);
or UO_2141 (O_2141,N_19953,N_19904);
or UO_2142 (O_2142,N_19898,N_19878);
or UO_2143 (O_2143,N_19812,N_19944);
xnor UO_2144 (O_2144,N_19912,N_19925);
nand UO_2145 (O_2145,N_19806,N_19819);
and UO_2146 (O_2146,N_19901,N_19896);
nor UO_2147 (O_2147,N_19930,N_19813);
xnor UO_2148 (O_2148,N_19913,N_19871);
nor UO_2149 (O_2149,N_19966,N_19888);
nand UO_2150 (O_2150,N_19853,N_19939);
nand UO_2151 (O_2151,N_19907,N_19887);
and UO_2152 (O_2152,N_19859,N_19876);
nand UO_2153 (O_2153,N_19926,N_19985);
nand UO_2154 (O_2154,N_19842,N_19909);
xor UO_2155 (O_2155,N_19887,N_19822);
nand UO_2156 (O_2156,N_19885,N_19851);
nand UO_2157 (O_2157,N_19918,N_19915);
and UO_2158 (O_2158,N_19920,N_19882);
nand UO_2159 (O_2159,N_19853,N_19992);
nor UO_2160 (O_2160,N_19837,N_19947);
nand UO_2161 (O_2161,N_19821,N_19881);
nand UO_2162 (O_2162,N_19873,N_19941);
or UO_2163 (O_2163,N_19866,N_19959);
xor UO_2164 (O_2164,N_19830,N_19967);
nor UO_2165 (O_2165,N_19800,N_19934);
and UO_2166 (O_2166,N_19959,N_19876);
nor UO_2167 (O_2167,N_19925,N_19805);
nand UO_2168 (O_2168,N_19949,N_19980);
nand UO_2169 (O_2169,N_19900,N_19997);
nand UO_2170 (O_2170,N_19821,N_19824);
and UO_2171 (O_2171,N_19923,N_19964);
and UO_2172 (O_2172,N_19812,N_19814);
or UO_2173 (O_2173,N_19802,N_19826);
or UO_2174 (O_2174,N_19998,N_19991);
and UO_2175 (O_2175,N_19942,N_19908);
xnor UO_2176 (O_2176,N_19896,N_19918);
or UO_2177 (O_2177,N_19945,N_19810);
nor UO_2178 (O_2178,N_19930,N_19856);
or UO_2179 (O_2179,N_19969,N_19939);
nand UO_2180 (O_2180,N_19961,N_19927);
nor UO_2181 (O_2181,N_19997,N_19807);
or UO_2182 (O_2182,N_19867,N_19806);
or UO_2183 (O_2183,N_19973,N_19995);
or UO_2184 (O_2184,N_19949,N_19987);
and UO_2185 (O_2185,N_19924,N_19972);
or UO_2186 (O_2186,N_19928,N_19984);
nor UO_2187 (O_2187,N_19948,N_19915);
nor UO_2188 (O_2188,N_19834,N_19903);
nand UO_2189 (O_2189,N_19828,N_19846);
or UO_2190 (O_2190,N_19825,N_19860);
nor UO_2191 (O_2191,N_19874,N_19837);
or UO_2192 (O_2192,N_19883,N_19829);
xor UO_2193 (O_2193,N_19805,N_19931);
xnor UO_2194 (O_2194,N_19836,N_19874);
nand UO_2195 (O_2195,N_19860,N_19944);
nand UO_2196 (O_2196,N_19965,N_19935);
and UO_2197 (O_2197,N_19959,N_19819);
nand UO_2198 (O_2198,N_19883,N_19984);
nand UO_2199 (O_2199,N_19861,N_19984);
nand UO_2200 (O_2200,N_19809,N_19966);
xnor UO_2201 (O_2201,N_19901,N_19981);
and UO_2202 (O_2202,N_19862,N_19971);
and UO_2203 (O_2203,N_19992,N_19944);
xor UO_2204 (O_2204,N_19892,N_19951);
nor UO_2205 (O_2205,N_19801,N_19876);
or UO_2206 (O_2206,N_19888,N_19961);
nor UO_2207 (O_2207,N_19950,N_19990);
or UO_2208 (O_2208,N_19957,N_19899);
nor UO_2209 (O_2209,N_19951,N_19939);
or UO_2210 (O_2210,N_19885,N_19931);
and UO_2211 (O_2211,N_19801,N_19896);
or UO_2212 (O_2212,N_19985,N_19990);
nor UO_2213 (O_2213,N_19935,N_19993);
nand UO_2214 (O_2214,N_19859,N_19851);
nor UO_2215 (O_2215,N_19975,N_19884);
or UO_2216 (O_2216,N_19975,N_19976);
and UO_2217 (O_2217,N_19902,N_19930);
xor UO_2218 (O_2218,N_19885,N_19938);
nor UO_2219 (O_2219,N_19857,N_19926);
nand UO_2220 (O_2220,N_19834,N_19879);
or UO_2221 (O_2221,N_19877,N_19874);
xnor UO_2222 (O_2222,N_19824,N_19976);
nor UO_2223 (O_2223,N_19939,N_19970);
or UO_2224 (O_2224,N_19872,N_19945);
xnor UO_2225 (O_2225,N_19906,N_19878);
or UO_2226 (O_2226,N_19970,N_19915);
or UO_2227 (O_2227,N_19924,N_19862);
and UO_2228 (O_2228,N_19827,N_19900);
and UO_2229 (O_2229,N_19843,N_19955);
and UO_2230 (O_2230,N_19871,N_19879);
nor UO_2231 (O_2231,N_19991,N_19921);
or UO_2232 (O_2232,N_19886,N_19888);
nor UO_2233 (O_2233,N_19968,N_19868);
or UO_2234 (O_2234,N_19991,N_19957);
nand UO_2235 (O_2235,N_19971,N_19938);
nand UO_2236 (O_2236,N_19890,N_19899);
or UO_2237 (O_2237,N_19997,N_19841);
and UO_2238 (O_2238,N_19974,N_19826);
nor UO_2239 (O_2239,N_19820,N_19868);
or UO_2240 (O_2240,N_19884,N_19993);
nand UO_2241 (O_2241,N_19839,N_19842);
nand UO_2242 (O_2242,N_19900,N_19971);
or UO_2243 (O_2243,N_19908,N_19978);
or UO_2244 (O_2244,N_19958,N_19939);
or UO_2245 (O_2245,N_19898,N_19806);
nor UO_2246 (O_2246,N_19844,N_19886);
nand UO_2247 (O_2247,N_19907,N_19802);
xor UO_2248 (O_2248,N_19878,N_19835);
xor UO_2249 (O_2249,N_19937,N_19927);
xor UO_2250 (O_2250,N_19812,N_19967);
and UO_2251 (O_2251,N_19857,N_19922);
and UO_2252 (O_2252,N_19915,N_19836);
nor UO_2253 (O_2253,N_19979,N_19982);
nand UO_2254 (O_2254,N_19909,N_19851);
xor UO_2255 (O_2255,N_19859,N_19914);
or UO_2256 (O_2256,N_19870,N_19919);
nor UO_2257 (O_2257,N_19982,N_19897);
nor UO_2258 (O_2258,N_19808,N_19997);
nand UO_2259 (O_2259,N_19832,N_19879);
xor UO_2260 (O_2260,N_19908,N_19894);
and UO_2261 (O_2261,N_19915,N_19830);
and UO_2262 (O_2262,N_19866,N_19873);
nand UO_2263 (O_2263,N_19804,N_19832);
xor UO_2264 (O_2264,N_19805,N_19876);
nor UO_2265 (O_2265,N_19879,N_19816);
or UO_2266 (O_2266,N_19845,N_19869);
xnor UO_2267 (O_2267,N_19855,N_19909);
xor UO_2268 (O_2268,N_19923,N_19811);
nand UO_2269 (O_2269,N_19859,N_19852);
and UO_2270 (O_2270,N_19931,N_19891);
or UO_2271 (O_2271,N_19868,N_19810);
xnor UO_2272 (O_2272,N_19971,N_19806);
xnor UO_2273 (O_2273,N_19971,N_19873);
or UO_2274 (O_2274,N_19812,N_19858);
and UO_2275 (O_2275,N_19842,N_19920);
and UO_2276 (O_2276,N_19838,N_19899);
xnor UO_2277 (O_2277,N_19965,N_19938);
xor UO_2278 (O_2278,N_19833,N_19977);
or UO_2279 (O_2279,N_19800,N_19955);
or UO_2280 (O_2280,N_19980,N_19898);
or UO_2281 (O_2281,N_19973,N_19996);
and UO_2282 (O_2282,N_19811,N_19942);
nand UO_2283 (O_2283,N_19835,N_19816);
xor UO_2284 (O_2284,N_19845,N_19917);
xor UO_2285 (O_2285,N_19965,N_19913);
nor UO_2286 (O_2286,N_19875,N_19963);
and UO_2287 (O_2287,N_19919,N_19891);
or UO_2288 (O_2288,N_19885,N_19803);
or UO_2289 (O_2289,N_19905,N_19800);
nor UO_2290 (O_2290,N_19914,N_19834);
and UO_2291 (O_2291,N_19801,N_19983);
nor UO_2292 (O_2292,N_19889,N_19934);
xor UO_2293 (O_2293,N_19839,N_19959);
nand UO_2294 (O_2294,N_19823,N_19831);
nor UO_2295 (O_2295,N_19916,N_19889);
or UO_2296 (O_2296,N_19935,N_19822);
nand UO_2297 (O_2297,N_19839,N_19977);
or UO_2298 (O_2298,N_19849,N_19812);
and UO_2299 (O_2299,N_19869,N_19928);
and UO_2300 (O_2300,N_19971,N_19999);
and UO_2301 (O_2301,N_19971,N_19951);
nand UO_2302 (O_2302,N_19869,N_19978);
nand UO_2303 (O_2303,N_19940,N_19811);
xnor UO_2304 (O_2304,N_19832,N_19900);
nor UO_2305 (O_2305,N_19938,N_19962);
and UO_2306 (O_2306,N_19951,N_19952);
nand UO_2307 (O_2307,N_19842,N_19889);
xor UO_2308 (O_2308,N_19991,N_19899);
nor UO_2309 (O_2309,N_19968,N_19935);
nor UO_2310 (O_2310,N_19929,N_19894);
nor UO_2311 (O_2311,N_19837,N_19881);
nor UO_2312 (O_2312,N_19990,N_19889);
nand UO_2313 (O_2313,N_19971,N_19943);
or UO_2314 (O_2314,N_19865,N_19887);
nor UO_2315 (O_2315,N_19982,N_19930);
nand UO_2316 (O_2316,N_19850,N_19930);
xor UO_2317 (O_2317,N_19962,N_19930);
nand UO_2318 (O_2318,N_19925,N_19803);
and UO_2319 (O_2319,N_19865,N_19846);
and UO_2320 (O_2320,N_19922,N_19900);
xor UO_2321 (O_2321,N_19886,N_19950);
nand UO_2322 (O_2322,N_19849,N_19953);
xor UO_2323 (O_2323,N_19822,N_19898);
nand UO_2324 (O_2324,N_19801,N_19875);
nor UO_2325 (O_2325,N_19886,N_19901);
xor UO_2326 (O_2326,N_19808,N_19904);
or UO_2327 (O_2327,N_19944,N_19942);
and UO_2328 (O_2328,N_19891,N_19818);
and UO_2329 (O_2329,N_19950,N_19865);
nand UO_2330 (O_2330,N_19931,N_19934);
nand UO_2331 (O_2331,N_19945,N_19868);
xor UO_2332 (O_2332,N_19860,N_19934);
nand UO_2333 (O_2333,N_19831,N_19927);
nor UO_2334 (O_2334,N_19877,N_19959);
and UO_2335 (O_2335,N_19873,N_19980);
nand UO_2336 (O_2336,N_19964,N_19872);
and UO_2337 (O_2337,N_19887,N_19814);
xnor UO_2338 (O_2338,N_19893,N_19998);
nand UO_2339 (O_2339,N_19894,N_19974);
xor UO_2340 (O_2340,N_19927,N_19814);
and UO_2341 (O_2341,N_19875,N_19944);
nand UO_2342 (O_2342,N_19979,N_19889);
or UO_2343 (O_2343,N_19885,N_19913);
nor UO_2344 (O_2344,N_19999,N_19828);
or UO_2345 (O_2345,N_19886,N_19838);
nor UO_2346 (O_2346,N_19933,N_19942);
nand UO_2347 (O_2347,N_19833,N_19954);
nor UO_2348 (O_2348,N_19808,N_19887);
or UO_2349 (O_2349,N_19990,N_19953);
nor UO_2350 (O_2350,N_19957,N_19958);
xor UO_2351 (O_2351,N_19938,N_19972);
xnor UO_2352 (O_2352,N_19837,N_19843);
and UO_2353 (O_2353,N_19877,N_19854);
xor UO_2354 (O_2354,N_19845,N_19934);
or UO_2355 (O_2355,N_19973,N_19942);
or UO_2356 (O_2356,N_19904,N_19954);
nor UO_2357 (O_2357,N_19880,N_19947);
nand UO_2358 (O_2358,N_19936,N_19837);
or UO_2359 (O_2359,N_19862,N_19839);
nor UO_2360 (O_2360,N_19971,N_19941);
or UO_2361 (O_2361,N_19927,N_19912);
xor UO_2362 (O_2362,N_19814,N_19852);
nand UO_2363 (O_2363,N_19869,N_19841);
or UO_2364 (O_2364,N_19952,N_19984);
xnor UO_2365 (O_2365,N_19812,N_19864);
xor UO_2366 (O_2366,N_19974,N_19867);
or UO_2367 (O_2367,N_19876,N_19828);
and UO_2368 (O_2368,N_19856,N_19925);
and UO_2369 (O_2369,N_19977,N_19937);
nor UO_2370 (O_2370,N_19823,N_19863);
and UO_2371 (O_2371,N_19841,N_19924);
xor UO_2372 (O_2372,N_19868,N_19848);
nor UO_2373 (O_2373,N_19982,N_19908);
xnor UO_2374 (O_2374,N_19818,N_19992);
and UO_2375 (O_2375,N_19904,N_19892);
and UO_2376 (O_2376,N_19915,N_19978);
or UO_2377 (O_2377,N_19850,N_19951);
xnor UO_2378 (O_2378,N_19938,N_19912);
xor UO_2379 (O_2379,N_19962,N_19863);
nor UO_2380 (O_2380,N_19834,N_19817);
or UO_2381 (O_2381,N_19821,N_19836);
or UO_2382 (O_2382,N_19932,N_19897);
nor UO_2383 (O_2383,N_19859,N_19940);
nor UO_2384 (O_2384,N_19828,N_19934);
and UO_2385 (O_2385,N_19809,N_19911);
nand UO_2386 (O_2386,N_19854,N_19824);
nor UO_2387 (O_2387,N_19870,N_19868);
or UO_2388 (O_2388,N_19927,N_19895);
xor UO_2389 (O_2389,N_19842,N_19945);
nor UO_2390 (O_2390,N_19984,N_19929);
and UO_2391 (O_2391,N_19938,N_19986);
and UO_2392 (O_2392,N_19999,N_19926);
nor UO_2393 (O_2393,N_19924,N_19949);
nand UO_2394 (O_2394,N_19840,N_19939);
and UO_2395 (O_2395,N_19936,N_19887);
and UO_2396 (O_2396,N_19848,N_19816);
and UO_2397 (O_2397,N_19873,N_19836);
xnor UO_2398 (O_2398,N_19843,N_19809);
nor UO_2399 (O_2399,N_19931,N_19894);
nor UO_2400 (O_2400,N_19867,N_19991);
xnor UO_2401 (O_2401,N_19874,N_19958);
nor UO_2402 (O_2402,N_19811,N_19965);
or UO_2403 (O_2403,N_19976,N_19874);
xor UO_2404 (O_2404,N_19833,N_19819);
xnor UO_2405 (O_2405,N_19809,N_19914);
nor UO_2406 (O_2406,N_19908,N_19935);
nor UO_2407 (O_2407,N_19942,N_19885);
xnor UO_2408 (O_2408,N_19958,N_19918);
or UO_2409 (O_2409,N_19983,N_19891);
and UO_2410 (O_2410,N_19934,N_19912);
nor UO_2411 (O_2411,N_19928,N_19930);
and UO_2412 (O_2412,N_19832,N_19970);
nand UO_2413 (O_2413,N_19918,N_19810);
nand UO_2414 (O_2414,N_19927,N_19903);
and UO_2415 (O_2415,N_19952,N_19871);
nand UO_2416 (O_2416,N_19876,N_19923);
and UO_2417 (O_2417,N_19868,N_19978);
and UO_2418 (O_2418,N_19884,N_19868);
nand UO_2419 (O_2419,N_19997,N_19806);
nand UO_2420 (O_2420,N_19937,N_19998);
nand UO_2421 (O_2421,N_19876,N_19891);
xor UO_2422 (O_2422,N_19962,N_19856);
nor UO_2423 (O_2423,N_19944,N_19971);
and UO_2424 (O_2424,N_19907,N_19901);
or UO_2425 (O_2425,N_19832,N_19935);
xnor UO_2426 (O_2426,N_19802,N_19810);
nor UO_2427 (O_2427,N_19862,N_19820);
nand UO_2428 (O_2428,N_19985,N_19836);
nand UO_2429 (O_2429,N_19824,N_19879);
and UO_2430 (O_2430,N_19951,N_19827);
nand UO_2431 (O_2431,N_19862,N_19811);
nor UO_2432 (O_2432,N_19836,N_19876);
nand UO_2433 (O_2433,N_19930,N_19875);
xnor UO_2434 (O_2434,N_19985,N_19825);
and UO_2435 (O_2435,N_19907,N_19996);
nand UO_2436 (O_2436,N_19972,N_19964);
nand UO_2437 (O_2437,N_19960,N_19997);
nand UO_2438 (O_2438,N_19900,N_19843);
xnor UO_2439 (O_2439,N_19857,N_19947);
or UO_2440 (O_2440,N_19977,N_19974);
xnor UO_2441 (O_2441,N_19992,N_19939);
nand UO_2442 (O_2442,N_19994,N_19920);
or UO_2443 (O_2443,N_19848,N_19907);
or UO_2444 (O_2444,N_19958,N_19878);
nor UO_2445 (O_2445,N_19809,N_19936);
or UO_2446 (O_2446,N_19905,N_19996);
or UO_2447 (O_2447,N_19911,N_19825);
nand UO_2448 (O_2448,N_19944,N_19831);
or UO_2449 (O_2449,N_19827,N_19894);
nor UO_2450 (O_2450,N_19874,N_19884);
xnor UO_2451 (O_2451,N_19947,N_19993);
and UO_2452 (O_2452,N_19945,N_19870);
or UO_2453 (O_2453,N_19840,N_19883);
or UO_2454 (O_2454,N_19854,N_19974);
nand UO_2455 (O_2455,N_19926,N_19938);
or UO_2456 (O_2456,N_19947,N_19893);
nand UO_2457 (O_2457,N_19936,N_19983);
and UO_2458 (O_2458,N_19884,N_19954);
xor UO_2459 (O_2459,N_19839,N_19818);
nand UO_2460 (O_2460,N_19934,N_19803);
xor UO_2461 (O_2461,N_19900,N_19842);
or UO_2462 (O_2462,N_19847,N_19874);
or UO_2463 (O_2463,N_19965,N_19869);
and UO_2464 (O_2464,N_19822,N_19966);
nand UO_2465 (O_2465,N_19801,N_19812);
or UO_2466 (O_2466,N_19956,N_19833);
nor UO_2467 (O_2467,N_19943,N_19975);
or UO_2468 (O_2468,N_19957,N_19874);
nor UO_2469 (O_2469,N_19973,N_19869);
nor UO_2470 (O_2470,N_19912,N_19902);
nand UO_2471 (O_2471,N_19996,N_19866);
and UO_2472 (O_2472,N_19987,N_19829);
and UO_2473 (O_2473,N_19800,N_19876);
or UO_2474 (O_2474,N_19932,N_19906);
and UO_2475 (O_2475,N_19938,N_19844);
nand UO_2476 (O_2476,N_19962,N_19946);
and UO_2477 (O_2477,N_19985,N_19877);
and UO_2478 (O_2478,N_19863,N_19884);
or UO_2479 (O_2479,N_19889,N_19822);
nor UO_2480 (O_2480,N_19896,N_19916);
xor UO_2481 (O_2481,N_19914,N_19989);
xor UO_2482 (O_2482,N_19928,N_19912);
and UO_2483 (O_2483,N_19975,N_19913);
nand UO_2484 (O_2484,N_19884,N_19870);
and UO_2485 (O_2485,N_19889,N_19945);
and UO_2486 (O_2486,N_19935,N_19840);
and UO_2487 (O_2487,N_19821,N_19943);
or UO_2488 (O_2488,N_19811,N_19854);
nand UO_2489 (O_2489,N_19861,N_19935);
nand UO_2490 (O_2490,N_19977,N_19998);
nor UO_2491 (O_2491,N_19839,N_19830);
nor UO_2492 (O_2492,N_19893,N_19956);
xor UO_2493 (O_2493,N_19921,N_19903);
xor UO_2494 (O_2494,N_19969,N_19928);
or UO_2495 (O_2495,N_19948,N_19921);
and UO_2496 (O_2496,N_19823,N_19801);
xor UO_2497 (O_2497,N_19862,N_19990);
nand UO_2498 (O_2498,N_19869,N_19890);
xnor UO_2499 (O_2499,N_19992,N_19803);
endmodule