module basic_2500_25000_3000_100_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
xnor U0 (N_0,In_2373,In_232);
and U1 (N_1,In_1419,In_936);
xnor U2 (N_2,In_443,In_1891);
nor U3 (N_3,In_2391,In_323);
nand U4 (N_4,In_1988,In_292);
nor U5 (N_5,In_568,In_2289);
or U6 (N_6,In_1072,In_2393);
and U7 (N_7,In_131,In_2185);
and U8 (N_8,In_1798,In_1390);
and U9 (N_9,In_836,In_894);
and U10 (N_10,In_1590,In_1909);
and U11 (N_11,In_522,In_286);
nand U12 (N_12,In_2330,In_2421);
and U13 (N_13,In_1217,In_576);
xnor U14 (N_14,In_351,In_1287);
nand U15 (N_15,In_2009,In_1858);
or U16 (N_16,In_1462,In_2323);
and U17 (N_17,In_1260,In_1520);
nor U18 (N_18,In_2285,In_1318);
or U19 (N_19,In_693,In_1888);
and U20 (N_20,In_841,In_1709);
nor U21 (N_21,In_1400,In_1621);
nand U22 (N_22,In_1420,In_1999);
xor U23 (N_23,In_220,In_1336);
and U24 (N_24,In_1296,In_630);
nand U25 (N_25,In_2075,In_1153);
nor U26 (N_26,In_2299,In_843);
and U27 (N_27,In_2275,In_477);
nand U28 (N_28,In_791,In_1130);
nand U29 (N_29,In_370,In_1345);
and U30 (N_30,In_2370,In_1223);
nor U31 (N_31,In_2423,In_1716);
nand U32 (N_32,In_2014,In_1529);
nand U33 (N_33,In_1134,In_618);
or U34 (N_34,In_119,In_672);
and U35 (N_35,In_1577,In_1768);
nor U36 (N_36,In_1237,In_2283);
nand U37 (N_37,In_2233,In_954);
nand U38 (N_38,In_668,In_752);
and U39 (N_39,In_1281,In_859);
xor U40 (N_40,In_1110,In_1450);
or U41 (N_41,In_1808,In_1763);
nor U42 (N_42,In_2415,In_2187);
nand U43 (N_43,In_1109,In_985);
nor U44 (N_44,In_1162,In_275);
xnor U45 (N_45,In_2427,In_1635);
nor U46 (N_46,In_1136,In_1949);
or U47 (N_47,In_747,In_2013);
or U48 (N_48,In_1322,In_1634);
xnor U49 (N_49,In_85,In_920);
nor U50 (N_50,In_792,In_1649);
nand U51 (N_51,In_1169,In_1492);
or U52 (N_52,In_529,In_498);
nor U53 (N_53,In_1044,In_338);
xnor U54 (N_54,In_1508,In_614);
nor U55 (N_55,In_1176,In_595);
and U56 (N_56,In_2206,In_136);
nor U57 (N_57,In_208,In_1405);
and U58 (N_58,In_188,In_2177);
nor U59 (N_59,In_1097,In_272);
nand U60 (N_60,In_611,In_999);
or U61 (N_61,In_678,In_949);
and U62 (N_62,In_2459,In_809);
nand U63 (N_63,In_1275,In_386);
or U64 (N_64,In_1922,In_1393);
or U65 (N_65,In_1025,In_1923);
xnor U66 (N_66,In_1631,In_723);
xnor U67 (N_67,In_2196,In_2113);
nand U68 (N_68,In_2496,In_24);
or U69 (N_69,In_2444,In_1997);
nand U70 (N_70,In_2062,In_337);
nor U71 (N_71,In_2153,In_1066);
or U72 (N_72,In_1510,In_1576);
nor U73 (N_73,In_74,In_2377);
or U74 (N_74,In_38,In_176);
and U75 (N_75,In_2333,In_589);
or U76 (N_76,In_459,In_1690);
nor U77 (N_77,In_1443,In_1158);
nand U78 (N_78,In_811,In_1863);
nor U79 (N_79,In_1561,In_2032);
nand U80 (N_80,In_2315,In_2350);
xor U81 (N_81,In_1804,In_264);
and U82 (N_82,In_1685,In_2202);
nor U83 (N_83,In_591,In_671);
or U84 (N_84,In_2473,In_1491);
xor U85 (N_85,In_265,In_1567);
nor U86 (N_86,In_1955,In_2383);
nand U87 (N_87,In_1924,In_1504);
nand U88 (N_88,In_2073,In_395);
nand U89 (N_89,In_1258,In_1411);
nand U90 (N_90,In_933,In_2448);
or U91 (N_91,In_2218,In_2263);
nand U92 (N_92,In_268,In_235);
nor U93 (N_93,In_1181,In_923);
nand U94 (N_94,In_2130,In_2428);
xor U95 (N_95,In_1712,In_285);
or U96 (N_96,In_783,In_510);
and U97 (N_97,In_1482,In_663);
nor U98 (N_98,In_1842,In_2029);
and U99 (N_99,In_1036,In_2392);
and U100 (N_100,In_1327,In_142);
nor U101 (N_101,In_1833,In_1422);
xnor U102 (N_102,In_1974,In_1885);
and U103 (N_103,In_1320,In_1063);
nand U104 (N_104,In_705,In_1156);
xor U105 (N_105,In_1371,In_206);
xnor U106 (N_106,In_883,In_2198);
xor U107 (N_107,In_2000,In_180);
and U108 (N_108,In_1195,In_2431);
or U109 (N_109,In_1672,In_2133);
nor U110 (N_110,In_353,In_694);
nor U111 (N_111,In_1172,In_280);
or U112 (N_112,In_955,In_1394);
and U113 (N_113,In_1428,In_1033);
nor U114 (N_114,In_1877,In_2320);
and U115 (N_115,In_1242,In_2264);
nand U116 (N_116,In_1090,In_1682);
nor U117 (N_117,In_1152,In_762);
nand U118 (N_118,In_2056,In_1103);
nand U119 (N_119,In_1361,In_2229);
nand U120 (N_120,In_1714,In_2027);
or U121 (N_121,In_789,In_730);
or U122 (N_122,In_14,In_1399);
nand U123 (N_123,In_330,In_1284);
and U124 (N_124,In_748,In_102);
or U125 (N_125,In_1416,In_556);
or U126 (N_126,In_506,In_1688);
or U127 (N_127,In_2397,In_1316);
and U128 (N_128,In_1933,In_1706);
or U129 (N_129,In_2197,In_807);
and U130 (N_130,In_1778,In_1585);
and U131 (N_131,In_1654,In_415);
nand U132 (N_132,In_1743,In_2463);
and U133 (N_133,In_967,In_1818);
and U134 (N_134,In_1802,In_1657);
nand U135 (N_135,In_2083,In_421);
xnor U136 (N_136,In_1012,In_1346);
or U137 (N_137,In_1465,In_2175);
xnor U138 (N_138,In_2118,In_1696);
and U139 (N_139,In_975,In_769);
xnor U140 (N_140,In_1574,In_114);
xnor U141 (N_141,In_781,In_1081);
nor U142 (N_142,In_1563,In_1961);
nand U143 (N_143,In_413,In_1832);
xnor U144 (N_144,In_2114,In_1190);
and U145 (N_145,In_638,In_1849);
or U146 (N_146,In_794,In_560);
xor U147 (N_147,In_44,In_743);
and U148 (N_148,In_2154,In_2340);
xnor U149 (N_149,In_227,In_2273);
xnor U150 (N_150,In_574,In_270);
nand U151 (N_151,In_2098,In_1000);
nor U152 (N_152,In_516,In_2184);
or U153 (N_153,In_1660,In_1835);
or U154 (N_154,In_1729,In_579);
and U155 (N_155,In_222,In_2212);
nand U156 (N_156,In_444,In_501);
xor U157 (N_157,In_1113,In_1203);
nor U158 (N_158,In_1836,In_2240);
and U159 (N_159,In_545,In_2410);
or U160 (N_160,In_866,In_193);
or U161 (N_161,In_1597,In_2244);
nand U162 (N_162,In_2077,In_2116);
or U163 (N_163,In_1377,In_1115);
nand U164 (N_164,In_1546,In_766);
or U165 (N_165,In_575,In_260);
nand U166 (N_166,In_332,In_1793);
nor U167 (N_167,In_1853,In_2477);
nor U168 (N_168,In_18,In_1698);
xnor U169 (N_169,In_1412,In_198);
and U170 (N_170,In_1487,In_348);
or U171 (N_171,In_0,In_755);
xnor U172 (N_172,In_1167,In_1363);
nor U173 (N_173,In_239,In_1993);
nor U174 (N_174,In_1898,In_1247);
nor U175 (N_175,In_2251,In_1904);
nor U176 (N_176,In_2443,In_930);
xnor U177 (N_177,In_2290,In_1104);
or U178 (N_178,In_988,In_89);
or U179 (N_179,In_785,In_1165);
and U180 (N_180,In_2360,In_118);
or U181 (N_181,In_91,In_1700);
nand U182 (N_182,In_1498,In_850);
xor U183 (N_183,In_1689,In_2188);
and U184 (N_184,In_643,In_1298);
and U185 (N_185,In_1248,In_2282);
nor U186 (N_186,In_1583,In_1338);
or U187 (N_187,In_1568,In_1668);
nor U188 (N_188,In_255,In_1274);
xnor U189 (N_189,In_2079,In_57);
and U190 (N_190,In_2007,In_863);
nand U191 (N_191,In_202,In_1582);
xor U192 (N_192,In_1548,In_1021);
nand U193 (N_193,In_761,In_488);
xor U194 (N_194,In_1945,In_346);
nand U195 (N_195,In_1356,In_1647);
or U196 (N_196,In_1079,In_290);
or U197 (N_197,In_2209,In_2484);
and U198 (N_198,In_284,In_271);
nor U199 (N_199,In_633,In_1116);
nand U200 (N_200,In_474,In_476);
or U201 (N_201,In_2446,In_986);
or U202 (N_202,In_1854,In_90);
nand U203 (N_203,In_2194,In_559);
nand U204 (N_204,In_9,In_2429);
xnor U205 (N_205,In_1687,In_902);
nand U206 (N_206,In_1524,In_962);
xor U207 (N_207,In_2037,In_234);
nand U208 (N_208,In_2139,In_1572);
nor U209 (N_209,In_1642,In_1928);
xor U210 (N_210,In_1321,In_1757);
xor U211 (N_211,In_645,In_660);
and U212 (N_212,In_1137,In_67);
nor U213 (N_213,In_2049,In_2310);
or U214 (N_214,In_2286,In_937);
and U215 (N_215,In_880,In_279);
and U216 (N_216,In_1086,In_2461);
xnor U217 (N_217,In_1463,In_1472);
nor U218 (N_218,In_151,In_786);
xnor U219 (N_219,In_165,In_1245);
xnor U220 (N_220,In_1900,In_2164);
nor U221 (N_221,In_735,In_893);
nand U222 (N_222,In_2199,In_313);
and U223 (N_223,In_1173,In_1906);
xnor U224 (N_224,In_306,In_2186);
or U225 (N_225,In_821,In_957);
nand U226 (N_226,In_511,In_1470);
and U227 (N_227,In_801,In_3);
nand U228 (N_228,In_1932,In_1008);
or U229 (N_229,In_2412,In_1624);
or U230 (N_230,In_185,In_544);
or U231 (N_231,In_223,In_1127);
nor U232 (N_232,In_329,In_1652);
and U233 (N_233,In_2277,In_1171);
nand U234 (N_234,In_523,In_721);
and U235 (N_235,In_2124,In_2126);
or U236 (N_236,In_363,In_2071);
or U237 (N_237,In_2211,In_812);
or U238 (N_238,In_434,In_2457);
and U239 (N_239,In_195,In_2163);
xor U240 (N_240,In_2024,In_2304);
xor U241 (N_241,In_1019,In_210);
nor U242 (N_242,In_6,In_1440);
nor U243 (N_243,In_1299,In_289);
nand U244 (N_244,In_205,In_661);
nand U245 (N_245,In_1351,In_1791);
nand U246 (N_246,In_1359,In_1307);
nand U247 (N_247,In_567,In_1522);
xor U248 (N_248,In_1114,In_321);
nor U249 (N_249,In_1882,In_2140);
nand U250 (N_250,In_108,In_1119);
nand U251 (N_251,In_266,N_106);
or U252 (N_252,In_228,In_1414);
or U253 (N_253,In_628,In_588);
nand U254 (N_254,In_16,In_867);
or U255 (N_255,N_137,In_20);
nand U256 (N_256,In_128,In_2216);
or U257 (N_257,In_602,In_1985);
nor U258 (N_258,In_1003,N_98);
and U259 (N_259,N_40,In_1725);
and U260 (N_260,In_2131,In_310);
and U261 (N_261,In_912,In_1051);
nand U262 (N_262,In_467,In_41);
or U263 (N_263,In_281,In_133);
and U264 (N_264,In_194,In_1141);
nor U265 (N_265,In_848,In_2308);
xnor U266 (N_266,In_1231,In_534);
and U267 (N_267,In_466,N_169);
xnor U268 (N_268,In_928,N_126);
nor U269 (N_269,In_1014,In_1294);
xnor U270 (N_270,In_857,In_824);
or U271 (N_271,In_2398,In_124);
nand U272 (N_272,N_194,In_2400);
and U273 (N_273,In_669,In_888);
and U274 (N_274,In_1558,In_2193);
xnor U275 (N_275,In_2318,In_518);
nand U276 (N_276,In_300,In_331);
nor U277 (N_277,In_787,In_293);
and U278 (N_278,In_2176,In_359);
and U279 (N_279,In_1333,In_1774);
and U280 (N_280,N_187,In_2353);
nor U281 (N_281,In_1212,N_138);
nand U282 (N_282,In_2348,In_1756);
or U283 (N_283,In_657,In_1352);
or U284 (N_284,In_1035,N_154);
and U285 (N_285,In_960,In_2028);
or U286 (N_286,In_1823,In_2380);
nand U287 (N_287,In_1002,N_201);
or U288 (N_288,In_1661,In_1500);
or U289 (N_289,In_1604,In_1755);
xnor U290 (N_290,In_606,In_50);
or U291 (N_291,In_480,In_297);
nand U292 (N_292,In_927,In_2493);
xnor U293 (N_293,In_2479,In_490);
xnor U294 (N_294,In_1809,N_78);
nor U295 (N_295,In_1028,In_1754);
and U296 (N_296,In_569,N_12);
or U297 (N_297,In_1154,In_681);
nand U298 (N_298,In_1565,In_1058);
nor U299 (N_299,N_71,In_1291);
nand U300 (N_300,In_725,In_2052);
xor U301 (N_301,N_96,In_1494);
nand U302 (N_302,In_2107,In_2325);
nor U303 (N_303,In_1088,In_2148);
xor U304 (N_304,In_1145,In_1770);
nand U305 (N_305,In_1735,In_1188);
or U306 (N_306,In_1375,In_1053);
nor U307 (N_307,In_1655,In_1140);
or U308 (N_308,In_1233,In_11);
nand U309 (N_309,In_238,In_1895);
and U310 (N_310,In_1719,In_527);
and U311 (N_311,N_7,In_489);
nand U312 (N_312,In_483,In_803);
and U313 (N_313,In_430,In_1753);
or U314 (N_314,In_356,In_684);
and U315 (N_315,In_604,In_1365);
and U316 (N_316,In_1252,In_315);
xor U317 (N_317,In_1705,In_951);
and U318 (N_318,In_1250,In_1787);
and U319 (N_319,In_1409,N_55);
and U320 (N_320,In_2364,In_771);
nor U321 (N_321,In_191,In_935);
xnor U322 (N_322,In_345,In_1160);
xnor U323 (N_323,In_388,In_1343);
nor U324 (N_324,In_585,In_833);
xor U325 (N_325,In_1599,In_1677);
and U326 (N_326,In_1975,In_2303);
nand U327 (N_327,In_759,In_1354);
and U328 (N_328,In_1221,In_2171);
nand U329 (N_329,In_779,In_1742);
xnor U330 (N_330,In_115,In_1550);
nand U331 (N_331,In_2091,In_712);
xor U332 (N_332,In_2437,In_1039);
nand U333 (N_333,In_2143,In_1966);
xnor U334 (N_334,In_2166,In_1224);
xor U335 (N_335,In_966,In_1177);
nor U336 (N_336,In_1612,In_891);
nor U337 (N_337,N_46,In_145);
nor U338 (N_338,In_1983,In_1573);
xor U339 (N_339,In_581,In_1082);
xor U340 (N_340,In_1942,In_2178);
nand U341 (N_341,In_1074,In_2357);
and U342 (N_342,In_865,In_819);
nor U343 (N_343,In_2088,In_675);
nand U344 (N_344,N_120,In_237);
nand U345 (N_345,N_76,In_2096);
and U346 (N_346,In_2368,In_1246);
nor U347 (N_347,In_2059,In_1857);
nand U348 (N_348,In_1484,In_418);
nor U349 (N_349,In_914,In_478);
and U350 (N_350,In_2468,In_1503);
and U351 (N_351,In_109,In_2135);
and U352 (N_352,In_2250,In_1444);
xnor U353 (N_353,In_189,In_619);
nand U354 (N_354,In_1551,In_1795);
nand U355 (N_355,In_1138,N_206);
and U356 (N_356,N_94,In_945);
or U357 (N_357,In_744,In_307);
nor U358 (N_358,In_1037,N_22);
nor U359 (N_359,In_1779,In_1976);
nor U360 (N_360,In_1232,N_37);
xor U361 (N_361,In_382,In_71);
xor U362 (N_362,N_178,In_1417);
or U363 (N_363,In_150,In_742);
nand U364 (N_364,In_910,In_55);
or U365 (N_365,In_2406,N_229);
nor U366 (N_366,In_259,In_393);
nand U367 (N_367,In_1870,In_507);
or U368 (N_368,N_70,In_646);
nand U369 (N_369,In_1916,In_2394);
nand U370 (N_370,In_2414,In_1471);
nand U371 (N_371,In_1151,In_2057);
and U372 (N_372,In_34,In_767);
nor U373 (N_373,In_827,N_16);
xor U374 (N_374,In_1117,In_887);
nor U375 (N_375,In_1027,In_547);
or U376 (N_376,In_834,In_2243);
or U377 (N_377,In_2356,N_100);
nand U378 (N_378,In_1135,In_1270);
or U379 (N_379,In_873,In_667);
xor U380 (N_380,In_1388,In_2201);
xor U381 (N_381,In_692,In_989);
and U382 (N_382,In_1531,In_773);
nand U383 (N_383,N_4,In_2352);
or U384 (N_384,In_1201,In_2111);
nand U385 (N_385,In_2345,In_1424);
nor U386 (N_386,In_424,In_899);
or U387 (N_387,In_199,In_1600);
or U388 (N_388,In_2046,In_944);
and U389 (N_389,In_861,N_147);
nor U390 (N_390,In_31,In_2097);
or U391 (N_391,In_521,In_814);
or U392 (N_392,In_1562,In_983);
xnor U393 (N_393,In_1429,In_1319);
xnor U394 (N_394,In_896,In_2104);
nand U395 (N_395,In_216,In_561);
nor U396 (N_396,In_2342,N_162);
and U397 (N_397,In_1785,N_80);
or U398 (N_398,In_1056,In_1474);
nor U399 (N_399,In_997,In_2346);
nor U400 (N_400,In_1326,In_813);
nand U401 (N_401,In_2092,In_1461);
or U402 (N_402,In_1289,In_2339);
and U403 (N_403,In_425,N_168);
or U404 (N_404,N_143,In_2256);
nor U405 (N_405,In_1641,In_1495);
xor U406 (N_406,In_1944,In_2441);
nor U407 (N_407,In_760,N_196);
or U408 (N_408,In_2039,In_155);
nand U409 (N_409,In_2061,In_978);
nand U410 (N_410,In_1089,In_1534);
xnor U411 (N_411,In_1971,N_153);
nor U412 (N_412,In_2121,In_1784);
or U413 (N_413,In_758,In_378);
or U414 (N_414,In_1030,N_79);
nor U415 (N_415,In_452,In_2288);
nand U416 (N_416,In_1805,In_1616);
xnor U417 (N_417,In_157,In_550);
or U418 (N_418,In_1889,In_2271);
and U419 (N_419,In_146,In_267);
nor U420 (N_420,In_2010,In_2294);
and U421 (N_421,In_1369,In_1048);
xor U422 (N_422,N_179,In_190);
xnor U423 (N_423,In_475,In_648);
or U424 (N_424,In_2074,In_1234);
nand U425 (N_425,In_810,In_152);
nor U426 (N_426,N_160,In_656);
and U427 (N_427,In_582,In_1329);
nor U428 (N_428,In_1178,N_11);
and U429 (N_429,In_2204,In_1230);
nor U430 (N_430,In_984,In_1507);
xnor U431 (N_431,In_603,In_183);
or U432 (N_432,In_1771,In_780);
xnor U433 (N_433,In_362,In_1249);
nor U434 (N_434,In_974,In_2322);
and U435 (N_435,N_54,In_1309);
and U436 (N_436,In_1383,In_1032);
nor U437 (N_437,In_379,In_1106);
or U438 (N_438,In_1179,In_2090);
nand U439 (N_439,In_2281,In_2372);
nor U440 (N_440,In_1728,In_1584);
and U441 (N_441,In_727,In_1925);
nor U442 (N_442,N_184,In_950);
or U443 (N_443,In_1914,In_1451);
and U444 (N_444,In_1391,In_2291);
or U445 (N_445,In_472,In_2376);
and U446 (N_446,In_457,In_2158);
and U447 (N_447,In_412,In_1239);
nor U448 (N_448,In_2362,N_66);
nor U449 (N_449,In_1713,In_2344);
nand U450 (N_450,In_1175,In_616);
nand U451 (N_451,In_1290,In_1168);
nor U452 (N_452,In_808,N_210);
nor U453 (N_453,In_77,In_1968);
nand U454 (N_454,In_217,In_2230);
nor U455 (N_455,In_765,In_508);
nor U456 (N_456,In_1007,In_495);
nand U457 (N_457,In_1038,In_1013);
nor U458 (N_458,In_1197,In_1701);
or U459 (N_459,N_18,In_1595);
or U460 (N_460,In_447,In_59);
or U461 (N_461,In_2045,N_205);
and U462 (N_462,In_221,In_5);
nand U463 (N_463,In_1166,N_202);
or U464 (N_464,N_75,N_69);
nand U465 (N_465,In_1332,In_1481);
nand U466 (N_466,In_2050,In_344);
nor U467 (N_467,In_2404,In_2048);
nor U468 (N_468,In_584,In_941);
xor U469 (N_469,In_795,In_2080);
and U470 (N_470,In_320,In_806);
xnor U471 (N_471,In_252,In_485);
nor U472 (N_472,In_2361,N_144);
nand U473 (N_473,In_1614,In_2167);
xnor U474 (N_474,In_493,In_654);
xnor U475 (N_475,N_36,In_1917);
or U476 (N_476,In_2274,In_1681);
nand U477 (N_477,In_2269,In_392);
xor U478 (N_478,In_2306,In_683);
xor U479 (N_479,N_49,In_187);
xnor U480 (N_480,In_361,In_1992);
and U481 (N_481,In_441,In_125);
nand U482 (N_482,In_1684,In_1257);
nor U483 (N_483,N_239,In_1650);
nand U484 (N_484,In_982,In_676);
or U485 (N_485,In_1436,In_971);
or U486 (N_486,In_86,In_845);
nand U487 (N_487,In_1840,In_428);
xor U488 (N_488,In_1202,In_2227);
nor U489 (N_489,In_254,In_815);
nor U490 (N_490,In_1490,In_246);
nand U491 (N_491,In_1220,In_1772);
xor U492 (N_492,In_1006,In_12);
and U493 (N_493,In_101,In_82);
or U494 (N_494,In_1293,N_116);
nor U495 (N_495,In_2490,In_2424);
xor U496 (N_496,In_1480,In_1827);
nor U497 (N_497,In_2261,In_182);
nand U498 (N_498,In_1302,In_666);
nand U499 (N_499,In_1355,In_134);
or U500 (N_500,In_1042,In_1609);
and U501 (N_501,N_83,In_1519);
nand U502 (N_502,In_1970,In_1552);
or U503 (N_503,In_994,In_470);
and U504 (N_504,N_339,In_583);
or U505 (N_505,In_167,N_414);
nand U506 (N_506,N_0,In_796);
nand U507 (N_507,N_473,In_1200);
xor U508 (N_508,In_741,In_1846);
nand U509 (N_509,N_407,In_1123);
xor U510 (N_510,N_447,In_405);
xor U511 (N_511,N_217,In_1732);
xor U512 (N_512,In_2179,In_2076);
xnor U513 (N_513,In_1887,In_1702);
nand U514 (N_514,In_2239,In_207);
nor U515 (N_515,In_1005,In_906);
xnor U516 (N_516,In_394,In_835);
and U517 (N_517,In_1398,In_898);
nand U518 (N_518,N_276,N_344);
nor U519 (N_519,N_499,In_1378);
xor U520 (N_520,In_1996,N_365);
xor U521 (N_521,In_431,In_1973);
nor U522 (N_522,In_2180,In_302);
xor U523 (N_523,In_2242,In_112);
or U524 (N_524,In_203,In_1415);
nor U525 (N_525,In_922,N_212);
or U526 (N_526,In_969,N_17);
or U527 (N_527,In_1344,In_243);
xnor U528 (N_528,In_2129,In_1357);
or U529 (N_529,In_110,In_1733);
or U530 (N_530,In_1253,In_1911);
nor U531 (N_531,In_2101,In_2381);
nand U532 (N_532,In_1538,In_129);
and U533 (N_533,In_63,In_903);
or U534 (N_534,In_2385,N_376);
and U535 (N_535,In_697,In_341);
xor U536 (N_536,In_1566,N_39);
nor U537 (N_537,N_309,N_431);
nand U538 (N_538,In_2040,In_1697);
xnor U539 (N_539,In_1781,In_1479);
nand U540 (N_540,N_332,In_1810);
xnor U541 (N_541,In_2301,N_10);
and U542 (N_542,In_1467,In_655);
xor U543 (N_543,In_1629,N_288);
xor U544 (N_544,In_2231,In_2150);
nand U545 (N_545,N_232,In_2287);
or U546 (N_546,In_1392,In_463);
nor U547 (N_547,In_263,In_1129);
xor U548 (N_548,In_1556,In_113);
or U549 (N_549,In_1536,N_273);
and U550 (N_550,In_1459,In_695);
and U551 (N_551,In_1666,In_2036);
xnor U552 (N_552,In_1589,In_737);
or U553 (N_553,In_700,In_251);
xor U554 (N_554,N_275,In_445);
nand U555 (N_555,In_2120,N_28);
nand U556 (N_556,N_242,In_2100);
nand U557 (N_557,In_640,In_1653);
xnor U558 (N_558,N_404,In_921);
or U559 (N_559,In_2481,N_384);
nand U560 (N_560,N_451,In_1972);
and U561 (N_561,In_670,N_263);
nor U562 (N_562,In_658,In_1737);
and U563 (N_563,In_1026,N_334);
nand U564 (N_564,In_2495,In_621);
or U565 (N_565,In_1844,In_719);
xnor U566 (N_566,In_1856,In_662);
or U567 (N_567,In_1523,N_77);
xor U568 (N_568,In_2054,In_2349);
and U569 (N_569,N_383,In_634);
and U570 (N_570,In_2145,In_736);
nor U571 (N_571,In_1069,In_2241);
and U572 (N_572,In_439,In_1073);
nor U573 (N_573,N_481,In_1822);
nand U574 (N_574,In_2203,N_397);
xor U575 (N_575,N_390,In_365);
nor U576 (N_576,In_104,In_548);
xor U577 (N_577,In_525,N_449);
xnor U578 (N_578,In_717,In_947);
and U579 (N_579,In_2138,In_87);
and U580 (N_580,In_625,In_1094);
and U581 (N_581,In_1532,In_533);
xor U582 (N_582,N_256,In_2359);
nor U583 (N_583,N_238,In_2375);
or U584 (N_584,In_2099,In_1850);
xnor U585 (N_585,In_1869,In_120);
nor U586 (N_586,N_220,In_1518);
xor U587 (N_587,N_164,In_4);
and U588 (N_588,In_2494,In_484);
or U589 (N_589,N_349,N_424);
nor U590 (N_590,In_714,N_409);
or U591 (N_591,N_459,N_361);
nor U592 (N_592,In_2109,In_2034);
or U593 (N_593,In_2245,In_2436);
and U594 (N_594,N_302,N_422);
or U595 (N_595,In_872,In_1297);
and U596 (N_596,In_1460,In_554);
nor U597 (N_597,In_1193,In_2365);
or U598 (N_598,In_2326,N_114);
nand U599 (N_599,In_376,In_1096);
or U600 (N_600,In_414,In_1268);
xnor U601 (N_601,In_287,In_2078);
xnor U602 (N_602,In_2316,In_1269);
or U603 (N_603,In_1111,In_1385);
and U604 (N_604,In_710,In_715);
nor U605 (N_605,In_2260,In_1847);
nor U606 (N_606,In_105,N_13);
nor U607 (N_607,In_1279,In_600);
nand U608 (N_608,In_276,In_1752);
nor U609 (N_609,In_1943,In_116);
or U610 (N_610,In_2319,N_243);
nand U611 (N_611,In_1662,In_1124);
or U612 (N_612,N_156,In_1905);
nand U613 (N_613,N_146,In_1594);
nand U614 (N_614,In_1206,In_626);
or U615 (N_615,In_2093,In_56);
nor U616 (N_616,In_1324,In_2051);
xor U617 (N_617,In_1893,N_483);
xnor U618 (N_618,In_2366,In_818);
nand U619 (N_619,In_689,In_541);
nand U620 (N_620,N_151,In_333);
or U621 (N_621,N_498,In_2396);
nand U622 (N_622,In_653,N_127);
and U623 (N_623,N_161,In_1308);
nand U624 (N_624,In_2307,In_1271);
or U625 (N_625,N_343,N_29);
or U626 (N_626,In_924,In_2152);
or U627 (N_627,In_1093,In_1376);
and U628 (N_628,In_855,In_1746);
or U629 (N_629,In_1204,In_21);
and U630 (N_630,In_2476,In_422);
xor U631 (N_631,In_734,In_925);
nor U632 (N_632,In_1121,N_199);
xnor U633 (N_633,In_486,In_1267);
and U634 (N_634,In_2491,In_411);
nor U635 (N_635,In_1617,N_461);
and U636 (N_636,In_980,In_860);
nand U637 (N_637,In_384,In_512);
and U638 (N_638,In_324,In_557);
nand U639 (N_639,In_1517,In_612);
and U640 (N_640,In_2215,In_578);
or U641 (N_641,In_745,N_59);
xnor U642 (N_642,In_423,In_1330);
xnor U643 (N_643,In_1978,N_307);
or U644 (N_644,In_291,In_158);
nor U645 (N_645,In_1300,In_1387);
xnor U646 (N_646,N_323,N_214);
or U647 (N_647,N_181,In_1816);
nor U648 (N_648,In_2247,In_1790);
or U649 (N_649,In_513,N_56);
nor U650 (N_650,N_150,In_2022);
or U651 (N_651,In_2460,In_369);
nor U652 (N_652,In_1717,In_8);
nand U653 (N_653,In_433,In_2254);
xor U654 (N_654,N_312,In_40);
xor U655 (N_655,In_389,In_2017);
xor U656 (N_656,N_482,In_2469);
xor U657 (N_657,In_1180,N_441);
xnor U658 (N_658,In_2489,In_2295);
nand U659 (N_659,In_1379,In_1184);
xnor U660 (N_660,N_231,In_1564);
nor U661 (N_661,In_130,In_1613);
or U662 (N_662,In_862,In_851);
or U663 (N_663,In_282,N_108);
nand U664 (N_664,In_1,In_2030);
xor U665 (N_665,In_1939,In_2136);
xnor U666 (N_666,In_959,In_1466);
xor U667 (N_667,In_1512,In_163);
nand U668 (N_668,In_305,In_2329);
and U669 (N_669,In_2492,In_2105);
and U670 (N_670,In_1723,N_367);
or U671 (N_671,In_2338,In_201);
xnor U672 (N_672,N_463,In_805);
nor U673 (N_673,In_2005,In_609);
xnor U674 (N_674,In_2082,In_127);
nor U675 (N_675,In_635,N_1);
and U676 (N_676,In_2207,In_776);
xnor U677 (N_677,In_1703,In_1229);
nand U678 (N_678,In_782,In_1948);
xnor U679 (N_679,In_856,N_381);
or U680 (N_680,N_313,In_357);
nand U681 (N_681,In_240,In_1087);
or U682 (N_682,In_551,In_1150);
or U683 (N_683,In_746,In_674);
nand U684 (N_684,In_2432,N_225);
nor U685 (N_685,In_519,In_391);
nor U686 (N_686,In_1159,In_250);
nor U687 (N_687,In_1867,In_335);
and U688 (N_688,In_78,N_111);
xor U689 (N_689,In_1699,N_62);
nor U690 (N_690,In_1813,In_1601);
xnor U691 (N_691,In_2095,In_2084);
xnor U692 (N_692,N_109,In_2403);
nand U693 (N_693,In_2069,In_1786);
xnor U694 (N_694,In_852,N_480);
and U695 (N_695,In_911,In_2472);
xnor U696 (N_696,In_2214,In_990);
or U697 (N_697,In_2248,In_1132);
and U698 (N_698,In_326,In_1575);
or U699 (N_699,In_2374,In_2435);
nand U700 (N_700,In_775,In_1963);
nor U701 (N_701,In_2081,In_2454);
xor U702 (N_702,In_631,N_466);
nor U703 (N_703,N_191,N_115);
nor U704 (N_704,In_2272,N_23);
and U705 (N_705,In_639,In_1432);
xor U706 (N_706,In_2317,In_837);
xor U707 (N_707,In_897,In_1632);
and U708 (N_708,N_68,In_278);
and U709 (N_709,N_311,In_1683);
xor U710 (N_710,N_97,In_99);
nor U711 (N_711,In_909,In_401);
or U712 (N_712,In_218,In_1744);
and U713 (N_713,N_378,In_2434);
or U714 (N_714,N_284,In_1255);
or U715 (N_715,In_1947,In_2311);
nand U716 (N_716,In_2213,In_1238);
nor U717 (N_717,In_1381,N_400);
or U718 (N_718,In_716,In_342);
nor U719 (N_719,In_528,N_155);
xnor U720 (N_720,In_28,In_1881);
and U721 (N_721,In_1402,In_1533);
nand U722 (N_722,In_1864,N_478);
or U723 (N_723,In_1364,In_1964);
xnor U724 (N_724,N_357,N_208);
and U725 (N_725,In_1143,In_2337);
xnor U726 (N_726,N_300,In_1986);
and U727 (N_727,N_280,In_1080);
nor U728 (N_728,In_247,In_665);
or U729 (N_729,In_1800,N_380);
and U730 (N_730,In_1210,In_750);
nand U731 (N_731,In_1695,In_2347);
xnor U732 (N_732,In_532,In_823);
and U733 (N_733,In_514,In_1310);
xor U734 (N_734,In_35,In_1049);
or U735 (N_735,In_1969,In_2146);
or U736 (N_736,In_137,In_1676);
and U737 (N_737,N_457,In_1041);
nor U738 (N_738,In_1240,In_479);
and U739 (N_739,In_2257,In_644);
nor U740 (N_740,N_286,In_2399);
nand U741 (N_741,In_241,In_409);
or U742 (N_742,N_436,In_961);
or U743 (N_743,In_905,In_2471);
or U744 (N_744,In_170,N_306);
nor U745 (N_745,In_1215,In_1674);
xnor U746 (N_746,In_1952,In_311);
and U747 (N_747,In_309,In_1883);
nor U748 (N_748,In_29,In_1506);
and U749 (N_749,In_52,In_2470);
nand U750 (N_750,In_555,N_412);
nor U751 (N_751,N_554,N_642);
and U752 (N_752,In_1052,In_680);
nand U753 (N_753,N_125,In_482);
nand U754 (N_754,N_166,In_166);
nor U755 (N_755,N_148,In_2462);
nor U756 (N_756,In_1852,In_1426);
nand U757 (N_757,N_602,In_1325);
nand U758 (N_758,N_614,In_1286);
nor U759 (N_759,N_465,N_450);
xnor U760 (N_760,In_1055,In_601);
nand U761 (N_761,N_656,N_625);
nor U762 (N_762,In_487,In_1903);
nand U763 (N_763,In_598,In_178);
or U764 (N_764,In_1669,In_352);
nand U765 (N_765,In_711,In_531);
xor U766 (N_766,In_1442,N_24);
nand U767 (N_767,In_2234,N_488);
or U768 (N_768,In_402,In_2015);
nand U769 (N_769,In_399,In_48);
nand U770 (N_770,N_277,In_2085);
nand U771 (N_771,In_2328,In_2386);
and U772 (N_772,N_45,N_686);
or U773 (N_773,In_417,In_1559);
xnor U774 (N_774,In_1236,In_1958);
or U775 (N_775,In_442,N_30);
xnor U776 (N_776,In_1261,In_93);
or U777 (N_777,In_2191,In_32);
or U778 (N_778,In_1693,N_446);
and U779 (N_779,N_289,In_764);
or U780 (N_780,In_1148,In_319);
xnor U781 (N_781,N_101,N_247);
nor U782 (N_782,N_224,In_1278);
and U783 (N_783,In_1819,In_2486);
and U784 (N_784,In_1886,N_335);
nor U785 (N_785,In_798,In_2447);
xor U786 (N_786,N_730,In_973);
and U787 (N_787,In_1667,N_437);
and U788 (N_788,In_2354,In_826);
or U789 (N_789,N_198,N_525);
nor U790 (N_790,N_226,In_869);
nand U791 (N_791,In_1776,In_538);
or U792 (N_792,In_304,In_726);
xor U793 (N_793,N_95,In_2210);
and U794 (N_794,In_97,In_1001);
and U795 (N_795,In_2012,In_1191);
and U796 (N_796,N_74,N_649);
or U797 (N_797,In_1644,N_132);
nand U798 (N_798,N_105,In_593);
and U799 (N_799,In_1128,In_1303);
or U800 (N_800,N_573,In_1636);
xnor U801 (N_801,In_977,In_1350);
nand U802 (N_802,In_184,In_2497);
xnor U803 (N_803,In_2020,In_2003);
nand U804 (N_804,In_1029,In_1704);
nor U805 (N_805,N_558,In_1010);
nor U806 (N_806,In_2482,In_607);
nand U807 (N_807,In_2043,In_846);
nor U808 (N_808,In_763,N_139);
xnor U809 (N_809,In_1446,In_1912);
nor U810 (N_810,In_1478,In_2363);
nand U811 (N_811,N_662,In_1349);
and U812 (N_812,In_979,In_53);
xnor U813 (N_813,N_467,N_269);
nor U814 (N_814,N_748,In_934);
or U815 (N_815,In_1543,In_1277);
xor U816 (N_816,In_1623,N_85);
and U817 (N_817,In_103,In_536);
or U818 (N_818,In_1711,In_832);
and U819 (N_819,N_703,In_261);
and U820 (N_820,In_1894,N_395);
nor U821 (N_821,In_790,In_1527);
nor U822 (N_822,N_699,N_657);
xnor U823 (N_823,In_1256,In_2483);
or U824 (N_824,In_1301,In_2169);
xor U825 (N_825,In_84,In_408);
xnor U826 (N_826,In_295,N_670);
and U827 (N_827,N_103,In_1855);
nand U828 (N_828,In_1722,In_1083);
and U829 (N_829,N_658,In_2343);
and U830 (N_830,N_274,In_739);
xnor U831 (N_831,In_2474,In_1061);
and U832 (N_832,In_1384,In_349);
or U833 (N_833,N_597,In_334);
or U834 (N_834,N_611,In_753);
or U835 (N_835,N_543,N_333);
xor U836 (N_836,In_1122,N_134);
xor U837 (N_837,In_46,In_1004);
nand U838 (N_838,N_676,In_1118);
or U839 (N_839,In_552,N_713);
nor U840 (N_840,N_705,N_310);
and U841 (N_841,In_907,In_938);
nand U842 (N_842,In_2006,N_486);
nand U843 (N_843,N_494,In_1227);
nor U844 (N_844,N_296,In_2485);
nand U845 (N_845,In_793,N_113);
nand U846 (N_846,In_1439,In_1112);
or U847 (N_847,In_2224,In_398);
nand U848 (N_848,N_423,In_2226);
xnor U849 (N_849,In_1637,N_324);
nor U850 (N_850,N_734,In_2419);
nand U851 (N_851,N_345,In_2021);
and U852 (N_852,In_2430,N_673);
nor U853 (N_853,In_1627,N_427);
nor U854 (N_854,In_688,In_2103);
or U855 (N_855,In_1608,N_580);
or U856 (N_856,N_67,In_42);
xor U857 (N_857,In_2159,In_1464);
nor U858 (N_858,In_740,In_225);
nand U859 (N_859,In_94,In_1921);
nor U860 (N_860,In_757,In_854);
and U861 (N_861,N_725,In_2065);
and U862 (N_862,N_632,N_544);
or U863 (N_863,N_43,In_995);
or U864 (N_864,In_1454,N_399);
xor U865 (N_865,N_245,In_1578);
or U866 (N_866,In_1673,In_62);
nand U867 (N_867,N_244,In_708);
xor U868 (N_868,In_171,In_1062);
and U869 (N_869,In_840,In_629);
and U870 (N_870,In_1890,N_351);
xor U871 (N_871,In_80,In_1946);
nand U872 (N_872,In_1995,In_2123);
xor U873 (N_873,In_1892,In_549);
nor U874 (N_874,N_643,In_991);
xnor U875 (N_875,In_1865,N_599);
xnor U876 (N_876,In_2297,N_123);
or U877 (N_877,In_778,In_1285);
and U878 (N_878,In_620,In_1401);
nand U879 (N_879,N_157,N_619);
and U880 (N_880,In_1456,In_1937);
nor U881 (N_881,In_1011,N_698);
xor U882 (N_882,N_413,N_552);
nand U883 (N_883,In_530,In_2122);
nand U884 (N_884,In_2384,In_1433);
nand U885 (N_885,In_54,N_696);
nor U886 (N_886,In_2174,In_1282);
nand U887 (N_887,In_2433,In_868);
nor U888 (N_888,In_135,In_1209);
and U889 (N_889,N_485,In_1315);
nor U890 (N_890,In_2382,In_733);
and U891 (N_891,N_561,N_258);
nand U892 (N_892,N_285,In_1710);
and U893 (N_893,N_316,In_1980);
nor U894 (N_894,In_1406,In_111);
xnor U895 (N_895,In_1929,N_320);
or U896 (N_896,In_1280,In_570);
nand U897 (N_897,N_726,N_557);
or U898 (N_898,In_1544,In_1765);
xnor U899 (N_899,N_476,N_31);
nand U900 (N_900,In_2292,In_1499);
nor U901 (N_901,In_682,In_881);
xor U902 (N_902,In_2449,N_608);
nor U903 (N_903,In_1362,In_1084);
or U904 (N_904,In_299,N_34);
nor U905 (N_905,In_2302,In_2422);
nand U906 (N_906,N_603,N_336);
or U907 (N_907,In_1875,In_2418);
and U908 (N_908,N_594,In_1782);
and U909 (N_909,In_1545,In_1453);
or U910 (N_910,In_1185,N_21);
or U911 (N_911,N_382,In_1457);
or U912 (N_912,In_1861,In_2417);
nor U913 (N_913,N_420,N_604);
nand U914 (N_914,In_366,In_2208);
nor U915 (N_915,In_502,In_2314);
and U916 (N_916,N_740,N_584);
xnor U917 (N_917,In_274,In_1934);
nor U918 (N_918,In_303,N_252);
xnor U919 (N_919,In_728,In_1016);
or U920 (N_920,In_213,In_1540);
nand U921 (N_921,In_1455,In_1108);
nand U922 (N_922,In_153,In_2456);
nor U923 (N_923,In_1157,In_1675);
nand U924 (N_924,In_1263,N_102);
nor U925 (N_925,In_1592,In_1775);
xnor U926 (N_926,In_1043,N_375);
nor U927 (N_927,N_732,N_565);
xnor U928 (N_928,N_607,In_890);
nor U929 (N_929,In_972,In_540);
xor U930 (N_930,In_226,In_1100);
xor U931 (N_931,In_256,In_61);
nor U932 (N_932,In_64,N_663);
or U933 (N_933,In_800,In_2409);
nand U934 (N_934,In_2222,N_359);
or U935 (N_935,In_2445,In_2170);
nand U936 (N_936,N_741,In_731);
nand U937 (N_937,N_610,In_1144);
nand U938 (N_938,In_1981,In_1815);
or U939 (N_939,In_407,N_523);
or U940 (N_940,In_436,In_2141);
nand U941 (N_941,In_258,N_362);
or U942 (N_942,N_355,In_1839);
or U943 (N_943,N_228,In_1192);
nand U944 (N_944,In_830,N_715);
or U945 (N_945,In_248,In_870);
or U946 (N_946,N_158,N_38);
and U947 (N_947,N_724,N_145);
and U948 (N_948,N_173,In_2004);
nand U949 (N_949,In_1908,In_871);
nand U950 (N_950,In_539,In_1560);
nor U951 (N_951,N_283,N_634);
nand U952 (N_952,In_106,N_240);
nand U953 (N_953,In_2147,N_272);
and U954 (N_954,N_235,In_713);
and U955 (N_955,In_427,N_508);
and U956 (N_956,In_1555,In_998);
nand U957 (N_957,N_301,N_72);
nand U958 (N_958,N_188,In_83);
and U959 (N_959,N_504,In_140);
nor U960 (N_960,N_556,N_321);
and U961 (N_961,N_530,In_563);
nand U962 (N_962,In_1207,N_42);
xnor U963 (N_963,N_331,In_2173);
or U964 (N_964,N_514,In_1645);
nor U965 (N_965,In_215,In_1736);
nor U966 (N_966,In_461,In_879);
and U967 (N_967,In_1761,In_1427);
xnor U968 (N_968,In_2161,N_563);
nor U969 (N_969,N_140,N_559);
and U970 (N_970,N_520,In_2267);
nand U971 (N_971,In_847,N_533);
nand U972 (N_972,In_1259,In_952);
nor U973 (N_973,In_1147,N_91);
xnor U974 (N_974,In_1235,In_1630);
nand U975 (N_975,In_1425,N_497);
nor U976 (N_976,In_592,In_1105);
nand U977 (N_977,In_169,In_2266);
and U978 (N_978,In_664,In_1602);
nand U979 (N_979,In_2458,In_964);
nand U980 (N_980,In_2467,In_492);
nand U981 (N_981,In_2183,N_667);
nand U982 (N_982,In_1715,In_249);
or U983 (N_983,In_294,In_1133);
and U984 (N_984,N_265,In_1831);
or U985 (N_985,In_864,In_802);
or U986 (N_986,In_1569,In_2205);
or U987 (N_987,In_159,In_2300);
nand U988 (N_988,In_1225,In_7);
nor U989 (N_989,N_64,In_1511);
nor U990 (N_990,In_1851,In_1824);
xnor U991 (N_991,In_1837,In_404);
nand U992 (N_992,N_503,In_2219);
nor U993 (N_993,In_1640,In_173);
nand U994 (N_994,In_141,In_1879);
nand U995 (N_995,In_449,N_492);
or U996 (N_996,In_1146,In_296);
nor U997 (N_997,In_1901,N_430);
xor U998 (N_998,N_261,N_453);
and U999 (N_999,In_844,In_231);
xor U1000 (N_1000,In_1628,In_316);
or U1001 (N_1001,In_542,In_1845);
nand U1002 (N_1002,N_974,N_903);
xnor U1003 (N_1003,In_168,N_500);
and U1004 (N_1004,In_1720,N_183);
xnor U1005 (N_1005,In_701,N_352);
xor U1006 (N_1006,In_1413,In_2451);
nand U1007 (N_1007,In_1880,N_719);
xnor U1008 (N_1008,N_26,N_562);
nand U1009 (N_1009,In_1208,N_426);
and U1010 (N_1010,N_983,N_689);
nor U1011 (N_1011,N_58,N_566);
xor U1012 (N_1012,In_419,N_405);
or U1013 (N_1013,In_1769,In_590);
nand U1014 (N_1014,N_495,In_1759);
nand U1015 (N_1015,In_931,In_829);
and U1016 (N_1016,In_1792,In_2067);
xnor U1017 (N_1017,In_1539,In_2455);
or U1018 (N_1018,In_718,N_510);
nor U1019 (N_1019,N_762,N_192);
nor U1020 (N_1020,N_363,In_1586);
xnor U1021 (N_1021,N_87,N_727);
nand U1022 (N_1022,In_1680,N_527);
xor U1023 (N_1023,N_964,N_479);
xor U1024 (N_1024,In_262,In_65);
nor U1025 (N_1025,In_72,In_462);
xnor U1026 (N_1026,In_312,N_124);
and U1027 (N_1027,N_876,In_1273);
or U1028 (N_1028,N_477,N_838);
nor U1029 (N_1029,N_775,N_353);
nor U1030 (N_1030,N_379,N_890);
nor U1031 (N_1031,N_176,N_297);
nand U1032 (N_1032,N_200,N_683);
xor U1033 (N_1033,In_1618,N_807);
nor U1034 (N_1034,In_1469,N_972);
and U1035 (N_1035,In_1542,In_1873);
nand U1036 (N_1036,In_481,In_2321);
and U1037 (N_1037,In_1334,N_165);
nand U1038 (N_1038,In_605,N_620);
and U1039 (N_1039,In_367,N_86);
nor U1040 (N_1040,In_1155,In_66);
or U1041 (N_1041,N_853,N_851);
and U1042 (N_1042,In_2018,N_325);
or U1043 (N_1043,N_170,N_856);
or U1044 (N_1044,N_84,N_955);
nor U1045 (N_1045,N_687,In_1727);
nand U1046 (N_1046,In_963,N_842);
or U1047 (N_1047,N_406,In_219);
xnor U1048 (N_1048,In_236,In_1423);
or U1049 (N_1049,N_891,In_2236);
or U1050 (N_1050,In_160,N_722);
and U1051 (N_1051,In_2332,In_1646);
nand U1052 (N_1052,N_292,In_1067);
and U1053 (N_1053,In_1395,N_710);
xor U1054 (N_1054,In_149,In_690);
nor U1055 (N_1055,N_743,N_588);
and U1056 (N_1056,N_454,In_2042);
xor U1057 (N_1057,In_2238,N_19);
and U1058 (N_1058,N_606,N_254);
or U1059 (N_1059,In_958,In_1335);
nand U1060 (N_1060,N_460,N_809);
nor U1061 (N_1061,In_92,In_831);
and U1062 (N_1062,N_402,In_81);
xnor U1063 (N_1063,In_1374,In_2094);
nand U1064 (N_1064,In_2252,N_968);
xor U1065 (N_1065,N_52,In_2355);
nand U1066 (N_1066,In_1161,In_328);
nand U1067 (N_1067,In_123,N_429);
or U1068 (N_1068,In_2452,In_679);
nor U1069 (N_1069,In_1826,N_560);
and U1070 (N_1070,In_1596,In_571);
or U1071 (N_1071,In_2313,N_299);
and U1072 (N_1072,In_916,N_763);
nor U1073 (N_1073,In_2008,N_965);
or U1074 (N_1074,In_1214,In_651);
nand U1075 (N_1075,In_143,In_1749);
nand U1076 (N_1076,N_957,In_2001);
or U1077 (N_1077,N_646,In_2087);
or U1078 (N_1078,N_308,In_2262);
and U1079 (N_1079,In_242,In_1670);
and U1080 (N_1080,N_759,N_505);
nor U1081 (N_1081,In_283,N_796);
xnor U1082 (N_1082,N_709,In_515);
and U1083 (N_1083,N_977,In_608);
or U1084 (N_1084,In_1458,N_171);
or U1085 (N_1085,N_452,In_1803);
xor U1086 (N_1086,N_8,In_277);
and U1087 (N_1087,N_623,In_842);
xor U1088 (N_1088,In_19,N_823);
xor U1089 (N_1089,In_876,In_2228);
nor U1090 (N_1090,N_874,N_389);
nand U1091 (N_1091,N_811,N_222);
nor U1092 (N_1092,In_1741,N_688);
nor U1093 (N_1093,N_577,In_200);
nand U1094 (N_1094,N_591,In_878);
nor U1095 (N_1095,N_526,In_374);
or U1096 (N_1096,N_535,In_1788);
xor U1097 (N_1097,In_2498,In_27);
nand U1098 (N_1098,N_519,In_1984);
xnor U1099 (N_1099,N_248,N_549);
and U1100 (N_1100,In_383,In_233);
nand U1101 (N_1101,N_578,N_769);
or U1102 (N_1102,N_618,N_660);
or U1103 (N_1103,In_1938,In_1077);
or U1104 (N_1104,N_35,In_1915);
xor U1105 (N_1105,In_192,In_2182);
nor U1106 (N_1106,N_513,N_904);
nor U1107 (N_1107,In_918,N_747);
or U1108 (N_1108,In_1724,In_229);
nand U1109 (N_1109,N_568,N_829);
nand U1110 (N_1110,In_1360,In_1820);
nand U1111 (N_1111,N_538,In_1730);
nand U1112 (N_1112,In_1530,N_923);
xor U1113 (N_1113,N_496,N_779);
or U1114 (N_1114,In_1068,In_1125);
and U1115 (N_1115,In_161,In_2023);
nor U1116 (N_1116,In_1120,In_1707);
xnor U1117 (N_1117,N_541,N_905);
and U1118 (N_1118,N_119,In_1622);
xor U1119 (N_1119,In_1306,In_1679);
nand U1120 (N_1120,In_1897,N_677);
nand U1121 (N_1121,N_822,In_520);
and U1122 (N_1122,N_51,In_641);
xnor U1123 (N_1123,In_148,In_410);
nand U1124 (N_1124,N_794,In_1018);
nand U1125 (N_1125,In_317,N_893);
or U1126 (N_1126,N_863,In_642);
xnor U1127 (N_1127,N_177,In_1570);
nor U1128 (N_1128,In_2189,In_464);
and U1129 (N_1129,N_949,In_777);
nor U1130 (N_1130,In_1541,N_781);
nand U1131 (N_1131,In_2106,N_628);
xnor U1132 (N_1132,N_844,N_692);
xnor U1133 (N_1133,N_484,In_2324);
nor U1134 (N_1134,In_1496,N_546);
nor U1135 (N_1135,In_2478,N_439);
or U1136 (N_1136,In_624,N_369);
xnor U1137 (N_1137,N_509,In_2440);
or U1138 (N_1138,N_861,N_553);
xnor U1139 (N_1139,N_391,N_491);
nand U1140 (N_1140,In_1603,In_2162);
nand U1141 (N_1141,In_1497,In_2305);
nand U1142 (N_1142,In_1196,In_1493);
or U1143 (N_1143,In_1070,In_1057);
and U1144 (N_1144,In_1838,N_879);
xor U1145 (N_1145,In_2038,N_415);
nand U1146 (N_1146,In_121,In_68);
or U1147 (N_1147,N_50,N_695);
nor U1148 (N_1148,In_2035,N_760);
nor U1149 (N_1149,In_1740,N_371);
or U1150 (N_1150,In_469,In_647);
nand U1151 (N_1151,N_962,N_14);
or U1152 (N_1152,N_574,In_1639);
or U1153 (N_1153,In_1186,In_1370);
xor U1154 (N_1154,In_2378,In_875);
nand U1155 (N_1155,In_43,In_650);
and U1156 (N_1156,N_587,In_1183);
nor U1157 (N_1157,N_678,In_186);
and U1158 (N_1158,In_703,In_504);
nor U1159 (N_1159,In_939,In_2358);
nand U1160 (N_1160,N_472,N_257);
or U1161 (N_1161,N_469,In_1859);
nand U1162 (N_1162,In_1515,N_279);
nand U1163 (N_1163,In_26,In_586);
and U1164 (N_1164,In_1606,N_792);
or U1165 (N_1165,N_979,In_1386);
xor U1166 (N_1166,N_487,N_776);
or U1167 (N_1167,N_271,In_1758);
and U1168 (N_1168,N_753,N_746);
nor U1169 (N_1169,N_934,In_904);
or U1170 (N_1170,In_1625,In_882);
nand U1171 (N_1171,In_2253,N_820);
xnor U1172 (N_1172,N_655,In_380);
nor U1173 (N_1173,N_711,In_1811);
nor U1174 (N_1174,In_738,N_630);
xor U1175 (N_1175,N_671,In_2011);
or U1176 (N_1176,In_107,N_777);
or U1177 (N_1177,In_1024,N_860);
nand U1178 (N_1178,N_720,In_1353);
nor U1179 (N_1179,N_850,N_315);
xor U1180 (N_1180,In_2442,In_1017);
nor U1181 (N_1181,N_733,In_573);
xor U1182 (N_1182,N_911,In_1262);
xnor U1183 (N_1183,N_669,N_490);
xnor U1184 (N_1184,In_2086,N_870);
xor U1185 (N_1185,In_1265,N_547);
xnor U1186 (N_1186,In_699,In_1516);
and U1187 (N_1187,N_819,In_245);
nand U1188 (N_1188,In_770,N_835);
xor U1189 (N_1189,N_598,N_648);
nor U1190 (N_1190,N_531,In_825);
or U1191 (N_1191,In_318,In_1501);
and U1192 (N_1192,N_987,In_1341);
xnor U1193 (N_1193,N_250,In_517);
xnor U1194 (N_1194,In_577,N_999);
and U1195 (N_1195,N_684,N_707);
nand U1196 (N_1196,In_1941,In_1404);
xor U1197 (N_1197,In_2200,In_1101);
xnor U1198 (N_1198,N_929,N_969);
or U1199 (N_1199,In_1040,N_918);
nor U1200 (N_1200,In_1991,In_1513);
or U1201 (N_1201,In_1860,N_282);
and U1202 (N_1202,N_932,N_990);
or U1203 (N_1203,In_354,In_1866);
xnor U1204 (N_1204,N_755,In_2487);
nor U1205 (N_1205,In_2298,N_203);
or U1206 (N_1206,In_162,In_1902);
nor U1207 (N_1207,N_230,In_497);
nand U1208 (N_1208,In_387,N_118);
nor U1209 (N_1209,N_159,In_340);
or U1210 (N_1210,N_121,N_907);
and U1211 (N_1211,N_374,N_867);
nand U1212 (N_1212,N_117,In_336);
xor U1213 (N_1213,In_2341,In_698);
nand U1214 (N_1214,N_295,In_2033);
and U1215 (N_1215,N_215,N_770);
or U1216 (N_1216,In_1418,N_570);
xor U1217 (N_1217,N_110,N_433);
or U1218 (N_1218,In_1745,N_89);
nor U1219 (N_1219,N_48,In_347);
nor U1220 (N_1220,N_700,In_2181);
or U1221 (N_1221,N_953,In_2420);
and U1222 (N_1222,In_2405,In_322);
xnor U1223 (N_1223,In_996,N_920);
or U1224 (N_1224,N_209,In_204);
or U1225 (N_1225,N_107,N_416);
nand U1226 (N_1226,In_1078,In_1806);
xnor U1227 (N_1227,In_76,N_392);
or U1228 (N_1228,In_1664,In_1977);
or U1229 (N_1229,In_179,N_612);
or U1230 (N_1230,In_1060,N_948);
xnor U1231 (N_1231,In_1762,N_988);
or U1232 (N_1232,N_659,In_17);
and U1233 (N_1233,In_147,In_1694);
and U1234 (N_1234,In_932,N_833);
and U1235 (N_1235,N_973,In_45);
and U1236 (N_1236,In_1485,N_635);
nand U1237 (N_1237,In_1174,In_375);
and U1238 (N_1238,In_2407,N_665);
nand U1239 (N_1239,In_1789,In_1205);
and U1240 (N_1240,In_610,In_2134);
or U1241 (N_1241,In_1751,In_2276);
and U1242 (N_1242,In_70,N_128);
or U1243 (N_1243,N_997,In_257);
and U1244 (N_1244,In_816,In_2151);
xnor U1245 (N_1245,N_825,In_2220);
or U1246 (N_1246,N_909,N_41);
nor U1247 (N_1247,In_1828,N_408);
nand U1248 (N_1248,In_36,In_2225);
or U1249 (N_1249,In_2280,In_79);
nor U1250 (N_1250,N_1056,N_294);
and U1251 (N_1251,In_623,In_1951);
xnor U1252 (N_1252,N_1148,N_1093);
and U1253 (N_1253,N_883,N_444);
nand U1254 (N_1254,N_142,In_1797);
xor U1255 (N_1255,In_301,N_875);
nand U1256 (N_1256,In_2335,N_782);
and U1257 (N_1257,In_2195,N_895);
and U1258 (N_1258,In_562,N_1075);
and U1259 (N_1259,N_92,N_135);
nor U1260 (N_1260,N_290,In_2327);
nor U1261 (N_1261,N_15,In_2278);
or U1262 (N_1262,In_1834,In_1020);
nand U1263 (N_1263,In_1876,N_1005);
or U1264 (N_1264,N_941,In_2031);
xnor U1265 (N_1265,In_1241,In_1899);
or U1266 (N_1266,N_1009,In_1940);
nand U1267 (N_1267,N_1141,In_1339);
or U1268 (N_1268,In_2270,N_1099);
xor U1269 (N_1269,N_1203,N_253);
or U1270 (N_1270,N_1080,N_637);
or U1271 (N_1271,In_1187,N_1140);
nand U1272 (N_1272,N_797,N_652);
nor U1273 (N_1273,In_117,In_2232);
or U1274 (N_1274,N_515,In_754);
or U1275 (N_1275,In_2371,N_865);
and U1276 (N_1276,In_1598,In_1783);
nor U1277 (N_1277,N_303,N_1090);
xor U1278 (N_1278,In_2064,N_993);
xnor U1279 (N_1279,In_1830,In_2336);
nor U1280 (N_1280,N_917,In_1965);
and U1281 (N_1281,N_1064,N_848);
xnor U1282 (N_1282,In_774,In_1486);
xor U1283 (N_1283,In_1528,In_1488);
or U1284 (N_1284,In_1382,In_919);
nand U1285 (N_1285,In_908,N_783);
xor U1286 (N_1286,N_641,N_1112);
xnor U1287 (N_1287,In_2047,N_858);
nor U1288 (N_1288,In_396,N_593);
or U1289 (N_1289,N_767,In_1218);
or U1290 (N_1290,N_627,N_317);
and U1291 (N_1291,In_25,N_1169);
xor U1292 (N_1292,In_1189,N_1149);
and U1293 (N_1293,N_246,In_1031);
or U1294 (N_1294,N_502,N_916);
nor U1295 (N_1295,N_839,N_3);
or U1296 (N_1296,In_970,In_2499);
or U1297 (N_1297,N_193,N_268);
or U1298 (N_1298,In_1421,In_2255);
nand U1299 (N_1299,In_546,N_945);
xor U1300 (N_1300,N_784,In_691);
nor U1301 (N_1301,N_757,In_1910);
or U1302 (N_1302,In_1015,N_1229);
and U1303 (N_1303,In_1182,N_702);
nand U1304 (N_1304,N_425,N_919);
xnor U1305 (N_1305,N_834,In_505);
nor U1306 (N_1306,N_859,N_849);
or U1307 (N_1307,N_731,N_1097);
xnor U1308 (N_1308,N_342,N_1173);
nand U1309 (N_1309,N_534,N_682);
nand U1310 (N_1310,N_1054,N_913);
or U1311 (N_1311,In_2068,N_1248);
and U1312 (N_1312,In_2413,In_1102);
xor U1313 (N_1313,In_1663,N_428);
nor U1314 (N_1314,In_553,In_1034);
and U1315 (N_1315,N_810,In_1194);
and U1316 (N_1316,N_190,In_587);
and U1317 (N_1317,N_1088,In_509);
and U1318 (N_1318,In_1957,N_458);
xor U1319 (N_1319,In_1452,N_1238);
xor U1320 (N_1320,N_708,In_381);
and U1321 (N_1321,In_946,N_401);
xnor U1322 (N_1322,In_687,In_273);
nor U1323 (N_1323,N_946,N_937);
xnor U1324 (N_1324,N_368,In_2475);
xnor U1325 (N_1325,N_185,N_1142);
nor U1326 (N_1326,In_1954,N_438);
and U1327 (N_1327,N_805,N_654);
xnor U1328 (N_1328,In_22,In_406);
and U1329 (N_1329,In_1244,N_639);
and U1330 (N_1330,In_1896,In_1367);
nand U1331 (N_1331,N_754,N_930);
xnor U1332 (N_1332,In_1777,N_621);
xnor U1333 (N_1333,N_881,N_1126);
xor U1334 (N_1334,N_129,N_975);
xnor U1335 (N_1335,N_1003,In_1331);
nand U1336 (N_1336,In_732,N_1035);
and U1337 (N_1337,N_804,N_892);
nand U1338 (N_1338,N_1228,In_987);
xnor U1339 (N_1339,N_772,N_1011);
nand U1340 (N_1340,In_1549,In_2387);
nand U1341 (N_1341,N_219,N_1013);
xor U1342 (N_1342,N_1123,In_2119);
and U1343 (N_1343,N_152,N_1086);
or U1344 (N_1344,N_443,N_1165);
and U1345 (N_1345,N_706,N_432);
or U1346 (N_1346,In_709,In_1389);
or U1347 (N_1347,In_768,In_1656);
or U1348 (N_1348,N_855,N_986);
and U1349 (N_1349,In_686,In_940);
nor U1350 (N_1350,N_421,In_397);
or U1351 (N_1351,N_358,N_221);
and U1352 (N_1352,N_951,N_522);
and U1353 (N_1353,In_1526,N_529);
and U1354 (N_1354,In_494,In_2246);
and U1355 (N_1355,In_772,In_96);
nor U1356 (N_1356,N_582,N_1199);
nand U1357 (N_1357,N_1130,N_651);
nor U1358 (N_1358,In_720,In_599);
or U1359 (N_1359,In_2149,N_1104);
nand U1360 (N_1360,In_1489,In_368);
and U1361 (N_1361,N_1083,N_197);
and U1362 (N_1362,N_846,In_1313);
nor U1363 (N_1363,In_1918,N_44);
nor U1364 (N_1364,In_1264,In_1050);
xnor U1365 (N_1365,In_884,N_862);
or U1366 (N_1366,N_195,In_1919);
or U1367 (N_1367,N_287,In_1213);
nand U1368 (N_1368,In_230,In_2160);
xnor U1369 (N_1369,N_396,N_524);
or U1370 (N_1370,In_652,In_1438);
or U1371 (N_1371,In_2439,N_1132);
and U1372 (N_1372,In_1648,N_756);
nand U1373 (N_1373,N_638,In_2041);
xnor U1374 (N_1374,N_633,In_1211);
nor U1375 (N_1375,In_1931,N_32);
nor U1376 (N_1376,In_288,N_1118);
nand U1377 (N_1377,N_938,In_1990);
and U1378 (N_1378,In_1998,In_1251);
xnor U1379 (N_1379,In_2249,N_251);
nor U1380 (N_1380,N_539,N_1098);
nor U1381 (N_1381,N_685,N_900);
nor U1382 (N_1382,In_2058,N_241);
or U1383 (N_1383,In_1691,N_1139);
xnor U1384 (N_1384,In_1936,N_785);
or U1385 (N_1385,N_1102,In_2334);
xor U1386 (N_1386,N_387,N_1200);
and U1387 (N_1387,N_1120,In_828);
or U1388 (N_1388,N_1197,N_99);
nand U1389 (N_1389,N_1135,N_278);
nand U1390 (N_1390,In_917,N_1241);
and U1391 (N_1391,N_1137,In_468);
and U1392 (N_1392,N_815,N_501);
and U1393 (N_1393,In_39,N_802);
xnor U1394 (N_1394,In_1441,N_1223);
nand U1395 (N_1395,In_1734,In_2063);
nand U1396 (N_1396,In_617,In_1718);
nand U1397 (N_1397,N_418,N_992);
nand U1398 (N_1398,In_1935,N_1084);
and U1399 (N_1399,In_2438,N_329);
nor U1400 (N_1400,N_931,N_764);
and U1401 (N_1401,N_1110,N_995);
nor U1402 (N_1402,N_1172,N_507);
nand U1403 (N_1403,N_749,In_2464);
and U1404 (N_1404,In_496,In_1292);
or U1405 (N_1405,In_144,N_370);
xor U1406 (N_1406,In_1579,In_564);
or U1407 (N_1407,In_901,N_259);
and U1408 (N_1408,In_1962,N_615);
nor U1409 (N_1409,N_1161,In_1659);
nor U1410 (N_1410,In_1408,N_411);
and U1411 (N_1411,In_88,N_82);
nor U1412 (N_1412,N_204,N_952);
nand U1413 (N_1413,N_233,In_60);
nor U1414 (N_1414,N_1021,In_122);
and U1415 (N_1415,In_1708,N_1089);
and U1416 (N_1416,N_927,In_2156);
nor U1417 (N_1417,In_2112,N_149);
and U1418 (N_1418,In_1447,In_1950);
xnor U1419 (N_1419,N_1121,N_419);
xnor U1420 (N_1420,In_377,In_702);
xor U1421 (N_1421,N_440,In_1611);
nand U1422 (N_1422,In_1314,N_435);
nor U1423 (N_1423,In_98,N_1201);
nor U1424 (N_1424,In_2465,N_576);
nand U1425 (N_1425,N_1008,In_15);
nor U1426 (N_1426,N_723,In_2401);
nor U1427 (N_1427,N_882,In_2019);
nand U1428 (N_1428,N_956,N_360);
or U1429 (N_1429,In_1638,N_866);
nand U1430 (N_1430,N_690,N_347);
and U1431 (N_1431,In_2388,N_1188);
nor U1432 (N_1432,N_1057,N_1063);
nor U1433 (N_1433,In_968,N_832);
or U1434 (N_1434,In_799,N_398);
or U1435 (N_1435,In_2117,N_889);
xnor U1436 (N_1436,In_453,N_1249);
nand U1437 (N_1437,N_589,N_1222);
or U1438 (N_1438,In_1437,N_234);
and U1439 (N_1439,In_1868,N_1065);
and U1440 (N_1440,In_1780,N_1074);
and U1441 (N_1441,In_784,N_1111);
or U1442 (N_1442,N_281,N_517);
nor U1443 (N_1443,N_1154,In_69);
nor U1444 (N_1444,In_1092,In_58);
xnor U1445 (N_1445,N_1208,In_1571);
or U1446 (N_1446,In_649,N_701);
xnor U1447 (N_1447,N_626,N_998);
and U1448 (N_1448,N_182,N_817);
xnor U1449 (N_1449,N_852,In_953);
nor U1450 (N_1450,In_1796,N_1000);
and U1451 (N_1451,N_1192,In_2115);
nand U1452 (N_1452,In_2217,In_1366);
nor U1453 (N_1453,N_47,In_2072);
xnor U1454 (N_1454,N_1167,In_1348);
or U1455 (N_1455,N_442,In_2453);
nor U1456 (N_1456,N_647,N_1240);
or U1457 (N_1457,N_824,N_122);
nor U1458 (N_1458,N_926,In_1164);
nor U1459 (N_1459,In_350,N_830);
and U1460 (N_1460,N_255,N_1217);
and U1461 (N_1461,N_774,In_2127);
nand U1462 (N_1462,In_849,N_806);
and U1463 (N_1463,N_966,In_196);
xor U1464 (N_1464,In_1620,N_887);
xnor U1465 (N_1465,N_864,N_338);
and U1466 (N_1466,In_915,N_167);
xor U1467 (N_1467,In_1091,N_1150);
nor U1468 (N_1468,N_1134,In_33);
nand U1469 (N_1469,N_1124,N_180);
nand U1470 (N_1470,N_672,N_1078);
and U1471 (N_1471,In_877,In_1821);
nand U1472 (N_1472,N_1204,In_1009);
or U1473 (N_1473,In_1283,N_1209);
and U1474 (N_1474,N_728,N_989);
nand U1475 (N_1475,N_958,N_267);
xor U1476 (N_1476,N_314,In_1615);
nand U1477 (N_1477,In_2137,N_1113);
or U1478 (N_1478,N_994,In_2060);
xor U1479 (N_1479,In_1581,In_596);
or U1480 (N_1480,In_2425,N_586);
nand U1481 (N_1481,N_795,In_1812);
nor U1482 (N_1482,N_213,N_629);
nor U1483 (N_1483,N_697,N_1230);
or U1484 (N_1484,N_330,N_1087);
or U1485 (N_1485,In_1927,N_174);
xnor U1486 (N_1486,In_1023,N_1038);
or U1487 (N_1487,N_978,In_1843);
and U1488 (N_1488,N_736,N_943);
xor U1489 (N_1489,N_1040,N_1092);
xor U1490 (N_1490,In_2402,In_2172);
or U1491 (N_1491,In_558,In_1505);
and U1492 (N_1492,N_694,In_885);
nor U1493 (N_1493,N_616,N_840);
nand U1494 (N_1494,N_1060,In_1760);
and U1495 (N_1495,N_65,N_1233);
and U1496 (N_1496,N_1061,In_2);
and U1497 (N_1497,In_2165,In_1445);
xor U1498 (N_1498,N_868,N_551);
or U1499 (N_1499,N_737,N_1195);
xnor U1500 (N_1500,N_1128,In_722);
nand U1501 (N_1501,In_460,In_2155);
xnor U1502 (N_1502,N_1376,In_1059);
and U1503 (N_1503,N_1409,In_1126);
nand U1504 (N_1504,In_437,N_1360);
or U1505 (N_1505,N_1423,In_1794);
nand U1506 (N_1506,In_181,N_1435);
and U1507 (N_1507,N_718,N_1107);
nor U1508 (N_1508,N_348,In_580);
nor U1509 (N_1509,In_1064,N_211);
nand U1510 (N_1510,N_1470,N_340);
nand U1511 (N_1511,N_1351,N_816);
nand U1512 (N_1512,In_126,N_1418);
xnor U1513 (N_1513,In_1987,N_1152);
nand U1514 (N_1514,N_1115,In_1098);
or U1515 (N_1515,N_1187,N_1477);
or U1516 (N_1516,N_304,N_1028);
xor U1517 (N_1517,N_1125,N_1295);
nand U1518 (N_1518,In_10,In_632);
xor U1519 (N_1519,N_1432,N_1498);
nor U1520 (N_1520,In_371,N_1037);
nor U1521 (N_1521,N_266,N_793);
nand U1522 (N_1522,In_543,N_1441);
xnor U1523 (N_1523,In_1403,In_572);
and U1524 (N_1524,N_518,N_1403);
and U1525 (N_1525,N_1309,N_896);
xor U1526 (N_1526,In_435,N_1181);
or U1527 (N_1527,In_2369,N_1373);
and U1528 (N_1528,N_721,N_354);
nand U1529 (N_1529,N_1308,In_465);
or U1530 (N_1530,In_1430,In_2265);
xnor U1531 (N_1531,N_1307,In_1956);
or U1532 (N_1532,In_212,In_454);
and U1533 (N_1533,N_1235,N_572);
nand U1534 (N_1534,N_1263,In_214);
and U1535 (N_1535,N_1273,N_1096);
or U1536 (N_1536,N_1243,N_1176);
nand U1537 (N_1537,N_751,N_1182);
nand U1538 (N_1538,In_1226,In_1243);
and U1539 (N_1539,N_1286,N_1396);
xnor U1540 (N_1540,In_1219,N_1268);
nand U1541 (N_1541,In_1926,In_1199);
or U1542 (N_1542,N_1393,In_1535);
and U1543 (N_1543,In_535,N_1114);
or U1544 (N_1544,N_366,N_1417);
or U1545 (N_1545,N_141,In_1372);
nand U1546 (N_1546,N_1299,In_756);
nand U1547 (N_1547,N_826,N_1472);
and U1548 (N_1548,N_915,N_1483);
nand U1549 (N_1549,In_2379,N_1290);
nand U1550 (N_1550,N_1339,N_1420);
nand U1551 (N_1551,N_516,In_943);
nor U1552 (N_1552,In_174,N_1219);
or U1553 (N_1553,N_914,N_1414);
nor U1554 (N_1554,N_1454,N_1305);
nand U1555 (N_1555,In_360,N_1412);
and U1556 (N_1556,N_1020,N_897);
nor U1557 (N_1557,N_1386,N_60);
and U1558 (N_1558,In_1449,N_1267);
nor U1559 (N_1559,N_1278,N_1265);
or U1560 (N_1560,N_942,In_839);
and U1561 (N_1561,In_1994,In_1272);
nor U1562 (N_1562,N_668,N_1287);
nand U1563 (N_1563,In_1547,N_1328);
or U1564 (N_1564,N_1363,N_1450);
nand U1565 (N_1565,In_1750,N_954);
xor U1566 (N_1566,N_1446,In_858);
or U1567 (N_1567,N_1499,N_1387);
or U1568 (N_1568,N_25,N_936);
nand U1569 (N_1569,N_1375,In_2055);
nand U1570 (N_1570,N_471,N_1391);
nor U1571 (N_1571,N_880,In_2268);
nor U1572 (N_1572,In_2168,In_707);
nor U1573 (N_1573,N_372,In_1907);
nand U1574 (N_1574,In_1884,N_1313);
nor U1575 (N_1575,In_2312,N_393);
and U1576 (N_1576,N_53,In_2108);
xor U1577 (N_1577,N_511,In_615);
xnor U1578 (N_1578,N_130,N_90);
or U1579 (N_1579,N_1103,In_2389);
nor U1580 (N_1580,In_139,N_322);
or U1581 (N_1581,In_1075,In_659);
nor U1582 (N_1582,N_1091,N_1459);
or U1583 (N_1583,N_1072,In_1825);
xor U1584 (N_1584,N_1304,N_944);
or U1585 (N_1585,N_1392,In_426);
nor U1586 (N_1586,N_1010,N_1030);
nor U1587 (N_1587,In_706,In_314);
or U1588 (N_1588,N_821,N_1429);
and U1589 (N_1589,N_1437,N_1453);
nor U1590 (N_1590,In_455,N_1369);
nor U1591 (N_1591,In_339,N_163);
or U1592 (N_1592,N_528,N_1133);
xnor U1593 (N_1593,N_841,N_1211);
or U1594 (N_1594,N_872,In_1397);
and U1595 (N_1595,N_1191,N_1046);
xor U1596 (N_1596,N_976,In_503);
or U1597 (N_1597,In_1448,N_899);
or U1598 (N_1598,N_645,In_1871);
nand U1599 (N_1599,N_445,N_1024);
xnor U1600 (N_1600,N_1257,In_2157);
and U1601 (N_1601,N_1471,In_1434);
xnor U1602 (N_1602,N_1105,N_1215);
nor U1603 (N_1603,N_293,In_1095);
nor U1604 (N_1604,N_1071,N_1279);
xnor U1605 (N_1605,In_429,N_1486);
xor U1606 (N_1606,N_1316,In_1311);
nor U1607 (N_1607,N_1400,N_9);
and U1608 (N_1608,In_1607,N_714);
nor U1609 (N_1609,In_2390,N_305);
and U1610 (N_1610,In_2309,N_1456);
nor U1611 (N_1611,N_877,In_874);
and U1612 (N_1612,N_327,N_1016);
xnor U1613 (N_1613,N_1070,In_1373);
nor U1614 (N_1614,N_959,In_1312);
nor U1615 (N_1615,In_364,In_2450);
or U1616 (N_1616,N_1157,N_675);
nand U1617 (N_1617,In_1288,N_752);
and U1618 (N_1618,N_537,N_1406);
xnor U1619 (N_1619,N_1006,In_500);
xnor U1620 (N_1620,In_1799,In_358);
and U1621 (N_1621,In_1358,N_984);
xor U1622 (N_1622,N_910,N_1293);
nor U1623 (N_1623,In_1473,N_1261);
nor U1624 (N_1624,N_1210,N_61);
nor U1625 (N_1625,N_186,N_27);
xor U1626 (N_1626,N_813,N_260);
or U1627 (N_1627,N_346,N_1216);
or U1628 (N_1628,N_1109,In_613);
xor U1629 (N_1629,N_1436,N_742);
nand U1630 (N_1630,N_104,N_1059);
or U1631 (N_1631,In_597,N_925);
nand U1632 (N_1632,N_1347,N_1255);
nand U1633 (N_1633,N_1467,N_548);
and U1634 (N_1634,In_175,N_506);
or U1635 (N_1635,In_1142,N_778);
nand U1636 (N_1636,N_456,In_325);
and U1637 (N_1637,N_1461,N_814);
nand U1638 (N_1638,In_471,N_262);
nor U1639 (N_1639,N_933,N_470);
nor U1640 (N_1640,In_1407,In_2488);
nand U1641 (N_1641,In_1817,N_1275);
and U1642 (N_1642,In_1514,N_1270);
or U1643 (N_1643,In_942,N_373);
xnor U1644 (N_1644,N_800,In_138);
or U1645 (N_1645,N_1345,N_799);
xnor U1646 (N_1646,In_211,N_264);
xor U1647 (N_1647,N_1050,N_1294);
and U1648 (N_1648,N_1002,N_1052);
nor U1649 (N_1649,In_2426,In_2132);
and U1650 (N_1650,N_1033,N_1053);
and U1651 (N_1651,In_1764,In_1198);
or U1652 (N_1652,In_1065,N_924);
nor U1653 (N_1653,In_1721,N_1399);
nor U1654 (N_1654,N_1462,N_1202);
and U1655 (N_1655,N_1321,N_1143);
and U1656 (N_1656,N_318,N_1326);
and U1657 (N_1657,In_473,N_786);
nor U1658 (N_1658,N_1079,N_270);
xnor U1659 (N_1659,In_895,N_33);
nand U1660 (N_1660,N_1205,In_729);
and U1661 (N_1661,N_940,In_372);
xnor U1662 (N_1662,N_613,N_249);
xor U1663 (N_1663,N_236,N_617);
nand U1664 (N_1664,N_1129,In_1580);
nor U1665 (N_1665,N_1319,N_462);
nand U1666 (N_1666,N_567,N_1213);
or U1667 (N_1667,N_1388,N_1022);
xor U1668 (N_1668,In_1671,In_981);
nand U1669 (N_1669,In_499,N_854);
xnor U1670 (N_1670,In_1807,In_913);
or U1671 (N_1671,In_2044,N_1254);
nor U1672 (N_1672,In_1731,In_2190);
and U1673 (N_1673,N_555,N_1315);
nand U1674 (N_1674,In_926,In_1149);
and U1675 (N_1675,In_2351,N_1193);
nor U1676 (N_1676,N_545,N_536);
nand U1677 (N_1677,N_636,In_636);
and U1678 (N_1678,In_1396,N_175);
nor U1679 (N_1679,N_761,N_475);
or U1680 (N_1680,In_172,N_1274);
or U1681 (N_1681,N_947,N_745);
nor U1682 (N_1682,In_2416,N_1122);
xor U1683 (N_1683,N_493,N_928);
nand U1684 (N_1684,N_1117,N_291);
or U1685 (N_1685,In_724,N_1482);
and U1686 (N_1686,N_789,N_227);
nand U1687 (N_1687,N_1468,In_1295);
nand U1688 (N_1688,In_1747,N_1252);
xor U1689 (N_1689,In_537,N_1138);
xor U1690 (N_1690,N_1001,N_337);
xnor U1691 (N_1691,N_791,In_2128);
nand U1692 (N_1692,N_1029,N_1421);
or U1693 (N_1693,N_1260,In_420);
nand U1694 (N_1694,N_878,N_1178);
and U1695 (N_1695,In_2367,In_2466);
xor U1696 (N_1696,N_716,N_1292);
or U1697 (N_1697,N_902,N_1171);
and U1698 (N_1698,N_1023,N_1452);
and U1699 (N_1699,N_1177,N_1395);
nand U1700 (N_1700,N_1492,N_922);
nor U1701 (N_1701,In_1328,In_1131);
nand U1702 (N_1702,N_1344,In_2089);
nand U1703 (N_1703,In_704,N_894);
nand U1704 (N_1704,N_1490,N_1302);
or U1705 (N_1705,N_1455,N_1425);
nor U1706 (N_1706,In_1979,In_1651);
nor U1707 (N_1707,In_1588,In_1814);
nor U1708 (N_1708,N_674,In_900);
xnor U1709 (N_1709,In_804,In_132);
nand U1710 (N_1710,N_1196,N_1410);
nor U1711 (N_1711,N_1296,In_1967);
xnor U1712 (N_1712,In_1989,N_1276);
nor U1713 (N_1713,N_653,N_1465);
or U1714 (N_1714,N_1258,N_1469);
nand U1715 (N_1715,N_961,N_542);
nor U1716 (N_1716,In_1626,In_1920);
xnor U1717 (N_1717,In_1468,N_1405);
xnor U1718 (N_1718,In_75,In_594);
nand U1719 (N_1719,N_1479,N_1367);
and U1720 (N_1720,N_1069,In_1748);
and U1721 (N_1721,N_1220,N_991);
nor U1722 (N_1722,N_63,N_985);
nor U1723 (N_1723,In_889,N_564);
or U1724 (N_1724,N_1127,N_1389);
or U1725 (N_1725,N_644,N_1198);
nor U1726 (N_1726,N_1004,In_1476);
and U1727 (N_1727,In_244,N_1424);
and U1728 (N_1728,N_735,In_526);
or U1729 (N_1729,N_1463,In_269);
nand U1730 (N_1730,In_47,N_888);
and U1731 (N_1731,N_1153,N_1350);
nor U1732 (N_1732,In_448,In_1380);
nand U1733 (N_1733,N_600,N_1170);
nor U1734 (N_1734,In_1170,N_1433);
and U1735 (N_1735,N_575,In_416);
nor U1736 (N_1736,N_1374,In_37);
nor U1737 (N_1737,N_1457,In_2258);
nand U1738 (N_1738,In_1878,N_464);
nand U1739 (N_1739,In_976,In_1848);
xnor U1740 (N_1740,N_1027,N_1018);
and U1741 (N_1741,N_1364,N_1151);
xor U1742 (N_1742,N_592,In_2293);
nor U1743 (N_1743,N_1048,N_93);
xor U1744 (N_1744,In_1410,N_765);
and U1745 (N_1745,N_650,N_218);
and U1746 (N_1746,N_1206,In_822);
nand U1747 (N_1747,In_2221,N_1180);
and U1748 (N_1748,N_1439,N_787);
nor U1749 (N_1749,In_1347,N_595);
nand U1750 (N_1750,N_1660,N_921);
or U1751 (N_1751,N_803,N_1729);
nand U1752 (N_1752,N_410,N_1572);
xor U1753 (N_1753,N_691,In_1593);
xor U1754 (N_1754,In_51,N_1545);
and U1755 (N_1755,N_1159,N_1478);
nand U1756 (N_1756,N_681,In_327);
or U1757 (N_1757,N_1697,In_2102);
nand U1758 (N_1758,N_1514,N_1160);
or U1759 (N_1759,N_1311,N_1523);
and U1760 (N_1760,In_177,N_1381);
and U1761 (N_1761,In_156,N_1303);
and U1762 (N_1762,In_2142,In_1340);
or U1763 (N_1763,N_1253,N_1357);
nor U1764 (N_1764,N_1535,In_2016);
nor U1765 (N_1765,N_1272,N_1608);
or U1766 (N_1766,N_1702,N_1047);
nand U1767 (N_1767,N_1166,N_768);
nand U1768 (N_1768,In_100,N_1485);
xnor U1769 (N_1769,N_1156,In_1738);
nor U1770 (N_1770,In_1605,N_1548);
xnor U1771 (N_1771,N_1227,In_446);
nor U1772 (N_1772,In_2331,N_836);
xor U1773 (N_1773,N_1378,N_1081);
and U1774 (N_1774,N_1571,In_209);
nand U1775 (N_1775,N_1636,N_1665);
xor U1776 (N_1776,N_1610,In_2144);
or U1777 (N_1777,N_1017,N_1542);
nand U1778 (N_1778,N_818,N_237);
and U1779 (N_1779,N_1672,In_308);
nand U1780 (N_1780,N_579,N_1224);
xnor U1781 (N_1781,N_1269,N_540);
nand U1782 (N_1782,In_1678,N_1489);
and U1783 (N_1783,N_1353,N_133);
nor U1784 (N_1784,N_1609,N_967);
or U1785 (N_1785,N_1318,N_1473);
or U1786 (N_1786,N_1558,N_583);
nor U1787 (N_1787,N_1012,N_1415);
or U1788 (N_1788,In_2279,In_993);
nor U1789 (N_1789,N_1551,N_1716);
nor U1790 (N_1790,N_1359,N_6);
and U1791 (N_1791,N_207,N_1236);
and U1792 (N_1792,N_1158,N_1266);
xnor U1793 (N_1793,In_1553,In_2026);
and U1794 (N_1794,N_970,N_1175);
xor U1795 (N_1795,N_1603,N_1051);
xor U1796 (N_1796,N_1427,In_817);
or U1797 (N_1797,N_1247,In_1521);
xor U1798 (N_1798,In_1801,In_1874);
and U1799 (N_1799,In_385,In_677);
xor U1800 (N_1800,In_1930,N_1563);
xnor U1801 (N_1801,N_1145,N_1034);
and U1802 (N_1802,N_1742,In_2002);
nor U1803 (N_1803,N_1717,N_950);
nand U1804 (N_1804,N_1179,N_1673);
or U1805 (N_1805,In_2125,N_1517);
and U1806 (N_1806,N_744,N_1271);
or U1807 (N_1807,In_2411,N_857);
xor U1808 (N_1808,In_1305,In_1107);
nand U1809 (N_1809,N_1566,N_908);
nor U1810 (N_1810,N_341,N_1668);
nor U1811 (N_1811,N_1163,N_1743);
xor U1812 (N_1812,N_1082,N_1509);
nor U1813 (N_1813,N_1361,N_394);
or U1814 (N_1814,N_57,N_1495);
and U1815 (N_1815,In_1557,N_326);
or U1816 (N_1816,N_1411,N_1448);
and U1817 (N_1817,In_1960,N_1657);
nor U1818 (N_1818,N_1595,N_1310);
and U1819 (N_1819,N_1264,N_1623);
nand U1820 (N_1820,N_812,In_2259);
xor U1821 (N_1821,N_1340,N_1282);
xnor U1822 (N_1822,N_1330,In_1841);
and U1823 (N_1823,N_1362,N_1358);
xnor U1824 (N_1824,N_1085,N_845);
and U1825 (N_1825,N_1333,In_1342);
nand U1826 (N_1826,N_1701,N_1640);
and U1827 (N_1827,N_1703,N_1648);
or U1828 (N_1828,N_1356,N_1671);
xnor U1829 (N_1829,N_1475,N_1190);
nor U1830 (N_1830,N_1505,N_1493);
or U1831 (N_1831,N_1385,In_1046);
or U1832 (N_1832,N_912,In_1766);
and U1833 (N_1833,In_1304,N_1066);
and U1834 (N_1834,N_906,N_1575);
xor U1835 (N_1835,In_95,N_1426);
or U1836 (N_1836,N_1407,N_417);
xor U1837 (N_1837,N_1068,In_1477);
and U1838 (N_1838,In_1913,N_1106);
or U1839 (N_1839,N_1183,N_1297);
and U1840 (N_1840,N_1488,N_1547);
or U1841 (N_1841,N_1042,N_1503);
xnor U1842 (N_1842,N_680,N_1639);
nand U1843 (N_1843,In_298,N_1402);
nor U1844 (N_1844,N_1334,N_1587);
nor U1845 (N_1845,N_1464,In_1862);
or U1846 (N_1846,N_1428,N_717);
xnor U1847 (N_1847,N_837,N_605);
xor U1848 (N_1848,N_1695,In_197);
and U1849 (N_1849,N_885,N_1250);
nand U1850 (N_1850,N_1522,N_1747);
nor U1851 (N_1851,N_1368,N_1629);
nand U1852 (N_1852,In_1254,N_1601);
or U1853 (N_1853,N_1622,N_981);
or U1854 (N_1854,N_1715,In_1619);
nor U1855 (N_1855,N_1589,N_1527);
and U1856 (N_1856,N_1588,N_1280);
or U1857 (N_1857,N_1283,N_766);
xor U1858 (N_1858,In_224,N_1323);
or U1859 (N_1859,In_1368,N_758);
xnor U1860 (N_1860,N_1604,N_1045);
nand U1861 (N_1861,N_1346,N_1076);
and U1862 (N_1862,N_172,N_512);
xnor U1863 (N_1863,N_729,In_1222);
or U1864 (N_1864,N_532,N_1533);
or U1865 (N_1865,N_1073,N_1515);
xnor U1866 (N_1866,In_1022,In_1591);
nor U1867 (N_1867,In_2070,N_1694);
and U1868 (N_1868,N_1683,In_1773);
or U1869 (N_1869,N_1658,N_455);
nand U1870 (N_1870,N_1447,N_1681);
or U1871 (N_1871,In_929,N_828);
or U1872 (N_1872,N_1733,N_884);
or U1873 (N_1873,N_1225,N_1371);
or U1874 (N_1874,N_1534,N_1590);
xnor U1875 (N_1875,N_1365,N_1707);
nand U1876 (N_1876,In_1076,In_1953);
xnor U1877 (N_1877,N_1725,In_30);
xnor U1878 (N_1878,N_1317,In_1228);
xnor U1879 (N_1879,N_1544,In_13);
or U1880 (N_1880,N_1430,N_1460);
nand U1881 (N_1881,N_1384,N_1131);
nand U1882 (N_1882,N_1625,N_1390);
and U1883 (N_1883,N_1422,N_1408);
and U1884 (N_1884,N_1557,N_1650);
or U1885 (N_1885,N_712,In_838);
or U1886 (N_1886,N_1049,N_661);
xor U1887 (N_1887,N_112,N_1458);
xnor U1888 (N_1888,N_1568,N_1329);
nand U1889 (N_1889,N_1559,N_386);
and U1890 (N_1890,N_1730,N_1713);
and U1891 (N_1891,N_590,N_1508);
or U1892 (N_1892,N_223,N_1724);
nand U1893 (N_1893,N_1584,N_1259);
nor U1894 (N_1894,N_521,N_1630);
nor U1895 (N_1895,N_622,N_1519);
nor U1896 (N_1896,In_749,In_1071);
or U1897 (N_1897,N_1095,In_1554);
and U1898 (N_1898,In_73,N_1289);
or U1899 (N_1899,In_1726,In_23);
xor U1900 (N_1900,N_1438,In_1686);
nor U1901 (N_1901,N_1506,N_640);
or U1902 (N_1902,N_1094,In_622);
or U1903 (N_1903,N_1643,N_1449);
and U1904 (N_1904,N_20,N_1667);
nor U1905 (N_1905,N_1306,In_1317);
or U1906 (N_1906,N_1136,N_1502);
and U1907 (N_1907,N_1100,N_1634);
or U1908 (N_1908,N_801,N_1256);
xor U1909 (N_1909,In_1502,N_1397);
nand U1910 (N_1910,N_1746,N_581);
nor U1911 (N_1911,In_2408,In_1658);
nor U1912 (N_1912,N_1670,N_1062);
or U1913 (N_1913,N_1612,N_1147);
and U1914 (N_1914,N_1019,N_1144);
or U1915 (N_1915,In_456,In_1483);
and U1916 (N_1916,N_1529,N_1585);
and U1917 (N_1917,N_1655,N_468);
xnor U1918 (N_1918,N_569,In_432);
nand U1919 (N_1919,N_1162,N_1741);
nand U1920 (N_1920,In_1829,N_1281);
nand U1921 (N_1921,N_1740,N_1491);
nor U1922 (N_1922,N_1524,N_1719);
xor U1923 (N_1923,N_1394,In_673);
xor U1924 (N_1924,N_798,In_373);
xor U1925 (N_1925,N_664,N_1526);
xnor U1926 (N_1926,N_1354,N_1659);
nand U1927 (N_1927,N_1687,N_1689);
nand U1928 (N_1928,N_1606,In_458);
nor U1929 (N_1929,N_1569,N_1581);
or U1930 (N_1930,N_1739,N_1647);
and U1931 (N_1931,N_1036,In_1435);
or U1932 (N_1932,N_1593,N_1416);
and U1933 (N_1933,N_1616,N_1582);
and U1934 (N_1934,N_739,N_1285);
or U1935 (N_1935,N_1732,N_1288);
nor U1936 (N_1936,N_1685,N_1349);
and U1937 (N_1937,N_1594,In_524);
or U1938 (N_1938,N_1641,N_1500);
nor U1939 (N_1939,N_1669,In_1692);
and U1940 (N_1940,N_1322,N_73);
nor U1941 (N_1941,N_871,N_1624);
xor U1942 (N_1942,N_1325,N_1413);
nand U1943 (N_1943,N_1301,N_1607);
nand U1944 (N_1944,N_1574,N_1684);
and U1945 (N_1945,N_1749,N_1564);
nor U1946 (N_1946,N_1664,N_1431);
nor U1947 (N_1947,In_1872,In_948);
nor U1948 (N_1948,N_571,N_1674);
nor U1949 (N_1949,In_1633,N_1735);
and U1950 (N_1950,N_1532,N_356);
xor U1951 (N_1951,N_1745,N_1619);
and U1952 (N_1952,N_1383,N_1737);
nand U1953 (N_1953,N_1244,N_1366);
and U1954 (N_1954,N_1580,N_609);
xnor U1955 (N_1955,N_1599,N_1212);
nor U1956 (N_1956,N_1442,N_1576);
and U1957 (N_1957,N_869,N_1718);
xnor U1958 (N_1958,N_1613,N_1679);
nor U1959 (N_1959,N_1675,N_1434);
or U1960 (N_1960,N_1277,In_343);
or U1961 (N_1961,N_980,N_1320);
or U1962 (N_1962,N_1627,N_1530);
and U1963 (N_1963,N_1677,In_400);
nand U1964 (N_1964,N_1015,N_1044);
and U1965 (N_1965,N_1714,N_935);
nor U1966 (N_1966,N_679,In_956);
and U1967 (N_1967,N_1600,In_1475);
or U1968 (N_1968,N_1680,N_1605);
nor U1969 (N_1969,In_2480,N_1487);
nand U1970 (N_1970,N_1645,N_1602);
nor U1971 (N_1971,N_1693,N_1646);
xor U1972 (N_1972,N_1543,N_1077);
or U1973 (N_1973,In_1739,In_1431);
and U1974 (N_1974,N_738,N_1642);
nor U1975 (N_1975,N_1690,In_1643);
or U1976 (N_1976,N_1734,N_1573);
nor U1977 (N_1977,In_390,N_1025);
and U1978 (N_1978,N_1704,In_965);
nand U1979 (N_1979,N_1398,N_771);
or U1980 (N_1980,N_873,N_1466);
xnor U1981 (N_1981,N_1401,N_1586);
nor U1982 (N_1982,N_1700,N_1300);
and U1983 (N_1983,N_1537,N_1218);
nand U1984 (N_1984,N_1168,N_1332);
or U1985 (N_1985,N_189,N_1652);
and U1986 (N_1986,N_1705,N_1214);
nand U1987 (N_1987,N_1440,N_1536);
xor U1988 (N_1988,N_1511,N_1338);
xnor U1989 (N_1989,N_1661,In_1216);
xor U1990 (N_1990,In_1323,N_550);
nor U1991 (N_1991,N_1101,N_1578);
nand U1992 (N_1992,In_2053,N_1184);
and U1993 (N_1993,N_1662,N_1342);
nor U1994 (N_1994,N_1521,N_1242);
or U1995 (N_1995,N_1239,In_788);
nand U1996 (N_1996,In_892,N_1380);
nor U1997 (N_1997,N_88,N_1370);
and U1998 (N_1998,N_631,N_1043);
xnor U1999 (N_1999,N_1480,In_751);
nand U2000 (N_2000,N_1520,N_1484);
or U2001 (N_2001,N_1829,N_1785);
xor U2002 (N_2002,N_1443,N_1644);
nand U2003 (N_2003,N_1839,N_1855);
nor U2004 (N_2004,N_1963,N_1251);
and U2005 (N_2005,N_1895,N_1805);
nor U2006 (N_2006,N_1404,N_1959);
and U2007 (N_2007,N_1540,N_1800);
xnor U2008 (N_2008,N_1744,N_1560);
xnor U2009 (N_2009,N_1858,In_1982);
and U2010 (N_2010,N_1245,N_1709);
and U2011 (N_2011,N_1961,N_1846);
nand U2012 (N_2012,N_1753,N_971);
or U2013 (N_2013,In_438,N_596);
nor U2014 (N_2014,N_1851,In_637);
nand U2015 (N_2015,N_1341,N_131);
or U2016 (N_2016,N_1174,N_1999);
nor U2017 (N_2017,N_1874,N_1894);
or U2018 (N_2018,In_1276,N_1696);
or U2019 (N_2019,N_319,N_1893);
or U2020 (N_2020,N_1859,N_1798);
or U2021 (N_2021,N_1723,N_1801);
and U2022 (N_2022,In_1337,In_1509);
and U2023 (N_2023,In_566,N_1828);
and U2024 (N_2024,N_1738,N_1981);
and U2025 (N_2025,N_1419,N_328);
and U2026 (N_2026,N_780,N_1312);
nand U2027 (N_2027,N_1754,N_1996);
or U2028 (N_2028,N_1885,N_1902);
nand U2029 (N_2029,N_1611,In_154);
or U2030 (N_2030,N_1884,N_1379);
xor U2031 (N_2031,N_1722,N_1862);
and U2032 (N_2032,N_1116,N_1780);
xnor U2033 (N_2033,N_1871,N_1567);
nand U2034 (N_2034,In_1959,N_1811);
nand U2035 (N_2035,N_827,N_1816);
nand U2036 (N_2036,N_1977,N_1790);
xnor U2037 (N_2037,N_1032,In_627);
xnor U2038 (N_2038,N_1878,N_1881);
xnor U2039 (N_2039,N_1776,N_1653);
nand U2040 (N_2040,N_1770,N_1583);
or U2041 (N_2041,N_1993,N_1194);
nand U2042 (N_2042,N_1866,N_1314);
and U2043 (N_2043,N_1982,N_1343);
xnor U2044 (N_2044,In_2066,N_1232);
nor U2045 (N_2045,N_1969,In_253);
or U2046 (N_2046,N_1970,N_1908);
and U2047 (N_2047,N_81,In_2025);
nand U2048 (N_2048,N_1539,N_1055);
xnor U2049 (N_2049,N_1731,N_1840);
nand U2050 (N_2050,N_1759,N_1663);
xor U2051 (N_2051,N_1951,N_963);
nand U2052 (N_2052,N_1799,In_1767);
nor U2053 (N_2053,N_1968,N_750);
xnor U2054 (N_2054,In_1047,N_1758);
and U2055 (N_2055,In_1587,N_1931);
or U2056 (N_2056,N_216,N_377);
nand U2057 (N_2057,In_1525,N_1854);
and U2058 (N_2058,N_1451,In_403);
xnor U2059 (N_2059,N_1974,N_1880);
nor U2060 (N_2060,N_1934,N_1284);
xor U2061 (N_2061,N_1992,N_1555);
xor U2062 (N_2062,N_1956,N_1591);
nor U2063 (N_2063,N_1789,N_1843);
nor U2064 (N_2064,N_1949,N_996);
or U2065 (N_2065,N_1980,N_1888);
nor U2066 (N_2066,N_1922,N_1875);
nand U2067 (N_2067,N_1649,N_1937);
nand U2068 (N_2068,N_474,N_1597);
xor U2069 (N_2069,N_1913,N_585);
nor U2070 (N_2070,In_49,N_1997);
or U2071 (N_2071,N_1676,N_1549);
xor U2072 (N_2072,N_1337,N_1771);
or U2073 (N_2073,N_1654,N_1822);
or U2074 (N_2074,In_440,N_1237);
and U2075 (N_2075,N_1155,N_1797);
nand U2076 (N_2076,In_491,N_693);
nor U2077 (N_2077,N_1942,N_1762);
nand U2078 (N_2078,In_1163,N_1955);
nand U2079 (N_2079,N_1510,N_1925);
and U2080 (N_2080,N_773,N_298);
xnor U2081 (N_2081,N_1765,N_1698);
and U2082 (N_2082,N_1755,N_1531);
nand U2083 (N_2083,N_1699,N_1058);
or U2084 (N_2084,N_1876,N_1474);
nor U2085 (N_2085,N_1528,N_1618);
nor U2086 (N_2086,N_1504,N_1892);
or U2087 (N_2087,N_1927,N_1826);
and U2088 (N_2088,N_1525,N_1932);
nand U2089 (N_2089,N_1807,N_1986);
xnor U2090 (N_2090,N_1164,In_1266);
and U2091 (N_2091,N_1818,N_1119);
nor U2092 (N_2092,In_2110,N_1031);
nand U2093 (N_2093,N_1995,N_1819);
xnor U2094 (N_2094,N_843,N_1513);
xor U2095 (N_2095,N_1146,N_1331);
and U2096 (N_2096,N_1838,N_1221);
nand U2097 (N_2097,N_1761,N_1912);
or U2098 (N_2098,N_1682,N_1945);
xor U2099 (N_2099,N_1561,N_1708);
nor U2100 (N_2100,N_1978,In_685);
nor U2101 (N_2101,N_1335,N_1928);
xnor U2102 (N_2102,N_1621,N_1631);
or U2103 (N_2103,N_385,N_403);
and U2104 (N_2104,N_1901,N_1896);
nand U2105 (N_2105,N_1727,In_2284);
xor U2106 (N_2106,N_1991,N_1596);
nand U2107 (N_2107,N_1935,N_1939);
xnor U2108 (N_2108,N_1845,N_1965);
and U2109 (N_2109,N_489,N_1633);
nand U2110 (N_2110,N_1910,In_992);
nand U2111 (N_2111,N_1953,N_1849);
or U2112 (N_2112,N_1900,N_1686);
and U2113 (N_2113,N_1924,N_1906);
and U2114 (N_2114,N_1481,N_1809);
or U2115 (N_2115,N_1907,N_704);
xor U2116 (N_2116,N_1706,N_1577);
xor U2117 (N_2117,N_1938,N_1947);
nand U2118 (N_2118,N_1553,N_1518);
or U2119 (N_2119,N_1444,N_1820);
and U2120 (N_2120,N_1766,N_939);
nand U2121 (N_2121,N_1920,In_853);
or U2122 (N_2122,N_1827,N_1887);
xnor U2123 (N_2123,N_1108,N_1445);
xnor U2124 (N_2124,N_1638,N_1786);
nand U2125 (N_2125,N_982,N_1973);
nor U2126 (N_2126,N_1833,N_1711);
nand U2127 (N_2127,N_1628,N_1796);
or U2128 (N_2128,N_901,N_1853);
nor U2129 (N_2129,N_1779,N_1760);
and U2130 (N_2130,N_1848,N_1909);
xor U2131 (N_2131,N_1857,N_1750);
or U2132 (N_2132,N_1911,N_1554);
and U2133 (N_2133,N_1940,N_1933);
and U2134 (N_2134,N_1964,N_1751);
xnor U2135 (N_2135,N_2,N_1975);
nand U2136 (N_2136,N_1842,N_1617);
or U2137 (N_2137,In_2296,N_808);
nand U2138 (N_2138,N_1792,N_1666);
nor U2139 (N_2139,N_1966,N_1494);
and U2140 (N_2140,N_1890,N_1579);
nand U2141 (N_2141,In_565,N_1943);
xnor U2142 (N_2142,N_1837,N_1752);
or U2143 (N_2143,N_1877,N_1728);
nor U2144 (N_2144,N_1757,N_1512);
nand U2145 (N_2145,N_1879,In_797);
nand U2146 (N_2146,N_388,N_1772);
xnor U2147 (N_2147,N_1836,N_1592);
or U2148 (N_2148,N_1615,N_1778);
xor U2149 (N_2149,N_1921,N_1841);
nand U2150 (N_2150,N_1941,N_1516);
xnor U2151 (N_2151,N_1773,N_1007);
and U2152 (N_2152,N_1355,N_1720);
nand U2153 (N_2153,N_1882,N_1787);
nor U2154 (N_2154,N_1919,In_820);
or U2155 (N_2155,N_601,N_1869);
xnor U2156 (N_2156,In_1537,N_1821);
nand U2157 (N_2157,N_1620,N_1844);
or U2158 (N_2158,N_1962,In_696);
and U2159 (N_2159,N_1507,N_1550);
and U2160 (N_2160,N_5,N_1352);
xor U2161 (N_2161,N_960,In_886);
or U2162 (N_2162,N_448,In_1054);
and U2163 (N_2163,N_1726,N_1972);
nor U2164 (N_2164,N_1998,In_2223);
nand U2165 (N_2165,N_1950,N_1791);
or U2166 (N_2166,N_1691,N_1823);
xor U2167 (N_2167,N_1915,N_1496);
xnor U2168 (N_2168,N_364,N_1777);
nand U2169 (N_2169,N_1039,N_1710);
xor U2170 (N_2170,N_1898,N_1763);
and U2171 (N_2171,N_1538,N_1944);
xnor U2172 (N_2172,In_355,N_1688);
nor U2173 (N_2173,In_450,N_1825);
xor U2174 (N_2174,N_1889,N_1546);
nor U2175 (N_2175,N_1541,N_1856);
and U2176 (N_2176,N_1979,N_1883);
and U2177 (N_2177,N_1501,N_1808);
xor U2178 (N_2178,N_1185,N_1867);
xor U2179 (N_2179,N_1656,N_1806);
and U2180 (N_2180,N_1863,N_1041);
nand U2181 (N_2181,In_2235,N_136);
or U2182 (N_2182,N_1067,N_1736);
nor U2183 (N_2183,N_1794,N_1917);
xnor U2184 (N_2184,N_1784,N_1954);
nor U2185 (N_2185,N_1983,N_1804);
xnor U2186 (N_2186,N_1767,N_1916);
nand U2187 (N_2187,N_1327,N_1476);
nand U2188 (N_2188,N_1336,N_1994);
xor U2189 (N_2189,N_1903,N_847);
and U2190 (N_2190,N_1298,N_1781);
xnor U2191 (N_2191,N_1930,N_624);
or U2192 (N_2192,In_164,N_1756);
xnor U2193 (N_2193,In_1610,In_2395);
or U2194 (N_2194,N_1960,N_1324);
nor U2195 (N_2195,In_1139,N_1865);
xnor U2196 (N_2196,N_1817,N_1872);
or U2197 (N_2197,N_1824,N_666);
nand U2198 (N_2198,N_1782,N_1774);
xor U2199 (N_2199,N_1764,N_831);
nand U2200 (N_2200,N_1860,N_1990);
or U2201 (N_2201,N_1886,N_1831);
and U2202 (N_2202,N_1793,N_1768);
or U2203 (N_2203,N_1946,N_1868);
or U2204 (N_2204,N_1186,N_350);
xor U2205 (N_2205,N_1899,N_1556);
nor U2206 (N_2206,N_1614,In_1085);
xor U2207 (N_2207,N_1812,N_1189);
nor U2208 (N_2208,N_1372,N_1598);
or U2209 (N_2209,N_1207,N_1815);
or U2210 (N_2210,In_1099,N_1923);
nand U2211 (N_2211,N_1957,N_1803);
or U2212 (N_2212,N_1897,N_1864);
or U2213 (N_2213,N_1904,N_1847);
xor U2214 (N_2214,N_1775,N_790);
nor U2215 (N_2215,N_1852,N_1246);
or U2216 (N_2216,N_1632,N_1795);
nor U2217 (N_2217,N_1948,In_1665);
or U2218 (N_2218,N_1637,In_2237);
or U2219 (N_2219,N_1226,N_1565);
nand U2220 (N_2220,N_886,N_1769);
and U2221 (N_2221,N_1873,N_434);
nor U2222 (N_2222,N_1626,N_1985);
nor U2223 (N_2223,N_1936,N_1984);
nand U2224 (N_2224,N_1989,N_1802);
xor U2225 (N_2225,N_1967,N_1497);
nor U2226 (N_2226,N_1234,N_1814);
nand U2227 (N_2227,N_1570,N_1952);
nand U2228 (N_2228,N_1721,N_1830);
nor U2229 (N_2229,N_788,N_1026);
or U2230 (N_2230,N_1712,N_1262);
xnor U2231 (N_2231,N_1748,N_1835);
nand U2232 (N_2232,N_1692,N_1905);
nand U2233 (N_2233,N_1926,N_1348);
and U2234 (N_2234,In_1045,N_1014);
or U2235 (N_2235,N_1988,N_1914);
and U2236 (N_2236,N_1870,N_898);
nand U2237 (N_2237,N_1929,N_1635);
nand U2238 (N_2238,N_1562,N_1987);
xor U2239 (N_2239,N_1231,N_1552);
and U2240 (N_2240,N_1291,N_1850);
and U2241 (N_2241,N_1678,N_1651);
and U2242 (N_2242,N_1861,N_1783);
xor U2243 (N_2243,N_1810,N_1788);
and U2244 (N_2244,N_1377,N_1918);
or U2245 (N_2245,In_451,N_1891);
and U2246 (N_2246,In_2192,N_1976);
nor U2247 (N_2247,N_1832,N_1958);
nand U2248 (N_2248,N_1971,N_1834);
nor U2249 (N_2249,N_1382,N_1813);
nor U2250 (N_2250,N_2166,N_2041);
xnor U2251 (N_2251,N_2104,N_2008);
xnor U2252 (N_2252,N_2034,N_2130);
and U2253 (N_2253,N_2098,N_2022);
nand U2254 (N_2254,N_2118,N_2047);
xor U2255 (N_2255,N_2190,N_2147);
nor U2256 (N_2256,N_2249,N_2197);
nand U2257 (N_2257,N_2066,N_2240);
xor U2258 (N_2258,N_2242,N_2173);
xor U2259 (N_2259,N_2110,N_2241);
nor U2260 (N_2260,N_2208,N_2164);
nor U2261 (N_2261,N_2096,N_2117);
nor U2262 (N_2262,N_2060,N_2079);
and U2263 (N_2263,N_2187,N_2089);
or U2264 (N_2264,N_2039,N_2019);
nand U2265 (N_2265,N_2140,N_2206);
or U2266 (N_2266,N_2188,N_2105);
xnor U2267 (N_2267,N_2185,N_2091);
xor U2268 (N_2268,N_2076,N_2014);
nor U2269 (N_2269,N_2239,N_2113);
or U2270 (N_2270,N_2026,N_2128);
or U2271 (N_2271,N_2148,N_2201);
nor U2272 (N_2272,N_2005,N_2044);
or U2273 (N_2273,N_2143,N_2061);
nand U2274 (N_2274,N_2040,N_2176);
and U2275 (N_2275,N_2112,N_2174);
and U2276 (N_2276,N_2013,N_2156);
xor U2277 (N_2277,N_2198,N_2139);
or U2278 (N_2278,N_2202,N_2043);
and U2279 (N_2279,N_2238,N_2230);
xnor U2280 (N_2280,N_2102,N_2232);
nor U2281 (N_2281,N_2015,N_2046);
or U2282 (N_2282,N_2036,N_2167);
or U2283 (N_2283,N_2215,N_2233);
nor U2284 (N_2284,N_2067,N_2161);
nand U2285 (N_2285,N_2035,N_2146);
xnor U2286 (N_2286,N_2149,N_2171);
and U2287 (N_2287,N_2042,N_2012);
or U2288 (N_2288,N_2010,N_2134);
or U2289 (N_2289,N_2062,N_2017);
and U2290 (N_2290,N_2184,N_2055);
or U2291 (N_2291,N_2109,N_2170);
xor U2292 (N_2292,N_2068,N_2065);
nand U2293 (N_2293,N_2211,N_2021);
nand U2294 (N_2294,N_2219,N_2051);
nor U2295 (N_2295,N_2237,N_2155);
nor U2296 (N_2296,N_2133,N_2119);
nand U2297 (N_2297,N_2037,N_2057);
nor U2298 (N_2298,N_2194,N_2003);
and U2299 (N_2299,N_2154,N_2178);
and U2300 (N_2300,N_2220,N_2050);
or U2301 (N_2301,N_2081,N_2231);
and U2302 (N_2302,N_2029,N_2053);
xor U2303 (N_2303,N_2214,N_2045);
and U2304 (N_2304,N_2180,N_2225);
nor U2305 (N_2305,N_2204,N_2024);
nand U2306 (N_2306,N_2120,N_2129);
nor U2307 (N_2307,N_2115,N_2209);
xnor U2308 (N_2308,N_2189,N_2123);
nor U2309 (N_2309,N_2028,N_2126);
and U2310 (N_2310,N_2131,N_2136);
and U2311 (N_2311,N_2116,N_2175);
or U2312 (N_2312,N_2049,N_2246);
nor U2313 (N_2313,N_2100,N_2199);
or U2314 (N_2314,N_2072,N_2210);
or U2315 (N_2315,N_2004,N_2226);
nor U2316 (N_2316,N_2075,N_2030);
nand U2317 (N_2317,N_2200,N_2111);
and U2318 (N_2318,N_2218,N_2077);
xor U2319 (N_2319,N_2088,N_2195);
nor U2320 (N_2320,N_2153,N_2070);
nand U2321 (N_2321,N_2172,N_2223);
nor U2322 (N_2322,N_2138,N_2092);
xor U2323 (N_2323,N_2179,N_2063);
nand U2324 (N_2324,N_2144,N_2157);
xor U2325 (N_2325,N_2247,N_2001);
nor U2326 (N_2326,N_2192,N_2141);
nor U2327 (N_2327,N_2058,N_2186);
and U2328 (N_2328,N_2074,N_2221);
nor U2329 (N_2329,N_2127,N_2248);
nor U2330 (N_2330,N_2064,N_2224);
nor U2331 (N_2331,N_2071,N_2243);
or U2332 (N_2332,N_2181,N_2083);
or U2333 (N_2333,N_2025,N_2011);
nand U2334 (N_2334,N_2033,N_2007);
nand U2335 (N_2335,N_2087,N_2158);
nand U2336 (N_2336,N_2016,N_2227);
and U2337 (N_2337,N_2152,N_2082);
nand U2338 (N_2338,N_2228,N_2205);
nor U2339 (N_2339,N_2160,N_2121);
and U2340 (N_2340,N_2142,N_2085);
xnor U2341 (N_2341,N_2137,N_2031);
nand U2342 (N_2342,N_2101,N_2132);
and U2343 (N_2343,N_2145,N_2073);
and U2344 (N_2344,N_2162,N_2163);
and U2345 (N_2345,N_2094,N_2222);
nor U2346 (N_2346,N_2125,N_2084);
and U2347 (N_2347,N_2108,N_2122);
or U2348 (N_2348,N_2165,N_2095);
and U2349 (N_2349,N_2207,N_2052);
and U2350 (N_2350,N_2135,N_2229);
or U2351 (N_2351,N_2032,N_2103);
and U2352 (N_2352,N_2234,N_2150);
xor U2353 (N_2353,N_2183,N_2099);
and U2354 (N_2354,N_2000,N_2245);
nand U2355 (N_2355,N_2023,N_2191);
and U2356 (N_2356,N_2054,N_2124);
or U2357 (N_2357,N_2107,N_2006);
nor U2358 (N_2358,N_2151,N_2217);
xor U2359 (N_2359,N_2193,N_2048);
and U2360 (N_2360,N_2086,N_2018);
and U2361 (N_2361,N_2114,N_2236);
and U2362 (N_2362,N_2027,N_2056);
nor U2363 (N_2363,N_2020,N_2213);
nand U2364 (N_2364,N_2168,N_2080);
or U2365 (N_2365,N_2009,N_2002);
and U2366 (N_2366,N_2097,N_2177);
xor U2367 (N_2367,N_2196,N_2159);
nor U2368 (N_2368,N_2203,N_2182);
nand U2369 (N_2369,N_2244,N_2078);
nand U2370 (N_2370,N_2106,N_2216);
nand U2371 (N_2371,N_2090,N_2069);
xor U2372 (N_2372,N_2235,N_2212);
nor U2373 (N_2373,N_2093,N_2169);
nor U2374 (N_2374,N_2059,N_2038);
and U2375 (N_2375,N_2213,N_2111);
or U2376 (N_2376,N_2210,N_2048);
nor U2377 (N_2377,N_2219,N_2099);
or U2378 (N_2378,N_2103,N_2156);
or U2379 (N_2379,N_2052,N_2159);
or U2380 (N_2380,N_2027,N_2124);
and U2381 (N_2381,N_2229,N_2161);
or U2382 (N_2382,N_2182,N_2004);
nand U2383 (N_2383,N_2074,N_2160);
nor U2384 (N_2384,N_2199,N_2237);
or U2385 (N_2385,N_2044,N_2086);
and U2386 (N_2386,N_2049,N_2182);
nand U2387 (N_2387,N_2052,N_2214);
xor U2388 (N_2388,N_2207,N_2233);
nand U2389 (N_2389,N_2189,N_2021);
xnor U2390 (N_2390,N_2206,N_2138);
xor U2391 (N_2391,N_2065,N_2004);
xnor U2392 (N_2392,N_2093,N_2136);
and U2393 (N_2393,N_2241,N_2048);
xnor U2394 (N_2394,N_2158,N_2016);
nand U2395 (N_2395,N_2103,N_2016);
or U2396 (N_2396,N_2144,N_2222);
xnor U2397 (N_2397,N_2153,N_2043);
nor U2398 (N_2398,N_2241,N_2002);
nor U2399 (N_2399,N_2115,N_2095);
and U2400 (N_2400,N_2045,N_2031);
or U2401 (N_2401,N_2227,N_2081);
nand U2402 (N_2402,N_2161,N_2021);
nor U2403 (N_2403,N_2220,N_2035);
xor U2404 (N_2404,N_2185,N_2105);
or U2405 (N_2405,N_2122,N_2106);
xor U2406 (N_2406,N_2147,N_2230);
or U2407 (N_2407,N_2001,N_2227);
nand U2408 (N_2408,N_2118,N_2040);
xnor U2409 (N_2409,N_2025,N_2040);
nor U2410 (N_2410,N_2060,N_2014);
or U2411 (N_2411,N_2242,N_2101);
or U2412 (N_2412,N_2158,N_2077);
xor U2413 (N_2413,N_2047,N_2014);
nor U2414 (N_2414,N_2184,N_2138);
nand U2415 (N_2415,N_2194,N_2114);
nor U2416 (N_2416,N_2064,N_2025);
and U2417 (N_2417,N_2032,N_2041);
xnor U2418 (N_2418,N_2206,N_2110);
and U2419 (N_2419,N_2194,N_2201);
or U2420 (N_2420,N_2127,N_2025);
and U2421 (N_2421,N_2188,N_2164);
nand U2422 (N_2422,N_2114,N_2046);
xnor U2423 (N_2423,N_2189,N_2197);
nand U2424 (N_2424,N_2143,N_2029);
and U2425 (N_2425,N_2186,N_2195);
nand U2426 (N_2426,N_2067,N_2014);
nor U2427 (N_2427,N_2078,N_2108);
and U2428 (N_2428,N_2241,N_2018);
nor U2429 (N_2429,N_2168,N_2079);
xnor U2430 (N_2430,N_2155,N_2214);
and U2431 (N_2431,N_2018,N_2056);
or U2432 (N_2432,N_2007,N_2129);
or U2433 (N_2433,N_2200,N_2244);
xor U2434 (N_2434,N_2175,N_2079);
and U2435 (N_2435,N_2144,N_2136);
or U2436 (N_2436,N_2239,N_2003);
and U2437 (N_2437,N_2235,N_2130);
nor U2438 (N_2438,N_2183,N_2234);
nand U2439 (N_2439,N_2190,N_2179);
or U2440 (N_2440,N_2095,N_2079);
and U2441 (N_2441,N_2058,N_2207);
nand U2442 (N_2442,N_2031,N_2127);
or U2443 (N_2443,N_2193,N_2091);
nor U2444 (N_2444,N_2040,N_2183);
xnor U2445 (N_2445,N_2070,N_2204);
and U2446 (N_2446,N_2025,N_2152);
or U2447 (N_2447,N_2144,N_2060);
nor U2448 (N_2448,N_2235,N_2018);
nor U2449 (N_2449,N_2001,N_2047);
xnor U2450 (N_2450,N_2070,N_2108);
xor U2451 (N_2451,N_2205,N_2240);
or U2452 (N_2452,N_2005,N_2199);
and U2453 (N_2453,N_2068,N_2187);
nand U2454 (N_2454,N_2028,N_2078);
or U2455 (N_2455,N_2178,N_2063);
nor U2456 (N_2456,N_2121,N_2224);
or U2457 (N_2457,N_2074,N_2205);
and U2458 (N_2458,N_2039,N_2027);
or U2459 (N_2459,N_2153,N_2000);
nor U2460 (N_2460,N_2244,N_2176);
nor U2461 (N_2461,N_2054,N_2120);
or U2462 (N_2462,N_2013,N_2000);
or U2463 (N_2463,N_2171,N_2148);
xnor U2464 (N_2464,N_2199,N_2115);
nand U2465 (N_2465,N_2004,N_2171);
nand U2466 (N_2466,N_2113,N_2068);
or U2467 (N_2467,N_2033,N_2166);
and U2468 (N_2468,N_2024,N_2009);
nand U2469 (N_2469,N_2068,N_2179);
and U2470 (N_2470,N_2184,N_2075);
xnor U2471 (N_2471,N_2230,N_2057);
nor U2472 (N_2472,N_2187,N_2201);
and U2473 (N_2473,N_2011,N_2073);
nor U2474 (N_2474,N_2177,N_2017);
nor U2475 (N_2475,N_2118,N_2135);
nand U2476 (N_2476,N_2230,N_2154);
and U2477 (N_2477,N_2065,N_2013);
nand U2478 (N_2478,N_2071,N_2111);
nand U2479 (N_2479,N_2172,N_2234);
nor U2480 (N_2480,N_2212,N_2036);
nor U2481 (N_2481,N_2091,N_2123);
xor U2482 (N_2482,N_2047,N_2150);
and U2483 (N_2483,N_2229,N_2151);
nor U2484 (N_2484,N_2235,N_2207);
nand U2485 (N_2485,N_2195,N_2096);
xnor U2486 (N_2486,N_2012,N_2143);
xor U2487 (N_2487,N_2109,N_2047);
nand U2488 (N_2488,N_2139,N_2212);
and U2489 (N_2489,N_2174,N_2040);
nor U2490 (N_2490,N_2227,N_2025);
and U2491 (N_2491,N_2015,N_2060);
xor U2492 (N_2492,N_2001,N_2093);
and U2493 (N_2493,N_2038,N_2064);
nor U2494 (N_2494,N_2140,N_2090);
xnor U2495 (N_2495,N_2241,N_2183);
nand U2496 (N_2496,N_2166,N_2072);
and U2497 (N_2497,N_2054,N_2101);
nor U2498 (N_2498,N_2206,N_2182);
or U2499 (N_2499,N_2061,N_2229);
or U2500 (N_2500,N_2286,N_2295);
and U2501 (N_2501,N_2478,N_2486);
and U2502 (N_2502,N_2407,N_2428);
nand U2503 (N_2503,N_2418,N_2458);
xnor U2504 (N_2504,N_2332,N_2391);
nand U2505 (N_2505,N_2450,N_2366);
and U2506 (N_2506,N_2386,N_2406);
and U2507 (N_2507,N_2467,N_2440);
xor U2508 (N_2508,N_2419,N_2466);
nand U2509 (N_2509,N_2349,N_2373);
nand U2510 (N_2510,N_2287,N_2359);
and U2511 (N_2511,N_2367,N_2452);
nor U2512 (N_2512,N_2446,N_2432);
and U2513 (N_2513,N_2459,N_2252);
or U2514 (N_2514,N_2380,N_2454);
and U2515 (N_2515,N_2263,N_2365);
or U2516 (N_2516,N_2494,N_2405);
nand U2517 (N_2517,N_2377,N_2370);
xnor U2518 (N_2518,N_2299,N_2338);
xnor U2519 (N_2519,N_2499,N_2296);
nand U2520 (N_2520,N_2308,N_2497);
nand U2521 (N_2521,N_2357,N_2465);
nand U2522 (N_2522,N_2268,N_2328);
xor U2523 (N_2523,N_2279,N_2425);
nand U2524 (N_2524,N_2256,N_2290);
xnor U2525 (N_2525,N_2480,N_2468);
xnor U2526 (N_2526,N_2420,N_2255);
nand U2527 (N_2527,N_2471,N_2309);
nand U2528 (N_2528,N_2430,N_2378);
or U2529 (N_2529,N_2444,N_2447);
or U2530 (N_2530,N_2489,N_2383);
xnor U2531 (N_2531,N_2475,N_2469);
nand U2532 (N_2532,N_2451,N_2395);
and U2533 (N_2533,N_2305,N_2384);
xor U2534 (N_2534,N_2336,N_2352);
nand U2535 (N_2535,N_2254,N_2498);
nand U2536 (N_2536,N_2262,N_2260);
and U2537 (N_2537,N_2462,N_2483);
or U2538 (N_2538,N_2368,N_2424);
or U2539 (N_2539,N_2429,N_2421);
xor U2540 (N_2540,N_2344,N_2341);
nand U2541 (N_2541,N_2314,N_2297);
and U2542 (N_2542,N_2481,N_2253);
xnor U2543 (N_2543,N_2404,N_2310);
xnor U2544 (N_2544,N_2283,N_2281);
and U2545 (N_2545,N_2294,N_2382);
xnor U2546 (N_2546,N_2449,N_2259);
nand U2547 (N_2547,N_2330,N_2251);
or U2548 (N_2548,N_2379,N_2324);
nor U2549 (N_2549,N_2398,N_2397);
nor U2550 (N_2550,N_2306,N_2414);
and U2551 (N_2551,N_2322,N_2453);
or U2552 (N_2552,N_2436,N_2304);
and U2553 (N_2553,N_2413,N_2394);
or U2554 (N_2554,N_2257,N_2291);
nor U2555 (N_2555,N_2474,N_2354);
nor U2556 (N_2556,N_2280,N_2327);
xor U2557 (N_2557,N_2312,N_2340);
nor U2558 (N_2558,N_2393,N_2445);
and U2559 (N_2559,N_2267,N_2288);
nor U2560 (N_2560,N_2434,N_2401);
nor U2561 (N_2561,N_2261,N_2250);
xor U2562 (N_2562,N_2316,N_2266);
and U2563 (N_2563,N_2361,N_2326);
nand U2564 (N_2564,N_2273,N_2301);
nor U2565 (N_2565,N_2318,N_2276);
or U2566 (N_2566,N_2388,N_2456);
nand U2567 (N_2567,N_2321,N_2369);
or U2568 (N_2568,N_2496,N_2319);
nor U2569 (N_2569,N_2493,N_2345);
nand U2570 (N_2570,N_2313,N_2325);
nand U2571 (N_2571,N_2356,N_2351);
nor U2572 (N_2572,N_2265,N_2409);
xor U2573 (N_2573,N_2358,N_2435);
nor U2574 (N_2574,N_2355,N_2311);
xnor U2575 (N_2575,N_2390,N_2392);
and U2576 (N_2576,N_2269,N_2285);
or U2577 (N_2577,N_2375,N_2270);
nor U2578 (N_2578,N_2300,N_2282);
nor U2579 (N_2579,N_2439,N_2289);
xnor U2580 (N_2580,N_2482,N_2426);
or U2581 (N_2581,N_2396,N_2350);
or U2582 (N_2582,N_2317,N_2362);
nand U2583 (N_2583,N_2277,N_2479);
xor U2584 (N_2584,N_2408,N_2463);
xnor U2585 (N_2585,N_2376,N_2477);
nand U2586 (N_2586,N_2353,N_2364);
or U2587 (N_2587,N_2472,N_2323);
nand U2588 (N_2588,N_2258,N_2455);
or U2589 (N_2589,N_2381,N_2272);
xnor U2590 (N_2590,N_2491,N_2416);
nand U2591 (N_2591,N_2422,N_2303);
and U2592 (N_2592,N_2410,N_2438);
nor U2593 (N_2593,N_2363,N_2320);
or U2594 (N_2594,N_2484,N_2389);
or U2595 (N_2595,N_2400,N_2271);
or U2596 (N_2596,N_2337,N_2315);
nor U2597 (N_2597,N_2431,N_2264);
and U2598 (N_2598,N_2293,N_2298);
or U2599 (N_2599,N_2448,N_2348);
xnor U2600 (N_2600,N_2307,N_2284);
nor U2601 (N_2601,N_2411,N_2490);
and U2602 (N_2602,N_2342,N_2360);
xor U2603 (N_2603,N_2335,N_2457);
xor U2604 (N_2604,N_2334,N_2331);
and U2605 (N_2605,N_2464,N_2415);
and U2606 (N_2606,N_2492,N_2274);
nand U2607 (N_2607,N_2488,N_2374);
nand U2608 (N_2608,N_2402,N_2371);
and U2609 (N_2609,N_2346,N_2433);
nand U2610 (N_2610,N_2372,N_2275);
or U2611 (N_2611,N_2403,N_2476);
nor U2612 (N_2612,N_2443,N_2302);
and U2613 (N_2613,N_2292,N_2495);
xnor U2614 (N_2614,N_2437,N_2427);
nor U2615 (N_2615,N_2470,N_2399);
nor U2616 (N_2616,N_2343,N_2333);
xor U2617 (N_2617,N_2485,N_2329);
and U2618 (N_2618,N_2347,N_2423);
nor U2619 (N_2619,N_2385,N_2487);
nor U2620 (N_2620,N_2412,N_2339);
xor U2621 (N_2621,N_2387,N_2442);
or U2622 (N_2622,N_2461,N_2417);
and U2623 (N_2623,N_2441,N_2473);
and U2624 (N_2624,N_2460,N_2278);
or U2625 (N_2625,N_2474,N_2337);
or U2626 (N_2626,N_2484,N_2347);
or U2627 (N_2627,N_2348,N_2485);
nand U2628 (N_2628,N_2373,N_2385);
or U2629 (N_2629,N_2281,N_2274);
nand U2630 (N_2630,N_2420,N_2402);
and U2631 (N_2631,N_2320,N_2269);
nand U2632 (N_2632,N_2378,N_2338);
or U2633 (N_2633,N_2297,N_2471);
nor U2634 (N_2634,N_2384,N_2298);
nand U2635 (N_2635,N_2341,N_2454);
and U2636 (N_2636,N_2433,N_2259);
or U2637 (N_2637,N_2372,N_2387);
nand U2638 (N_2638,N_2250,N_2424);
or U2639 (N_2639,N_2371,N_2422);
xnor U2640 (N_2640,N_2258,N_2320);
or U2641 (N_2641,N_2267,N_2394);
nor U2642 (N_2642,N_2412,N_2291);
xor U2643 (N_2643,N_2314,N_2443);
xor U2644 (N_2644,N_2325,N_2266);
or U2645 (N_2645,N_2285,N_2275);
xnor U2646 (N_2646,N_2404,N_2352);
nand U2647 (N_2647,N_2484,N_2447);
or U2648 (N_2648,N_2255,N_2443);
xor U2649 (N_2649,N_2414,N_2402);
or U2650 (N_2650,N_2391,N_2395);
nor U2651 (N_2651,N_2462,N_2396);
xor U2652 (N_2652,N_2261,N_2492);
nor U2653 (N_2653,N_2313,N_2395);
xor U2654 (N_2654,N_2316,N_2445);
and U2655 (N_2655,N_2360,N_2434);
and U2656 (N_2656,N_2340,N_2472);
nand U2657 (N_2657,N_2487,N_2287);
xnor U2658 (N_2658,N_2457,N_2303);
nand U2659 (N_2659,N_2272,N_2368);
xor U2660 (N_2660,N_2277,N_2320);
and U2661 (N_2661,N_2382,N_2340);
and U2662 (N_2662,N_2380,N_2363);
and U2663 (N_2663,N_2322,N_2314);
nor U2664 (N_2664,N_2388,N_2404);
nand U2665 (N_2665,N_2337,N_2466);
nand U2666 (N_2666,N_2419,N_2474);
nand U2667 (N_2667,N_2447,N_2264);
xor U2668 (N_2668,N_2420,N_2496);
xnor U2669 (N_2669,N_2383,N_2403);
or U2670 (N_2670,N_2260,N_2449);
and U2671 (N_2671,N_2272,N_2359);
nor U2672 (N_2672,N_2312,N_2390);
or U2673 (N_2673,N_2287,N_2486);
xnor U2674 (N_2674,N_2371,N_2349);
nand U2675 (N_2675,N_2379,N_2436);
or U2676 (N_2676,N_2356,N_2419);
nand U2677 (N_2677,N_2268,N_2337);
xnor U2678 (N_2678,N_2464,N_2325);
nor U2679 (N_2679,N_2489,N_2317);
nand U2680 (N_2680,N_2389,N_2408);
and U2681 (N_2681,N_2312,N_2333);
or U2682 (N_2682,N_2364,N_2259);
nand U2683 (N_2683,N_2492,N_2377);
or U2684 (N_2684,N_2435,N_2498);
xor U2685 (N_2685,N_2268,N_2359);
nand U2686 (N_2686,N_2460,N_2363);
nand U2687 (N_2687,N_2346,N_2438);
xor U2688 (N_2688,N_2297,N_2269);
nor U2689 (N_2689,N_2351,N_2489);
and U2690 (N_2690,N_2352,N_2422);
nand U2691 (N_2691,N_2357,N_2425);
and U2692 (N_2692,N_2419,N_2338);
nand U2693 (N_2693,N_2426,N_2430);
xor U2694 (N_2694,N_2264,N_2479);
xnor U2695 (N_2695,N_2349,N_2329);
nand U2696 (N_2696,N_2465,N_2344);
nand U2697 (N_2697,N_2423,N_2331);
and U2698 (N_2698,N_2301,N_2492);
or U2699 (N_2699,N_2428,N_2429);
nand U2700 (N_2700,N_2270,N_2372);
nor U2701 (N_2701,N_2446,N_2442);
xnor U2702 (N_2702,N_2408,N_2282);
or U2703 (N_2703,N_2349,N_2359);
xnor U2704 (N_2704,N_2365,N_2439);
xor U2705 (N_2705,N_2278,N_2410);
nand U2706 (N_2706,N_2427,N_2250);
nand U2707 (N_2707,N_2334,N_2290);
or U2708 (N_2708,N_2344,N_2260);
and U2709 (N_2709,N_2365,N_2479);
nand U2710 (N_2710,N_2409,N_2411);
nor U2711 (N_2711,N_2383,N_2379);
nand U2712 (N_2712,N_2445,N_2262);
or U2713 (N_2713,N_2475,N_2442);
nand U2714 (N_2714,N_2424,N_2299);
and U2715 (N_2715,N_2356,N_2263);
nand U2716 (N_2716,N_2442,N_2406);
xor U2717 (N_2717,N_2288,N_2339);
and U2718 (N_2718,N_2449,N_2464);
and U2719 (N_2719,N_2494,N_2265);
xor U2720 (N_2720,N_2440,N_2348);
xnor U2721 (N_2721,N_2267,N_2386);
xnor U2722 (N_2722,N_2354,N_2255);
nor U2723 (N_2723,N_2274,N_2266);
or U2724 (N_2724,N_2299,N_2479);
or U2725 (N_2725,N_2404,N_2372);
nand U2726 (N_2726,N_2390,N_2374);
nor U2727 (N_2727,N_2418,N_2282);
nor U2728 (N_2728,N_2481,N_2379);
or U2729 (N_2729,N_2352,N_2324);
nor U2730 (N_2730,N_2314,N_2409);
xnor U2731 (N_2731,N_2326,N_2388);
and U2732 (N_2732,N_2303,N_2382);
nor U2733 (N_2733,N_2369,N_2354);
nor U2734 (N_2734,N_2343,N_2444);
nor U2735 (N_2735,N_2300,N_2478);
or U2736 (N_2736,N_2364,N_2466);
or U2737 (N_2737,N_2443,N_2490);
nand U2738 (N_2738,N_2464,N_2421);
and U2739 (N_2739,N_2332,N_2483);
nor U2740 (N_2740,N_2260,N_2308);
xor U2741 (N_2741,N_2478,N_2396);
and U2742 (N_2742,N_2317,N_2426);
or U2743 (N_2743,N_2433,N_2287);
nor U2744 (N_2744,N_2292,N_2277);
xor U2745 (N_2745,N_2385,N_2360);
nand U2746 (N_2746,N_2456,N_2283);
and U2747 (N_2747,N_2308,N_2467);
xor U2748 (N_2748,N_2300,N_2464);
or U2749 (N_2749,N_2300,N_2426);
and U2750 (N_2750,N_2691,N_2528);
nand U2751 (N_2751,N_2696,N_2652);
nand U2752 (N_2752,N_2705,N_2697);
xor U2753 (N_2753,N_2559,N_2560);
nand U2754 (N_2754,N_2586,N_2719);
or U2755 (N_2755,N_2737,N_2583);
or U2756 (N_2756,N_2684,N_2722);
or U2757 (N_2757,N_2510,N_2748);
and U2758 (N_2758,N_2610,N_2533);
or U2759 (N_2759,N_2595,N_2516);
nand U2760 (N_2760,N_2596,N_2635);
nand U2761 (N_2761,N_2524,N_2725);
xnor U2762 (N_2762,N_2709,N_2732);
nor U2763 (N_2763,N_2633,N_2518);
and U2764 (N_2764,N_2541,N_2517);
nor U2765 (N_2765,N_2542,N_2745);
nor U2766 (N_2766,N_2642,N_2543);
xnor U2767 (N_2767,N_2508,N_2630);
nand U2768 (N_2768,N_2694,N_2550);
nand U2769 (N_2769,N_2599,N_2655);
or U2770 (N_2770,N_2706,N_2601);
or U2771 (N_2771,N_2502,N_2673);
nor U2772 (N_2772,N_2628,N_2643);
nor U2773 (N_2773,N_2576,N_2572);
and U2774 (N_2774,N_2639,N_2519);
and U2775 (N_2775,N_2648,N_2733);
or U2776 (N_2776,N_2615,N_2536);
xor U2777 (N_2777,N_2638,N_2581);
and U2778 (N_2778,N_2570,N_2677);
nand U2779 (N_2779,N_2703,N_2564);
xnor U2780 (N_2780,N_2501,N_2651);
and U2781 (N_2781,N_2503,N_2580);
or U2782 (N_2782,N_2558,N_2627);
or U2783 (N_2783,N_2674,N_2568);
xor U2784 (N_2784,N_2654,N_2623);
and U2785 (N_2785,N_2529,N_2688);
xor U2786 (N_2786,N_2574,N_2571);
and U2787 (N_2787,N_2675,N_2613);
nand U2788 (N_2788,N_2577,N_2511);
nand U2789 (N_2789,N_2585,N_2681);
xnor U2790 (N_2790,N_2605,N_2515);
xnor U2791 (N_2791,N_2620,N_2552);
or U2792 (N_2792,N_2584,N_2589);
nor U2793 (N_2793,N_2742,N_2665);
nor U2794 (N_2794,N_2602,N_2726);
xor U2795 (N_2795,N_2637,N_2707);
nand U2796 (N_2796,N_2539,N_2606);
xnor U2797 (N_2797,N_2693,N_2700);
nor U2798 (N_2798,N_2640,N_2649);
and U2799 (N_2799,N_2616,N_2553);
or U2800 (N_2800,N_2666,N_2522);
xnor U2801 (N_2801,N_2582,N_2561);
nor U2802 (N_2802,N_2590,N_2715);
or U2803 (N_2803,N_2658,N_2540);
or U2804 (N_2804,N_2532,N_2609);
or U2805 (N_2805,N_2721,N_2668);
or U2806 (N_2806,N_2617,N_2634);
nand U2807 (N_2807,N_2593,N_2548);
xnor U2808 (N_2808,N_2619,N_2743);
and U2809 (N_2809,N_2685,N_2738);
or U2810 (N_2810,N_2611,N_2514);
xnor U2811 (N_2811,N_2579,N_2641);
or U2812 (N_2812,N_2698,N_2664);
or U2813 (N_2813,N_2712,N_2736);
xor U2814 (N_2814,N_2672,N_2646);
and U2815 (N_2815,N_2746,N_2573);
nand U2816 (N_2816,N_2505,N_2661);
or U2817 (N_2817,N_2520,N_2594);
or U2818 (N_2818,N_2671,N_2740);
nor U2819 (N_2819,N_2718,N_2538);
and U2820 (N_2820,N_2592,N_2667);
nand U2821 (N_2821,N_2544,N_2534);
nor U2822 (N_2822,N_2565,N_2631);
and U2823 (N_2823,N_2527,N_2720);
nand U2824 (N_2824,N_2625,N_2555);
xor U2825 (N_2825,N_2551,N_2608);
nand U2826 (N_2826,N_2699,N_2506);
xnor U2827 (N_2827,N_2702,N_2566);
xor U2828 (N_2828,N_2537,N_2734);
nor U2829 (N_2829,N_2717,N_2644);
or U2830 (N_2830,N_2670,N_2597);
nor U2831 (N_2831,N_2530,N_2682);
xnor U2832 (N_2832,N_2679,N_2730);
nand U2833 (N_2833,N_2744,N_2612);
nor U2834 (N_2834,N_2728,N_2741);
and U2835 (N_2835,N_2739,N_2632);
and U2836 (N_2836,N_2687,N_2624);
or U2837 (N_2837,N_2735,N_2607);
or U2838 (N_2838,N_2513,N_2567);
or U2839 (N_2839,N_2680,N_2659);
xnor U2840 (N_2840,N_2747,N_2525);
nand U2841 (N_2841,N_2692,N_2587);
nand U2842 (N_2842,N_2531,N_2678);
nor U2843 (N_2843,N_2621,N_2663);
nor U2844 (N_2844,N_2500,N_2588);
xor U2845 (N_2845,N_2556,N_2554);
and U2846 (N_2846,N_2669,N_2727);
nand U2847 (N_2847,N_2578,N_2563);
and U2848 (N_2848,N_2729,N_2504);
or U2849 (N_2849,N_2662,N_2686);
or U2850 (N_2850,N_2710,N_2690);
and U2851 (N_2851,N_2647,N_2521);
xor U2852 (N_2852,N_2749,N_2598);
or U2853 (N_2853,N_2731,N_2545);
or U2854 (N_2854,N_2626,N_2660);
or U2855 (N_2855,N_2603,N_2557);
nand U2856 (N_2856,N_2509,N_2512);
nor U2857 (N_2857,N_2629,N_2591);
or U2858 (N_2858,N_2657,N_2711);
xnor U2859 (N_2859,N_2604,N_2683);
or U2860 (N_2860,N_2562,N_2704);
nand U2861 (N_2861,N_2645,N_2546);
or U2862 (N_2862,N_2714,N_2653);
xor U2863 (N_2863,N_2689,N_2575);
nand U2864 (N_2864,N_2614,N_2600);
xor U2865 (N_2865,N_2656,N_2724);
nand U2866 (N_2866,N_2547,N_2708);
or U2867 (N_2867,N_2526,N_2535);
and U2868 (N_2868,N_2622,N_2676);
xor U2869 (N_2869,N_2650,N_2716);
nand U2870 (N_2870,N_2507,N_2695);
xnor U2871 (N_2871,N_2569,N_2549);
and U2872 (N_2872,N_2701,N_2636);
xor U2873 (N_2873,N_2618,N_2523);
nor U2874 (N_2874,N_2723,N_2713);
nor U2875 (N_2875,N_2639,N_2602);
xnor U2876 (N_2876,N_2583,N_2604);
nand U2877 (N_2877,N_2704,N_2620);
nand U2878 (N_2878,N_2617,N_2736);
nor U2879 (N_2879,N_2613,N_2506);
or U2880 (N_2880,N_2537,N_2716);
and U2881 (N_2881,N_2541,N_2731);
nor U2882 (N_2882,N_2681,N_2588);
xor U2883 (N_2883,N_2599,N_2564);
xnor U2884 (N_2884,N_2686,N_2530);
and U2885 (N_2885,N_2722,N_2713);
or U2886 (N_2886,N_2500,N_2657);
nor U2887 (N_2887,N_2725,N_2531);
nor U2888 (N_2888,N_2693,N_2554);
nor U2889 (N_2889,N_2711,N_2505);
nor U2890 (N_2890,N_2722,N_2579);
nor U2891 (N_2891,N_2674,N_2678);
and U2892 (N_2892,N_2557,N_2606);
xnor U2893 (N_2893,N_2665,N_2647);
xnor U2894 (N_2894,N_2645,N_2713);
and U2895 (N_2895,N_2500,N_2624);
nand U2896 (N_2896,N_2567,N_2733);
nor U2897 (N_2897,N_2669,N_2700);
nand U2898 (N_2898,N_2606,N_2611);
nand U2899 (N_2899,N_2585,N_2616);
nand U2900 (N_2900,N_2525,N_2542);
xnor U2901 (N_2901,N_2644,N_2576);
nand U2902 (N_2902,N_2587,N_2715);
xnor U2903 (N_2903,N_2651,N_2652);
nor U2904 (N_2904,N_2506,N_2720);
nand U2905 (N_2905,N_2621,N_2716);
or U2906 (N_2906,N_2673,N_2672);
and U2907 (N_2907,N_2631,N_2670);
xnor U2908 (N_2908,N_2679,N_2646);
nand U2909 (N_2909,N_2606,N_2640);
or U2910 (N_2910,N_2726,N_2501);
xnor U2911 (N_2911,N_2714,N_2676);
nor U2912 (N_2912,N_2577,N_2657);
nand U2913 (N_2913,N_2605,N_2568);
xnor U2914 (N_2914,N_2572,N_2557);
or U2915 (N_2915,N_2738,N_2587);
and U2916 (N_2916,N_2702,N_2742);
or U2917 (N_2917,N_2537,N_2502);
or U2918 (N_2918,N_2647,N_2505);
nor U2919 (N_2919,N_2647,N_2704);
or U2920 (N_2920,N_2700,N_2505);
nor U2921 (N_2921,N_2592,N_2523);
or U2922 (N_2922,N_2647,N_2509);
or U2923 (N_2923,N_2550,N_2625);
nand U2924 (N_2924,N_2738,N_2743);
xor U2925 (N_2925,N_2664,N_2715);
xnor U2926 (N_2926,N_2523,N_2694);
or U2927 (N_2927,N_2577,N_2559);
or U2928 (N_2928,N_2703,N_2714);
or U2929 (N_2929,N_2508,N_2600);
nand U2930 (N_2930,N_2582,N_2646);
or U2931 (N_2931,N_2603,N_2658);
and U2932 (N_2932,N_2746,N_2618);
and U2933 (N_2933,N_2528,N_2588);
nor U2934 (N_2934,N_2564,N_2663);
xor U2935 (N_2935,N_2732,N_2617);
xor U2936 (N_2936,N_2597,N_2669);
nand U2937 (N_2937,N_2531,N_2726);
and U2938 (N_2938,N_2519,N_2682);
xnor U2939 (N_2939,N_2570,N_2608);
or U2940 (N_2940,N_2671,N_2652);
nor U2941 (N_2941,N_2507,N_2543);
and U2942 (N_2942,N_2637,N_2739);
nor U2943 (N_2943,N_2586,N_2707);
nand U2944 (N_2944,N_2673,N_2725);
and U2945 (N_2945,N_2643,N_2600);
nand U2946 (N_2946,N_2545,N_2500);
xor U2947 (N_2947,N_2549,N_2583);
or U2948 (N_2948,N_2684,N_2627);
nor U2949 (N_2949,N_2577,N_2528);
xor U2950 (N_2950,N_2715,N_2537);
nand U2951 (N_2951,N_2515,N_2607);
and U2952 (N_2952,N_2629,N_2668);
and U2953 (N_2953,N_2636,N_2676);
nor U2954 (N_2954,N_2527,N_2573);
xor U2955 (N_2955,N_2525,N_2748);
xor U2956 (N_2956,N_2630,N_2593);
and U2957 (N_2957,N_2548,N_2545);
xnor U2958 (N_2958,N_2617,N_2661);
and U2959 (N_2959,N_2706,N_2720);
and U2960 (N_2960,N_2741,N_2637);
and U2961 (N_2961,N_2592,N_2710);
and U2962 (N_2962,N_2710,N_2707);
nand U2963 (N_2963,N_2546,N_2730);
nand U2964 (N_2964,N_2652,N_2615);
and U2965 (N_2965,N_2616,N_2686);
xnor U2966 (N_2966,N_2712,N_2701);
nand U2967 (N_2967,N_2653,N_2505);
xnor U2968 (N_2968,N_2560,N_2543);
xnor U2969 (N_2969,N_2539,N_2643);
and U2970 (N_2970,N_2737,N_2643);
nand U2971 (N_2971,N_2706,N_2656);
nor U2972 (N_2972,N_2703,N_2745);
or U2973 (N_2973,N_2638,N_2564);
or U2974 (N_2974,N_2564,N_2525);
nand U2975 (N_2975,N_2567,N_2517);
nor U2976 (N_2976,N_2686,N_2540);
and U2977 (N_2977,N_2711,N_2703);
xnor U2978 (N_2978,N_2598,N_2726);
nor U2979 (N_2979,N_2665,N_2550);
and U2980 (N_2980,N_2552,N_2555);
and U2981 (N_2981,N_2538,N_2705);
xnor U2982 (N_2982,N_2711,N_2552);
xnor U2983 (N_2983,N_2647,N_2645);
nand U2984 (N_2984,N_2628,N_2621);
and U2985 (N_2985,N_2547,N_2747);
nor U2986 (N_2986,N_2589,N_2535);
and U2987 (N_2987,N_2684,N_2713);
xnor U2988 (N_2988,N_2659,N_2583);
xor U2989 (N_2989,N_2600,N_2576);
nor U2990 (N_2990,N_2528,N_2525);
nor U2991 (N_2991,N_2700,N_2603);
xnor U2992 (N_2992,N_2554,N_2689);
xnor U2993 (N_2993,N_2613,N_2536);
nor U2994 (N_2994,N_2596,N_2653);
xor U2995 (N_2995,N_2722,N_2584);
and U2996 (N_2996,N_2680,N_2596);
xor U2997 (N_2997,N_2532,N_2522);
xor U2998 (N_2998,N_2587,N_2663);
xnor U2999 (N_2999,N_2720,N_2636);
nand U3000 (N_3000,N_2991,N_2973);
and U3001 (N_3001,N_2768,N_2901);
xnor U3002 (N_3002,N_2845,N_2877);
or U3003 (N_3003,N_2856,N_2880);
or U3004 (N_3004,N_2859,N_2970);
and U3005 (N_3005,N_2923,N_2964);
and U3006 (N_3006,N_2808,N_2751);
or U3007 (N_3007,N_2777,N_2934);
and U3008 (N_3008,N_2852,N_2779);
xnor U3009 (N_3009,N_2840,N_2847);
or U3010 (N_3010,N_2885,N_2913);
nand U3011 (N_3011,N_2952,N_2818);
nor U3012 (N_3012,N_2884,N_2920);
nand U3013 (N_3013,N_2906,N_2869);
xnor U3014 (N_3014,N_2796,N_2989);
and U3015 (N_3015,N_2902,N_2876);
nand U3016 (N_3016,N_2921,N_2870);
xor U3017 (N_3017,N_2947,N_2780);
or U3018 (N_3018,N_2760,N_2834);
nand U3019 (N_3019,N_2763,N_2863);
nand U3020 (N_3020,N_2810,N_2839);
nand U3021 (N_3021,N_2850,N_2937);
nand U3022 (N_3022,N_2925,N_2787);
xnor U3023 (N_3023,N_2953,N_2995);
or U3024 (N_3024,N_2811,N_2844);
nand U3025 (N_3025,N_2871,N_2967);
nor U3026 (N_3026,N_2762,N_2754);
xor U3027 (N_3027,N_2927,N_2928);
nand U3028 (N_3028,N_2832,N_2959);
or U3029 (N_3029,N_2978,N_2764);
xnor U3030 (N_3030,N_2949,N_2875);
nand U3031 (N_3031,N_2817,N_2756);
and U3032 (N_3032,N_2940,N_2790);
nand U3033 (N_3033,N_2893,N_2954);
or U3034 (N_3034,N_2882,N_2969);
nor U3035 (N_3035,N_2938,N_2957);
or U3036 (N_3036,N_2807,N_2828);
nand U3037 (N_3037,N_2912,N_2892);
xor U3038 (N_3038,N_2766,N_2750);
nor U3039 (N_3039,N_2799,N_2965);
xnor U3040 (N_3040,N_2917,N_2890);
nand U3041 (N_3041,N_2771,N_2908);
nor U3042 (N_3042,N_2905,N_2857);
and U3043 (N_3043,N_2775,N_2803);
and U3044 (N_3044,N_2948,N_2895);
nand U3045 (N_3045,N_2753,N_2886);
xor U3046 (N_3046,N_2889,N_2776);
or U3047 (N_3047,N_2769,N_2897);
nor U3048 (N_3048,N_2974,N_2891);
nor U3049 (N_3049,N_2958,N_2909);
and U3050 (N_3050,N_2931,N_2757);
nand U3051 (N_3051,N_2843,N_2903);
nor U3052 (N_3052,N_2961,N_2819);
or U3053 (N_3053,N_2981,N_2907);
and U3054 (N_3054,N_2977,N_2822);
nand U3055 (N_3055,N_2836,N_2941);
and U3056 (N_3056,N_2944,N_2888);
nor U3057 (N_3057,N_2783,N_2820);
or U3058 (N_3058,N_2951,N_2855);
and U3059 (N_3059,N_2914,N_2994);
nor U3060 (N_3060,N_2900,N_2926);
xnor U3061 (N_3061,N_2813,N_2976);
and U3062 (N_3062,N_2831,N_2864);
nand U3063 (N_3063,N_2792,N_2963);
or U3064 (N_3064,N_2781,N_2975);
nor U3065 (N_3065,N_2804,N_2998);
xnor U3066 (N_3066,N_2767,N_2791);
nand U3067 (N_3067,N_2881,N_2933);
nor U3068 (N_3068,N_2761,N_2812);
or U3069 (N_3069,N_2786,N_2825);
or U3070 (N_3070,N_2835,N_2930);
or U3071 (N_3071,N_2867,N_2830);
nand U3072 (N_3072,N_2833,N_2824);
nor U3073 (N_3073,N_2814,N_2983);
xnor U3074 (N_3074,N_2988,N_2996);
nor U3075 (N_3075,N_2883,N_2943);
nor U3076 (N_3076,N_2910,N_2987);
xnor U3077 (N_3077,N_2922,N_2801);
xor U3078 (N_3078,N_2955,N_2800);
or U3079 (N_3079,N_2924,N_2849);
nor U3080 (N_3080,N_2966,N_2915);
or U3081 (N_3081,N_2872,N_2874);
xnor U3082 (N_3082,N_2999,N_2815);
and U3083 (N_3083,N_2848,N_2782);
and U3084 (N_3084,N_2778,N_2950);
and U3085 (N_3085,N_2837,N_2789);
or U3086 (N_3086,N_2853,N_2990);
xnor U3087 (N_3087,N_2968,N_2841);
xnor U3088 (N_3088,N_2794,N_2972);
xnor U3089 (N_3089,N_2854,N_2752);
or U3090 (N_3090,N_2755,N_2993);
nor U3091 (N_3091,N_2873,N_2986);
nand U3092 (N_3092,N_2896,N_2851);
nand U3093 (N_3093,N_2919,N_2971);
xnor U3094 (N_3094,N_2798,N_2758);
nor U3095 (N_3095,N_2860,N_2946);
nor U3096 (N_3096,N_2936,N_2774);
xnor U3097 (N_3097,N_2868,N_2985);
nor U3098 (N_3098,N_2862,N_2979);
nor U3099 (N_3099,N_2911,N_2838);
and U3100 (N_3100,N_2899,N_2929);
nand U3101 (N_3101,N_2802,N_2945);
and U3102 (N_3102,N_2894,N_2797);
nor U3103 (N_3103,N_2829,N_2942);
nor U3104 (N_3104,N_2878,N_2984);
or U3105 (N_3105,N_2770,N_2784);
nor U3106 (N_3106,N_2997,N_2865);
xor U3107 (N_3107,N_2918,N_2826);
nand U3108 (N_3108,N_2935,N_2805);
nand U3109 (N_3109,N_2904,N_2898);
nand U3110 (N_3110,N_2821,N_2887);
and U3111 (N_3111,N_2956,N_2772);
nor U3112 (N_3112,N_2879,N_2759);
or U3113 (N_3113,N_2861,N_2960);
and U3114 (N_3114,N_2992,N_2816);
xor U3115 (N_3115,N_2793,N_2765);
nand U3116 (N_3116,N_2962,N_2939);
or U3117 (N_3117,N_2866,N_2858);
or U3118 (N_3118,N_2788,N_2795);
xnor U3119 (N_3119,N_2773,N_2982);
xor U3120 (N_3120,N_2827,N_2809);
xor U3121 (N_3121,N_2932,N_2980);
nand U3122 (N_3122,N_2823,N_2842);
nand U3123 (N_3123,N_2916,N_2785);
nor U3124 (N_3124,N_2846,N_2806);
or U3125 (N_3125,N_2970,N_2816);
nor U3126 (N_3126,N_2839,N_2911);
nand U3127 (N_3127,N_2848,N_2905);
nand U3128 (N_3128,N_2938,N_2995);
nand U3129 (N_3129,N_2862,N_2792);
and U3130 (N_3130,N_2778,N_2999);
xnor U3131 (N_3131,N_2981,N_2924);
and U3132 (N_3132,N_2776,N_2778);
xor U3133 (N_3133,N_2859,N_2880);
xor U3134 (N_3134,N_2885,N_2763);
nor U3135 (N_3135,N_2818,N_2959);
and U3136 (N_3136,N_2901,N_2915);
nand U3137 (N_3137,N_2848,N_2847);
nor U3138 (N_3138,N_2964,N_2842);
xnor U3139 (N_3139,N_2863,N_2810);
nor U3140 (N_3140,N_2950,N_2838);
nand U3141 (N_3141,N_2853,N_2863);
nand U3142 (N_3142,N_2944,N_2927);
and U3143 (N_3143,N_2858,N_2901);
or U3144 (N_3144,N_2992,N_2942);
and U3145 (N_3145,N_2921,N_2843);
xor U3146 (N_3146,N_2974,N_2949);
nor U3147 (N_3147,N_2889,N_2830);
and U3148 (N_3148,N_2891,N_2900);
nor U3149 (N_3149,N_2779,N_2885);
and U3150 (N_3150,N_2968,N_2824);
and U3151 (N_3151,N_2913,N_2846);
xnor U3152 (N_3152,N_2945,N_2851);
or U3153 (N_3153,N_2792,N_2763);
or U3154 (N_3154,N_2808,N_2846);
nand U3155 (N_3155,N_2786,N_2956);
nand U3156 (N_3156,N_2773,N_2881);
or U3157 (N_3157,N_2909,N_2918);
nand U3158 (N_3158,N_2874,N_2873);
nor U3159 (N_3159,N_2778,N_2869);
and U3160 (N_3160,N_2842,N_2932);
and U3161 (N_3161,N_2868,N_2776);
and U3162 (N_3162,N_2799,N_2769);
or U3163 (N_3163,N_2955,N_2916);
nor U3164 (N_3164,N_2773,N_2936);
xor U3165 (N_3165,N_2884,N_2839);
nand U3166 (N_3166,N_2785,N_2943);
nor U3167 (N_3167,N_2814,N_2923);
xor U3168 (N_3168,N_2750,N_2922);
xor U3169 (N_3169,N_2968,N_2934);
xor U3170 (N_3170,N_2991,N_2938);
or U3171 (N_3171,N_2819,N_2890);
or U3172 (N_3172,N_2891,N_2844);
nor U3173 (N_3173,N_2913,N_2784);
nand U3174 (N_3174,N_2779,N_2830);
nand U3175 (N_3175,N_2855,N_2969);
or U3176 (N_3176,N_2815,N_2798);
nand U3177 (N_3177,N_2942,N_2995);
nand U3178 (N_3178,N_2784,N_2924);
nand U3179 (N_3179,N_2850,N_2915);
xor U3180 (N_3180,N_2809,N_2799);
and U3181 (N_3181,N_2965,N_2918);
and U3182 (N_3182,N_2920,N_2867);
nor U3183 (N_3183,N_2982,N_2751);
and U3184 (N_3184,N_2907,N_2942);
or U3185 (N_3185,N_2969,N_2891);
and U3186 (N_3186,N_2874,N_2941);
xnor U3187 (N_3187,N_2844,N_2810);
nand U3188 (N_3188,N_2972,N_2801);
or U3189 (N_3189,N_2761,N_2947);
nor U3190 (N_3190,N_2939,N_2752);
nand U3191 (N_3191,N_2918,N_2892);
nor U3192 (N_3192,N_2777,N_2769);
or U3193 (N_3193,N_2958,N_2974);
and U3194 (N_3194,N_2987,N_2936);
xor U3195 (N_3195,N_2985,N_2892);
xor U3196 (N_3196,N_2948,N_2993);
xor U3197 (N_3197,N_2962,N_2981);
nand U3198 (N_3198,N_2925,N_2868);
nand U3199 (N_3199,N_2756,N_2761);
xor U3200 (N_3200,N_2938,N_2912);
and U3201 (N_3201,N_2959,N_2821);
and U3202 (N_3202,N_2872,N_2824);
nand U3203 (N_3203,N_2827,N_2931);
nor U3204 (N_3204,N_2765,N_2974);
and U3205 (N_3205,N_2870,N_2885);
nor U3206 (N_3206,N_2929,N_2836);
nand U3207 (N_3207,N_2846,N_2915);
nand U3208 (N_3208,N_2805,N_2919);
nor U3209 (N_3209,N_2854,N_2883);
or U3210 (N_3210,N_2871,N_2768);
or U3211 (N_3211,N_2865,N_2853);
nand U3212 (N_3212,N_2780,N_2826);
nand U3213 (N_3213,N_2934,N_2885);
nor U3214 (N_3214,N_2930,N_2983);
or U3215 (N_3215,N_2963,N_2885);
nand U3216 (N_3216,N_2952,N_2957);
or U3217 (N_3217,N_2778,N_2834);
or U3218 (N_3218,N_2926,N_2819);
nand U3219 (N_3219,N_2973,N_2790);
xor U3220 (N_3220,N_2802,N_2848);
xor U3221 (N_3221,N_2922,N_2897);
or U3222 (N_3222,N_2948,N_2921);
and U3223 (N_3223,N_2981,N_2861);
xor U3224 (N_3224,N_2814,N_2960);
and U3225 (N_3225,N_2772,N_2771);
and U3226 (N_3226,N_2989,N_2996);
xnor U3227 (N_3227,N_2772,N_2796);
and U3228 (N_3228,N_2933,N_2854);
or U3229 (N_3229,N_2972,N_2858);
nor U3230 (N_3230,N_2758,N_2991);
nor U3231 (N_3231,N_2912,N_2813);
and U3232 (N_3232,N_2989,N_2925);
xnor U3233 (N_3233,N_2845,N_2879);
xor U3234 (N_3234,N_2839,N_2946);
nor U3235 (N_3235,N_2986,N_2964);
and U3236 (N_3236,N_2873,N_2802);
xor U3237 (N_3237,N_2760,N_2853);
xnor U3238 (N_3238,N_2941,N_2829);
and U3239 (N_3239,N_2995,N_2977);
nand U3240 (N_3240,N_2821,N_2878);
xnor U3241 (N_3241,N_2930,N_2912);
and U3242 (N_3242,N_2950,N_2817);
nand U3243 (N_3243,N_2891,N_2836);
or U3244 (N_3244,N_2951,N_2772);
and U3245 (N_3245,N_2782,N_2825);
xnor U3246 (N_3246,N_2976,N_2871);
xnor U3247 (N_3247,N_2824,N_2773);
xnor U3248 (N_3248,N_2890,N_2770);
nand U3249 (N_3249,N_2832,N_2987);
nor U3250 (N_3250,N_3193,N_3145);
nand U3251 (N_3251,N_3001,N_3026);
or U3252 (N_3252,N_3228,N_3128);
and U3253 (N_3253,N_3165,N_3035);
xor U3254 (N_3254,N_3086,N_3152);
or U3255 (N_3255,N_3096,N_3091);
and U3256 (N_3256,N_3075,N_3117);
or U3257 (N_3257,N_3019,N_3221);
nand U3258 (N_3258,N_3194,N_3039);
nor U3259 (N_3259,N_3083,N_3003);
nor U3260 (N_3260,N_3072,N_3048);
and U3261 (N_3261,N_3240,N_3089);
xor U3262 (N_3262,N_3130,N_3110);
nand U3263 (N_3263,N_3006,N_3051);
nor U3264 (N_3264,N_3021,N_3212);
xnor U3265 (N_3265,N_3232,N_3078);
or U3266 (N_3266,N_3027,N_3069);
nand U3267 (N_3267,N_3201,N_3202);
xnor U3268 (N_3268,N_3023,N_3033);
nor U3269 (N_3269,N_3198,N_3104);
and U3270 (N_3270,N_3149,N_3060);
nor U3271 (N_3271,N_3045,N_3199);
or U3272 (N_3272,N_3044,N_3239);
nand U3273 (N_3273,N_3184,N_3182);
nand U3274 (N_3274,N_3205,N_3178);
and U3275 (N_3275,N_3009,N_3008);
or U3276 (N_3276,N_3237,N_3061);
nand U3277 (N_3277,N_3057,N_3148);
xnor U3278 (N_3278,N_3140,N_3097);
or U3279 (N_3279,N_3190,N_3047);
nand U3280 (N_3280,N_3064,N_3220);
nor U3281 (N_3281,N_3192,N_3231);
nor U3282 (N_3282,N_3093,N_3055);
or U3283 (N_3283,N_3107,N_3095);
nor U3284 (N_3284,N_3007,N_3123);
and U3285 (N_3285,N_3084,N_3063);
and U3286 (N_3286,N_3210,N_3041);
nor U3287 (N_3287,N_3109,N_3218);
nor U3288 (N_3288,N_3187,N_3214);
nor U3289 (N_3289,N_3243,N_3090);
xnor U3290 (N_3290,N_3206,N_3166);
nand U3291 (N_3291,N_3038,N_3070);
and U3292 (N_3292,N_3151,N_3010);
nand U3293 (N_3293,N_3219,N_3098);
nand U3294 (N_3294,N_3147,N_3106);
and U3295 (N_3295,N_3118,N_3241);
or U3296 (N_3296,N_3032,N_3042);
xor U3297 (N_3297,N_3211,N_3004);
or U3298 (N_3298,N_3233,N_3196);
and U3299 (N_3299,N_3142,N_3133);
nand U3300 (N_3300,N_3122,N_3170);
or U3301 (N_3301,N_3203,N_3216);
nand U3302 (N_3302,N_3005,N_3013);
xnor U3303 (N_3303,N_3222,N_3082);
xor U3304 (N_3304,N_3167,N_3209);
nor U3305 (N_3305,N_3085,N_3120);
or U3306 (N_3306,N_3238,N_3073);
or U3307 (N_3307,N_3100,N_3080);
xor U3308 (N_3308,N_3015,N_3011);
and U3309 (N_3309,N_3012,N_3054);
xnor U3310 (N_3310,N_3188,N_3144);
and U3311 (N_3311,N_3087,N_3103);
or U3312 (N_3312,N_3179,N_3177);
xnor U3313 (N_3313,N_3146,N_3230);
nand U3314 (N_3314,N_3245,N_3105);
or U3315 (N_3315,N_3043,N_3094);
or U3316 (N_3316,N_3071,N_3134);
xnor U3317 (N_3317,N_3036,N_3161);
nand U3318 (N_3318,N_3226,N_3129);
nand U3319 (N_3319,N_3236,N_3079);
nand U3320 (N_3320,N_3197,N_3076);
or U3321 (N_3321,N_3074,N_3116);
xnor U3322 (N_3322,N_3156,N_3217);
nand U3323 (N_3323,N_3126,N_3248);
nand U3324 (N_3324,N_3066,N_3050);
or U3325 (N_3325,N_3017,N_3135);
or U3326 (N_3326,N_3227,N_3185);
nor U3327 (N_3327,N_3139,N_3059);
or U3328 (N_3328,N_3025,N_3138);
nor U3329 (N_3329,N_3159,N_3030);
nand U3330 (N_3330,N_3157,N_3215);
xnor U3331 (N_3331,N_3204,N_3127);
and U3332 (N_3332,N_3173,N_3121);
or U3333 (N_3333,N_3154,N_3213);
or U3334 (N_3334,N_3189,N_3223);
xnor U3335 (N_3335,N_3065,N_3029);
and U3336 (N_3336,N_3153,N_3132);
nand U3337 (N_3337,N_3014,N_3141);
nor U3338 (N_3338,N_3099,N_3175);
nor U3339 (N_3339,N_3163,N_3031);
nor U3340 (N_3340,N_3229,N_3249);
nand U3341 (N_3341,N_3235,N_3191);
and U3342 (N_3342,N_3053,N_3049);
xnor U3343 (N_3343,N_3125,N_3046);
nor U3344 (N_3344,N_3037,N_3234);
or U3345 (N_3345,N_3242,N_3018);
nor U3346 (N_3346,N_3244,N_3186);
nand U3347 (N_3347,N_3195,N_3062);
nor U3348 (N_3348,N_3158,N_3208);
and U3349 (N_3349,N_3034,N_3247);
nand U3350 (N_3350,N_3040,N_3168);
and U3351 (N_3351,N_3174,N_3067);
and U3352 (N_3352,N_3000,N_3155);
or U3353 (N_3353,N_3052,N_3246);
nor U3354 (N_3354,N_3150,N_3024);
or U3355 (N_3355,N_3160,N_3111);
or U3356 (N_3356,N_3002,N_3020);
nor U3357 (N_3357,N_3183,N_3102);
xor U3358 (N_3358,N_3124,N_3114);
or U3359 (N_3359,N_3028,N_3143);
and U3360 (N_3360,N_3169,N_3131);
nor U3361 (N_3361,N_3077,N_3176);
and U3362 (N_3362,N_3164,N_3171);
nand U3363 (N_3363,N_3113,N_3181);
xor U3364 (N_3364,N_3115,N_3022);
and U3365 (N_3365,N_3172,N_3101);
or U3366 (N_3366,N_3180,N_3081);
and U3367 (N_3367,N_3092,N_3162);
nor U3368 (N_3368,N_3088,N_3136);
nor U3369 (N_3369,N_3207,N_3056);
or U3370 (N_3370,N_3058,N_3225);
xor U3371 (N_3371,N_3068,N_3224);
and U3372 (N_3372,N_3112,N_3200);
or U3373 (N_3373,N_3119,N_3016);
nand U3374 (N_3374,N_3108,N_3137);
nand U3375 (N_3375,N_3172,N_3063);
nand U3376 (N_3376,N_3215,N_3219);
nand U3377 (N_3377,N_3098,N_3106);
xnor U3378 (N_3378,N_3008,N_3026);
or U3379 (N_3379,N_3138,N_3043);
xnor U3380 (N_3380,N_3189,N_3236);
nor U3381 (N_3381,N_3000,N_3223);
or U3382 (N_3382,N_3187,N_3028);
nand U3383 (N_3383,N_3190,N_3158);
or U3384 (N_3384,N_3226,N_3141);
nor U3385 (N_3385,N_3083,N_3244);
and U3386 (N_3386,N_3053,N_3121);
nand U3387 (N_3387,N_3077,N_3025);
xnor U3388 (N_3388,N_3092,N_3034);
nor U3389 (N_3389,N_3217,N_3092);
xor U3390 (N_3390,N_3035,N_3249);
and U3391 (N_3391,N_3154,N_3125);
and U3392 (N_3392,N_3225,N_3147);
or U3393 (N_3393,N_3039,N_3051);
and U3394 (N_3394,N_3228,N_3065);
nand U3395 (N_3395,N_3092,N_3104);
xnor U3396 (N_3396,N_3225,N_3172);
and U3397 (N_3397,N_3192,N_3244);
nand U3398 (N_3398,N_3108,N_3213);
and U3399 (N_3399,N_3017,N_3114);
or U3400 (N_3400,N_3006,N_3089);
xor U3401 (N_3401,N_3001,N_3138);
nand U3402 (N_3402,N_3102,N_3239);
nand U3403 (N_3403,N_3002,N_3094);
and U3404 (N_3404,N_3020,N_3142);
nor U3405 (N_3405,N_3083,N_3095);
and U3406 (N_3406,N_3107,N_3048);
or U3407 (N_3407,N_3232,N_3100);
nand U3408 (N_3408,N_3021,N_3191);
xor U3409 (N_3409,N_3230,N_3083);
nand U3410 (N_3410,N_3186,N_3171);
nand U3411 (N_3411,N_3100,N_3083);
or U3412 (N_3412,N_3069,N_3228);
and U3413 (N_3413,N_3029,N_3172);
xnor U3414 (N_3414,N_3061,N_3062);
or U3415 (N_3415,N_3150,N_3199);
nand U3416 (N_3416,N_3031,N_3069);
xor U3417 (N_3417,N_3126,N_3107);
xor U3418 (N_3418,N_3052,N_3223);
xor U3419 (N_3419,N_3107,N_3207);
nor U3420 (N_3420,N_3048,N_3227);
and U3421 (N_3421,N_3012,N_3067);
or U3422 (N_3422,N_3041,N_3035);
nor U3423 (N_3423,N_3141,N_3206);
or U3424 (N_3424,N_3000,N_3110);
nand U3425 (N_3425,N_3102,N_3113);
nand U3426 (N_3426,N_3246,N_3146);
nor U3427 (N_3427,N_3112,N_3053);
and U3428 (N_3428,N_3189,N_3042);
xor U3429 (N_3429,N_3192,N_3039);
nor U3430 (N_3430,N_3103,N_3024);
and U3431 (N_3431,N_3104,N_3143);
and U3432 (N_3432,N_3009,N_3102);
nand U3433 (N_3433,N_3240,N_3105);
xnor U3434 (N_3434,N_3174,N_3106);
nand U3435 (N_3435,N_3012,N_3058);
or U3436 (N_3436,N_3084,N_3167);
nand U3437 (N_3437,N_3101,N_3086);
nor U3438 (N_3438,N_3246,N_3230);
and U3439 (N_3439,N_3014,N_3032);
nor U3440 (N_3440,N_3240,N_3106);
nand U3441 (N_3441,N_3071,N_3137);
xor U3442 (N_3442,N_3041,N_3135);
nand U3443 (N_3443,N_3170,N_3193);
nor U3444 (N_3444,N_3148,N_3074);
nand U3445 (N_3445,N_3215,N_3172);
or U3446 (N_3446,N_3170,N_3188);
nor U3447 (N_3447,N_3154,N_3031);
and U3448 (N_3448,N_3123,N_3068);
or U3449 (N_3449,N_3095,N_3194);
nand U3450 (N_3450,N_3178,N_3156);
or U3451 (N_3451,N_3247,N_3232);
nand U3452 (N_3452,N_3011,N_3177);
or U3453 (N_3453,N_3010,N_3139);
and U3454 (N_3454,N_3187,N_3064);
nor U3455 (N_3455,N_3149,N_3187);
xnor U3456 (N_3456,N_3094,N_3197);
and U3457 (N_3457,N_3190,N_3156);
nand U3458 (N_3458,N_3182,N_3045);
xor U3459 (N_3459,N_3037,N_3170);
nand U3460 (N_3460,N_3208,N_3201);
xor U3461 (N_3461,N_3052,N_3168);
nor U3462 (N_3462,N_3036,N_3071);
and U3463 (N_3463,N_3202,N_3056);
or U3464 (N_3464,N_3078,N_3238);
nand U3465 (N_3465,N_3019,N_3116);
xnor U3466 (N_3466,N_3237,N_3180);
and U3467 (N_3467,N_3089,N_3148);
nor U3468 (N_3468,N_3084,N_3222);
xnor U3469 (N_3469,N_3080,N_3127);
nand U3470 (N_3470,N_3046,N_3236);
nor U3471 (N_3471,N_3128,N_3222);
nor U3472 (N_3472,N_3007,N_3087);
nand U3473 (N_3473,N_3113,N_3093);
nand U3474 (N_3474,N_3006,N_3023);
or U3475 (N_3475,N_3233,N_3068);
nor U3476 (N_3476,N_3216,N_3145);
nand U3477 (N_3477,N_3094,N_3072);
and U3478 (N_3478,N_3016,N_3214);
xor U3479 (N_3479,N_3128,N_3156);
nor U3480 (N_3480,N_3025,N_3067);
or U3481 (N_3481,N_3204,N_3212);
or U3482 (N_3482,N_3025,N_3068);
or U3483 (N_3483,N_3159,N_3147);
nand U3484 (N_3484,N_3098,N_3099);
xnor U3485 (N_3485,N_3011,N_3076);
and U3486 (N_3486,N_3148,N_3180);
nand U3487 (N_3487,N_3096,N_3070);
nor U3488 (N_3488,N_3160,N_3110);
and U3489 (N_3489,N_3057,N_3227);
or U3490 (N_3490,N_3190,N_3143);
and U3491 (N_3491,N_3239,N_3117);
nand U3492 (N_3492,N_3064,N_3133);
or U3493 (N_3493,N_3129,N_3115);
nor U3494 (N_3494,N_3085,N_3103);
nor U3495 (N_3495,N_3024,N_3048);
and U3496 (N_3496,N_3062,N_3105);
nand U3497 (N_3497,N_3051,N_3001);
and U3498 (N_3498,N_3149,N_3042);
nand U3499 (N_3499,N_3133,N_3001);
nor U3500 (N_3500,N_3281,N_3336);
xor U3501 (N_3501,N_3371,N_3490);
nor U3502 (N_3502,N_3301,N_3308);
xnor U3503 (N_3503,N_3359,N_3404);
nand U3504 (N_3504,N_3448,N_3346);
or U3505 (N_3505,N_3487,N_3278);
nor U3506 (N_3506,N_3435,N_3398);
xnor U3507 (N_3507,N_3458,N_3498);
nor U3508 (N_3508,N_3262,N_3275);
nor U3509 (N_3509,N_3377,N_3461);
xor U3510 (N_3510,N_3290,N_3323);
or U3511 (N_3511,N_3470,N_3297);
and U3512 (N_3512,N_3303,N_3492);
xnor U3513 (N_3513,N_3347,N_3272);
nor U3514 (N_3514,N_3373,N_3311);
or U3515 (N_3515,N_3376,N_3496);
nor U3516 (N_3516,N_3357,N_3427);
xor U3517 (N_3517,N_3274,N_3318);
xnor U3518 (N_3518,N_3326,N_3285);
nand U3519 (N_3519,N_3405,N_3356);
or U3520 (N_3520,N_3329,N_3399);
nand U3521 (N_3521,N_3423,N_3299);
xor U3522 (N_3522,N_3322,N_3302);
xnor U3523 (N_3523,N_3429,N_3372);
nor U3524 (N_3524,N_3387,N_3374);
and U3525 (N_3525,N_3462,N_3413);
xor U3526 (N_3526,N_3460,N_3366);
or U3527 (N_3527,N_3397,N_3294);
or U3528 (N_3528,N_3390,N_3475);
nand U3529 (N_3529,N_3471,N_3402);
and U3530 (N_3530,N_3345,N_3416);
xnor U3531 (N_3531,N_3447,N_3330);
or U3532 (N_3532,N_3419,N_3282);
and U3533 (N_3533,N_3408,N_3289);
and U3534 (N_3534,N_3436,N_3484);
or U3535 (N_3535,N_3383,N_3327);
nor U3536 (N_3536,N_3361,N_3332);
and U3537 (N_3537,N_3328,N_3381);
or U3538 (N_3538,N_3307,N_3375);
nand U3539 (N_3539,N_3368,N_3292);
xor U3540 (N_3540,N_3263,N_3250);
and U3541 (N_3541,N_3493,N_3384);
and U3542 (N_3542,N_3264,N_3414);
nor U3543 (N_3543,N_3352,N_3320);
nand U3544 (N_3544,N_3449,N_3273);
and U3545 (N_3545,N_3364,N_3442);
or U3546 (N_3546,N_3425,N_3454);
and U3547 (N_3547,N_3463,N_3338);
nor U3548 (N_3548,N_3270,N_3488);
xor U3549 (N_3549,N_3392,N_3296);
nand U3550 (N_3550,N_3256,N_3465);
xnor U3551 (N_3551,N_3450,N_3410);
nand U3552 (N_3552,N_3446,N_3421);
xor U3553 (N_3553,N_3431,N_3315);
or U3554 (N_3554,N_3258,N_3255);
or U3555 (N_3555,N_3483,N_3276);
nor U3556 (N_3556,N_3474,N_3467);
xnor U3557 (N_3557,N_3389,N_3426);
nand U3558 (N_3558,N_3331,N_3340);
xor U3559 (N_3559,N_3486,N_3300);
or U3560 (N_3560,N_3485,N_3464);
nor U3561 (N_3561,N_3266,N_3333);
nor U3562 (N_3562,N_3451,N_3499);
or U3563 (N_3563,N_3260,N_3388);
nor U3564 (N_3564,N_3283,N_3469);
or U3565 (N_3565,N_3358,N_3444);
or U3566 (N_3566,N_3351,N_3253);
nor U3567 (N_3567,N_3453,N_3418);
and U3568 (N_3568,N_3481,N_3365);
xnor U3569 (N_3569,N_3355,N_3482);
nor U3570 (N_3570,N_3288,N_3433);
nand U3571 (N_3571,N_3417,N_3494);
and U3572 (N_3572,N_3324,N_3312);
nand U3573 (N_3573,N_3265,N_3295);
or U3574 (N_3574,N_3452,N_3400);
nand U3575 (N_3575,N_3251,N_3316);
nor U3576 (N_3576,N_3268,N_3439);
xnor U3577 (N_3577,N_3489,N_3385);
nor U3578 (N_3578,N_3386,N_3434);
nor U3579 (N_3579,N_3319,N_3370);
and U3580 (N_3580,N_3280,N_3252);
nand U3581 (N_3581,N_3286,N_3348);
or U3582 (N_3582,N_3437,N_3304);
xor U3583 (N_3583,N_3382,N_3342);
or U3584 (N_3584,N_3363,N_3335);
or U3585 (N_3585,N_3362,N_3394);
or U3586 (N_3586,N_3473,N_3456);
nand U3587 (N_3587,N_3380,N_3468);
nand U3588 (N_3588,N_3305,N_3267);
nor U3589 (N_3589,N_3350,N_3424);
and U3590 (N_3590,N_3438,N_3271);
or U3591 (N_3591,N_3334,N_3480);
xnor U3592 (N_3592,N_3401,N_3349);
and U3593 (N_3593,N_3430,N_3309);
nand U3594 (N_3594,N_3459,N_3395);
nor U3595 (N_3595,N_3441,N_3353);
xnor U3596 (N_3596,N_3379,N_3497);
nor U3597 (N_3597,N_3337,N_3495);
nor U3598 (N_3598,N_3317,N_3391);
xnor U3599 (N_3599,N_3310,N_3306);
or U3600 (N_3600,N_3440,N_3321);
nand U3601 (N_3601,N_3443,N_3412);
nor U3602 (N_3602,N_3339,N_3254);
and U3603 (N_3603,N_3277,N_3279);
nand U3604 (N_3604,N_3325,N_3466);
xnor U3605 (N_3605,N_3341,N_3455);
nand U3606 (N_3606,N_3396,N_3284);
and U3607 (N_3607,N_3428,N_3313);
nand U3608 (N_3608,N_3409,N_3360);
xnor U3609 (N_3609,N_3476,N_3407);
and U3610 (N_3610,N_3422,N_3367);
and U3611 (N_3611,N_3472,N_3393);
or U3612 (N_3612,N_3287,N_3261);
and U3613 (N_3613,N_3344,N_3491);
nor U3614 (N_3614,N_3411,N_3259);
nand U3615 (N_3615,N_3457,N_3445);
xnor U3616 (N_3616,N_3369,N_3314);
xor U3617 (N_3617,N_3415,N_3298);
or U3618 (N_3618,N_3420,N_3257);
or U3619 (N_3619,N_3269,N_3378);
nor U3620 (N_3620,N_3478,N_3354);
xnor U3621 (N_3621,N_3403,N_3343);
nand U3622 (N_3622,N_3479,N_3477);
nand U3623 (N_3623,N_3406,N_3293);
nor U3624 (N_3624,N_3432,N_3291);
nor U3625 (N_3625,N_3386,N_3273);
nand U3626 (N_3626,N_3374,N_3470);
or U3627 (N_3627,N_3457,N_3446);
xor U3628 (N_3628,N_3471,N_3419);
or U3629 (N_3629,N_3401,N_3373);
and U3630 (N_3630,N_3426,N_3478);
or U3631 (N_3631,N_3462,N_3420);
or U3632 (N_3632,N_3458,N_3456);
xnor U3633 (N_3633,N_3393,N_3394);
nand U3634 (N_3634,N_3468,N_3323);
nor U3635 (N_3635,N_3342,N_3353);
nand U3636 (N_3636,N_3361,N_3260);
nor U3637 (N_3637,N_3430,N_3496);
and U3638 (N_3638,N_3449,N_3343);
nand U3639 (N_3639,N_3354,N_3276);
nand U3640 (N_3640,N_3342,N_3488);
xor U3641 (N_3641,N_3333,N_3429);
and U3642 (N_3642,N_3419,N_3414);
and U3643 (N_3643,N_3335,N_3387);
xor U3644 (N_3644,N_3278,N_3296);
and U3645 (N_3645,N_3349,N_3441);
nor U3646 (N_3646,N_3325,N_3484);
or U3647 (N_3647,N_3292,N_3254);
and U3648 (N_3648,N_3444,N_3279);
and U3649 (N_3649,N_3496,N_3490);
nor U3650 (N_3650,N_3411,N_3475);
nor U3651 (N_3651,N_3434,N_3499);
nor U3652 (N_3652,N_3343,N_3398);
or U3653 (N_3653,N_3355,N_3284);
nand U3654 (N_3654,N_3433,N_3477);
nand U3655 (N_3655,N_3366,N_3335);
or U3656 (N_3656,N_3262,N_3252);
xnor U3657 (N_3657,N_3297,N_3435);
or U3658 (N_3658,N_3466,N_3301);
and U3659 (N_3659,N_3468,N_3499);
or U3660 (N_3660,N_3474,N_3290);
nor U3661 (N_3661,N_3474,N_3420);
nand U3662 (N_3662,N_3254,N_3393);
xor U3663 (N_3663,N_3301,N_3385);
xnor U3664 (N_3664,N_3460,N_3259);
or U3665 (N_3665,N_3364,N_3283);
xor U3666 (N_3666,N_3464,N_3398);
and U3667 (N_3667,N_3376,N_3440);
nand U3668 (N_3668,N_3472,N_3462);
xnor U3669 (N_3669,N_3491,N_3416);
nor U3670 (N_3670,N_3394,N_3443);
and U3671 (N_3671,N_3412,N_3464);
nand U3672 (N_3672,N_3408,N_3327);
nor U3673 (N_3673,N_3486,N_3418);
nand U3674 (N_3674,N_3344,N_3388);
nand U3675 (N_3675,N_3420,N_3362);
and U3676 (N_3676,N_3377,N_3326);
nand U3677 (N_3677,N_3351,N_3384);
nand U3678 (N_3678,N_3478,N_3404);
or U3679 (N_3679,N_3444,N_3291);
nand U3680 (N_3680,N_3418,N_3402);
xnor U3681 (N_3681,N_3464,N_3468);
nor U3682 (N_3682,N_3402,N_3337);
xnor U3683 (N_3683,N_3472,N_3488);
nand U3684 (N_3684,N_3484,N_3396);
nor U3685 (N_3685,N_3342,N_3456);
xor U3686 (N_3686,N_3351,N_3355);
or U3687 (N_3687,N_3408,N_3281);
or U3688 (N_3688,N_3251,N_3344);
and U3689 (N_3689,N_3304,N_3484);
xor U3690 (N_3690,N_3412,N_3383);
or U3691 (N_3691,N_3325,N_3334);
or U3692 (N_3692,N_3363,N_3410);
xnor U3693 (N_3693,N_3280,N_3301);
nor U3694 (N_3694,N_3288,N_3454);
xnor U3695 (N_3695,N_3419,N_3352);
nand U3696 (N_3696,N_3263,N_3381);
nand U3697 (N_3697,N_3254,N_3361);
xor U3698 (N_3698,N_3444,N_3423);
nand U3699 (N_3699,N_3349,N_3397);
xor U3700 (N_3700,N_3291,N_3453);
xnor U3701 (N_3701,N_3320,N_3391);
xnor U3702 (N_3702,N_3276,N_3339);
xnor U3703 (N_3703,N_3384,N_3494);
nor U3704 (N_3704,N_3427,N_3434);
nor U3705 (N_3705,N_3358,N_3366);
nand U3706 (N_3706,N_3302,N_3311);
nor U3707 (N_3707,N_3309,N_3496);
nand U3708 (N_3708,N_3390,N_3294);
nor U3709 (N_3709,N_3462,N_3361);
nand U3710 (N_3710,N_3278,N_3457);
or U3711 (N_3711,N_3386,N_3254);
nand U3712 (N_3712,N_3369,N_3401);
nor U3713 (N_3713,N_3413,N_3385);
and U3714 (N_3714,N_3262,N_3469);
nor U3715 (N_3715,N_3350,N_3307);
xnor U3716 (N_3716,N_3447,N_3338);
or U3717 (N_3717,N_3445,N_3270);
and U3718 (N_3718,N_3378,N_3447);
or U3719 (N_3719,N_3484,N_3377);
nand U3720 (N_3720,N_3469,N_3488);
and U3721 (N_3721,N_3385,N_3272);
and U3722 (N_3722,N_3284,N_3251);
xor U3723 (N_3723,N_3255,N_3431);
nor U3724 (N_3724,N_3387,N_3263);
nor U3725 (N_3725,N_3257,N_3341);
nor U3726 (N_3726,N_3397,N_3411);
and U3727 (N_3727,N_3258,N_3307);
nor U3728 (N_3728,N_3311,N_3466);
xnor U3729 (N_3729,N_3257,N_3375);
nor U3730 (N_3730,N_3313,N_3378);
xor U3731 (N_3731,N_3297,N_3277);
xnor U3732 (N_3732,N_3262,N_3277);
nand U3733 (N_3733,N_3296,N_3283);
nand U3734 (N_3734,N_3485,N_3401);
or U3735 (N_3735,N_3379,N_3320);
nor U3736 (N_3736,N_3309,N_3258);
or U3737 (N_3737,N_3302,N_3351);
or U3738 (N_3738,N_3422,N_3370);
nor U3739 (N_3739,N_3452,N_3467);
and U3740 (N_3740,N_3445,N_3329);
and U3741 (N_3741,N_3299,N_3437);
xor U3742 (N_3742,N_3439,N_3374);
and U3743 (N_3743,N_3492,N_3271);
nor U3744 (N_3744,N_3414,N_3423);
or U3745 (N_3745,N_3468,N_3430);
or U3746 (N_3746,N_3282,N_3468);
nand U3747 (N_3747,N_3417,N_3305);
nand U3748 (N_3748,N_3265,N_3332);
and U3749 (N_3749,N_3329,N_3470);
nand U3750 (N_3750,N_3728,N_3746);
or U3751 (N_3751,N_3656,N_3524);
nor U3752 (N_3752,N_3749,N_3662);
nand U3753 (N_3753,N_3709,N_3520);
and U3754 (N_3754,N_3676,N_3504);
nor U3755 (N_3755,N_3645,N_3682);
nand U3756 (N_3756,N_3665,N_3693);
nor U3757 (N_3757,N_3711,N_3632);
nor U3758 (N_3758,N_3510,N_3516);
or U3759 (N_3759,N_3578,N_3560);
nand U3760 (N_3760,N_3678,N_3668);
xnor U3761 (N_3761,N_3585,N_3590);
and U3762 (N_3762,N_3705,N_3553);
xor U3763 (N_3763,N_3694,N_3624);
nand U3764 (N_3764,N_3597,N_3556);
or U3765 (N_3765,N_3538,N_3708);
nand U3766 (N_3766,N_3503,N_3661);
or U3767 (N_3767,N_3514,N_3589);
xnor U3768 (N_3768,N_3534,N_3639);
or U3769 (N_3769,N_3549,N_3716);
nand U3770 (N_3770,N_3614,N_3715);
or U3771 (N_3771,N_3544,N_3684);
and U3772 (N_3772,N_3506,N_3652);
and U3773 (N_3773,N_3622,N_3500);
or U3774 (N_3774,N_3733,N_3685);
xor U3775 (N_3775,N_3660,N_3601);
or U3776 (N_3776,N_3535,N_3558);
or U3777 (N_3777,N_3604,N_3568);
nor U3778 (N_3778,N_3546,N_3699);
xor U3779 (N_3779,N_3593,N_3689);
or U3780 (N_3780,N_3517,N_3648);
nor U3781 (N_3781,N_3629,N_3569);
nor U3782 (N_3782,N_3521,N_3547);
or U3783 (N_3783,N_3505,N_3673);
nand U3784 (N_3784,N_3743,N_3653);
and U3785 (N_3785,N_3714,N_3518);
and U3786 (N_3786,N_3515,N_3586);
or U3787 (N_3787,N_3532,N_3721);
nor U3788 (N_3788,N_3598,N_3666);
and U3789 (N_3789,N_3557,N_3696);
or U3790 (N_3790,N_3640,N_3536);
or U3791 (N_3791,N_3621,N_3611);
nand U3792 (N_3792,N_3643,N_3508);
or U3793 (N_3793,N_3595,N_3579);
or U3794 (N_3794,N_3695,N_3594);
nand U3795 (N_3795,N_3683,N_3607);
and U3796 (N_3796,N_3634,N_3548);
xor U3797 (N_3797,N_3727,N_3651);
nand U3798 (N_3798,N_3550,N_3596);
nor U3799 (N_3799,N_3576,N_3541);
nor U3800 (N_3800,N_3512,N_3735);
xor U3801 (N_3801,N_3738,N_3628);
nor U3802 (N_3802,N_3613,N_3582);
and U3803 (N_3803,N_3667,N_3664);
nand U3804 (N_3804,N_3719,N_3572);
or U3805 (N_3805,N_3744,N_3531);
and U3806 (N_3806,N_3574,N_3600);
nand U3807 (N_3807,N_3539,N_3713);
nand U3808 (N_3808,N_3740,N_3729);
and U3809 (N_3809,N_3599,N_3573);
xnor U3810 (N_3810,N_3525,N_3543);
and U3811 (N_3811,N_3633,N_3575);
nor U3812 (N_3812,N_3565,N_3663);
and U3813 (N_3813,N_3670,N_3702);
nand U3814 (N_3814,N_3731,N_3567);
and U3815 (N_3815,N_3561,N_3644);
nand U3816 (N_3816,N_3507,N_3566);
or U3817 (N_3817,N_3583,N_3509);
or U3818 (N_3818,N_3584,N_3712);
xor U3819 (N_3819,N_3703,N_3623);
xor U3820 (N_3820,N_3502,N_3739);
nor U3821 (N_3821,N_3698,N_3537);
and U3822 (N_3822,N_3642,N_3625);
nand U3823 (N_3823,N_3737,N_3542);
xnor U3824 (N_3824,N_3707,N_3527);
xor U3825 (N_3825,N_3618,N_3615);
nor U3826 (N_3826,N_3616,N_3501);
nor U3827 (N_3827,N_3649,N_3747);
nor U3828 (N_3828,N_3552,N_3617);
and U3829 (N_3829,N_3559,N_3641);
or U3830 (N_3830,N_3669,N_3671);
and U3831 (N_3831,N_3706,N_3674);
nand U3832 (N_3832,N_3717,N_3647);
and U3833 (N_3833,N_3554,N_3655);
and U3834 (N_3834,N_3730,N_3697);
nor U3835 (N_3835,N_3700,N_3687);
or U3836 (N_3836,N_3533,N_3522);
or U3837 (N_3837,N_3636,N_3690);
nor U3838 (N_3838,N_3686,N_3608);
xor U3839 (N_3839,N_3732,N_3724);
nor U3840 (N_3840,N_3609,N_3606);
xnor U3841 (N_3841,N_3602,N_3701);
or U3842 (N_3842,N_3511,N_3741);
or U3843 (N_3843,N_3726,N_3675);
or U3844 (N_3844,N_3605,N_3637);
and U3845 (N_3845,N_3654,N_3734);
nand U3846 (N_3846,N_3610,N_3545);
nor U3847 (N_3847,N_3603,N_3745);
and U3848 (N_3848,N_3627,N_3526);
nand U3849 (N_3849,N_3620,N_3681);
xor U3850 (N_3850,N_3562,N_3580);
nand U3851 (N_3851,N_3592,N_3551);
nand U3852 (N_3852,N_3680,N_3555);
xnor U3853 (N_3853,N_3748,N_3672);
xor U3854 (N_3854,N_3657,N_3619);
and U3855 (N_3855,N_3723,N_3742);
or U3856 (N_3856,N_3677,N_3679);
and U3857 (N_3857,N_3650,N_3588);
and U3858 (N_3858,N_3736,N_3530);
xor U3859 (N_3859,N_3570,N_3591);
and U3860 (N_3860,N_3577,N_3513);
xor U3861 (N_3861,N_3563,N_3631);
or U3862 (N_3862,N_3691,N_3581);
xnor U3863 (N_3863,N_3528,N_3722);
nor U3864 (N_3864,N_3523,N_3612);
nor U3865 (N_3865,N_3587,N_3630);
nand U3866 (N_3866,N_3659,N_3718);
or U3867 (N_3867,N_3571,N_3710);
xor U3868 (N_3868,N_3635,N_3658);
nor U3869 (N_3869,N_3564,N_3688);
nand U3870 (N_3870,N_3519,N_3692);
nor U3871 (N_3871,N_3725,N_3540);
nand U3872 (N_3872,N_3720,N_3704);
and U3873 (N_3873,N_3529,N_3646);
nor U3874 (N_3874,N_3626,N_3638);
nand U3875 (N_3875,N_3614,N_3626);
nand U3876 (N_3876,N_3718,N_3554);
nand U3877 (N_3877,N_3742,N_3692);
nor U3878 (N_3878,N_3694,N_3586);
xor U3879 (N_3879,N_3600,N_3737);
nor U3880 (N_3880,N_3542,N_3658);
xnor U3881 (N_3881,N_3728,N_3749);
nor U3882 (N_3882,N_3724,N_3558);
nand U3883 (N_3883,N_3629,N_3566);
nand U3884 (N_3884,N_3671,N_3710);
or U3885 (N_3885,N_3602,N_3546);
and U3886 (N_3886,N_3676,N_3654);
and U3887 (N_3887,N_3689,N_3698);
and U3888 (N_3888,N_3636,N_3670);
or U3889 (N_3889,N_3666,N_3575);
nand U3890 (N_3890,N_3656,N_3681);
or U3891 (N_3891,N_3642,N_3671);
xnor U3892 (N_3892,N_3604,N_3666);
or U3893 (N_3893,N_3662,N_3538);
and U3894 (N_3894,N_3575,N_3675);
and U3895 (N_3895,N_3581,N_3571);
nand U3896 (N_3896,N_3665,N_3582);
xor U3897 (N_3897,N_3617,N_3734);
nor U3898 (N_3898,N_3680,N_3544);
or U3899 (N_3899,N_3555,N_3721);
or U3900 (N_3900,N_3543,N_3738);
or U3901 (N_3901,N_3533,N_3535);
nor U3902 (N_3902,N_3726,N_3576);
nand U3903 (N_3903,N_3633,N_3707);
nand U3904 (N_3904,N_3667,N_3546);
and U3905 (N_3905,N_3602,N_3527);
nor U3906 (N_3906,N_3706,N_3540);
or U3907 (N_3907,N_3535,N_3629);
or U3908 (N_3908,N_3562,N_3732);
and U3909 (N_3909,N_3716,N_3663);
nor U3910 (N_3910,N_3557,N_3552);
nand U3911 (N_3911,N_3641,N_3597);
or U3912 (N_3912,N_3690,N_3747);
and U3913 (N_3913,N_3530,N_3554);
xnor U3914 (N_3914,N_3714,N_3525);
xnor U3915 (N_3915,N_3529,N_3561);
and U3916 (N_3916,N_3741,N_3541);
and U3917 (N_3917,N_3635,N_3732);
xnor U3918 (N_3918,N_3610,N_3572);
and U3919 (N_3919,N_3700,N_3642);
or U3920 (N_3920,N_3642,N_3727);
or U3921 (N_3921,N_3652,N_3573);
or U3922 (N_3922,N_3622,N_3623);
or U3923 (N_3923,N_3628,N_3505);
xor U3924 (N_3924,N_3534,N_3571);
and U3925 (N_3925,N_3532,N_3523);
or U3926 (N_3926,N_3594,N_3710);
nor U3927 (N_3927,N_3717,N_3619);
nor U3928 (N_3928,N_3663,N_3610);
and U3929 (N_3929,N_3558,N_3621);
nand U3930 (N_3930,N_3670,N_3666);
xor U3931 (N_3931,N_3696,N_3515);
and U3932 (N_3932,N_3718,N_3739);
xnor U3933 (N_3933,N_3590,N_3749);
xor U3934 (N_3934,N_3691,N_3636);
and U3935 (N_3935,N_3703,N_3709);
nor U3936 (N_3936,N_3503,N_3695);
nor U3937 (N_3937,N_3506,N_3610);
and U3938 (N_3938,N_3710,N_3609);
xnor U3939 (N_3939,N_3663,N_3566);
nand U3940 (N_3940,N_3631,N_3693);
or U3941 (N_3941,N_3592,N_3730);
xnor U3942 (N_3942,N_3541,N_3603);
xor U3943 (N_3943,N_3519,N_3696);
nand U3944 (N_3944,N_3665,N_3617);
or U3945 (N_3945,N_3662,N_3608);
nor U3946 (N_3946,N_3514,N_3707);
xnor U3947 (N_3947,N_3602,N_3637);
nor U3948 (N_3948,N_3671,N_3738);
and U3949 (N_3949,N_3648,N_3548);
xor U3950 (N_3950,N_3669,N_3548);
and U3951 (N_3951,N_3590,N_3624);
xor U3952 (N_3952,N_3731,N_3681);
or U3953 (N_3953,N_3505,N_3634);
nand U3954 (N_3954,N_3561,N_3508);
or U3955 (N_3955,N_3633,N_3621);
or U3956 (N_3956,N_3583,N_3508);
nor U3957 (N_3957,N_3657,N_3709);
and U3958 (N_3958,N_3730,N_3657);
xnor U3959 (N_3959,N_3505,N_3530);
or U3960 (N_3960,N_3678,N_3557);
xnor U3961 (N_3961,N_3707,N_3513);
and U3962 (N_3962,N_3597,N_3681);
nand U3963 (N_3963,N_3747,N_3517);
or U3964 (N_3964,N_3575,N_3725);
nor U3965 (N_3965,N_3724,N_3563);
or U3966 (N_3966,N_3620,N_3727);
xnor U3967 (N_3967,N_3559,N_3685);
nand U3968 (N_3968,N_3746,N_3617);
nand U3969 (N_3969,N_3606,N_3505);
or U3970 (N_3970,N_3633,N_3706);
nor U3971 (N_3971,N_3736,N_3659);
nand U3972 (N_3972,N_3581,N_3531);
xnor U3973 (N_3973,N_3713,N_3503);
or U3974 (N_3974,N_3567,N_3624);
or U3975 (N_3975,N_3590,N_3611);
xnor U3976 (N_3976,N_3630,N_3715);
nor U3977 (N_3977,N_3746,N_3531);
xor U3978 (N_3978,N_3530,N_3523);
xor U3979 (N_3979,N_3599,N_3604);
nand U3980 (N_3980,N_3602,N_3599);
nand U3981 (N_3981,N_3740,N_3589);
nor U3982 (N_3982,N_3561,N_3586);
xor U3983 (N_3983,N_3578,N_3682);
or U3984 (N_3984,N_3526,N_3582);
nand U3985 (N_3985,N_3567,N_3527);
and U3986 (N_3986,N_3587,N_3579);
nand U3987 (N_3987,N_3598,N_3719);
nor U3988 (N_3988,N_3654,N_3666);
nor U3989 (N_3989,N_3519,N_3534);
nand U3990 (N_3990,N_3723,N_3719);
and U3991 (N_3991,N_3530,N_3586);
nor U3992 (N_3992,N_3515,N_3529);
xor U3993 (N_3993,N_3529,N_3660);
xnor U3994 (N_3994,N_3647,N_3516);
or U3995 (N_3995,N_3598,N_3566);
xnor U3996 (N_3996,N_3673,N_3621);
nand U3997 (N_3997,N_3708,N_3529);
nand U3998 (N_3998,N_3676,N_3530);
and U3999 (N_3999,N_3506,N_3691);
nand U4000 (N_4000,N_3923,N_3903);
or U4001 (N_4001,N_3803,N_3882);
xor U4002 (N_4002,N_3999,N_3811);
or U4003 (N_4003,N_3754,N_3928);
nor U4004 (N_4004,N_3891,N_3935);
nand U4005 (N_4005,N_3852,N_3820);
xor U4006 (N_4006,N_3915,N_3981);
xnor U4007 (N_4007,N_3775,N_3782);
nor U4008 (N_4008,N_3830,N_3792);
xnor U4009 (N_4009,N_3844,N_3819);
or U4010 (N_4010,N_3965,N_3990);
or U4011 (N_4011,N_3791,N_3900);
or U4012 (N_4012,N_3894,N_3950);
xor U4013 (N_4013,N_3947,N_3925);
nor U4014 (N_4014,N_3941,N_3851);
or U4015 (N_4015,N_3765,N_3942);
nand U4016 (N_4016,N_3822,N_3829);
nand U4017 (N_4017,N_3808,N_3798);
and U4018 (N_4018,N_3847,N_3889);
and U4019 (N_4019,N_3839,N_3868);
or U4020 (N_4020,N_3899,N_3908);
nand U4021 (N_4021,N_3979,N_3897);
xor U4022 (N_4022,N_3895,N_3930);
xor U4023 (N_4023,N_3859,N_3773);
xnor U4024 (N_4024,N_3848,N_3814);
nor U4025 (N_4025,N_3837,N_3813);
nand U4026 (N_4026,N_3910,N_3907);
or U4027 (N_4027,N_3783,N_3956);
or U4028 (N_4028,N_3969,N_3764);
nand U4029 (N_4029,N_3939,N_3761);
and U4030 (N_4030,N_3875,N_3784);
nand U4031 (N_4031,N_3809,N_3790);
nand U4032 (N_4032,N_3873,N_3821);
xor U4033 (N_4033,N_3975,N_3867);
nor U4034 (N_4034,N_3805,N_3982);
and U4035 (N_4035,N_3849,N_3824);
nand U4036 (N_4036,N_3856,N_3924);
xnor U4037 (N_4037,N_3962,N_3948);
and U4038 (N_4038,N_3788,N_3978);
nand U4039 (N_4039,N_3931,N_3926);
nor U4040 (N_4040,N_3957,N_3911);
xnor U4041 (N_4041,N_3817,N_3758);
or U4042 (N_4042,N_3987,N_3943);
and U4043 (N_4043,N_3976,N_3878);
nor U4044 (N_4044,N_3883,N_3785);
xnor U4045 (N_4045,N_3920,N_3946);
nor U4046 (N_4046,N_3906,N_3996);
xnor U4047 (N_4047,N_3905,N_3973);
nor U4048 (N_4048,N_3917,N_3855);
nand U4049 (N_4049,N_3961,N_3995);
and U4050 (N_4050,N_3879,N_3834);
xor U4051 (N_4051,N_3968,N_3967);
nand U4052 (N_4052,N_3789,N_3771);
and U4053 (N_4053,N_3832,N_3945);
nor U4054 (N_4054,N_3958,N_3760);
nand U4055 (N_4055,N_3767,N_3794);
and U4056 (N_4056,N_3870,N_3826);
and U4057 (N_4057,N_3853,N_3985);
nand U4058 (N_4058,N_3971,N_3828);
nand U4059 (N_4059,N_3772,N_3901);
and U4060 (N_4060,N_3762,N_3777);
xnor U4061 (N_4061,N_3862,N_3838);
and U4062 (N_4062,N_3833,N_3921);
xor U4063 (N_4063,N_3866,N_3937);
xnor U4064 (N_4064,N_3993,N_3984);
xnor U4065 (N_4065,N_3970,N_3904);
or U4066 (N_4066,N_3845,N_3799);
nor U4067 (N_4067,N_3932,N_3869);
and U4068 (N_4068,N_3954,N_3831);
nor U4069 (N_4069,N_3994,N_3843);
and U4070 (N_4070,N_3780,N_3887);
and U4071 (N_4071,N_3888,N_3877);
or U4072 (N_4072,N_3840,N_3757);
nor U4073 (N_4073,N_3779,N_3774);
nand U4074 (N_4074,N_3801,N_3919);
and U4075 (N_4075,N_3896,N_3863);
nor U4076 (N_4076,N_3865,N_3763);
and U4077 (N_4077,N_3796,N_3854);
or U4078 (N_4078,N_3955,N_3909);
and U4079 (N_4079,N_3972,N_3850);
xor U4080 (N_4080,N_3823,N_3871);
or U4081 (N_4081,N_3934,N_3997);
or U4082 (N_4082,N_3918,N_3912);
nor U4083 (N_4083,N_3940,N_3818);
xor U4084 (N_4084,N_3781,N_3806);
xor U4085 (N_4085,N_3766,N_3890);
and U4086 (N_4086,N_3751,N_3927);
nor U4087 (N_4087,N_3756,N_3815);
nand U4088 (N_4088,N_3989,N_3768);
or U4089 (N_4089,N_3892,N_3846);
or U4090 (N_4090,N_3860,N_3963);
xnor U4091 (N_4091,N_3872,N_3960);
xnor U4092 (N_4092,N_3770,N_3835);
and U4093 (N_4093,N_3816,N_3842);
nand U4094 (N_4094,N_3884,N_3755);
or U4095 (N_4095,N_3793,N_3800);
or U4096 (N_4096,N_3812,N_3752);
or U4097 (N_4097,N_3759,N_3953);
nand U4098 (N_4098,N_3880,N_3836);
nand U4099 (N_4099,N_3876,N_3974);
nand U4100 (N_4100,N_3913,N_3857);
and U4101 (N_4101,N_3949,N_3776);
or U4102 (N_4102,N_3750,N_3914);
or U4103 (N_4103,N_3804,N_3988);
nand U4104 (N_4104,N_3786,N_3886);
or U4105 (N_4105,N_3810,N_3902);
nor U4106 (N_4106,N_3861,N_3922);
xor U4107 (N_4107,N_3769,N_3898);
nand U4108 (N_4108,N_3797,N_3980);
nand U4109 (N_4109,N_3959,N_3795);
or U4110 (N_4110,N_3753,N_3936);
or U4111 (N_4111,N_3944,N_3807);
or U4112 (N_4112,N_3933,N_3964);
and U4113 (N_4113,N_3841,N_3983);
nand U4114 (N_4114,N_3929,N_3874);
or U4115 (N_4115,N_3825,N_3778);
nand U4116 (N_4116,N_3977,N_3858);
xnor U4117 (N_4117,N_3893,N_3992);
nor U4118 (N_4118,N_3951,N_3938);
nor U4119 (N_4119,N_3991,N_3986);
nand U4120 (N_4120,N_3881,N_3998);
and U4121 (N_4121,N_3885,N_3802);
xor U4122 (N_4122,N_3864,N_3966);
xor U4123 (N_4123,N_3787,N_3916);
nand U4124 (N_4124,N_3952,N_3827);
and U4125 (N_4125,N_3801,N_3867);
or U4126 (N_4126,N_3795,N_3803);
and U4127 (N_4127,N_3855,N_3766);
and U4128 (N_4128,N_3926,N_3943);
and U4129 (N_4129,N_3754,N_3964);
nand U4130 (N_4130,N_3808,N_3986);
and U4131 (N_4131,N_3822,N_3981);
nand U4132 (N_4132,N_3911,N_3821);
and U4133 (N_4133,N_3977,N_3760);
xor U4134 (N_4134,N_3839,N_3781);
or U4135 (N_4135,N_3870,N_3818);
xnor U4136 (N_4136,N_3920,N_3918);
xor U4137 (N_4137,N_3836,N_3898);
xor U4138 (N_4138,N_3828,N_3939);
nand U4139 (N_4139,N_3808,N_3900);
or U4140 (N_4140,N_3880,N_3988);
or U4141 (N_4141,N_3947,N_3858);
xnor U4142 (N_4142,N_3920,N_3907);
nor U4143 (N_4143,N_3948,N_3820);
nand U4144 (N_4144,N_3838,N_3822);
nor U4145 (N_4145,N_3876,N_3853);
xor U4146 (N_4146,N_3801,N_3845);
or U4147 (N_4147,N_3932,N_3773);
xor U4148 (N_4148,N_3907,N_3924);
and U4149 (N_4149,N_3920,N_3992);
and U4150 (N_4150,N_3833,N_3866);
nand U4151 (N_4151,N_3755,N_3891);
and U4152 (N_4152,N_3815,N_3941);
and U4153 (N_4153,N_3968,N_3884);
nand U4154 (N_4154,N_3953,N_3819);
and U4155 (N_4155,N_3841,N_3996);
and U4156 (N_4156,N_3756,N_3861);
nand U4157 (N_4157,N_3895,N_3918);
or U4158 (N_4158,N_3757,N_3835);
and U4159 (N_4159,N_3991,N_3792);
and U4160 (N_4160,N_3937,N_3973);
and U4161 (N_4161,N_3978,N_3998);
xor U4162 (N_4162,N_3924,N_3898);
nand U4163 (N_4163,N_3860,N_3896);
or U4164 (N_4164,N_3858,N_3950);
nor U4165 (N_4165,N_3865,N_3858);
nand U4166 (N_4166,N_3883,N_3763);
nand U4167 (N_4167,N_3982,N_3903);
xnor U4168 (N_4168,N_3993,N_3792);
nand U4169 (N_4169,N_3988,N_3839);
or U4170 (N_4170,N_3775,N_3889);
or U4171 (N_4171,N_3917,N_3901);
nor U4172 (N_4172,N_3970,N_3807);
nand U4173 (N_4173,N_3851,N_3936);
xor U4174 (N_4174,N_3828,N_3959);
nand U4175 (N_4175,N_3803,N_3841);
xnor U4176 (N_4176,N_3984,N_3813);
nand U4177 (N_4177,N_3961,N_3999);
nand U4178 (N_4178,N_3876,N_3787);
nor U4179 (N_4179,N_3972,N_3779);
or U4180 (N_4180,N_3824,N_3828);
or U4181 (N_4181,N_3821,N_3954);
and U4182 (N_4182,N_3920,N_3820);
or U4183 (N_4183,N_3861,N_3991);
and U4184 (N_4184,N_3790,N_3929);
nor U4185 (N_4185,N_3847,N_3885);
or U4186 (N_4186,N_3877,N_3850);
and U4187 (N_4187,N_3897,N_3787);
nor U4188 (N_4188,N_3950,N_3762);
xnor U4189 (N_4189,N_3923,N_3762);
or U4190 (N_4190,N_3839,N_3885);
xnor U4191 (N_4191,N_3879,N_3856);
nor U4192 (N_4192,N_3899,N_3946);
nor U4193 (N_4193,N_3904,N_3821);
and U4194 (N_4194,N_3902,N_3899);
nand U4195 (N_4195,N_3816,N_3807);
and U4196 (N_4196,N_3824,N_3894);
nor U4197 (N_4197,N_3936,N_3876);
nor U4198 (N_4198,N_3964,N_3941);
and U4199 (N_4199,N_3978,N_3759);
or U4200 (N_4200,N_3786,N_3835);
or U4201 (N_4201,N_3754,N_3981);
nor U4202 (N_4202,N_3841,N_3773);
or U4203 (N_4203,N_3872,N_3813);
xor U4204 (N_4204,N_3915,N_3824);
nor U4205 (N_4205,N_3817,N_3777);
nand U4206 (N_4206,N_3794,N_3797);
and U4207 (N_4207,N_3809,N_3978);
nor U4208 (N_4208,N_3755,N_3999);
and U4209 (N_4209,N_3860,N_3858);
nand U4210 (N_4210,N_3939,N_3908);
and U4211 (N_4211,N_3932,N_3944);
and U4212 (N_4212,N_3874,N_3882);
xor U4213 (N_4213,N_3858,N_3857);
nor U4214 (N_4214,N_3876,N_3867);
xor U4215 (N_4215,N_3780,N_3752);
nand U4216 (N_4216,N_3760,N_3995);
nand U4217 (N_4217,N_3894,N_3819);
xnor U4218 (N_4218,N_3951,N_3830);
nor U4219 (N_4219,N_3881,N_3811);
and U4220 (N_4220,N_3995,N_3976);
nor U4221 (N_4221,N_3761,N_3947);
and U4222 (N_4222,N_3813,N_3753);
and U4223 (N_4223,N_3892,N_3972);
nor U4224 (N_4224,N_3827,N_3804);
nand U4225 (N_4225,N_3990,N_3874);
and U4226 (N_4226,N_3842,N_3921);
nor U4227 (N_4227,N_3958,N_3791);
and U4228 (N_4228,N_3824,N_3830);
or U4229 (N_4229,N_3911,N_3885);
and U4230 (N_4230,N_3811,N_3853);
nor U4231 (N_4231,N_3826,N_3859);
or U4232 (N_4232,N_3761,N_3940);
and U4233 (N_4233,N_3831,N_3803);
or U4234 (N_4234,N_3805,N_3847);
nand U4235 (N_4235,N_3928,N_3860);
and U4236 (N_4236,N_3910,N_3900);
and U4237 (N_4237,N_3944,N_3894);
nand U4238 (N_4238,N_3885,N_3979);
or U4239 (N_4239,N_3999,N_3889);
xnor U4240 (N_4240,N_3978,N_3811);
or U4241 (N_4241,N_3781,N_3818);
and U4242 (N_4242,N_3769,N_3876);
nand U4243 (N_4243,N_3947,N_3780);
nand U4244 (N_4244,N_3811,N_3816);
or U4245 (N_4245,N_3858,N_3990);
xnor U4246 (N_4246,N_3868,N_3892);
nand U4247 (N_4247,N_3846,N_3916);
nor U4248 (N_4248,N_3931,N_3903);
xor U4249 (N_4249,N_3961,N_3898);
and U4250 (N_4250,N_4058,N_4205);
xnor U4251 (N_4251,N_4004,N_4007);
and U4252 (N_4252,N_4233,N_4193);
nor U4253 (N_4253,N_4024,N_4075);
nand U4254 (N_4254,N_4104,N_4034);
or U4255 (N_4255,N_4150,N_4141);
xnor U4256 (N_4256,N_4006,N_4207);
nor U4257 (N_4257,N_4076,N_4210);
or U4258 (N_4258,N_4026,N_4091);
xnor U4259 (N_4259,N_4096,N_4227);
or U4260 (N_4260,N_4135,N_4018);
nand U4261 (N_4261,N_4171,N_4070);
nand U4262 (N_4262,N_4093,N_4248);
or U4263 (N_4263,N_4048,N_4125);
nor U4264 (N_4264,N_4116,N_4161);
xnor U4265 (N_4265,N_4221,N_4173);
nand U4266 (N_4266,N_4149,N_4169);
or U4267 (N_4267,N_4080,N_4202);
and U4268 (N_4268,N_4234,N_4030);
and U4269 (N_4269,N_4201,N_4158);
or U4270 (N_4270,N_4164,N_4146);
xnor U4271 (N_4271,N_4130,N_4177);
xor U4272 (N_4272,N_4047,N_4072);
and U4273 (N_4273,N_4245,N_4203);
and U4274 (N_4274,N_4056,N_4038);
nor U4275 (N_4275,N_4153,N_4224);
nand U4276 (N_4276,N_4138,N_4215);
or U4277 (N_4277,N_4021,N_4032);
xor U4278 (N_4278,N_4217,N_4228);
xnor U4279 (N_4279,N_4157,N_4129);
or U4280 (N_4280,N_4092,N_4049);
and U4281 (N_4281,N_4073,N_4220);
or U4282 (N_4282,N_4187,N_4074);
nor U4283 (N_4283,N_4112,N_4022);
nand U4284 (N_4284,N_4062,N_4102);
or U4285 (N_4285,N_4110,N_4154);
and U4286 (N_4286,N_4106,N_4059);
nand U4287 (N_4287,N_4061,N_4023);
and U4288 (N_4288,N_4136,N_4063);
and U4289 (N_4289,N_4140,N_4042);
nor U4290 (N_4290,N_4185,N_4095);
xnor U4291 (N_4291,N_4176,N_4094);
xnor U4292 (N_4292,N_4001,N_4015);
or U4293 (N_4293,N_4077,N_4081);
or U4294 (N_4294,N_4238,N_4100);
or U4295 (N_4295,N_4151,N_4208);
and U4296 (N_4296,N_4053,N_4046);
nand U4297 (N_4297,N_4108,N_4137);
or U4298 (N_4298,N_4060,N_4163);
nor U4299 (N_4299,N_4000,N_4249);
xor U4300 (N_4300,N_4064,N_4044);
and U4301 (N_4301,N_4120,N_4019);
and U4302 (N_4302,N_4170,N_4231);
xnor U4303 (N_4303,N_4243,N_4127);
nand U4304 (N_4304,N_4237,N_4174);
or U4305 (N_4305,N_4068,N_4065);
nor U4306 (N_4306,N_4118,N_4098);
nand U4307 (N_4307,N_4235,N_4230);
nand U4308 (N_4308,N_4041,N_4086);
nand U4309 (N_4309,N_4020,N_4197);
and U4310 (N_4310,N_4155,N_4101);
nand U4311 (N_4311,N_4142,N_4051);
nand U4312 (N_4312,N_4111,N_4114);
nand U4313 (N_4313,N_4082,N_4180);
xor U4314 (N_4314,N_4036,N_4222);
and U4315 (N_4315,N_4010,N_4219);
and U4316 (N_4316,N_4045,N_4186);
nor U4317 (N_4317,N_4002,N_4078);
or U4318 (N_4318,N_4126,N_4239);
xnor U4319 (N_4319,N_4226,N_4121);
or U4320 (N_4320,N_4028,N_4069);
and U4321 (N_4321,N_4009,N_4213);
xor U4322 (N_4322,N_4206,N_4159);
nand U4323 (N_4323,N_4122,N_4160);
nand U4324 (N_4324,N_4216,N_4033);
xnor U4325 (N_4325,N_4218,N_4200);
nand U4326 (N_4326,N_4166,N_4017);
nor U4327 (N_4327,N_4040,N_4192);
nor U4328 (N_4328,N_4145,N_4131);
and U4329 (N_4329,N_4152,N_4223);
nor U4330 (N_4330,N_4172,N_4246);
or U4331 (N_4331,N_4052,N_4005);
and U4332 (N_4332,N_4128,N_4109);
and U4333 (N_4333,N_4247,N_4008);
or U4334 (N_4334,N_4117,N_4241);
or U4335 (N_4335,N_4167,N_4242);
nand U4336 (N_4336,N_4043,N_4057);
xor U4337 (N_4337,N_4012,N_4194);
or U4338 (N_4338,N_4212,N_4105);
nor U4339 (N_4339,N_4025,N_4211);
nor U4340 (N_4340,N_4236,N_4147);
nand U4341 (N_4341,N_4123,N_4035);
and U4342 (N_4342,N_4144,N_4079);
xor U4343 (N_4343,N_4156,N_4067);
xnor U4344 (N_4344,N_4087,N_4085);
and U4345 (N_4345,N_4099,N_4209);
or U4346 (N_4346,N_4179,N_4011);
and U4347 (N_4347,N_4133,N_4182);
xnor U4348 (N_4348,N_4016,N_4013);
and U4349 (N_4349,N_4071,N_4214);
or U4350 (N_4350,N_4066,N_4240);
nand U4351 (N_4351,N_4103,N_4083);
and U4352 (N_4352,N_4029,N_4175);
nand U4353 (N_4353,N_4119,N_4014);
and U4354 (N_4354,N_4148,N_4181);
nand U4355 (N_4355,N_4055,N_4027);
and U4356 (N_4356,N_4031,N_4037);
xor U4357 (N_4357,N_4039,N_4139);
and U4358 (N_4358,N_4184,N_4143);
and U4359 (N_4359,N_4232,N_4188);
nor U4360 (N_4360,N_4089,N_4189);
or U4361 (N_4361,N_4050,N_4178);
nand U4362 (N_4362,N_4124,N_4225);
and U4363 (N_4363,N_4244,N_4191);
and U4364 (N_4364,N_4183,N_4003);
xor U4365 (N_4365,N_4134,N_4090);
and U4366 (N_4366,N_4165,N_4054);
nor U4367 (N_4367,N_4107,N_4229);
and U4368 (N_4368,N_4195,N_4088);
and U4369 (N_4369,N_4113,N_4196);
and U4370 (N_4370,N_4198,N_4168);
xnor U4371 (N_4371,N_4162,N_4204);
or U4372 (N_4372,N_4084,N_4199);
nor U4373 (N_4373,N_4115,N_4097);
and U4374 (N_4374,N_4132,N_4190);
nor U4375 (N_4375,N_4159,N_4201);
nor U4376 (N_4376,N_4028,N_4146);
or U4377 (N_4377,N_4083,N_4126);
nor U4378 (N_4378,N_4033,N_4098);
nand U4379 (N_4379,N_4085,N_4138);
nand U4380 (N_4380,N_4197,N_4019);
nor U4381 (N_4381,N_4108,N_4202);
and U4382 (N_4382,N_4184,N_4017);
and U4383 (N_4383,N_4121,N_4006);
xnor U4384 (N_4384,N_4207,N_4024);
nor U4385 (N_4385,N_4143,N_4188);
or U4386 (N_4386,N_4013,N_4179);
xor U4387 (N_4387,N_4002,N_4191);
or U4388 (N_4388,N_4098,N_4141);
and U4389 (N_4389,N_4228,N_4235);
nand U4390 (N_4390,N_4102,N_4115);
xnor U4391 (N_4391,N_4139,N_4172);
and U4392 (N_4392,N_4124,N_4183);
or U4393 (N_4393,N_4141,N_4060);
nand U4394 (N_4394,N_4001,N_4073);
nor U4395 (N_4395,N_4155,N_4158);
nor U4396 (N_4396,N_4194,N_4061);
and U4397 (N_4397,N_4043,N_4210);
or U4398 (N_4398,N_4086,N_4139);
xor U4399 (N_4399,N_4017,N_4173);
xor U4400 (N_4400,N_4093,N_4084);
or U4401 (N_4401,N_4165,N_4238);
or U4402 (N_4402,N_4219,N_4030);
or U4403 (N_4403,N_4103,N_4097);
or U4404 (N_4404,N_4095,N_4023);
nor U4405 (N_4405,N_4068,N_4154);
nand U4406 (N_4406,N_4216,N_4234);
xnor U4407 (N_4407,N_4116,N_4009);
xor U4408 (N_4408,N_4036,N_4093);
and U4409 (N_4409,N_4037,N_4197);
and U4410 (N_4410,N_4128,N_4091);
xnor U4411 (N_4411,N_4076,N_4200);
or U4412 (N_4412,N_4059,N_4014);
nor U4413 (N_4413,N_4037,N_4167);
nor U4414 (N_4414,N_4080,N_4174);
nand U4415 (N_4415,N_4111,N_4004);
nand U4416 (N_4416,N_4242,N_4155);
or U4417 (N_4417,N_4005,N_4023);
and U4418 (N_4418,N_4181,N_4099);
nor U4419 (N_4419,N_4193,N_4028);
and U4420 (N_4420,N_4111,N_4229);
nor U4421 (N_4421,N_4121,N_4120);
xnor U4422 (N_4422,N_4233,N_4077);
and U4423 (N_4423,N_4218,N_4060);
or U4424 (N_4424,N_4086,N_4082);
xnor U4425 (N_4425,N_4152,N_4164);
nand U4426 (N_4426,N_4209,N_4157);
or U4427 (N_4427,N_4046,N_4200);
nand U4428 (N_4428,N_4224,N_4183);
and U4429 (N_4429,N_4223,N_4117);
xnor U4430 (N_4430,N_4125,N_4045);
or U4431 (N_4431,N_4065,N_4175);
or U4432 (N_4432,N_4177,N_4131);
and U4433 (N_4433,N_4195,N_4029);
nand U4434 (N_4434,N_4198,N_4047);
nor U4435 (N_4435,N_4110,N_4227);
or U4436 (N_4436,N_4176,N_4044);
nor U4437 (N_4437,N_4248,N_4051);
nand U4438 (N_4438,N_4148,N_4059);
or U4439 (N_4439,N_4153,N_4204);
or U4440 (N_4440,N_4092,N_4151);
and U4441 (N_4441,N_4101,N_4099);
or U4442 (N_4442,N_4074,N_4184);
xor U4443 (N_4443,N_4238,N_4019);
xor U4444 (N_4444,N_4215,N_4240);
nand U4445 (N_4445,N_4086,N_4170);
or U4446 (N_4446,N_4077,N_4183);
nor U4447 (N_4447,N_4202,N_4102);
and U4448 (N_4448,N_4226,N_4072);
nand U4449 (N_4449,N_4233,N_4107);
or U4450 (N_4450,N_4221,N_4147);
nand U4451 (N_4451,N_4077,N_4197);
or U4452 (N_4452,N_4035,N_4033);
nor U4453 (N_4453,N_4031,N_4081);
nand U4454 (N_4454,N_4093,N_4034);
or U4455 (N_4455,N_4044,N_4018);
xor U4456 (N_4456,N_4084,N_4070);
xor U4457 (N_4457,N_4008,N_4055);
and U4458 (N_4458,N_4024,N_4176);
nor U4459 (N_4459,N_4009,N_4138);
xnor U4460 (N_4460,N_4153,N_4134);
nand U4461 (N_4461,N_4237,N_4033);
xor U4462 (N_4462,N_4149,N_4002);
xor U4463 (N_4463,N_4217,N_4175);
and U4464 (N_4464,N_4224,N_4002);
and U4465 (N_4465,N_4235,N_4180);
xor U4466 (N_4466,N_4052,N_4102);
xnor U4467 (N_4467,N_4159,N_4207);
and U4468 (N_4468,N_4152,N_4249);
xnor U4469 (N_4469,N_4137,N_4192);
nor U4470 (N_4470,N_4150,N_4133);
or U4471 (N_4471,N_4028,N_4023);
and U4472 (N_4472,N_4216,N_4198);
xor U4473 (N_4473,N_4207,N_4214);
or U4474 (N_4474,N_4093,N_4216);
nand U4475 (N_4475,N_4206,N_4232);
or U4476 (N_4476,N_4215,N_4181);
nor U4477 (N_4477,N_4021,N_4066);
and U4478 (N_4478,N_4113,N_4152);
nor U4479 (N_4479,N_4150,N_4232);
nor U4480 (N_4480,N_4156,N_4008);
or U4481 (N_4481,N_4019,N_4218);
nand U4482 (N_4482,N_4004,N_4012);
nor U4483 (N_4483,N_4148,N_4131);
nor U4484 (N_4484,N_4000,N_4136);
xnor U4485 (N_4485,N_4049,N_4187);
xnor U4486 (N_4486,N_4071,N_4133);
nand U4487 (N_4487,N_4078,N_4083);
and U4488 (N_4488,N_4059,N_4156);
nor U4489 (N_4489,N_4021,N_4104);
nor U4490 (N_4490,N_4032,N_4241);
nand U4491 (N_4491,N_4091,N_4114);
nand U4492 (N_4492,N_4175,N_4197);
nand U4493 (N_4493,N_4075,N_4051);
and U4494 (N_4494,N_4135,N_4046);
nand U4495 (N_4495,N_4222,N_4164);
or U4496 (N_4496,N_4070,N_4028);
nand U4497 (N_4497,N_4149,N_4088);
nor U4498 (N_4498,N_4062,N_4213);
or U4499 (N_4499,N_4193,N_4245);
xnor U4500 (N_4500,N_4456,N_4417);
nand U4501 (N_4501,N_4477,N_4382);
nand U4502 (N_4502,N_4325,N_4426);
and U4503 (N_4503,N_4469,N_4364);
nand U4504 (N_4504,N_4420,N_4395);
or U4505 (N_4505,N_4479,N_4357);
or U4506 (N_4506,N_4435,N_4460);
or U4507 (N_4507,N_4307,N_4498);
and U4508 (N_4508,N_4428,N_4402);
and U4509 (N_4509,N_4371,N_4302);
xnor U4510 (N_4510,N_4271,N_4370);
xor U4511 (N_4511,N_4368,N_4401);
nor U4512 (N_4512,N_4259,N_4438);
and U4513 (N_4513,N_4481,N_4267);
xnor U4514 (N_4514,N_4335,N_4303);
xnor U4515 (N_4515,N_4390,N_4366);
nand U4516 (N_4516,N_4471,N_4377);
or U4517 (N_4517,N_4457,N_4251);
xnor U4518 (N_4518,N_4496,N_4486);
and U4519 (N_4519,N_4447,N_4403);
or U4520 (N_4520,N_4353,N_4262);
or U4521 (N_4521,N_4375,N_4332);
xnor U4522 (N_4522,N_4295,N_4491);
nand U4523 (N_4523,N_4387,N_4478);
and U4524 (N_4524,N_4425,N_4298);
nor U4525 (N_4525,N_4441,N_4328);
and U4526 (N_4526,N_4293,N_4421);
or U4527 (N_4527,N_4274,N_4299);
xnor U4528 (N_4528,N_4378,N_4288);
xor U4529 (N_4529,N_4495,N_4367);
nor U4530 (N_4530,N_4482,N_4446);
nor U4531 (N_4531,N_4424,N_4484);
nor U4532 (N_4532,N_4489,N_4392);
nor U4533 (N_4533,N_4316,N_4397);
and U4534 (N_4534,N_4338,N_4289);
nand U4535 (N_4535,N_4407,N_4343);
or U4536 (N_4536,N_4376,N_4359);
nor U4537 (N_4537,N_4297,N_4347);
or U4538 (N_4538,N_4444,N_4396);
xor U4539 (N_4539,N_4345,N_4315);
and U4540 (N_4540,N_4334,N_4344);
xor U4541 (N_4541,N_4280,N_4342);
and U4542 (N_4542,N_4459,N_4453);
nor U4543 (N_4543,N_4494,N_4388);
or U4544 (N_4544,N_4306,N_4410);
and U4545 (N_4545,N_4451,N_4254);
xnor U4546 (N_4546,N_4458,N_4252);
xor U4547 (N_4547,N_4304,N_4399);
nor U4548 (N_4548,N_4432,N_4260);
and U4549 (N_4549,N_4331,N_4309);
xnor U4550 (N_4550,N_4406,N_4348);
and U4551 (N_4551,N_4337,N_4433);
nor U4552 (N_4552,N_4250,N_4419);
or U4553 (N_4553,N_4487,N_4430);
nor U4554 (N_4554,N_4291,N_4281);
or U4555 (N_4555,N_4330,N_4270);
nand U4556 (N_4556,N_4266,N_4324);
nand U4557 (N_4557,N_4386,N_4400);
or U4558 (N_4558,N_4286,N_4322);
and U4559 (N_4559,N_4414,N_4422);
nor U4560 (N_4560,N_4379,N_4372);
and U4561 (N_4561,N_4365,N_4312);
nand U4562 (N_4562,N_4314,N_4300);
and U4563 (N_4563,N_4283,N_4265);
xnor U4564 (N_4564,N_4340,N_4268);
or U4565 (N_4565,N_4323,N_4415);
xnor U4566 (N_4566,N_4409,N_4470);
nand U4567 (N_4567,N_4360,N_4462);
xor U4568 (N_4568,N_4336,N_4255);
and U4569 (N_4569,N_4448,N_4354);
or U4570 (N_4570,N_4294,N_4427);
nand U4571 (N_4571,N_4256,N_4463);
nand U4572 (N_4572,N_4391,N_4355);
nand U4573 (N_4573,N_4356,N_4321);
nor U4574 (N_4574,N_4464,N_4490);
nor U4575 (N_4575,N_4454,N_4461);
xnor U4576 (N_4576,N_4389,N_4499);
or U4577 (N_4577,N_4341,N_4276);
nand U4578 (N_4578,N_4290,N_4319);
nand U4579 (N_4579,N_4466,N_4318);
or U4580 (N_4580,N_4442,N_4416);
nor U4581 (N_4581,N_4257,N_4326);
or U4582 (N_4582,N_4277,N_4253);
xnor U4583 (N_4583,N_4349,N_4369);
xnor U4584 (N_4584,N_4445,N_4404);
and U4585 (N_4585,N_4275,N_4339);
nand U4586 (N_4586,N_4394,N_4362);
nand U4587 (N_4587,N_4320,N_4380);
and U4588 (N_4588,N_4310,N_4385);
nand U4589 (N_4589,N_4273,N_4434);
or U4590 (N_4590,N_4405,N_4363);
nand U4591 (N_4591,N_4439,N_4413);
and U4592 (N_4592,N_4493,N_4258);
nand U4593 (N_4593,N_4333,N_4329);
xor U4594 (N_4594,N_4311,N_4383);
and U4595 (N_4595,N_4285,N_4450);
nor U4596 (N_4596,N_4497,N_4412);
and U4597 (N_4597,N_4488,N_4408);
and U4598 (N_4598,N_4440,N_4473);
nand U4599 (N_4599,N_4292,N_4476);
nor U4600 (N_4600,N_4346,N_4278);
xor U4601 (N_4601,N_4472,N_4296);
or U4602 (N_4602,N_4418,N_4351);
and U4603 (N_4603,N_4263,N_4452);
and U4604 (N_4604,N_4358,N_4468);
xor U4605 (N_4605,N_4465,N_4443);
and U4606 (N_4606,N_4480,N_4374);
xnor U4607 (N_4607,N_4350,N_4431);
or U4608 (N_4608,N_4361,N_4264);
nand U4609 (N_4609,N_4373,N_4384);
nor U4610 (N_4610,N_4381,N_4393);
xor U4611 (N_4611,N_4411,N_4327);
or U4612 (N_4612,N_4492,N_4429);
nand U4613 (N_4613,N_4305,N_4483);
and U4614 (N_4614,N_4301,N_4436);
and U4615 (N_4615,N_4279,N_4485);
nand U4616 (N_4616,N_4282,N_4467);
and U4617 (N_4617,N_4475,N_4449);
nor U4618 (N_4618,N_4313,N_4284);
or U4619 (N_4619,N_4398,N_4287);
or U4620 (N_4620,N_4455,N_4308);
xnor U4621 (N_4621,N_4352,N_4269);
or U4622 (N_4622,N_4474,N_4272);
nor U4623 (N_4623,N_4261,N_4423);
nand U4624 (N_4624,N_4437,N_4317);
or U4625 (N_4625,N_4287,N_4353);
nor U4626 (N_4626,N_4298,N_4276);
nand U4627 (N_4627,N_4332,N_4415);
and U4628 (N_4628,N_4355,N_4324);
and U4629 (N_4629,N_4286,N_4484);
or U4630 (N_4630,N_4293,N_4255);
and U4631 (N_4631,N_4370,N_4389);
nor U4632 (N_4632,N_4456,N_4256);
or U4633 (N_4633,N_4491,N_4255);
or U4634 (N_4634,N_4422,N_4372);
or U4635 (N_4635,N_4438,N_4433);
xor U4636 (N_4636,N_4363,N_4291);
xnor U4637 (N_4637,N_4466,N_4346);
xnor U4638 (N_4638,N_4313,N_4495);
and U4639 (N_4639,N_4297,N_4284);
and U4640 (N_4640,N_4431,N_4338);
xnor U4641 (N_4641,N_4467,N_4376);
nor U4642 (N_4642,N_4271,N_4255);
nand U4643 (N_4643,N_4486,N_4457);
or U4644 (N_4644,N_4318,N_4491);
and U4645 (N_4645,N_4453,N_4302);
nand U4646 (N_4646,N_4287,N_4264);
nand U4647 (N_4647,N_4278,N_4410);
and U4648 (N_4648,N_4264,N_4482);
nor U4649 (N_4649,N_4360,N_4378);
nor U4650 (N_4650,N_4480,N_4336);
and U4651 (N_4651,N_4416,N_4303);
and U4652 (N_4652,N_4420,N_4497);
nand U4653 (N_4653,N_4423,N_4305);
and U4654 (N_4654,N_4376,N_4289);
and U4655 (N_4655,N_4318,N_4476);
and U4656 (N_4656,N_4432,N_4368);
nand U4657 (N_4657,N_4290,N_4312);
and U4658 (N_4658,N_4467,N_4365);
and U4659 (N_4659,N_4430,N_4271);
or U4660 (N_4660,N_4309,N_4301);
or U4661 (N_4661,N_4478,N_4399);
and U4662 (N_4662,N_4447,N_4328);
nor U4663 (N_4663,N_4305,N_4480);
nor U4664 (N_4664,N_4422,N_4412);
and U4665 (N_4665,N_4451,N_4382);
and U4666 (N_4666,N_4250,N_4398);
nor U4667 (N_4667,N_4450,N_4269);
nor U4668 (N_4668,N_4280,N_4434);
and U4669 (N_4669,N_4462,N_4479);
and U4670 (N_4670,N_4339,N_4401);
or U4671 (N_4671,N_4392,N_4322);
nand U4672 (N_4672,N_4433,N_4307);
or U4673 (N_4673,N_4458,N_4401);
or U4674 (N_4674,N_4442,N_4411);
or U4675 (N_4675,N_4455,N_4336);
xor U4676 (N_4676,N_4272,N_4445);
nand U4677 (N_4677,N_4334,N_4451);
nor U4678 (N_4678,N_4371,N_4431);
nand U4679 (N_4679,N_4447,N_4474);
xnor U4680 (N_4680,N_4388,N_4267);
nand U4681 (N_4681,N_4400,N_4312);
or U4682 (N_4682,N_4293,N_4278);
and U4683 (N_4683,N_4493,N_4379);
nor U4684 (N_4684,N_4375,N_4262);
nand U4685 (N_4685,N_4331,N_4356);
and U4686 (N_4686,N_4291,N_4310);
xor U4687 (N_4687,N_4444,N_4334);
and U4688 (N_4688,N_4265,N_4475);
and U4689 (N_4689,N_4455,N_4371);
nand U4690 (N_4690,N_4342,N_4413);
nand U4691 (N_4691,N_4368,N_4385);
or U4692 (N_4692,N_4477,N_4320);
xor U4693 (N_4693,N_4409,N_4314);
nor U4694 (N_4694,N_4462,N_4429);
or U4695 (N_4695,N_4487,N_4325);
or U4696 (N_4696,N_4310,N_4492);
and U4697 (N_4697,N_4498,N_4286);
or U4698 (N_4698,N_4258,N_4464);
xnor U4699 (N_4699,N_4391,N_4260);
or U4700 (N_4700,N_4348,N_4484);
or U4701 (N_4701,N_4349,N_4321);
nor U4702 (N_4702,N_4479,N_4342);
and U4703 (N_4703,N_4421,N_4488);
xor U4704 (N_4704,N_4302,N_4273);
nor U4705 (N_4705,N_4256,N_4466);
nand U4706 (N_4706,N_4349,N_4423);
and U4707 (N_4707,N_4341,N_4289);
xnor U4708 (N_4708,N_4320,N_4427);
nand U4709 (N_4709,N_4385,N_4433);
xor U4710 (N_4710,N_4355,N_4270);
and U4711 (N_4711,N_4347,N_4432);
nand U4712 (N_4712,N_4393,N_4280);
and U4713 (N_4713,N_4490,N_4424);
xor U4714 (N_4714,N_4280,N_4294);
xnor U4715 (N_4715,N_4276,N_4287);
nand U4716 (N_4716,N_4386,N_4410);
and U4717 (N_4717,N_4253,N_4365);
and U4718 (N_4718,N_4415,N_4339);
and U4719 (N_4719,N_4344,N_4492);
and U4720 (N_4720,N_4463,N_4265);
or U4721 (N_4721,N_4253,N_4421);
nor U4722 (N_4722,N_4454,N_4301);
nor U4723 (N_4723,N_4486,N_4428);
and U4724 (N_4724,N_4365,N_4295);
xor U4725 (N_4725,N_4341,N_4400);
xor U4726 (N_4726,N_4309,N_4287);
nand U4727 (N_4727,N_4286,N_4355);
nor U4728 (N_4728,N_4309,N_4297);
and U4729 (N_4729,N_4291,N_4339);
or U4730 (N_4730,N_4270,N_4439);
and U4731 (N_4731,N_4320,N_4354);
nor U4732 (N_4732,N_4312,N_4445);
and U4733 (N_4733,N_4383,N_4252);
or U4734 (N_4734,N_4333,N_4281);
nand U4735 (N_4735,N_4386,N_4331);
and U4736 (N_4736,N_4470,N_4396);
or U4737 (N_4737,N_4429,N_4255);
nor U4738 (N_4738,N_4456,N_4491);
nor U4739 (N_4739,N_4492,N_4425);
nor U4740 (N_4740,N_4307,N_4394);
nor U4741 (N_4741,N_4377,N_4250);
nand U4742 (N_4742,N_4407,N_4398);
nor U4743 (N_4743,N_4268,N_4464);
or U4744 (N_4744,N_4413,N_4284);
nor U4745 (N_4745,N_4273,N_4482);
xnor U4746 (N_4746,N_4354,N_4344);
xor U4747 (N_4747,N_4415,N_4309);
nand U4748 (N_4748,N_4313,N_4468);
nand U4749 (N_4749,N_4498,N_4366);
and U4750 (N_4750,N_4646,N_4725);
xor U4751 (N_4751,N_4592,N_4587);
and U4752 (N_4752,N_4739,N_4690);
nand U4753 (N_4753,N_4665,N_4668);
and U4754 (N_4754,N_4595,N_4663);
nor U4755 (N_4755,N_4559,N_4673);
nand U4756 (N_4756,N_4521,N_4637);
and U4757 (N_4757,N_4659,N_4544);
nor U4758 (N_4758,N_4612,N_4580);
nand U4759 (N_4759,N_4512,N_4629);
xnor U4760 (N_4760,N_4555,N_4740);
and U4761 (N_4761,N_4604,N_4723);
nand U4762 (N_4762,N_4624,N_4609);
and U4763 (N_4763,N_4554,N_4516);
nor U4764 (N_4764,N_4603,N_4530);
nand U4765 (N_4765,N_4616,N_4669);
or U4766 (N_4766,N_4570,N_4718);
nor U4767 (N_4767,N_4531,N_4611);
and U4768 (N_4768,N_4648,N_4571);
or U4769 (N_4769,N_4707,N_4656);
nand U4770 (N_4770,N_4550,N_4613);
xnor U4771 (N_4771,N_4691,N_4503);
or U4772 (N_4772,N_4638,N_4596);
nand U4773 (N_4773,N_4749,N_4647);
nand U4774 (N_4774,N_4508,N_4532);
nand U4775 (N_4775,N_4677,N_4643);
and U4776 (N_4776,N_4676,N_4650);
nor U4777 (N_4777,N_4632,N_4682);
nand U4778 (N_4778,N_4608,N_4704);
nor U4779 (N_4779,N_4680,N_4543);
xor U4780 (N_4780,N_4526,N_4639);
nor U4781 (N_4781,N_4713,N_4698);
xnor U4782 (N_4782,N_4716,N_4664);
nor U4783 (N_4783,N_4642,N_4599);
xor U4784 (N_4784,N_4715,N_4649);
nor U4785 (N_4785,N_4699,N_4561);
nor U4786 (N_4786,N_4722,N_4567);
or U4787 (N_4787,N_4667,N_4692);
or U4788 (N_4788,N_4514,N_4625);
nand U4789 (N_4789,N_4505,N_4510);
or U4790 (N_4790,N_4600,N_4737);
xor U4791 (N_4791,N_4515,N_4672);
xnor U4792 (N_4792,N_4683,N_4535);
and U4793 (N_4793,N_4605,N_4708);
nor U4794 (N_4794,N_4689,N_4744);
xnor U4795 (N_4795,N_4651,N_4743);
nor U4796 (N_4796,N_4574,N_4547);
nand U4797 (N_4797,N_4536,N_4586);
xnor U4798 (N_4798,N_4504,N_4548);
nand U4799 (N_4799,N_4655,N_4719);
xor U4800 (N_4800,N_4614,N_4590);
or U4801 (N_4801,N_4562,N_4636);
and U4802 (N_4802,N_4720,N_4675);
or U4803 (N_4803,N_4635,N_4581);
nor U4804 (N_4804,N_4721,N_4578);
xnor U4805 (N_4805,N_4712,N_4618);
or U4806 (N_4806,N_4593,N_4585);
nor U4807 (N_4807,N_4519,N_4545);
and U4808 (N_4808,N_4674,N_4741);
xnor U4809 (N_4809,N_4588,N_4644);
and U4810 (N_4810,N_4745,N_4534);
or U4811 (N_4811,N_4686,N_4617);
or U4812 (N_4812,N_4598,N_4709);
nor U4813 (N_4813,N_4724,N_4627);
nor U4814 (N_4814,N_4634,N_4678);
nor U4815 (N_4815,N_4517,N_4540);
and U4816 (N_4816,N_4670,N_4657);
nor U4817 (N_4817,N_4524,N_4702);
and U4818 (N_4818,N_4693,N_4513);
and U4819 (N_4819,N_4735,N_4738);
and U4820 (N_4820,N_4584,N_4557);
xor U4821 (N_4821,N_4717,N_4607);
or U4822 (N_4822,N_4502,N_4660);
or U4823 (N_4823,N_4729,N_4507);
nand U4824 (N_4824,N_4703,N_4563);
and U4825 (N_4825,N_4583,N_4522);
nor U4826 (N_4826,N_4685,N_4538);
or U4827 (N_4827,N_4546,N_4658);
nor U4828 (N_4828,N_4573,N_4553);
or U4829 (N_4829,N_4734,N_4564);
or U4830 (N_4830,N_4631,N_4576);
nand U4831 (N_4831,N_4518,N_4727);
nor U4832 (N_4832,N_4623,N_4736);
nor U4833 (N_4833,N_4696,N_4528);
or U4834 (N_4834,N_4652,N_4594);
nand U4835 (N_4835,N_4633,N_4640);
and U4836 (N_4836,N_4748,N_4732);
nor U4837 (N_4837,N_4566,N_4610);
nor U4838 (N_4838,N_4577,N_4697);
and U4839 (N_4839,N_4662,N_4601);
nand U4840 (N_4840,N_4746,N_4710);
xnor U4841 (N_4841,N_4541,N_4747);
xnor U4842 (N_4842,N_4621,N_4597);
and U4843 (N_4843,N_4619,N_4591);
nand U4844 (N_4844,N_4565,N_4742);
nand U4845 (N_4845,N_4552,N_4626);
and U4846 (N_4846,N_4527,N_4681);
nand U4847 (N_4847,N_4558,N_4560);
nand U4848 (N_4848,N_4569,N_4714);
and U4849 (N_4849,N_4645,N_4706);
and U4850 (N_4850,N_4589,N_4501);
xnor U4851 (N_4851,N_4509,N_4537);
nand U4852 (N_4852,N_4622,N_4726);
nand U4853 (N_4853,N_4695,N_4511);
and U4854 (N_4854,N_4568,N_4572);
and U4855 (N_4855,N_4694,N_4641);
xor U4856 (N_4856,N_4529,N_4705);
nand U4857 (N_4857,N_4506,N_4551);
nand U4858 (N_4858,N_4575,N_4688);
xnor U4859 (N_4859,N_4602,N_4653);
nand U4860 (N_4860,N_4630,N_4701);
xnor U4861 (N_4861,N_4731,N_4556);
xnor U4862 (N_4862,N_4615,N_4500);
xor U4863 (N_4863,N_4606,N_4684);
nand U4864 (N_4864,N_4525,N_4579);
nand U4865 (N_4865,N_4549,N_4620);
nand U4866 (N_4866,N_4730,N_4666);
and U4867 (N_4867,N_4539,N_4533);
nor U4868 (N_4868,N_4523,N_4520);
xnor U4869 (N_4869,N_4542,N_4654);
xor U4870 (N_4870,N_4687,N_4711);
xnor U4871 (N_4871,N_4679,N_4628);
nor U4872 (N_4872,N_4582,N_4700);
and U4873 (N_4873,N_4728,N_4733);
nor U4874 (N_4874,N_4671,N_4661);
xor U4875 (N_4875,N_4529,N_4653);
or U4876 (N_4876,N_4745,N_4590);
nand U4877 (N_4877,N_4589,N_4626);
nor U4878 (N_4878,N_4664,N_4639);
nand U4879 (N_4879,N_4574,N_4511);
and U4880 (N_4880,N_4596,N_4578);
or U4881 (N_4881,N_4624,N_4736);
nor U4882 (N_4882,N_4708,N_4626);
nor U4883 (N_4883,N_4556,N_4734);
nor U4884 (N_4884,N_4664,N_4500);
and U4885 (N_4885,N_4731,N_4605);
or U4886 (N_4886,N_4551,N_4641);
and U4887 (N_4887,N_4660,N_4731);
nand U4888 (N_4888,N_4509,N_4517);
and U4889 (N_4889,N_4561,N_4746);
and U4890 (N_4890,N_4726,N_4579);
xor U4891 (N_4891,N_4520,N_4745);
xnor U4892 (N_4892,N_4550,N_4555);
and U4893 (N_4893,N_4597,N_4716);
and U4894 (N_4894,N_4507,N_4610);
xnor U4895 (N_4895,N_4684,N_4581);
nand U4896 (N_4896,N_4619,N_4632);
or U4897 (N_4897,N_4695,N_4518);
and U4898 (N_4898,N_4641,N_4646);
or U4899 (N_4899,N_4574,N_4715);
and U4900 (N_4900,N_4666,N_4583);
and U4901 (N_4901,N_4703,N_4646);
nand U4902 (N_4902,N_4669,N_4679);
xnor U4903 (N_4903,N_4597,N_4525);
nor U4904 (N_4904,N_4582,N_4513);
and U4905 (N_4905,N_4609,N_4679);
xor U4906 (N_4906,N_4651,N_4586);
and U4907 (N_4907,N_4708,N_4500);
xnor U4908 (N_4908,N_4719,N_4737);
nor U4909 (N_4909,N_4553,N_4580);
and U4910 (N_4910,N_4625,N_4618);
xor U4911 (N_4911,N_4611,N_4549);
nor U4912 (N_4912,N_4586,N_4613);
nand U4913 (N_4913,N_4594,N_4728);
and U4914 (N_4914,N_4648,N_4515);
and U4915 (N_4915,N_4524,N_4687);
and U4916 (N_4916,N_4553,N_4563);
and U4917 (N_4917,N_4535,N_4613);
xor U4918 (N_4918,N_4722,N_4560);
nand U4919 (N_4919,N_4587,N_4654);
nor U4920 (N_4920,N_4676,N_4572);
xor U4921 (N_4921,N_4587,N_4594);
and U4922 (N_4922,N_4707,N_4607);
xnor U4923 (N_4923,N_4602,N_4587);
nand U4924 (N_4924,N_4527,N_4505);
xor U4925 (N_4925,N_4743,N_4571);
nor U4926 (N_4926,N_4606,N_4723);
xor U4927 (N_4927,N_4651,N_4697);
or U4928 (N_4928,N_4692,N_4504);
xnor U4929 (N_4929,N_4635,N_4538);
nand U4930 (N_4930,N_4668,N_4539);
nand U4931 (N_4931,N_4523,N_4550);
and U4932 (N_4932,N_4618,N_4616);
or U4933 (N_4933,N_4664,N_4581);
xnor U4934 (N_4934,N_4623,N_4576);
or U4935 (N_4935,N_4622,N_4711);
nor U4936 (N_4936,N_4529,N_4592);
nor U4937 (N_4937,N_4707,N_4504);
or U4938 (N_4938,N_4747,N_4646);
xor U4939 (N_4939,N_4641,N_4740);
nor U4940 (N_4940,N_4690,N_4550);
or U4941 (N_4941,N_4590,N_4573);
xor U4942 (N_4942,N_4609,N_4723);
nand U4943 (N_4943,N_4608,N_4745);
and U4944 (N_4944,N_4730,N_4715);
nand U4945 (N_4945,N_4618,N_4626);
nand U4946 (N_4946,N_4537,N_4695);
nand U4947 (N_4947,N_4546,N_4710);
xor U4948 (N_4948,N_4676,N_4527);
or U4949 (N_4949,N_4606,N_4689);
or U4950 (N_4950,N_4636,N_4675);
nand U4951 (N_4951,N_4667,N_4592);
or U4952 (N_4952,N_4640,N_4539);
or U4953 (N_4953,N_4543,N_4520);
and U4954 (N_4954,N_4508,N_4574);
or U4955 (N_4955,N_4548,N_4691);
or U4956 (N_4956,N_4714,N_4530);
nor U4957 (N_4957,N_4580,N_4694);
nand U4958 (N_4958,N_4747,N_4691);
xnor U4959 (N_4959,N_4660,N_4645);
or U4960 (N_4960,N_4745,N_4566);
nand U4961 (N_4961,N_4671,N_4668);
or U4962 (N_4962,N_4718,N_4506);
nand U4963 (N_4963,N_4712,N_4525);
and U4964 (N_4964,N_4507,N_4705);
or U4965 (N_4965,N_4611,N_4628);
nor U4966 (N_4966,N_4667,N_4588);
nor U4967 (N_4967,N_4565,N_4571);
and U4968 (N_4968,N_4675,N_4589);
nand U4969 (N_4969,N_4700,N_4675);
or U4970 (N_4970,N_4670,N_4535);
xor U4971 (N_4971,N_4569,N_4549);
or U4972 (N_4972,N_4586,N_4679);
xnor U4973 (N_4973,N_4575,N_4558);
or U4974 (N_4974,N_4625,N_4574);
nand U4975 (N_4975,N_4688,N_4663);
xnor U4976 (N_4976,N_4660,N_4625);
nand U4977 (N_4977,N_4619,N_4730);
xnor U4978 (N_4978,N_4679,N_4712);
nand U4979 (N_4979,N_4738,N_4746);
and U4980 (N_4980,N_4681,N_4732);
and U4981 (N_4981,N_4725,N_4693);
xor U4982 (N_4982,N_4693,N_4574);
nand U4983 (N_4983,N_4642,N_4522);
or U4984 (N_4984,N_4637,N_4716);
nor U4985 (N_4985,N_4654,N_4729);
or U4986 (N_4986,N_4650,N_4678);
nor U4987 (N_4987,N_4708,N_4714);
xor U4988 (N_4988,N_4541,N_4658);
or U4989 (N_4989,N_4626,N_4567);
nand U4990 (N_4990,N_4543,N_4659);
xnor U4991 (N_4991,N_4718,N_4622);
xor U4992 (N_4992,N_4660,N_4679);
nand U4993 (N_4993,N_4699,N_4610);
nand U4994 (N_4994,N_4660,N_4527);
xor U4995 (N_4995,N_4637,N_4644);
and U4996 (N_4996,N_4533,N_4578);
nor U4997 (N_4997,N_4531,N_4625);
nand U4998 (N_4998,N_4705,N_4698);
nand U4999 (N_4999,N_4598,N_4674);
and U5000 (N_5000,N_4924,N_4943);
or U5001 (N_5001,N_4914,N_4971);
nand U5002 (N_5002,N_4790,N_4951);
nand U5003 (N_5003,N_4903,N_4796);
and U5004 (N_5004,N_4922,N_4909);
nor U5005 (N_5005,N_4894,N_4750);
and U5006 (N_5006,N_4807,N_4862);
and U5007 (N_5007,N_4937,N_4978);
xor U5008 (N_5008,N_4842,N_4847);
and U5009 (N_5009,N_4770,N_4848);
nor U5010 (N_5010,N_4826,N_4964);
and U5011 (N_5011,N_4830,N_4936);
nor U5012 (N_5012,N_4835,N_4858);
xnor U5013 (N_5013,N_4915,N_4899);
and U5014 (N_5014,N_4851,N_4992);
nand U5015 (N_5015,N_4892,N_4864);
and U5016 (N_5016,N_4872,N_4965);
nand U5017 (N_5017,N_4893,N_4814);
xnor U5018 (N_5018,N_4928,N_4968);
nand U5019 (N_5019,N_4753,N_4947);
nor U5020 (N_5020,N_4809,N_4788);
xnor U5021 (N_5021,N_4844,N_4787);
nor U5022 (N_5022,N_4776,N_4831);
and U5023 (N_5023,N_4785,N_4884);
xor U5024 (N_5024,N_4886,N_4925);
nand U5025 (N_5025,N_4756,N_4856);
or U5026 (N_5026,N_4885,N_4775);
or U5027 (N_5027,N_4958,N_4765);
nor U5028 (N_5028,N_4933,N_4904);
xnor U5029 (N_5029,N_4760,N_4939);
or U5030 (N_5030,N_4763,N_4876);
or U5031 (N_5031,N_4865,N_4912);
nor U5032 (N_5032,N_4952,N_4956);
and U5033 (N_5033,N_4838,N_4950);
or U5034 (N_5034,N_4993,N_4762);
or U5035 (N_5035,N_4895,N_4784);
or U5036 (N_5036,N_4970,N_4853);
or U5037 (N_5037,N_4755,N_4861);
or U5038 (N_5038,N_4857,N_4781);
nor U5039 (N_5039,N_4940,N_4832);
nand U5040 (N_5040,N_4778,N_4897);
nand U5041 (N_5041,N_4932,N_4859);
nand U5042 (N_5042,N_4877,N_4977);
nor U5043 (N_5043,N_4811,N_4946);
xor U5044 (N_5044,N_4767,N_4982);
nor U5045 (N_5045,N_4969,N_4949);
or U5046 (N_5046,N_4754,N_4772);
nor U5047 (N_5047,N_4891,N_4927);
xor U5048 (N_5048,N_4817,N_4930);
nor U5049 (N_5049,N_4955,N_4918);
or U5050 (N_5050,N_4846,N_4873);
or U5051 (N_5051,N_4855,N_4878);
xnor U5052 (N_5052,N_4988,N_4759);
xor U5053 (N_5053,N_4780,N_4828);
nand U5054 (N_5054,N_4942,N_4783);
or U5055 (N_5055,N_4866,N_4902);
or U5056 (N_5056,N_4802,N_4959);
nand U5057 (N_5057,N_4761,N_4983);
xor U5058 (N_5058,N_4883,N_4995);
and U5059 (N_5059,N_4797,N_4829);
xor U5060 (N_5060,N_4997,N_4896);
nand U5061 (N_5061,N_4908,N_4757);
nand U5062 (N_5062,N_4999,N_4870);
nor U5063 (N_5063,N_4769,N_4773);
xor U5064 (N_5064,N_4989,N_4833);
nor U5065 (N_5065,N_4813,N_4868);
or U5066 (N_5066,N_4919,N_4889);
nor U5067 (N_5067,N_4822,N_4823);
nor U5068 (N_5068,N_4898,N_4879);
xor U5069 (N_5069,N_4984,N_4843);
xor U5070 (N_5070,N_4845,N_4820);
nand U5071 (N_5071,N_4973,N_4917);
nand U5072 (N_5072,N_4808,N_4938);
and U5073 (N_5073,N_4967,N_4803);
and U5074 (N_5074,N_4966,N_4911);
nand U5075 (N_5075,N_4907,N_4852);
nor U5076 (N_5076,N_4818,N_4929);
or U5077 (N_5077,N_4800,N_4782);
nor U5078 (N_5078,N_4887,N_4985);
nor U5079 (N_5079,N_4931,N_4824);
nor U5080 (N_5080,N_4980,N_4901);
xnor U5081 (N_5081,N_4900,N_4752);
or U5082 (N_5082,N_4996,N_4766);
nor U5083 (N_5083,N_4953,N_4854);
or U5084 (N_5084,N_4841,N_4871);
xnor U5085 (N_5085,N_4906,N_4888);
and U5086 (N_5086,N_4758,N_4972);
xnor U5087 (N_5087,N_4957,N_4987);
nand U5088 (N_5088,N_4961,N_4768);
nand U5089 (N_5089,N_4990,N_4810);
or U5090 (N_5090,N_4850,N_4812);
xnor U5091 (N_5091,N_4805,N_4920);
nor U5092 (N_5092,N_4981,N_4994);
xnor U5093 (N_5093,N_4774,N_4840);
or U5094 (N_5094,N_4921,N_4934);
nand U5095 (N_5095,N_4880,N_4863);
nor U5096 (N_5096,N_4849,N_4948);
xnor U5097 (N_5097,N_4890,N_4976);
and U5098 (N_5098,N_4804,N_4792);
or U5099 (N_5099,N_4801,N_4825);
and U5100 (N_5100,N_4963,N_4764);
and U5101 (N_5101,N_4806,N_4875);
and U5102 (N_5102,N_4979,N_4923);
xnor U5103 (N_5103,N_4837,N_4819);
or U5104 (N_5104,N_4998,N_4905);
or U5105 (N_5105,N_4926,N_4834);
and U5106 (N_5106,N_4867,N_4869);
nor U5107 (N_5107,N_4882,N_4821);
xnor U5108 (N_5108,N_4779,N_4991);
nor U5109 (N_5109,N_4836,N_4935);
nor U5110 (N_5110,N_4910,N_4974);
or U5111 (N_5111,N_4799,N_4771);
nor U5112 (N_5112,N_4777,N_4786);
xnor U5113 (N_5113,N_4881,N_4874);
or U5114 (N_5114,N_4815,N_4945);
and U5115 (N_5115,N_4793,N_4798);
and U5116 (N_5116,N_4975,N_4795);
xnor U5117 (N_5117,N_4789,N_4794);
nand U5118 (N_5118,N_4954,N_4860);
nor U5119 (N_5119,N_4986,N_4960);
xnor U5120 (N_5120,N_4916,N_4941);
nand U5121 (N_5121,N_4791,N_4816);
xor U5122 (N_5122,N_4751,N_4962);
nand U5123 (N_5123,N_4827,N_4839);
or U5124 (N_5124,N_4944,N_4913);
xnor U5125 (N_5125,N_4772,N_4786);
and U5126 (N_5126,N_4760,N_4872);
nand U5127 (N_5127,N_4793,N_4848);
and U5128 (N_5128,N_4968,N_4916);
or U5129 (N_5129,N_4913,N_4899);
nor U5130 (N_5130,N_4960,N_4758);
and U5131 (N_5131,N_4832,N_4967);
and U5132 (N_5132,N_4976,N_4871);
xnor U5133 (N_5133,N_4775,N_4919);
nor U5134 (N_5134,N_4936,N_4809);
xor U5135 (N_5135,N_4779,N_4811);
nor U5136 (N_5136,N_4999,N_4761);
or U5137 (N_5137,N_4755,N_4805);
xor U5138 (N_5138,N_4891,N_4852);
nor U5139 (N_5139,N_4972,N_4766);
nand U5140 (N_5140,N_4918,N_4875);
nor U5141 (N_5141,N_4981,N_4926);
or U5142 (N_5142,N_4954,N_4912);
xor U5143 (N_5143,N_4918,N_4967);
or U5144 (N_5144,N_4846,N_4757);
nor U5145 (N_5145,N_4821,N_4878);
nand U5146 (N_5146,N_4758,N_4898);
and U5147 (N_5147,N_4891,N_4779);
and U5148 (N_5148,N_4799,N_4832);
nand U5149 (N_5149,N_4887,N_4910);
nand U5150 (N_5150,N_4851,N_4763);
xor U5151 (N_5151,N_4781,N_4776);
xor U5152 (N_5152,N_4761,N_4780);
nor U5153 (N_5153,N_4978,N_4848);
or U5154 (N_5154,N_4758,N_4788);
nor U5155 (N_5155,N_4799,N_4972);
and U5156 (N_5156,N_4760,N_4837);
nor U5157 (N_5157,N_4750,N_4965);
nand U5158 (N_5158,N_4979,N_4838);
nor U5159 (N_5159,N_4924,N_4982);
xnor U5160 (N_5160,N_4818,N_4766);
xor U5161 (N_5161,N_4757,N_4811);
and U5162 (N_5162,N_4843,N_4991);
xnor U5163 (N_5163,N_4927,N_4984);
nand U5164 (N_5164,N_4818,N_4776);
and U5165 (N_5165,N_4976,N_4791);
and U5166 (N_5166,N_4786,N_4788);
xnor U5167 (N_5167,N_4882,N_4950);
or U5168 (N_5168,N_4762,N_4984);
xor U5169 (N_5169,N_4864,N_4975);
or U5170 (N_5170,N_4975,N_4981);
nand U5171 (N_5171,N_4909,N_4910);
nor U5172 (N_5172,N_4776,N_4941);
nand U5173 (N_5173,N_4841,N_4867);
nand U5174 (N_5174,N_4879,N_4998);
nand U5175 (N_5175,N_4995,N_4865);
xor U5176 (N_5176,N_4862,N_4990);
nor U5177 (N_5177,N_4995,N_4857);
or U5178 (N_5178,N_4934,N_4750);
nor U5179 (N_5179,N_4953,N_4899);
nand U5180 (N_5180,N_4980,N_4767);
and U5181 (N_5181,N_4750,N_4819);
nor U5182 (N_5182,N_4965,N_4875);
nor U5183 (N_5183,N_4979,N_4821);
nor U5184 (N_5184,N_4901,N_4757);
or U5185 (N_5185,N_4834,N_4974);
nor U5186 (N_5186,N_4935,N_4850);
nor U5187 (N_5187,N_4750,N_4915);
and U5188 (N_5188,N_4860,N_4816);
xnor U5189 (N_5189,N_4903,N_4752);
nor U5190 (N_5190,N_4780,N_4850);
xnor U5191 (N_5191,N_4786,N_4879);
xor U5192 (N_5192,N_4906,N_4757);
nand U5193 (N_5193,N_4816,N_4978);
nor U5194 (N_5194,N_4828,N_4961);
and U5195 (N_5195,N_4915,N_4950);
nand U5196 (N_5196,N_4965,N_4861);
or U5197 (N_5197,N_4860,N_4793);
and U5198 (N_5198,N_4785,N_4928);
xnor U5199 (N_5199,N_4873,N_4971);
xnor U5200 (N_5200,N_4947,N_4751);
and U5201 (N_5201,N_4788,N_4852);
nand U5202 (N_5202,N_4839,N_4786);
nor U5203 (N_5203,N_4949,N_4925);
and U5204 (N_5204,N_4936,N_4851);
or U5205 (N_5205,N_4962,N_4874);
xor U5206 (N_5206,N_4995,N_4967);
nand U5207 (N_5207,N_4825,N_4917);
and U5208 (N_5208,N_4845,N_4759);
or U5209 (N_5209,N_4953,N_4817);
nand U5210 (N_5210,N_4759,N_4827);
or U5211 (N_5211,N_4805,N_4931);
and U5212 (N_5212,N_4815,N_4809);
nor U5213 (N_5213,N_4863,N_4900);
nand U5214 (N_5214,N_4862,N_4984);
nor U5215 (N_5215,N_4935,N_4875);
and U5216 (N_5216,N_4919,N_4886);
xnor U5217 (N_5217,N_4868,N_4992);
nor U5218 (N_5218,N_4900,N_4834);
or U5219 (N_5219,N_4819,N_4958);
xor U5220 (N_5220,N_4952,N_4858);
and U5221 (N_5221,N_4901,N_4987);
nand U5222 (N_5222,N_4765,N_4942);
or U5223 (N_5223,N_4925,N_4960);
or U5224 (N_5224,N_4903,N_4850);
nor U5225 (N_5225,N_4877,N_4997);
xor U5226 (N_5226,N_4964,N_4959);
nand U5227 (N_5227,N_4880,N_4761);
and U5228 (N_5228,N_4919,N_4812);
xnor U5229 (N_5229,N_4919,N_4921);
or U5230 (N_5230,N_4761,N_4907);
or U5231 (N_5231,N_4834,N_4998);
nor U5232 (N_5232,N_4839,N_4798);
nor U5233 (N_5233,N_4796,N_4870);
and U5234 (N_5234,N_4783,N_4951);
and U5235 (N_5235,N_4973,N_4959);
nor U5236 (N_5236,N_4957,N_4965);
and U5237 (N_5237,N_4802,N_4957);
nand U5238 (N_5238,N_4780,N_4995);
nor U5239 (N_5239,N_4984,N_4853);
or U5240 (N_5240,N_4775,N_4848);
or U5241 (N_5241,N_4971,N_4848);
xor U5242 (N_5242,N_4853,N_4763);
and U5243 (N_5243,N_4882,N_4835);
xor U5244 (N_5244,N_4910,N_4864);
nor U5245 (N_5245,N_4795,N_4849);
nor U5246 (N_5246,N_4815,N_4912);
nor U5247 (N_5247,N_4994,N_4966);
or U5248 (N_5248,N_4840,N_4996);
nand U5249 (N_5249,N_4771,N_4780);
nand U5250 (N_5250,N_5109,N_5030);
or U5251 (N_5251,N_5159,N_5057);
or U5252 (N_5252,N_5234,N_5189);
nor U5253 (N_5253,N_5184,N_5138);
nand U5254 (N_5254,N_5064,N_5041);
nand U5255 (N_5255,N_5087,N_5187);
xor U5256 (N_5256,N_5073,N_5160);
nor U5257 (N_5257,N_5246,N_5106);
nor U5258 (N_5258,N_5089,N_5132);
and U5259 (N_5259,N_5185,N_5112);
xnor U5260 (N_5260,N_5009,N_5034);
nor U5261 (N_5261,N_5179,N_5026);
xnor U5262 (N_5262,N_5149,N_5228);
nand U5263 (N_5263,N_5051,N_5152);
nand U5264 (N_5264,N_5125,N_5216);
nor U5265 (N_5265,N_5163,N_5061);
xor U5266 (N_5266,N_5151,N_5053);
xor U5267 (N_5267,N_5186,N_5209);
nand U5268 (N_5268,N_5119,N_5081);
nor U5269 (N_5269,N_5094,N_5108);
nand U5270 (N_5270,N_5215,N_5050);
xnor U5271 (N_5271,N_5102,N_5084);
and U5272 (N_5272,N_5178,N_5023);
or U5273 (N_5273,N_5117,N_5122);
and U5274 (N_5274,N_5223,N_5201);
or U5275 (N_5275,N_5193,N_5227);
xor U5276 (N_5276,N_5166,N_5110);
xnor U5277 (N_5277,N_5194,N_5036);
nand U5278 (N_5278,N_5222,N_5180);
or U5279 (N_5279,N_5033,N_5190);
xor U5280 (N_5280,N_5200,N_5097);
nand U5281 (N_5281,N_5062,N_5044);
nor U5282 (N_5282,N_5143,N_5188);
or U5283 (N_5283,N_5226,N_5249);
and U5284 (N_5284,N_5065,N_5150);
xor U5285 (N_5285,N_5075,N_5177);
and U5286 (N_5286,N_5017,N_5091);
nand U5287 (N_5287,N_5114,N_5131);
xnor U5288 (N_5288,N_5086,N_5219);
xor U5289 (N_5289,N_5220,N_5020);
and U5290 (N_5290,N_5213,N_5191);
nand U5291 (N_5291,N_5165,N_5146);
xor U5292 (N_5292,N_5205,N_5211);
and U5293 (N_5293,N_5028,N_5148);
or U5294 (N_5294,N_5043,N_5123);
and U5295 (N_5295,N_5092,N_5074);
nand U5296 (N_5296,N_5248,N_5105);
and U5297 (N_5297,N_5042,N_5140);
nor U5298 (N_5298,N_5083,N_5046);
or U5299 (N_5299,N_5098,N_5198);
nand U5300 (N_5300,N_5101,N_5022);
or U5301 (N_5301,N_5055,N_5129);
and U5302 (N_5302,N_5155,N_5002);
xnor U5303 (N_5303,N_5170,N_5208);
and U5304 (N_5304,N_5134,N_5144);
nor U5305 (N_5305,N_5124,N_5142);
and U5306 (N_5306,N_5004,N_5233);
nor U5307 (N_5307,N_5225,N_5118);
nor U5308 (N_5308,N_5076,N_5013);
xnor U5309 (N_5309,N_5052,N_5007);
nand U5310 (N_5310,N_5058,N_5231);
xor U5311 (N_5311,N_5095,N_5192);
nor U5312 (N_5312,N_5011,N_5162);
nor U5313 (N_5313,N_5049,N_5016);
xor U5314 (N_5314,N_5217,N_5136);
xnor U5315 (N_5315,N_5199,N_5090);
or U5316 (N_5316,N_5048,N_5203);
nor U5317 (N_5317,N_5128,N_5060);
and U5318 (N_5318,N_5172,N_5072);
and U5319 (N_5319,N_5088,N_5247);
nor U5320 (N_5320,N_5175,N_5082);
and U5321 (N_5321,N_5054,N_5196);
xnor U5322 (N_5322,N_5229,N_5113);
nand U5323 (N_5323,N_5232,N_5242);
and U5324 (N_5324,N_5243,N_5080);
nor U5325 (N_5325,N_5068,N_5182);
or U5326 (N_5326,N_5018,N_5099);
nand U5327 (N_5327,N_5156,N_5014);
nor U5328 (N_5328,N_5130,N_5063);
and U5329 (N_5329,N_5210,N_5005);
nor U5330 (N_5330,N_5221,N_5010);
nand U5331 (N_5331,N_5167,N_5207);
and U5332 (N_5332,N_5212,N_5157);
nand U5333 (N_5333,N_5107,N_5224);
nor U5334 (N_5334,N_5104,N_5169);
nor U5335 (N_5335,N_5015,N_5093);
xor U5336 (N_5336,N_5003,N_5111);
xnor U5337 (N_5337,N_5120,N_5218);
and U5338 (N_5338,N_5145,N_5241);
nand U5339 (N_5339,N_5079,N_5066);
and U5340 (N_5340,N_5040,N_5085);
or U5341 (N_5341,N_5100,N_5206);
and U5342 (N_5342,N_5059,N_5176);
xor U5343 (N_5343,N_5027,N_5230);
and U5344 (N_5344,N_5025,N_5147);
nand U5345 (N_5345,N_5133,N_5038);
nor U5346 (N_5346,N_5245,N_5235);
or U5347 (N_5347,N_5158,N_5244);
and U5348 (N_5348,N_5067,N_5071);
nor U5349 (N_5349,N_5197,N_5045);
xor U5350 (N_5350,N_5135,N_5056);
and U5351 (N_5351,N_5153,N_5037);
xor U5352 (N_5352,N_5039,N_5238);
or U5353 (N_5353,N_5126,N_5001);
and U5354 (N_5354,N_5171,N_5021);
xnor U5355 (N_5355,N_5006,N_5183);
and U5356 (N_5356,N_5174,N_5202);
nor U5357 (N_5357,N_5103,N_5195);
nand U5358 (N_5358,N_5164,N_5141);
or U5359 (N_5359,N_5173,N_5029);
or U5360 (N_5360,N_5127,N_5239);
xor U5361 (N_5361,N_5237,N_5115);
nand U5362 (N_5362,N_5070,N_5121);
nand U5363 (N_5363,N_5032,N_5137);
nand U5364 (N_5364,N_5008,N_5078);
xor U5365 (N_5365,N_5116,N_5236);
nor U5366 (N_5366,N_5069,N_5181);
nor U5367 (N_5367,N_5154,N_5047);
nor U5368 (N_5368,N_5096,N_5240);
or U5369 (N_5369,N_5204,N_5012);
nor U5370 (N_5370,N_5024,N_5077);
nor U5371 (N_5371,N_5168,N_5031);
nand U5372 (N_5372,N_5019,N_5161);
or U5373 (N_5373,N_5214,N_5139);
nand U5374 (N_5374,N_5000,N_5035);
nand U5375 (N_5375,N_5047,N_5000);
xor U5376 (N_5376,N_5122,N_5142);
xor U5377 (N_5377,N_5147,N_5162);
nor U5378 (N_5378,N_5246,N_5198);
nor U5379 (N_5379,N_5023,N_5012);
xor U5380 (N_5380,N_5050,N_5240);
and U5381 (N_5381,N_5175,N_5056);
or U5382 (N_5382,N_5162,N_5158);
nand U5383 (N_5383,N_5124,N_5010);
xnor U5384 (N_5384,N_5224,N_5133);
and U5385 (N_5385,N_5245,N_5002);
xnor U5386 (N_5386,N_5163,N_5216);
xnor U5387 (N_5387,N_5162,N_5144);
and U5388 (N_5388,N_5217,N_5102);
xnor U5389 (N_5389,N_5144,N_5059);
or U5390 (N_5390,N_5003,N_5107);
xnor U5391 (N_5391,N_5191,N_5139);
xor U5392 (N_5392,N_5032,N_5089);
nand U5393 (N_5393,N_5061,N_5140);
and U5394 (N_5394,N_5187,N_5205);
xnor U5395 (N_5395,N_5114,N_5032);
nor U5396 (N_5396,N_5168,N_5071);
nand U5397 (N_5397,N_5161,N_5150);
nor U5398 (N_5398,N_5183,N_5207);
or U5399 (N_5399,N_5248,N_5173);
and U5400 (N_5400,N_5147,N_5165);
nand U5401 (N_5401,N_5019,N_5102);
xor U5402 (N_5402,N_5248,N_5030);
and U5403 (N_5403,N_5146,N_5224);
nor U5404 (N_5404,N_5198,N_5021);
and U5405 (N_5405,N_5196,N_5145);
xnor U5406 (N_5406,N_5096,N_5114);
nand U5407 (N_5407,N_5222,N_5229);
or U5408 (N_5408,N_5227,N_5163);
and U5409 (N_5409,N_5235,N_5141);
xor U5410 (N_5410,N_5143,N_5136);
xnor U5411 (N_5411,N_5061,N_5101);
nor U5412 (N_5412,N_5091,N_5185);
and U5413 (N_5413,N_5059,N_5218);
nand U5414 (N_5414,N_5182,N_5102);
or U5415 (N_5415,N_5239,N_5124);
nand U5416 (N_5416,N_5140,N_5144);
nand U5417 (N_5417,N_5221,N_5162);
xnor U5418 (N_5418,N_5089,N_5156);
nand U5419 (N_5419,N_5234,N_5181);
nand U5420 (N_5420,N_5034,N_5067);
or U5421 (N_5421,N_5245,N_5188);
and U5422 (N_5422,N_5001,N_5190);
nand U5423 (N_5423,N_5130,N_5178);
or U5424 (N_5424,N_5228,N_5182);
and U5425 (N_5425,N_5203,N_5121);
nand U5426 (N_5426,N_5042,N_5073);
or U5427 (N_5427,N_5185,N_5183);
xnor U5428 (N_5428,N_5191,N_5138);
nor U5429 (N_5429,N_5024,N_5144);
xor U5430 (N_5430,N_5091,N_5071);
nor U5431 (N_5431,N_5101,N_5074);
nand U5432 (N_5432,N_5222,N_5047);
or U5433 (N_5433,N_5138,N_5050);
and U5434 (N_5434,N_5242,N_5003);
xor U5435 (N_5435,N_5014,N_5010);
nand U5436 (N_5436,N_5120,N_5142);
xor U5437 (N_5437,N_5182,N_5237);
nor U5438 (N_5438,N_5205,N_5063);
nand U5439 (N_5439,N_5211,N_5016);
and U5440 (N_5440,N_5058,N_5038);
and U5441 (N_5441,N_5190,N_5135);
nand U5442 (N_5442,N_5009,N_5177);
nor U5443 (N_5443,N_5099,N_5065);
and U5444 (N_5444,N_5188,N_5039);
nand U5445 (N_5445,N_5131,N_5074);
xor U5446 (N_5446,N_5165,N_5068);
nand U5447 (N_5447,N_5228,N_5238);
nand U5448 (N_5448,N_5240,N_5051);
xnor U5449 (N_5449,N_5053,N_5134);
nand U5450 (N_5450,N_5242,N_5104);
nand U5451 (N_5451,N_5050,N_5180);
xnor U5452 (N_5452,N_5126,N_5089);
and U5453 (N_5453,N_5110,N_5189);
nor U5454 (N_5454,N_5030,N_5217);
nand U5455 (N_5455,N_5158,N_5064);
nand U5456 (N_5456,N_5190,N_5049);
or U5457 (N_5457,N_5132,N_5068);
and U5458 (N_5458,N_5063,N_5084);
or U5459 (N_5459,N_5040,N_5069);
xnor U5460 (N_5460,N_5145,N_5005);
or U5461 (N_5461,N_5059,N_5159);
or U5462 (N_5462,N_5072,N_5074);
nor U5463 (N_5463,N_5242,N_5135);
xor U5464 (N_5464,N_5216,N_5104);
nor U5465 (N_5465,N_5107,N_5193);
xor U5466 (N_5466,N_5125,N_5016);
nand U5467 (N_5467,N_5076,N_5199);
nor U5468 (N_5468,N_5168,N_5104);
xnor U5469 (N_5469,N_5198,N_5147);
xnor U5470 (N_5470,N_5161,N_5048);
and U5471 (N_5471,N_5056,N_5032);
or U5472 (N_5472,N_5179,N_5045);
nand U5473 (N_5473,N_5035,N_5108);
or U5474 (N_5474,N_5111,N_5088);
or U5475 (N_5475,N_5064,N_5066);
or U5476 (N_5476,N_5186,N_5242);
xnor U5477 (N_5477,N_5114,N_5150);
and U5478 (N_5478,N_5155,N_5222);
or U5479 (N_5479,N_5238,N_5011);
nor U5480 (N_5480,N_5112,N_5062);
xnor U5481 (N_5481,N_5003,N_5051);
and U5482 (N_5482,N_5149,N_5232);
nand U5483 (N_5483,N_5009,N_5210);
and U5484 (N_5484,N_5176,N_5209);
or U5485 (N_5485,N_5229,N_5100);
nand U5486 (N_5486,N_5066,N_5018);
nor U5487 (N_5487,N_5095,N_5093);
nor U5488 (N_5488,N_5095,N_5127);
or U5489 (N_5489,N_5036,N_5065);
and U5490 (N_5490,N_5179,N_5248);
or U5491 (N_5491,N_5092,N_5008);
nor U5492 (N_5492,N_5143,N_5116);
nor U5493 (N_5493,N_5019,N_5205);
xnor U5494 (N_5494,N_5046,N_5222);
nand U5495 (N_5495,N_5142,N_5048);
nor U5496 (N_5496,N_5237,N_5045);
nor U5497 (N_5497,N_5244,N_5023);
or U5498 (N_5498,N_5194,N_5126);
or U5499 (N_5499,N_5085,N_5067);
nand U5500 (N_5500,N_5432,N_5324);
or U5501 (N_5501,N_5404,N_5300);
or U5502 (N_5502,N_5344,N_5463);
nand U5503 (N_5503,N_5414,N_5423);
xor U5504 (N_5504,N_5489,N_5455);
xnor U5505 (N_5505,N_5498,N_5292);
xor U5506 (N_5506,N_5367,N_5488);
nor U5507 (N_5507,N_5269,N_5296);
and U5508 (N_5508,N_5291,N_5471);
and U5509 (N_5509,N_5415,N_5469);
and U5510 (N_5510,N_5263,N_5381);
or U5511 (N_5511,N_5451,N_5456);
and U5512 (N_5512,N_5407,N_5287);
nand U5513 (N_5513,N_5478,N_5363);
xor U5514 (N_5514,N_5319,N_5290);
nand U5515 (N_5515,N_5312,N_5316);
nor U5516 (N_5516,N_5295,N_5412);
and U5517 (N_5517,N_5462,N_5443);
and U5518 (N_5518,N_5356,N_5258);
or U5519 (N_5519,N_5399,N_5409);
and U5520 (N_5520,N_5476,N_5271);
or U5521 (N_5521,N_5400,N_5314);
or U5522 (N_5522,N_5477,N_5354);
nor U5523 (N_5523,N_5441,N_5482);
and U5524 (N_5524,N_5307,N_5388);
and U5525 (N_5525,N_5332,N_5440);
or U5526 (N_5526,N_5322,N_5436);
nand U5527 (N_5527,N_5346,N_5361);
nand U5528 (N_5528,N_5416,N_5475);
and U5529 (N_5529,N_5311,N_5438);
or U5530 (N_5530,N_5470,N_5317);
or U5531 (N_5531,N_5250,N_5278);
or U5532 (N_5532,N_5283,N_5386);
and U5533 (N_5533,N_5329,N_5347);
or U5534 (N_5534,N_5277,N_5282);
and U5535 (N_5535,N_5398,N_5351);
xnor U5536 (N_5536,N_5293,N_5431);
or U5537 (N_5537,N_5371,N_5421);
nand U5538 (N_5538,N_5288,N_5392);
xnor U5539 (N_5539,N_5397,N_5357);
nor U5540 (N_5540,N_5497,N_5486);
and U5541 (N_5541,N_5362,N_5474);
and U5542 (N_5542,N_5370,N_5430);
xnor U5543 (N_5543,N_5256,N_5484);
nand U5544 (N_5544,N_5480,N_5457);
nand U5545 (N_5545,N_5483,N_5402);
or U5546 (N_5546,N_5369,N_5270);
nand U5547 (N_5547,N_5289,N_5259);
or U5548 (N_5548,N_5377,N_5396);
nor U5549 (N_5549,N_5422,N_5275);
and U5550 (N_5550,N_5395,N_5366);
xor U5551 (N_5551,N_5403,N_5360);
nand U5552 (N_5552,N_5251,N_5389);
xnor U5553 (N_5553,N_5331,N_5375);
xor U5554 (N_5554,N_5336,N_5445);
xor U5555 (N_5555,N_5461,N_5450);
xnor U5556 (N_5556,N_5447,N_5297);
and U5557 (N_5557,N_5301,N_5434);
nor U5558 (N_5558,N_5350,N_5303);
and U5559 (N_5559,N_5429,N_5338);
and U5560 (N_5560,N_5328,N_5424);
and U5561 (N_5561,N_5284,N_5299);
and U5562 (N_5562,N_5453,N_5320);
nor U5563 (N_5563,N_5254,N_5279);
nand U5564 (N_5564,N_5267,N_5379);
nand U5565 (N_5565,N_5257,N_5365);
nor U5566 (N_5566,N_5264,N_5262);
nor U5567 (N_5567,N_5401,N_5458);
xor U5568 (N_5568,N_5349,N_5466);
nor U5569 (N_5569,N_5353,N_5417);
nand U5570 (N_5570,N_5425,N_5376);
and U5571 (N_5571,N_5446,N_5352);
nor U5572 (N_5572,N_5286,N_5408);
xnor U5573 (N_5573,N_5487,N_5339);
nor U5574 (N_5574,N_5368,N_5494);
xnor U5575 (N_5575,N_5285,N_5315);
xnor U5576 (N_5576,N_5437,N_5467);
nor U5577 (N_5577,N_5490,N_5473);
nor U5578 (N_5578,N_5495,N_5280);
or U5579 (N_5579,N_5444,N_5406);
nor U5580 (N_5580,N_5413,N_5493);
nor U5581 (N_5581,N_5266,N_5492);
nor U5582 (N_5582,N_5449,N_5298);
nand U5583 (N_5583,N_5454,N_5309);
nand U5584 (N_5584,N_5318,N_5428);
xor U5585 (N_5585,N_5372,N_5378);
and U5586 (N_5586,N_5394,N_5265);
nor U5587 (N_5587,N_5333,N_5260);
or U5588 (N_5588,N_5281,N_5439);
nand U5589 (N_5589,N_5334,N_5253);
or U5590 (N_5590,N_5335,N_5464);
and U5591 (N_5591,N_5459,N_5383);
or U5592 (N_5592,N_5405,N_5273);
or U5593 (N_5593,N_5419,N_5433);
nor U5594 (N_5594,N_5330,N_5341);
xor U5595 (N_5595,N_5355,N_5325);
nand U5596 (N_5596,N_5442,N_5435);
nand U5597 (N_5597,N_5268,N_5321);
xor U5598 (N_5598,N_5420,N_5418);
nor U5599 (N_5599,N_5343,N_5364);
and U5600 (N_5600,N_5272,N_5472);
xnor U5601 (N_5601,N_5340,N_5382);
xnor U5602 (N_5602,N_5306,N_5261);
nand U5603 (N_5603,N_5323,N_5374);
and U5604 (N_5604,N_5491,N_5387);
xor U5605 (N_5605,N_5385,N_5479);
and U5606 (N_5606,N_5305,N_5499);
xnor U5607 (N_5607,N_5380,N_5410);
nor U5608 (N_5608,N_5481,N_5342);
or U5609 (N_5609,N_5448,N_5390);
or U5610 (N_5610,N_5411,N_5302);
xor U5611 (N_5611,N_5373,N_5384);
nor U5612 (N_5612,N_5465,N_5313);
or U5613 (N_5613,N_5252,N_5327);
nand U5614 (N_5614,N_5304,N_5294);
nor U5615 (N_5615,N_5359,N_5427);
or U5616 (N_5616,N_5337,N_5468);
nand U5617 (N_5617,N_5393,N_5358);
or U5618 (N_5618,N_5485,N_5348);
or U5619 (N_5619,N_5452,N_5496);
and U5620 (N_5620,N_5276,N_5255);
or U5621 (N_5621,N_5391,N_5310);
xnor U5622 (N_5622,N_5345,N_5308);
xnor U5623 (N_5623,N_5426,N_5326);
or U5624 (N_5624,N_5460,N_5274);
nor U5625 (N_5625,N_5440,N_5413);
nor U5626 (N_5626,N_5433,N_5420);
xnor U5627 (N_5627,N_5495,N_5492);
nand U5628 (N_5628,N_5390,N_5322);
or U5629 (N_5629,N_5498,N_5321);
or U5630 (N_5630,N_5438,N_5495);
and U5631 (N_5631,N_5396,N_5434);
xnor U5632 (N_5632,N_5440,N_5481);
nand U5633 (N_5633,N_5312,N_5309);
nor U5634 (N_5634,N_5460,N_5473);
and U5635 (N_5635,N_5258,N_5325);
nand U5636 (N_5636,N_5319,N_5335);
xnor U5637 (N_5637,N_5486,N_5351);
nand U5638 (N_5638,N_5443,N_5422);
xor U5639 (N_5639,N_5475,N_5303);
nand U5640 (N_5640,N_5333,N_5262);
or U5641 (N_5641,N_5276,N_5391);
xor U5642 (N_5642,N_5376,N_5337);
xor U5643 (N_5643,N_5425,N_5256);
and U5644 (N_5644,N_5286,N_5342);
nand U5645 (N_5645,N_5257,N_5373);
or U5646 (N_5646,N_5372,N_5298);
nand U5647 (N_5647,N_5349,N_5493);
nand U5648 (N_5648,N_5453,N_5464);
xor U5649 (N_5649,N_5311,N_5316);
or U5650 (N_5650,N_5295,N_5311);
nand U5651 (N_5651,N_5264,N_5437);
nand U5652 (N_5652,N_5373,N_5288);
and U5653 (N_5653,N_5342,N_5470);
nor U5654 (N_5654,N_5292,N_5374);
or U5655 (N_5655,N_5314,N_5497);
or U5656 (N_5656,N_5295,N_5340);
nor U5657 (N_5657,N_5458,N_5351);
xor U5658 (N_5658,N_5410,N_5467);
xor U5659 (N_5659,N_5347,N_5309);
and U5660 (N_5660,N_5483,N_5362);
and U5661 (N_5661,N_5297,N_5336);
nor U5662 (N_5662,N_5435,N_5292);
nor U5663 (N_5663,N_5286,N_5411);
or U5664 (N_5664,N_5286,N_5387);
nor U5665 (N_5665,N_5320,N_5389);
and U5666 (N_5666,N_5291,N_5465);
nor U5667 (N_5667,N_5434,N_5304);
xor U5668 (N_5668,N_5305,N_5326);
nor U5669 (N_5669,N_5417,N_5456);
and U5670 (N_5670,N_5332,N_5403);
and U5671 (N_5671,N_5488,N_5252);
and U5672 (N_5672,N_5430,N_5267);
and U5673 (N_5673,N_5403,N_5280);
xor U5674 (N_5674,N_5397,N_5371);
and U5675 (N_5675,N_5322,N_5369);
or U5676 (N_5676,N_5430,N_5306);
or U5677 (N_5677,N_5372,N_5266);
nand U5678 (N_5678,N_5250,N_5421);
xnor U5679 (N_5679,N_5288,N_5267);
and U5680 (N_5680,N_5418,N_5483);
nand U5681 (N_5681,N_5343,N_5496);
nor U5682 (N_5682,N_5426,N_5352);
nor U5683 (N_5683,N_5305,N_5417);
nand U5684 (N_5684,N_5478,N_5295);
nand U5685 (N_5685,N_5485,N_5496);
nor U5686 (N_5686,N_5276,N_5359);
xnor U5687 (N_5687,N_5393,N_5460);
nor U5688 (N_5688,N_5263,N_5408);
xor U5689 (N_5689,N_5369,N_5289);
or U5690 (N_5690,N_5443,N_5499);
nand U5691 (N_5691,N_5475,N_5492);
or U5692 (N_5692,N_5385,N_5364);
nand U5693 (N_5693,N_5298,N_5368);
nor U5694 (N_5694,N_5328,N_5288);
or U5695 (N_5695,N_5469,N_5377);
nor U5696 (N_5696,N_5295,N_5377);
nand U5697 (N_5697,N_5345,N_5449);
or U5698 (N_5698,N_5431,N_5477);
nand U5699 (N_5699,N_5305,N_5475);
and U5700 (N_5700,N_5356,N_5399);
nor U5701 (N_5701,N_5439,N_5452);
nand U5702 (N_5702,N_5391,N_5279);
xor U5703 (N_5703,N_5279,N_5418);
nand U5704 (N_5704,N_5442,N_5342);
xnor U5705 (N_5705,N_5345,N_5378);
nor U5706 (N_5706,N_5336,N_5479);
nand U5707 (N_5707,N_5339,N_5480);
nor U5708 (N_5708,N_5377,N_5432);
or U5709 (N_5709,N_5258,N_5471);
nor U5710 (N_5710,N_5444,N_5409);
nor U5711 (N_5711,N_5345,N_5491);
and U5712 (N_5712,N_5398,N_5448);
and U5713 (N_5713,N_5462,N_5488);
nor U5714 (N_5714,N_5339,N_5271);
or U5715 (N_5715,N_5335,N_5337);
xnor U5716 (N_5716,N_5387,N_5461);
or U5717 (N_5717,N_5398,N_5429);
nor U5718 (N_5718,N_5472,N_5365);
nor U5719 (N_5719,N_5442,N_5474);
nand U5720 (N_5720,N_5265,N_5466);
nand U5721 (N_5721,N_5412,N_5372);
nand U5722 (N_5722,N_5307,N_5326);
nand U5723 (N_5723,N_5455,N_5393);
and U5724 (N_5724,N_5447,N_5441);
nor U5725 (N_5725,N_5322,N_5346);
or U5726 (N_5726,N_5298,N_5463);
nand U5727 (N_5727,N_5395,N_5457);
xor U5728 (N_5728,N_5366,N_5427);
xnor U5729 (N_5729,N_5328,N_5457);
nor U5730 (N_5730,N_5420,N_5417);
nor U5731 (N_5731,N_5474,N_5410);
xor U5732 (N_5732,N_5379,N_5497);
xor U5733 (N_5733,N_5356,N_5340);
nor U5734 (N_5734,N_5334,N_5388);
or U5735 (N_5735,N_5302,N_5378);
nor U5736 (N_5736,N_5296,N_5425);
nand U5737 (N_5737,N_5336,N_5393);
and U5738 (N_5738,N_5499,N_5262);
and U5739 (N_5739,N_5360,N_5324);
nand U5740 (N_5740,N_5414,N_5445);
and U5741 (N_5741,N_5392,N_5366);
xnor U5742 (N_5742,N_5268,N_5443);
nor U5743 (N_5743,N_5443,N_5321);
nor U5744 (N_5744,N_5405,N_5252);
or U5745 (N_5745,N_5454,N_5296);
nand U5746 (N_5746,N_5289,N_5414);
nand U5747 (N_5747,N_5346,N_5451);
nand U5748 (N_5748,N_5338,N_5310);
or U5749 (N_5749,N_5298,N_5387);
and U5750 (N_5750,N_5565,N_5502);
nor U5751 (N_5751,N_5606,N_5736);
nand U5752 (N_5752,N_5612,N_5568);
nand U5753 (N_5753,N_5540,N_5599);
or U5754 (N_5754,N_5547,N_5585);
nand U5755 (N_5755,N_5653,N_5644);
nand U5756 (N_5756,N_5594,N_5588);
and U5757 (N_5757,N_5596,N_5580);
nand U5758 (N_5758,N_5514,N_5741);
xnor U5759 (N_5759,N_5522,N_5687);
xor U5760 (N_5760,N_5627,N_5717);
and U5761 (N_5761,N_5551,N_5508);
nor U5762 (N_5762,N_5680,N_5593);
or U5763 (N_5763,N_5509,N_5639);
and U5764 (N_5764,N_5692,N_5590);
nor U5765 (N_5765,N_5711,N_5507);
and U5766 (N_5766,N_5578,N_5607);
and U5767 (N_5767,N_5631,N_5564);
xor U5768 (N_5768,N_5729,N_5661);
xnor U5769 (N_5769,N_5684,N_5690);
and U5770 (N_5770,N_5724,N_5703);
xnor U5771 (N_5771,N_5604,N_5586);
xnor U5772 (N_5772,N_5681,N_5746);
nand U5773 (N_5773,N_5732,N_5542);
nand U5774 (N_5774,N_5519,N_5698);
nand U5775 (N_5775,N_5669,N_5714);
nor U5776 (N_5776,N_5674,N_5614);
nor U5777 (N_5777,N_5647,N_5621);
nand U5778 (N_5778,N_5572,N_5728);
and U5779 (N_5779,N_5738,N_5634);
nand U5780 (N_5780,N_5718,N_5628);
xnor U5781 (N_5781,N_5595,N_5506);
nand U5782 (N_5782,N_5529,N_5528);
nor U5783 (N_5783,N_5570,N_5613);
and U5784 (N_5784,N_5615,N_5662);
nor U5785 (N_5785,N_5598,N_5641);
nor U5786 (N_5786,N_5739,N_5555);
nor U5787 (N_5787,N_5510,N_5575);
xnor U5788 (N_5788,N_5707,N_5525);
nor U5789 (N_5789,N_5747,N_5679);
xnor U5790 (N_5790,N_5642,N_5638);
xor U5791 (N_5791,N_5640,N_5597);
xor U5792 (N_5792,N_5643,N_5582);
nand U5793 (N_5793,N_5589,N_5699);
or U5794 (N_5794,N_5715,N_5683);
xor U5795 (N_5795,N_5544,N_5671);
nand U5796 (N_5796,N_5696,N_5516);
nand U5797 (N_5797,N_5676,N_5523);
nand U5798 (N_5798,N_5533,N_5501);
or U5799 (N_5799,N_5546,N_5592);
nand U5800 (N_5800,N_5670,N_5550);
nor U5801 (N_5801,N_5538,N_5623);
nor U5802 (N_5802,N_5712,N_5743);
nand U5803 (N_5803,N_5625,N_5733);
nand U5804 (N_5804,N_5720,N_5695);
nor U5805 (N_5805,N_5652,N_5742);
nor U5806 (N_5806,N_5622,N_5563);
nor U5807 (N_5807,N_5536,N_5633);
and U5808 (N_5808,N_5531,N_5554);
nand U5809 (N_5809,N_5504,N_5503);
or U5810 (N_5810,N_5745,N_5527);
or U5811 (N_5811,N_5620,N_5734);
nor U5812 (N_5812,N_5559,N_5664);
xor U5813 (N_5813,N_5658,N_5672);
and U5814 (N_5814,N_5629,N_5524);
xnor U5815 (N_5815,N_5610,N_5710);
xor U5816 (N_5816,N_5657,N_5654);
nand U5817 (N_5817,N_5505,N_5584);
nor U5818 (N_5818,N_5624,N_5637);
xor U5819 (N_5819,N_5583,N_5727);
and U5820 (N_5820,N_5602,N_5665);
nor U5821 (N_5821,N_5691,N_5571);
or U5822 (N_5822,N_5539,N_5689);
xor U5823 (N_5823,N_5512,N_5705);
or U5824 (N_5824,N_5731,N_5579);
nand U5825 (N_5825,N_5557,N_5721);
or U5826 (N_5826,N_5726,N_5603);
and U5827 (N_5827,N_5673,N_5520);
and U5828 (N_5828,N_5682,N_5740);
nor U5829 (N_5829,N_5697,N_5737);
and U5830 (N_5830,N_5735,N_5630);
or U5831 (N_5831,N_5635,N_5675);
and U5832 (N_5832,N_5655,N_5611);
nor U5833 (N_5833,N_5706,N_5744);
and U5834 (N_5834,N_5618,N_5659);
xor U5835 (N_5835,N_5651,N_5561);
and U5836 (N_5836,N_5701,N_5619);
and U5837 (N_5837,N_5632,N_5685);
xor U5838 (N_5838,N_5660,N_5515);
nor U5839 (N_5839,N_5581,N_5648);
or U5840 (N_5840,N_5521,N_5713);
xnor U5841 (N_5841,N_5560,N_5537);
and U5842 (N_5842,N_5667,N_5656);
nand U5843 (N_5843,N_5723,N_5549);
xor U5844 (N_5844,N_5716,N_5693);
nand U5845 (N_5845,N_5543,N_5636);
nand U5846 (N_5846,N_5608,N_5562);
nor U5847 (N_5847,N_5649,N_5722);
nand U5848 (N_5848,N_5666,N_5567);
nor U5849 (N_5849,N_5605,N_5650);
nor U5850 (N_5850,N_5545,N_5709);
nand U5851 (N_5851,N_5748,N_5500);
nand U5852 (N_5852,N_5730,N_5576);
and U5853 (N_5853,N_5663,N_5573);
xor U5854 (N_5854,N_5688,N_5574);
nor U5855 (N_5855,N_5616,N_5534);
xor U5856 (N_5856,N_5558,N_5569);
and U5857 (N_5857,N_5511,N_5541);
nor U5858 (N_5858,N_5702,N_5645);
and U5859 (N_5859,N_5587,N_5601);
and U5860 (N_5860,N_5532,N_5725);
xnor U5861 (N_5861,N_5646,N_5678);
xnor U5862 (N_5862,N_5600,N_5694);
and U5863 (N_5863,N_5552,N_5548);
xnor U5864 (N_5864,N_5553,N_5526);
or U5865 (N_5865,N_5535,N_5704);
nor U5866 (N_5866,N_5617,N_5556);
and U5867 (N_5867,N_5518,N_5708);
or U5868 (N_5868,N_5686,N_5719);
nand U5869 (N_5869,N_5626,N_5577);
nand U5870 (N_5870,N_5513,N_5517);
or U5871 (N_5871,N_5677,N_5609);
xnor U5872 (N_5872,N_5530,N_5591);
or U5873 (N_5873,N_5700,N_5566);
and U5874 (N_5874,N_5668,N_5749);
nand U5875 (N_5875,N_5506,N_5707);
nor U5876 (N_5876,N_5639,N_5576);
nand U5877 (N_5877,N_5611,N_5608);
nand U5878 (N_5878,N_5513,N_5686);
or U5879 (N_5879,N_5526,N_5619);
and U5880 (N_5880,N_5589,N_5608);
nand U5881 (N_5881,N_5636,N_5642);
or U5882 (N_5882,N_5507,N_5529);
xor U5883 (N_5883,N_5674,N_5541);
nor U5884 (N_5884,N_5520,N_5503);
or U5885 (N_5885,N_5610,N_5681);
nor U5886 (N_5886,N_5707,N_5729);
or U5887 (N_5887,N_5690,N_5565);
and U5888 (N_5888,N_5668,N_5561);
nor U5889 (N_5889,N_5636,N_5648);
nor U5890 (N_5890,N_5741,N_5594);
xor U5891 (N_5891,N_5718,N_5627);
xor U5892 (N_5892,N_5502,N_5531);
xnor U5893 (N_5893,N_5650,N_5557);
nor U5894 (N_5894,N_5564,N_5726);
nand U5895 (N_5895,N_5719,N_5731);
and U5896 (N_5896,N_5667,N_5699);
xor U5897 (N_5897,N_5582,N_5701);
xor U5898 (N_5898,N_5670,N_5545);
and U5899 (N_5899,N_5618,N_5620);
nand U5900 (N_5900,N_5615,N_5604);
nor U5901 (N_5901,N_5637,N_5646);
xnor U5902 (N_5902,N_5713,N_5744);
and U5903 (N_5903,N_5503,N_5643);
nand U5904 (N_5904,N_5532,N_5679);
xnor U5905 (N_5905,N_5736,N_5653);
and U5906 (N_5906,N_5567,N_5695);
xor U5907 (N_5907,N_5551,N_5714);
nor U5908 (N_5908,N_5523,N_5698);
or U5909 (N_5909,N_5606,N_5666);
or U5910 (N_5910,N_5570,N_5553);
and U5911 (N_5911,N_5626,N_5547);
nor U5912 (N_5912,N_5551,N_5596);
xor U5913 (N_5913,N_5739,N_5661);
xnor U5914 (N_5914,N_5685,N_5545);
and U5915 (N_5915,N_5689,N_5520);
or U5916 (N_5916,N_5566,N_5731);
and U5917 (N_5917,N_5749,N_5632);
nor U5918 (N_5918,N_5564,N_5575);
and U5919 (N_5919,N_5563,N_5562);
xnor U5920 (N_5920,N_5677,N_5718);
nor U5921 (N_5921,N_5524,N_5747);
nand U5922 (N_5922,N_5543,N_5541);
and U5923 (N_5923,N_5524,N_5621);
nor U5924 (N_5924,N_5707,N_5621);
and U5925 (N_5925,N_5674,N_5700);
xnor U5926 (N_5926,N_5626,N_5675);
or U5927 (N_5927,N_5636,N_5571);
or U5928 (N_5928,N_5736,N_5546);
nor U5929 (N_5929,N_5658,N_5701);
nand U5930 (N_5930,N_5604,N_5535);
nand U5931 (N_5931,N_5514,N_5707);
or U5932 (N_5932,N_5509,N_5703);
nand U5933 (N_5933,N_5704,N_5618);
or U5934 (N_5934,N_5570,N_5555);
or U5935 (N_5935,N_5732,N_5526);
xor U5936 (N_5936,N_5513,N_5515);
nor U5937 (N_5937,N_5605,N_5727);
xnor U5938 (N_5938,N_5668,N_5632);
or U5939 (N_5939,N_5611,N_5539);
xnor U5940 (N_5940,N_5660,N_5713);
and U5941 (N_5941,N_5589,N_5678);
and U5942 (N_5942,N_5581,N_5631);
nor U5943 (N_5943,N_5740,N_5727);
nand U5944 (N_5944,N_5599,N_5657);
and U5945 (N_5945,N_5554,N_5745);
nand U5946 (N_5946,N_5522,N_5736);
xnor U5947 (N_5947,N_5544,N_5549);
nor U5948 (N_5948,N_5549,N_5558);
or U5949 (N_5949,N_5530,N_5598);
nand U5950 (N_5950,N_5558,N_5573);
and U5951 (N_5951,N_5688,N_5597);
or U5952 (N_5952,N_5559,N_5504);
nor U5953 (N_5953,N_5511,N_5732);
nand U5954 (N_5954,N_5600,N_5671);
or U5955 (N_5955,N_5674,N_5715);
xnor U5956 (N_5956,N_5742,N_5731);
and U5957 (N_5957,N_5601,N_5700);
and U5958 (N_5958,N_5531,N_5542);
and U5959 (N_5959,N_5669,N_5610);
xor U5960 (N_5960,N_5709,N_5697);
and U5961 (N_5961,N_5542,N_5565);
nand U5962 (N_5962,N_5564,N_5540);
nor U5963 (N_5963,N_5701,N_5633);
xor U5964 (N_5964,N_5644,N_5693);
xor U5965 (N_5965,N_5564,N_5637);
nor U5966 (N_5966,N_5655,N_5534);
nand U5967 (N_5967,N_5642,N_5532);
nor U5968 (N_5968,N_5709,N_5736);
xnor U5969 (N_5969,N_5747,N_5564);
nand U5970 (N_5970,N_5674,N_5723);
and U5971 (N_5971,N_5700,N_5746);
nor U5972 (N_5972,N_5746,N_5740);
and U5973 (N_5973,N_5728,N_5691);
or U5974 (N_5974,N_5685,N_5672);
or U5975 (N_5975,N_5607,N_5728);
and U5976 (N_5976,N_5698,N_5508);
xor U5977 (N_5977,N_5552,N_5541);
nor U5978 (N_5978,N_5698,N_5613);
nand U5979 (N_5979,N_5671,N_5693);
xnor U5980 (N_5980,N_5700,N_5513);
and U5981 (N_5981,N_5666,N_5626);
or U5982 (N_5982,N_5570,N_5742);
nand U5983 (N_5983,N_5623,N_5616);
nand U5984 (N_5984,N_5550,N_5647);
nand U5985 (N_5985,N_5633,N_5729);
xnor U5986 (N_5986,N_5668,N_5597);
and U5987 (N_5987,N_5663,N_5521);
xor U5988 (N_5988,N_5598,N_5534);
xor U5989 (N_5989,N_5679,N_5631);
and U5990 (N_5990,N_5679,N_5696);
nor U5991 (N_5991,N_5543,N_5621);
xor U5992 (N_5992,N_5712,N_5713);
or U5993 (N_5993,N_5663,N_5611);
nor U5994 (N_5994,N_5628,N_5713);
and U5995 (N_5995,N_5632,N_5740);
and U5996 (N_5996,N_5529,N_5639);
nand U5997 (N_5997,N_5666,N_5519);
nand U5998 (N_5998,N_5624,N_5718);
nand U5999 (N_5999,N_5534,N_5587);
nor U6000 (N_6000,N_5812,N_5910);
nor U6001 (N_6001,N_5999,N_5886);
nand U6002 (N_6002,N_5839,N_5797);
nor U6003 (N_6003,N_5976,N_5768);
or U6004 (N_6004,N_5933,N_5905);
or U6005 (N_6005,N_5810,N_5777);
xor U6006 (N_6006,N_5757,N_5780);
nand U6007 (N_6007,N_5907,N_5982);
xnor U6008 (N_6008,N_5852,N_5921);
xor U6009 (N_6009,N_5965,N_5860);
nand U6010 (N_6010,N_5826,N_5937);
nor U6011 (N_6011,N_5952,N_5991);
xor U6012 (N_6012,N_5775,N_5916);
and U6013 (N_6013,N_5786,N_5846);
nor U6014 (N_6014,N_5863,N_5875);
nor U6015 (N_6015,N_5801,N_5960);
and U6016 (N_6016,N_5998,N_5803);
xor U6017 (N_6017,N_5844,N_5945);
nor U6018 (N_6018,N_5782,N_5977);
nand U6019 (N_6019,N_5861,N_5979);
nor U6020 (N_6020,N_5963,N_5829);
nand U6021 (N_6021,N_5908,N_5843);
nor U6022 (N_6022,N_5769,N_5848);
nand U6023 (N_6023,N_5867,N_5823);
xor U6024 (N_6024,N_5834,N_5988);
or U6025 (N_6025,N_5888,N_5955);
nor U6026 (N_6026,N_5943,N_5840);
or U6027 (N_6027,N_5898,N_5983);
or U6028 (N_6028,N_5940,N_5959);
xnor U6029 (N_6029,N_5900,N_5774);
nand U6030 (N_6030,N_5750,N_5809);
nor U6031 (N_6031,N_5752,N_5990);
and U6032 (N_6032,N_5909,N_5985);
nor U6033 (N_6033,N_5891,N_5760);
or U6034 (N_6034,N_5927,N_5767);
and U6035 (N_6035,N_5854,N_5997);
nor U6036 (N_6036,N_5974,N_5948);
and U6037 (N_6037,N_5805,N_5785);
nor U6038 (N_6038,N_5773,N_5831);
and U6039 (N_6039,N_5939,N_5830);
nand U6040 (N_6040,N_5930,N_5971);
nand U6041 (N_6041,N_5894,N_5987);
and U6042 (N_6042,N_5765,N_5795);
xor U6043 (N_6043,N_5996,N_5928);
and U6044 (N_6044,N_5804,N_5827);
nor U6045 (N_6045,N_5808,N_5904);
or U6046 (N_6046,N_5756,N_5980);
nor U6047 (N_6047,N_5942,N_5766);
and U6048 (N_6048,N_5876,N_5871);
nor U6049 (N_6049,N_5889,N_5869);
nor U6050 (N_6050,N_5978,N_5895);
nand U6051 (N_6051,N_5878,N_5903);
xor U6052 (N_6052,N_5883,N_5864);
or U6053 (N_6053,N_5944,N_5761);
nor U6054 (N_6054,N_5970,N_5936);
xnor U6055 (N_6055,N_5914,N_5759);
xor U6056 (N_6056,N_5851,N_5794);
or U6057 (N_6057,N_5918,N_5778);
or U6058 (N_6058,N_5992,N_5956);
nor U6059 (N_6059,N_5814,N_5923);
xnor U6060 (N_6060,N_5853,N_5873);
xor U6061 (N_6061,N_5981,N_5802);
nor U6062 (N_6062,N_5995,N_5882);
or U6063 (N_6063,N_5967,N_5920);
xor U6064 (N_6064,N_5941,N_5820);
or U6065 (N_6065,N_5924,N_5932);
nand U6066 (N_6066,N_5799,N_5790);
and U6067 (N_6067,N_5817,N_5946);
nor U6068 (N_6068,N_5962,N_5807);
nand U6069 (N_6069,N_5954,N_5806);
and U6070 (N_6070,N_5925,N_5881);
nor U6071 (N_6071,N_5969,N_5847);
xor U6072 (N_6072,N_5911,N_5776);
or U6073 (N_6073,N_5865,N_5961);
or U6074 (N_6074,N_5929,N_5815);
or U6075 (N_6075,N_5993,N_5841);
and U6076 (N_6076,N_5788,N_5800);
xnor U6077 (N_6077,N_5947,N_5835);
and U6078 (N_6078,N_5789,N_5966);
and U6079 (N_6079,N_5922,N_5949);
nand U6080 (N_6080,N_5850,N_5866);
nand U6081 (N_6081,N_5915,N_5912);
nor U6082 (N_6082,N_5906,N_5816);
nand U6083 (N_6083,N_5935,N_5934);
nor U6084 (N_6084,N_5870,N_5836);
and U6085 (N_6085,N_5825,N_5938);
nor U6086 (N_6086,N_5872,N_5771);
nor U6087 (N_6087,N_5887,N_5770);
or U6088 (N_6088,N_5845,N_5796);
or U6089 (N_6089,N_5896,N_5899);
nor U6090 (N_6090,N_5951,N_5833);
or U6091 (N_6091,N_5855,N_5986);
nor U6092 (N_6092,N_5975,N_5885);
nand U6093 (N_6093,N_5751,N_5755);
or U6094 (N_6094,N_5994,N_5818);
xnor U6095 (N_6095,N_5781,N_5931);
or U6096 (N_6096,N_5784,N_5917);
and U6097 (N_6097,N_5792,N_5838);
and U6098 (N_6098,N_5972,N_5824);
or U6099 (N_6099,N_5849,N_5879);
or U6100 (N_6100,N_5821,N_5763);
nand U6101 (N_6101,N_5779,N_5764);
xnor U6102 (N_6102,N_5884,N_5811);
nor U6103 (N_6103,N_5842,N_5791);
xor U6104 (N_6104,N_5968,N_5819);
nor U6105 (N_6105,N_5813,N_5957);
nor U6106 (N_6106,N_5926,N_5973);
nand U6107 (N_6107,N_5754,N_5877);
nor U6108 (N_6108,N_5893,N_5989);
nor U6109 (N_6109,N_5832,N_5880);
nor U6110 (N_6110,N_5758,N_5953);
nor U6111 (N_6111,N_5868,N_5753);
or U6112 (N_6112,N_5772,N_5874);
and U6113 (N_6113,N_5897,N_5901);
nand U6114 (N_6114,N_5913,N_5890);
nand U6115 (N_6115,N_5902,N_5857);
nand U6116 (N_6116,N_5762,N_5858);
or U6117 (N_6117,N_5787,N_5822);
xor U6118 (N_6118,N_5793,N_5950);
nor U6119 (N_6119,N_5798,N_5856);
nand U6120 (N_6120,N_5964,N_5958);
xor U6121 (N_6121,N_5837,N_5859);
xnor U6122 (N_6122,N_5892,N_5862);
nor U6123 (N_6123,N_5828,N_5783);
xor U6124 (N_6124,N_5919,N_5984);
nand U6125 (N_6125,N_5981,N_5886);
and U6126 (N_6126,N_5911,N_5822);
and U6127 (N_6127,N_5886,N_5764);
nor U6128 (N_6128,N_5990,N_5780);
or U6129 (N_6129,N_5894,N_5898);
or U6130 (N_6130,N_5924,N_5786);
nand U6131 (N_6131,N_5767,N_5783);
nand U6132 (N_6132,N_5893,N_5863);
nand U6133 (N_6133,N_5910,N_5997);
or U6134 (N_6134,N_5773,N_5931);
nand U6135 (N_6135,N_5909,N_5847);
nand U6136 (N_6136,N_5900,N_5985);
nor U6137 (N_6137,N_5886,N_5880);
nand U6138 (N_6138,N_5906,N_5984);
nand U6139 (N_6139,N_5894,N_5861);
or U6140 (N_6140,N_5956,N_5837);
or U6141 (N_6141,N_5808,N_5771);
xor U6142 (N_6142,N_5889,N_5779);
nor U6143 (N_6143,N_5984,N_5852);
or U6144 (N_6144,N_5787,N_5869);
xor U6145 (N_6145,N_5774,N_5916);
and U6146 (N_6146,N_5927,N_5906);
xor U6147 (N_6147,N_5827,N_5840);
nor U6148 (N_6148,N_5978,N_5795);
or U6149 (N_6149,N_5790,N_5997);
or U6150 (N_6150,N_5818,N_5967);
or U6151 (N_6151,N_5973,N_5960);
nor U6152 (N_6152,N_5884,N_5765);
and U6153 (N_6153,N_5779,N_5906);
nand U6154 (N_6154,N_5935,N_5761);
and U6155 (N_6155,N_5811,N_5774);
nand U6156 (N_6156,N_5762,N_5842);
nand U6157 (N_6157,N_5902,N_5792);
nand U6158 (N_6158,N_5934,N_5779);
nand U6159 (N_6159,N_5822,N_5842);
and U6160 (N_6160,N_5974,N_5815);
xor U6161 (N_6161,N_5897,N_5769);
xnor U6162 (N_6162,N_5877,N_5867);
nor U6163 (N_6163,N_5779,N_5892);
nor U6164 (N_6164,N_5873,N_5867);
nand U6165 (N_6165,N_5782,N_5829);
xor U6166 (N_6166,N_5852,N_5956);
and U6167 (N_6167,N_5936,N_5858);
nor U6168 (N_6168,N_5803,N_5824);
and U6169 (N_6169,N_5897,N_5961);
and U6170 (N_6170,N_5870,N_5923);
nand U6171 (N_6171,N_5993,N_5839);
or U6172 (N_6172,N_5879,N_5775);
nor U6173 (N_6173,N_5923,N_5933);
nand U6174 (N_6174,N_5796,N_5777);
xor U6175 (N_6175,N_5940,N_5782);
and U6176 (N_6176,N_5979,N_5996);
nor U6177 (N_6177,N_5814,N_5966);
or U6178 (N_6178,N_5926,N_5855);
and U6179 (N_6179,N_5835,N_5811);
and U6180 (N_6180,N_5759,N_5906);
or U6181 (N_6181,N_5997,N_5753);
nand U6182 (N_6182,N_5833,N_5787);
nor U6183 (N_6183,N_5792,N_5997);
and U6184 (N_6184,N_5830,N_5836);
xor U6185 (N_6185,N_5759,N_5962);
nor U6186 (N_6186,N_5940,N_5824);
nand U6187 (N_6187,N_5975,N_5953);
nor U6188 (N_6188,N_5782,N_5819);
nand U6189 (N_6189,N_5792,N_5996);
nor U6190 (N_6190,N_5796,N_5919);
or U6191 (N_6191,N_5999,N_5798);
nand U6192 (N_6192,N_5878,N_5776);
and U6193 (N_6193,N_5989,N_5971);
and U6194 (N_6194,N_5889,N_5875);
nor U6195 (N_6195,N_5795,N_5948);
nand U6196 (N_6196,N_5863,N_5945);
or U6197 (N_6197,N_5814,N_5919);
and U6198 (N_6198,N_5894,N_5790);
or U6199 (N_6199,N_5945,N_5906);
nand U6200 (N_6200,N_5909,N_5753);
or U6201 (N_6201,N_5967,N_5857);
xor U6202 (N_6202,N_5873,N_5849);
or U6203 (N_6203,N_5883,N_5959);
or U6204 (N_6204,N_5829,N_5836);
nand U6205 (N_6205,N_5769,N_5879);
xor U6206 (N_6206,N_5911,N_5989);
nor U6207 (N_6207,N_5980,N_5856);
nand U6208 (N_6208,N_5828,N_5814);
nand U6209 (N_6209,N_5825,N_5905);
or U6210 (N_6210,N_5938,N_5932);
or U6211 (N_6211,N_5818,N_5788);
and U6212 (N_6212,N_5779,N_5916);
xnor U6213 (N_6213,N_5895,N_5853);
xor U6214 (N_6214,N_5817,N_5771);
and U6215 (N_6215,N_5791,N_5928);
nand U6216 (N_6216,N_5757,N_5853);
xor U6217 (N_6217,N_5872,N_5858);
xor U6218 (N_6218,N_5940,N_5846);
nand U6219 (N_6219,N_5961,N_5782);
nor U6220 (N_6220,N_5790,N_5755);
xor U6221 (N_6221,N_5950,N_5773);
nor U6222 (N_6222,N_5893,N_5768);
nor U6223 (N_6223,N_5990,N_5875);
nand U6224 (N_6224,N_5942,N_5904);
xor U6225 (N_6225,N_5910,N_5948);
nand U6226 (N_6226,N_5821,N_5751);
and U6227 (N_6227,N_5895,N_5797);
xnor U6228 (N_6228,N_5871,N_5829);
nor U6229 (N_6229,N_5819,N_5996);
nor U6230 (N_6230,N_5911,N_5953);
or U6231 (N_6231,N_5787,N_5872);
xnor U6232 (N_6232,N_5797,N_5914);
or U6233 (N_6233,N_5992,N_5803);
or U6234 (N_6234,N_5805,N_5974);
nand U6235 (N_6235,N_5983,N_5814);
nor U6236 (N_6236,N_5951,N_5911);
and U6237 (N_6237,N_5998,N_5890);
or U6238 (N_6238,N_5817,N_5870);
and U6239 (N_6239,N_5785,N_5764);
xnor U6240 (N_6240,N_5992,N_5901);
nand U6241 (N_6241,N_5760,N_5949);
nand U6242 (N_6242,N_5974,N_5966);
xor U6243 (N_6243,N_5925,N_5942);
nand U6244 (N_6244,N_5898,N_5967);
nand U6245 (N_6245,N_5993,N_5800);
and U6246 (N_6246,N_5797,N_5946);
xnor U6247 (N_6247,N_5785,N_5973);
nand U6248 (N_6248,N_5791,N_5798);
nor U6249 (N_6249,N_5900,N_5753);
and U6250 (N_6250,N_6051,N_6049);
nand U6251 (N_6251,N_6151,N_6142);
and U6252 (N_6252,N_6196,N_6247);
xor U6253 (N_6253,N_6188,N_6123);
nor U6254 (N_6254,N_6175,N_6086);
xor U6255 (N_6255,N_6139,N_6232);
xor U6256 (N_6256,N_6120,N_6143);
or U6257 (N_6257,N_6007,N_6066);
xor U6258 (N_6258,N_6116,N_6203);
nand U6259 (N_6259,N_6003,N_6119);
nor U6260 (N_6260,N_6057,N_6226);
and U6261 (N_6261,N_6213,N_6117);
and U6262 (N_6262,N_6233,N_6236);
and U6263 (N_6263,N_6046,N_6174);
xnor U6264 (N_6264,N_6092,N_6228);
nand U6265 (N_6265,N_6054,N_6141);
or U6266 (N_6266,N_6004,N_6109);
or U6267 (N_6267,N_6069,N_6208);
or U6268 (N_6268,N_6146,N_6118);
nand U6269 (N_6269,N_6210,N_6005);
nand U6270 (N_6270,N_6212,N_6091);
nand U6271 (N_6271,N_6076,N_6112);
or U6272 (N_6272,N_6240,N_6101);
or U6273 (N_6273,N_6144,N_6053);
nand U6274 (N_6274,N_6088,N_6100);
and U6275 (N_6275,N_6089,N_6098);
and U6276 (N_6276,N_6055,N_6105);
nand U6277 (N_6277,N_6068,N_6081);
or U6278 (N_6278,N_6052,N_6031);
and U6279 (N_6279,N_6245,N_6215);
xor U6280 (N_6280,N_6164,N_6234);
nand U6281 (N_6281,N_6063,N_6130);
xnor U6282 (N_6282,N_6201,N_6248);
nand U6283 (N_6283,N_6166,N_6000);
or U6284 (N_6284,N_6029,N_6173);
xnor U6285 (N_6285,N_6114,N_6168);
xor U6286 (N_6286,N_6161,N_6194);
or U6287 (N_6287,N_6061,N_6097);
nor U6288 (N_6288,N_6195,N_6067);
and U6289 (N_6289,N_6036,N_6012);
or U6290 (N_6290,N_6186,N_6157);
nand U6291 (N_6291,N_6011,N_6206);
or U6292 (N_6292,N_6178,N_6059);
and U6293 (N_6293,N_6093,N_6246);
xor U6294 (N_6294,N_6034,N_6028);
nand U6295 (N_6295,N_6043,N_6115);
nor U6296 (N_6296,N_6140,N_6223);
nand U6297 (N_6297,N_6087,N_6138);
or U6298 (N_6298,N_6129,N_6229);
nor U6299 (N_6299,N_6024,N_6113);
and U6300 (N_6300,N_6017,N_6176);
xnor U6301 (N_6301,N_6127,N_6102);
xnor U6302 (N_6302,N_6227,N_6207);
and U6303 (N_6303,N_6071,N_6077);
or U6304 (N_6304,N_6183,N_6243);
and U6305 (N_6305,N_6056,N_6058);
nor U6306 (N_6306,N_6211,N_6122);
and U6307 (N_6307,N_6185,N_6009);
or U6308 (N_6308,N_6078,N_6008);
nand U6309 (N_6309,N_6225,N_6108);
nand U6310 (N_6310,N_6182,N_6099);
or U6311 (N_6311,N_6191,N_6190);
nand U6312 (N_6312,N_6065,N_6047);
nor U6313 (N_6313,N_6096,N_6032);
or U6314 (N_6314,N_6060,N_6027);
and U6315 (N_6315,N_6180,N_6220);
xor U6316 (N_6316,N_6222,N_6241);
nor U6317 (N_6317,N_6133,N_6103);
nor U6318 (N_6318,N_6167,N_6231);
or U6319 (N_6319,N_6082,N_6015);
nor U6320 (N_6320,N_6132,N_6170);
xor U6321 (N_6321,N_6001,N_6070);
xor U6322 (N_6322,N_6218,N_6237);
and U6323 (N_6323,N_6209,N_6171);
or U6324 (N_6324,N_6050,N_6073);
nand U6325 (N_6325,N_6149,N_6104);
or U6326 (N_6326,N_6181,N_6165);
nor U6327 (N_6327,N_6016,N_6090);
nand U6328 (N_6328,N_6107,N_6010);
xnor U6329 (N_6329,N_6162,N_6064);
or U6330 (N_6330,N_6013,N_6199);
nor U6331 (N_6331,N_6037,N_6221);
or U6332 (N_6332,N_6075,N_6153);
nand U6333 (N_6333,N_6084,N_6192);
or U6334 (N_6334,N_6124,N_6026);
nor U6335 (N_6335,N_6177,N_6189);
nand U6336 (N_6336,N_6147,N_6074);
and U6337 (N_6337,N_6235,N_6169);
nor U6338 (N_6338,N_6111,N_6038);
xor U6339 (N_6339,N_6020,N_6238);
or U6340 (N_6340,N_6244,N_6224);
nand U6341 (N_6341,N_6085,N_6021);
and U6342 (N_6342,N_6137,N_6150);
or U6343 (N_6343,N_6048,N_6072);
xor U6344 (N_6344,N_6042,N_6006);
xor U6345 (N_6345,N_6014,N_6179);
nor U6346 (N_6346,N_6035,N_6040);
nor U6347 (N_6347,N_6136,N_6152);
nor U6348 (N_6348,N_6023,N_6018);
nand U6349 (N_6349,N_6160,N_6204);
or U6350 (N_6350,N_6249,N_6041);
and U6351 (N_6351,N_6156,N_6030);
and U6352 (N_6352,N_6135,N_6214);
or U6353 (N_6353,N_6044,N_6125);
nor U6354 (N_6354,N_6155,N_6094);
xor U6355 (N_6355,N_6022,N_6095);
nor U6356 (N_6356,N_6230,N_6148);
nand U6357 (N_6357,N_6145,N_6039);
or U6358 (N_6358,N_6079,N_6193);
xnor U6359 (N_6359,N_6200,N_6205);
and U6360 (N_6360,N_6121,N_6080);
and U6361 (N_6361,N_6131,N_6239);
or U6362 (N_6362,N_6128,N_6163);
xor U6363 (N_6363,N_6106,N_6019);
nand U6364 (N_6364,N_6172,N_6062);
and U6365 (N_6365,N_6158,N_6219);
and U6366 (N_6366,N_6202,N_6045);
or U6367 (N_6367,N_6110,N_6083);
or U6368 (N_6368,N_6126,N_6217);
or U6369 (N_6369,N_6187,N_6134);
nor U6370 (N_6370,N_6216,N_6025);
nand U6371 (N_6371,N_6002,N_6154);
or U6372 (N_6372,N_6197,N_6184);
nor U6373 (N_6373,N_6159,N_6198);
xor U6374 (N_6374,N_6242,N_6033);
and U6375 (N_6375,N_6195,N_6013);
or U6376 (N_6376,N_6030,N_6088);
xnor U6377 (N_6377,N_6213,N_6202);
and U6378 (N_6378,N_6093,N_6088);
and U6379 (N_6379,N_6036,N_6038);
nand U6380 (N_6380,N_6041,N_6029);
and U6381 (N_6381,N_6049,N_6008);
nor U6382 (N_6382,N_6173,N_6135);
xnor U6383 (N_6383,N_6102,N_6129);
nor U6384 (N_6384,N_6182,N_6195);
and U6385 (N_6385,N_6218,N_6034);
xor U6386 (N_6386,N_6165,N_6031);
nor U6387 (N_6387,N_6077,N_6233);
nor U6388 (N_6388,N_6021,N_6135);
and U6389 (N_6389,N_6187,N_6145);
nor U6390 (N_6390,N_6024,N_6094);
nor U6391 (N_6391,N_6227,N_6194);
nand U6392 (N_6392,N_6091,N_6245);
or U6393 (N_6393,N_6095,N_6195);
or U6394 (N_6394,N_6057,N_6173);
nor U6395 (N_6395,N_6196,N_6015);
nor U6396 (N_6396,N_6179,N_6130);
nor U6397 (N_6397,N_6006,N_6230);
and U6398 (N_6398,N_6056,N_6069);
nand U6399 (N_6399,N_6233,N_6208);
or U6400 (N_6400,N_6129,N_6056);
nor U6401 (N_6401,N_6218,N_6026);
or U6402 (N_6402,N_6063,N_6076);
xnor U6403 (N_6403,N_6153,N_6069);
nor U6404 (N_6404,N_6207,N_6175);
nand U6405 (N_6405,N_6014,N_6040);
nand U6406 (N_6406,N_6189,N_6155);
xnor U6407 (N_6407,N_6072,N_6234);
or U6408 (N_6408,N_6167,N_6208);
and U6409 (N_6409,N_6140,N_6214);
xor U6410 (N_6410,N_6069,N_6102);
and U6411 (N_6411,N_6196,N_6010);
nor U6412 (N_6412,N_6050,N_6026);
xor U6413 (N_6413,N_6190,N_6197);
xor U6414 (N_6414,N_6140,N_6186);
nor U6415 (N_6415,N_6003,N_6112);
nand U6416 (N_6416,N_6095,N_6027);
and U6417 (N_6417,N_6149,N_6111);
xor U6418 (N_6418,N_6035,N_6195);
xnor U6419 (N_6419,N_6203,N_6062);
xor U6420 (N_6420,N_6137,N_6100);
and U6421 (N_6421,N_6145,N_6029);
and U6422 (N_6422,N_6182,N_6106);
xnor U6423 (N_6423,N_6030,N_6229);
or U6424 (N_6424,N_6012,N_6190);
and U6425 (N_6425,N_6074,N_6236);
and U6426 (N_6426,N_6109,N_6230);
and U6427 (N_6427,N_6170,N_6085);
and U6428 (N_6428,N_6017,N_6227);
nor U6429 (N_6429,N_6073,N_6009);
and U6430 (N_6430,N_6000,N_6219);
nand U6431 (N_6431,N_6039,N_6245);
and U6432 (N_6432,N_6107,N_6246);
and U6433 (N_6433,N_6230,N_6214);
nor U6434 (N_6434,N_6233,N_6076);
nor U6435 (N_6435,N_6176,N_6046);
nor U6436 (N_6436,N_6012,N_6163);
nand U6437 (N_6437,N_6155,N_6246);
xor U6438 (N_6438,N_6035,N_6130);
xnor U6439 (N_6439,N_6060,N_6209);
or U6440 (N_6440,N_6199,N_6114);
or U6441 (N_6441,N_6138,N_6081);
or U6442 (N_6442,N_6239,N_6223);
and U6443 (N_6443,N_6080,N_6054);
xor U6444 (N_6444,N_6244,N_6043);
xor U6445 (N_6445,N_6083,N_6218);
or U6446 (N_6446,N_6188,N_6214);
nand U6447 (N_6447,N_6135,N_6241);
nor U6448 (N_6448,N_6198,N_6002);
xor U6449 (N_6449,N_6198,N_6216);
xor U6450 (N_6450,N_6077,N_6155);
nor U6451 (N_6451,N_6067,N_6093);
nand U6452 (N_6452,N_6132,N_6223);
or U6453 (N_6453,N_6183,N_6135);
nand U6454 (N_6454,N_6089,N_6180);
xnor U6455 (N_6455,N_6108,N_6000);
nor U6456 (N_6456,N_6206,N_6151);
nor U6457 (N_6457,N_6023,N_6197);
or U6458 (N_6458,N_6006,N_6190);
nor U6459 (N_6459,N_6012,N_6069);
nand U6460 (N_6460,N_6073,N_6047);
and U6461 (N_6461,N_6185,N_6201);
xnor U6462 (N_6462,N_6144,N_6225);
or U6463 (N_6463,N_6174,N_6171);
nand U6464 (N_6464,N_6143,N_6248);
nor U6465 (N_6465,N_6037,N_6065);
or U6466 (N_6466,N_6152,N_6124);
nor U6467 (N_6467,N_6041,N_6224);
xor U6468 (N_6468,N_6025,N_6163);
and U6469 (N_6469,N_6117,N_6095);
nand U6470 (N_6470,N_6078,N_6015);
xor U6471 (N_6471,N_6193,N_6167);
and U6472 (N_6472,N_6136,N_6202);
or U6473 (N_6473,N_6095,N_6129);
and U6474 (N_6474,N_6200,N_6225);
nor U6475 (N_6475,N_6086,N_6181);
or U6476 (N_6476,N_6139,N_6080);
xnor U6477 (N_6477,N_6063,N_6024);
and U6478 (N_6478,N_6003,N_6086);
nor U6479 (N_6479,N_6056,N_6216);
and U6480 (N_6480,N_6207,N_6040);
or U6481 (N_6481,N_6189,N_6239);
xor U6482 (N_6482,N_6238,N_6168);
and U6483 (N_6483,N_6174,N_6218);
nor U6484 (N_6484,N_6051,N_6164);
nand U6485 (N_6485,N_6006,N_6229);
xnor U6486 (N_6486,N_6017,N_6024);
and U6487 (N_6487,N_6166,N_6129);
nor U6488 (N_6488,N_6116,N_6068);
and U6489 (N_6489,N_6135,N_6142);
xor U6490 (N_6490,N_6082,N_6153);
and U6491 (N_6491,N_6102,N_6174);
or U6492 (N_6492,N_6115,N_6199);
nand U6493 (N_6493,N_6167,N_6200);
xor U6494 (N_6494,N_6242,N_6227);
nand U6495 (N_6495,N_6005,N_6104);
and U6496 (N_6496,N_6219,N_6229);
nor U6497 (N_6497,N_6085,N_6240);
nor U6498 (N_6498,N_6038,N_6078);
nand U6499 (N_6499,N_6249,N_6051);
and U6500 (N_6500,N_6469,N_6312);
xor U6501 (N_6501,N_6277,N_6446);
nand U6502 (N_6502,N_6353,N_6282);
or U6503 (N_6503,N_6360,N_6358);
nand U6504 (N_6504,N_6269,N_6430);
and U6505 (N_6505,N_6324,N_6288);
and U6506 (N_6506,N_6302,N_6256);
xnor U6507 (N_6507,N_6348,N_6291);
and U6508 (N_6508,N_6252,N_6434);
xnor U6509 (N_6509,N_6251,N_6262);
and U6510 (N_6510,N_6411,N_6383);
nand U6511 (N_6511,N_6280,N_6495);
or U6512 (N_6512,N_6419,N_6369);
nand U6513 (N_6513,N_6297,N_6479);
nor U6514 (N_6514,N_6349,N_6308);
and U6515 (N_6515,N_6400,N_6403);
xnor U6516 (N_6516,N_6265,N_6490);
nor U6517 (N_6517,N_6323,N_6373);
nor U6518 (N_6518,N_6330,N_6452);
or U6519 (N_6519,N_6498,N_6418);
nor U6520 (N_6520,N_6426,N_6260);
nand U6521 (N_6521,N_6285,N_6465);
xor U6522 (N_6522,N_6420,N_6341);
and U6523 (N_6523,N_6259,N_6384);
nand U6524 (N_6524,N_6334,N_6255);
or U6525 (N_6525,N_6301,N_6450);
nand U6526 (N_6526,N_6470,N_6332);
and U6527 (N_6527,N_6402,N_6437);
nor U6528 (N_6528,N_6365,N_6336);
nand U6529 (N_6529,N_6423,N_6471);
nand U6530 (N_6530,N_6363,N_6344);
nor U6531 (N_6531,N_6499,N_6389);
and U6532 (N_6532,N_6414,N_6431);
and U6533 (N_6533,N_6339,N_6325);
nand U6534 (N_6534,N_6326,N_6295);
nor U6535 (N_6535,N_6393,N_6333);
xor U6536 (N_6536,N_6435,N_6484);
nor U6537 (N_6537,N_6335,N_6307);
nand U6538 (N_6538,N_6309,N_6355);
nand U6539 (N_6539,N_6351,N_6364);
xor U6540 (N_6540,N_6340,N_6454);
or U6541 (N_6541,N_6440,N_6428);
and U6542 (N_6542,N_6395,N_6476);
nand U6543 (N_6543,N_6433,N_6381);
or U6544 (N_6544,N_6268,N_6493);
and U6545 (N_6545,N_6409,N_6274);
or U6546 (N_6546,N_6394,N_6250);
xnor U6547 (N_6547,N_6284,N_6375);
nand U6548 (N_6548,N_6457,N_6408);
nand U6549 (N_6549,N_6480,N_6441);
and U6550 (N_6550,N_6391,N_6468);
or U6551 (N_6551,N_6387,N_6281);
nor U6552 (N_6552,N_6464,N_6398);
xnor U6553 (N_6553,N_6292,N_6407);
and U6554 (N_6554,N_6397,N_6385);
xnor U6555 (N_6555,N_6315,N_6258);
or U6556 (N_6556,N_6346,N_6416);
or U6557 (N_6557,N_6311,N_6254);
or U6558 (N_6558,N_6405,N_6496);
xnor U6559 (N_6559,N_6412,N_6371);
xnor U6560 (N_6560,N_6319,N_6460);
or U6561 (N_6561,N_6267,N_6449);
xor U6562 (N_6562,N_6357,N_6456);
nor U6563 (N_6563,N_6316,N_6329);
xor U6564 (N_6564,N_6492,N_6366);
xnor U6565 (N_6565,N_6374,N_6487);
xnor U6566 (N_6566,N_6475,N_6310);
and U6567 (N_6567,N_6317,N_6261);
and U6568 (N_6568,N_6293,N_6376);
xor U6569 (N_6569,N_6392,N_6350);
xor U6570 (N_6570,N_6379,N_6410);
or U6571 (N_6571,N_6273,N_6290);
nand U6572 (N_6572,N_6270,N_6463);
or U6573 (N_6573,N_6474,N_6266);
nand U6574 (N_6574,N_6396,N_6271);
and U6575 (N_6575,N_6466,N_6415);
or U6576 (N_6576,N_6472,N_6305);
nor U6577 (N_6577,N_6367,N_6283);
nor U6578 (N_6578,N_6427,N_6486);
nand U6579 (N_6579,N_6424,N_6448);
and U6580 (N_6580,N_6343,N_6327);
nand U6581 (N_6581,N_6370,N_6488);
and U6582 (N_6582,N_6276,N_6362);
or U6583 (N_6583,N_6342,N_6287);
and U6584 (N_6584,N_6372,N_6485);
or U6585 (N_6585,N_6303,N_6455);
or U6586 (N_6586,N_6447,N_6337);
nand U6587 (N_6587,N_6483,N_6289);
nand U6588 (N_6588,N_6286,N_6299);
xnor U6589 (N_6589,N_6331,N_6356);
and U6590 (N_6590,N_6461,N_6473);
or U6591 (N_6591,N_6451,N_6482);
or U6592 (N_6592,N_6377,N_6304);
xor U6593 (N_6593,N_6306,N_6432);
and U6594 (N_6594,N_6368,N_6388);
nor U6595 (N_6595,N_6378,N_6497);
nand U6596 (N_6596,N_6354,N_6421);
and U6597 (N_6597,N_6338,N_6478);
nor U6598 (N_6598,N_6443,N_6328);
nor U6599 (N_6599,N_6453,N_6382);
nor U6600 (N_6600,N_6445,N_6386);
nor U6601 (N_6601,N_6359,N_6458);
and U6602 (N_6602,N_6494,N_6298);
or U6603 (N_6603,N_6361,N_6444);
nor U6604 (N_6604,N_6436,N_6314);
nor U6605 (N_6605,N_6272,N_6425);
and U6606 (N_6606,N_6406,N_6413);
xor U6607 (N_6607,N_6417,N_6462);
nand U6608 (N_6608,N_6320,N_6253);
or U6609 (N_6609,N_6390,N_6429);
nor U6610 (N_6610,N_6352,N_6399);
xnor U6611 (N_6611,N_6422,N_6439);
xor U6612 (N_6612,N_6318,N_6380);
nor U6613 (N_6613,N_6467,N_6257);
and U6614 (N_6614,N_6491,N_6294);
xor U6615 (N_6615,N_6296,N_6300);
xnor U6616 (N_6616,N_6279,N_6442);
or U6617 (N_6617,N_6275,N_6347);
nor U6618 (N_6618,N_6489,N_6477);
and U6619 (N_6619,N_6264,N_6321);
xnor U6620 (N_6620,N_6459,N_6278);
nor U6621 (N_6621,N_6313,N_6481);
xnor U6622 (N_6622,N_6401,N_6322);
or U6623 (N_6623,N_6263,N_6438);
xor U6624 (N_6624,N_6345,N_6404);
nand U6625 (N_6625,N_6494,N_6376);
or U6626 (N_6626,N_6439,N_6373);
xor U6627 (N_6627,N_6425,N_6346);
xor U6628 (N_6628,N_6491,N_6380);
nor U6629 (N_6629,N_6253,N_6357);
or U6630 (N_6630,N_6486,N_6270);
and U6631 (N_6631,N_6302,N_6435);
xnor U6632 (N_6632,N_6298,N_6495);
nand U6633 (N_6633,N_6497,N_6395);
or U6634 (N_6634,N_6374,N_6486);
nand U6635 (N_6635,N_6279,N_6441);
and U6636 (N_6636,N_6389,N_6481);
or U6637 (N_6637,N_6255,N_6457);
and U6638 (N_6638,N_6481,N_6339);
nand U6639 (N_6639,N_6312,N_6416);
and U6640 (N_6640,N_6465,N_6497);
nor U6641 (N_6641,N_6452,N_6324);
and U6642 (N_6642,N_6456,N_6412);
and U6643 (N_6643,N_6392,N_6477);
nand U6644 (N_6644,N_6371,N_6319);
xnor U6645 (N_6645,N_6276,N_6413);
nor U6646 (N_6646,N_6394,N_6459);
and U6647 (N_6647,N_6384,N_6287);
or U6648 (N_6648,N_6437,N_6472);
nand U6649 (N_6649,N_6336,N_6341);
nand U6650 (N_6650,N_6406,N_6277);
and U6651 (N_6651,N_6366,N_6359);
nand U6652 (N_6652,N_6431,N_6437);
nand U6653 (N_6653,N_6428,N_6318);
or U6654 (N_6654,N_6283,N_6292);
xnor U6655 (N_6655,N_6379,N_6411);
and U6656 (N_6656,N_6494,N_6309);
nand U6657 (N_6657,N_6262,N_6343);
nand U6658 (N_6658,N_6256,N_6495);
xnor U6659 (N_6659,N_6385,N_6401);
and U6660 (N_6660,N_6330,N_6281);
nor U6661 (N_6661,N_6369,N_6269);
nand U6662 (N_6662,N_6466,N_6319);
nor U6663 (N_6663,N_6308,N_6457);
and U6664 (N_6664,N_6293,N_6426);
or U6665 (N_6665,N_6447,N_6330);
xor U6666 (N_6666,N_6377,N_6267);
or U6667 (N_6667,N_6314,N_6258);
or U6668 (N_6668,N_6326,N_6339);
xor U6669 (N_6669,N_6353,N_6473);
nor U6670 (N_6670,N_6398,N_6388);
nand U6671 (N_6671,N_6474,N_6256);
xnor U6672 (N_6672,N_6261,N_6403);
or U6673 (N_6673,N_6398,N_6439);
or U6674 (N_6674,N_6428,N_6401);
and U6675 (N_6675,N_6450,N_6374);
nand U6676 (N_6676,N_6407,N_6270);
xnor U6677 (N_6677,N_6475,N_6254);
xor U6678 (N_6678,N_6403,N_6330);
xnor U6679 (N_6679,N_6358,N_6255);
or U6680 (N_6680,N_6482,N_6391);
xor U6681 (N_6681,N_6294,N_6374);
nor U6682 (N_6682,N_6466,N_6384);
or U6683 (N_6683,N_6317,N_6390);
nor U6684 (N_6684,N_6358,N_6434);
xor U6685 (N_6685,N_6430,N_6357);
nor U6686 (N_6686,N_6426,N_6450);
nor U6687 (N_6687,N_6319,N_6254);
and U6688 (N_6688,N_6357,N_6387);
or U6689 (N_6689,N_6496,N_6346);
or U6690 (N_6690,N_6276,N_6354);
and U6691 (N_6691,N_6290,N_6416);
and U6692 (N_6692,N_6456,N_6493);
or U6693 (N_6693,N_6365,N_6436);
xnor U6694 (N_6694,N_6395,N_6350);
or U6695 (N_6695,N_6286,N_6400);
or U6696 (N_6696,N_6374,N_6347);
or U6697 (N_6697,N_6354,N_6295);
nor U6698 (N_6698,N_6257,N_6354);
nand U6699 (N_6699,N_6255,N_6342);
and U6700 (N_6700,N_6390,N_6352);
and U6701 (N_6701,N_6291,N_6287);
and U6702 (N_6702,N_6368,N_6369);
nor U6703 (N_6703,N_6294,N_6462);
nand U6704 (N_6704,N_6339,N_6301);
nor U6705 (N_6705,N_6282,N_6291);
nor U6706 (N_6706,N_6301,N_6250);
nand U6707 (N_6707,N_6391,N_6361);
or U6708 (N_6708,N_6321,N_6408);
nand U6709 (N_6709,N_6426,N_6468);
or U6710 (N_6710,N_6447,N_6485);
and U6711 (N_6711,N_6371,N_6259);
xor U6712 (N_6712,N_6368,N_6277);
and U6713 (N_6713,N_6473,N_6338);
xor U6714 (N_6714,N_6319,N_6342);
and U6715 (N_6715,N_6393,N_6268);
nand U6716 (N_6716,N_6444,N_6377);
xnor U6717 (N_6717,N_6268,N_6457);
xor U6718 (N_6718,N_6278,N_6341);
nand U6719 (N_6719,N_6438,N_6261);
and U6720 (N_6720,N_6267,N_6400);
nand U6721 (N_6721,N_6489,N_6372);
nor U6722 (N_6722,N_6292,N_6335);
or U6723 (N_6723,N_6354,N_6250);
and U6724 (N_6724,N_6310,N_6334);
or U6725 (N_6725,N_6302,N_6296);
or U6726 (N_6726,N_6294,N_6492);
or U6727 (N_6727,N_6301,N_6285);
nor U6728 (N_6728,N_6427,N_6354);
or U6729 (N_6729,N_6496,N_6392);
and U6730 (N_6730,N_6336,N_6272);
nand U6731 (N_6731,N_6448,N_6313);
or U6732 (N_6732,N_6427,N_6314);
or U6733 (N_6733,N_6390,N_6434);
nor U6734 (N_6734,N_6459,N_6472);
xor U6735 (N_6735,N_6446,N_6264);
nor U6736 (N_6736,N_6390,N_6418);
nor U6737 (N_6737,N_6352,N_6365);
or U6738 (N_6738,N_6260,N_6374);
xor U6739 (N_6739,N_6492,N_6439);
xor U6740 (N_6740,N_6351,N_6395);
or U6741 (N_6741,N_6413,N_6369);
xor U6742 (N_6742,N_6476,N_6401);
xnor U6743 (N_6743,N_6258,N_6433);
nand U6744 (N_6744,N_6411,N_6467);
nand U6745 (N_6745,N_6294,N_6428);
nand U6746 (N_6746,N_6453,N_6261);
or U6747 (N_6747,N_6257,N_6321);
or U6748 (N_6748,N_6486,N_6257);
nor U6749 (N_6749,N_6385,N_6279);
nand U6750 (N_6750,N_6714,N_6696);
and U6751 (N_6751,N_6574,N_6643);
or U6752 (N_6752,N_6600,N_6688);
or U6753 (N_6753,N_6588,N_6673);
nand U6754 (N_6754,N_6505,N_6630);
and U6755 (N_6755,N_6544,N_6517);
xnor U6756 (N_6756,N_6741,N_6685);
and U6757 (N_6757,N_6732,N_6611);
xnor U6758 (N_6758,N_6651,N_6746);
nand U6759 (N_6759,N_6536,N_6649);
xor U6760 (N_6760,N_6698,N_6516);
nor U6761 (N_6761,N_6690,N_6532);
and U6762 (N_6762,N_6653,N_6676);
nand U6763 (N_6763,N_6557,N_6576);
or U6764 (N_6764,N_6697,N_6580);
xnor U6765 (N_6765,N_6632,N_6612);
xnor U6766 (N_6766,N_6527,N_6603);
nand U6767 (N_6767,N_6682,N_6736);
nor U6768 (N_6768,N_6601,N_6669);
xnor U6769 (N_6769,N_6569,N_6507);
nor U6770 (N_6770,N_6738,N_6726);
or U6771 (N_6771,N_6559,N_6512);
nor U6772 (N_6772,N_6558,N_6594);
nand U6773 (N_6773,N_6735,N_6729);
or U6774 (N_6774,N_6706,N_6589);
and U6775 (N_6775,N_6618,N_6679);
nor U6776 (N_6776,N_6502,N_6662);
and U6777 (N_6777,N_6657,N_6519);
xnor U6778 (N_6778,N_6501,N_6522);
and U6779 (N_6779,N_6724,N_6587);
xnor U6780 (N_6780,N_6638,N_6704);
and U6781 (N_6781,N_6709,N_6530);
or U6782 (N_6782,N_6528,N_6712);
or U6783 (N_6783,N_6586,N_6565);
and U6784 (N_6784,N_6699,N_6675);
or U6785 (N_6785,N_6607,N_6547);
xnor U6786 (N_6786,N_6645,N_6624);
xnor U6787 (N_6787,N_6731,N_6694);
and U6788 (N_6788,N_6553,N_6680);
nand U6789 (N_6789,N_6610,N_6743);
xor U6790 (N_6790,N_6693,N_6566);
xor U6791 (N_6791,N_6560,N_6717);
or U6792 (N_6792,N_6652,N_6552);
nor U6793 (N_6793,N_6633,N_6689);
nor U6794 (N_6794,N_6748,N_6615);
xnor U6795 (N_6795,N_6551,N_6749);
or U6796 (N_6796,N_6556,N_6523);
xnor U6797 (N_6797,N_6713,N_6681);
and U6798 (N_6798,N_6616,N_6504);
xor U6799 (N_6799,N_6708,N_6617);
nand U6800 (N_6800,N_6641,N_6684);
xor U6801 (N_6801,N_6639,N_6613);
nor U6802 (N_6802,N_6526,N_6664);
nor U6803 (N_6803,N_6578,N_6722);
nand U6804 (N_6804,N_6604,N_6570);
xor U6805 (N_6805,N_6625,N_6614);
or U6806 (N_6806,N_6668,N_6591);
nor U6807 (N_6807,N_6564,N_6609);
and U6808 (N_6808,N_6718,N_6503);
nand U6809 (N_6809,N_6647,N_6514);
and U6810 (N_6810,N_6535,N_6597);
nor U6811 (N_6811,N_6703,N_6571);
xnor U6812 (N_6812,N_6555,N_6747);
xnor U6813 (N_6813,N_6602,N_6642);
nor U6814 (N_6814,N_6742,N_6541);
nand U6815 (N_6815,N_6695,N_6648);
xor U6816 (N_6816,N_6734,N_6740);
xnor U6817 (N_6817,N_6672,N_6744);
nor U6818 (N_6818,N_6721,N_6581);
nand U6819 (N_6819,N_6521,N_6691);
and U6820 (N_6820,N_6575,N_6550);
and U6821 (N_6821,N_6739,N_6542);
xor U6822 (N_6822,N_6733,N_6562);
and U6823 (N_6823,N_6595,N_6592);
or U6824 (N_6824,N_6661,N_6646);
or U6825 (N_6825,N_6593,N_6692);
nor U6826 (N_6826,N_6656,N_6660);
nand U6827 (N_6827,N_6678,N_6666);
xnor U6828 (N_6828,N_6723,N_6687);
xnor U6829 (N_6829,N_6534,N_6508);
nor U6830 (N_6830,N_6515,N_6710);
nor U6831 (N_6831,N_6537,N_6650);
xnor U6832 (N_6832,N_6658,N_6719);
nand U6833 (N_6833,N_6640,N_6520);
and U6834 (N_6834,N_6509,N_6631);
and U6835 (N_6835,N_6577,N_6671);
or U6836 (N_6836,N_6540,N_6525);
or U6837 (N_6837,N_6572,N_6590);
nor U6838 (N_6838,N_6511,N_6619);
nand U6839 (N_6839,N_6725,N_6582);
xor U6840 (N_6840,N_6513,N_6626);
or U6841 (N_6841,N_6677,N_6629);
nor U6842 (N_6842,N_6711,N_6545);
nand U6843 (N_6843,N_6644,N_6573);
xnor U6844 (N_6844,N_6727,N_6599);
nand U6845 (N_6845,N_6605,N_6524);
xnor U6846 (N_6846,N_6655,N_6745);
nor U6847 (N_6847,N_6554,N_6715);
nor U6848 (N_6848,N_6728,N_6634);
xor U6849 (N_6849,N_6659,N_6636);
nor U6850 (N_6850,N_6567,N_6546);
xor U6851 (N_6851,N_6683,N_6548);
or U6852 (N_6852,N_6539,N_6533);
and U6853 (N_6853,N_6702,N_6596);
and U6854 (N_6854,N_6500,N_6620);
nor U6855 (N_6855,N_6737,N_6510);
or U6856 (N_6856,N_6720,N_6707);
nand U6857 (N_6857,N_6623,N_6583);
or U6858 (N_6858,N_6579,N_6716);
nor U6859 (N_6859,N_6621,N_6531);
nor U6860 (N_6860,N_6518,N_6598);
or U6861 (N_6861,N_6563,N_6538);
or U6862 (N_6862,N_6730,N_6686);
and U6863 (N_6863,N_6529,N_6561);
nor U6864 (N_6864,N_6670,N_6608);
nor U6865 (N_6865,N_6568,N_6663);
nor U6866 (N_6866,N_6543,N_6674);
nor U6867 (N_6867,N_6584,N_6506);
or U6868 (N_6868,N_6700,N_6585);
nor U6869 (N_6869,N_6667,N_6701);
nand U6870 (N_6870,N_6705,N_6665);
nand U6871 (N_6871,N_6637,N_6606);
and U6872 (N_6872,N_6627,N_6635);
or U6873 (N_6873,N_6654,N_6549);
xnor U6874 (N_6874,N_6622,N_6628);
and U6875 (N_6875,N_6635,N_6638);
nand U6876 (N_6876,N_6680,N_6591);
xor U6877 (N_6877,N_6731,N_6535);
and U6878 (N_6878,N_6636,N_6511);
and U6879 (N_6879,N_6541,N_6608);
or U6880 (N_6880,N_6693,N_6740);
nand U6881 (N_6881,N_6619,N_6679);
xnor U6882 (N_6882,N_6503,N_6527);
nand U6883 (N_6883,N_6694,N_6636);
nand U6884 (N_6884,N_6525,N_6635);
xnor U6885 (N_6885,N_6588,N_6721);
xor U6886 (N_6886,N_6632,N_6667);
nor U6887 (N_6887,N_6582,N_6577);
xnor U6888 (N_6888,N_6632,N_6684);
nor U6889 (N_6889,N_6736,N_6735);
xnor U6890 (N_6890,N_6501,N_6731);
nand U6891 (N_6891,N_6749,N_6651);
nand U6892 (N_6892,N_6588,N_6675);
and U6893 (N_6893,N_6633,N_6563);
or U6894 (N_6894,N_6676,N_6638);
xor U6895 (N_6895,N_6742,N_6645);
or U6896 (N_6896,N_6748,N_6646);
nand U6897 (N_6897,N_6711,N_6697);
nor U6898 (N_6898,N_6586,N_6674);
nor U6899 (N_6899,N_6656,N_6611);
and U6900 (N_6900,N_6740,N_6514);
nand U6901 (N_6901,N_6657,N_6608);
or U6902 (N_6902,N_6676,N_6533);
nor U6903 (N_6903,N_6639,N_6654);
xor U6904 (N_6904,N_6593,N_6670);
nor U6905 (N_6905,N_6700,N_6514);
xor U6906 (N_6906,N_6596,N_6591);
nor U6907 (N_6907,N_6521,N_6745);
or U6908 (N_6908,N_6694,N_6656);
xor U6909 (N_6909,N_6603,N_6594);
nand U6910 (N_6910,N_6667,N_6631);
nand U6911 (N_6911,N_6582,N_6673);
and U6912 (N_6912,N_6693,N_6602);
and U6913 (N_6913,N_6713,N_6731);
nor U6914 (N_6914,N_6511,N_6748);
xnor U6915 (N_6915,N_6714,N_6710);
nand U6916 (N_6916,N_6536,N_6544);
and U6917 (N_6917,N_6560,N_6687);
xnor U6918 (N_6918,N_6658,N_6559);
nor U6919 (N_6919,N_6657,N_6652);
nor U6920 (N_6920,N_6662,N_6505);
nand U6921 (N_6921,N_6624,N_6655);
xor U6922 (N_6922,N_6727,N_6600);
nor U6923 (N_6923,N_6515,N_6525);
and U6924 (N_6924,N_6691,N_6510);
and U6925 (N_6925,N_6684,N_6725);
nand U6926 (N_6926,N_6554,N_6584);
nand U6927 (N_6927,N_6582,N_6708);
xor U6928 (N_6928,N_6648,N_6608);
nor U6929 (N_6929,N_6691,N_6623);
xor U6930 (N_6930,N_6563,N_6672);
nor U6931 (N_6931,N_6588,N_6728);
nor U6932 (N_6932,N_6691,N_6683);
and U6933 (N_6933,N_6731,N_6724);
or U6934 (N_6934,N_6558,N_6579);
xnor U6935 (N_6935,N_6642,N_6671);
or U6936 (N_6936,N_6626,N_6520);
or U6937 (N_6937,N_6721,N_6548);
or U6938 (N_6938,N_6622,N_6726);
and U6939 (N_6939,N_6560,N_6574);
nand U6940 (N_6940,N_6644,N_6601);
and U6941 (N_6941,N_6524,N_6552);
or U6942 (N_6942,N_6512,N_6541);
xor U6943 (N_6943,N_6724,N_6607);
xor U6944 (N_6944,N_6722,N_6726);
xor U6945 (N_6945,N_6742,N_6649);
xnor U6946 (N_6946,N_6727,N_6711);
nand U6947 (N_6947,N_6549,N_6724);
xor U6948 (N_6948,N_6628,N_6509);
nor U6949 (N_6949,N_6667,N_6669);
nor U6950 (N_6950,N_6562,N_6701);
or U6951 (N_6951,N_6682,N_6654);
and U6952 (N_6952,N_6561,N_6632);
and U6953 (N_6953,N_6578,N_6737);
nand U6954 (N_6954,N_6748,N_6602);
xor U6955 (N_6955,N_6673,N_6577);
nor U6956 (N_6956,N_6697,N_6530);
nand U6957 (N_6957,N_6652,N_6672);
nand U6958 (N_6958,N_6621,N_6727);
xor U6959 (N_6959,N_6531,N_6709);
nand U6960 (N_6960,N_6549,N_6558);
or U6961 (N_6961,N_6510,N_6613);
xnor U6962 (N_6962,N_6612,N_6618);
or U6963 (N_6963,N_6577,N_6590);
xnor U6964 (N_6964,N_6699,N_6715);
or U6965 (N_6965,N_6526,N_6670);
nor U6966 (N_6966,N_6535,N_6713);
xor U6967 (N_6967,N_6655,N_6525);
xnor U6968 (N_6968,N_6609,N_6542);
and U6969 (N_6969,N_6588,N_6625);
and U6970 (N_6970,N_6598,N_6712);
nor U6971 (N_6971,N_6594,N_6676);
nor U6972 (N_6972,N_6522,N_6659);
xor U6973 (N_6973,N_6560,N_6679);
nand U6974 (N_6974,N_6725,N_6591);
nor U6975 (N_6975,N_6697,N_6651);
or U6976 (N_6976,N_6730,N_6734);
and U6977 (N_6977,N_6668,N_6677);
nor U6978 (N_6978,N_6739,N_6680);
and U6979 (N_6979,N_6681,N_6737);
xor U6980 (N_6980,N_6617,N_6567);
and U6981 (N_6981,N_6523,N_6532);
nand U6982 (N_6982,N_6568,N_6675);
nor U6983 (N_6983,N_6567,N_6669);
xor U6984 (N_6984,N_6562,N_6672);
nand U6985 (N_6985,N_6570,N_6631);
and U6986 (N_6986,N_6680,N_6707);
nor U6987 (N_6987,N_6575,N_6647);
or U6988 (N_6988,N_6749,N_6573);
or U6989 (N_6989,N_6590,N_6729);
xnor U6990 (N_6990,N_6680,N_6512);
or U6991 (N_6991,N_6606,N_6578);
and U6992 (N_6992,N_6530,N_6644);
nor U6993 (N_6993,N_6504,N_6587);
or U6994 (N_6994,N_6703,N_6590);
or U6995 (N_6995,N_6715,N_6716);
or U6996 (N_6996,N_6580,N_6530);
or U6997 (N_6997,N_6671,N_6520);
nor U6998 (N_6998,N_6723,N_6600);
nor U6999 (N_6999,N_6739,N_6527);
nor U7000 (N_7000,N_6996,N_6955);
nand U7001 (N_7001,N_6891,N_6991);
and U7002 (N_7002,N_6956,N_6840);
nor U7003 (N_7003,N_6819,N_6757);
and U7004 (N_7004,N_6963,N_6990);
nand U7005 (N_7005,N_6874,N_6782);
nand U7006 (N_7006,N_6947,N_6865);
or U7007 (N_7007,N_6964,N_6787);
or U7008 (N_7008,N_6952,N_6982);
xor U7009 (N_7009,N_6841,N_6784);
nor U7010 (N_7010,N_6950,N_6892);
nand U7011 (N_7011,N_6870,N_6960);
xnor U7012 (N_7012,N_6910,N_6808);
and U7013 (N_7013,N_6820,N_6814);
nor U7014 (N_7014,N_6771,N_6863);
and U7015 (N_7015,N_6926,N_6922);
nor U7016 (N_7016,N_6998,N_6989);
xor U7017 (N_7017,N_6920,N_6951);
or U7018 (N_7018,N_6916,N_6761);
and U7019 (N_7019,N_6795,N_6961);
or U7020 (N_7020,N_6766,N_6908);
xnor U7021 (N_7021,N_6978,N_6890);
xnor U7022 (N_7022,N_6983,N_6842);
and U7023 (N_7023,N_6886,N_6853);
nor U7024 (N_7024,N_6806,N_6867);
and U7025 (N_7025,N_6792,N_6753);
nand U7026 (N_7026,N_6793,N_6826);
or U7027 (N_7027,N_6958,N_6941);
and U7028 (N_7028,N_6872,N_6830);
xnor U7029 (N_7029,N_6929,N_6932);
and U7030 (N_7030,N_6786,N_6828);
nor U7031 (N_7031,N_6860,N_6946);
xor U7032 (N_7032,N_6760,N_6871);
xor U7033 (N_7033,N_6827,N_6781);
nand U7034 (N_7034,N_6977,N_6949);
or U7035 (N_7035,N_6931,N_6809);
xor U7036 (N_7036,N_6822,N_6918);
xnor U7037 (N_7037,N_6783,N_6899);
nor U7038 (N_7038,N_6804,N_6843);
nand U7039 (N_7039,N_6992,N_6844);
or U7040 (N_7040,N_6759,N_6852);
xor U7041 (N_7041,N_6751,N_6770);
nor U7042 (N_7042,N_6923,N_6758);
or U7043 (N_7043,N_6796,N_6925);
nand U7044 (N_7044,N_6815,N_6881);
or U7045 (N_7045,N_6954,N_6911);
nand U7046 (N_7046,N_6778,N_6772);
nand U7047 (N_7047,N_6893,N_6845);
xor U7048 (N_7048,N_6837,N_6797);
nand U7049 (N_7049,N_6868,N_6934);
and U7050 (N_7050,N_6810,N_6805);
or U7051 (N_7051,N_6789,N_6776);
and U7052 (N_7052,N_6988,N_6930);
nor U7053 (N_7053,N_6856,N_6769);
nand U7054 (N_7054,N_6875,N_6833);
xor U7055 (N_7055,N_6948,N_6777);
nor U7056 (N_7056,N_6773,N_6942);
or U7057 (N_7057,N_6879,N_6905);
xnor U7058 (N_7058,N_6834,N_6913);
or U7059 (N_7059,N_6752,N_6800);
xor U7060 (N_7060,N_6903,N_6900);
xor U7061 (N_7061,N_6953,N_6980);
nand U7062 (N_7062,N_6972,N_6799);
or U7063 (N_7063,N_6854,N_6775);
nand U7064 (N_7064,N_6921,N_6851);
nand U7065 (N_7065,N_6801,N_6817);
nand U7066 (N_7066,N_6885,N_6866);
nor U7067 (N_7067,N_6750,N_6968);
and U7068 (N_7068,N_6807,N_6975);
xor U7069 (N_7069,N_6979,N_6894);
and U7070 (N_7070,N_6765,N_6970);
nor U7071 (N_7071,N_6764,N_6887);
nor U7072 (N_7072,N_6888,N_6829);
or U7073 (N_7073,N_6962,N_6816);
xor U7074 (N_7074,N_6974,N_6993);
and U7075 (N_7075,N_6754,N_6987);
or U7076 (N_7076,N_6882,N_6780);
and U7077 (N_7077,N_6973,N_6902);
nor U7078 (N_7078,N_6914,N_6994);
or U7079 (N_7079,N_6901,N_6861);
xnor U7080 (N_7080,N_6763,N_6984);
nor U7081 (N_7081,N_6924,N_6848);
nand U7082 (N_7082,N_6896,N_6825);
nor U7083 (N_7083,N_6944,N_6909);
and U7084 (N_7084,N_6859,N_6847);
nor U7085 (N_7085,N_6966,N_6767);
nor U7086 (N_7086,N_6755,N_6971);
xnor U7087 (N_7087,N_6768,N_6936);
or U7088 (N_7088,N_6774,N_6876);
and U7089 (N_7089,N_6821,N_6981);
or U7090 (N_7090,N_6836,N_6928);
nand U7091 (N_7091,N_6937,N_6938);
xnor U7092 (N_7092,N_6855,N_6785);
xnor U7093 (N_7093,N_6985,N_6864);
nand U7094 (N_7094,N_6917,N_6823);
or U7095 (N_7095,N_6945,N_6790);
and U7096 (N_7096,N_6846,N_6940);
and U7097 (N_7097,N_6791,N_6884);
nor U7098 (N_7098,N_6798,N_6959);
nand U7099 (N_7099,N_6933,N_6831);
and U7100 (N_7100,N_6832,N_6898);
nand U7101 (N_7101,N_6907,N_6862);
nand U7102 (N_7102,N_6835,N_6927);
xnor U7103 (N_7103,N_6995,N_6997);
nand U7104 (N_7104,N_6897,N_6858);
and U7105 (N_7105,N_6802,N_6873);
and U7106 (N_7106,N_6986,N_6813);
xnor U7107 (N_7107,N_6880,N_6919);
nor U7108 (N_7108,N_6912,N_6965);
and U7109 (N_7109,N_6779,N_6969);
xor U7110 (N_7110,N_6915,N_6906);
nor U7111 (N_7111,N_6803,N_6999);
and U7112 (N_7112,N_6839,N_6943);
nand U7113 (N_7113,N_6878,N_6857);
or U7114 (N_7114,N_6976,N_6824);
nand U7115 (N_7115,N_6788,N_6849);
nand U7116 (N_7116,N_6756,N_6811);
and U7117 (N_7117,N_6869,N_6967);
nand U7118 (N_7118,N_6939,N_6850);
nor U7119 (N_7119,N_6957,N_6883);
nand U7120 (N_7120,N_6794,N_6935);
nor U7121 (N_7121,N_6762,N_6895);
nor U7122 (N_7122,N_6818,N_6838);
and U7123 (N_7123,N_6889,N_6812);
and U7124 (N_7124,N_6904,N_6877);
xor U7125 (N_7125,N_6976,N_6845);
and U7126 (N_7126,N_6926,N_6793);
nand U7127 (N_7127,N_6928,N_6900);
xor U7128 (N_7128,N_6927,N_6996);
nand U7129 (N_7129,N_6830,N_6867);
nand U7130 (N_7130,N_6944,N_6893);
or U7131 (N_7131,N_6885,N_6868);
nor U7132 (N_7132,N_6930,N_6952);
nor U7133 (N_7133,N_6874,N_6866);
nand U7134 (N_7134,N_6974,N_6808);
or U7135 (N_7135,N_6790,N_6932);
nand U7136 (N_7136,N_6937,N_6840);
or U7137 (N_7137,N_6930,N_6804);
nand U7138 (N_7138,N_6801,N_6815);
nand U7139 (N_7139,N_6825,N_6861);
nand U7140 (N_7140,N_6760,N_6866);
nor U7141 (N_7141,N_6966,N_6984);
or U7142 (N_7142,N_6939,N_6889);
nand U7143 (N_7143,N_6752,N_6986);
and U7144 (N_7144,N_6856,N_6874);
or U7145 (N_7145,N_6996,N_6869);
and U7146 (N_7146,N_6755,N_6939);
nor U7147 (N_7147,N_6750,N_6893);
or U7148 (N_7148,N_6905,N_6872);
and U7149 (N_7149,N_6956,N_6944);
xor U7150 (N_7150,N_6832,N_6965);
or U7151 (N_7151,N_6896,N_6830);
nor U7152 (N_7152,N_6785,N_6942);
or U7153 (N_7153,N_6790,N_6900);
and U7154 (N_7154,N_6767,N_6934);
xor U7155 (N_7155,N_6935,N_6912);
xnor U7156 (N_7156,N_6884,N_6801);
and U7157 (N_7157,N_6783,N_6859);
xor U7158 (N_7158,N_6842,N_6947);
nand U7159 (N_7159,N_6875,N_6759);
nor U7160 (N_7160,N_6803,N_6902);
and U7161 (N_7161,N_6907,N_6754);
and U7162 (N_7162,N_6908,N_6777);
nor U7163 (N_7163,N_6842,N_6775);
nor U7164 (N_7164,N_6811,N_6829);
xnor U7165 (N_7165,N_6860,N_6897);
or U7166 (N_7166,N_6997,N_6855);
nor U7167 (N_7167,N_6966,N_6922);
nand U7168 (N_7168,N_6962,N_6760);
and U7169 (N_7169,N_6845,N_6996);
and U7170 (N_7170,N_6956,N_6895);
nor U7171 (N_7171,N_6866,N_6838);
xnor U7172 (N_7172,N_6817,N_6974);
nor U7173 (N_7173,N_6781,N_6884);
nand U7174 (N_7174,N_6894,N_6795);
and U7175 (N_7175,N_6862,N_6838);
and U7176 (N_7176,N_6769,N_6786);
nor U7177 (N_7177,N_6966,N_6963);
and U7178 (N_7178,N_6999,N_6858);
xnor U7179 (N_7179,N_6794,N_6768);
nand U7180 (N_7180,N_6893,N_6979);
or U7181 (N_7181,N_6805,N_6893);
or U7182 (N_7182,N_6824,N_6832);
nand U7183 (N_7183,N_6806,N_6941);
and U7184 (N_7184,N_6976,N_6933);
nand U7185 (N_7185,N_6985,N_6852);
xnor U7186 (N_7186,N_6776,N_6994);
and U7187 (N_7187,N_6983,N_6922);
and U7188 (N_7188,N_6876,N_6967);
or U7189 (N_7189,N_6929,N_6817);
or U7190 (N_7190,N_6912,N_6765);
and U7191 (N_7191,N_6863,N_6995);
xnor U7192 (N_7192,N_6800,N_6889);
xnor U7193 (N_7193,N_6850,N_6775);
and U7194 (N_7194,N_6771,N_6793);
or U7195 (N_7195,N_6911,N_6777);
nand U7196 (N_7196,N_6987,N_6753);
and U7197 (N_7197,N_6807,N_6799);
and U7198 (N_7198,N_6833,N_6867);
or U7199 (N_7199,N_6753,N_6763);
nand U7200 (N_7200,N_6933,N_6999);
and U7201 (N_7201,N_6931,N_6924);
or U7202 (N_7202,N_6774,N_6753);
nor U7203 (N_7203,N_6851,N_6880);
nand U7204 (N_7204,N_6836,N_6939);
or U7205 (N_7205,N_6878,N_6796);
nor U7206 (N_7206,N_6844,N_6841);
xor U7207 (N_7207,N_6986,N_6917);
nand U7208 (N_7208,N_6993,N_6936);
nand U7209 (N_7209,N_6937,N_6873);
nor U7210 (N_7210,N_6790,N_6981);
and U7211 (N_7211,N_6790,N_6824);
nor U7212 (N_7212,N_6750,N_6905);
or U7213 (N_7213,N_6838,N_6881);
nand U7214 (N_7214,N_6880,N_6909);
or U7215 (N_7215,N_6796,N_6896);
and U7216 (N_7216,N_6798,N_6788);
nand U7217 (N_7217,N_6887,N_6766);
nor U7218 (N_7218,N_6783,N_6768);
and U7219 (N_7219,N_6794,N_6802);
and U7220 (N_7220,N_6861,N_6992);
nand U7221 (N_7221,N_6809,N_6913);
nor U7222 (N_7222,N_6873,N_6952);
or U7223 (N_7223,N_6912,N_6992);
nand U7224 (N_7224,N_6912,N_6767);
and U7225 (N_7225,N_6874,N_6832);
nand U7226 (N_7226,N_6911,N_6985);
or U7227 (N_7227,N_6899,N_6901);
or U7228 (N_7228,N_6934,N_6967);
nor U7229 (N_7229,N_6883,N_6959);
nor U7230 (N_7230,N_6964,N_6911);
or U7231 (N_7231,N_6995,N_6981);
nor U7232 (N_7232,N_6843,N_6854);
nor U7233 (N_7233,N_6790,N_6876);
xor U7234 (N_7234,N_6986,N_6844);
nor U7235 (N_7235,N_6888,N_6989);
and U7236 (N_7236,N_6838,N_6904);
or U7237 (N_7237,N_6831,N_6930);
and U7238 (N_7238,N_6935,N_6915);
xnor U7239 (N_7239,N_6869,N_6795);
nand U7240 (N_7240,N_6999,N_6945);
nand U7241 (N_7241,N_6800,N_6883);
and U7242 (N_7242,N_6967,N_6765);
xnor U7243 (N_7243,N_6938,N_6869);
or U7244 (N_7244,N_6894,N_6987);
nand U7245 (N_7245,N_6973,N_6753);
nand U7246 (N_7246,N_6846,N_6990);
nor U7247 (N_7247,N_6822,N_6832);
nand U7248 (N_7248,N_6902,N_6826);
xnor U7249 (N_7249,N_6811,N_6953);
nand U7250 (N_7250,N_7104,N_7034);
nor U7251 (N_7251,N_7037,N_7185);
and U7252 (N_7252,N_7144,N_7049);
and U7253 (N_7253,N_7113,N_7089);
nand U7254 (N_7254,N_7236,N_7002);
nand U7255 (N_7255,N_7217,N_7135);
nor U7256 (N_7256,N_7241,N_7150);
nand U7257 (N_7257,N_7181,N_7030);
nand U7258 (N_7258,N_7134,N_7159);
nor U7259 (N_7259,N_7069,N_7022);
and U7260 (N_7260,N_7175,N_7248);
nand U7261 (N_7261,N_7023,N_7087);
or U7262 (N_7262,N_7059,N_7109);
nand U7263 (N_7263,N_7006,N_7190);
and U7264 (N_7264,N_7077,N_7208);
xor U7265 (N_7265,N_7133,N_7053);
nand U7266 (N_7266,N_7029,N_7076);
and U7267 (N_7267,N_7170,N_7165);
and U7268 (N_7268,N_7106,N_7005);
nand U7269 (N_7269,N_7176,N_7224);
nand U7270 (N_7270,N_7240,N_7148);
nand U7271 (N_7271,N_7244,N_7167);
or U7272 (N_7272,N_7136,N_7228);
xnor U7273 (N_7273,N_7163,N_7040);
or U7274 (N_7274,N_7225,N_7179);
or U7275 (N_7275,N_7213,N_7050);
xor U7276 (N_7276,N_7191,N_7085);
nand U7277 (N_7277,N_7214,N_7079);
nand U7278 (N_7278,N_7035,N_7239);
and U7279 (N_7279,N_7245,N_7215);
xor U7280 (N_7280,N_7147,N_7220);
nor U7281 (N_7281,N_7070,N_7007);
nand U7282 (N_7282,N_7108,N_7010);
nor U7283 (N_7283,N_7116,N_7102);
xnor U7284 (N_7284,N_7209,N_7160);
nand U7285 (N_7285,N_7041,N_7054);
nand U7286 (N_7286,N_7008,N_7092);
nand U7287 (N_7287,N_7161,N_7099);
nand U7288 (N_7288,N_7201,N_7025);
nand U7289 (N_7289,N_7074,N_7200);
nor U7290 (N_7290,N_7098,N_7062);
nand U7291 (N_7291,N_7067,N_7157);
or U7292 (N_7292,N_7166,N_7028);
and U7293 (N_7293,N_7186,N_7064);
nor U7294 (N_7294,N_7122,N_7171);
and U7295 (N_7295,N_7233,N_7036);
xnor U7296 (N_7296,N_7048,N_7212);
xnor U7297 (N_7297,N_7111,N_7055);
or U7298 (N_7298,N_7097,N_7203);
nand U7299 (N_7299,N_7207,N_7078);
xor U7300 (N_7300,N_7012,N_7145);
nand U7301 (N_7301,N_7105,N_7218);
xor U7302 (N_7302,N_7221,N_7013);
and U7303 (N_7303,N_7047,N_7044);
nand U7304 (N_7304,N_7130,N_7016);
nand U7305 (N_7305,N_7032,N_7095);
xnor U7306 (N_7306,N_7014,N_7018);
or U7307 (N_7307,N_7011,N_7121);
xor U7308 (N_7308,N_7232,N_7198);
nor U7309 (N_7309,N_7229,N_7138);
nand U7310 (N_7310,N_7088,N_7183);
or U7311 (N_7311,N_7158,N_7020);
nor U7312 (N_7312,N_7019,N_7177);
xor U7313 (N_7313,N_7107,N_7066);
and U7314 (N_7314,N_7132,N_7249);
or U7315 (N_7315,N_7091,N_7237);
xor U7316 (N_7316,N_7180,N_7100);
nand U7317 (N_7317,N_7045,N_7120);
and U7318 (N_7318,N_7103,N_7112);
nor U7319 (N_7319,N_7182,N_7126);
or U7320 (N_7320,N_7151,N_7242);
nand U7321 (N_7321,N_7184,N_7068);
or U7322 (N_7322,N_7216,N_7004);
nand U7323 (N_7323,N_7204,N_7247);
nand U7324 (N_7324,N_7139,N_7093);
or U7325 (N_7325,N_7154,N_7082);
nor U7326 (N_7326,N_7071,N_7058);
or U7327 (N_7327,N_7114,N_7231);
and U7328 (N_7328,N_7046,N_7075);
nand U7329 (N_7329,N_7131,N_7061);
xor U7330 (N_7330,N_7003,N_7235);
xnor U7331 (N_7331,N_7189,N_7063);
or U7332 (N_7332,N_7129,N_7118);
xnor U7333 (N_7333,N_7033,N_7057);
or U7334 (N_7334,N_7015,N_7024);
or U7335 (N_7335,N_7192,N_7195);
xor U7336 (N_7336,N_7060,N_7199);
xnor U7337 (N_7337,N_7031,N_7172);
and U7338 (N_7338,N_7110,N_7205);
nor U7339 (N_7339,N_7065,N_7042);
xnor U7340 (N_7340,N_7234,N_7178);
and U7341 (N_7341,N_7123,N_7021);
nor U7342 (N_7342,N_7127,N_7238);
xor U7343 (N_7343,N_7083,N_7197);
xor U7344 (N_7344,N_7039,N_7153);
xor U7345 (N_7345,N_7096,N_7230);
xnor U7346 (N_7346,N_7017,N_7117);
or U7347 (N_7347,N_7219,N_7149);
nor U7348 (N_7348,N_7094,N_7187);
and U7349 (N_7349,N_7227,N_7115);
or U7350 (N_7350,N_7128,N_7156);
xor U7351 (N_7351,N_7223,N_7152);
xnor U7352 (N_7352,N_7169,N_7090);
or U7353 (N_7353,N_7222,N_7211);
and U7354 (N_7354,N_7246,N_7137);
nand U7355 (N_7355,N_7226,N_7026);
nor U7356 (N_7356,N_7101,N_7140);
or U7357 (N_7357,N_7125,N_7164);
nand U7358 (N_7358,N_7146,N_7124);
or U7359 (N_7359,N_7202,N_7196);
nand U7360 (N_7360,N_7056,N_7174);
or U7361 (N_7361,N_7173,N_7141);
nand U7362 (N_7362,N_7142,N_7168);
or U7363 (N_7363,N_7072,N_7043);
nor U7364 (N_7364,N_7081,N_7155);
nor U7365 (N_7365,N_7073,N_7210);
or U7366 (N_7366,N_7193,N_7243);
or U7367 (N_7367,N_7143,N_7051);
nand U7368 (N_7368,N_7038,N_7052);
nor U7369 (N_7369,N_7001,N_7188);
nand U7370 (N_7370,N_7080,N_7206);
xnor U7371 (N_7371,N_7000,N_7027);
nand U7372 (N_7372,N_7119,N_7009);
nand U7373 (N_7373,N_7086,N_7194);
nor U7374 (N_7374,N_7084,N_7162);
nor U7375 (N_7375,N_7046,N_7119);
xnor U7376 (N_7376,N_7039,N_7151);
and U7377 (N_7377,N_7141,N_7067);
xor U7378 (N_7378,N_7121,N_7101);
nor U7379 (N_7379,N_7218,N_7180);
xnor U7380 (N_7380,N_7183,N_7070);
or U7381 (N_7381,N_7243,N_7196);
and U7382 (N_7382,N_7151,N_7188);
or U7383 (N_7383,N_7124,N_7155);
xor U7384 (N_7384,N_7109,N_7183);
nor U7385 (N_7385,N_7041,N_7153);
or U7386 (N_7386,N_7122,N_7066);
and U7387 (N_7387,N_7112,N_7120);
or U7388 (N_7388,N_7104,N_7236);
xor U7389 (N_7389,N_7224,N_7119);
and U7390 (N_7390,N_7182,N_7052);
and U7391 (N_7391,N_7001,N_7074);
and U7392 (N_7392,N_7162,N_7033);
nand U7393 (N_7393,N_7080,N_7126);
xor U7394 (N_7394,N_7052,N_7024);
xor U7395 (N_7395,N_7001,N_7206);
or U7396 (N_7396,N_7226,N_7213);
nor U7397 (N_7397,N_7137,N_7231);
xor U7398 (N_7398,N_7175,N_7238);
nor U7399 (N_7399,N_7171,N_7199);
or U7400 (N_7400,N_7014,N_7096);
nor U7401 (N_7401,N_7062,N_7110);
and U7402 (N_7402,N_7163,N_7133);
or U7403 (N_7403,N_7146,N_7151);
and U7404 (N_7404,N_7178,N_7152);
xnor U7405 (N_7405,N_7077,N_7076);
and U7406 (N_7406,N_7037,N_7085);
and U7407 (N_7407,N_7021,N_7146);
and U7408 (N_7408,N_7234,N_7035);
nand U7409 (N_7409,N_7096,N_7005);
nor U7410 (N_7410,N_7156,N_7060);
nor U7411 (N_7411,N_7234,N_7089);
or U7412 (N_7412,N_7214,N_7179);
nor U7413 (N_7413,N_7155,N_7005);
nor U7414 (N_7414,N_7186,N_7148);
or U7415 (N_7415,N_7064,N_7135);
nand U7416 (N_7416,N_7127,N_7204);
nand U7417 (N_7417,N_7154,N_7072);
xor U7418 (N_7418,N_7006,N_7155);
xor U7419 (N_7419,N_7192,N_7079);
or U7420 (N_7420,N_7217,N_7210);
xor U7421 (N_7421,N_7241,N_7042);
nand U7422 (N_7422,N_7087,N_7110);
nand U7423 (N_7423,N_7243,N_7046);
nor U7424 (N_7424,N_7238,N_7036);
xnor U7425 (N_7425,N_7201,N_7077);
xor U7426 (N_7426,N_7231,N_7167);
nor U7427 (N_7427,N_7020,N_7137);
nand U7428 (N_7428,N_7155,N_7118);
and U7429 (N_7429,N_7221,N_7078);
and U7430 (N_7430,N_7064,N_7123);
nand U7431 (N_7431,N_7055,N_7243);
or U7432 (N_7432,N_7065,N_7239);
nor U7433 (N_7433,N_7044,N_7246);
and U7434 (N_7434,N_7082,N_7245);
xor U7435 (N_7435,N_7000,N_7180);
or U7436 (N_7436,N_7146,N_7037);
nor U7437 (N_7437,N_7066,N_7105);
nor U7438 (N_7438,N_7134,N_7139);
xor U7439 (N_7439,N_7151,N_7063);
or U7440 (N_7440,N_7223,N_7084);
xor U7441 (N_7441,N_7248,N_7100);
nand U7442 (N_7442,N_7100,N_7163);
or U7443 (N_7443,N_7078,N_7147);
nand U7444 (N_7444,N_7137,N_7067);
nand U7445 (N_7445,N_7109,N_7078);
xnor U7446 (N_7446,N_7048,N_7116);
or U7447 (N_7447,N_7129,N_7162);
or U7448 (N_7448,N_7013,N_7116);
and U7449 (N_7449,N_7014,N_7147);
or U7450 (N_7450,N_7174,N_7238);
nand U7451 (N_7451,N_7155,N_7059);
or U7452 (N_7452,N_7057,N_7179);
nor U7453 (N_7453,N_7042,N_7184);
xor U7454 (N_7454,N_7015,N_7087);
nand U7455 (N_7455,N_7042,N_7239);
nor U7456 (N_7456,N_7144,N_7186);
nand U7457 (N_7457,N_7188,N_7039);
and U7458 (N_7458,N_7141,N_7113);
nand U7459 (N_7459,N_7057,N_7145);
xor U7460 (N_7460,N_7154,N_7153);
nand U7461 (N_7461,N_7164,N_7067);
xnor U7462 (N_7462,N_7212,N_7183);
nand U7463 (N_7463,N_7058,N_7117);
nand U7464 (N_7464,N_7187,N_7098);
and U7465 (N_7465,N_7181,N_7074);
or U7466 (N_7466,N_7113,N_7184);
xnor U7467 (N_7467,N_7241,N_7248);
and U7468 (N_7468,N_7093,N_7144);
nor U7469 (N_7469,N_7089,N_7172);
nand U7470 (N_7470,N_7215,N_7201);
and U7471 (N_7471,N_7082,N_7065);
nand U7472 (N_7472,N_7231,N_7100);
nor U7473 (N_7473,N_7201,N_7125);
nand U7474 (N_7474,N_7056,N_7249);
xor U7475 (N_7475,N_7085,N_7052);
xnor U7476 (N_7476,N_7181,N_7137);
xor U7477 (N_7477,N_7152,N_7085);
nand U7478 (N_7478,N_7231,N_7084);
xnor U7479 (N_7479,N_7079,N_7136);
or U7480 (N_7480,N_7208,N_7187);
nor U7481 (N_7481,N_7038,N_7081);
xnor U7482 (N_7482,N_7052,N_7071);
or U7483 (N_7483,N_7122,N_7084);
and U7484 (N_7484,N_7144,N_7060);
xor U7485 (N_7485,N_7071,N_7131);
and U7486 (N_7486,N_7009,N_7202);
xor U7487 (N_7487,N_7152,N_7016);
and U7488 (N_7488,N_7024,N_7214);
or U7489 (N_7489,N_7010,N_7205);
and U7490 (N_7490,N_7078,N_7197);
nand U7491 (N_7491,N_7201,N_7039);
xnor U7492 (N_7492,N_7241,N_7080);
nor U7493 (N_7493,N_7034,N_7153);
and U7494 (N_7494,N_7069,N_7210);
xnor U7495 (N_7495,N_7091,N_7047);
nor U7496 (N_7496,N_7009,N_7131);
nand U7497 (N_7497,N_7052,N_7104);
xor U7498 (N_7498,N_7096,N_7114);
and U7499 (N_7499,N_7079,N_7245);
nand U7500 (N_7500,N_7480,N_7465);
and U7501 (N_7501,N_7270,N_7487);
or U7502 (N_7502,N_7316,N_7473);
or U7503 (N_7503,N_7260,N_7392);
nor U7504 (N_7504,N_7351,N_7364);
nand U7505 (N_7505,N_7376,N_7268);
and U7506 (N_7506,N_7464,N_7322);
nor U7507 (N_7507,N_7405,N_7422);
xor U7508 (N_7508,N_7410,N_7475);
and U7509 (N_7509,N_7290,N_7365);
nor U7510 (N_7510,N_7257,N_7263);
nor U7511 (N_7511,N_7252,N_7299);
and U7512 (N_7512,N_7462,N_7324);
or U7513 (N_7513,N_7310,N_7354);
nand U7514 (N_7514,N_7319,N_7467);
xor U7515 (N_7515,N_7417,N_7439);
xor U7516 (N_7516,N_7388,N_7363);
xnor U7517 (N_7517,N_7420,N_7497);
nand U7518 (N_7518,N_7303,N_7336);
or U7519 (N_7519,N_7321,N_7353);
nand U7520 (N_7520,N_7330,N_7343);
nor U7521 (N_7521,N_7483,N_7395);
xnor U7522 (N_7522,N_7424,N_7498);
xor U7523 (N_7523,N_7358,N_7393);
nor U7524 (N_7524,N_7391,N_7261);
and U7525 (N_7525,N_7381,N_7399);
nand U7526 (N_7526,N_7385,N_7367);
xor U7527 (N_7527,N_7470,N_7433);
and U7528 (N_7528,N_7426,N_7412);
nor U7529 (N_7529,N_7409,N_7356);
nor U7530 (N_7530,N_7347,N_7271);
and U7531 (N_7531,N_7423,N_7496);
xor U7532 (N_7532,N_7396,N_7284);
nor U7533 (N_7533,N_7253,N_7281);
nor U7534 (N_7534,N_7489,N_7382);
xor U7535 (N_7535,N_7380,N_7300);
xnor U7536 (N_7536,N_7430,N_7262);
or U7537 (N_7537,N_7461,N_7339);
and U7538 (N_7538,N_7297,N_7397);
nor U7539 (N_7539,N_7312,N_7302);
xor U7540 (N_7540,N_7408,N_7273);
or U7541 (N_7541,N_7334,N_7458);
xor U7542 (N_7542,N_7447,N_7311);
and U7543 (N_7543,N_7349,N_7404);
and U7544 (N_7544,N_7400,N_7411);
or U7545 (N_7545,N_7280,N_7277);
nor U7546 (N_7546,N_7267,N_7377);
and U7547 (N_7547,N_7459,N_7337);
xnor U7548 (N_7548,N_7301,N_7387);
and U7549 (N_7549,N_7373,N_7471);
nand U7550 (N_7550,N_7389,N_7463);
or U7551 (N_7551,N_7272,N_7256);
or U7552 (N_7552,N_7414,N_7278);
and U7553 (N_7553,N_7425,N_7289);
nand U7554 (N_7554,N_7275,N_7350);
or U7555 (N_7555,N_7355,N_7360);
nand U7556 (N_7556,N_7251,N_7352);
xor U7557 (N_7557,N_7384,N_7478);
or U7558 (N_7558,N_7481,N_7394);
xnor U7559 (N_7559,N_7413,N_7383);
and U7560 (N_7560,N_7361,N_7468);
and U7561 (N_7561,N_7269,N_7274);
and U7562 (N_7562,N_7482,N_7366);
nor U7563 (N_7563,N_7402,N_7431);
and U7564 (N_7564,N_7436,N_7437);
nand U7565 (N_7565,N_7443,N_7307);
xnor U7566 (N_7566,N_7315,N_7419);
and U7567 (N_7567,N_7286,N_7466);
or U7568 (N_7568,N_7428,N_7341);
nand U7569 (N_7569,N_7340,N_7288);
xor U7570 (N_7570,N_7308,N_7485);
and U7571 (N_7571,N_7318,N_7492);
nor U7572 (N_7572,N_7305,N_7346);
nand U7573 (N_7573,N_7345,N_7287);
and U7574 (N_7574,N_7294,N_7327);
nor U7575 (N_7575,N_7285,N_7418);
and U7576 (N_7576,N_7460,N_7495);
or U7577 (N_7577,N_7484,N_7452);
xor U7578 (N_7578,N_7313,N_7266);
nand U7579 (N_7579,N_7357,N_7491);
and U7580 (N_7580,N_7429,N_7314);
or U7581 (N_7581,N_7421,N_7333);
nand U7582 (N_7582,N_7292,N_7390);
nor U7583 (N_7583,N_7320,N_7407);
nand U7584 (N_7584,N_7344,N_7317);
and U7585 (N_7585,N_7499,N_7264);
and U7586 (N_7586,N_7276,N_7435);
nand U7587 (N_7587,N_7490,N_7469);
xor U7588 (N_7588,N_7474,N_7374);
or U7589 (N_7589,N_7282,N_7476);
nand U7590 (N_7590,N_7359,N_7304);
or U7591 (N_7591,N_7442,N_7259);
xnor U7592 (N_7592,N_7432,N_7494);
xnor U7593 (N_7593,N_7254,N_7453);
nand U7594 (N_7594,N_7454,N_7451);
nor U7595 (N_7595,N_7342,N_7306);
nand U7596 (N_7596,N_7372,N_7296);
nand U7597 (N_7597,N_7493,N_7362);
or U7598 (N_7598,N_7427,N_7434);
or U7599 (N_7599,N_7295,N_7265);
or U7600 (N_7600,N_7416,N_7456);
nand U7601 (N_7601,N_7348,N_7401);
and U7602 (N_7602,N_7332,N_7309);
xnor U7603 (N_7603,N_7440,N_7446);
or U7604 (N_7604,N_7255,N_7326);
and U7605 (N_7605,N_7378,N_7258);
or U7606 (N_7606,N_7329,N_7477);
xnor U7607 (N_7607,N_7331,N_7379);
or U7608 (N_7608,N_7369,N_7371);
xnor U7609 (N_7609,N_7406,N_7328);
or U7610 (N_7610,N_7472,N_7279);
and U7611 (N_7611,N_7438,N_7370);
nand U7612 (N_7612,N_7323,N_7368);
nand U7613 (N_7613,N_7293,N_7449);
nand U7614 (N_7614,N_7450,N_7457);
xnor U7615 (N_7615,N_7298,N_7398);
or U7616 (N_7616,N_7403,N_7444);
xor U7617 (N_7617,N_7486,N_7375);
xor U7618 (N_7618,N_7291,N_7283);
xnor U7619 (N_7619,N_7250,N_7325);
or U7620 (N_7620,N_7338,N_7386);
and U7621 (N_7621,N_7441,N_7445);
nor U7622 (N_7622,N_7448,N_7335);
nor U7623 (N_7623,N_7455,N_7479);
nand U7624 (N_7624,N_7415,N_7488);
xnor U7625 (N_7625,N_7425,N_7260);
xnor U7626 (N_7626,N_7444,N_7261);
or U7627 (N_7627,N_7470,N_7304);
nor U7628 (N_7628,N_7459,N_7387);
nand U7629 (N_7629,N_7296,N_7319);
or U7630 (N_7630,N_7363,N_7290);
nand U7631 (N_7631,N_7421,N_7457);
or U7632 (N_7632,N_7405,N_7470);
nor U7633 (N_7633,N_7408,N_7342);
and U7634 (N_7634,N_7389,N_7286);
nand U7635 (N_7635,N_7265,N_7358);
and U7636 (N_7636,N_7353,N_7278);
or U7637 (N_7637,N_7417,N_7404);
xnor U7638 (N_7638,N_7262,N_7323);
nor U7639 (N_7639,N_7257,N_7315);
and U7640 (N_7640,N_7283,N_7419);
and U7641 (N_7641,N_7288,N_7303);
nor U7642 (N_7642,N_7377,N_7408);
or U7643 (N_7643,N_7363,N_7431);
nor U7644 (N_7644,N_7431,N_7253);
and U7645 (N_7645,N_7449,N_7411);
nor U7646 (N_7646,N_7454,N_7394);
nand U7647 (N_7647,N_7297,N_7354);
nor U7648 (N_7648,N_7454,N_7498);
or U7649 (N_7649,N_7376,N_7364);
or U7650 (N_7650,N_7334,N_7463);
nor U7651 (N_7651,N_7257,N_7396);
or U7652 (N_7652,N_7444,N_7365);
xnor U7653 (N_7653,N_7397,N_7253);
and U7654 (N_7654,N_7282,N_7434);
nand U7655 (N_7655,N_7312,N_7494);
and U7656 (N_7656,N_7348,N_7453);
nor U7657 (N_7657,N_7465,N_7385);
and U7658 (N_7658,N_7344,N_7331);
nor U7659 (N_7659,N_7339,N_7440);
and U7660 (N_7660,N_7448,N_7411);
or U7661 (N_7661,N_7319,N_7393);
and U7662 (N_7662,N_7461,N_7375);
and U7663 (N_7663,N_7352,N_7303);
xor U7664 (N_7664,N_7456,N_7332);
or U7665 (N_7665,N_7392,N_7272);
nor U7666 (N_7666,N_7325,N_7258);
nor U7667 (N_7667,N_7424,N_7419);
nand U7668 (N_7668,N_7413,N_7443);
or U7669 (N_7669,N_7273,N_7418);
and U7670 (N_7670,N_7466,N_7260);
xor U7671 (N_7671,N_7413,N_7456);
nand U7672 (N_7672,N_7337,N_7325);
nand U7673 (N_7673,N_7291,N_7353);
nor U7674 (N_7674,N_7386,N_7420);
or U7675 (N_7675,N_7492,N_7416);
xnor U7676 (N_7676,N_7478,N_7287);
or U7677 (N_7677,N_7405,N_7427);
nor U7678 (N_7678,N_7339,N_7289);
nor U7679 (N_7679,N_7346,N_7470);
xnor U7680 (N_7680,N_7459,N_7380);
or U7681 (N_7681,N_7319,N_7452);
nor U7682 (N_7682,N_7336,N_7276);
xor U7683 (N_7683,N_7497,N_7462);
or U7684 (N_7684,N_7325,N_7388);
xor U7685 (N_7685,N_7499,N_7449);
and U7686 (N_7686,N_7462,N_7303);
nor U7687 (N_7687,N_7295,N_7401);
nand U7688 (N_7688,N_7354,N_7336);
nand U7689 (N_7689,N_7499,N_7493);
nor U7690 (N_7690,N_7393,N_7344);
or U7691 (N_7691,N_7471,N_7371);
xor U7692 (N_7692,N_7453,N_7390);
or U7693 (N_7693,N_7454,N_7449);
xnor U7694 (N_7694,N_7366,N_7475);
and U7695 (N_7695,N_7290,N_7413);
nand U7696 (N_7696,N_7478,N_7332);
nand U7697 (N_7697,N_7357,N_7408);
and U7698 (N_7698,N_7408,N_7469);
and U7699 (N_7699,N_7401,N_7449);
and U7700 (N_7700,N_7495,N_7457);
nand U7701 (N_7701,N_7326,N_7315);
xnor U7702 (N_7702,N_7321,N_7388);
nor U7703 (N_7703,N_7459,N_7468);
and U7704 (N_7704,N_7250,N_7319);
and U7705 (N_7705,N_7257,N_7251);
nor U7706 (N_7706,N_7432,N_7434);
or U7707 (N_7707,N_7490,N_7398);
and U7708 (N_7708,N_7395,N_7282);
and U7709 (N_7709,N_7434,N_7341);
xor U7710 (N_7710,N_7455,N_7443);
and U7711 (N_7711,N_7408,N_7392);
or U7712 (N_7712,N_7497,N_7307);
nand U7713 (N_7713,N_7284,N_7459);
nor U7714 (N_7714,N_7476,N_7272);
and U7715 (N_7715,N_7271,N_7325);
nand U7716 (N_7716,N_7367,N_7384);
or U7717 (N_7717,N_7314,N_7273);
or U7718 (N_7718,N_7396,N_7407);
nor U7719 (N_7719,N_7263,N_7484);
and U7720 (N_7720,N_7335,N_7332);
nand U7721 (N_7721,N_7348,N_7273);
nand U7722 (N_7722,N_7479,N_7284);
nand U7723 (N_7723,N_7292,N_7445);
nor U7724 (N_7724,N_7278,N_7341);
nand U7725 (N_7725,N_7440,N_7406);
nand U7726 (N_7726,N_7361,N_7313);
xor U7727 (N_7727,N_7389,N_7378);
xnor U7728 (N_7728,N_7326,N_7417);
or U7729 (N_7729,N_7376,N_7356);
and U7730 (N_7730,N_7448,N_7488);
xor U7731 (N_7731,N_7459,N_7480);
or U7732 (N_7732,N_7405,N_7396);
and U7733 (N_7733,N_7426,N_7416);
or U7734 (N_7734,N_7472,N_7287);
nand U7735 (N_7735,N_7286,N_7473);
xnor U7736 (N_7736,N_7319,N_7358);
nor U7737 (N_7737,N_7363,N_7329);
nor U7738 (N_7738,N_7323,N_7442);
nor U7739 (N_7739,N_7321,N_7473);
and U7740 (N_7740,N_7340,N_7380);
nand U7741 (N_7741,N_7465,N_7301);
nand U7742 (N_7742,N_7274,N_7452);
nor U7743 (N_7743,N_7327,N_7367);
or U7744 (N_7744,N_7272,N_7394);
nor U7745 (N_7745,N_7457,N_7402);
nor U7746 (N_7746,N_7309,N_7470);
nor U7747 (N_7747,N_7333,N_7335);
nand U7748 (N_7748,N_7494,N_7417);
and U7749 (N_7749,N_7476,N_7315);
nand U7750 (N_7750,N_7553,N_7645);
xnor U7751 (N_7751,N_7698,N_7706);
nor U7752 (N_7752,N_7686,N_7525);
or U7753 (N_7753,N_7615,N_7533);
or U7754 (N_7754,N_7624,N_7605);
xnor U7755 (N_7755,N_7544,N_7649);
or U7756 (N_7756,N_7683,N_7537);
nand U7757 (N_7757,N_7639,N_7586);
nor U7758 (N_7758,N_7551,N_7648);
nand U7759 (N_7759,N_7581,N_7567);
and U7760 (N_7760,N_7731,N_7628);
and U7761 (N_7761,N_7536,N_7743);
or U7762 (N_7762,N_7590,N_7550);
or U7763 (N_7763,N_7737,N_7647);
nor U7764 (N_7764,N_7502,N_7524);
nor U7765 (N_7765,N_7642,N_7509);
nor U7766 (N_7766,N_7671,N_7687);
xnor U7767 (N_7767,N_7704,N_7644);
xor U7768 (N_7768,N_7664,N_7727);
and U7769 (N_7769,N_7702,N_7679);
nor U7770 (N_7770,N_7629,N_7626);
xnor U7771 (N_7771,N_7701,N_7577);
xor U7772 (N_7772,N_7715,N_7508);
or U7773 (N_7773,N_7714,N_7747);
xnor U7774 (N_7774,N_7610,N_7543);
or U7775 (N_7775,N_7599,N_7657);
nor U7776 (N_7776,N_7717,N_7658);
xnor U7777 (N_7777,N_7589,N_7726);
or U7778 (N_7778,N_7580,N_7689);
or U7779 (N_7779,N_7622,N_7596);
nor U7780 (N_7780,N_7614,N_7584);
or U7781 (N_7781,N_7646,N_7637);
and U7782 (N_7782,N_7719,N_7660);
or U7783 (N_7783,N_7548,N_7670);
nor U7784 (N_7784,N_7549,N_7510);
xnor U7785 (N_7785,N_7598,N_7588);
or U7786 (N_7786,N_7542,N_7557);
xor U7787 (N_7787,N_7541,N_7675);
nand U7788 (N_7788,N_7620,N_7709);
nor U7789 (N_7789,N_7538,N_7652);
or U7790 (N_7790,N_7560,N_7554);
nor U7791 (N_7791,N_7676,N_7690);
xnor U7792 (N_7792,N_7523,N_7625);
nor U7793 (N_7793,N_7742,N_7749);
or U7794 (N_7794,N_7569,N_7619);
or U7795 (N_7795,N_7566,N_7655);
nor U7796 (N_7796,N_7656,N_7653);
or U7797 (N_7797,N_7516,N_7638);
or U7798 (N_7798,N_7568,N_7712);
nand U7799 (N_7799,N_7640,N_7735);
nor U7800 (N_7800,N_7733,N_7713);
and U7801 (N_7801,N_7722,N_7505);
xor U7802 (N_7802,N_7711,N_7562);
nand U7803 (N_7803,N_7650,N_7604);
nand U7804 (N_7804,N_7707,N_7504);
and U7805 (N_7805,N_7678,N_7730);
nor U7806 (N_7806,N_7745,N_7728);
nand U7807 (N_7807,N_7535,N_7613);
xnor U7808 (N_7808,N_7710,N_7695);
nor U7809 (N_7809,N_7587,N_7534);
and U7810 (N_7810,N_7659,N_7684);
and U7811 (N_7811,N_7597,N_7531);
xor U7812 (N_7812,N_7558,N_7691);
xor U7813 (N_7813,N_7705,N_7685);
nor U7814 (N_7814,N_7514,N_7739);
nor U7815 (N_7815,N_7555,N_7623);
xnor U7816 (N_7816,N_7521,N_7627);
or U7817 (N_7817,N_7547,N_7700);
xnor U7818 (N_7818,N_7602,N_7621);
or U7819 (N_7819,N_7725,N_7545);
nand U7820 (N_7820,N_7736,N_7616);
and U7821 (N_7821,N_7631,N_7672);
and U7822 (N_7822,N_7633,N_7559);
and U7823 (N_7823,N_7519,N_7643);
nand U7824 (N_7824,N_7608,N_7517);
xor U7825 (N_7825,N_7692,N_7716);
and U7826 (N_7826,N_7723,N_7738);
or U7827 (N_7827,N_7575,N_7574);
and U7828 (N_7828,N_7540,N_7618);
or U7829 (N_7829,N_7703,N_7666);
or U7830 (N_7830,N_7546,N_7669);
xnor U7831 (N_7831,N_7673,N_7539);
xor U7832 (N_7832,N_7732,N_7699);
xor U7833 (N_7833,N_7529,N_7518);
nand U7834 (N_7834,N_7708,N_7593);
and U7835 (N_7835,N_7688,N_7583);
and U7836 (N_7836,N_7552,N_7630);
nand U7837 (N_7837,N_7563,N_7667);
or U7838 (N_7838,N_7661,N_7665);
or U7839 (N_7839,N_7740,N_7724);
xor U7840 (N_7840,N_7578,N_7572);
xnor U7841 (N_7841,N_7532,N_7696);
xor U7842 (N_7842,N_7503,N_7641);
xnor U7843 (N_7843,N_7697,N_7609);
nor U7844 (N_7844,N_7677,N_7561);
or U7845 (N_7845,N_7526,N_7662);
xnor U7846 (N_7846,N_7564,N_7612);
or U7847 (N_7847,N_7741,N_7746);
nand U7848 (N_7848,N_7694,N_7668);
or U7849 (N_7849,N_7601,N_7682);
nand U7850 (N_7850,N_7527,N_7654);
nand U7851 (N_7851,N_7681,N_7636);
nor U7852 (N_7852,N_7528,N_7585);
and U7853 (N_7853,N_7634,N_7607);
or U7854 (N_7854,N_7595,N_7576);
nor U7855 (N_7855,N_7680,N_7571);
nand U7856 (N_7856,N_7606,N_7520);
xnor U7857 (N_7857,N_7500,N_7603);
nor U7858 (N_7858,N_7582,N_7635);
or U7859 (N_7859,N_7594,N_7718);
or U7860 (N_7860,N_7693,N_7512);
xor U7861 (N_7861,N_7611,N_7729);
nor U7862 (N_7862,N_7513,N_7632);
and U7863 (N_7863,N_7734,N_7674);
nand U7864 (N_7864,N_7507,N_7506);
and U7865 (N_7865,N_7515,N_7720);
nand U7866 (N_7866,N_7579,N_7744);
nor U7867 (N_7867,N_7522,N_7600);
nand U7868 (N_7868,N_7592,N_7573);
or U7869 (N_7869,N_7663,N_7530);
and U7870 (N_7870,N_7511,N_7591);
and U7871 (N_7871,N_7748,N_7565);
xnor U7872 (N_7872,N_7651,N_7721);
nor U7873 (N_7873,N_7501,N_7556);
xor U7874 (N_7874,N_7570,N_7617);
nor U7875 (N_7875,N_7503,N_7724);
and U7876 (N_7876,N_7683,N_7588);
and U7877 (N_7877,N_7527,N_7675);
and U7878 (N_7878,N_7732,N_7684);
nand U7879 (N_7879,N_7563,N_7529);
xor U7880 (N_7880,N_7693,N_7746);
or U7881 (N_7881,N_7584,N_7724);
nor U7882 (N_7882,N_7545,N_7575);
xnor U7883 (N_7883,N_7597,N_7711);
xor U7884 (N_7884,N_7600,N_7530);
or U7885 (N_7885,N_7657,N_7542);
xnor U7886 (N_7886,N_7522,N_7687);
nor U7887 (N_7887,N_7727,N_7638);
xor U7888 (N_7888,N_7608,N_7690);
or U7889 (N_7889,N_7536,N_7533);
or U7890 (N_7890,N_7551,N_7695);
or U7891 (N_7891,N_7548,N_7697);
xnor U7892 (N_7892,N_7678,N_7621);
or U7893 (N_7893,N_7594,N_7730);
nand U7894 (N_7894,N_7661,N_7531);
nand U7895 (N_7895,N_7530,N_7670);
and U7896 (N_7896,N_7735,N_7641);
xnor U7897 (N_7897,N_7735,N_7525);
or U7898 (N_7898,N_7594,N_7536);
or U7899 (N_7899,N_7704,N_7569);
nor U7900 (N_7900,N_7717,N_7534);
nand U7901 (N_7901,N_7737,N_7556);
nand U7902 (N_7902,N_7636,N_7550);
nor U7903 (N_7903,N_7645,N_7577);
and U7904 (N_7904,N_7668,N_7740);
or U7905 (N_7905,N_7663,N_7536);
nand U7906 (N_7906,N_7709,N_7651);
or U7907 (N_7907,N_7556,N_7635);
xor U7908 (N_7908,N_7737,N_7645);
and U7909 (N_7909,N_7737,N_7653);
xnor U7910 (N_7910,N_7607,N_7532);
or U7911 (N_7911,N_7543,N_7704);
or U7912 (N_7912,N_7516,N_7552);
nor U7913 (N_7913,N_7567,N_7697);
or U7914 (N_7914,N_7659,N_7733);
nor U7915 (N_7915,N_7654,N_7592);
and U7916 (N_7916,N_7663,N_7552);
and U7917 (N_7917,N_7545,N_7563);
or U7918 (N_7918,N_7630,N_7734);
xor U7919 (N_7919,N_7665,N_7646);
nand U7920 (N_7920,N_7615,N_7514);
and U7921 (N_7921,N_7502,N_7650);
and U7922 (N_7922,N_7555,N_7567);
xnor U7923 (N_7923,N_7682,N_7558);
xnor U7924 (N_7924,N_7597,N_7533);
nor U7925 (N_7925,N_7628,N_7646);
nor U7926 (N_7926,N_7600,N_7665);
nand U7927 (N_7927,N_7560,N_7545);
or U7928 (N_7928,N_7543,N_7540);
nor U7929 (N_7929,N_7664,N_7653);
and U7930 (N_7930,N_7686,N_7638);
and U7931 (N_7931,N_7605,N_7632);
xor U7932 (N_7932,N_7616,N_7604);
nand U7933 (N_7933,N_7536,N_7728);
xnor U7934 (N_7934,N_7733,N_7676);
nand U7935 (N_7935,N_7719,N_7517);
and U7936 (N_7936,N_7667,N_7518);
or U7937 (N_7937,N_7746,N_7733);
nand U7938 (N_7938,N_7618,N_7577);
xor U7939 (N_7939,N_7591,N_7536);
nand U7940 (N_7940,N_7742,N_7548);
xnor U7941 (N_7941,N_7658,N_7518);
or U7942 (N_7942,N_7537,N_7677);
nor U7943 (N_7943,N_7615,N_7732);
and U7944 (N_7944,N_7662,N_7628);
or U7945 (N_7945,N_7642,N_7582);
nand U7946 (N_7946,N_7525,N_7639);
xnor U7947 (N_7947,N_7513,N_7504);
nand U7948 (N_7948,N_7520,N_7705);
nor U7949 (N_7949,N_7665,N_7729);
nand U7950 (N_7950,N_7501,N_7618);
nor U7951 (N_7951,N_7598,N_7550);
and U7952 (N_7952,N_7625,N_7695);
xor U7953 (N_7953,N_7558,N_7553);
or U7954 (N_7954,N_7508,N_7512);
nor U7955 (N_7955,N_7693,N_7656);
nand U7956 (N_7956,N_7674,N_7675);
or U7957 (N_7957,N_7613,N_7701);
or U7958 (N_7958,N_7649,N_7581);
and U7959 (N_7959,N_7674,N_7611);
nand U7960 (N_7960,N_7516,N_7630);
xor U7961 (N_7961,N_7653,N_7574);
or U7962 (N_7962,N_7664,N_7564);
and U7963 (N_7963,N_7586,N_7708);
nor U7964 (N_7964,N_7679,N_7594);
and U7965 (N_7965,N_7577,N_7562);
or U7966 (N_7966,N_7714,N_7592);
nor U7967 (N_7967,N_7557,N_7555);
or U7968 (N_7968,N_7717,N_7610);
xor U7969 (N_7969,N_7606,N_7749);
nor U7970 (N_7970,N_7598,N_7587);
nor U7971 (N_7971,N_7591,N_7589);
nor U7972 (N_7972,N_7663,N_7632);
and U7973 (N_7973,N_7691,N_7552);
nand U7974 (N_7974,N_7558,N_7542);
or U7975 (N_7975,N_7566,N_7641);
nor U7976 (N_7976,N_7711,N_7746);
or U7977 (N_7977,N_7684,N_7693);
nor U7978 (N_7978,N_7533,N_7587);
nand U7979 (N_7979,N_7725,N_7645);
xnor U7980 (N_7980,N_7666,N_7699);
nand U7981 (N_7981,N_7715,N_7720);
xnor U7982 (N_7982,N_7739,N_7552);
nand U7983 (N_7983,N_7563,N_7591);
nor U7984 (N_7984,N_7637,N_7730);
nor U7985 (N_7985,N_7695,N_7706);
xnor U7986 (N_7986,N_7532,N_7617);
xnor U7987 (N_7987,N_7655,N_7633);
xnor U7988 (N_7988,N_7673,N_7613);
nor U7989 (N_7989,N_7557,N_7605);
xor U7990 (N_7990,N_7688,N_7578);
xnor U7991 (N_7991,N_7647,N_7518);
and U7992 (N_7992,N_7611,N_7588);
nor U7993 (N_7993,N_7526,N_7589);
xor U7994 (N_7994,N_7601,N_7652);
nand U7995 (N_7995,N_7641,N_7643);
xor U7996 (N_7996,N_7607,N_7676);
or U7997 (N_7997,N_7530,N_7593);
nor U7998 (N_7998,N_7663,N_7547);
nor U7999 (N_7999,N_7547,N_7715);
nand U8000 (N_8000,N_7798,N_7849);
nor U8001 (N_8001,N_7984,N_7949);
nor U8002 (N_8002,N_7942,N_7969);
xor U8003 (N_8003,N_7892,N_7906);
xor U8004 (N_8004,N_7924,N_7922);
or U8005 (N_8005,N_7888,N_7845);
nand U8006 (N_8006,N_7805,N_7960);
xor U8007 (N_8007,N_7935,N_7860);
or U8008 (N_8008,N_7936,N_7948);
xor U8009 (N_8009,N_7777,N_7870);
and U8010 (N_8010,N_7867,N_7901);
and U8011 (N_8011,N_7894,N_7873);
and U8012 (N_8012,N_7868,N_7891);
or U8013 (N_8013,N_7784,N_7752);
nor U8014 (N_8014,N_7972,N_7934);
nor U8015 (N_8015,N_7778,N_7751);
and U8016 (N_8016,N_7826,N_7963);
or U8017 (N_8017,N_7863,N_7895);
or U8018 (N_8018,N_7874,N_7928);
and U8019 (N_8019,N_7834,N_7846);
xnor U8020 (N_8020,N_7783,N_7915);
xnor U8021 (N_8021,N_7918,N_7768);
nor U8022 (N_8022,N_7802,N_7831);
xor U8023 (N_8023,N_7989,N_7961);
or U8024 (N_8024,N_7925,N_7799);
xnor U8025 (N_8025,N_7985,N_7885);
and U8026 (N_8026,N_7824,N_7780);
or U8027 (N_8027,N_7793,N_7847);
and U8028 (N_8028,N_7996,N_7764);
xnor U8029 (N_8029,N_7902,N_7825);
and U8030 (N_8030,N_7787,N_7986);
and U8031 (N_8031,N_7995,N_7794);
xor U8032 (N_8032,N_7788,N_7856);
and U8033 (N_8033,N_7758,N_7759);
xnor U8034 (N_8034,N_7843,N_7980);
and U8035 (N_8035,N_7931,N_7818);
nor U8036 (N_8036,N_7842,N_7887);
xnor U8037 (N_8037,N_7875,N_7998);
or U8038 (N_8038,N_7904,N_7757);
nand U8039 (N_8039,N_7871,N_7903);
nor U8040 (N_8040,N_7755,N_7907);
nor U8041 (N_8041,N_7872,N_7859);
or U8042 (N_8042,N_7968,N_7938);
or U8043 (N_8043,N_7916,N_7750);
nand U8044 (N_8044,N_7880,N_7862);
nand U8045 (N_8045,N_7990,N_7781);
nand U8046 (N_8046,N_7866,N_7886);
and U8047 (N_8047,N_7965,N_7993);
xnor U8048 (N_8048,N_7978,N_7970);
xor U8049 (N_8049,N_7876,N_7954);
xor U8050 (N_8050,N_7806,N_7837);
and U8051 (N_8051,N_7911,N_7910);
xnor U8052 (N_8052,N_7800,N_7797);
and U8053 (N_8053,N_7878,N_7857);
nor U8054 (N_8054,N_7850,N_7973);
nand U8055 (N_8055,N_7814,N_7956);
and U8056 (N_8056,N_7765,N_7991);
or U8057 (N_8057,N_7900,N_7763);
and U8058 (N_8058,N_7789,N_7905);
xor U8059 (N_8059,N_7877,N_7861);
nand U8060 (N_8060,N_7767,N_7829);
nand U8061 (N_8061,N_7955,N_7950);
nand U8062 (N_8062,N_7812,N_7770);
nand U8063 (N_8063,N_7813,N_7959);
and U8064 (N_8064,N_7908,N_7801);
xor U8065 (N_8065,N_7774,N_7939);
nor U8066 (N_8066,N_7761,N_7945);
or U8067 (N_8067,N_7881,N_7835);
nand U8068 (N_8068,N_7941,N_7756);
and U8069 (N_8069,N_7795,N_7773);
nand U8070 (N_8070,N_7827,N_7760);
nor U8071 (N_8071,N_7943,N_7952);
nor U8072 (N_8072,N_7772,N_7909);
nand U8073 (N_8073,N_7883,N_7988);
and U8074 (N_8074,N_7896,N_7809);
and U8075 (N_8075,N_7839,N_7766);
and U8076 (N_8076,N_7994,N_7917);
and U8077 (N_8077,N_7967,N_7944);
nor U8078 (N_8078,N_7869,N_7975);
nor U8079 (N_8079,N_7937,N_7786);
xnor U8080 (N_8080,N_7841,N_7853);
xnor U8081 (N_8081,N_7840,N_7971);
and U8082 (N_8082,N_7792,N_7890);
and U8083 (N_8083,N_7962,N_7811);
xnor U8084 (N_8084,N_7893,N_7782);
xnor U8085 (N_8085,N_7753,N_7929);
or U8086 (N_8086,N_7833,N_7912);
or U8087 (N_8087,N_7803,N_7854);
and U8088 (N_8088,N_7884,N_7977);
nand U8089 (N_8089,N_7852,N_7848);
and U8090 (N_8090,N_7923,N_7864);
and U8091 (N_8091,N_7983,N_7790);
xor U8092 (N_8092,N_7775,N_7920);
nand U8093 (N_8093,N_7879,N_7796);
and U8094 (N_8094,N_7940,N_7844);
and U8095 (N_8095,N_7776,N_7951);
nor U8096 (N_8096,N_7930,N_7855);
or U8097 (N_8097,N_7964,N_7919);
nor U8098 (N_8098,N_7815,N_7769);
nand U8099 (N_8099,N_7882,N_7851);
nor U8100 (N_8100,N_7821,N_7974);
nand U8101 (N_8101,N_7810,N_7865);
nand U8102 (N_8102,N_7817,N_7933);
xor U8103 (N_8103,N_7992,N_7823);
nor U8104 (N_8104,N_7804,N_7899);
xnor U8105 (N_8105,N_7999,N_7957);
nor U8106 (N_8106,N_7807,N_7966);
or U8107 (N_8107,N_7947,N_7932);
nand U8108 (N_8108,N_7897,N_7987);
nand U8109 (N_8109,N_7820,N_7946);
nor U8110 (N_8110,N_7979,N_7913);
or U8111 (N_8111,N_7976,N_7981);
nand U8112 (N_8112,N_7958,N_7982);
or U8113 (N_8113,N_7926,N_7858);
and U8114 (N_8114,N_7836,N_7779);
or U8115 (N_8115,N_7754,N_7808);
nand U8116 (N_8116,N_7898,N_7822);
nand U8117 (N_8117,N_7889,N_7921);
nor U8118 (N_8118,N_7791,N_7832);
or U8119 (N_8119,N_7819,N_7953);
nand U8120 (N_8120,N_7838,N_7816);
nor U8121 (N_8121,N_7785,N_7830);
nor U8122 (N_8122,N_7828,N_7762);
or U8123 (N_8123,N_7771,N_7927);
nor U8124 (N_8124,N_7914,N_7997);
or U8125 (N_8125,N_7835,N_7915);
and U8126 (N_8126,N_7875,N_7938);
xnor U8127 (N_8127,N_7842,N_7988);
xor U8128 (N_8128,N_7805,N_7916);
or U8129 (N_8129,N_7786,N_7950);
nand U8130 (N_8130,N_7888,N_7771);
xnor U8131 (N_8131,N_7964,N_7848);
and U8132 (N_8132,N_7765,N_7904);
or U8133 (N_8133,N_7930,N_7751);
xnor U8134 (N_8134,N_7933,N_7824);
nor U8135 (N_8135,N_7821,N_7943);
nor U8136 (N_8136,N_7985,N_7979);
nor U8137 (N_8137,N_7967,N_7848);
nand U8138 (N_8138,N_7860,N_7926);
nand U8139 (N_8139,N_7947,N_7780);
xor U8140 (N_8140,N_7816,N_7854);
xor U8141 (N_8141,N_7956,N_7761);
and U8142 (N_8142,N_7903,N_7999);
and U8143 (N_8143,N_7785,N_7833);
or U8144 (N_8144,N_7753,N_7756);
nor U8145 (N_8145,N_7768,N_7783);
nor U8146 (N_8146,N_7856,N_7892);
nand U8147 (N_8147,N_7830,N_7817);
nand U8148 (N_8148,N_7985,N_7836);
nor U8149 (N_8149,N_7886,N_7777);
nand U8150 (N_8150,N_7763,N_7863);
nand U8151 (N_8151,N_7997,N_7891);
and U8152 (N_8152,N_7927,N_7834);
xnor U8153 (N_8153,N_7776,N_7958);
xnor U8154 (N_8154,N_7805,N_7797);
xor U8155 (N_8155,N_7818,N_7830);
nand U8156 (N_8156,N_7883,N_7840);
or U8157 (N_8157,N_7982,N_7960);
nor U8158 (N_8158,N_7786,N_7951);
nand U8159 (N_8159,N_7814,N_7935);
and U8160 (N_8160,N_7971,N_7842);
xnor U8161 (N_8161,N_7876,N_7753);
nor U8162 (N_8162,N_7879,N_7857);
or U8163 (N_8163,N_7932,N_7829);
or U8164 (N_8164,N_7969,N_7932);
nand U8165 (N_8165,N_7769,N_7857);
and U8166 (N_8166,N_7755,N_7958);
xnor U8167 (N_8167,N_7800,N_7880);
nor U8168 (N_8168,N_7806,N_7864);
and U8169 (N_8169,N_7756,N_7946);
and U8170 (N_8170,N_7985,N_7969);
nand U8171 (N_8171,N_7769,N_7797);
xnor U8172 (N_8172,N_7860,N_7784);
nor U8173 (N_8173,N_7784,N_7805);
or U8174 (N_8174,N_7902,N_7914);
nor U8175 (N_8175,N_7774,N_7791);
or U8176 (N_8176,N_7750,N_7836);
xor U8177 (N_8177,N_7889,N_7975);
nand U8178 (N_8178,N_7844,N_7937);
and U8179 (N_8179,N_7961,N_7995);
nor U8180 (N_8180,N_7892,N_7963);
or U8181 (N_8181,N_7793,N_7922);
xor U8182 (N_8182,N_7947,N_7766);
nor U8183 (N_8183,N_7771,N_7837);
xor U8184 (N_8184,N_7902,N_7762);
or U8185 (N_8185,N_7940,N_7814);
and U8186 (N_8186,N_7915,N_7993);
xor U8187 (N_8187,N_7924,N_7849);
nand U8188 (N_8188,N_7950,N_7875);
and U8189 (N_8189,N_7968,N_7917);
xor U8190 (N_8190,N_7930,N_7868);
nor U8191 (N_8191,N_7872,N_7815);
nand U8192 (N_8192,N_7758,N_7936);
nand U8193 (N_8193,N_7865,N_7934);
or U8194 (N_8194,N_7961,N_7885);
nand U8195 (N_8195,N_7908,N_7944);
nand U8196 (N_8196,N_7791,N_7937);
and U8197 (N_8197,N_7883,N_7819);
nor U8198 (N_8198,N_7878,N_7803);
xnor U8199 (N_8199,N_7789,N_7922);
or U8200 (N_8200,N_7857,N_7793);
and U8201 (N_8201,N_7757,N_7835);
xor U8202 (N_8202,N_7752,N_7953);
xnor U8203 (N_8203,N_7960,N_7975);
nand U8204 (N_8204,N_7849,N_7774);
and U8205 (N_8205,N_7907,N_7794);
nand U8206 (N_8206,N_7791,N_7902);
or U8207 (N_8207,N_7877,N_7995);
and U8208 (N_8208,N_7936,N_7990);
nand U8209 (N_8209,N_7924,N_7862);
nor U8210 (N_8210,N_7908,N_7823);
xnor U8211 (N_8211,N_7837,N_7935);
xor U8212 (N_8212,N_7803,N_7965);
xor U8213 (N_8213,N_7994,N_7858);
nor U8214 (N_8214,N_7877,N_7989);
xnor U8215 (N_8215,N_7953,N_7924);
nor U8216 (N_8216,N_7894,N_7804);
nand U8217 (N_8217,N_7966,N_7967);
and U8218 (N_8218,N_7853,N_7769);
xnor U8219 (N_8219,N_7996,N_7787);
and U8220 (N_8220,N_7759,N_7847);
or U8221 (N_8221,N_7975,N_7796);
xor U8222 (N_8222,N_7923,N_7854);
or U8223 (N_8223,N_7858,N_7949);
nand U8224 (N_8224,N_7858,N_7937);
and U8225 (N_8225,N_7875,N_7972);
and U8226 (N_8226,N_7783,N_7995);
nor U8227 (N_8227,N_7840,N_7789);
and U8228 (N_8228,N_7756,N_7811);
nor U8229 (N_8229,N_7905,N_7919);
nand U8230 (N_8230,N_7850,N_7949);
or U8231 (N_8231,N_7984,N_7782);
xnor U8232 (N_8232,N_7974,N_7997);
or U8233 (N_8233,N_7924,N_7958);
or U8234 (N_8234,N_7821,N_7910);
nand U8235 (N_8235,N_7872,N_7869);
or U8236 (N_8236,N_7961,N_7752);
or U8237 (N_8237,N_7984,N_7834);
nand U8238 (N_8238,N_7929,N_7897);
nand U8239 (N_8239,N_7837,N_7939);
or U8240 (N_8240,N_7811,N_7999);
xnor U8241 (N_8241,N_7925,N_7997);
nand U8242 (N_8242,N_7753,N_7862);
or U8243 (N_8243,N_7969,N_7777);
xor U8244 (N_8244,N_7896,N_7866);
nor U8245 (N_8245,N_7883,N_7907);
xnor U8246 (N_8246,N_7872,N_7837);
nand U8247 (N_8247,N_7784,N_7918);
or U8248 (N_8248,N_7895,N_7955);
and U8249 (N_8249,N_7840,N_7791);
xnor U8250 (N_8250,N_8243,N_8063);
or U8251 (N_8251,N_8075,N_8224);
xnor U8252 (N_8252,N_8107,N_8039);
nand U8253 (N_8253,N_8122,N_8021);
and U8254 (N_8254,N_8031,N_8093);
xnor U8255 (N_8255,N_8111,N_8053);
nand U8256 (N_8256,N_8114,N_8097);
and U8257 (N_8257,N_8110,N_8038);
xor U8258 (N_8258,N_8001,N_8159);
xor U8259 (N_8259,N_8035,N_8043);
nor U8260 (N_8260,N_8189,N_8149);
nand U8261 (N_8261,N_8119,N_8181);
nor U8262 (N_8262,N_8142,N_8085);
and U8263 (N_8263,N_8147,N_8005);
and U8264 (N_8264,N_8092,N_8227);
xor U8265 (N_8265,N_8208,N_8015);
nand U8266 (N_8266,N_8161,N_8121);
and U8267 (N_8267,N_8176,N_8140);
and U8268 (N_8268,N_8061,N_8009);
xor U8269 (N_8269,N_8222,N_8100);
or U8270 (N_8270,N_8120,N_8150);
nor U8271 (N_8271,N_8192,N_8145);
or U8272 (N_8272,N_8198,N_8070);
or U8273 (N_8273,N_8249,N_8203);
or U8274 (N_8274,N_8175,N_8076);
nand U8275 (N_8275,N_8101,N_8073);
or U8276 (N_8276,N_8058,N_8086);
nor U8277 (N_8277,N_8012,N_8083);
nand U8278 (N_8278,N_8104,N_8199);
nor U8279 (N_8279,N_8131,N_8116);
xnor U8280 (N_8280,N_8064,N_8052);
nand U8281 (N_8281,N_8095,N_8055);
nor U8282 (N_8282,N_8229,N_8182);
nor U8283 (N_8283,N_8187,N_8210);
nand U8284 (N_8284,N_8117,N_8197);
xnor U8285 (N_8285,N_8193,N_8123);
or U8286 (N_8286,N_8235,N_8242);
or U8287 (N_8287,N_8071,N_8088);
and U8288 (N_8288,N_8136,N_8153);
nand U8289 (N_8289,N_8004,N_8002);
xnor U8290 (N_8290,N_8172,N_8056);
nand U8291 (N_8291,N_8084,N_8194);
xor U8292 (N_8292,N_8216,N_8118);
nor U8293 (N_8293,N_8127,N_8003);
xor U8294 (N_8294,N_8183,N_8163);
xor U8295 (N_8295,N_8047,N_8205);
xnor U8296 (N_8296,N_8139,N_8000);
nand U8297 (N_8297,N_8013,N_8178);
nor U8298 (N_8298,N_8184,N_8166);
nand U8299 (N_8299,N_8225,N_8233);
nor U8300 (N_8300,N_8022,N_8045);
and U8301 (N_8301,N_8232,N_8155);
nand U8302 (N_8302,N_8244,N_8200);
and U8303 (N_8303,N_8081,N_8141);
nand U8304 (N_8304,N_8019,N_8195);
and U8305 (N_8305,N_8134,N_8007);
nand U8306 (N_8306,N_8029,N_8125);
and U8307 (N_8307,N_8190,N_8068);
and U8308 (N_8308,N_8024,N_8011);
xnor U8309 (N_8309,N_8091,N_8236);
or U8310 (N_8310,N_8126,N_8204);
or U8311 (N_8311,N_8060,N_8078);
and U8312 (N_8312,N_8165,N_8206);
or U8313 (N_8313,N_8102,N_8173);
nand U8314 (N_8314,N_8219,N_8098);
and U8315 (N_8315,N_8037,N_8241);
and U8316 (N_8316,N_8143,N_8240);
xor U8317 (N_8317,N_8228,N_8167);
xnor U8318 (N_8318,N_8032,N_8246);
xnor U8319 (N_8319,N_8105,N_8212);
or U8320 (N_8320,N_8202,N_8023);
xnor U8321 (N_8321,N_8066,N_8169);
and U8322 (N_8322,N_8177,N_8248);
or U8323 (N_8323,N_8162,N_8221);
and U8324 (N_8324,N_8016,N_8089);
xor U8325 (N_8325,N_8094,N_8154);
nand U8326 (N_8326,N_8214,N_8026);
nand U8327 (N_8327,N_8239,N_8008);
and U8328 (N_8328,N_8062,N_8191);
nand U8329 (N_8329,N_8087,N_8157);
or U8330 (N_8330,N_8170,N_8112);
and U8331 (N_8331,N_8074,N_8196);
and U8332 (N_8332,N_8049,N_8158);
nor U8333 (N_8333,N_8027,N_8090);
and U8334 (N_8334,N_8168,N_8014);
or U8335 (N_8335,N_8077,N_8234);
and U8336 (N_8336,N_8059,N_8188);
or U8337 (N_8337,N_8124,N_8223);
nor U8338 (N_8338,N_8231,N_8115);
xor U8339 (N_8339,N_8207,N_8051);
nand U8340 (N_8340,N_8017,N_8042);
nand U8341 (N_8341,N_8171,N_8030);
xor U8342 (N_8342,N_8185,N_8186);
nand U8343 (N_8343,N_8137,N_8160);
nor U8344 (N_8344,N_8151,N_8006);
or U8345 (N_8345,N_8018,N_8072);
xor U8346 (N_8346,N_8148,N_8057);
nand U8347 (N_8347,N_8129,N_8033);
xnor U8348 (N_8348,N_8096,N_8130);
xor U8349 (N_8349,N_8099,N_8065);
xor U8350 (N_8350,N_8044,N_8152);
and U8351 (N_8351,N_8010,N_8025);
nor U8352 (N_8352,N_8226,N_8144);
or U8353 (N_8353,N_8237,N_8201);
nor U8354 (N_8354,N_8179,N_8174);
nand U8355 (N_8355,N_8213,N_8164);
and U8356 (N_8356,N_8238,N_8048);
nor U8357 (N_8357,N_8080,N_8069);
xor U8358 (N_8358,N_8133,N_8247);
nand U8359 (N_8359,N_8050,N_8215);
or U8360 (N_8360,N_8067,N_8046);
xnor U8361 (N_8361,N_8113,N_8041);
nand U8362 (N_8362,N_8103,N_8146);
nand U8363 (N_8363,N_8138,N_8020);
and U8364 (N_8364,N_8079,N_8220);
nor U8365 (N_8365,N_8109,N_8218);
and U8366 (N_8366,N_8211,N_8135);
nand U8367 (N_8367,N_8217,N_8036);
or U8368 (N_8368,N_8245,N_8034);
and U8369 (N_8369,N_8082,N_8156);
xor U8370 (N_8370,N_8209,N_8108);
xor U8371 (N_8371,N_8106,N_8040);
nor U8372 (N_8372,N_8180,N_8128);
xor U8373 (N_8373,N_8230,N_8132);
nand U8374 (N_8374,N_8028,N_8054);
and U8375 (N_8375,N_8118,N_8097);
nor U8376 (N_8376,N_8100,N_8115);
and U8377 (N_8377,N_8101,N_8068);
nor U8378 (N_8378,N_8117,N_8136);
and U8379 (N_8379,N_8231,N_8199);
xor U8380 (N_8380,N_8174,N_8123);
nor U8381 (N_8381,N_8006,N_8122);
xnor U8382 (N_8382,N_8001,N_8113);
nor U8383 (N_8383,N_8039,N_8196);
and U8384 (N_8384,N_8150,N_8189);
nor U8385 (N_8385,N_8027,N_8169);
and U8386 (N_8386,N_8142,N_8156);
nor U8387 (N_8387,N_8097,N_8210);
and U8388 (N_8388,N_8034,N_8171);
nand U8389 (N_8389,N_8161,N_8028);
nand U8390 (N_8390,N_8036,N_8243);
and U8391 (N_8391,N_8164,N_8246);
nor U8392 (N_8392,N_8228,N_8141);
nand U8393 (N_8393,N_8235,N_8145);
xor U8394 (N_8394,N_8156,N_8202);
nor U8395 (N_8395,N_8017,N_8039);
and U8396 (N_8396,N_8161,N_8020);
xnor U8397 (N_8397,N_8139,N_8180);
or U8398 (N_8398,N_8143,N_8003);
xor U8399 (N_8399,N_8097,N_8235);
or U8400 (N_8400,N_8225,N_8211);
and U8401 (N_8401,N_8220,N_8105);
or U8402 (N_8402,N_8114,N_8159);
nor U8403 (N_8403,N_8209,N_8117);
and U8404 (N_8404,N_8143,N_8069);
and U8405 (N_8405,N_8044,N_8227);
nand U8406 (N_8406,N_8192,N_8027);
nand U8407 (N_8407,N_8120,N_8211);
nor U8408 (N_8408,N_8167,N_8079);
and U8409 (N_8409,N_8030,N_8088);
or U8410 (N_8410,N_8109,N_8058);
or U8411 (N_8411,N_8187,N_8191);
or U8412 (N_8412,N_8202,N_8241);
xor U8413 (N_8413,N_8098,N_8228);
xnor U8414 (N_8414,N_8016,N_8237);
or U8415 (N_8415,N_8125,N_8048);
nor U8416 (N_8416,N_8181,N_8240);
or U8417 (N_8417,N_8023,N_8172);
and U8418 (N_8418,N_8120,N_8086);
nand U8419 (N_8419,N_8211,N_8029);
or U8420 (N_8420,N_8108,N_8237);
and U8421 (N_8421,N_8161,N_8199);
nand U8422 (N_8422,N_8159,N_8094);
nand U8423 (N_8423,N_8232,N_8194);
xnor U8424 (N_8424,N_8225,N_8216);
or U8425 (N_8425,N_8083,N_8212);
or U8426 (N_8426,N_8000,N_8065);
and U8427 (N_8427,N_8249,N_8134);
and U8428 (N_8428,N_8102,N_8133);
xnor U8429 (N_8429,N_8080,N_8235);
nand U8430 (N_8430,N_8065,N_8019);
xnor U8431 (N_8431,N_8182,N_8167);
or U8432 (N_8432,N_8016,N_8151);
nand U8433 (N_8433,N_8180,N_8047);
nand U8434 (N_8434,N_8185,N_8106);
nand U8435 (N_8435,N_8164,N_8241);
nor U8436 (N_8436,N_8037,N_8144);
or U8437 (N_8437,N_8246,N_8009);
and U8438 (N_8438,N_8011,N_8021);
and U8439 (N_8439,N_8089,N_8159);
or U8440 (N_8440,N_8204,N_8161);
and U8441 (N_8441,N_8150,N_8037);
xor U8442 (N_8442,N_8042,N_8019);
nand U8443 (N_8443,N_8097,N_8101);
nand U8444 (N_8444,N_8037,N_8162);
or U8445 (N_8445,N_8041,N_8197);
and U8446 (N_8446,N_8047,N_8050);
or U8447 (N_8447,N_8063,N_8037);
or U8448 (N_8448,N_8190,N_8242);
xnor U8449 (N_8449,N_8016,N_8188);
and U8450 (N_8450,N_8242,N_8076);
or U8451 (N_8451,N_8051,N_8141);
nand U8452 (N_8452,N_8128,N_8082);
xnor U8453 (N_8453,N_8118,N_8044);
nor U8454 (N_8454,N_8032,N_8147);
or U8455 (N_8455,N_8203,N_8047);
xnor U8456 (N_8456,N_8026,N_8042);
nand U8457 (N_8457,N_8148,N_8047);
and U8458 (N_8458,N_8100,N_8056);
xnor U8459 (N_8459,N_8092,N_8249);
nand U8460 (N_8460,N_8059,N_8245);
nand U8461 (N_8461,N_8156,N_8116);
xnor U8462 (N_8462,N_8018,N_8080);
nand U8463 (N_8463,N_8183,N_8014);
or U8464 (N_8464,N_8120,N_8210);
nand U8465 (N_8465,N_8248,N_8012);
xnor U8466 (N_8466,N_8069,N_8041);
xor U8467 (N_8467,N_8116,N_8237);
nand U8468 (N_8468,N_8002,N_8006);
nor U8469 (N_8469,N_8073,N_8132);
and U8470 (N_8470,N_8019,N_8060);
or U8471 (N_8471,N_8201,N_8077);
nand U8472 (N_8472,N_8211,N_8160);
nor U8473 (N_8473,N_8244,N_8000);
and U8474 (N_8474,N_8231,N_8061);
or U8475 (N_8475,N_8206,N_8168);
nand U8476 (N_8476,N_8071,N_8001);
nor U8477 (N_8477,N_8084,N_8057);
or U8478 (N_8478,N_8085,N_8157);
xnor U8479 (N_8479,N_8080,N_8077);
nor U8480 (N_8480,N_8085,N_8039);
nand U8481 (N_8481,N_8159,N_8210);
nand U8482 (N_8482,N_8167,N_8222);
xor U8483 (N_8483,N_8000,N_8062);
xor U8484 (N_8484,N_8231,N_8208);
xnor U8485 (N_8485,N_8123,N_8236);
xor U8486 (N_8486,N_8121,N_8027);
nand U8487 (N_8487,N_8010,N_8120);
or U8488 (N_8488,N_8074,N_8158);
or U8489 (N_8489,N_8170,N_8055);
or U8490 (N_8490,N_8160,N_8205);
nor U8491 (N_8491,N_8106,N_8021);
xor U8492 (N_8492,N_8010,N_8078);
nor U8493 (N_8493,N_8108,N_8227);
nor U8494 (N_8494,N_8191,N_8123);
xnor U8495 (N_8495,N_8089,N_8097);
or U8496 (N_8496,N_8181,N_8009);
nand U8497 (N_8497,N_8238,N_8006);
nor U8498 (N_8498,N_8182,N_8178);
and U8499 (N_8499,N_8242,N_8237);
xor U8500 (N_8500,N_8252,N_8339);
nor U8501 (N_8501,N_8463,N_8396);
nor U8502 (N_8502,N_8462,N_8406);
xor U8503 (N_8503,N_8495,N_8288);
nand U8504 (N_8504,N_8378,N_8416);
and U8505 (N_8505,N_8390,N_8344);
nor U8506 (N_8506,N_8284,N_8392);
nand U8507 (N_8507,N_8349,N_8274);
xor U8508 (N_8508,N_8366,N_8329);
nand U8509 (N_8509,N_8469,N_8404);
nor U8510 (N_8510,N_8418,N_8335);
and U8511 (N_8511,N_8261,N_8374);
nor U8512 (N_8512,N_8336,N_8389);
or U8513 (N_8513,N_8306,N_8379);
nor U8514 (N_8514,N_8403,N_8270);
or U8515 (N_8515,N_8386,N_8259);
and U8516 (N_8516,N_8408,N_8452);
or U8517 (N_8517,N_8393,N_8399);
and U8518 (N_8518,N_8364,N_8485);
and U8519 (N_8519,N_8251,N_8486);
nor U8520 (N_8520,N_8303,N_8254);
and U8521 (N_8521,N_8347,N_8474);
nand U8522 (N_8522,N_8465,N_8280);
or U8523 (N_8523,N_8441,N_8457);
and U8524 (N_8524,N_8295,N_8409);
or U8525 (N_8525,N_8415,N_8311);
nand U8526 (N_8526,N_8296,N_8494);
nor U8527 (N_8527,N_8262,N_8377);
nand U8528 (N_8528,N_8314,N_8285);
nand U8529 (N_8529,N_8273,N_8267);
nand U8530 (N_8530,N_8310,N_8454);
or U8531 (N_8531,N_8438,N_8313);
nand U8532 (N_8532,N_8286,N_8269);
nand U8533 (N_8533,N_8496,N_8498);
xnor U8534 (N_8534,N_8351,N_8304);
nand U8535 (N_8535,N_8343,N_8394);
nor U8536 (N_8536,N_8425,N_8384);
nor U8537 (N_8537,N_8302,N_8472);
or U8538 (N_8538,N_8411,N_8317);
or U8539 (N_8539,N_8354,N_8460);
xor U8540 (N_8540,N_8445,N_8299);
or U8541 (N_8541,N_8291,N_8467);
and U8542 (N_8542,N_8289,N_8375);
xor U8543 (N_8543,N_8401,N_8308);
nand U8544 (N_8544,N_8466,N_8279);
nand U8545 (N_8545,N_8435,N_8468);
xnor U8546 (N_8546,N_8423,N_8447);
nand U8547 (N_8547,N_8440,N_8437);
nor U8548 (N_8548,N_8405,N_8400);
and U8549 (N_8549,N_8464,N_8350);
nor U8550 (N_8550,N_8282,N_8353);
or U8551 (N_8551,N_8357,N_8397);
or U8552 (N_8552,N_8298,N_8410);
or U8553 (N_8553,N_8414,N_8258);
nand U8554 (N_8554,N_8356,N_8348);
nand U8555 (N_8555,N_8491,N_8337);
and U8556 (N_8556,N_8385,N_8319);
nand U8557 (N_8557,N_8361,N_8431);
nand U8558 (N_8558,N_8489,N_8265);
and U8559 (N_8559,N_8430,N_8432);
xor U8560 (N_8560,N_8439,N_8272);
nand U8561 (N_8561,N_8434,N_8278);
or U8562 (N_8562,N_8388,N_8448);
nor U8563 (N_8563,N_8358,N_8250);
nand U8564 (N_8564,N_8484,N_8476);
nand U8565 (N_8565,N_8422,N_8479);
xnor U8566 (N_8566,N_8455,N_8478);
nor U8567 (N_8567,N_8459,N_8473);
nor U8568 (N_8568,N_8324,N_8305);
and U8569 (N_8569,N_8382,N_8419);
xnor U8570 (N_8570,N_8487,N_8497);
xnor U8571 (N_8571,N_8475,N_8490);
xnor U8572 (N_8572,N_8321,N_8312);
xnor U8573 (N_8573,N_8307,N_8301);
and U8574 (N_8574,N_8499,N_8362);
nor U8575 (N_8575,N_8268,N_8446);
nor U8576 (N_8576,N_8407,N_8322);
nand U8577 (N_8577,N_8309,N_8290);
or U8578 (N_8578,N_8277,N_8331);
nor U8579 (N_8579,N_8297,N_8424);
nor U8580 (N_8580,N_8266,N_8417);
and U8581 (N_8581,N_8355,N_8481);
or U8582 (N_8582,N_8387,N_8294);
and U8583 (N_8583,N_8333,N_8367);
or U8584 (N_8584,N_8257,N_8426);
or U8585 (N_8585,N_8391,N_8334);
and U8586 (N_8586,N_8402,N_8345);
or U8587 (N_8587,N_8255,N_8341);
xor U8588 (N_8588,N_8275,N_8300);
nor U8589 (N_8589,N_8369,N_8352);
and U8590 (N_8590,N_8363,N_8480);
or U8591 (N_8591,N_8293,N_8380);
nor U8592 (N_8592,N_8492,N_8330);
or U8593 (N_8593,N_8338,N_8281);
or U8594 (N_8594,N_8287,N_8342);
xor U8595 (N_8595,N_8471,N_8458);
and U8596 (N_8596,N_8477,N_8263);
and U8597 (N_8597,N_8372,N_8420);
xor U8598 (N_8598,N_8453,N_8451);
xnor U8599 (N_8599,N_8271,N_8421);
nor U8600 (N_8600,N_8253,N_8443);
nand U8601 (N_8601,N_8264,N_8456);
and U8602 (N_8602,N_8332,N_8376);
and U8603 (N_8603,N_8427,N_8470);
nand U8604 (N_8604,N_8381,N_8260);
and U8605 (N_8605,N_8365,N_8368);
and U8606 (N_8606,N_8315,N_8316);
and U8607 (N_8607,N_8433,N_8383);
nand U8608 (N_8608,N_8283,N_8461);
xnor U8609 (N_8609,N_8256,N_8450);
xor U8610 (N_8610,N_8412,N_8327);
nand U8611 (N_8611,N_8398,N_8292);
xor U8612 (N_8612,N_8482,N_8442);
xor U8613 (N_8613,N_8370,N_8371);
nand U8614 (N_8614,N_8413,N_8493);
and U8615 (N_8615,N_8276,N_8488);
and U8616 (N_8616,N_8328,N_8318);
nand U8617 (N_8617,N_8320,N_8323);
xor U8618 (N_8618,N_8395,N_8340);
nor U8619 (N_8619,N_8326,N_8428);
nand U8620 (N_8620,N_8444,N_8360);
or U8621 (N_8621,N_8346,N_8429);
nor U8622 (N_8622,N_8449,N_8483);
xor U8623 (N_8623,N_8436,N_8373);
nand U8624 (N_8624,N_8325,N_8359);
nor U8625 (N_8625,N_8408,N_8458);
and U8626 (N_8626,N_8419,N_8320);
nor U8627 (N_8627,N_8259,N_8414);
xnor U8628 (N_8628,N_8390,N_8423);
xor U8629 (N_8629,N_8297,N_8435);
nand U8630 (N_8630,N_8337,N_8295);
xnor U8631 (N_8631,N_8462,N_8491);
nand U8632 (N_8632,N_8452,N_8395);
nand U8633 (N_8633,N_8456,N_8439);
xor U8634 (N_8634,N_8414,N_8444);
or U8635 (N_8635,N_8404,N_8483);
nor U8636 (N_8636,N_8285,N_8417);
xor U8637 (N_8637,N_8496,N_8455);
nor U8638 (N_8638,N_8291,N_8318);
or U8639 (N_8639,N_8432,N_8326);
nand U8640 (N_8640,N_8331,N_8450);
nor U8641 (N_8641,N_8315,N_8258);
nand U8642 (N_8642,N_8383,N_8480);
xor U8643 (N_8643,N_8490,N_8268);
nand U8644 (N_8644,N_8419,N_8388);
and U8645 (N_8645,N_8402,N_8411);
nor U8646 (N_8646,N_8326,N_8400);
nor U8647 (N_8647,N_8337,N_8308);
and U8648 (N_8648,N_8346,N_8333);
nand U8649 (N_8649,N_8338,N_8470);
nand U8650 (N_8650,N_8458,N_8487);
nor U8651 (N_8651,N_8454,N_8359);
nand U8652 (N_8652,N_8418,N_8406);
and U8653 (N_8653,N_8314,N_8294);
and U8654 (N_8654,N_8339,N_8333);
nor U8655 (N_8655,N_8396,N_8485);
or U8656 (N_8656,N_8258,N_8288);
and U8657 (N_8657,N_8263,N_8454);
or U8658 (N_8658,N_8440,N_8405);
or U8659 (N_8659,N_8273,N_8284);
and U8660 (N_8660,N_8395,N_8299);
nor U8661 (N_8661,N_8252,N_8441);
nor U8662 (N_8662,N_8409,N_8293);
and U8663 (N_8663,N_8431,N_8478);
nand U8664 (N_8664,N_8330,N_8475);
nor U8665 (N_8665,N_8342,N_8322);
and U8666 (N_8666,N_8371,N_8488);
nor U8667 (N_8667,N_8372,N_8264);
and U8668 (N_8668,N_8309,N_8397);
xor U8669 (N_8669,N_8481,N_8268);
or U8670 (N_8670,N_8371,N_8455);
nand U8671 (N_8671,N_8324,N_8393);
nor U8672 (N_8672,N_8481,N_8496);
nand U8673 (N_8673,N_8299,N_8358);
nor U8674 (N_8674,N_8269,N_8273);
xnor U8675 (N_8675,N_8390,N_8451);
nor U8676 (N_8676,N_8493,N_8386);
or U8677 (N_8677,N_8433,N_8400);
nand U8678 (N_8678,N_8309,N_8307);
nor U8679 (N_8679,N_8451,N_8291);
or U8680 (N_8680,N_8313,N_8341);
xnor U8681 (N_8681,N_8490,N_8297);
and U8682 (N_8682,N_8457,N_8254);
nor U8683 (N_8683,N_8469,N_8359);
or U8684 (N_8684,N_8311,N_8383);
and U8685 (N_8685,N_8488,N_8422);
nor U8686 (N_8686,N_8380,N_8456);
nor U8687 (N_8687,N_8327,N_8460);
nand U8688 (N_8688,N_8407,N_8431);
and U8689 (N_8689,N_8488,N_8445);
or U8690 (N_8690,N_8287,N_8457);
or U8691 (N_8691,N_8318,N_8379);
and U8692 (N_8692,N_8456,N_8262);
nor U8693 (N_8693,N_8276,N_8408);
nor U8694 (N_8694,N_8444,N_8474);
or U8695 (N_8695,N_8274,N_8454);
xor U8696 (N_8696,N_8474,N_8395);
nand U8697 (N_8697,N_8453,N_8424);
nand U8698 (N_8698,N_8399,N_8275);
and U8699 (N_8699,N_8285,N_8371);
xor U8700 (N_8700,N_8321,N_8494);
xor U8701 (N_8701,N_8325,N_8440);
and U8702 (N_8702,N_8263,N_8358);
nor U8703 (N_8703,N_8267,N_8447);
or U8704 (N_8704,N_8490,N_8414);
and U8705 (N_8705,N_8406,N_8482);
nand U8706 (N_8706,N_8367,N_8261);
xor U8707 (N_8707,N_8252,N_8282);
xor U8708 (N_8708,N_8312,N_8260);
nand U8709 (N_8709,N_8435,N_8448);
or U8710 (N_8710,N_8397,N_8422);
nand U8711 (N_8711,N_8471,N_8374);
or U8712 (N_8712,N_8286,N_8431);
xnor U8713 (N_8713,N_8281,N_8365);
xnor U8714 (N_8714,N_8433,N_8486);
nor U8715 (N_8715,N_8353,N_8438);
and U8716 (N_8716,N_8481,N_8472);
xor U8717 (N_8717,N_8449,N_8272);
nand U8718 (N_8718,N_8295,N_8497);
and U8719 (N_8719,N_8343,N_8458);
and U8720 (N_8720,N_8386,N_8291);
nor U8721 (N_8721,N_8349,N_8271);
nand U8722 (N_8722,N_8459,N_8475);
or U8723 (N_8723,N_8404,N_8482);
xor U8724 (N_8724,N_8284,N_8311);
nor U8725 (N_8725,N_8254,N_8393);
and U8726 (N_8726,N_8442,N_8409);
xnor U8727 (N_8727,N_8468,N_8349);
or U8728 (N_8728,N_8388,N_8420);
nand U8729 (N_8729,N_8362,N_8460);
nor U8730 (N_8730,N_8330,N_8416);
xor U8731 (N_8731,N_8355,N_8407);
or U8732 (N_8732,N_8461,N_8392);
nor U8733 (N_8733,N_8418,N_8369);
nor U8734 (N_8734,N_8417,N_8328);
nand U8735 (N_8735,N_8319,N_8263);
nand U8736 (N_8736,N_8330,N_8463);
nor U8737 (N_8737,N_8419,N_8426);
nand U8738 (N_8738,N_8405,N_8448);
or U8739 (N_8739,N_8270,N_8423);
nand U8740 (N_8740,N_8390,N_8488);
nor U8741 (N_8741,N_8327,N_8345);
or U8742 (N_8742,N_8296,N_8443);
and U8743 (N_8743,N_8290,N_8442);
or U8744 (N_8744,N_8327,N_8257);
or U8745 (N_8745,N_8377,N_8394);
xnor U8746 (N_8746,N_8416,N_8482);
and U8747 (N_8747,N_8402,N_8408);
xor U8748 (N_8748,N_8456,N_8447);
xnor U8749 (N_8749,N_8254,N_8490);
nor U8750 (N_8750,N_8633,N_8521);
nor U8751 (N_8751,N_8628,N_8707);
nand U8752 (N_8752,N_8640,N_8672);
xnor U8753 (N_8753,N_8613,N_8583);
xnor U8754 (N_8754,N_8559,N_8509);
and U8755 (N_8755,N_8673,N_8742);
nor U8756 (N_8756,N_8632,N_8724);
nand U8757 (N_8757,N_8556,N_8681);
nand U8758 (N_8758,N_8530,N_8537);
nand U8759 (N_8759,N_8591,N_8693);
and U8760 (N_8760,N_8720,N_8717);
and U8761 (N_8761,N_8695,N_8580);
nand U8762 (N_8762,N_8739,N_8533);
xnor U8763 (N_8763,N_8728,N_8502);
nor U8764 (N_8764,N_8526,N_8539);
nand U8765 (N_8765,N_8546,N_8549);
xnor U8766 (N_8766,N_8518,N_8595);
or U8767 (N_8767,N_8571,N_8726);
nor U8768 (N_8768,N_8642,N_8588);
or U8769 (N_8769,N_8531,N_8691);
nand U8770 (N_8770,N_8631,N_8500);
or U8771 (N_8771,N_8620,N_8596);
and U8772 (N_8772,N_8510,N_8586);
or U8773 (N_8773,N_8519,N_8678);
nor U8774 (N_8774,N_8582,N_8507);
nand U8775 (N_8775,N_8542,N_8748);
nor U8776 (N_8776,N_8505,N_8513);
xnor U8777 (N_8777,N_8705,N_8609);
xnor U8778 (N_8778,N_8696,N_8587);
nand U8779 (N_8779,N_8655,N_8653);
xnor U8780 (N_8780,N_8608,N_8698);
nor U8781 (N_8781,N_8687,N_8711);
or U8782 (N_8782,N_8567,N_8685);
nand U8783 (N_8783,N_8560,N_8700);
nand U8784 (N_8784,N_8575,N_8714);
nand U8785 (N_8785,N_8736,N_8611);
and U8786 (N_8786,N_8644,N_8654);
or U8787 (N_8787,N_8532,N_8503);
and U8788 (N_8788,N_8699,N_8585);
and U8789 (N_8789,N_8744,N_8598);
and U8790 (N_8790,N_8554,N_8543);
nor U8791 (N_8791,N_8683,N_8605);
or U8792 (N_8792,N_8501,N_8704);
nor U8793 (N_8793,N_8656,N_8740);
and U8794 (N_8794,N_8593,N_8718);
or U8795 (N_8795,N_8722,N_8675);
and U8796 (N_8796,N_8627,N_8721);
nor U8797 (N_8797,N_8630,N_8688);
nor U8798 (N_8798,N_8517,N_8636);
nor U8799 (N_8799,N_8729,N_8573);
and U8800 (N_8800,N_8527,N_8639);
nor U8801 (N_8801,N_8743,N_8663);
or U8802 (N_8802,N_8734,N_8525);
nor U8803 (N_8803,N_8650,N_8572);
or U8804 (N_8804,N_8679,N_8647);
or U8805 (N_8805,N_8523,N_8566);
nor U8806 (N_8806,N_8594,N_8702);
or U8807 (N_8807,N_8694,N_8658);
and U8808 (N_8808,N_8610,N_8619);
nand U8809 (N_8809,N_8689,N_8684);
xor U8810 (N_8810,N_8520,N_8738);
xnor U8811 (N_8811,N_8564,N_8599);
xor U8812 (N_8812,N_8731,N_8514);
xor U8813 (N_8813,N_8600,N_8657);
nand U8814 (N_8814,N_8651,N_8552);
and U8815 (N_8815,N_8727,N_8622);
nor U8816 (N_8816,N_8550,N_8579);
and U8817 (N_8817,N_8592,N_8607);
or U8818 (N_8818,N_8522,N_8601);
nand U8819 (N_8819,N_8645,N_8666);
xor U8820 (N_8820,N_8581,N_8618);
nor U8821 (N_8821,N_8561,N_8661);
nand U8822 (N_8822,N_8506,N_8528);
or U8823 (N_8823,N_8606,N_8735);
or U8824 (N_8824,N_8612,N_8545);
or U8825 (N_8825,N_8652,N_8646);
and U8826 (N_8826,N_8524,N_8569);
nor U8827 (N_8827,N_8625,N_8534);
and U8828 (N_8828,N_8697,N_8665);
or U8829 (N_8829,N_8590,N_8710);
xor U8830 (N_8830,N_8538,N_8741);
and U8831 (N_8831,N_8745,N_8547);
nand U8832 (N_8832,N_8648,N_8701);
or U8833 (N_8833,N_8617,N_8706);
nand U8834 (N_8834,N_8634,N_8643);
nand U8835 (N_8835,N_8548,N_8563);
and U8836 (N_8836,N_8703,N_8725);
or U8837 (N_8837,N_8529,N_8649);
nor U8838 (N_8838,N_8568,N_8659);
nand U8839 (N_8839,N_8623,N_8624);
and U8840 (N_8840,N_8574,N_8551);
nor U8841 (N_8841,N_8667,N_8716);
nand U8842 (N_8842,N_8709,N_8577);
xor U8843 (N_8843,N_8570,N_8616);
xor U8844 (N_8844,N_8638,N_8565);
and U8845 (N_8845,N_8746,N_8715);
or U8846 (N_8846,N_8737,N_8584);
and U8847 (N_8847,N_8749,N_8660);
xnor U8848 (N_8848,N_8671,N_8557);
nand U8849 (N_8849,N_8692,N_8668);
nand U8850 (N_8850,N_8578,N_8544);
and U8851 (N_8851,N_8597,N_8712);
and U8852 (N_8852,N_8615,N_8637);
and U8853 (N_8853,N_8515,N_8732);
nand U8854 (N_8854,N_8553,N_8662);
and U8855 (N_8855,N_8516,N_8669);
nand U8856 (N_8856,N_8677,N_8723);
nor U8857 (N_8857,N_8626,N_8733);
xnor U8858 (N_8858,N_8562,N_8558);
nand U8859 (N_8859,N_8641,N_8690);
nand U8860 (N_8860,N_8504,N_8664);
or U8861 (N_8861,N_8730,N_8719);
and U8862 (N_8862,N_8713,N_8708);
nor U8863 (N_8863,N_8614,N_8555);
xor U8864 (N_8864,N_8604,N_8535);
xor U8865 (N_8865,N_8682,N_8635);
or U8866 (N_8866,N_8629,N_8508);
nor U8867 (N_8867,N_8680,N_8747);
nor U8868 (N_8868,N_8621,N_8670);
nand U8869 (N_8869,N_8674,N_8676);
and U8870 (N_8870,N_8576,N_8603);
xnor U8871 (N_8871,N_8686,N_8589);
xnor U8872 (N_8872,N_8512,N_8602);
and U8873 (N_8873,N_8536,N_8511);
nand U8874 (N_8874,N_8541,N_8540);
or U8875 (N_8875,N_8563,N_8567);
xor U8876 (N_8876,N_8648,N_8589);
or U8877 (N_8877,N_8591,N_8689);
and U8878 (N_8878,N_8678,N_8571);
xor U8879 (N_8879,N_8693,N_8636);
and U8880 (N_8880,N_8591,N_8546);
xor U8881 (N_8881,N_8534,N_8546);
and U8882 (N_8882,N_8526,N_8730);
nor U8883 (N_8883,N_8630,N_8626);
nand U8884 (N_8884,N_8710,N_8629);
or U8885 (N_8885,N_8590,N_8550);
xnor U8886 (N_8886,N_8594,N_8642);
or U8887 (N_8887,N_8712,N_8643);
or U8888 (N_8888,N_8516,N_8596);
nor U8889 (N_8889,N_8653,N_8519);
or U8890 (N_8890,N_8545,N_8738);
and U8891 (N_8891,N_8506,N_8663);
or U8892 (N_8892,N_8546,N_8537);
nor U8893 (N_8893,N_8566,N_8549);
or U8894 (N_8894,N_8660,N_8626);
xnor U8895 (N_8895,N_8516,N_8575);
xor U8896 (N_8896,N_8606,N_8627);
or U8897 (N_8897,N_8691,N_8506);
or U8898 (N_8898,N_8718,N_8609);
xnor U8899 (N_8899,N_8534,N_8577);
or U8900 (N_8900,N_8631,N_8699);
nand U8901 (N_8901,N_8580,N_8712);
xor U8902 (N_8902,N_8617,N_8659);
nand U8903 (N_8903,N_8585,N_8515);
or U8904 (N_8904,N_8586,N_8709);
and U8905 (N_8905,N_8564,N_8678);
and U8906 (N_8906,N_8641,N_8650);
nor U8907 (N_8907,N_8590,N_8635);
or U8908 (N_8908,N_8648,N_8527);
nand U8909 (N_8909,N_8540,N_8700);
or U8910 (N_8910,N_8709,N_8693);
nor U8911 (N_8911,N_8588,N_8506);
xnor U8912 (N_8912,N_8679,N_8621);
nand U8913 (N_8913,N_8697,N_8714);
nor U8914 (N_8914,N_8540,N_8598);
or U8915 (N_8915,N_8628,N_8679);
nor U8916 (N_8916,N_8656,N_8708);
nor U8917 (N_8917,N_8590,N_8534);
nor U8918 (N_8918,N_8530,N_8618);
nand U8919 (N_8919,N_8599,N_8634);
or U8920 (N_8920,N_8573,N_8522);
nand U8921 (N_8921,N_8545,N_8670);
nand U8922 (N_8922,N_8557,N_8621);
nand U8923 (N_8923,N_8583,N_8716);
nor U8924 (N_8924,N_8533,N_8585);
nor U8925 (N_8925,N_8556,N_8651);
and U8926 (N_8926,N_8628,N_8503);
xnor U8927 (N_8927,N_8584,N_8605);
and U8928 (N_8928,N_8594,N_8625);
xnor U8929 (N_8929,N_8713,N_8552);
xnor U8930 (N_8930,N_8646,N_8726);
and U8931 (N_8931,N_8675,N_8569);
xnor U8932 (N_8932,N_8641,N_8623);
and U8933 (N_8933,N_8743,N_8520);
or U8934 (N_8934,N_8595,N_8544);
nand U8935 (N_8935,N_8613,N_8746);
and U8936 (N_8936,N_8549,N_8604);
or U8937 (N_8937,N_8749,N_8692);
nor U8938 (N_8938,N_8675,N_8696);
and U8939 (N_8939,N_8694,N_8552);
nor U8940 (N_8940,N_8578,N_8536);
and U8941 (N_8941,N_8667,N_8575);
and U8942 (N_8942,N_8563,N_8645);
and U8943 (N_8943,N_8698,N_8687);
or U8944 (N_8944,N_8702,N_8627);
or U8945 (N_8945,N_8727,N_8601);
nand U8946 (N_8946,N_8603,N_8614);
nand U8947 (N_8947,N_8749,N_8588);
or U8948 (N_8948,N_8727,N_8563);
nor U8949 (N_8949,N_8595,N_8527);
and U8950 (N_8950,N_8532,N_8596);
nand U8951 (N_8951,N_8692,N_8681);
xor U8952 (N_8952,N_8672,N_8620);
or U8953 (N_8953,N_8735,N_8622);
nand U8954 (N_8954,N_8680,N_8646);
and U8955 (N_8955,N_8717,N_8679);
and U8956 (N_8956,N_8600,N_8500);
or U8957 (N_8957,N_8705,N_8689);
or U8958 (N_8958,N_8560,N_8587);
or U8959 (N_8959,N_8525,N_8589);
or U8960 (N_8960,N_8582,N_8642);
nor U8961 (N_8961,N_8621,N_8702);
or U8962 (N_8962,N_8684,N_8548);
nand U8963 (N_8963,N_8604,N_8670);
or U8964 (N_8964,N_8554,N_8620);
or U8965 (N_8965,N_8596,N_8603);
and U8966 (N_8966,N_8622,N_8642);
or U8967 (N_8967,N_8601,N_8542);
xor U8968 (N_8968,N_8581,N_8723);
and U8969 (N_8969,N_8681,N_8685);
nand U8970 (N_8970,N_8555,N_8527);
xor U8971 (N_8971,N_8516,N_8580);
nor U8972 (N_8972,N_8509,N_8650);
or U8973 (N_8973,N_8588,N_8654);
nor U8974 (N_8974,N_8506,N_8744);
nand U8975 (N_8975,N_8587,N_8717);
nand U8976 (N_8976,N_8635,N_8693);
xor U8977 (N_8977,N_8681,N_8690);
nor U8978 (N_8978,N_8645,N_8745);
or U8979 (N_8979,N_8717,N_8594);
and U8980 (N_8980,N_8527,N_8659);
xnor U8981 (N_8981,N_8549,N_8631);
nand U8982 (N_8982,N_8553,N_8651);
or U8983 (N_8983,N_8585,N_8722);
nor U8984 (N_8984,N_8563,N_8547);
nor U8985 (N_8985,N_8634,N_8638);
nor U8986 (N_8986,N_8533,N_8551);
nand U8987 (N_8987,N_8738,N_8524);
nor U8988 (N_8988,N_8682,N_8620);
nand U8989 (N_8989,N_8639,N_8541);
nand U8990 (N_8990,N_8511,N_8560);
and U8991 (N_8991,N_8656,N_8528);
or U8992 (N_8992,N_8653,N_8533);
and U8993 (N_8993,N_8683,N_8663);
nand U8994 (N_8994,N_8516,N_8609);
xnor U8995 (N_8995,N_8526,N_8626);
xnor U8996 (N_8996,N_8740,N_8542);
or U8997 (N_8997,N_8641,N_8594);
or U8998 (N_8998,N_8677,N_8628);
and U8999 (N_8999,N_8720,N_8632);
and U9000 (N_9000,N_8865,N_8849);
and U9001 (N_9001,N_8836,N_8978);
or U9002 (N_9002,N_8795,N_8843);
nand U9003 (N_9003,N_8854,N_8835);
and U9004 (N_9004,N_8827,N_8871);
or U9005 (N_9005,N_8841,N_8907);
nor U9006 (N_9006,N_8816,N_8965);
nand U9007 (N_9007,N_8851,N_8863);
and U9008 (N_9008,N_8903,N_8959);
nand U9009 (N_9009,N_8869,N_8757);
and U9010 (N_9010,N_8796,N_8777);
nor U9011 (N_9011,N_8797,N_8824);
or U9012 (N_9012,N_8887,N_8801);
nor U9013 (N_9013,N_8883,N_8769);
nand U9014 (N_9014,N_8756,N_8894);
nor U9015 (N_9015,N_8780,N_8791);
nand U9016 (N_9016,N_8805,N_8804);
xor U9017 (N_9017,N_8826,N_8977);
and U9018 (N_9018,N_8954,N_8867);
and U9019 (N_9019,N_8917,N_8866);
nor U9020 (N_9020,N_8955,N_8789);
or U9021 (N_9021,N_8776,N_8808);
or U9022 (N_9022,N_8892,N_8957);
xor U9023 (N_9023,N_8817,N_8859);
nand U9024 (N_9024,N_8951,N_8833);
xor U9025 (N_9025,N_8874,N_8987);
nand U9026 (N_9026,N_8919,N_8885);
xor U9027 (N_9027,N_8834,N_8912);
or U9028 (N_9028,N_8927,N_8967);
nand U9029 (N_9029,N_8822,N_8914);
nor U9030 (N_9030,N_8971,N_8973);
and U9031 (N_9031,N_8992,N_8774);
nor U9032 (N_9032,N_8872,N_8985);
or U9033 (N_9033,N_8900,N_8782);
nor U9034 (N_9034,N_8750,N_8860);
or U9035 (N_9035,N_8794,N_8989);
and U9036 (N_9036,N_8921,N_8832);
and U9037 (N_9037,N_8825,N_8988);
and U9038 (N_9038,N_8788,N_8787);
and U9039 (N_9039,N_8831,N_8751);
or U9040 (N_9040,N_8844,N_8922);
or U9041 (N_9041,N_8845,N_8878);
or U9042 (N_9042,N_8966,N_8968);
nor U9043 (N_9043,N_8932,N_8870);
and U9044 (N_9044,N_8928,N_8896);
or U9045 (N_9045,N_8877,N_8908);
xnor U9046 (N_9046,N_8939,N_8862);
and U9047 (N_9047,N_8850,N_8775);
nor U9048 (N_9048,N_8924,N_8949);
nand U9049 (N_9049,N_8895,N_8781);
nand U9050 (N_9050,N_8884,N_8998);
xnor U9051 (N_9051,N_8893,N_8980);
or U9052 (N_9052,N_8864,N_8898);
and U9053 (N_9053,N_8943,N_8846);
nand U9054 (N_9054,N_8837,N_8948);
nand U9055 (N_9055,N_8760,N_8911);
or U9056 (N_9056,N_8848,N_8950);
and U9057 (N_9057,N_8940,N_8888);
nor U9058 (N_9058,N_8961,N_8991);
nor U9059 (N_9059,N_8983,N_8942);
nor U9060 (N_9060,N_8926,N_8875);
nand U9061 (N_9061,N_8937,N_8925);
or U9062 (N_9062,N_8916,N_8952);
and U9063 (N_9063,N_8963,N_8953);
nor U9064 (N_9064,N_8856,N_8993);
nor U9065 (N_9065,N_8990,N_8807);
and U9066 (N_9066,N_8838,N_8821);
and U9067 (N_9067,N_8785,N_8934);
xnor U9068 (N_9068,N_8800,N_8897);
nor U9069 (N_9069,N_8829,N_8913);
or U9070 (N_9070,N_8981,N_8938);
and U9071 (N_9071,N_8886,N_8759);
nand U9072 (N_9072,N_8812,N_8802);
xnor U9073 (N_9073,N_8999,N_8882);
nor U9074 (N_9074,N_8997,N_8899);
xnor U9075 (N_9075,N_8920,N_8762);
and U9076 (N_9076,N_8984,N_8935);
nand U9077 (N_9077,N_8770,N_8881);
or U9078 (N_9078,N_8861,N_8815);
nand U9079 (N_9079,N_8814,N_8960);
nor U9080 (N_9080,N_8929,N_8858);
and U9081 (N_9081,N_8873,N_8958);
nor U9082 (N_9082,N_8758,N_8974);
or U9083 (N_9083,N_8853,N_8975);
nor U9084 (N_9084,N_8778,N_8764);
nand U9085 (N_9085,N_8810,N_8910);
or U9086 (N_9086,N_8763,N_8779);
or U9087 (N_9087,N_8902,N_8793);
nor U9088 (N_9088,N_8772,N_8847);
or U9089 (N_9089,N_8755,N_8923);
xor U9090 (N_9090,N_8905,N_8972);
nand U9091 (N_9091,N_8809,N_8813);
nand U9092 (N_9092,N_8868,N_8996);
and U9093 (N_9093,N_8904,N_8964);
nand U9094 (N_9094,N_8799,N_8931);
xor U9095 (N_9095,N_8823,N_8930);
and U9096 (N_9096,N_8969,N_8818);
nand U9097 (N_9097,N_8995,N_8976);
and U9098 (N_9098,N_8947,N_8752);
or U9099 (N_9099,N_8891,N_8820);
or U9100 (N_9100,N_8962,N_8806);
or U9101 (N_9101,N_8784,N_8889);
or U9102 (N_9102,N_8819,N_8840);
and U9103 (N_9103,N_8790,N_8909);
xor U9104 (N_9104,N_8852,N_8944);
and U9105 (N_9105,N_8798,N_8766);
nand U9106 (N_9106,N_8876,N_8945);
xor U9107 (N_9107,N_8828,N_8970);
xnor U9108 (N_9108,N_8842,N_8906);
xnor U9109 (N_9109,N_8933,N_8918);
or U9110 (N_9110,N_8786,N_8761);
nor U9111 (N_9111,N_8890,N_8915);
nor U9112 (N_9112,N_8767,N_8941);
xnor U9113 (N_9113,N_8946,N_8754);
xor U9114 (N_9114,N_8986,N_8768);
and U9115 (N_9115,N_8879,N_8773);
nand U9116 (N_9116,N_8857,N_8936);
xor U9117 (N_9117,N_8811,N_8880);
nor U9118 (N_9118,N_8979,N_8792);
or U9119 (N_9119,N_8855,N_8765);
nand U9120 (N_9120,N_8982,N_8830);
nand U9121 (N_9121,N_8753,N_8803);
and U9122 (N_9122,N_8956,N_8839);
and U9123 (N_9123,N_8771,N_8994);
nor U9124 (N_9124,N_8901,N_8783);
nand U9125 (N_9125,N_8989,N_8973);
and U9126 (N_9126,N_8821,N_8964);
xnor U9127 (N_9127,N_8931,N_8891);
nand U9128 (N_9128,N_8899,N_8954);
nor U9129 (N_9129,N_8935,N_8897);
or U9130 (N_9130,N_8785,N_8957);
nand U9131 (N_9131,N_8936,N_8904);
nor U9132 (N_9132,N_8865,N_8834);
or U9133 (N_9133,N_8934,N_8888);
and U9134 (N_9134,N_8868,N_8940);
xor U9135 (N_9135,N_8811,N_8976);
xnor U9136 (N_9136,N_8858,N_8878);
nand U9137 (N_9137,N_8880,N_8898);
or U9138 (N_9138,N_8955,N_8821);
nand U9139 (N_9139,N_8999,N_8879);
nor U9140 (N_9140,N_8824,N_8933);
or U9141 (N_9141,N_8993,N_8858);
nor U9142 (N_9142,N_8818,N_8959);
and U9143 (N_9143,N_8918,N_8907);
or U9144 (N_9144,N_8818,N_8875);
and U9145 (N_9145,N_8751,N_8990);
nand U9146 (N_9146,N_8789,N_8995);
nor U9147 (N_9147,N_8780,N_8923);
nand U9148 (N_9148,N_8971,N_8772);
nor U9149 (N_9149,N_8757,N_8843);
and U9150 (N_9150,N_8797,N_8928);
and U9151 (N_9151,N_8887,N_8821);
and U9152 (N_9152,N_8991,N_8933);
xnor U9153 (N_9153,N_8970,N_8834);
and U9154 (N_9154,N_8792,N_8887);
nand U9155 (N_9155,N_8925,N_8896);
xor U9156 (N_9156,N_8965,N_8821);
nand U9157 (N_9157,N_8905,N_8894);
nor U9158 (N_9158,N_8980,N_8829);
and U9159 (N_9159,N_8773,N_8769);
nand U9160 (N_9160,N_8935,N_8902);
and U9161 (N_9161,N_8901,N_8992);
nor U9162 (N_9162,N_8822,N_8897);
xor U9163 (N_9163,N_8948,N_8945);
nor U9164 (N_9164,N_8908,N_8882);
or U9165 (N_9165,N_8955,N_8962);
and U9166 (N_9166,N_8802,N_8904);
and U9167 (N_9167,N_8919,N_8847);
xnor U9168 (N_9168,N_8804,N_8864);
and U9169 (N_9169,N_8841,N_8875);
nand U9170 (N_9170,N_8823,N_8820);
xnor U9171 (N_9171,N_8850,N_8854);
nand U9172 (N_9172,N_8965,N_8753);
or U9173 (N_9173,N_8848,N_8818);
or U9174 (N_9174,N_8849,N_8783);
nor U9175 (N_9175,N_8775,N_8833);
nor U9176 (N_9176,N_8999,N_8889);
xor U9177 (N_9177,N_8842,N_8792);
or U9178 (N_9178,N_8984,N_8965);
and U9179 (N_9179,N_8833,N_8937);
nand U9180 (N_9180,N_8771,N_8819);
or U9181 (N_9181,N_8795,N_8785);
or U9182 (N_9182,N_8934,N_8988);
xnor U9183 (N_9183,N_8902,N_8946);
nand U9184 (N_9184,N_8760,N_8984);
xor U9185 (N_9185,N_8750,N_8765);
and U9186 (N_9186,N_8946,N_8960);
and U9187 (N_9187,N_8881,N_8774);
or U9188 (N_9188,N_8930,N_8955);
and U9189 (N_9189,N_8769,N_8757);
or U9190 (N_9190,N_8923,N_8778);
or U9191 (N_9191,N_8825,N_8828);
and U9192 (N_9192,N_8827,N_8900);
or U9193 (N_9193,N_8891,N_8796);
nand U9194 (N_9194,N_8936,N_8983);
and U9195 (N_9195,N_8987,N_8897);
nor U9196 (N_9196,N_8793,N_8893);
or U9197 (N_9197,N_8819,N_8905);
nand U9198 (N_9198,N_8852,N_8754);
nor U9199 (N_9199,N_8943,N_8802);
and U9200 (N_9200,N_8932,N_8818);
and U9201 (N_9201,N_8760,N_8953);
nor U9202 (N_9202,N_8913,N_8948);
and U9203 (N_9203,N_8877,N_8886);
or U9204 (N_9204,N_8793,N_8826);
nand U9205 (N_9205,N_8771,N_8925);
xnor U9206 (N_9206,N_8986,N_8851);
nor U9207 (N_9207,N_8927,N_8854);
nand U9208 (N_9208,N_8980,N_8813);
xnor U9209 (N_9209,N_8821,N_8803);
nand U9210 (N_9210,N_8954,N_8756);
and U9211 (N_9211,N_8911,N_8789);
or U9212 (N_9212,N_8753,N_8816);
nor U9213 (N_9213,N_8983,N_8766);
and U9214 (N_9214,N_8827,N_8860);
xor U9215 (N_9215,N_8917,N_8812);
nand U9216 (N_9216,N_8786,N_8983);
xnor U9217 (N_9217,N_8950,N_8901);
xor U9218 (N_9218,N_8778,N_8900);
or U9219 (N_9219,N_8870,N_8785);
nand U9220 (N_9220,N_8821,N_8890);
nand U9221 (N_9221,N_8801,N_8824);
or U9222 (N_9222,N_8830,N_8968);
nand U9223 (N_9223,N_8822,N_8943);
xor U9224 (N_9224,N_8899,N_8968);
xnor U9225 (N_9225,N_8940,N_8810);
or U9226 (N_9226,N_8797,N_8926);
or U9227 (N_9227,N_8896,N_8904);
nor U9228 (N_9228,N_8959,N_8784);
nor U9229 (N_9229,N_8967,N_8785);
nor U9230 (N_9230,N_8759,N_8884);
nor U9231 (N_9231,N_8773,N_8761);
or U9232 (N_9232,N_8785,N_8826);
xor U9233 (N_9233,N_8872,N_8765);
nand U9234 (N_9234,N_8869,N_8805);
nand U9235 (N_9235,N_8847,N_8907);
or U9236 (N_9236,N_8927,N_8928);
and U9237 (N_9237,N_8996,N_8805);
and U9238 (N_9238,N_8842,N_8938);
nand U9239 (N_9239,N_8931,N_8766);
xnor U9240 (N_9240,N_8938,N_8839);
nand U9241 (N_9241,N_8985,N_8995);
or U9242 (N_9242,N_8914,N_8885);
or U9243 (N_9243,N_8928,N_8826);
nor U9244 (N_9244,N_8765,N_8821);
and U9245 (N_9245,N_8916,N_8812);
xnor U9246 (N_9246,N_8968,N_8832);
nand U9247 (N_9247,N_8861,N_8980);
or U9248 (N_9248,N_8984,N_8798);
nor U9249 (N_9249,N_8930,N_8977);
and U9250 (N_9250,N_9032,N_9147);
and U9251 (N_9251,N_9082,N_9109);
nor U9252 (N_9252,N_9214,N_9155);
or U9253 (N_9253,N_9093,N_9189);
and U9254 (N_9254,N_9160,N_9039);
or U9255 (N_9255,N_9102,N_9111);
nor U9256 (N_9256,N_9050,N_9004);
or U9257 (N_9257,N_9203,N_9121);
nor U9258 (N_9258,N_9126,N_9108);
or U9259 (N_9259,N_9092,N_9249);
nor U9260 (N_9260,N_9038,N_9088);
and U9261 (N_9261,N_9045,N_9059);
nand U9262 (N_9262,N_9187,N_9163);
and U9263 (N_9263,N_9218,N_9112);
or U9264 (N_9264,N_9028,N_9210);
nand U9265 (N_9265,N_9058,N_9242);
nor U9266 (N_9266,N_9070,N_9106);
or U9267 (N_9267,N_9083,N_9068);
xor U9268 (N_9268,N_9179,N_9029);
nor U9269 (N_9269,N_9167,N_9177);
nor U9270 (N_9270,N_9193,N_9033);
xnor U9271 (N_9271,N_9144,N_9199);
or U9272 (N_9272,N_9094,N_9002);
or U9273 (N_9273,N_9086,N_9031);
and U9274 (N_9274,N_9145,N_9003);
nand U9275 (N_9275,N_9128,N_9209);
or U9276 (N_9276,N_9204,N_9046);
nand U9277 (N_9277,N_9194,N_9156);
xor U9278 (N_9278,N_9183,N_9150);
xnor U9279 (N_9279,N_9116,N_9162);
xor U9280 (N_9280,N_9175,N_9178);
and U9281 (N_9281,N_9247,N_9005);
nand U9282 (N_9282,N_9018,N_9165);
or U9283 (N_9283,N_9008,N_9117);
nor U9284 (N_9284,N_9076,N_9011);
xor U9285 (N_9285,N_9164,N_9014);
and U9286 (N_9286,N_9080,N_9065);
xnor U9287 (N_9287,N_9051,N_9021);
nor U9288 (N_9288,N_9030,N_9152);
or U9289 (N_9289,N_9235,N_9101);
xor U9290 (N_9290,N_9107,N_9173);
nor U9291 (N_9291,N_9007,N_9232);
nor U9292 (N_9292,N_9159,N_9140);
nand U9293 (N_9293,N_9228,N_9224);
and U9294 (N_9294,N_9157,N_9123);
nand U9295 (N_9295,N_9133,N_9026);
nor U9296 (N_9296,N_9205,N_9115);
xnor U9297 (N_9297,N_9091,N_9085);
or U9298 (N_9298,N_9171,N_9132);
nor U9299 (N_9299,N_9020,N_9191);
and U9300 (N_9300,N_9110,N_9089);
xnor U9301 (N_9301,N_9061,N_9148);
xnor U9302 (N_9302,N_9053,N_9015);
nand U9303 (N_9303,N_9119,N_9146);
nand U9304 (N_9304,N_9222,N_9137);
nor U9305 (N_9305,N_9190,N_9024);
and U9306 (N_9306,N_9064,N_9069);
and U9307 (N_9307,N_9138,N_9196);
and U9308 (N_9308,N_9198,N_9067);
or U9309 (N_9309,N_9236,N_9166);
and U9310 (N_9310,N_9221,N_9048);
nor U9311 (N_9311,N_9043,N_9248);
nor U9312 (N_9312,N_9034,N_9142);
or U9313 (N_9313,N_9216,N_9184);
or U9314 (N_9314,N_9040,N_9013);
nand U9315 (N_9315,N_9154,N_9139);
nor U9316 (N_9316,N_9239,N_9097);
or U9317 (N_9317,N_9079,N_9237);
or U9318 (N_9318,N_9245,N_9225);
nor U9319 (N_9319,N_9240,N_9114);
nand U9320 (N_9320,N_9136,N_9169);
xor U9321 (N_9321,N_9072,N_9118);
or U9322 (N_9322,N_9201,N_9151);
and U9323 (N_9323,N_9104,N_9042);
and U9324 (N_9324,N_9087,N_9100);
and U9325 (N_9325,N_9230,N_9044);
nand U9326 (N_9326,N_9016,N_9153);
nor U9327 (N_9327,N_9006,N_9027);
nor U9328 (N_9328,N_9023,N_9186);
xnor U9329 (N_9329,N_9066,N_9010);
nor U9330 (N_9330,N_9056,N_9226);
xnor U9331 (N_9331,N_9176,N_9081);
nor U9332 (N_9332,N_9130,N_9057);
xnor U9333 (N_9333,N_9241,N_9244);
nand U9334 (N_9334,N_9170,N_9096);
and U9335 (N_9335,N_9212,N_9054);
nor U9336 (N_9336,N_9062,N_9217);
nor U9337 (N_9337,N_9223,N_9161);
nand U9338 (N_9338,N_9095,N_9197);
and U9339 (N_9339,N_9049,N_9143);
xnor U9340 (N_9340,N_9055,N_9246);
nand U9341 (N_9341,N_9125,N_9229);
or U9342 (N_9342,N_9090,N_9036);
nor U9343 (N_9343,N_9022,N_9060);
nor U9344 (N_9344,N_9000,N_9172);
or U9345 (N_9345,N_9025,N_9105);
xor U9346 (N_9346,N_9149,N_9238);
or U9347 (N_9347,N_9129,N_9134);
or U9348 (N_9348,N_9180,N_9052);
xnor U9349 (N_9349,N_9185,N_9202);
nor U9350 (N_9350,N_9207,N_9124);
xnor U9351 (N_9351,N_9113,N_9041);
and U9352 (N_9352,N_9019,N_9084);
nand U9353 (N_9353,N_9127,N_9174);
xnor U9354 (N_9354,N_9141,N_9231);
nand U9355 (N_9355,N_9099,N_9200);
or U9356 (N_9356,N_9234,N_9035);
or U9357 (N_9357,N_9168,N_9211);
and U9358 (N_9358,N_9075,N_9195);
nor U9359 (N_9359,N_9233,N_9181);
nor U9360 (N_9360,N_9243,N_9227);
and U9361 (N_9361,N_9037,N_9074);
or U9362 (N_9362,N_9047,N_9213);
xnor U9363 (N_9363,N_9017,N_9098);
or U9364 (N_9364,N_9103,N_9071);
nor U9365 (N_9365,N_9009,N_9001);
nor U9366 (N_9366,N_9182,N_9077);
and U9367 (N_9367,N_9078,N_9220);
and U9368 (N_9368,N_9208,N_9219);
and U9369 (N_9369,N_9192,N_9215);
or U9370 (N_9370,N_9012,N_9158);
or U9371 (N_9371,N_9073,N_9122);
or U9372 (N_9372,N_9120,N_9206);
nor U9373 (N_9373,N_9063,N_9135);
and U9374 (N_9374,N_9188,N_9131);
xnor U9375 (N_9375,N_9213,N_9025);
or U9376 (N_9376,N_9074,N_9023);
or U9377 (N_9377,N_9240,N_9179);
or U9378 (N_9378,N_9125,N_9104);
and U9379 (N_9379,N_9101,N_9098);
nand U9380 (N_9380,N_9222,N_9000);
nor U9381 (N_9381,N_9027,N_9073);
or U9382 (N_9382,N_9214,N_9158);
and U9383 (N_9383,N_9073,N_9215);
nand U9384 (N_9384,N_9205,N_9207);
or U9385 (N_9385,N_9193,N_9075);
and U9386 (N_9386,N_9237,N_9220);
xnor U9387 (N_9387,N_9206,N_9033);
xor U9388 (N_9388,N_9181,N_9175);
or U9389 (N_9389,N_9026,N_9221);
nand U9390 (N_9390,N_9213,N_9040);
xnor U9391 (N_9391,N_9195,N_9072);
nand U9392 (N_9392,N_9247,N_9086);
xor U9393 (N_9393,N_9079,N_9033);
nor U9394 (N_9394,N_9086,N_9063);
and U9395 (N_9395,N_9174,N_9100);
and U9396 (N_9396,N_9171,N_9142);
and U9397 (N_9397,N_9011,N_9013);
xor U9398 (N_9398,N_9165,N_9200);
nor U9399 (N_9399,N_9064,N_9040);
or U9400 (N_9400,N_9207,N_9111);
and U9401 (N_9401,N_9193,N_9115);
nor U9402 (N_9402,N_9190,N_9032);
nor U9403 (N_9403,N_9114,N_9111);
xor U9404 (N_9404,N_9247,N_9025);
xor U9405 (N_9405,N_9218,N_9092);
and U9406 (N_9406,N_9106,N_9214);
xnor U9407 (N_9407,N_9015,N_9234);
and U9408 (N_9408,N_9055,N_9119);
xor U9409 (N_9409,N_9002,N_9224);
nand U9410 (N_9410,N_9153,N_9013);
or U9411 (N_9411,N_9134,N_9116);
and U9412 (N_9412,N_9202,N_9097);
nor U9413 (N_9413,N_9172,N_9012);
nand U9414 (N_9414,N_9010,N_9128);
xnor U9415 (N_9415,N_9183,N_9056);
and U9416 (N_9416,N_9218,N_9131);
or U9417 (N_9417,N_9049,N_9216);
or U9418 (N_9418,N_9064,N_9071);
xor U9419 (N_9419,N_9040,N_9043);
nand U9420 (N_9420,N_9105,N_9014);
and U9421 (N_9421,N_9110,N_9150);
and U9422 (N_9422,N_9174,N_9177);
nor U9423 (N_9423,N_9132,N_9081);
nand U9424 (N_9424,N_9132,N_9064);
and U9425 (N_9425,N_9109,N_9021);
nand U9426 (N_9426,N_9195,N_9071);
and U9427 (N_9427,N_9177,N_9206);
nor U9428 (N_9428,N_9069,N_9110);
nand U9429 (N_9429,N_9105,N_9242);
or U9430 (N_9430,N_9111,N_9201);
xor U9431 (N_9431,N_9029,N_9070);
or U9432 (N_9432,N_9013,N_9065);
nor U9433 (N_9433,N_9084,N_9057);
nand U9434 (N_9434,N_9006,N_9124);
nand U9435 (N_9435,N_9013,N_9223);
and U9436 (N_9436,N_9157,N_9041);
xor U9437 (N_9437,N_9164,N_9020);
xor U9438 (N_9438,N_9008,N_9026);
nor U9439 (N_9439,N_9100,N_9054);
or U9440 (N_9440,N_9116,N_9169);
and U9441 (N_9441,N_9127,N_9090);
nand U9442 (N_9442,N_9049,N_9228);
and U9443 (N_9443,N_9006,N_9162);
xnor U9444 (N_9444,N_9245,N_9234);
nor U9445 (N_9445,N_9247,N_9214);
nor U9446 (N_9446,N_9225,N_9147);
or U9447 (N_9447,N_9098,N_9173);
nand U9448 (N_9448,N_9228,N_9182);
nor U9449 (N_9449,N_9126,N_9053);
xnor U9450 (N_9450,N_9085,N_9231);
nor U9451 (N_9451,N_9175,N_9018);
xor U9452 (N_9452,N_9149,N_9136);
and U9453 (N_9453,N_9090,N_9073);
or U9454 (N_9454,N_9216,N_9074);
nand U9455 (N_9455,N_9040,N_9192);
nand U9456 (N_9456,N_9213,N_9245);
nor U9457 (N_9457,N_9040,N_9038);
nor U9458 (N_9458,N_9177,N_9122);
or U9459 (N_9459,N_9012,N_9243);
nand U9460 (N_9460,N_9057,N_9220);
nor U9461 (N_9461,N_9123,N_9125);
and U9462 (N_9462,N_9247,N_9227);
and U9463 (N_9463,N_9011,N_9052);
and U9464 (N_9464,N_9112,N_9155);
and U9465 (N_9465,N_9133,N_9166);
nand U9466 (N_9466,N_9013,N_9017);
and U9467 (N_9467,N_9130,N_9072);
nor U9468 (N_9468,N_9001,N_9021);
xnor U9469 (N_9469,N_9141,N_9217);
nor U9470 (N_9470,N_9032,N_9013);
nand U9471 (N_9471,N_9040,N_9093);
and U9472 (N_9472,N_9033,N_9142);
nand U9473 (N_9473,N_9183,N_9218);
nand U9474 (N_9474,N_9014,N_9247);
or U9475 (N_9475,N_9121,N_9221);
or U9476 (N_9476,N_9090,N_9060);
nand U9477 (N_9477,N_9107,N_9222);
or U9478 (N_9478,N_9185,N_9115);
or U9479 (N_9479,N_9129,N_9031);
and U9480 (N_9480,N_9022,N_9073);
nor U9481 (N_9481,N_9103,N_9213);
nor U9482 (N_9482,N_9119,N_9157);
nor U9483 (N_9483,N_9070,N_9213);
nand U9484 (N_9484,N_9114,N_9172);
or U9485 (N_9485,N_9132,N_9098);
or U9486 (N_9486,N_9228,N_9024);
nand U9487 (N_9487,N_9089,N_9223);
nand U9488 (N_9488,N_9120,N_9138);
nand U9489 (N_9489,N_9216,N_9039);
or U9490 (N_9490,N_9151,N_9205);
nor U9491 (N_9491,N_9205,N_9210);
nand U9492 (N_9492,N_9001,N_9121);
nor U9493 (N_9493,N_9237,N_9106);
nand U9494 (N_9494,N_9088,N_9065);
nor U9495 (N_9495,N_9193,N_9129);
nand U9496 (N_9496,N_9139,N_9009);
xor U9497 (N_9497,N_9147,N_9077);
or U9498 (N_9498,N_9061,N_9186);
xor U9499 (N_9499,N_9142,N_9219);
xnor U9500 (N_9500,N_9393,N_9492);
nor U9501 (N_9501,N_9337,N_9370);
nand U9502 (N_9502,N_9487,N_9360);
xor U9503 (N_9503,N_9356,N_9412);
or U9504 (N_9504,N_9489,N_9343);
nor U9505 (N_9505,N_9289,N_9403);
and U9506 (N_9506,N_9365,N_9257);
or U9507 (N_9507,N_9355,N_9270);
and U9508 (N_9508,N_9452,N_9335);
or U9509 (N_9509,N_9394,N_9474);
nor U9510 (N_9510,N_9274,N_9253);
nor U9511 (N_9511,N_9451,N_9287);
and U9512 (N_9512,N_9288,N_9381);
xor U9513 (N_9513,N_9303,N_9454);
and U9514 (N_9514,N_9349,N_9329);
nand U9515 (N_9515,N_9496,N_9433);
and U9516 (N_9516,N_9357,N_9493);
nand U9517 (N_9517,N_9392,N_9453);
nor U9518 (N_9518,N_9427,N_9256);
nand U9519 (N_9519,N_9376,N_9327);
nand U9520 (N_9520,N_9374,N_9295);
xor U9521 (N_9521,N_9345,N_9318);
or U9522 (N_9522,N_9362,N_9417);
xnor U9523 (N_9523,N_9450,N_9398);
nor U9524 (N_9524,N_9435,N_9461);
or U9525 (N_9525,N_9494,N_9275);
nand U9526 (N_9526,N_9304,N_9354);
nand U9527 (N_9527,N_9254,N_9294);
nand U9528 (N_9528,N_9292,N_9322);
xnor U9529 (N_9529,N_9438,N_9323);
nand U9530 (N_9530,N_9383,N_9437);
xnor U9531 (N_9531,N_9305,N_9375);
xnor U9532 (N_9532,N_9434,N_9382);
nand U9533 (N_9533,N_9359,N_9466);
and U9534 (N_9534,N_9480,N_9273);
or U9535 (N_9535,N_9348,N_9324);
nand U9536 (N_9536,N_9314,N_9346);
or U9537 (N_9537,N_9291,N_9440);
or U9538 (N_9538,N_9262,N_9363);
nor U9539 (N_9539,N_9286,N_9421);
nand U9540 (N_9540,N_9473,N_9312);
nor U9541 (N_9541,N_9321,N_9252);
or U9542 (N_9542,N_9407,N_9366);
nand U9543 (N_9543,N_9410,N_9317);
xor U9544 (N_9544,N_9467,N_9261);
nor U9545 (N_9545,N_9499,N_9416);
or U9546 (N_9546,N_9455,N_9290);
nor U9547 (N_9547,N_9491,N_9276);
or U9548 (N_9548,N_9373,N_9353);
xor U9549 (N_9549,N_9409,N_9456);
and U9550 (N_9550,N_9478,N_9444);
nand U9551 (N_9551,N_9272,N_9255);
nand U9552 (N_9552,N_9358,N_9411);
or U9553 (N_9553,N_9333,N_9468);
and U9554 (N_9554,N_9300,N_9457);
nor U9555 (N_9555,N_9388,N_9309);
xor U9556 (N_9556,N_9250,N_9342);
or U9557 (N_9557,N_9470,N_9483);
xnor U9558 (N_9558,N_9367,N_9284);
nand U9559 (N_9559,N_9399,N_9344);
and U9560 (N_9560,N_9386,N_9296);
xnor U9561 (N_9561,N_9271,N_9269);
xnor U9562 (N_9562,N_9377,N_9465);
nor U9563 (N_9563,N_9278,N_9404);
xor U9564 (N_9564,N_9445,N_9326);
and U9565 (N_9565,N_9315,N_9330);
and U9566 (N_9566,N_9432,N_9319);
nor U9567 (N_9567,N_9280,N_9334);
and U9568 (N_9568,N_9441,N_9371);
nor U9569 (N_9569,N_9299,N_9397);
nand U9570 (N_9570,N_9482,N_9351);
or U9571 (N_9571,N_9472,N_9372);
xor U9572 (N_9572,N_9422,N_9378);
nor U9573 (N_9573,N_9268,N_9379);
xnor U9574 (N_9574,N_9396,N_9385);
nand U9575 (N_9575,N_9313,N_9395);
nand U9576 (N_9576,N_9310,N_9459);
nand U9577 (N_9577,N_9361,N_9476);
or U9578 (N_9578,N_9264,N_9419);
and U9579 (N_9579,N_9469,N_9497);
nand U9580 (N_9580,N_9259,N_9267);
nor U9581 (N_9581,N_9460,N_9265);
nand U9582 (N_9582,N_9448,N_9258);
and U9583 (N_9583,N_9443,N_9263);
nor U9584 (N_9584,N_9266,N_9339);
and U9585 (N_9585,N_9429,N_9477);
nor U9586 (N_9586,N_9402,N_9484);
xnor U9587 (N_9587,N_9281,N_9390);
or U9588 (N_9588,N_9307,N_9325);
nor U9589 (N_9589,N_9308,N_9277);
nand U9590 (N_9590,N_9302,N_9481);
or U9591 (N_9591,N_9418,N_9336);
nand U9592 (N_9592,N_9293,N_9479);
or U9593 (N_9593,N_9406,N_9340);
and U9594 (N_9594,N_9400,N_9446);
and U9595 (N_9595,N_9320,N_9331);
nor U9596 (N_9596,N_9279,N_9306);
and U9597 (N_9597,N_9369,N_9498);
or U9598 (N_9598,N_9449,N_9424);
and U9599 (N_9599,N_9486,N_9251);
nand U9600 (N_9600,N_9447,N_9408);
and U9601 (N_9601,N_9414,N_9462);
or U9602 (N_9602,N_9338,N_9436);
nand U9603 (N_9603,N_9282,N_9425);
nand U9604 (N_9604,N_9415,N_9471);
nand U9605 (N_9605,N_9328,N_9495);
nor U9606 (N_9606,N_9458,N_9389);
or U9607 (N_9607,N_9488,N_9439);
or U9608 (N_9608,N_9431,N_9332);
xor U9609 (N_9609,N_9463,N_9380);
nand U9610 (N_9610,N_9283,N_9364);
and U9611 (N_9611,N_9426,N_9285);
and U9612 (N_9612,N_9413,N_9260);
and U9613 (N_9613,N_9391,N_9347);
nor U9614 (N_9614,N_9352,N_9298);
xnor U9615 (N_9615,N_9405,N_9297);
xnor U9616 (N_9616,N_9384,N_9485);
nor U9617 (N_9617,N_9464,N_9475);
nand U9618 (N_9618,N_9350,N_9423);
or U9619 (N_9619,N_9442,N_9401);
nor U9620 (N_9620,N_9387,N_9316);
nor U9621 (N_9621,N_9430,N_9420);
nor U9622 (N_9622,N_9428,N_9368);
nor U9623 (N_9623,N_9301,N_9490);
nand U9624 (N_9624,N_9341,N_9311);
and U9625 (N_9625,N_9442,N_9340);
nor U9626 (N_9626,N_9497,N_9403);
or U9627 (N_9627,N_9308,N_9353);
nand U9628 (N_9628,N_9488,N_9478);
nand U9629 (N_9629,N_9295,N_9426);
nand U9630 (N_9630,N_9258,N_9351);
nor U9631 (N_9631,N_9293,N_9414);
and U9632 (N_9632,N_9308,N_9375);
xnor U9633 (N_9633,N_9460,N_9307);
xor U9634 (N_9634,N_9304,N_9270);
xor U9635 (N_9635,N_9346,N_9364);
xnor U9636 (N_9636,N_9457,N_9253);
or U9637 (N_9637,N_9378,N_9476);
or U9638 (N_9638,N_9328,N_9360);
nand U9639 (N_9639,N_9279,N_9295);
nand U9640 (N_9640,N_9459,N_9305);
nor U9641 (N_9641,N_9306,N_9451);
xnor U9642 (N_9642,N_9469,N_9428);
xnor U9643 (N_9643,N_9446,N_9336);
and U9644 (N_9644,N_9303,N_9446);
and U9645 (N_9645,N_9360,N_9409);
nor U9646 (N_9646,N_9447,N_9450);
xor U9647 (N_9647,N_9475,N_9311);
or U9648 (N_9648,N_9396,N_9337);
nor U9649 (N_9649,N_9466,N_9307);
nand U9650 (N_9650,N_9473,N_9392);
nand U9651 (N_9651,N_9313,N_9319);
xnor U9652 (N_9652,N_9366,N_9445);
or U9653 (N_9653,N_9271,N_9406);
nand U9654 (N_9654,N_9271,N_9426);
nor U9655 (N_9655,N_9426,N_9344);
and U9656 (N_9656,N_9459,N_9401);
xnor U9657 (N_9657,N_9320,N_9364);
nor U9658 (N_9658,N_9392,N_9427);
nor U9659 (N_9659,N_9455,N_9335);
xor U9660 (N_9660,N_9471,N_9462);
nand U9661 (N_9661,N_9460,N_9459);
or U9662 (N_9662,N_9455,N_9278);
and U9663 (N_9663,N_9404,N_9414);
or U9664 (N_9664,N_9268,N_9466);
xor U9665 (N_9665,N_9351,N_9436);
nor U9666 (N_9666,N_9416,N_9354);
or U9667 (N_9667,N_9274,N_9316);
nor U9668 (N_9668,N_9309,N_9255);
nor U9669 (N_9669,N_9326,N_9260);
nand U9670 (N_9670,N_9443,N_9459);
xnor U9671 (N_9671,N_9408,N_9378);
or U9672 (N_9672,N_9254,N_9472);
nor U9673 (N_9673,N_9261,N_9294);
nor U9674 (N_9674,N_9492,N_9317);
or U9675 (N_9675,N_9374,N_9296);
xnor U9676 (N_9676,N_9480,N_9452);
nor U9677 (N_9677,N_9405,N_9421);
or U9678 (N_9678,N_9341,N_9344);
or U9679 (N_9679,N_9454,N_9274);
or U9680 (N_9680,N_9423,N_9488);
xor U9681 (N_9681,N_9323,N_9370);
nor U9682 (N_9682,N_9438,N_9449);
nor U9683 (N_9683,N_9468,N_9345);
nand U9684 (N_9684,N_9432,N_9360);
xor U9685 (N_9685,N_9415,N_9342);
xor U9686 (N_9686,N_9352,N_9456);
xor U9687 (N_9687,N_9388,N_9253);
xor U9688 (N_9688,N_9412,N_9432);
nand U9689 (N_9689,N_9469,N_9433);
or U9690 (N_9690,N_9373,N_9407);
nor U9691 (N_9691,N_9328,N_9269);
nand U9692 (N_9692,N_9340,N_9496);
and U9693 (N_9693,N_9266,N_9475);
xnor U9694 (N_9694,N_9339,N_9414);
xor U9695 (N_9695,N_9361,N_9278);
nand U9696 (N_9696,N_9318,N_9483);
and U9697 (N_9697,N_9284,N_9309);
nand U9698 (N_9698,N_9433,N_9281);
nand U9699 (N_9699,N_9325,N_9439);
and U9700 (N_9700,N_9258,N_9363);
or U9701 (N_9701,N_9395,N_9376);
nor U9702 (N_9702,N_9423,N_9401);
and U9703 (N_9703,N_9442,N_9353);
and U9704 (N_9704,N_9390,N_9329);
nand U9705 (N_9705,N_9494,N_9327);
xor U9706 (N_9706,N_9261,N_9365);
and U9707 (N_9707,N_9369,N_9408);
xor U9708 (N_9708,N_9464,N_9445);
nor U9709 (N_9709,N_9496,N_9252);
nand U9710 (N_9710,N_9346,N_9456);
nand U9711 (N_9711,N_9451,N_9461);
nor U9712 (N_9712,N_9304,N_9424);
nand U9713 (N_9713,N_9276,N_9421);
and U9714 (N_9714,N_9331,N_9426);
or U9715 (N_9715,N_9338,N_9272);
or U9716 (N_9716,N_9452,N_9453);
or U9717 (N_9717,N_9437,N_9415);
and U9718 (N_9718,N_9332,N_9294);
or U9719 (N_9719,N_9417,N_9489);
xor U9720 (N_9720,N_9476,N_9451);
or U9721 (N_9721,N_9480,N_9413);
and U9722 (N_9722,N_9345,N_9284);
xnor U9723 (N_9723,N_9383,N_9484);
xor U9724 (N_9724,N_9362,N_9420);
xor U9725 (N_9725,N_9432,N_9351);
xnor U9726 (N_9726,N_9383,N_9260);
xnor U9727 (N_9727,N_9468,N_9365);
and U9728 (N_9728,N_9309,N_9297);
nand U9729 (N_9729,N_9381,N_9482);
and U9730 (N_9730,N_9479,N_9390);
xnor U9731 (N_9731,N_9344,N_9384);
nor U9732 (N_9732,N_9493,N_9431);
nand U9733 (N_9733,N_9323,N_9297);
nor U9734 (N_9734,N_9465,N_9288);
or U9735 (N_9735,N_9377,N_9275);
and U9736 (N_9736,N_9428,N_9426);
xor U9737 (N_9737,N_9253,N_9475);
or U9738 (N_9738,N_9272,N_9421);
and U9739 (N_9739,N_9407,N_9393);
and U9740 (N_9740,N_9456,N_9471);
or U9741 (N_9741,N_9439,N_9289);
nand U9742 (N_9742,N_9263,N_9271);
nand U9743 (N_9743,N_9465,N_9297);
and U9744 (N_9744,N_9327,N_9408);
or U9745 (N_9745,N_9435,N_9279);
and U9746 (N_9746,N_9495,N_9443);
and U9747 (N_9747,N_9405,N_9373);
xor U9748 (N_9748,N_9291,N_9427);
nand U9749 (N_9749,N_9491,N_9313);
xnor U9750 (N_9750,N_9541,N_9689);
or U9751 (N_9751,N_9570,N_9700);
or U9752 (N_9752,N_9563,N_9710);
and U9753 (N_9753,N_9698,N_9505);
and U9754 (N_9754,N_9509,N_9666);
and U9755 (N_9755,N_9667,N_9711);
nor U9756 (N_9756,N_9506,N_9669);
xnor U9757 (N_9757,N_9683,N_9713);
nand U9758 (N_9758,N_9718,N_9609);
nand U9759 (N_9759,N_9625,N_9673);
and U9760 (N_9760,N_9661,N_9626);
nor U9761 (N_9761,N_9548,N_9603);
nand U9762 (N_9762,N_9672,N_9627);
nand U9763 (N_9763,N_9720,N_9599);
and U9764 (N_9764,N_9679,N_9643);
nand U9765 (N_9765,N_9724,N_9630);
xor U9766 (N_9766,N_9633,N_9567);
and U9767 (N_9767,N_9604,N_9642);
xnor U9768 (N_9768,N_9629,N_9534);
or U9769 (N_9769,N_9547,N_9621);
or U9770 (N_9770,N_9613,N_9516);
xor U9771 (N_9771,N_9717,N_9656);
xnor U9772 (N_9772,N_9631,N_9514);
nor U9773 (N_9773,N_9701,N_9746);
nand U9774 (N_9774,N_9727,N_9688);
nand U9775 (N_9775,N_9686,N_9645);
xor U9776 (N_9776,N_9678,N_9602);
nand U9777 (N_9777,N_9663,N_9530);
xnor U9778 (N_9778,N_9576,N_9716);
nor U9779 (N_9779,N_9522,N_9564);
and U9780 (N_9780,N_9634,N_9691);
or U9781 (N_9781,N_9612,N_9513);
nand U9782 (N_9782,N_9674,N_9715);
nor U9783 (N_9783,N_9702,N_9590);
xor U9784 (N_9784,N_9744,N_9502);
nand U9785 (N_9785,N_9741,N_9620);
and U9786 (N_9786,N_9580,N_9721);
nor U9787 (N_9787,N_9649,N_9521);
xnor U9788 (N_9788,N_9740,N_9670);
nor U9789 (N_9789,N_9703,N_9664);
xor U9790 (N_9790,N_9719,N_9519);
and U9791 (N_9791,N_9520,N_9552);
nand U9792 (N_9792,N_9550,N_9589);
xor U9793 (N_9793,N_9668,N_9592);
nor U9794 (N_9794,N_9704,N_9554);
nor U9795 (N_9795,N_9714,N_9615);
nand U9796 (N_9796,N_9601,N_9595);
xnor U9797 (N_9797,N_9648,N_9729);
or U9798 (N_9798,N_9539,N_9690);
xor U9799 (N_9799,N_9597,N_9532);
nand U9800 (N_9800,N_9560,N_9680);
nand U9801 (N_9801,N_9579,N_9685);
and U9802 (N_9802,N_9538,N_9739);
and U9803 (N_9803,N_9556,N_9731);
nor U9804 (N_9804,N_9503,N_9583);
and U9805 (N_9805,N_9593,N_9549);
or U9806 (N_9806,N_9641,N_9693);
xor U9807 (N_9807,N_9571,N_9684);
or U9808 (N_9808,N_9518,N_9640);
and U9809 (N_9809,N_9585,N_9540);
xor U9810 (N_9810,N_9591,N_9699);
nor U9811 (N_9811,N_9543,N_9728);
and U9812 (N_9812,N_9558,N_9695);
xor U9813 (N_9813,N_9588,N_9551);
or U9814 (N_9814,N_9510,N_9594);
xnor U9815 (N_9815,N_9737,N_9681);
and U9816 (N_9816,N_9565,N_9608);
xor U9817 (N_9817,N_9676,N_9636);
nor U9818 (N_9818,N_9742,N_9722);
xnor U9819 (N_9819,N_9557,N_9586);
xor U9820 (N_9820,N_9660,N_9692);
or U9821 (N_9821,N_9525,N_9581);
and U9822 (N_9822,N_9677,N_9638);
or U9823 (N_9823,N_9652,N_9682);
and U9824 (N_9824,N_9651,N_9561);
or U9825 (N_9825,N_9524,N_9584);
and U9826 (N_9826,N_9743,N_9533);
and U9827 (N_9827,N_9568,N_9712);
nor U9828 (N_9828,N_9596,N_9528);
or U9829 (N_9829,N_9536,N_9733);
xor U9830 (N_9830,N_9734,N_9500);
or U9831 (N_9831,N_9559,N_9607);
xnor U9832 (N_9832,N_9578,N_9515);
nor U9833 (N_9833,N_9706,N_9582);
or U9834 (N_9834,N_9575,N_9738);
and U9835 (N_9835,N_9749,N_9555);
or U9836 (N_9836,N_9696,N_9605);
xnor U9837 (N_9837,N_9598,N_9523);
nand U9838 (N_9838,N_9730,N_9527);
xor U9839 (N_9839,N_9616,N_9647);
nor U9840 (N_9840,N_9635,N_9507);
or U9841 (N_9841,N_9657,N_9619);
nand U9842 (N_9842,N_9512,N_9707);
nand U9843 (N_9843,N_9662,N_9517);
or U9844 (N_9844,N_9573,N_9725);
or U9845 (N_9845,N_9735,N_9617);
and U9846 (N_9846,N_9600,N_9610);
xnor U9847 (N_9847,N_9542,N_9697);
nand U9848 (N_9848,N_9562,N_9659);
and U9849 (N_9849,N_9709,N_9569);
nor U9850 (N_9850,N_9732,N_9526);
and U9851 (N_9851,N_9611,N_9574);
nand U9852 (N_9852,N_9748,N_9622);
and U9853 (N_9853,N_9535,N_9726);
xnor U9854 (N_9854,N_9618,N_9665);
and U9855 (N_9855,N_9504,N_9546);
nand U9856 (N_9856,N_9694,N_9736);
nand U9857 (N_9857,N_9658,N_9646);
xnor U9858 (N_9858,N_9614,N_9708);
and U9859 (N_9859,N_9537,N_9587);
and U9860 (N_9860,N_9637,N_9644);
xnor U9861 (N_9861,N_9531,N_9639);
xor U9862 (N_9862,N_9747,N_9529);
and U9863 (N_9863,N_9654,N_9553);
and U9864 (N_9864,N_9671,N_9705);
or U9865 (N_9865,N_9508,N_9572);
nand U9866 (N_9866,N_9544,N_9687);
or U9867 (N_9867,N_9511,N_9566);
and U9868 (N_9868,N_9745,N_9545);
nor U9869 (N_9869,N_9632,N_9675);
and U9870 (N_9870,N_9606,N_9623);
nor U9871 (N_9871,N_9501,N_9655);
nor U9872 (N_9872,N_9723,N_9650);
nand U9873 (N_9873,N_9653,N_9624);
nand U9874 (N_9874,N_9577,N_9628);
nand U9875 (N_9875,N_9606,N_9636);
xnor U9876 (N_9876,N_9565,N_9630);
xnor U9877 (N_9877,N_9593,N_9628);
and U9878 (N_9878,N_9503,N_9661);
nand U9879 (N_9879,N_9721,N_9734);
xnor U9880 (N_9880,N_9702,N_9555);
xor U9881 (N_9881,N_9708,N_9707);
nor U9882 (N_9882,N_9678,N_9627);
nand U9883 (N_9883,N_9513,N_9663);
nor U9884 (N_9884,N_9636,N_9526);
nand U9885 (N_9885,N_9748,N_9559);
nand U9886 (N_9886,N_9535,N_9540);
or U9887 (N_9887,N_9582,N_9720);
nand U9888 (N_9888,N_9607,N_9503);
or U9889 (N_9889,N_9540,N_9732);
xnor U9890 (N_9890,N_9716,N_9617);
nor U9891 (N_9891,N_9560,N_9723);
or U9892 (N_9892,N_9661,N_9720);
nand U9893 (N_9893,N_9613,N_9673);
nand U9894 (N_9894,N_9540,N_9740);
xor U9895 (N_9895,N_9504,N_9595);
nand U9896 (N_9896,N_9684,N_9575);
or U9897 (N_9897,N_9688,N_9612);
or U9898 (N_9898,N_9552,N_9648);
and U9899 (N_9899,N_9511,N_9525);
and U9900 (N_9900,N_9635,N_9506);
and U9901 (N_9901,N_9740,N_9657);
nand U9902 (N_9902,N_9746,N_9687);
nor U9903 (N_9903,N_9529,N_9594);
and U9904 (N_9904,N_9717,N_9636);
xor U9905 (N_9905,N_9669,N_9524);
and U9906 (N_9906,N_9713,N_9523);
or U9907 (N_9907,N_9701,N_9623);
nand U9908 (N_9908,N_9555,N_9618);
nand U9909 (N_9909,N_9695,N_9692);
and U9910 (N_9910,N_9609,N_9746);
nor U9911 (N_9911,N_9675,N_9536);
and U9912 (N_9912,N_9602,N_9720);
nor U9913 (N_9913,N_9514,N_9523);
or U9914 (N_9914,N_9529,N_9552);
xor U9915 (N_9915,N_9706,N_9665);
xor U9916 (N_9916,N_9660,N_9557);
or U9917 (N_9917,N_9715,N_9694);
or U9918 (N_9918,N_9704,N_9583);
xor U9919 (N_9919,N_9578,N_9671);
and U9920 (N_9920,N_9662,N_9714);
or U9921 (N_9921,N_9564,N_9682);
nor U9922 (N_9922,N_9546,N_9614);
nand U9923 (N_9923,N_9607,N_9606);
and U9924 (N_9924,N_9575,N_9560);
xor U9925 (N_9925,N_9706,N_9608);
nand U9926 (N_9926,N_9656,N_9700);
and U9927 (N_9927,N_9605,N_9692);
or U9928 (N_9928,N_9607,N_9692);
xor U9929 (N_9929,N_9740,N_9638);
xnor U9930 (N_9930,N_9598,N_9603);
xnor U9931 (N_9931,N_9567,N_9716);
xor U9932 (N_9932,N_9572,N_9714);
or U9933 (N_9933,N_9666,N_9637);
and U9934 (N_9934,N_9528,N_9577);
or U9935 (N_9935,N_9695,N_9669);
nand U9936 (N_9936,N_9585,N_9559);
or U9937 (N_9937,N_9590,N_9555);
and U9938 (N_9938,N_9574,N_9737);
or U9939 (N_9939,N_9742,N_9601);
xnor U9940 (N_9940,N_9606,N_9661);
and U9941 (N_9941,N_9674,N_9698);
nor U9942 (N_9942,N_9670,N_9563);
and U9943 (N_9943,N_9609,N_9557);
and U9944 (N_9944,N_9667,N_9547);
xnor U9945 (N_9945,N_9640,N_9646);
and U9946 (N_9946,N_9532,N_9518);
and U9947 (N_9947,N_9548,N_9642);
nand U9948 (N_9948,N_9545,N_9719);
xor U9949 (N_9949,N_9634,N_9637);
xnor U9950 (N_9950,N_9691,N_9669);
nand U9951 (N_9951,N_9690,N_9671);
xnor U9952 (N_9952,N_9695,N_9630);
or U9953 (N_9953,N_9528,N_9626);
nor U9954 (N_9954,N_9574,N_9681);
xor U9955 (N_9955,N_9537,N_9720);
nand U9956 (N_9956,N_9515,N_9723);
and U9957 (N_9957,N_9566,N_9625);
nand U9958 (N_9958,N_9604,N_9510);
nand U9959 (N_9959,N_9614,N_9633);
or U9960 (N_9960,N_9569,N_9727);
and U9961 (N_9961,N_9510,N_9533);
xor U9962 (N_9962,N_9689,N_9539);
and U9963 (N_9963,N_9748,N_9679);
or U9964 (N_9964,N_9568,N_9540);
xnor U9965 (N_9965,N_9692,N_9703);
nor U9966 (N_9966,N_9564,N_9698);
nand U9967 (N_9967,N_9675,N_9542);
and U9968 (N_9968,N_9563,N_9611);
nor U9969 (N_9969,N_9566,N_9675);
xor U9970 (N_9970,N_9587,N_9584);
and U9971 (N_9971,N_9664,N_9545);
nor U9972 (N_9972,N_9619,N_9637);
and U9973 (N_9973,N_9578,N_9530);
nand U9974 (N_9974,N_9515,N_9646);
or U9975 (N_9975,N_9612,N_9678);
or U9976 (N_9976,N_9670,N_9637);
xor U9977 (N_9977,N_9737,N_9630);
nand U9978 (N_9978,N_9555,N_9685);
nor U9979 (N_9979,N_9725,N_9669);
xor U9980 (N_9980,N_9673,N_9594);
nor U9981 (N_9981,N_9541,N_9745);
and U9982 (N_9982,N_9611,N_9687);
nor U9983 (N_9983,N_9695,N_9656);
and U9984 (N_9984,N_9569,N_9572);
nand U9985 (N_9985,N_9665,N_9579);
nand U9986 (N_9986,N_9583,N_9684);
nor U9987 (N_9987,N_9655,N_9558);
xnor U9988 (N_9988,N_9724,N_9685);
nand U9989 (N_9989,N_9603,N_9617);
nand U9990 (N_9990,N_9623,N_9745);
nand U9991 (N_9991,N_9729,N_9587);
nand U9992 (N_9992,N_9602,N_9598);
nand U9993 (N_9993,N_9549,N_9672);
xor U9994 (N_9994,N_9609,N_9627);
xor U9995 (N_9995,N_9632,N_9664);
and U9996 (N_9996,N_9733,N_9644);
and U9997 (N_9997,N_9663,N_9644);
nand U9998 (N_9998,N_9649,N_9539);
or U9999 (N_9999,N_9737,N_9529);
or U10000 (N_10000,N_9799,N_9946);
xnor U10001 (N_10001,N_9967,N_9778);
or U10002 (N_10002,N_9986,N_9810);
or U10003 (N_10003,N_9786,N_9871);
nor U10004 (N_10004,N_9954,N_9836);
nand U10005 (N_10005,N_9848,N_9780);
and U10006 (N_10006,N_9856,N_9789);
xnor U10007 (N_10007,N_9842,N_9998);
and U10008 (N_10008,N_9797,N_9942);
and U10009 (N_10009,N_9760,N_9866);
or U10010 (N_10010,N_9944,N_9765);
nor U10011 (N_10011,N_9817,N_9870);
nor U10012 (N_10012,N_9880,N_9812);
xor U10013 (N_10013,N_9827,N_9968);
and U10014 (N_10014,N_9845,N_9888);
nor U10015 (N_10015,N_9966,N_9941);
nand U10016 (N_10016,N_9805,N_9816);
nand U10017 (N_10017,N_9793,N_9985);
nor U10018 (N_10018,N_9838,N_9791);
nand U10019 (N_10019,N_9973,N_9847);
or U10020 (N_10020,N_9914,N_9751);
nor U10021 (N_10021,N_9795,N_9806);
or U10022 (N_10022,N_9863,N_9932);
and U10023 (N_10023,N_9950,N_9821);
or U10024 (N_10024,N_9775,N_9777);
nand U10025 (N_10025,N_9965,N_9908);
xor U10026 (N_10026,N_9918,N_9983);
xnor U10027 (N_10027,N_9974,N_9811);
or U10028 (N_10028,N_9926,N_9959);
nor U10029 (N_10029,N_9996,N_9921);
nor U10030 (N_10030,N_9882,N_9952);
xor U10031 (N_10031,N_9898,N_9976);
nand U10032 (N_10032,N_9879,N_9840);
nand U10033 (N_10033,N_9909,N_9906);
xnor U10034 (N_10034,N_9872,N_9958);
nor U10035 (N_10035,N_9955,N_9960);
and U10036 (N_10036,N_9802,N_9990);
and U10037 (N_10037,N_9864,N_9970);
or U10038 (N_10038,N_9943,N_9800);
xor U10039 (N_10039,N_9972,N_9759);
xnor U10040 (N_10040,N_9766,N_9887);
or U10041 (N_10041,N_9915,N_9770);
nor U10042 (N_10042,N_9991,N_9815);
nor U10043 (N_10043,N_9822,N_9999);
and U10044 (N_10044,N_9979,N_9889);
xor U10045 (N_10045,N_9782,N_9831);
or U10046 (N_10046,N_9933,N_9892);
nor U10047 (N_10047,N_9884,N_9792);
and U10048 (N_10048,N_9774,N_9833);
xnor U10049 (N_10049,N_9935,N_9794);
nand U10050 (N_10050,N_9784,N_9773);
nand U10051 (N_10051,N_9807,N_9790);
nand U10052 (N_10052,N_9982,N_9953);
nor U10053 (N_10053,N_9993,N_9891);
xor U10054 (N_10054,N_9750,N_9895);
nand U10055 (N_10055,N_9951,N_9803);
and U10056 (N_10056,N_9936,N_9772);
nor U10057 (N_10057,N_9981,N_9910);
nor U10058 (N_10058,N_9828,N_9969);
xor U10059 (N_10059,N_9861,N_9937);
nand U10060 (N_10060,N_9930,N_9894);
and U10061 (N_10061,N_9855,N_9896);
and U10062 (N_10062,N_9992,N_9925);
nor U10063 (N_10063,N_9885,N_9850);
xor U10064 (N_10064,N_9771,N_9754);
or U10065 (N_10065,N_9874,N_9913);
or U10066 (N_10066,N_9801,N_9901);
xnor U10067 (N_10067,N_9826,N_9940);
nor U10068 (N_10068,N_9897,N_9912);
nor U10069 (N_10069,N_9938,N_9758);
xor U10070 (N_10070,N_9869,N_9858);
nand U10071 (N_10071,N_9929,N_9988);
xor U10072 (N_10072,N_9776,N_9862);
nand U10073 (N_10073,N_9948,N_9767);
nor U10074 (N_10074,N_9907,N_9829);
and U10075 (N_10075,N_9779,N_9798);
nand U10076 (N_10076,N_9964,N_9867);
or U10077 (N_10077,N_9824,N_9919);
xnor U10078 (N_10078,N_9844,N_9788);
and U10079 (N_10079,N_9752,N_9939);
nand U10080 (N_10080,N_9813,N_9804);
and U10081 (N_10081,N_9873,N_9865);
nor U10082 (N_10082,N_9934,N_9823);
xnor U10083 (N_10083,N_9854,N_9947);
nor U10084 (N_10084,N_9753,N_9890);
nand U10085 (N_10085,N_9984,N_9920);
and U10086 (N_10086,N_9860,N_9927);
and U10087 (N_10087,N_9846,N_9837);
or U10088 (N_10088,N_9785,N_9851);
or U10089 (N_10089,N_9928,N_9916);
xnor U10090 (N_10090,N_9899,N_9963);
xnor U10091 (N_10091,N_9841,N_9980);
and U10092 (N_10092,N_9769,N_9755);
nor U10093 (N_10093,N_9905,N_9849);
xor U10094 (N_10094,N_9975,N_9878);
and U10095 (N_10095,N_9764,N_9995);
and U10096 (N_10096,N_9768,N_9757);
or U10097 (N_10097,N_9917,N_9922);
xor U10098 (N_10098,N_9971,N_9904);
nor U10099 (N_10099,N_9814,N_9977);
and U10100 (N_10100,N_9957,N_9818);
xnor U10101 (N_10101,N_9994,N_9945);
nor U10102 (N_10102,N_9809,N_9883);
nor U10103 (N_10103,N_9881,N_9911);
and U10104 (N_10104,N_9808,N_9825);
xor U10105 (N_10105,N_9893,N_9877);
nor U10106 (N_10106,N_9857,N_9781);
or U10107 (N_10107,N_9819,N_9834);
xor U10108 (N_10108,N_9761,N_9832);
nand U10109 (N_10109,N_9839,N_9859);
nand U10110 (N_10110,N_9989,N_9949);
or U10111 (N_10111,N_9853,N_9820);
nand U10112 (N_10112,N_9987,N_9835);
nand U10113 (N_10113,N_9924,N_9783);
nand U10114 (N_10114,N_9868,N_9763);
xnor U10115 (N_10115,N_9900,N_9796);
nor U10116 (N_10116,N_9956,N_9903);
or U10117 (N_10117,N_9852,N_9876);
nor U10118 (N_10118,N_9931,N_9978);
and U10119 (N_10119,N_9830,N_9962);
or U10120 (N_10120,N_9787,N_9886);
nor U10121 (N_10121,N_9762,N_9997);
nor U10122 (N_10122,N_9923,N_9843);
xnor U10123 (N_10123,N_9756,N_9875);
nor U10124 (N_10124,N_9902,N_9961);
nor U10125 (N_10125,N_9760,N_9751);
nor U10126 (N_10126,N_9933,N_9887);
xnor U10127 (N_10127,N_9795,N_9778);
nor U10128 (N_10128,N_9986,N_9870);
or U10129 (N_10129,N_9989,N_9856);
nor U10130 (N_10130,N_9751,N_9997);
and U10131 (N_10131,N_9902,N_9916);
and U10132 (N_10132,N_9876,N_9939);
or U10133 (N_10133,N_9891,N_9814);
nand U10134 (N_10134,N_9859,N_9808);
and U10135 (N_10135,N_9909,N_9903);
and U10136 (N_10136,N_9842,N_9841);
or U10137 (N_10137,N_9955,N_9863);
and U10138 (N_10138,N_9840,N_9959);
and U10139 (N_10139,N_9756,N_9806);
or U10140 (N_10140,N_9852,N_9917);
and U10141 (N_10141,N_9786,N_9800);
nand U10142 (N_10142,N_9754,N_9855);
and U10143 (N_10143,N_9810,N_9816);
or U10144 (N_10144,N_9838,N_9970);
nand U10145 (N_10145,N_9890,N_9997);
xnor U10146 (N_10146,N_9965,N_9822);
xnor U10147 (N_10147,N_9771,N_9979);
and U10148 (N_10148,N_9779,N_9807);
or U10149 (N_10149,N_9812,N_9855);
nor U10150 (N_10150,N_9975,N_9949);
nand U10151 (N_10151,N_9866,N_9972);
nor U10152 (N_10152,N_9925,N_9926);
xnor U10153 (N_10153,N_9791,N_9830);
xor U10154 (N_10154,N_9998,N_9860);
nor U10155 (N_10155,N_9916,N_9917);
and U10156 (N_10156,N_9783,N_9804);
xnor U10157 (N_10157,N_9918,N_9807);
or U10158 (N_10158,N_9765,N_9842);
xor U10159 (N_10159,N_9922,N_9942);
and U10160 (N_10160,N_9867,N_9757);
and U10161 (N_10161,N_9886,N_9999);
nand U10162 (N_10162,N_9784,N_9968);
nor U10163 (N_10163,N_9840,N_9798);
and U10164 (N_10164,N_9863,N_9815);
nor U10165 (N_10165,N_9891,N_9750);
or U10166 (N_10166,N_9750,N_9784);
nor U10167 (N_10167,N_9939,N_9773);
nor U10168 (N_10168,N_9930,N_9803);
and U10169 (N_10169,N_9776,N_9757);
and U10170 (N_10170,N_9831,N_9936);
nand U10171 (N_10171,N_9912,N_9777);
or U10172 (N_10172,N_9783,N_9981);
or U10173 (N_10173,N_9838,N_9968);
nor U10174 (N_10174,N_9886,N_9829);
or U10175 (N_10175,N_9976,N_9961);
nand U10176 (N_10176,N_9910,N_9813);
or U10177 (N_10177,N_9906,N_9960);
or U10178 (N_10178,N_9908,N_9907);
nor U10179 (N_10179,N_9893,N_9968);
nor U10180 (N_10180,N_9849,N_9933);
and U10181 (N_10181,N_9800,N_9878);
or U10182 (N_10182,N_9938,N_9772);
xnor U10183 (N_10183,N_9993,N_9999);
xnor U10184 (N_10184,N_9825,N_9759);
and U10185 (N_10185,N_9790,N_9776);
nand U10186 (N_10186,N_9808,N_9915);
or U10187 (N_10187,N_9975,N_9753);
nand U10188 (N_10188,N_9756,N_9757);
xor U10189 (N_10189,N_9783,N_9939);
nor U10190 (N_10190,N_9823,N_9965);
nor U10191 (N_10191,N_9957,N_9779);
nand U10192 (N_10192,N_9931,N_9909);
nand U10193 (N_10193,N_9903,N_9846);
nor U10194 (N_10194,N_9756,N_9853);
nand U10195 (N_10195,N_9824,N_9938);
xor U10196 (N_10196,N_9885,N_9897);
and U10197 (N_10197,N_9758,N_9815);
nand U10198 (N_10198,N_9876,N_9930);
nor U10199 (N_10199,N_9872,N_9877);
xor U10200 (N_10200,N_9975,N_9866);
nor U10201 (N_10201,N_9916,N_9980);
nor U10202 (N_10202,N_9829,N_9929);
nand U10203 (N_10203,N_9831,N_9859);
or U10204 (N_10204,N_9815,N_9929);
xnor U10205 (N_10205,N_9929,N_9883);
and U10206 (N_10206,N_9827,N_9880);
or U10207 (N_10207,N_9946,N_9944);
or U10208 (N_10208,N_9916,N_9752);
and U10209 (N_10209,N_9921,N_9760);
or U10210 (N_10210,N_9997,N_9945);
or U10211 (N_10211,N_9860,N_9880);
nor U10212 (N_10212,N_9851,N_9857);
nand U10213 (N_10213,N_9781,N_9923);
or U10214 (N_10214,N_9790,N_9829);
or U10215 (N_10215,N_9758,N_9817);
or U10216 (N_10216,N_9755,N_9910);
and U10217 (N_10217,N_9874,N_9991);
and U10218 (N_10218,N_9952,N_9775);
and U10219 (N_10219,N_9872,N_9873);
xnor U10220 (N_10220,N_9982,N_9906);
xnor U10221 (N_10221,N_9815,N_9789);
and U10222 (N_10222,N_9973,N_9878);
xnor U10223 (N_10223,N_9944,N_9791);
nand U10224 (N_10224,N_9965,N_9918);
or U10225 (N_10225,N_9966,N_9958);
nor U10226 (N_10226,N_9990,N_9873);
and U10227 (N_10227,N_9913,N_9947);
nor U10228 (N_10228,N_9810,N_9824);
nor U10229 (N_10229,N_9911,N_9988);
and U10230 (N_10230,N_9934,N_9871);
nand U10231 (N_10231,N_9948,N_9991);
nor U10232 (N_10232,N_9811,N_9822);
nor U10233 (N_10233,N_9781,N_9888);
nor U10234 (N_10234,N_9935,N_9767);
xnor U10235 (N_10235,N_9987,N_9818);
or U10236 (N_10236,N_9755,N_9967);
nand U10237 (N_10237,N_9852,N_9943);
and U10238 (N_10238,N_9755,N_9875);
and U10239 (N_10239,N_9900,N_9982);
nor U10240 (N_10240,N_9858,N_9911);
or U10241 (N_10241,N_9876,N_9842);
or U10242 (N_10242,N_9823,N_9762);
nand U10243 (N_10243,N_9884,N_9891);
nor U10244 (N_10244,N_9917,N_9809);
or U10245 (N_10245,N_9940,N_9873);
xor U10246 (N_10246,N_9808,N_9792);
nand U10247 (N_10247,N_9773,N_9956);
xor U10248 (N_10248,N_9889,N_9918);
nand U10249 (N_10249,N_9887,N_9968);
or U10250 (N_10250,N_10062,N_10193);
xnor U10251 (N_10251,N_10150,N_10156);
xnor U10252 (N_10252,N_10124,N_10011);
and U10253 (N_10253,N_10007,N_10036);
nand U10254 (N_10254,N_10227,N_10096);
or U10255 (N_10255,N_10022,N_10089);
nand U10256 (N_10256,N_10132,N_10231);
or U10257 (N_10257,N_10017,N_10186);
or U10258 (N_10258,N_10087,N_10113);
and U10259 (N_10259,N_10091,N_10063);
nor U10260 (N_10260,N_10086,N_10243);
nand U10261 (N_10261,N_10176,N_10056);
or U10262 (N_10262,N_10126,N_10211);
nor U10263 (N_10263,N_10027,N_10230);
nor U10264 (N_10264,N_10109,N_10141);
or U10265 (N_10265,N_10078,N_10170);
xor U10266 (N_10266,N_10065,N_10127);
nor U10267 (N_10267,N_10025,N_10019);
nand U10268 (N_10268,N_10135,N_10202);
nor U10269 (N_10269,N_10140,N_10210);
nand U10270 (N_10270,N_10146,N_10072);
nand U10271 (N_10271,N_10052,N_10131);
xor U10272 (N_10272,N_10160,N_10178);
xnor U10273 (N_10273,N_10249,N_10067);
nor U10274 (N_10274,N_10004,N_10058);
or U10275 (N_10275,N_10026,N_10246);
xor U10276 (N_10276,N_10165,N_10028);
nor U10277 (N_10277,N_10204,N_10155);
or U10278 (N_10278,N_10020,N_10023);
nand U10279 (N_10279,N_10203,N_10185);
and U10280 (N_10280,N_10112,N_10125);
or U10281 (N_10281,N_10081,N_10181);
nand U10282 (N_10282,N_10094,N_10157);
and U10283 (N_10283,N_10054,N_10130);
nor U10284 (N_10284,N_10162,N_10082);
xnor U10285 (N_10285,N_10044,N_10158);
nand U10286 (N_10286,N_10198,N_10134);
and U10287 (N_10287,N_10201,N_10092);
nand U10288 (N_10288,N_10048,N_10171);
and U10289 (N_10289,N_10049,N_10166);
and U10290 (N_10290,N_10111,N_10079);
nor U10291 (N_10291,N_10104,N_10161);
or U10292 (N_10292,N_10245,N_10115);
nand U10293 (N_10293,N_10199,N_10235);
nor U10294 (N_10294,N_10122,N_10241);
or U10295 (N_10295,N_10217,N_10233);
or U10296 (N_10296,N_10205,N_10090);
nand U10297 (N_10297,N_10148,N_10110);
xor U10298 (N_10298,N_10064,N_10190);
or U10299 (N_10299,N_10041,N_10183);
nand U10300 (N_10300,N_10207,N_10038);
xnor U10301 (N_10301,N_10219,N_10239);
or U10302 (N_10302,N_10014,N_10191);
nor U10303 (N_10303,N_10060,N_10013);
nor U10304 (N_10304,N_10214,N_10221);
nand U10305 (N_10305,N_10075,N_10105);
xnor U10306 (N_10306,N_10120,N_10169);
xnor U10307 (N_10307,N_10189,N_10173);
nand U10308 (N_10308,N_10143,N_10145);
and U10309 (N_10309,N_10024,N_10128);
xnor U10310 (N_10310,N_10192,N_10206);
xor U10311 (N_10311,N_10047,N_10200);
xor U10312 (N_10312,N_10084,N_10240);
xnor U10313 (N_10313,N_10144,N_10172);
nor U10314 (N_10314,N_10061,N_10077);
and U10315 (N_10315,N_10224,N_10142);
or U10316 (N_10316,N_10010,N_10175);
and U10317 (N_10317,N_10008,N_10196);
and U10318 (N_10318,N_10238,N_10103);
or U10319 (N_10319,N_10030,N_10147);
and U10320 (N_10320,N_10001,N_10118);
xnor U10321 (N_10321,N_10129,N_10194);
and U10322 (N_10322,N_10042,N_10153);
nand U10323 (N_10323,N_10248,N_10133);
nand U10324 (N_10324,N_10182,N_10216);
xnor U10325 (N_10325,N_10114,N_10034);
nand U10326 (N_10326,N_10039,N_10225);
or U10327 (N_10327,N_10102,N_10098);
xnor U10328 (N_10328,N_10040,N_10016);
and U10329 (N_10329,N_10237,N_10119);
or U10330 (N_10330,N_10074,N_10123);
nand U10331 (N_10331,N_10076,N_10244);
nand U10332 (N_10332,N_10003,N_10242);
xnor U10333 (N_10333,N_10232,N_10220);
nor U10334 (N_10334,N_10117,N_10021);
nor U10335 (N_10335,N_10197,N_10050);
nor U10336 (N_10336,N_10136,N_10159);
nand U10337 (N_10337,N_10223,N_10187);
xor U10338 (N_10338,N_10057,N_10121);
xor U10339 (N_10339,N_10035,N_10138);
or U10340 (N_10340,N_10149,N_10229);
and U10341 (N_10341,N_10000,N_10071);
nand U10342 (N_10342,N_10085,N_10095);
or U10343 (N_10343,N_10107,N_10116);
nand U10344 (N_10344,N_10046,N_10099);
xnor U10345 (N_10345,N_10073,N_10066);
nand U10346 (N_10346,N_10208,N_10247);
nand U10347 (N_10347,N_10051,N_10083);
and U10348 (N_10348,N_10033,N_10228);
and U10349 (N_10349,N_10222,N_10002);
and U10350 (N_10350,N_10031,N_10045);
and U10351 (N_10351,N_10101,N_10195);
xnor U10352 (N_10352,N_10100,N_10218);
nor U10353 (N_10353,N_10088,N_10069);
nor U10354 (N_10354,N_10009,N_10108);
nand U10355 (N_10355,N_10037,N_10137);
and U10356 (N_10356,N_10032,N_10070);
or U10357 (N_10357,N_10180,N_10012);
nand U10358 (N_10358,N_10093,N_10053);
or U10359 (N_10359,N_10018,N_10188);
nor U10360 (N_10360,N_10163,N_10055);
nand U10361 (N_10361,N_10029,N_10209);
or U10362 (N_10362,N_10080,N_10213);
or U10363 (N_10363,N_10179,N_10152);
nor U10364 (N_10364,N_10015,N_10068);
nor U10365 (N_10365,N_10215,N_10097);
or U10366 (N_10366,N_10184,N_10005);
or U10367 (N_10367,N_10168,N_10164);
nor U10368 (N_10368,N_10139,N_10043);
xor U10369 (N_10369,N_10226,N_10059);
nor U10370 (N_10370,N_10212,N_10006);
nand U10371 (N_10371,N_10151,N_10177);
or U10372 (N_10372,N_10234,N_10167);
nand U10373 (N_10373,N_10154,N_10174);
or U10374 (N_10374,N_10236,N_10106);
nand U10375 (N_10375,N_10050,N_10205);
nor U10376 (N_10376,N_10034,N_10187);
and U10377 (N_10377,N_10180,N_10249);
xor U10378 (N_10378,N_10222,N_10163);
and U10379 (N_10379,N_10240,N_10159);
xor U10380 (N_10380,N_10095,N_10030);
or U10381 (N_10381,N_10183,N_10026);
xnor U10382 (N_10382,N_10217,N_10062);
nor U10383 (N_10383,N_10198,N_10035);
nand U10384 (N_10384,N_10203,N_10009);
xnor U10385 (N_10385,N_10094,N_10002);
xor U10386 (N_10386,N_10131,N_10030);
and U10387 (N_10387,N_10108,N_10159);
nor U10388 (N_10388,N_10118,N_10211);
nor U10389 (N_10389,N_10233,N_10246);
xor U10390 (N_10390,N_10134,N_10203);
and U10391 (N_10391,N_10146,N_10189);
nor U10392 (N_10392,N_10141,N_10123);
xnor U10393 (N_10393,N_10203,N_10019);
and U10394 (N_10394,N_10143,N_10140);
nor U10395 (N_10395,N_10050,N_10238);
or U10396 (N_10396,N_10026,N_10162);
xor U10397 (N_10397,N_10086,N_10043);
or U10398 (N_10398,N_10002,N_10173);
nor U10399 (N_10399,N_10241,N_10213);
nor U10400 (N_10400,N_10014,N_10229);
or U10401 (N_10401,N_10021,N_10146);
or U10402 (N_10402,N_10100,N_10121);
nor U10403 (N_10403,N_10241,N_10113);
and U10404 (N_10404,N_10248,N_10041);
or U10405 (N_10405,N_10070,N_10065);
xor U10406 (N_10406,N_10243,N_10146);
nand U10407 (N_10407,N_10156,N_10127);
or U10408 (N_10408,N_10052,N_10233);
nor U10409 (N_10409,N_10043,N_10057);
xor U10410 (N_10410,N_10110,N_10009);
nor U10411 (N_10411,N_10116,N_10225);
or U10412 (N_10412,N_10085,N_10143);
nor U10413 (N_10413,N_10014,N_10146);
nor U10414 (N_10414,N_10218,N_10081);
or U10415 (N_10415,N_10157,N_10036);
nor U10416 (N_10416,N_10063,N_10130);
and U10417 (N_10417,N_10166,N_10199);
or U10418 (N_10418,N_10179,N_10223);
and U10419 (N_10419,N_10114,N_10046);
nand U10420 (N_10420,N_10135,N_10099);
xor U10421 (N_10421,N_10215,N_10214);
and U10422 (N_10422,N_10087,N_10245);
or U10423 (N_10423,N_10184,N_10057);
nor U10424 (N_10424,N_10220,N_10150);
or U10425 (N_10425,N_10144,N_10064);
or U10426 (N_10426,N_10103,N_10030);
or U10427 (N_10427,N_10205,N_10169);
xnor U10428 (N_10428,N_10190,N_10162);
and U10429 (N_10429,N_10060,N_10235);
nor U10430 (N_10430,N_10128,N_10199);
or U10431 (N_10431,N_10062,N_10008);
and U10432 (N_10432,N_10234,N_10010);
and U10433 (N_10433,N_10022,N_10010);
and U10434 (N_10434,N_10122,N_10197);
xnor U10435 (N_10435,N_10177,N_10057);
xnor U10436 (N_10436,N_10130,N_10002);
xor U10437 (N_10437,N_10091,N_10155);
xnor U10438 (N_10438,N_10234,N_10079);
xor U10439 (N_10439,N_10000,N_10053);
nand U10440 (N_10440,N_10222,N_10160);
xnor U10441 (N_10441,N_10063,N_10203);
or U10442 (N_10442,N_10049,N_10160);
nor U10443 (N_10443,N_10092,N_10004);
nand U10444 (N_10444,N_10050,N_10224);
xor U10445 (N_10445,N_10070,N_10181);
nor U10446 (N_10446,N_10174,N_10078);
xnor U10447 (N_10447,N_10173,N_10100);
xnor U10448 (N_10448,N_10243,N_10125);
or U10449 (N_10449,N_10005,N_10035);
or U10450 (N_10450,N_10020,N_10028);
nand U10451 (N_10451,N_10081,N_10121);
nor U10452 (N_10452,N_10177,N_10058);
and U10453 (N_10453,N_10048,N_10142);
nor U10454 (N_10454,N_10175,N_10000);
xnor U10455 (N_10455,N_10196,N_10004);
xor U10456 (N_10456,N_10126,N_10202);
or U10457 (N_10457,N_10096,N_10046);
xor U10458 (N_10458,N_10124,N_10131);
xnor U10459 (N_10459,N_10101,N_10236);
nor U10460 (N_10460,N_10025,N_10102);
and U10461 (N_10461,N_10046,N_10183);
and U10462 (N_10462,N_10078,N_10121);
and U10463 (N_10463,N_10178,N_10119);
nor U10464 (N_10464,N_10019,N_10057);
nor U10465 (N_10465,N_10082,N_10081);
nand U10466 (N_10466,N_10172,N_10080);
or U10467 (N_10467,N_10096,N_10025);
nand U10468 (N_10468,N_10124,N_10129);
nor U10469 (N_10469,N_10238,N_10093);
or U10470 (N_10470,N_10040,N_10005);
nand U10471 (N_10471,N_10228,N_10078);
or U10472 (N_10472,N_10224,N_10172);
and U10473 (N_10473,N_10158,N_10228);
xor U10474 (N_10474,N_10131,N_10070);
nor U10475 (N_10475,N_10044,N_10211);
and U10476 (N_10476,N_10006,N_10177);
and U10477 (N_10477,N_10103,N_10118);
or U10478 (N_10478,N_10118,N_10133);
or U10479 (N_10479,N_10169,N_10171);
nor U10480 (N_10480,N_10218,N_10206);
xnor U10481 (N_10481,N_10234,N_10084);
or U10482 (N_10482,N_10242,N_10018);
nand U10483 (N_10483,N_10050,N_10249);
nor U10484 (N_10484,N_10227,N_10211);
nor U10485 (N_10485,N_10168,N_10045);
nand U10486 (N_10486,N_10211,N_10106);
nand U10487 (N_10487,N_10149,N_10051);
xor U10488 (N_10488,N_10057,N_10225);
nor U10489 (N_10489,N_10182,N_10013);
or U10490 (N_10490,N_10076,N_10220);
and U10491 (N_10491,N_10034,N_10103);
or U10492 (N_10492,N_10173,N_10160);
xnor U10493 (N_10493,N_10200,N_10128);
or U10494 (N_10494,N_10162,N_10027);
xnor U10495 (N_10495,N_10054,N_10116);
nor U10496 (N_10496,N_10023,N_10142);
xnor U10497 (N_10497,N_10175,N_10195);
nand U10498 (N_10498,N_10014,N_10227);
or U10499 (N_10499,N_10128,N_10249);
xnor U10500 (N_10500,N_10353,N_10413);
nand U10501 (N_10501,N_10380,N_10439);
or U10502 (N_10502,N_10473,N_10316);
and U10503 (N_10503,N_10369,N_10376);
nor U10504 (N_10504,N_10362,N_10284);
nor U10505 (N_10505,N_10474,N_10400);
nor U10506 (N_10506,N_10270,N_10281);
or U10507 (N_10507,N_10414,N_10455);
nor U10508 (N_10508,N_10258,N_10336);
or U10509 (N_10509,N_10467,N_10348);
and U10510 (N_10510,N_10437,N_10373);
or U10511 (N_10511,N_10299,N_10429);
or U10512 (N_10512,N_10321,N_10485);
nand U10513 (N_10513,N_10290,N_10289);
nor U10514 (N_10514,N_10423,N_10344);
and U10515 (N_10515,N_10392,N_10463);
and U10516 (N_10516,N_10418,N_10411);
or U10517 (N_10517,N_10350,N_10441);
nor U10518 (N_10518,N_10261,N_10273);
xnor U10519 (N_10519,N_10499,N_10378);
and U10520 (N_10520,N_10438,N_10271);
nor U10521 (N_10521,N_10309,N_10372);
nand U10522 (N_10522,N_10297,N_10375);
or U10523 (N_10523,N_10282,N_10268);
and U10524 (N_10524,N_10476,N_10453);
xor U10525 (N_10525,N_10356,N_10374);
and U10526 (N_10526,N_10267,N_10492);
xor U10527 (N_10527,N_10409,N_10331);
or U10528 (N_10528,N_10365,N_10488);
xor U10529 (N_10529,N_10388,N_10421);
xor U10530 (N_10530,N_10448,N_10340);
nand U10531 (N_10531,N_10498,N_10406);
nor U10532 (N_10532,N_10456,N_10252);
and U10533 (N_10533,N_10457,N_10296);
nand U10534 (N_10534,N_10458,N_10315);
and U10535 (N_10535,N_10325,N_10276);
xnor U10536 (N_10536,N_10433,N_10481);
nor U10537 (N_10537,N_10338,N_10327);
or U10538 (N_10538,N_10322,N_10478);
nor U10539 (N_10539,N_10472,N_10415);
nor U10540 (N_10540,N_10295,N_10487);
and U10541 (N_10541,N_10263,N_10293);
nor U10542 (N_10542,N_10253,N_10494);
nand U10543 (N_10543,N_10401,N_10454);
nand U10544 (N_10544,N_10332,N_10496);
nor U10545 (N_10545,N_10442,N_10363);
nand U10546 (N_10546,N_10355,N_10425);
and U10547 (N_10547,N_10447,N_10434);
nand U10548 (N_10548,N_10286,N_10475);
xor U10549 (N_10549,N_10343,N_10279);
xnor U10550 (N_10550,N_10342,N_10287);
and U10551 (N_10551,N_10334,N_10254);
xnor U10552 (N_10552,N_10395,N_10339);
nor U10553 (N_10553,N_10495,N_10314);
or U10554 (N_10554,N_10484,N_10366);
and U10555 (N_10555,N_10398,N_10430);
or U10556 (N_10556,N_10391,N_10311);
nand U10557 (N_10557,N_10451,N_10403);
xor U10558 (N_10558,N_10352,N_10399);
nor U10559 (N_10559,N_10377,N_10435);
nand U10560 (N_10560,N_10305,N_10266);
or U10561 (N_10561,N_10346,N_10264);
nor U10562 (N_10562,N_10444,N_10449);
and U10563 (N_10563,N_10379,N_10464);
or U10564 (N_10564,N_10470,N_10445);
and U10565 (N_10565,N_10387,N_10324);
xor U10566 (N_10566,N_10318,N_10275);
and U10567 (N_10567,N_10294,N_10328);
xor U10568 (N_10568,N_10466,N_10477);
nand U10569 (N_10569,N_10420,N_10359);
or U10570 (N_10570,N_10490,N_10424);
or U10571 (N_10571,N_10381,N_10402);
nand U10572 (N_10572,N_10303,N_10250);
nor U10573 (N_10573,N_10436,N_10300);
nor U10574 (N_10574,N_10278,N_10256);
nand U10575 (N_10575,N_10446,N_10427);
nand U10576 (N_10576,N_10308,N_10357);
nand U10577 (N_10577,N_10419,N_10469);
nor U10578 (N_10578,N_10396,N_10404);
nor U10579 (N_10579,N_10277,N_10265);
or U10580 (N_10580,N_10341,N_10407);
and U10581 (N_10581,N_10260,N_10360);
or U10582 (N_10582,N_10259,N_10428);
nor U10583 (N_10583,N_10288,N_10384);
or U10584 (N_10584,N_10480,N_10390);
xnor U10585 (N_10585,N_10367,N_10383);
or U10586 (N_10586,N_10302,N_10426);
xnor U10587 (N_10587,N_10333,N_10479);
and U10588 (N_10588,N_10482,N_10405);
and U10589 (N_10589,N_10431,N_10298);
or U10590 (N_10590,N_10408,N_10301);
and U10591 (N_10591,N_10382,N_10274);
xor U10592 (N_10592,N_10262,N_10422);
and U10593 (N_10593,N_10307,N_10385);
or U10594 (N_10594,N_10329,N_10335);
and U10595 (N_10595,N_10417,N_10410);
nand U10596 (N_10596,N_10368,N_10459);
nor U10597 (N_10597,N_10292,N_10491);
nand U10598 (N_10598,N_10312,N_10371);
nand U10599 (N_10599,N_10291,N_10393);
xor U10600 (N_10600,N_10358,N_10330);
nand U10601 (N_10601,N_10323,N_10347);
or U10602 (N_10602,N_10460,N_10432);
nor U10603 (N_10603,N_10354,N_10255);
xor U10604 (N_10604,N_10416,N_10452);
nand U10605 (N_10605,N_10351,N_10280);
nor U10606 (N_10606,N_10306,N_10389);
xor U10607 (N_10607,N_10497,N_10394);
nor U10608 (N_10608,N_10361,N_10283);
xnor U10609 (N_10609,N_10304,N_10269);
xor U10610 (N_10610,N_10468,N_10310);
and U10611 (N_10611,N_10465,N_10251);
nor U10612 (N_10612,N_10493,N_10440);
and U10613 (N_10613,N_10285,N_10489);
nand U10614 (N_10614,N_10483,N_10257);
nand U10615 (N_10615,N_10471,N_10397);
nor U10616 (N_10616,N_10345,N_10337);
and U10617 (N_10617,N_10370,N_10462);
nor U10618 (N_10618,N_10450,N_10272);
and U10619 (N_10619,N_10461,N_10486);
or U10620 (N_10620,N_10386,N_10412);
nor U10621 (N_10621,N_10326,N_10320);
nor U10622 (N_10622,N_10349,N_10443);
nand U10623 (N_10623,N_10319,N_10364);
or U10624 (N_10624,N_10313,N_10317);
nor U10625 (N_10625,N_10423,N_10387);
and U10626 (N_10626,N_10414,N_10399);
and U10627 (N_10627,N_10472,N_10277);
xnor U10628 (N_10628,N_10473,N_10289);
or U10629 (N_10629,N_10492,N_10337);
and U10630 (N_10630,N_10305,N_10270);
xnor U10631 (N_10631,N_10485,N_10406);
or U10632 (N_10632,N_10362,N_10352);
nand U10633 (N_10633,N_10250,N_10392);
xor U10634 (N_10634,N_10401,N_10345);
and U10635 (N_10635,N_10330,N_10350);
or U10636 (N_10636,N_10287,N_10281);
and U10637 (N_10637,N_10343,N_10277);
or U10638 (N_10638,N_10477,N_10304);
xnor U10639 (N_10639,N_10405,N_10379);
and U10640 (N_10640,N_10393,N_10364);
nand U10641 (N_10641,N_10395,N_10487);
or U10642 (N_10642,N_10464,N_10370);
nor U10643 (N_10643,N_10496,N_10470);
or U10644 (N_10644,N_10297,N_10340);
or U10645 (N_10645,N_10388,N_10267);
or U10646 (N_10646,N_10477,N_10377);
nor U10647 (N_10647,N_10272,N_10267);
or U10648 (N_10648,N_10369,N_10499);
and U10649 (N_10649,N_10438,N_10349);
xnor U10650 (N_10650,N_10333,N_10442);
or U10651 (N_10651,N_10463,N_10400);
or U10652 (N_10652,N_10267,N_10293);
nor U10653 (N_10653,N_10461,N_10261);
or U10654 (N_10654,N_10375,N_10413);
and U10655 (N_10655,N_10442,N_10287);
or U10656 (N_10656,N_10321,N_10299);
xnor U10657 (N_10657,N_10427,N_10481);
nand U10658 (N_10658,N_10389,N_10441);
nand U10659 (N_10659,N_10371,N_10290);
nand U10660 (N_10660,N_10356,N_10266);
nor U10661 (N_10661,N_10418,N_10369);
nand U10662 (N_10662,N_10423,N_10268);
and U10663 (N_10663,N_10493,N_10478);
or U10664 (N_10664,N_10366,N_10380);
nand U10665 (N_10665,N_10465,N_10297);
xnor U10666 (N_10666,N_10391,N_10312);
xnor U10667 (N_10667,N_10321,N_10359);
nor U10668 (N_10668,N_10366,N_10264);
nand U10669 (N_10669,N_10344,N_10440);
or U10670 (N_10670,N_10307,N_10438);
or U10671 (N_10671,N_10450,N_10410);
xor U10672 (N_10672,N_10253,N_10348);
and U10673 (N_10673,N_10438,N_10435);
nor U10674 (N_10674,N_10314,N_10485);
xor U10675 (N_10675,N_10440,N_10473);
xor U10676 (N_10676,N_10345,N_10360);
nand U10677 (N_10677,N_10344,N_10329);
or U10678 (N_10678,N_10492,N_10437);
or U10679 (N_10679,N_10261,N_10265);
or U10680 (N_10680,N_10275,N_10498);
nor U10681 (N_10681,N_10351,N_10303);
or U10682 (N_10682,N_10304,N_10278);
or U10683 (N_10683,N_10452,N_10445);
or U10684 (N_10684,N_10463,N_10348);
xnor U10685 (N_10685,N_10495,N_10416);
nor U10686 (N_10686,N_10489,N_10476);
xnor U10687 (N_10687,N_10343,N_10300);
or U10688 (N_10688,N_10257,N_10468);
xnor U10689 (N_10689,N_10427,N_10321);
nor U10690 (N_10690,N_10477,N_10335);
and U10691 (N_10691,N_10457,N_10349);
nand U10692 (N_10692,N_10335,N_10297);
xnor U10693 (N_10693,N_10267,N_10324);
xnor U10694 (N_10694,N_10478,N_10458);
nand U10695 (N_10695,N_10319,N_10482);
nor U10696 (N_10696,N_10301,N_10286);
nand U10697 (N_10697,N_10424,N_10355);
nand U10698 (N_10698,N_10490,N_10464);
nand U10699 (N_10699,N_10449,N_10491);
xor U10700 (N_10700,N_10313,N_10432);
and U10701 (N_10701,N_10265,N_10320);
nor U10702 (N_10702,N_10396,N_10327);
nor U10703 (N_10703,N_10292,N_10396);
or U10704 (N_10704,N_10381,N_10385);
nand U10705 (N_10705,N_10423,N_10300);
nor U10706 (N_10706,N_10479,N_10411);
and U10707 (N_10707,N_10416,N_10264);
and U10708 (N_10708,N_10499,N_10385);
nand U10709 (N_10709,N_10450,N_10333);
nand U10710 (N_10710,N_10322,N_10251);
and U10711 (N_10711,N_10310,N_10295);
nor U10712 (N_10712,N_10436,N_10396);
xor U10713 (N_10713,N_10432,N_10384);
or U10714 (N_10714,N_10292,N_10451);
or U10715 (N_10715,N_10278,N_10344);
xnor U10716 (N_10716,N_10332,N_10457);
nor U10717 (N_10717,N_10471,N_10442);
and U10718 (N_10718,N_10287,N_10485);
nand U10719 (N_10719,N_10250,N_10406);
or U10720 (N_10720,N_10325,N_10412);
and U10721 (N_10721,N_10250,N_10285);
nor U10722 (N_10722,N_10299,N_10432);
xnor U10723 (N_10723,N_10473,N_10288);
nor U10724 (N_10724,N_10477,N_10268);
nand U10725 (N_10725,N_10338,N_10451);
nor U10726 (N_10726,N_10398,N_10284);
and U10727 (N_10727,N_10260,N_10430);
or U10728 (N_10728,N_10348,N_10476);
and U10729 (N_10729,N_10420,N_10397);
or U10730 (N_10730,N_10479,N_10287);
nand U10731 (N_10731,N_10254,N_10442);
xnor U10732 (N_10732,N_10451,N_10425);
nor U10733 (N_10733,N_10340,N_10386);
nor U10734 (N_10734,N_10356,N_10394);
xor U10735 (N_10735,N_10446,N_10434);
nand U10736 (N_10736,N_10357,N_10304);
and U10737 (N_10737,N_10294,N_10382);
and U10738 (N_10738,N_10309,N_10337);
nor U10739 (N_10739,N_10252,N_10288);
nand U10740 (N_10740,N_10481,N_10497);
nand U10741 (N_10741,N_10351,N_10498);
nand U10742 (N_10742,N_10308,N_10439);
and U10743 (N_10743,N_10409,N_10257);
nor U10744 (N_10744,N_10325,N_10292);
or U10745 (N_10745,N_10379,N_10429);
nand U10746 (N_10746,N_10333,N_10466);
and U10747 (N_10747,N_10277,N_10271);
or U10748 (N_10748,N_10468,N_10330);
and U10749 (N_10749,N_10388,N_10390);
nand U10750 (N_10750,N_10732,N_10539);
and U10751 (N_10751,N_10697,N_10660);
and U10752 (N_10752,N_10742,N_10556);
or U10753 (N_10753,N_10622,N_10701);
nand U10754 (N_10754,N_10598,N_10696);
or U10755 (N_10755,N_10553,N_10537);
nand U10756 (N_10756,N_10678,N_10748);
nor U10757 (N_10757,N_10724,N_10698);
or U10758 (N_10758,N_10649,N_10526);
and U10759 (N_10759,N_10636,N_10746);
nor U10760 (N_10760,N_10576,N_10740);
xnor U10761 (N_10761,N_10567,N_10568);
and U10762 (N_10762,N_10523,N_10578);
nand U10763 (N_10763,N_10703,N_10735);
nand U10764 (N_10764,N_10500,N_10546);
nor U10765 (N_10765,N_10533,N_10586);
and U10766 (N_10766,N_10626,N_10525);
and U10767 (N_10767,N_10672,N_10702);
and U10768 (N_10768,N_10670,N_10579);
or U10769 (N_10769,N_10723,N_10739);
nor U10770 (N_10770,N_10625,N_10656);
and U10771 (N_10771,N_10590,N_10587);
and U10772 (N_10772,N_10575,N_10544);
nor U10773 (N_10773,N_10518,N_10628);
nor U10774 (N_10774,N_10506,N_10617);
and U10775 (N_10775,N_10534,N_10507);
xnor U10776 (N_10776,N_10563,N_10595);
xnor U10777 (N_10777,N_10540,N_10619);
xnor U10778 (N_10778,N_10684,N_10704);
nand U10779 (N_10779,N_10705,N_10725);
nand U10780 (N_10780,N_10733,N_10527);
xnor U10781 (N_10781,N_10606,N_10535);
or U10782 (N_10782,N_10543,N_10646);
xor U10783 (N_10783,N_10550,N_10612);
or U10784 (N_10784,N_10727,N_10699);
nor U10785 (N_10785,N_10505,N_10736);
xor U10786 (N_10786,N_10630,N_10585);
and U10787 (N_10787,N_10747,N_10706);
and U10788 (N_10788,N_10712,N_10528);
nand U10789 (N_10789,N_10611,N_10669);
nor U10790 (N_10790,N_10682,N_10503);
nor U10791 (N_10791,N_10618,N_10597);
nand U10792 (N_10792,N_10613,N_10651);
nand U10793 (N_10793,N_10666,N_10547);
and U10794 (N_10794,N_10531,N_10570);
xor U10795 (N_10795,N_10592,N_10726);
nor U10796 (N_10796,N_10675,N_10560);
nand U10797 (N_10797,N_10709,N_10718);
nand U10798 (N_10798,N_10594,N_10596);
and U10799 (N_10799,N_10624,N_10645);
xnor U10800 (N_10800,N_10730,N_10708);
nor U10801 (N_10801,N_10734,N_10583);
or U10802 (N_10802,N_10639,N_10609);
nor U10803 (N_10803,N_10510,N_10520);
or U10804 (N_10804,N_10688,N_10504);
and U10805 (N_10805,N_10744,N_10693);
nor U10806 (N_10806,N_10635,N_10502);
nor U10807 (N_10807,N_10659,N_10582);
or U10808 (N_10808,N_10581,N_10519);
xor U10809 (N_10809,N_10572,N_10549);
nand U10810 (N_10810,N_10720,N_10593);
or U10811 (N_10811,N_10644,N_10642);
and U10812 (N_10812,N_10654,N_10513);
and U10813 (N_10813,N_10512,N_10623);
or U10814 (N_10814,N_10691,N_10667);
or U10815 (N_10815,N_10648,N_10640);
nor U10816 (N_10816,N_10721,N_10588);
or U10817 (N_10817,N_10524,N_10728);
nor U10818 (N_10818,N_10632,N_10552);
xnor U10819 (N_10819,N_10710,N_10653);
or U10820 (N_10820,N_10658,N_10616);
and U10821 (N_10821,N_10584,N_10621);
or U10822 (N_10822,N_10631,N_10650);
and U10823 (N_10823,N_10664,N_10738);
nand U10824 (N_10824,N_10610,N_10529);
and U10825 (N_10825,N_10605,N_10674);
xor U10826 (N_10826,N_10687,N_10603);
xnor U10827 (N_10827,N_10686,N_10555);
nand U10828 (N_10828,N_10677,N_10574);
and U10829 (N_10829,N_10511,N_10508);
xnor U10830 (N_10830,N_10569,N_10711);
or U10831 (N_10831,N_10509,N_10722);
and U10832 (N_10832,N_10741,N_10690);
nand U10833 (N_10833,N_10600,N_10634);
xnor U10834 (N_10834,N_10737,N_10561);
nand U10835 (N_10835,N_10538,N_10548);
nor U10836 (N_10836,N_10565,N_10679);
nand U10837 (N_10837,N_10638,N_10713);
nor U10838 (N_10838,N_10557,N_10662);
or U10839 (N_10839,N_10580,N_10577);
nand U10840 (N_10840,N_10559,N_10633);
xnor U10841 (N_10841,N_10608,N_10599);
or U10842 (N_10842,N_10637,N_10607);
nor U10843 (N_10843,N_10671,N_10573);
or U10844 (N_10844,N_10541,N_10652);
xor U10845 (N_10845,N_10685,N_10558);
nand U10846 (N_10846,N_10661,N_10663);
xnor U10847 (N_10847,N_10681,N_10521);
xor U10848 (N_10848,N_10647,N_10536);
xor U10849 (N_10849,N_10532,N_10657);
and U10850 (N_10850,N_10714,N_10695);
nand U10851 (N_10851,N_10501,N_10601);
nor U10852 (N_10852,N_10515,N_10668);
nor U10853 (N_10853,N_10719,N_10629);
or U10854 (N_10854,N_10715,N_10614);
nor U10855 (N_10855,N_10641,N_10514);
nor U10856 (N_10856,N_10676,N_10743);
nand U10857 (N_10857,N_10643,N_10680);
nor U10858 (N_10858,N_10731,N_10562);
xor U10859 (N_10859,N_10566,N_10694);
and U10860 (N_10860,N_10517,N_10545);
and U10861 (N_10861,N_10683,N_10530);
nor U10862 (N_10862,N_10516,N_10665);
xnor U10863 (N_10863,N_10542,N_10551);
or U10864 (N_10864,N_10716,N_10564);
or U10865 (N_10865,N_10591,N_10729);
xnor U10866 (N_10866,N_10627,N_10749);
nor U10867 (N_10867,N_10571,N_10655);
or U10868 (N_10868,N_10602,N_10707);
or U10869 (N_10869,N_10745,N_10673);
nand U10870 (N_10870,N_10589,N_10554);
and U10871 (N_10871,N_10717,N_10604);
and U10872 (N_10872,N_10700,N_10522);
or U10873 (N_10873,N_10615,N_10692);
and U10874 (N_10874,N_10689,N_10620);
and U10875 (N_10875,N_10674,N_10672);
xor U10876 (N_10876,N_10679,N_10656);
or U10877 (N_10877,N_10643,N_10675);
xor U10878 (N_10878,N_10618,N_10746);
nor U10879 (N_10879,N_10704,N_10508);
and U10880 (N_10880,N_10534,N_10509);
or U10881 (N_10881,N_10680,N_10590);
or U10882 (N_10882,N_10506,N_10615);
xnor U10883 (N_10883,N_10622,N_10673);
nand U10884 (N_10884,N_10733,N_10609);
and U10885 (N_10885,N_10741,N_10569);
nand U10886 (N_10886,N_10585,N_10621);
xor U10887 (N_10887,N_10698,N_10645);
nor U10888 (N_10888,N_10533,N_10747);
nor U10889 (N_10889,N_10728,N_10740);
xnor U10890 (N_10890,N_10635,N_10722);
nand U10891 (N_10891,N_10680,N_10690);
or U10892 (N_10892,N_10534,N_10654);
and U10893 (N_10893,N_10663,N_10679);
and U10894 (N_10894,N_10596,N_10560);
and U10895 (N_10895,N_10598,N_10652);
and U10896 (N_10896,N_10598,N_10713);
and U10897 (N_10897,N_10508,N_10741);
nor U10898 (N_10898,N_10695,N_10676);
nand U10899 (N_10899,N_10727,N_10743);
nor U10900 (N_10900,N_10644,N_10728);
nor U10901 (N_10901,N_10660,N_10691);
nor U10902 (N_10902,N_10591,N_10511);
xnor U10903 (N_10903,N_10649,N_10547);
and U10904 (N_10904,N_10536,N_10562);
or U10905 (N_10905,N_10501,N_10727);
nand U10906 (N_10906,N_10546,N_10670);
nand U10907 (N_10907,N_10560,N_10719);
xor U10908 (N_10908,N_10648,N_10702);
or U10909 (N_10909,N_10709,N_10510);
xnor U10910 (N_10910,N_10608,N_10555);
xnor U10911 (N_10911,N_10707,N_10726);
nand U10912 (N_10912,N_10681,N_10717);
or U10913 (N_10913,N_10631,N_10699);
nand U10914 (N_10914,N_10643,N_10540);
xnor U10915 (N_10915,N_10605,N_10714);
xor U10916 (N_10916,N_10626,N_10700);
or U10917 (N_10917,N_10589,N_10502);
xor U10918 (N_10918,N_10589,N_10696);
or U10919 (N_10919,N_10619,N_10620);
nor U10920 (N_10920,N_10593,N_10664);
xnor U10921 (N_10921,N_10622,N_10532);
xor U10922 (N_10922,N_10648,N_10531);
nor U10923 (N_10923,N_10733,N_10546);
nand U10924 (N_10924,N_10682,N_10711);
nor U10925 (N_10925,N_10715,N_10582);
nand U10926 (N_10926,N_10664,N_10655);
or U10927 (N_10927,N_10533,N_10689);
and U10928 (N_10928,N_10599,N_10568);
nand U10929 (N_10929,N_10686,N_10602);
nand U10930 (N_10930,N_10578,N_10508);
and U10931 (N_10931,N_10596,N_10670);
nand U10932 (N_10932,N_10641,N_10563);
xnor U10933 (N_10933,N_10667,N_10700);
nor U10934 (N_10934,N_10546,N_10620);
nand U10935 (N_10935,N_10578,N_10675);
and U10936 (N_10936,N_10608,N_10554);
nor U10937 (N_10937,N_10650,N_10664);
or U10938 (N_10938,N_10682,N_10690);
nand U10939 (N_10939,N_10691,N_10580);
or U10940 (N_10940,N_10635,N_10599);
xor U10941 (N_10941,N_10579,N_10516);
or U10942 (N_10942,N_10500,N_10672);
nand U10943 (N_10943,N_10707,N_10603);
xor U10944 (N_10944,N_10605,N_10737);
and U10945 (N_10945,N_10662,N_10711);
or U10946 (N_10946,N_10657,N_10643);
nand U10947 (N_10947,N_10722,N_10608);
and U10948 (N_10948,N_10567,N_10691);
nand U10949 (N_10949,N_10515,N_10565);
and U10950 (N_10950,N_10520,N_10599);
and U10951 (N_10951,N_10617,N_10611);
nand U10952 (N_10952,N_10587,N_10519);
and U10953 (N_10953,N_10657,N_10539);
nor U10954 (N_10954,N_10725,N_10603);
nor U10955 (N_10955,N_10642,N_10584);
nor U10956 (N_10956,N_10709,N_10740);
and U10957 (N_10957,N_10665,N_10676);
and U10958 (N_10958,N_10736,N_10683);
nand U10959 (N_10959,N_10581,N_10609);
xnor U10960 (N_10960,N_10563,N_10600);
and U10961 (N_10961,N_10503,N_10651);
xnor U10962 (N_10962,N_10712,N_10602);
xnor U10963 (N_10963,N_10706,N_10651);
nor U10964 (N_10964,N_10713,N_10654);
and U10965 (N_10965,N_10503,N_10596);
or U10966 (N_10966,N_10722,N_10627);
xor U10967 (N_10967,N_10542,N_10510);
nand U10968 (N_10968,N_10534,N_10603);
nor U10969 (N_10969,N_10636,N_10663);
or U10970 (N_10970,N_10506,N_10641);
or U10971 (N_10971,N_10524,N_10513);
nand U10972 (N_10972,N_10733,N_10577);
nor U10973 (N_10973,N_10520,N_10585);
xor U10974 (N_10974,N_10584,N_10617);
and U10975 (N_10975,N_10719,N_10590);
and U10976 (N_10976,N_10653,N_10725);
nand U10977 (N_10977,N_10549,N_10711);
nor U10978 (N_10978,N_10632,N_10589);
xor U10979 (N_10979,N_10565,N_10741);
nand U10980 (N_10980,N_10705,N_10575);
xnor U10981 (N_10981,N_10570,N_10556);
nor U10982 (N_10982,N_10601,N_10580);
nand U10983 (N_10983,N_10661,N_10562);
nor U10984 (N_10984,N_10569,N_10608);
or U10985 (N_10985,N_10587,N_10702);
and U10986 (N_10986,N_10698,N_10500);
xor U10987 (N_10987,N_10547,N_10655);
nand U10988 (N_10988,N_10583,N_10638);
and U10989 (N_10989,N_10666,N_10676);
xor U10990 (N_10990,N_10637,N_10719);
and U10991 (N_10991,N_10560,N_10545);
nor U10992 (N_10992,N_10598,N_10536);
and U10993 (N_10993,N_10725,N_10735);
nor U10994 (N_10994,N_10701,N_10659);
nor U10995 (N_10995,N_10623,N_10727);
nor U10996 (N_10996,N_10672,N_10677);
nor U10997 (N_10997,N_10713,N_10608);
and U10998 (N_10998,N_10564,N_10669);
or U10999 (N_10999,N_10683,N_10568);
nor U11000 (N_11000,N_10802,N_10811);
nor U11001 (N_11001,N_10944,N_10760);
nor U11002 (N_11002,N_10959,N_10865);
nor U11003 (N_11003,N_10953,N_10925);
and U11004 (N_11004,N_10861,N_10785);
or U11005 (N_11005,N_10869,N_10875);
and U11006 (N_11006,N_10934,N_10879);
and U11007 (N_11007,N_10906,N_10967);
and U11008 (N_11008,N_10890,N_10895);
nand U11009 (N_11009,N_10850,N_10857);
or U11010 (N_11010,N_10844,N_10926);
nor U11011 (N_11011,N_10988,N_10939);
xnor U11012 (N_11012,N_10966,N_10845);
nor U11013 (N_11013,N_10784,N_10770);
and U11014 (N_11014,N_10955,N_10825);
nand U11015 (N_11015,N_10989,N_10794);
and U11016 (N_11016,N_10913,N_10927);
and U11017 (N_11017,N_10853,N_10956);
nor U11018 (N_11018,N_10804,N_10924);
nor U11019 (N_11019,N_10991,N_10851);
nand U11020 (N_11020,N_10821,N_10759);
and U11021 (N_11021,N_10948,N_10874);
nor U11022 (N_11022,N_10904,N_10848);
nor U11023 (N_11023,N_10867,N_10807);
or U11024 (N_11024,N_10993,N_10949);
and U11025 (N_11025,N_10951,N_10887);
or U11026 (N_11026,N_10883,N_10805);
or U11027 (N_11027,N_10781,N_10872);
and U11028 (N_11028,N_10981,N_10986);
or U11029 (N_11029,N_10864,N_10787);
or U11030 (N_11030,N_10958,N_10833);
nor U11031 (N_11031,N_10756,N_10928);
nor U11032 (N_11032,N_10982,N_10909);
nand U11033 (N_11033,N_10894,N_10929);
nor U11034 (N_11034,N_10970,N_10751);
nand U11035 (N_11035,N_10810,N_10996);
xnor U11036 (N_11036,N_10942,N_10808);
or U11037 (N_11037,N_10963,N_10830);
or U11038 (N_11038,N_10754,N_10915);
nand U11039 (N_11039,N_10892,N_10941);
nand U11040 (N_11040,N_10968,N_10778);
and U11041 (N_11041,N_10871,N_10773);
nor U11042 (N_11042,N_10774,N_10987);
xnor U11043 (N_11043,N_10791,N_10900);
or U11044 (N_11044,N_10873,N_10856);
or U11045 (N_11045,N_10801,N_10828);
and U11046 (N_11046,N_10772,N_10999);
xnor U11047 (N_11047,N_10782,N_10814);
and U11048 (N_11048,N_10923,N_10995);
and U11049 (N_11049,N_10973,N_10972);
nand U11050 (N_11050,N_10876,N_10832);
nand U11051 (N_11051,N_10975,N_10868);
and U11052 (N_11052,N_10863,N_10943);
xor U11053 (N_11053,N_10893,N_10750);
and U11054 (N_11054,N_10891,N_10885);
and U11055 (N_11055,N_10767,N_10919);
and U11056 (N_11056,N_10837,N_10954);
or U11057 (N_11057,N_10945,N_10843);
nor U11058 (N_11058,N_10809,N_10799);
xor U11059 (N_11059,N_10888,N_10783);
nor U11060 (N_11060,N_10903,N_10870);
xor U11061 (N_11061,N_10858,N_10979);
or U11062 (N_11062,N_10940,N_10839);
nor U11063 (N_11063,N_10902,N_10788);
xor U11064 (N_11064,N_10947,N_10997);
and U11065 (N_11065,N_10884,N_10914);
xor U11066 (N_11066,N_10806,N_10898);
nand U11067 (N_11067,N_10950,N_10921);
and U11068 (N_11068,N_10961,N_10765);
and U11069 (N_11069,N_10769,N_10836);
nor U11070 (N_11070,N_10916,N_10881);
xnor U11071 (N_11071,N_10755,N_10918);
nor U11072 (N_11072,N_10860,N_10930);
xnor U11073 (N_11073,N_10786,N_10766);
or U11074 (N_11074,N_10964,N_10820);
or U11075 (N_11075,N_10812,N_10790);
and U11076 (N_11076,N_10795,N_10803);
nor U11077 (N_11077,N_10937,N_10777);
nand U11078 (N_11078,N_10912,N_10908);
nand U11079 (N_11079,N_10880,N_10822);
xnor U11080 (N_11080,N_10849,N_10905);
xnor U11081 (N_11081,N_10776,N_10907);
nor U11082 (N_11082,N_10882,N_10840);
or U11083 (N_11083,N_10932,N_10969);
nand U11084 (N_11084,N_10962,N_10771);
and U11085 (N_11085,N_10957,N_10976);
or U11086 (N_11086,N_10838,N_10800);
nor U11087 (N_11087,N_10946,N_10978);
nand U11088 (N_11088,N_10757,N_10817);
and U11089 (N_11089,N_10753,N_10977);
xor U11090 (N_11090,N_10789,N_10819);
nand U11091 (N_11091,N_10813,N_10971);
and U11092 (N_11092,N_10911,N_10931);
nand U11093 (N_11093,N_10793,N_10775);
nor U11094 (N_11094,N_10846,N_10960);
or U11095 (N_11095,N_10752,N_10829);
xor U11096 (N_11096,N_10965,N_10998);
xnor U11097 (N_11097,N_10854,N_10889);
nor U11098 (N_11098,N_10761,N_10936);
and U11099 (N_11099,N_10792,N_10763);
or U11100 (N_11100,N_10797,N_10935);
nand U11101 (N_11101,N_10985,N_10901);
xor U11102 (N_11102,N_10980,N_10922);
or U11103 (N_11103,N_10859,N_10827);
xor U11104 (N_11104,N_10780,N_10762);
and U11105 (N_11105,N_10933,N_10816);
nor U11106 (N_11106,N_10798,N_10834);
nand U11107 (N_11107,N_10992,N_10938);
nor U11108 (N_11108,N_10835,N_10796);
nor U11109 (N_11109,N_10764,N_10899);
nand U11110 (N_11110,N_10910,N_10952);
nor U11111 (N_11111,N_10920,N_10862);
and U11112 (N_11112,N_10815,N_10994);
and U11113 (N_11113,N_10855,N_10877);
nand U11114 (N_11114,N_10974,N_10878);
and U11115 (N_11115,N_10841,N_10896);
nand U11116 (N_11116,N_10847,N_10897);
and U11117 (N_11117,N_10831,N_10818);
or U11118 (N_11118,N_10990,N_10824);
and U11119 (N_11119,N_10842,N_10823);
and U11120 (N_11120,N_10983,N_10866);
nor U11121 (N_11121,N_10779,N_10758);
and U11122 (N_11122,N_10886,N_10984);
xor U11123 (N_11123,N_10768,N_10826);
or U11124 (N_11124,N_10917,N_10852);
and U11125 (N_11125,N_10911,N_10912);
nor U11126 (N_11126,N_10758,N_10861);
xnor U11127 (N_11127,N_10771,N_10956);
nand U11128 (N_11128,N_10799,N_10953);
and U11129 (N_11129,N_10884,N_10782);
and U11130 (N_11130,N_10961,N_10795);
nor U11131 (N_11131,N_10860,N_10791);
or U11132 (N_11132,N_10789,N_10779);
xnor U11133 (N_11133,N_10781,N_10825);
xor U11134 (N_11134,N_10990,N_10788);
or U11135 (N_11135,N_10957,N_10809);
xnor U11136 (N_11136,N_10816,N_10868);
xnor U11137 (N_11137,N_10873,N_10870);
nand U11138 (N_11138,N_10778,N_10783);
and U11139 (N_11139,N_10834,N_10791);
nand U11140 (N_11140,N_10827,N_10785);
nor U11141 (N_11141,N_10785,N_10750);
nor U11142 (N_11142,N_10812,N_10915);
nand U11143 (N_11143,N_10848,N_10856);
xor U11144 (N_11144,N_10913,N_10798);
or U11145 (N_11145,N_10904,N_10783);
or U11146 (N_11146,N_10872,N_10804);
or U11147 (N_11147,N_10897,N_10893);
nor U11148 (N_11148,N_10834,N_10829);
and U11149 (N_11149,N_10871,N_10966);
or U11150 (N_11150,N_10841,N_10820);
or U11151 (N_11151,N_10812,N_10760);
and U11152 (N_11152,N_10865,N_10994);
nand U11153 (N_11153,N_10920,N_10778);
and U11154 (N_11154,N_10806,N_10765);
or U11155 (N_11155,N_10781,N_10839);
and U11156 (N_11156,N_10984,N_10865);
or U11157 (N_11157,N_10953,N_10875);
or U11158 (N_11158,N_10922,N_10861);
nor U11159 (N_11159,N_10789,N_10900);
xnor U11160 (N_11160,N_10810,N_10994);
nand U11161 (N_11161,N_10977,N_10969);
xnor U11162 (N_11162,N_10929,N_10872);
xor U11163 (N_11163,N_10934,N_10836);
nand U11164 (N_11164,N_10814,N_10755);
nor U11165 (N_11165,N_10848,N_10884);
and U11166 (N_11166,N_10797,N_10909);
and U11167 (N_11167,N_10992,N_10880);
or U11168 (N_11168,N_10753,N_10819);
nor U11169 (N_11169,N_10903,N_10969);
or U11170 (N_11170,N_10917,N_10760);
or U11171 (N_11171,N_10762,N_10798);
xnor U11172 (N_11172,N_10802,N_10997);
xor U11173 (N_11173,N_10759,N_10912);
nor U11174 (N_11174,N_10907,N_10843);
nor U11175 (N_11175,N_10899,N_10775);
nand U11176 (N_11176,N_10891,N_10799);
and U11177 (N_11177,N_10781,N_10942);
or U11178 (N_11178,N_10838,N_10766);
nand U11179 (N_11179,N_10947,N_10821);
nand U11180 (N_11180,N_10980,N_10954);
nor U11181 (N_11181,N_10762,N_10829);
and U11182 (N_11182,N_10771,N_10998);
xor U11183 (N_11183,N_10841,N_10799);
xor U11184 (N_11184,N_10830,N_10860);
nor U11185 (N_11185,N_10928,N_10806);
xnor U11186 (N_11186,N_10864,N_10824);
and U11187 (N_11187,N_10786,N_10991);
xor U11188 (N_11188,N_10988,N_10966);
nand U11189 (N_11189,N_10985,N_10950);
nor U11190 (N_11190,N_10817,N_10805);
nor U11191 (N_11191,N_10795,N_10919);
nor U11192 (N_11192,N_10978,N_10939);
xnor U11193 (N_11193,N_10794,N_10926);
and U11194 (N_11194,N_10907,N_10974);
nand U11195 (N_11195,N_10826,N_10947);
xnor U11196 (N_11196,N_10998,N_10981);
and U11197 (N_11197,N_10814,N_10929);
xnor U11198 (N_11198,N_10886,N_10972);
or U11199 (N_11199,N_10930,N_10915);
and U11200 (N_11200,N_10771,N_10809);
nor U11201 (N_11201,N_10800,N_10895);
and U11202 (N_11202,N_10789,N_10950);
xnor U11203 (N_11203,N_10884,N_10996);
nor U11204 (N_11204,N_10991,N_10815);
or U11205 (N_11205,N_10765,N_10927);
or U11206 (N_11206,N_10871,N_10908);
or U11207 (N_11207,N_10910,N_10848);
or U11208 (N_11208,N_10855,N_10830);
nand U11209 (N_11209,N_10923,N_10989);
and U11210 (N_11210,N_10903,N_10862);
and U11211 (N_11211,N_10773,N_10848);
and U11212 (N_11212,N_10863,N_10960);
and U11213 (N_11213,N_10795,N_10778);
nor U11214 (N_11214,N_10869,N_10985);
nand U11215 (N_11215,N_10875,N_10811);
nor U11216 (N_11216,N_10809,N_10901);
xnor U11217 (N_11217,N_10966,N_10929);
xor U11218 (N_11218,N_10852,N_10764);
or U11219 (N_11219,N_10859,N_10891);
nor U11220 (N_11220,N_10879,N_10925);
nor U11221 (N_11221,N_10959,N_10987);
and U11222 (N_11222,N_10755,N_10835);
nand U11223 (N_11223,N_10835,N_10941);
xor U11224 (N_11224,N_10982,N_10880);
nand U11225 (N_11225,N_10988,N_10931);
xor U11226 (N_11226,N_10908,N_10852);
xor U11227 (N_11227,N_10755,N_10834);
nor U11228 (N_11228,N_10912,N_10832);
xnor U11229 (N_11229,N_10778,N_10963);
nand U11230 (N_11230,N_10959,N_10856);
or U11231 (N_11231,N_10835,N_10759);
and U11232 (N_11232,N_10815,N_10987);
or U11233 (N_11233,N_10974,N_10775);
nand U11234 (N_11234,N_10781,N_10870);
or U11235 (N_11235,N_10880,N_10968);
xor U11236 (N_11236,N_10960,N_10923);
xor U11237 (N_11237,N_10892,N_10997);
xor U11238 (N_11238,N_10875,N_10862);
nor U11239 (N_11239,N_10810,N_10831);
xnor U11240 (N_11240,N_10824,N_10807);
nor U11241 (N_11241,N_10828,N_10820);
and U11242 (N_11242,N_10938,N_10776);
nand U11243 (N_11243,N_10829,N_10923);
nor U11244 (N_11244,N_10955,N_10839);
xor U11245 (N_11245,N_10916,N_10832);
and U11246 (N_11246,N_10906,N_10968);
and U11247 (N_11247,N_10757,N_10955);
xnor U11248 (N_11248,N_10937,N_10855);
or U11249 (N_11249,N_10979,N_10901);
nor U11250 (N_11250,N_11013,N_11218);
nor U11251 (N_11251,N_11019,N_11030);
xor U11252 (N_11252,N_11109,N_11118);
nand U11253 (N_11253,N_11003,N_11131);
and U11254 (N_11254,N_11159,N_11130);
xor U11255 (N_11255,N_11193,N_11084);
xnor U11256 (N_11256,N_11066,N_11001);
nor U11257 (N_11257,N_11047,N_11140);
xnor U11258 (N_11258,N_11008,N_11240);
nand U11259 (N_11259,N_11075,N_11201);
xnor U11260 (N_11260,N_11239,N_11242);
nand U11261 (N_11261,N_11198,N_11234);
and U11262 (N_11262,N_11028,N_11195);
xor U11263 (N_11263,N_11007,N_11196);
xnor U11264 (N_11264,N_11022,N_11093);
and U11265 (N_11265,N_11162,N_11054);
nor U11266 (N_11266,N_11231,N_11059);
and U11267 (N_11267,N_11112,N_11135);
and U11268 (N_11268,N_11205,N_11191);
nor U11269 (N_11269,N_11045,N_11023);
nor U11270 (N_11270,N_11098,N_11186);
nand U11271 (N_11271,N_11136,N_11236);
or U11272 (N_11272,N_11115,N_11128);
and U11273 (N_11273,N_11002,N_11061);
xor U11274 (N_11274,N_11202,N_11173);
and U11275 (N_11275,N_11033,N_11151);
nand U11276 (N_11276,N_11228,N_11249);
or U11277 (N_11277,N_11086,N_11143);
and U11278 (N_11278,N_11025,N_11104);
and U11279 (N_11279,N_11081,N_11089);
xnor U11280 (N_11280,N_11035,N_11248);
xor U11281 (N_11281,N_11020,N_11216);
and U11282 (N_11282,N_11048,N_11122);
and U11283 (N_11283,N_11042,N_11126);
nor U11284 (N_11284,N_11150,N_11102);
nand U11285 (N_11285,N_11206,N_11044);
nand U11286 (N_11286,N_11096,N_11145);
nand U11287 (N_11287,N_11217,N_11064);
xor U11288 (N_11288,N_11107,N_11114);
and U11289 (N_11289,N_11214,N_11091);
xor U11290 (N_11290,N_11247,N_11032);
xnor U11291 (N_11291,N_11055,N_11026);
nand U11292 (N_11292,N_11188,N_11027);
nor U11293 (N_11293,N_11060,N_11233);
nand U11294 (N_11294,N_11094,N_11199);
nor U11295 (N_11295,N_11180,N_11229);
and U11296 (N_11296,N_11110,N_11170);
nor U11297 (N_11297,N_11051,N_11220);
or U11298 (N_11298,N_11052,N_11245);
nor U11299 (N_11299,N_11176,N_11071);
nand U11300 (N_11300,N_11190,N_11015);
and U11301 (N_11301,N_11034,N_11031);
and U11302 (N_11302,N_11073,N_11204);
nor U11303 (N_11303,N_11085,N_11076);
and U11304 (N_11304,N_11213,N_11222);
nand U11305 (N_11305,N_11133,N_11123);
and U11306 (N_11306,N_11010,N_11155);
or U11307 (N_11307,N_11153,N_11164);
and U11308 (N_11308,N_11241,N_11215);
xnor U11309 (N_11309,N_11097,N_11018);
xnor U11310 (N_11310,N_11158,N_11132);
or U11311 (N_11311,N_11221,N_11014);
nand U11312 (N_11312,N_11046,N_11038);
nand U11313 (N_11313,N_11111,N_11141);
xor U11314 (N_11314,N_11121,N_11117);
nand U11315 (N_11315,N_11120,N_11012);
xnor U11316 (N_11316,N_11134,N_11223);
and U11317 (N_11317,N_11056,N_11004);
and U11318 (N_11318,N_11208,N_11088);
nand U11319 (N_11319,N_11040,N_11041);
nor U11320 (N_11320,N_11080,N_11039);
nor U11321 (N_11321,N_11192,N_11219);
nand U11322 (N_11322,N_11183,N_11050);
xnor U11323 (N_11323,N_11149,N_11172);
nor U11324 (N_11324,N_11138,N_11062);
nand U11325 (N_11325,N_11016,N_11057);
or U11326 (N_11326,N_11127,N_11144);
or U11327 (N_11327,N_11113,N_11244);
or U11328 (N_11328,N_11163,N_11137);
nand U11329 (N_11329,N_11232,N_11212);
and U11330 (N_11330,N_11237,N_11211);
and U11331 (N_11331,N_11129,N_11246);
nand U11332 (N_11332,N_11043,N_11203);
xnor U11333 (N_11333,N_11021,N_11147);
or U11334 (N_11334,N_11181,N_11227);
nor U11335 (N_11335,N_11171,N_11157);
nor U11336 (N_11336,N_11197,N_11074);
xor U11337 (N_11337,N_11029,N_11226);
nor U11338 (N_11338,N_11156,N_11177);
or U11339 (N_11339,N_11103,N_11166);
or U11340 (N_11340,N_11017,N_11024);
and U11341 (N_11341,N_11243,N_11182);
and U11342 (N_11342,N_11077,N_11179);
nand U11343 (N_11343,N_11070,N_11072);
or U11344 (N_11344,N_11011,N_11090);
or U11345 (N_11345,N_11189,N_11210);
and U11346 (N_11346,N_11125,N_11083);
or U11347 (N_11347,N_11063,N_11108);
xor U11348 (N_11348,N_11168,N_11207);
xnor U11349 (N_11349,N_11067,N_11225);
nor U11350 (N_11350,N_11142,N_11000);
xor U11351 (N_11351,N_11082,N_11146);
or U11352 (N_11352,N_11224,N_11100);
nor U11353 (N_11353,N_11095,N_11036);
or U11354 (N_11354,N_11184,N_11101);
nor U11355 (N_11355,N_11053,N_11194);
or U11356 (N_11356,N_11079,N_11209);
or U11357 (N_11357,N_11175,N_11235);
nor U11358 (N_11358,N_11005,N_11174);
and U11359 (N_11359,N_11119,N_11092);
nand U11360 (N_11360,N_11169,N_11152);
xor U11361 (N_11361,N_11105,N_11116);
or U11362 (N_11362,N_11087,N_11065);
nand U11363 (N_11363,N_11068,N_11148);
xnor U11364 (N_11364,N_11161,N_11230);
nor U11365 (N_11365,N_11099,N_11238);
or U11366 (N_11366,N_11069,N_11006);
and U11367 (N_11367,N_11167,N_11124);
nand U11368 (N_11368,N_11037,N_11009);
xor U11369 (N_11369,N_11154,N_11160);
or U11370 (N_11370,N_11187,N_11200);
nor U11371 (N_11371,N_11078,N_11049);
nand U11372 (N_11372,N_11165,N_11058);
nand U11373 (N_11373,N_11106,N_11178);
nand U11374 (N_11374,N_11185,N_11139);
xnor U11375 (N_11375,N_11194,N_11089);
xnor U11376 (N_11376,N_11178,N_11101);
xor U11377 (N_11377,N_11001,N_11122);
and U11378 (N_11378,N_11159,N_11157);
or U11379 (N_11379,N_11172,N_11093);
nor U11380 (N_11380,N_11180,N_11047);
and U11381 (N_11381,N_11132,N_11199);
nor U11382 (N_11382,N_11212,N_11135);
nand U11383 (N_11383,N_11231,N_11235);
or U11384 (N_11384,N_11091,N_11103);
or U11385 (N_11385,N_11143,N_11077);
nand U11386 (N_11386,N_11005,N_11028);
nor U11387 (N_11387,N_11116,N_11118);
or U11388 (N_11388,N_11001,N_11235);
or U11389 (N_11389,N_11219,N_11048);
nand U11390 (N_11390,N_11087,N_11086);
nand U11391 (N_11391,N_11172,N_11163);
xnor U11392 (N_11392,N_11197,N_11149);
nand U11393 (N_11393,N_11240,N_11034);
nor U11394 (N_11394,N_11019,N_11035);
nor U11395 (N_11395,N_11004,N_11245);
nand U11396 (N_11396,N_11175,N_11216);
or U11397 (N_11397,N_11167,N_11095);
or U11398 (N_11398,N_11034,N_11148);
xor U11399 (N_11399,N_11159,N_11132);
nor U11400 (N_11400,N_11135,N_11005);
and U11401 (N_11401,N_11242,N_11054);
xnor U11402 (N_11402,N_11210,N_11173);
xnor U11403 (N_11403,N_11153,N_11055);
or U11404 (N_11404,N_11162,N_11173);
and U11405 (N_11405,N_11241,N_11183);
nand U11406 (N_11406,N_11002,N_11213);
nor U11407 (N_11407,N_11207,N_11043);
xor U11408 (N_11408,N_11077,N_11025);
xnor U11409 (N_11409,N_11103,N_11133);
or U11410 (N_11410,N_11225,N_11195);
nor U11411 (N_11411,N_11041,N_11021);
or U11412 (N_11412,N_11201,N_11127);
nand U11413 (N_11413,N_11183,N_11073);
nand U11414 (N_11414,N_11215,N_11047);
or U11415 (N_11415,N_11047,N_11178);
nor U11416 (N_11416,N_11152,N_11180);
nand U11417 (N_11417,N_11146,N_11159);
and U11418 (N_11418,N_11032,N_11102);
or U11419 (N_11419,N_11180,N_11059);
and U11420 (N_11420,N_11206,N_11076);
and U11421 (N_11421,N_11158,N_11215);
nor U11422 (N_11422,N_11050,N_11157);
or U11423 (N_11423,N_11101,N_11135);
nand U11424 (N_11424,N_11051,N_11193);
xnor U11425 (N_11425,N_11044,N_11141);
nand U11426 (N_11426,N_11105,N_11012);
or U11427 (N_11427,N_11152,N_11112);
or U11428 (N_11428,N_11084,N_11227);
nand U11429 (N_11429,N_11202,N_11201);
xnor U11430 (N_11430,N_11208,N_11075);
or U11431 (N_11431,N_11133,N_11204);
and U11432 (N_11432,N_11138,N_11083);
xnor U11433 (N_11433,N_11190,N_11198);
nand U11434 (N_11434,N_11155,N_11016);
and U11435 (N_11435,N_11161,N_11001);
xor U11436 (N_11436,N_11079,N_11234);
nor U11437 (N_11437,N_11000,N_11029);
nand U11438 (N_11438,N_11097,N_11002);
or U11439 (N_11439,N_11000,N_11150);
xor U11440 (N_11440,N_11084,N_11210);
or U11441 (N_11441,N_11065,N_11179);
nand U11442 (N_11442,N_11012,N_11141);
nor U11443 (N_11443,N_11187,N_11155);
xnor U11444 (N_11444,N_11247,N_11200);
nand U11445 (N_11445,N_11083,N_11072);
xnor U11446 (N_11446,N_11053,N_11092);
or U11447 (N_11447,N_11045,N_11040);
nand U11448 (N_11448,N_11158,N_11195);
and U11449 (N_11449,N_11238,N_11087);
and U11450 (N_11450,N_11096,N_11066);
or U11451 (N_11451,N_11130,N_11076);
nor U11452 (N_11452,N_11205,N_11080);
or U11453 (N_11453,N_11041,N_11107);
and U11454 (N_11454,N_11164,N_11177);
nor U11455 (N_11455,N_11007,N_11006);
nand U11456 (N_11456,N_11215,N_11022);
nor U11457 (N_11457,N_11006,N_11151);
nand U11458 (N_11458,N_11241,N_11033);
nor U11459 (N_11459,N_11151,N_11236);
nor U11460 (N_11460,N_11184,N_11067);
and U11461 (N_11461,N_11030,N_11102);
nand U11462 (N_11462,N_11245,N_11143);
xnor U11463 (N_11463,N_11235,N_11193);
nand U11464 (N_11464,N_11244,N_11045);
and U11465 (N_11465,N_11011,N_11226);
nand U11466 (N_11466,N_11076,N_11249);
and U11467 (N_11467,N_11173,N_11205);
xor U11468 (N_11468,N_11047,N_11111);
xor U11469 (N_11469,N_11090,N_11002);
xor U11470 (N_11470,N_11006,N_11033);
nand U11471 (N_11471,N_11067,N_11020);
xor U11472 (N_11472,N_11232,N_11096);
xnor U11473 (N_11473,N_11075,N_11157);
xnor U11474 (N_11474,N_11179,N_11152);
nand U11475 (N_11475,N_11078,N_11067);
and U11476 (N_11476,N_11050,N_11111);
nor U11477 (N_11477,N_11108,N_11094);
nand U11478 (N_11478,N_11153,N_11068);
nand U11479 (N_11479,N_11128,N_11071);
or U11480 (N_11480,N_11069,N_11062);
nor U11481 (N_11481,N_11115,N_11151);
nor U11482 (N_11482,N_11003,N_11162);
and U11483 (N_11483,N_11161,N_11133);
and U11484 (N_11484,N_11134,N_11160);
nand U11485 (N_11485,N_11185,N_11083);
nand U11486 (N_11486,N_11116,N_11124);
nand U11487 (N_11487,N_11019,N_11139);
or U11488 (N_11488,N_11192,N_11118);
nor U11489 (N_11489,N_11169,N_11050);
nor U11490 (N_11490,N_11040,N_11197);
nor U11491 (N_11491,N_11193,N_11082);
or U11492 (N_11492,N_11125,N_11169);
nand U11493 (N_11493,N_11002,N_11029);
and U11494 (N_11494,N_11066,N_11019);
or U11495 (N_11495,N_11189,N_11219);
and U11496 (N_11496,N_11241,N_11063);
or U11497 (N_11497,N_11244,N_11091);
nand U11498 (N_11498,N_11041,N_11234);
xnor U11499 (N_11499,N_11101,N_11069);
and U11500 (N_11500,N_11485,N_11398);
nor U11501 (N_11501,N_11495,N_11352);
nand U11502 (N_11502,N_11256,N_11371);
and U11503 (N_11503,N_11311,N_11300);
nand U11504 (N_11504,N_11356,N_11444);
and U11505 (N_11505,N_11323,N_11291);
nand U11506 (N_11506,N_11309,N_11331);
nand U11507 (N_11507,N_11379,N_11457);
or U11508 (N_11508,N_11378,N_11325);
or U11509 (N_11509,N_11345,N_11433);
or U11510 (N_11510,N_11357,N_11429);
nand U11511 (N_11511,N_11389,N_11264);
nor U11512 (N_11512,N_11497,N_11287);
and U11513 (N_11513,N_11475,N_11401);
nor U11514 (N_11514,N_11326,N_11377);
nor U11515 (N_11515,N_11308,N_11299);
xor U11516 (N_11516,N_11259,N_11471);
nor U11517 (N_11517,N_11280,N_11418);
nor U11518 (N_11518,N_11448,N_11430);
and U11519 (N_11519,N_11346,N_11310);
xor U11520 (N_11520,N_11402,N_11406);
and U11521 (N_11521,N_11409,N_11404);
or U11522 (N_11522,N_11293,N_11286);
nor U11523 (N_11523,N_11373,N_11257);
and U11524 (N_11524,N_11327,N_11423);
nand U11525 (N_11525,N_11440,N_11476);
xnor U11526 (N_11526,N_11274,N_11255);
and U11527 (N_11527,N_11426,N_11496);
and U11528 (N_11528,N_11353,N_11302);
or U11529 (N_11529,N_11303,N_11278);
and U11530 (N_11530,N_11481,N_11499);
xor U11531 (N_11531,N_11470,N_11453);
nor U11532 (N_11532,N_11443,N_11321);
nand U11533 (N_11533,N_11474,N_11392);
nor U11534 (N_11534,N_11296,N_11416);
xnor U11535 (N_11535,N_11472,N_11432);
xor U11536 (N_11536,N_11307,N_11276);
nor U11537 (N_11537,N_11450,N_11253);
nand U11538 (N_11538,N_11313,N_11295);
xor U11539 (N_11539,N_11330,N_11337);
or U11540 (N_11540,N_11320,N_11268);
and U11541 (N_11541,N_11354,N_11284);
xor U11542 (N_11542,N_11410,N_11351);
nand U11543 (N_11543,N_11362,N_11387);
nor U11544 (N_11544,N_11266,N_11396);
nor U11545 (N_11545,N_11460,N_11380);
xnor U11546 (N_11546,N_11332,N_11348);
nor U11547 (N_11547,N_11455,N_11262);
xor U11548 (N_11548,N_11382,N_11458);
xor U11549 (N_11549,N_11322,N_11358);
and U11550 (N_11550,N_11366,N_11273);
xor U11551 (N_11551,N_11408,N_11361);
nor U11552 (N_11552,N_11384,N_11372);
and U11553 (N_11553,N_11400,N_11388);
or U11554 (N_11554,N_11427,N_11288);
and U11555 (N_11555,N_11316,N_11304);
nor U11556 (N_11556,N_11492,N_11317);
nor U11557 (N_11557,N_11431,N_11467);
nor U11558 (N_11558,N_11491,N_11441);
or U11559 (N_11559,N_11462,N_11424);
or U11560 (N_11560,N_11340,N_11258);
nand U11561 (N_11561,N_11281,N_11411);
and U11562 (N_11562,N_11261,N_11318);
or U11563 (N_11563,N_11428,N_11381);
nand U11564 (N_11564,N_11403,N_11370);
xor U11565 (N_11565,N_11263,N_11483);
xor U11566 (N_11566,N_11490,N_11477);
nand U11567 (N_11567,N_11333,N_11368);
nand U11568 (N_11568,N_11267,N_11363);
xor U11569 (N_11569,N_11315,N_11489);
and U11570 (N_11570,N_11463,N_11265);
nand U11571 (N_11571,N_11438,N_11487);
nand U11572 (N_11572,N_11367,N_11260);
nor U11573 (N_11573,N_11482,N_11461);
or U11574 (N_11574,N_11494,N_11399);
nand U11575 (N_11575,N_11415,N_11254);
and U11576 (N_11576,N_11334,N_11290);
nand U11577 (N_11577,N_11272,N_11386);
xor U11578 (N_11578,N_11336,N_11446);
xnor U11579 (N_11579,N_11269,N_11421);
nand U11580 (N_11580,N_11298,N_11279);
nor U11581 (N_11581,N_11270,N_11473);
or U11582 (N_11582,N_11312,N_11420);
nand U11583 (N_11583,N_11375,N_11349);
or U11584 (N_11584,N_11436,N_11412);
nand U11585 (N_11585,N_11397,N_11282);
and U11586 (N_11586,N_11391,N_11447);
nor U11587 (N_11587,N_11466,N_11435);
nand U11588 (N_11588,N_11271,N_11335);
or U11589 (N_11589,N_11297,N_11252);
xnor U11590 (N_11590,N_11341,N_11407);
xnor U11591 (N_11591,N_11289,N_11413);
or U11592 (N_11592,N_11451,N_11342);
nand U11593 (N_11593,N_11285,N_11479);
and U11594 (N_11594,N_11442,N_11301);
nor U11595 (N_11595,N_11484,N_11294);
nor U11596 (N_11596,N_11454,N_11394);
nand U11597 (N_11597,N_11464,N_11385);
nor U11598 (N_11598,N_11364,N_11344);
and U11599 (N_11599,N_11355,N_11324);
or U11600 (N_11600,N_11414,N_11306);
or U11601 (N_11601,N_11350,N_11437);
nand U11602 (N_11602,N_11376,N_11277);
and U11603 (N_11603,N_11347,N_11250);
and U11604 (N_11604,N_11393,N_11343);
nor U11605 (N_11605,N_11425,N_11417);
or U11606 (N_11606,N_11275,N_11405);
xnor U11607 (N_11607,N_11488,N_11422);
or U11608 (N_11608,N_11365,N_11339);
or U11609 (N_11609,N_11434,N_11456);
xnor U11610 (N_11610,N_11465,N_11390);
xor U11611 (N_11611,N_11283,N_11493);
or U11612 (N_11612,N_11329,N_11468);
and U11613 (N_11613,N_11338,N_11305);
nand U11614 (N_11614,N_11439,N_11449);
nand U11615 (N_11615,N_11459,N_11419);
xor U11616 (N_11616,N_11359,N_11369);
nor U11617 (N_11617,N_11452,N_11374);
nand U11618 (N_11618,N_11480,N_11319);
and U11619 (N_11619,N_11314,N_11498);
xnor U11620 (N_11620,N_11251,N_11360);
nand U11621 (N_11621,N_11395,N_11328);
nand U11622 (N_11622,N_11445,N_11292);
and U11623 (N_11623,N_11486,N_11478);
nor U11624 (N_11624,N_11383,N_11469);
and U11625 (N_11625,N_11411,N_11448);
or U11626 (N_11626,N_11329,N_11259);
xor U11627 (N_11627,N_11272,N_11359);
or U11628 (N_11628,N_11358,N_11259);
xnor U11629 (N_11629,N_11488,N_11379);
or U11630 (N_11630,N_11382,N_11338);
nand U11631 (N_11631,N_11273,N_11282);
and U11632 (N_11632,N_11345,N_11340);
nand U11633 (N_11633,N_11480,N_11253);
or U11634 (N_11634,N_11468,N_11295);
xnor U11635 (N_11635,N_11483,N_11470);
or U11636 (N_11636,N_11314,N_11252);
or U11637 (N_11637,N_11336,N_11409);
or U11638 (N_11638,N_11259,N_11391);
and U11639 (N_11639,N_11445,N_11279);
or U11640 (N_11640,N_11362,N_11421);
nor U11641 (N_11641,N_11486,N_11379);
nand U11642 (N_11642,N_11365,N_11480);
and U11643 (N_11643,N_11391,N_11303);
nand U11644 (N_11644,N_11459,N_11485);
xnor U11645 (N_11645,N_11429,N_11411);
xnor U11646 (N_11646,N_11421,N_11354);
or U11647 (N_11647,N_11329,N_11457);
or U11648 (N_11648,N_11330,N_11488);
nor U11649 (N_11649,N_11310,N_11441);
nand U11650 (N_11650,N_11296,N_11288);
nand U11651 (N_11651,N_11262,N_11436);
xnor U11652 (N_11652,N_11297,N_11344);
xor U11653 (N_11653,N_11293,N_11376);
xnor U11654 (N_11654,N_11258,N_11261);
and U11655 (N_11655,N_11318,N_11381);
or U11656 (N_11656,N_11421,N_11406);
nor U11657 (N_11657,N_11280,N_11482);
xor U11658 (N_11658,N_11281,N_11497);
nor U11659 (N_11659,N_11450,N_11438);
nor U11660 (N_11660,N_11338,N_11319);
nor U11661 (N_11661,N_11374,N_11379);
nor U11662 (N_11662,N_11321,N_11417);
nor U11663 (N_11663,N_11453,N_11491);
or U11664 (N_11664,N_11478,N_11298);
nor U11665 (N_11665,N_11259,N_11410);
xor U11666 (N_11666,N_11455,N_11470);
and U11667 (N_11667,N_11322,N_11338);
xor U11668 (N_11668,N_11424,N_11480);
or U11669 (N_11669,N_11345,N_11348);
xnor U11670 (N_11670,N_11386,N_11301);
nand U11671 (N_11671,N_11474,N_11357);
or U11672 (N_11672,N_11415,N_11317);
and U11673 (N_11673,N_11409,N_11388);
or U11674 (N_11674,N_11252,N_11260);
nand U11675 (N_11675,N_11321,N_11271);
and U11676 (N_11676,N_11473,N_11369);
or U11677 (N_11677,N_11434,N_11420);
xor U11678 (N_11678,N_11371,N_11384);
or U11679 (N_11679,N_11438,N_11425);
or U11680 (N_11680,N_11463,N_11415);
xnor U11681 (N_11681,N_11251,N_11488);
xnor U11682 (N_11682,N_11354,N_11385);
and U11683 (N_11683,N_11306,N_11420);
nand U11684 (N_11684,N_11339,N_11481);
and U11685 (N_11685,N_11408,N_11480);
nand U11686 (N_11686,N_11287,N_11289);
and U11687 (N_11687,N_11341,N_11396);
nand U11688 (N_11688,N_11405,N_11336);
or U11689 (N_11689,N_11413,N_11460);
xnor U11690 (N_11690,N_11431,N_11261);
nand U11691 (N_11691,N_11297,N_11370);
and U11692 (N_11692,N_11367,N_11253);
xor U11693 (N_11693,N_11315,N_11469);
xnor U11694 (N_11694,N_11307,N_11405);
or U11695 (N_11695,N_11407,N_11381);
and U11696 (N_11696,N_11460,N_11392);
or U11697 (N_11697,N_11331,N_11332);
nand U11698 (N_11698,N_11296,N_11323);
nand U11699 (N_11699,N_11276,N_11337);
xnor U11700 (N_11700,N_11397,N_11311);
nor U11701 (N_11701,N_11383,N_11437);
nand U11702 (N_11702,N_11463,N_11409);
nor U11703 (N_11703,N_11355,N_11480);
and U11704 (N_11704,N_11366,N_11483);
nor U11705 (N_11705,N_11328,N_11375);
xor U11706 (N_11706,N_11324,N_11291);
and U11707 (N_11707,N_11435,N_11337);
nand U11708 (N_11708,N_11400,N_11459);
or U11709 (N_11709,N_11328,N_11286);
nand U11710 (N_11710,N_11476,N_11379);
or U11711 (N_11711,N_11424,N_11256);
nand U11712 (N_11712,N_11338,N_11263);
nand U11713 (N_11713,N_11373,N_11250);
and U11714 (N_11714,N_11407,N_11393);
or U11715 (N_11715,N_11441,N_11396);
xor U11716 (N_11716,N_11390,N_11347);
nor U11717 (N_11717,N_11399,N_11335);
xnor U11718 (N_11718,N_11261,N_11453);
nor U11719 (N_11719,N_11368,N_11315);
or U11720 (N_11720,N_11420,N_11282);
or U11721 (N_11721,N_11273,N_11365);
xor U11722 (N_11722,N_11287,N_11252);
nor U11723 (N_11723,N_11304,N_11454);
or U11724 (N_11724,N_11402,N_11264);
xnor U11725 (N_11725,N_11331,N_11374);
nor U11726 (N_11726,N_11450,N_11339);
xnor U11727 (N_11727,N_11492,N_11257);
nor U11728 (N_11728,N_11382,N_11287);
nand U11729 (N_11729,N_11450,N_11269);
and U11730 (N_11730,N_11266,N_11331);
or U11731 (N_11731,N_11488,N_11407);
or U11732 (N_11732,N_11372,N_11374);
nand U11733 (N_11733,N_11311,N_11490);
xor U11734 (N_11734,N_11358,N_11337);
xnor U11735 (N_11735,N_11463,N_11313);
xnor U11736 (N_11736,N_11355,N_11395);
or U11737 (N_11737,N_11262,N_11461);
nand U11738 (N_11738,N_11313,N_11256);
nor U11739 (N_11739,N_11338,N_11422);
or U11740 (N_11740,N_11346,N_11317);
or U11741 (N_11741,N_11286,N_11499);
and U11742 (N_11742,N_11428,N_11329);
and U11743 (N_11743,N_11364,N_11482);
and U11744 (N_11744,N_11349,N_11266);
or U11745 (N_11745,N_11381,N_11304);
xnor U11746 (N_11746,N_11335,N_11421);
nand U11747 (N_11747,N_11480,N_11277);
or U11748 (N_11748,N_11353,N_11358);
or U11749 (N_11749,N_11365,N_11319);
and U11750 (N_11750,N_11526,N_11715);
or U11751 (N_11751,N_11663,N_11542);
xor U11752 (N_11752,N_11732,N_11712);
nand U11753 (N_11753,N_11703,N_11520);
xnor U11754 (N_11754,N_11672,N_11648);
xor U11755 (N_11755,N_11702,N_11619);
or U11756 (N_11756,N_11581,N_11639);
nor U11757 (N_11757,N_11711,N_11691);
and U11758 (N_11758,N_11610,N_11667);
nand U11759 (N_11759,N_11530,N_11737);
xnor U11760 (N_11760,N_11660,N_11503);
or U11761 (N_11761,N_11586,N_11652);
xnor U11762 (N_11762,N_11541,N_11707);
or U11763 (N_11763,N_11690,N_11678);
xnor U11764 (N_11764,N_11749,N_11731);
and U11765 (N_11765,N_11537,N_11563);
xnor U11766 (N_11766,N_11558,N_11576);
or U11767 (N_11767,N_11545,N_11512);
and U11768 (N_11768,N_11714,N_11535);
or U11769 (N_11769,N_11739,N_11710);
xor U11770 (N_11770,N_11516,N_11655);
and U11771 (N_11771,N_11525,N_11741);
xor U11772 (N_11772,N_11510,N_11719);
and U11773 (N_11773,N_11736,N_11509);
or U11774 (N_11774,N_11676,N_11556);
nor U11775 (N_11775,N_11500,N_11721);
or U11776 (N_11776,N_11649,N_11553);
and U11777 (N_11777,N_11653,N_11596);
nor U11778 (N_11778,N_11521,N_11677);
nor U11779 (N_11779,N_11573,N_11692);
and U11780 (N_11780,N_11585,N_11602);
xnor U11781 (N_11781,N_11594,N_11728);
or U11782 (N_11782,N_11668,N_11567);
and U11783 (N_11783,N_11633,N_11616);
nand U11784 (N_11784,N_11716,N_11701);
nor U11785 (N_11785,N_11515,N_11513);
and U11786 (N_11786,N_11607,N_11587);
nor U11787 (N_11787,N_11625,N_11745);
nor U11788 (N_11788,N_11675,N_11688);
nand U11789 (N_11789,N_11502,N_11704);
xnor U11790 (N_11790,N_11546,N_11566);
and U11791 (N_11791,N_11571,N_11599);
nor U11792 (N_11792,N_11523,N_11651);
nand U11793 (N_11793,N_11600,N_11726);
nor U11794 (N_11794,N_11624,N_11577);
or U11795 (N_11795,N_11729,N_11679);
nand U11796 (N_11796,N_11578,N_11614);
nand U11797 (N_11797,N_11575,N_11684);
nand U11798 (N_11798,N_11682,N_11548);
and U11799 (N_11799,N_11748,N_11713);
or U11800 (N_11800,N_11501,N_11557);
nand U11801 (N_11801,N_11685,N_11519);
xnor U11802 (N_11802,N_11611,N_11540);
nand U11803 (N_11803,N_11645,N_11559);
nand U11804 (N_11804,N_11696,N_11669);
xnor U11805 (N_11805,N_11555,N_11572);
and U11806 (N_11806,N_11640,N_11584);
nor U11807 (N_11807,N_11671,N_11593);
nor U11808 (N_11808,N_11699,N_11642);
or U11809 (N_11809,N_11720,N_11562);
and U11810 (N_11810,N_11533,N_11681);
nand U11811 (N_11811,N_11673,N_11643);
and U11812 (N_11812,N_11529,N_11524);
and U11813 (N_11813,N_11622,N_11536);
or U11814 (N_11814,N_11511,N_11595);
xor U11815 (N_11815,N_11606,N_11658);
xnor U11816 (N_11816,N_11644,N_11574);
nand U11817 (N_11817,N_11708,N_11592);
nor U11818 (N_11818,N_11664,N_11661);
or U11819 (N_11819,N_11733,N_11626);
nor U11820 (N_11820,N_11608,N_11544);
or U11821 (N_11821,N_11693,N_11665);
and U11822 (N_11822,N_11654,N_11734);
and U11823 (N_11823,N_11740,N_11638);
nand U11824 (N_11824,N_11507,N_11589);
and U11825 (N_11825,N_11518,N_11538);
xnor U11826 (N_11826,N_11659,N_11580);
xnor U11827 (N_11827,N_11723,N_11612);
nor U11828 (N_11828,N_11746,N_11632);
and U11829 (N_11829,N_11583,N_11522);
nor U11830 (N_11830,N_11547,N_11647);
nor U11831 (N_11831,N_11637,N_11700);
or U11832 (N_11832,N_11590,N_11550);
or U11833 (N_11833,N_11743,N_11694);
xnor U11834 (N_11834,N_11709,N_11695);
or U11835 (N_11835,N_11683,N_11514);
nor U11836 (N_11836,N_11698,N_11552);
or U11837 (N_11837,N_11598,N_11747);
or U11838 (N_11838,N_11569,N_11738);
or U11839 (N_11839,N_11724,N_11623);
or U11840 (N_11840,N_11551,N_11539);
xnor U11841 (N_11841,N_11722,N_11628);
nand U11842 (N_11842,N_11735,N_11657);
or U11843 (N_11843,N_11579,N_11630);
nand U11844 (N_11844,N_11670,N_11705);
nand U11845 (N_11845,N_11528,N_11725);
nor U11846 (N_11846,N_11527,N_11508);
and U11847 (N_11847,N_11609,N_11564);
or U11848 (N_11848,N_11727,N_11615);
and U11849 (N_11849,N_11531,N_11718);
and U11850 (N_11850,N_11656,N_11634);
nor U11851 (N_11851,N_11706,N_11565);
or U11852 (N_11852,N_11662,N_11568);
nor U11853 (N_11853,N_11635,N_11686);
nor U11854 (N_11854,N_11597,N_11601);
and U11855 (N_11855,N_11603,N_11582);
or U11856 (N_11856,N_11687,N_11605);
or U11857 (N_11857,N_11532,N_11591);
and U11858 (N_11858,N_11620,N_11641);
xnor U11859 (N_11859,N_11517,N_11561);
or U11860 (N_11860,N_11570,N_11621);
nor U11861 (N_11861,N_11627,N_11689);
and U11862 (N_11862,N_11646,N_11560);
or U11863 (N_11863,N_11742,N_11617);
xor U11864 (N_11864,N_11618,N_11534);
xnor U11865 (N_11865,N_11680,N_11613);
xor U11866 (N_11866,N_11674,N_11744);
and U11867 (N_11867,N_11549,N_11506);
nand U11868 (N_11868,N_11554,N_11650);
nand U11869 (N_11869,N_11631,N_11604);
nand U11870 (N_11870,N_11717,N_11588);
and U11871 (N_11871,N_11730,N_11666);
nor U11872 (N_11872,N_11543,N_11697);
nand U11873 (N_11873,N_11636,N_11629);
or U11874 (N_11874,N_11504,N_11505);
xor U11875 (N_11875,N_11567,N_11692);
or U11876 (N_11876,N_11571,N_11527);
nor U11877 (N_11877,N_11542,N_11569);
nand U11878 (N_11878,N_11503,N_11571);
or U11879 (N_11879,N_11703,N_11580);
nor U11880 (N_11880,N_11742,N_11653);
xor U11881 (N_11881,N_11564,N_11684);
nand U11882 (N_11882,N_11732,N_11588);
xor U11883 (N_11883,N_11721,N_11735);
and U11884 (N_11884,N_11528,N_11665);
nor U11885 (N_11885,N_11703,N_11730);
nand U11886 (N_11886,N_11675,N_11731);
or U11887 (N_11887,N_11595,N_11520);
and U11888 (N_11888,N_11577,N_11691);
nor U11889 (N_11889,N_11643,N_11746);
xor U11890 (N_11890,N_11742,N_11669);
nand U11891 (N_11891,N_11525,N_11701);
and U11892 (N_11892,N_11579,N_11595);
or U11893 (N_11893,N_11690,N_11680);
xnor U11894 (N_11894,N_11695,N_11587);
and U11895 (N_11895,N_11576,N_11660);
nand U11896 (N_11896,N_11589,N_11567);
nor U11897 (N_11897,N_11705,N_11542);
nor U11898 (N_11898,N_11661,N_11569);
nand U11899 (N_11899,N_11602,N_11598);
nand U11900 (N_11900,N_11512,N_11535);
nor U11901 (N_11901,N_11617,N_11655);
nand U11902 (N_11902,N_11516,N_11551);
and U11903 (N_11903,N_11743,N_11596);
nand U11904 (N_11904,N_11579,N_11745);
and U11905 (N_11905,N_11688,N_11611);
nand U11906 (N_11906,N_11646,N_11715);
or U11907 (N_11907,N_11595,N_11557);
nand U11908 (N_11908,N_11688,N_11731);
nand U11909 (N_11909,N_11740,N_11655);
and U11910 (N_11910,N_11713,N_11711);
xor U11911 (N_11911,N_11575,N_11666);
xnor U11912 (N_11912,N_11667,N_11647);
xor U11913 (N_11913,N_11697,N_11749);
and U11914 (N_11914,N_11689,N_11725);
nor U11915 (N_11915,N_11622,N_11631);
xor U11916 (N_11916,N_11638,N_11549);
xnor U11917 (N_11917,N_11561,N_11510);
or U11918 (N_11918,N_11640,N_11571);
xor U11919 (N_11919,N_11630,N_11687);
or U11920 (N_11920,N_11708,N_11555);
nor U11921 (N_11921,N_11560,N_11648);
or U11922 (N_11922,N_11729,N_11583);
and U11923 (N_11923,N_11583,N_11740);
nand U11924 (N_11924,N_11528,N_11536);
xnor U11925 (N_11925,N_11688,N_11698);
nor U11926 (N_11926,N_11737,N_11677);
and U11927 (N_11927,N_11600,N_11566);
nand U11928 (N_11928,N_11509,N_11676);
or U11929 (N_11929,N_11732,N_11674);
nor U11930 (N_11930,N_11635,N_11636);
and U11931 (N_11931,N_11567,N_11621);
and U11932 (N_11932,N_11692,N_11543);
xor U11933 (N_11933,N_11629,N_11734);
or U11934 (N_11934,N_11656,N_11516);
nor U11935 (N_11935,N_11694,N_11560);
and U11936 (N_11936,N_11724,N_11502);
xor U11937 (N_11937,N_11514,N_11602);
or U11938 (N_11938,N_11662,N_11676);
xnor U11939 (N_11939,N_11719,N_11636);
xnor U11940 (N_11940,N_11560,N_11735);
nand U11941 (N_11941,N_11527,N_11717);
xnor U11942 (N_11942,N_11621,N_11507);
nor U11943 (N_11943,N_11603,N_11699);
or U11944 (N_11944,N_11664,N_11741);
or U11945 (N_11945,N_11704,N_11597);
nor U11946 (N_11946,N_11553,N_11634);
nor U11947 (N_11947,N_11668,N_11613);
xor U11948 (N_11948,N_11583,N_11625);
nor U11949 (N_11949,N_11560,N_11691);
or U11950 (N_11950,N_11709,N_11604);
and U11951 (N_11951,N_11613,N_11505);
or U11952 (N_11952,N_11607,N_11501);
xor U11953 (N_11953,N_11687,N_11506);
xnor U11954 (N_11954,N_11588,N_11710);
xnor U11955 (N_11955,N_11617,N_11564);
xor U11956 (N_11956,N_11593,N_11659);
and U11957 (N_11957,N_11569,N_11562);
xnor U11958 (N_11958,N_11629,N_11550);
xnor U11959 (N_11959,N_11719,N_11523);
and U11960 (N_11960,N_11682,N_11538);
and U11961 (N_11961,N_11675,N_11597);
nor U11962 (N_11962,N_11573,N_11624);
or U11963 (N_11963,N_11572,N_11551);
and U11964 (N_11964,N_11686,N_11618);
or U11965 (N_11965,N_11546,N_11746);
nor U11966 (N_11966,N_11741,N_11562);
and U11967 (N_11967,N_11635,N_11564);
nand U11968 (N_11968,N_11600,N_11723);
or U11969 (N_11969,N_11664,N_11708);
or U11970 (N_11970,N_11700,N_11718);
nand U11971 (N_11971,N_11512,N_11665);
xor U11972 (N_11972,N_11516,N_11619);
nand U11973 (N_11973,N_11668,N_11558);
xnor U11974 (N_11974,N_11506,N_11587);
nor U11975 (N_11975,N_11515,N_11526);
nor U11976 (N_11976,N_11599,N_11738);
and U11977 (N_11977,N_11745,N_11696);
or U11978 (N_11978,N_11735,N_11701);
xnor U11979 (N_11979,N_11609,N_11518);
and U11980 (N_11980,N_11682,N_11566);
nand U11981 (N_11981,N_11735,N_11571);
nor U11982 (N_11982,N_11721,N_11590);
or U11983 (N_11983,N_11517,N_11737);
nand U11984 (N_11984,N_11686,N_11674);
and U11985 (N_11985,N_11712,N_11675);
and U11986 (N_11986,N_11732,N_11713);
or U11987 (N_11987,N_11748,N_11701);
nand U11988 (N_11988,N_11732,N_11660);
and U11989 (N_11989,N_11610,N_11524);
nor U11990 (N_11990,N_11706,N_11637);
nor U11991 (N_11991,N_11675,N_11600);
nand U11992 (N_11992,N_11698,N_11672);
nor U11993 (N_11993,N_11744,N_11723);
or U11994 (N_11994,N_11603,N_11658);
nor U11995 (N_11995,N_11749,N_11584);
xor U11996 (N_11996,N_11506,N_11545);
nand U11997 (N_11997,N_11581,N_11663);
nand U11998 (N_11998,N_11522,N_11591);
nand U11999 (N_11999,N_11718,N_11735);
and U12000 (N_12000,N_11806,N_11898);
or U12001 (N_12001,N_11942,N_11950);
nand U12002 (N_12002,N_11975,N_11818);
nor U12003 (N_12003,N_11982,N_11993);
or U12004 (N_12004,N_11903,N_11966);
nand U12005 (N_12005,N_11880,N_11754);
xnor U12006 (N_12006,N_11976,N_11838);
nor U12007 (N_12007,N_11855,N_11790);
and U12008 (N_12008,N_11949,N_11894);
xor U12009 (N_12009,N_11986,N_11809);
or U12010 (N_12010,N_11786,N_11829);
nand U12011 (N_12011,N_11781,N_11791);
or U12012 (N_12012,N_11863,N_11867);
xnor U12013 (N_12013,N_11803,N_11778);
nand U12014 (N_12014,N_11774,N_11890);
nor U12015 (N_12015,N_11813,N_11879);
nand U12016 (N_12016,N_11826,N_11914);
xor U12017 (N_12017,N_11875,N_11891);
nand U12018 (N_12018,N_11892,N_11797);
or U12019 (N_12019,N_11854,N_11977);
or U12020 (N_12020,N_11856,N_11761);
or U12021 (N_12021,N_11868,N_11938);
or U12022 (N_12022,N_11870,N_11864);
nor U12023 (N_12023,N_11817,N_11918);
xor U12024 (N_12024,N_11753,N_11767);
xor U12025 (N_12025,N_11971,N_11845);
nand U12026 (N_12026,N_11980,N_11897);
xnor U12027 (N_12027,N_11853,N_11835);
nand U12028 (N_12028,N_11902,N_11848);
and U12029 (N_12029,N_11936,N_11847);
xnor U12030 (N_12030,N_11978,N_11924);
xnor U12031 (N_12031,N_11758,N_11860);
xor U12032 (N_12032,N_11851,N_11805);
or U12033 (N_12033,N_11810,N_11849);
nor U12034 (N_12034,N_11766,N_11850);
nand U12035 (N_12035,N_11765,N_11959);
xnor U12036 (N_12036,N_11908,N_11955);
nor U12037 (N_12037,N_11901,N_11878);
xnor U12038 (N_12038,N_11907,N_11899);
and U12039 (N_12039,N_11906,N_11915);
or U12040 (N_12040,N_11904,N_11945);
nor U12041 (N_12041,N_11769,N_11931);
or U12042 (N_12042,N_11777,N_11815);
nor U12043 (N_12043,N_11954,N_11947);
and U12044 (N_12044,N_11872,N_11909);
or U12045 (N_12045,N_11820,N_11884);
and U12046 (N_12046,N_11926,N_11784);
nor U12047 (N_12047,N_11752,N_11923);
or U12048 (N_12048,N_11846,N_11999);
or U12049 (N_12049,N_11772,N_11830);
nand U12050 (N_12050,N_11920,N_11973);
nor U12051 (N_12051,N_11819,N_11824);
xor U12052 (N_12052,N_11943,N_11996);
xnor U12053 (N_12053,N_11771,N_11750);
xnor U12054 (N_12054,N_11808,N_11827);
or U12055 (N_12055,N_11921,N_11968);
xnor U12056 (N_12056,N_11958,N_11957);
nand U12057 (N_12057,N_11811,N_11912);
nand U12058 (N_12058,N_11930,N_11991);
nand U12059 (N_12059,N_11799,N_11967);
nand U12060 (N_12060,N_11961,N_11814);
xnor U12061 (N_12061,N_11944,N_11939);
nand U12062 (N_12062,N_11842,N_11756);
nand U12063 (N_12063,N_11989,N_11893);
xor U12064 (N_12064,N_11937,N_11965);
nand U12065 (N_12065,N_11916,N_11768);
nand U12066 (N_12066,N_11836,N_11773);
or U12067 (N_12067,N_11940,N_11877);
or U12068 (N_12068,N_11833,N_11964);
and U12069 (N_12069,N_11793,N_11828);
and U12070 (N_12070,N_11946,N_11816);
and U12071 (N_12071,N_11785,N_11922);
xor U12072 (N_12072,N_11843,N_11800);
and U12073 (N_12073,N_11974,N_11987);
nor U12074 (N_12074,N_11841,N_11876);
nand U12075 (N_12075,N_11783,N_11852);
and U12076 (N_12076,N_11956,N_11887);
xor U12077 (N_12077,N_11871,N_11911);
xnor U12078 (N_12078,N_11981,N_11757);
nand U12079 (N_12079,N_11927,N_11792);
or U12080 (N_12080,N_11821,N_11919);
or U12081 (N_12081,N_11928,N_11760);
and U12082 (N_12082,N_11992,N_11985);
or U12083 (N_12083,N_11776,N_11755);
nor U12084 (N_12084,N_11900,N_11859);
or U12085 (N_12085,N_11751,N_11801);
xor U12086 (N_12086,N_11831,N_11990);
xor U12087 (N_12087,N_11822,N_11881);
and U12088 (N_12088,N_11866,N_11759);
and U12089 (N_12089,N_11804,N_11888);
xor U12090 (N_12090,N_11840,N_11862);
nand U12091 (N_12091,N_11839,N_11934);
nand U12092 (N_12092,N_11969,N_11832);
xor U12093 (N_12093,N_11995,N_11935);
and U12094 (N_12094,N_11913,N_11948);
nand U12095 (N_12095,N_11960,N_11796);
or U12096 (N_12096,N_11886,N_11795);
xnor U12097 (N_12097,N_11798,N_11857);
and U12098 (N_12098,N_11910,N_11979);
nor U12099 (N_12099,N_11825,N_11789);
or U12100 (N_12100,N_11953,N_11764);
or U12101 (N_12101,N_11837,N_11963);
or U12102 (N_12102,N_11823,N_11874);
nor U12103 (N_12103,N_11997,N_11788);
nor U12104 (N_12104,N_11775,N_11763);
nand U12105 (N_12105,N_11873,N_11988);
or U12106 (N_12106,N_11896,N_11770);
and U12107 (N_12107,N_11962,N_11802);
or U12108 (N_12108,N_11858,N_11865);
nand U12109 (N_12109,N_11972,N_11998);
or U12110 (N_12110,N_11882,N_11869);
and U12111 (N_12111,N_11794,N_11807);
and U12112 (N_12112,N_11885,N_11812);
and U12113 (N_12113,N_11779,N_11970);
nand U12114 (N_12114,N_11994,N_11941);
nand U12115 (N_12115,N_11844,N_11983);
xnor U12116 (N_12116,N_11762,N_11984);
or U12117 (N_12117,N_11780,N_11883);
and U12118 (N_12118,N_11787,N_11895);
nor U12119 (N_12119,N_11905,N_11952);
nand U12120 (N_12120,N_11932,N_11861);
and U12121 (N_12121,N_11889,N_11951);
xor U12122 (N_12122,N_11929,N_11834);
nand U12123 (N_12123,N_11925,N_11782);
nor U12124 (N_12124,N_11917,N_11933);
nand U12125 (N_12125,N_11782,N_11995);
nand U12126 (N_12126,N_11836,N_11899);
and U12127 (N_12127,N_11920,N_11922);
xor U12128 (N_12128,N_11868,N_11876);
nand U12129 (N_12129,N_11915,N_11843);
or U12130 (N_12130,N_11842,N_11873);
and U12131 (N_12131,N_11992,N_11924);
nor U12132 (N_12132,N_11951,N_11799);
nand U12133 (N_12133,N_11800,N_11989);
nor U12134 (N_12134,N_11845,N_11766);
nor U12135 (N_12135,N_11914,N_11946);
xnor U12136 (N_12136,N_11916,N_11761);
or U12137 (N_12137,N_11870,N_11752);
or U12138 (N_12138,N_11846,N_11884);
and U12139 (N_12139,N_11837,N_11857);
nor U12140 (N_12140,N_11934,N_11845);
nand U12141 (N_12141,N_11923,N_11877);
or U12142 (N_12142,N_11939,N_11867);
nand U12143 (N_12143,N_11840,N_11958);
and U12144 (N_12144,N_11877,N_11936);
nand U12145 (N_12145,N_11971,N_11883);
nand U12146 (N_12146,N_11861,N_11838);
or U12147 (N_12147,N_11814,N_11934);
and U12148 (N_12148,N_11891,N_11779);
xnor U12149 (N_12149,N_11768,N_11900);
or U12150 (N_12150,N_11772,N_11799);
or U12151 (N_12151,N_11844,N_11895);
and U12152 (N_12152,N_11854,N_11964);
and U12153 (N_12153,N_11922,N_11843);
nand U12154 (N_12154,N_11959,N_11890);
or U12155 (N_12155,N_11952,N_11831);
or U12156 (N_12156,N_11846,N_11852);
and U12157 (N_12157,N_11819,N_11963);
xor U12158 (N_12158,N_11822,N_11782);
nand U12159 (N_12159,N_11983,N_11787);
and U12160 (N_12160,N_11761,N_11782);
nor U12161 (N_12161,N_11894,N_11966);
and U12162 (N_12162,N_11915,N_11848);
xnor U12163 (N_12163,N_11771,N_11861);
or U12164 (N_12164,N_11803,N_11831);
nand U12165 (N_12165,N_11935,N_11840);
xnor U12166 (N_12166,N_11782,N_11948);
and U12167 (N_12167,N_11996,N_11783);
nor U12168 (N_12168,N_11900,N_11788);
xor U12169 (N_12169,N_11926,N_11858);
nor U12170 (N_12170,N_11761,N_11925);
nor U12171 (N_12171,N_11991,N_11994);
nand U12172 (N_12172,N_11882,N_11818);
nand U12173 (N_12173,N_11783,N_11804);
nand U12174 (N_12174,N_11965,N_11779);
or U12175 (N_12175,N_11836,N_11880);
nand U12176 (N_12176,N_11775,N_11978);
and U12177 (N_12177,N_11990,N_11962);
xor U12178 (N_12178,N_11951,N_11781);
nand U12179 (N_12179,N_11954,N_11993);
xnor U12180 (N_12180,N_11910,N_11772);
nor U12181 (N_12181,N_11802,N_11755);
and U12182 (N_12182,N_11832,N_11906);
or U12183 (N_12183,N_11754,N_11750);
nand U12184 (N_12184,N_11825,N_11819);
and U12185 (N_12185,N_11818,N_11770);
and U12186 (N_12186,N_11985,N_11870);
nor U12187 (N_12187,N_11924,N_11866);
and U12188 (N_12188,N_11940,N_11929);
xnor U12189 (N_12189,N_11990,N_11754);
nand U12190 (N_12190,N_11894,N_11767);
nand U12191 (N_12191,N_11899,N_11970);
and U12192 (N_12192,N_11844,N_11925);
xnor U12193 (N_12193,N_11926,N_11984);
nand U12194 (N_12194,N_11899,N_11859);
nor U12195 (N_12195,N_11832,N_11885);
nand U12196 (N_12196,N_11940,N_11784);
nand U12197 (N_12197,N_11978,N_11897);
xor U12198 (N_12198,N_11879,N_11834);
nand U12199 (N_12199,N_11968,N_11913);
or U12200 (N_12200,N_11848,N_11850);
nand U12201 (N_12201,N_11800,N_11958);
nor U12202 (N_12202,N_11761,N_11792);
nor U12203 (N_12203,N_11804,N_11983);
nor U12204 (N_12204,N_11954,N_11751);
nand U12205 (N_12205,N_11931,N_11932);
or U12206 (N_12206,N_11874,N_11972);
and U12207 (N_12207,N_11867,N_11799);
nand U12208 (N_12208,N_11830,N_11804);
and U12209 (N_12209,N_11870,N_11917);
and U12210 (N_12210,N_11766,N_11750);
xnor U12211 (N_12211,N_11900,N_11784);
nand U12212 (N_12212,N_11996,N_11810);
nor U12213 (N_12213,N_11812,N_11905);
or U12214 (N_12214,N_11823,N_11827);
and U12215 (N_12215,N_11782,N_11911);
nand U12216 (N_12216,N_11901,N_11922);
and U12217 (N_12217,N_11840,N_11849);
nand U12218 (N_12218,N_11862,N_11922);
and U12219 (N_12219,N_11991,N_11948);
nand U12220 (N_12220,N_11817,N_11832);
or U12221 (N_12221,N_11898,N_11913);
nand U12222 (N_12222,N_11896,N_11833);
nand U12223 (N_12223,N_11871,N_11949);
or U12224 (N_12224,N_11874,N_11963);
nand U12225 (N_12225,N_11987,N_11889);
and U12226 (N_12226,N_11847,N_11960);
xnor U12227 (N_12227,N_11856,N_11798);
nand U12228 (N_12228,N_11986,N_11975);
and U12229 (N_12229,N_11885,N_11758);
nand U12230 (N_12230,N_11909,N_11930);
xor U12231 (N_12231,N_11999,N_11960);
or U12232 (N_12232,N_11846,N_11753);
or U12233 (N_12233,N_11902,N_11821);
nand U12234 (N_12234,N_11833,N_11762);
nor U12235 (N_12235,N_11800,N_11832);
nand U12236 (N_12236,N_11804,N_11753);
nand U12237 (N_12237,N_11893,N_11995);
nor U12238 (N_12238,N_11899,N_11935);
nand U12239 (N_12239,N_11855,N_11831);
and U12240 (N_12240,N_11914,N_11855);
or U12241 (N_12241,N_11821,N_11992);
and U12242 (N_12242,N_11759,N_11780);
nor U12243 (N_12243,N_11801,N_11971);
nor U12244 (N_12244,N_11758,N_11980);
and U12245 (N_12245,N_11750,N_11899);
and U12246 (N_12246,N_11849,N_11918);
xor U12247 (N_12247,N_11912,N_11783);
nand U12248 (N_12248,N_11971,N_11755);
nand U12249 (N_12249,N_11870,N_11976);
xnor U12250 (N_12250,N_12132,N_12085);
xnor U12251 (N_12251,N_12246,N_12107);
nand U12252 (N_12252,N_12176,N_12032);
xnor U12253 (N_12253,N_12030,N_12216);
or U12254 (N_12254,N_12009,N_12086);
nor U12255 (N_12255,N_12233,N_12073);
nor U12256 (N_12256,N_12114,N_12131);
and U12257 (N_12257,N_12024,N_12014);
or U12258 (N_12258,N_12047,N_12244);
nand U12259 (N_12259,N_12128,N_12170);
and U12260 (N_12260,N_12046,N_12089);
nor U12261 (N_12261,N_12044,N_12210);
nor U12262 (N_12262,N_12074,N_12197);
or U12263 (N_12263,N_12020,N_12237);
nand U12264 (N_12264,N_12016,N_12125);
and U12265 (N_12265,N_12177,N_12108);
or U12266 (N_12266,N_12178,N_12143);
nand U12267 (N_12267,N_12162,N_12069);
xnor U12268 (N_12268,N_12070,N_12241);
nor U12269 (N_12269,N_12208,N_12139);
and U12270 (N_12270,N_12027,N_12072);
and U12271 (N_12271,N_12117,N_12242);
xor U12272 (N_12272,N_12181,N_12213);
nor U12273 (N_12273,N_12167,N_12105);
xnor U12274 (N_12274,N_12059,N_12007);
or U12275 (N_12275,N_12054,N_12037);
nor U12276 (N_12276,N_12075,N_12211);
xnor U12277 (N_12277,N_12102,N_12051);
and U12278 (N_12278,N_12022,N_12110);
nor U12279 (N_12279,N_12228,N_12225);
xnor U12280 (N_12280,N_12091,N_12004);
xor U12281 (N_12281,N_12183,N_12062);
or U12282 (N_12282,N_12207,N_12238);
xor U12283 (N_12283,N_12104,N_12193);
and U12284 (N_12284,N_12093,N_12231);
xor U12285 (N_12285,N_12119,N_12101);
and U12286 (N_12286,N_12112,N_12088);
xnor U12287 (N_12287,N_12190,N_12226);
and U12288 (N_12288,N_12189,N_12191);
nor U12289 (N_12289,N_12099,N_12214);
nand U12290 (N_12290,N_12169,N_12063);
xor U12291 (N_12291,N_12227,N_12168);
nand U12292 (N_12292,N_12160,N_12036);
xor U12293 (N_12293,N_12081,N_12100);
nor U12294 (N_12294,N_12080,N_12221);
or U12295 (N_12295,N_12078,N_12017);
xor U12296 (N_12296,N_12234,N_12229);
nor U12297 (N_12297,N_12049,N_12068);
or U12298 (N_12298,N_12147,N_12205);
and U12299 (N_12299,N_12103,N_12011);
or U12300 (N_12300,N_12052,N_12135);
nor U12301 (N_12301,N_12155,N_12028);
nor U12302 (N_12302,N_12196,N_12240);
xor U12303 (N_12303,N_12094,N_12120);
xnor U12304 (N_12304,N_12133,N_12247);
or U12305 (N_12305,N_12066,N_12060);
nor U12306 (N_12306,N_12146,N_12179);
or U12307 (N_12307,N_12106,N_12209);
nor U12308 (N_12308,N_12087,N_12113);
nand U12309 (N_12309,N_12008,N_12029);
nor U12310 (N_12310,N_12023,N_12116);
and U12311 (N_12311,N_12111,N_12163);
and U12312 (N_12312,N_12067,N_12019);
nand U12313 (N_12313,N_12061,N_12172);
nand U12314 (N_12314,N_12137,N_12180);
nor U12315 (N_12315,N_12220,N_12026);
nor U12316 (N_12316,N_12230,N_12122);
xor U12317 (N_12317,N_12136,N_12015);
xnor U12318 (N_12318,N_12152,N_12200);
nor U12319 (N_12319,N_12035,N_12041);
and U12320 (N_12320,N_12006,N_12204);
nor U12321 (N_12321,N_12033,N_12175);
or U12322 (N_12322,N_12043,N_12159);
nor U12323 (N_12323,N_12127,N_12161);
xor U12324 (N_12324,N_12077,N_12144);
and U12325 (N_12325,N_12005,N_12050);
xor U12326 (N_12326,N_12215,N_12065);
nand U12327 (N_12327,N_12118,N_12224);
xnor U12328 (N_12328,N_12243,N_12218);
and U12329 (N_12329,N_12140,N_12000);
nor U12330 (N_12330,N_12239,N_12048);
nor U12331 (N_12331,N_12042,N_12186);
and U12332 (N_12332,N_12012,N_12192);
nand U12333 (N_12333,N_12153,N_12056);
nand U12334 (N_12334,N_12212,N_12222);
nand U12335 (N_12335,N_12090,N_12115);
nand U12336 (N_12336,N_12129,N_12002);
nor U12337 (N_12337,N_12217,N_12203);
nor U12338 (N_12338,N_12034,N_12154);
or U12339 (N_12339,N_12018,N_12223);
and U12340 (N_12340,N_12236,N_12039);
nor U12341 (N_12341,N_12188,N_12138);
xor U12342 (N_12342,N_12134,N_12201);
nand U12343 (N_12343,N_12092,N_12055);
nor U12344 (N_12344,N_12083,N_12064);
or U12345 (N_12345,N_12095,N_12053);
xnor U12346 (N_12346,N_12071,N_12151);
or U12347 (N_12347,N_12123,N_12057);
xor U12348 (N_12348,N_12149,N_12249);
or U12349 (N_12349,N_12079,N_12165);
or U12350 (N_12350,N_12098,N_12150);
nor U12351 (N_12351,N_12202,N_12038);
nor U12352 (N_12352,N_12130,N_12126);
and U12353 (N_12353,N_12187,N_12082);
nand U12354 (N_12354,N_12145,N_12158);
nor U12355 (N_12355,N_12198,N_12248);
xnor U12356 (N_12356,N_12021,N_12013);
and U12357 (N_12357,N_12010,N_12097);
xnor U12358 (N_12358,N_12185,N_12001);
or U12359 (N_12359,N_12148,N_12124);
or U12360 (N_12360,N_12040,N_12025);
xnor U12361 (N_12361,N_12173,N_12121);
nand U12362 (N_12362,N_12182,N_12171);
or U12363 (N_12363,N_12199,N_12194);
xor U12364 (N_12364,N_12003,N_12084);
nor U12365 (N_12365,N_12031,N_12235);
nor U12366 (N_12366,N_12045,N_12166);
nand U12367 (N_12367,N_12219,N_12157);
or U12368 (N_12368,N_12058,N_12096);
or U12369 (N_12369,N_12206,N_12141);
xnor U12370 (N_12370,N_12076,N_12156);
and U12371 (N_12371,N_12195,N_12109);
and U12372 (N_12372,N_12184,N_12232);
and U12373 (N_12373,N_12245,N_12164);
nor U12374 (N_12374,N_12142,N_12174);
and U12375 (N_12375,N_12229,N_12204);
or U12376 (N_12376,N_12037,N_12017);
and U12377 (N_12377,N_12095,N_12206);
xor U12378 (N_12378,N_12012,N_12092);
or U12379 (N_12379,N_12044,N_12199);
and U12380 (N_12380,N_12236,N_12128);
and U12381 (N_12381,N_12147,N_12098);
nor U12382 (N_12382,N_12149,N_12035);
nand U12383 (N_12383,N_12025,N_12217);
and U12384 (N_12384,N_12011,N_12115);
nand U12385 (N_12385,N_12184,N_12147);
xor U12386 (N_12386,N_12234,N_12154);
xor U12387 (N_12387,N_12247,N_12244);
nor U12388 (N_12388,N_12232,N_12013);
xor U12389 (N_12389,N_12077,N_12045);
nand U12390 (N_12390,N_12140,N_12059);
xnor U12391 (N_12391,N_12206,N_12192);
and U12392 (N_12392,N_12159,N_12183);
and U12393 (N_12393,N_12024,N_12138);
xor U12394 (N_12394,N_12032,N_12067);
or U12395 (N_12395,N_12000,N_12126);
xnor U12396 (N_12396,N_12241,N_12118);
and U12397 (N_12397,N_12234,N_12100);
xor U12398 (N_12398,N_12203,N_12004);
nand U12399 (N_12399,N_12184,N_12100);
and U12400 (N_12400,N_12098,N_12157);
xnor U12401 (N_12401,N_12096,N_12153);
or U12402 (N_12402,N_12017,N_12127);
nand U12403 (N_12403,N_12034,N_12204);
nor U12404 (N_12404,N_12137,N_12103);
xor U12405 (N_12405,N_12015,N_12024);
nor U12406 (N_12406,N_12190,N_12161);
and U12407 (N_12407,N_12237,N_12194);
nor U12408 (N_12408,N_12034,N_12107);
nor U12409 (N_12409,N_12153,N_12168);
and U12410 (N_12410,N_12152,N_12095);
nand U12411 (N_12411,N_12159,N_12112);
or U12412 (N_12412,N_12131,N_12133);
and U12413 (N_12413,N_12185,N_12182);
nand U12414 (N_12414,N_12087,N_12137);
and U12415 (N_12415,N_12113,N_12228);
xnor U12416 (N_12416,N_12127,N_12142);
xnor U12417 (N_12417,N_12034,N_12072);
nand U12418 (N_12418,N_12142,N_12007);
or U12419 (N_12419,N_12111,N_12041);
and U12420 (N_12420,N_12097,N_12202);
and U12421 (N_12421,N_12042,N_12034);
xor U12422 (N_12422,N_12072,N_12235);
nand U12423 (N_12423,N_12203,N_12087);
and U12424 (N_12424,N_12047,N_12087);
and U12425 (N_12425,N_12123,N_12071);
and U12426 (N_12426,N_12045,N_12191);
or U12427 (N_12427,N_12147,N_12198);
and U12428 (N_12428,N_12006,N_12109);
nand U12429 (N_12429,N_12183,N_12114);
xor U12430 (N_12430,N_12158,N_12012);
nor U12431 (N_12431,N_12116,N_12105);
xnor U12432 (N_12432,N_12215,N_12056);
or U12433 (N_12433,N_12008,N_12244);
xnor U12434 (N_12434,N_12150,N_12141);
or U12435 (N_12435,N_12172,N_12161);
nand U12436 (N_12436,N_12037,N_12025);
or U12437 (N_12437,N_12217,N_12059);
xnor U12438 (N_12438,N_12060,N_12092);
nor U12439 (N_12439,N_12066,N_12117);
nand U12440 (N_12440,N_12055,N_12087);
nand U12441 (N_12441,N_12177,N_12054);
nand U12442 (N_12442,N_12068,N_12203);
and U12443 (N_12443,N_12209,N_12195);
xnor U12444 (N_12444,N_12219,N_12118);
nor U12445 (N_12445,N_12180,N_12007);
or U12446 (N_12446,N_12015,N_12113);
nand U12447 (N_12447,N_12165,N_12020);
nand U12448 (N_12448,N_12148,N_12093);
nand U12449 (N_12449,N_12150,N_12116);
and U12450 (N_12450,N_12096,N_12165);
xnor U12451 (N_12451,N_12043,N_12137);
xnor U12452 (N_12452,N_12119,N_12023);
nor U12453 (N_12453,N_12008,N_12057);
nand U12454 (N_12454,N_12149,N_12116);
nand U12455 (N_12455,N_12142,N_12209);
xnor U12456 (N_12456,N_12077,N_12241);
nand U12457 (N_12457,N_12008,N_12101);
xnor U12458 (N_12458,N_12123,N_12078);
nand U12459 (N_12459,N_12163,N_12242);
nor U12460 (N_12460,N_12238,N_12113);
nor U12461 (N_12461,N_12142,N_12064);
and U12462 (N_12462,N_12107,N_12124);
and U12463 (N_12463,N_12228,N_12208);
or U12464 (N_12464,N_12103,N_12205);
xor U12465 (N_12465,N_12199,N_12018);
xor U12466 (N_12466,N_12120,N_12084);
xnor U12467 (N_12467,N_12036,N_12048);
nand U12468 (N_12468,N_12164,N_12181);
xor U12469 (N_12469,N_12018,N_12242);
and U12470 (N_12470,N_12086,N_12075);
nand U12471 (N_12471,N_12092,N_12066);
xnor U12472 (N_12472,N_12016,N_12149);
nor U12473 (N_12473,N_12081,N_12119);
xor U12474 (N_12474,N_12022,N_12001);
xnor U12475 (N_12475,N_12193,N_12094);
or U12476 (N_12476,N_12098,N_12054);
nor U12477 (N_12477,N_12157,N_12248);
and U12478 (N_12478,N_12205,N_12066);
or U12479 (N_12479,N_12081,N_12236);
xor U12480 (N_12480,N_12231,N_12212);
and U12481 (N_12481,N_12199,N_12050);
or U12482 (N_12482,N_12241,N_12027);
and U12483 (N_12483,N_12197,N_12162);
nor U12484 (N_12484,N_12132,N_12152);
or U12485 (N_12485,N_12241,N_12231);
xnor U12486 (N_12486,N_12030,N_12224);
xnor U12487 (N_12487,N_12042,N_12007);
or U12488 (N_12488,N_12044,N_12146);
and U12489 (N_12489,N_12238,N_12209);
xnor U12490 (N_12490,N_12146,N_12038);
and U12491 (N_12491,N_12120,N_12072);
nand U12492 (N_12492,N_12190,N_12069);
nand U12493 (N_12493,N_12164,N_12075);
nor U12494 (N_12494,N_12060,N_12078);
and U12495 (N_12495,N_12194,N_12066);
nand U12496 (N_12496,N_12182,N_12241);
nand U12497 (N_12497,N_12104,N_12217);
xnor U12498 (N_12498,N_12106,N_12225);
nor U12499 (N_12499,N_12136,N_12045);
or U12500 (N_12500,N_12361,N_12377);
nand U12501 (N_12501,N_12486,N_12442);
nand U12502 (N_12502,N_12408,N_12311);
or U12503 (N_12503,N_12402,N_12265);
xnor U12504 (N_12504,N_12288,N_12465);
and U12505 (N_12505,N_12464,N_12365);
nand U12506 (N_12506,N_12400,N_12478);
and U12507 (N_12507,N_12329,N_12429);
or U12508 (N_12508,N_12299,N_12324);
nor U12509 (N_12509,N_12315,N_12414);
nand U12510 (N_12510,N_12335,N_12273);
nor U12511 (N_12511,N_12373,N_12390);
or U12512 (N_12512,N_12268,N_12491);
nand U12513 (N_12513,N_12443,N_12428);
and U12514 (N_12514,N_12289,N_12317);
and U12515 (N_12515,N_12405,N_12308);
nor U12516 (N_12516,N_12480,N_12275);
nor U12517 (N_12517,N_12399,N_12497);
nor U12518 (N_12518,N_12459,N_12292);
nor U12519 (N_12519,N_12333,N_12492);
and U12520 (N_12520,N_12318,N_12267);
nand U12521 (N_12521,N_12363,N_12295);
xnor U12522 (N_12522,N_12391,N_12293);
xnor U12523 (N_12523,N_12355,N_12294);
xnor U12524 (N_12524,N_12291,N_12416);
nand U12525 (N_12525,N_12300,N_12372);
xnor U12526 (N_12526,N_12309,N_12407);
nor U12527 (N_12527,N_12276,N_12419);
nand U12528 (N_12528,N_12487,N_12353);
and U12529 (N_12529,N_12298,N_12446);
and U12530 (N_12530,N_12266,N_12452);
or U12531 (N_12531,N_12313,N_12250);
xnor U12532 (N_12532,N_12489,N_12339);
xor U12533 (N_12533,N_12471,N_12296);
nor U12534 (N_12534,N_12457,N_12332);
nand U12535 (N_12535,N_12322,N_12270);
or U12536 (N_12536,N_12398,N_12424);
or U12537 (N_12537,N_12279,N_12327);
nand U12538 (N_12538,N_12254,N_12302);
or U12539 (N_12539,N_12403,N_12352);
xor U12540 (N_12540,N_12432,N_12348);
xor U12541 (N_12541,N_12338,N_12297);
xnor U12542 (N_12542,N_12447,N_12427);
nor U12543 (N_12543,N_12436,N_12358);
nor U12544 (N_12544,N_12470,N_12351);
nand U12545 (N_12545,N_12259,N_12437);
nor U12546 (N_12546,N_12382,N_12421);
and U12547 (N_12547,N_12345,N_12380);
and U12548 (N_12548,N_12354,N_12422);
nand U12549 (N_12549,N_12425,N_12357);
nor U12550 (N_12550,N_12321,N_12462);
nand U12551 (N_12551,N_12325,N_12258);
nor U12552 (N_12552,N_12406,N_12385);
nand U12553 (N_12553,N_12269,N_12411);
nor U12554 (N_12554,N_12316,N_12434);
xnor U12555 (N_12555,N_12349,N_12320);
or U12556 (N_12556,N_12412,N_12448);
nand U12557 (N_12557,N_12444,N_12376);
nor U12558 (N_12558,N_12395,N_12496);
and U12559 (N_12559,N_12393,N_12346);
or U12560 (N_12560,N_12473,N_12342);
and U12561 (N_12561,N_12368,N_12445);
nand U12562 (N_12562,N_12262,N_12394);
nor U12563 (N_12563,N_12477,N_12344);
xor U12564 (N_12564,N_12413,N_12364);
nor U12565 (N_12565,N_12255,N_12341);
and U12566 (N_12566,N_12485,N_12435);
nor U12567 (N_12567,N_12326,N_12263);
and U12568 (N_12568,N_12453,N_12387);
or U12569 (N_12569,N_12347,N_12280);
nor U12570 (N_12570,N_12369,N_12306);
and U12571 (N_12571,N_12277,N_12483);
xor U12572 (N_12572,N_12493,N_12409);
xor U12573 (N_12573,N_12384,N_12456);
or U12574 (N_12574,N_12479,N_12467);
or U12575 (N_12575,N_12449,N_12334);
and U12576 (N_12576,N_12482,N_12397);
xor U12577 (N_12577,N_12307,N_12389);
xor U12578 (N_12578,N_12301,N_12451);
xor U12579 (N_12579,N_12433,N_12371);
nand U12580 (N_12580,N_12415,N_12439);
or U12581 (N_12581,N_12356,N_12495);
nand U12582 (N_12582,N_12460,N_12367);
nor U12583 (N_12583,N_12418,N_12392);
nand U12584 (N_12584,N_12466,N_12374);
nor U12585 (N_12585,N_12441,N_12383);
and U12586 (N_12586,N_12417,N_12274);
nand U12587 (N_12587,N_12252,N_12396);
or U12588 (N_12588,N_12350,N_12488);
or U12589 (N_12589,N_12378,N_12430);
and U12590 (N_12590,N_12458,N_12463);
or U12591 (N_12591,N_12314,N_12319);
nand U12592 (N_12592,N_12450,N_12271);
and U12593 (N_12593,N_12499,N_12257);
xor U12594 (N_12594,N_12474,N_12328);
nor U12595 (N_12595,N_12386,N_12330);
nor U12596 (N_12596,N_12423,N_12336);
or U12597 (N_12597,N_12476,N_12404);
nor U12598 (N_12598,N_12256,N_12469);
xnor U12599 (N_12599,N_12438,N_12251);
or U12600 (N_12600,N_12310,N_12331);
and U12601 (N_12601,N_12323,N_12484);
and U12602 (N_12602,N_12305,N_12303);
and U12603 (N_12603,N_12253,N_12472);
or U12604 (N_12604,N_12278,N_12401);
or U12605 (N_12605,N_12343,N_12284);
nand U12606 (N_12606,N_12312,N_12454);
or U12607 (N_12607,N_12286,N_12272);
nand U12608 (N_12608,N_12426,N_12283);
and U12609 (N_12609,N_12360,N_12379);
and U12610 (N_12610,N_12337,N_12304);
or U12611 (N_12611,N_12281,N_12264);
or U12612 (N_12612,N_12290,N_12481);
xor U12613 (N_12613,N_12440,N_12381);
xor U12614 (N_12614,N_12261,N_12260);
xor U12615 (N_12615,N_12468,N_12498);
xor U12616 (N_12616,N_12359,N_12287);
and U12617 (N_12617,N_12410,N_12475);
nand U12618 (N_12618,N_12455,N_12375);
nand U12619 (N_12619,N_12282,N_12370);
nand U12620 (N_12620,N_12366,N_12431);
and U12621 (N_12621,N_12490,N_12340);
or U12622 (N_12622,N_12494,N_12388);
nand U12623 (N_12623,N_12362,N_12285);
or U12624 (N_12624,N_12420,N_12461);
or U12625 (N_12625,N_12461,N_12257);
and U12626 (N_12626,N_12373,N_12292);
nor U12627 (N_12627,N_12326,N_12394);
nand U12628 (N_12628,N_12477,N_12315);
nor U12629 (N_12629,N_12287,N_12260);
xnor U12630 (N_12630,N_12465,N_12406);
and U12631 (N_12631,N_12265,N_12268);
nor U12632 (N_12632,N_12431,N_12284);
or U12633 (N_12633,N_12336,N_12346);
nand U12634 (N_12634,N_12454,N_12311);
and U12635 (N_12635,N_12308,N_12320);
nor U12636 (N_12636,N_12475,N_12403);
xor U12637 (N_12637,N_12331,N_12279);
or U12638 (N_12638,N_12320,N_12490);
nand U12639 (N_12639,N_12381,N_12443);
nand U12640 (N_12640,N_12419,N_12349);
xor U12641 (N_12641,N_12275,N_12330);
xor U12642 (N_12642,N_12253,N_12268);
and U12643 (N_12643,N_12424,N_12421);
xnor U12644 (N_12644,N_12348,N_12484);
nor U12645 (N_12645,N_12430,N_12396);
xnor U12646 (N_12646,N_12430,N_12465);
nor U12647 (N_12647,N_12334,N_12280);
or U12648 (N_12648,N_12419,N_12372);
or U12649 (N_12649,N_12345,N_12422);
nand U12650 (N_12650,N_12489,N_12360);
and U12651 (N_12651,N_12264,N_12401);
nor U12652 (N_12652,N_12422,N_12331);
nor U12653 (N_12653,N_12435,N_12448);
nor U12654 (N_12654,N_12287,N_12331);
xnor U12655 (N_12655,N_12309,N_12443);
nor U12656 (N_12656,N_12499,N_12437);
and U12657 (N_12657,N_12281,N_12377);
xor U12658 (N_12658,N_12379,N_12310);
and U12659 (N_12659,N_12255,N_12371);
or U12660 (N_12660,N_12301,N_12357);
or U12661 (N_12661,N_12308,N_12410);
or U12662 (N_12662,N_12421,N_12499);
nand U12663 (N_12663,N_12255,N_12450);
nor U12664 (N_12664,N_12322,N_12292);
or U12665 (N_12665,N_12314,N_12421);
nor U12666 (N_12666,N_12279,N_12485);
and U12667 (N_12667,N_12431,N_12375);
or U12668 (N_12668,N_12312,N_12499);
and U12669 (N_12669,N_12372,N_12457);
xnor U12670 (N_12670,N_12250,N_12459);
and U12671 (N_12671,N_12315,N_12494);
or U12672 (N_12672,N_12319,N_12434);
and U12673 (N_12673,N_12340,N_12368);
nand U12674 (N_12674,N_12260,N_12354);
and U12675 (N_12675,N_12312,N_12428);
and U12676 (N_12676,N_12492,N_12372);
nor U12677 (N_12677,N_12463,N_12411);
nor U12678 (N_12678,N_12424,N_12282);
or U12679 (N_12679,N_12348,N_12469);
xor U12680 (N_12680,N_12253,N_12373);
nor U12681 (N_12681,N_12362,N_12427);
xnor U12682 (N_12682,N_12404,N_12372);
and U12683 (N_12683,N_12374,N_12378);
or U12684 (N_12684,N_12348,N_12496);
xor U12685 (N_12685,N_12266,N_12401);
and U12686 (N_12686,N_12317,N_12327);
xnor U12687 (N_12687,N_12476,N_12458);
nand U12688 (N_12688,N_12264,N_12293);
xnor U12689 (N_12689,N_12322,N_12280);
or U12690 (N_12690,N_12273,N_12257);
xnor U12691 (N_12691,N_12306,N_12384);
or U12692 (N_12692,N_12308,N_12386);
nor U12693 (N_12693,N_12374,N_12433);
xor U12694 (N_12694,N_12488,N_12254);
nor U12695 (N_12695,N_12374,N_12298);
nor U12696 (N_12696,N_12272,N_12293);
and U12697 (N_12697,N_12338,N_12387);
nor U12698 (N_12698,N_12429,N_12420);
nor U12699 (N_12699,N_12353,N_12288);
xor U12700 (N_12700,N_12491,N_12298);
or U12701 (N_12701,N_12319,N_12386);
nor U12702 (N_12702,N_12417,N_12464);
nand U12703 (N_12703,N_12465,N_12267);
nand U12704 (N_12704,N_12372,N_12274);
nand U12705 (N_12705,N_12266,N_12297);
or U12706 (N_12706,N_12375,N_12463);
nand U12707 (N_12707,N_12371,N_12431);
and U12708 (N_12708,N_12361,N_12436);
or U12709 (N_12709,N_12396,N_12331);
and U12710 (N_12710,N_12493,N_12413);
xor U12711 (N_12711,N_12278,N_12276);
nor U12712 (N_12712,N_12430,N_12488);
or U12713 (N_12713,N_12454,N_12400);
and U12714 (N_12714,N_12255,N_12363);
and U12715 (N_12715,N_12280,N_12486);
nand U12716 (N_12716,N_12350,N_12258);
or U12717 (N_12717,N_12308,N_12302);
and U12718 (N_12718,N_12440,N_12277);
nor U12719 (N_12719,N_12283,N_12468);
xor U12720 (N_12720,N_12279,N_12398);
and U12721 (N_12721,N_12399,N_12480);
or U12722 (N_12722,N_12269,N_12308);
xor U12723 (N_12723,N_12367,N_12426);
and U12724 (N_12724,N_12323,N_12364);
and U12725 (N_12725,N_12400,N_12358);
xnor U12726 (N_12726,N_12416,N_12348);
nand U12727 (N_12727,N_12341,N_12314);
nand U12728 (N_12728,N_12277,N_12460);
and U12729 (N_12729,N_12368,N_12339);
and U12730 (N_12730,N_12389,N_12342);
and U12731 (N_12731,N_12458,N_12498);
and U12732 (N_12732,N_12411,N_12429);
xor U12733 (N_12733,N_12278,N_12498);
nor U12734 (N_12734,N_12491,N_12316);
nand U12735 (N_12735,N_12303,N_12273);
nand U12736 (N_12736,N_12299,N_12465);
or U12737 (N_12737,N_12388,N_12452);
nand U12738 (N_12738,N_12468,N_12289);
or U12739 (N_12739,N_12349,N_12484);
nor U12740 (N_12740,N_12414,N_12258);
nor U12741 (N_12741,N_12282,N_12387);
nor U12742 (N_12742,N_12460,N_12267);
xor U12743 (N_12743,N_12293,N_12325);
nor U12744 (N_12744,N_12353,N_12417);
nor U12745 (N_12745,N_12328,N_12332);
xnor U12746 (N_12746,N_12485,N_12269);
or U12747 (N_12747,N_12295,N_12414);
and U12748 (N_12748,N_12444,N_12449);
nand U12749 (N_12749,N_12401,N_12253);
xnor U12750 (N_12750,N_12635,N_12514);
nor U12751 (N_12751,N_12720,N_12622);
nand U12752 (N_12752,N_12505,N_12539);
xor U12753 (N_12753,N_12680,N_12709);
nand U12754 (N_12754,N_12699,N_12733);
nand U12755 (N_12755,N_12511,N_12577);
nand U12756 (N_12756,N_12633,N_12670);
nand U12757 (N_12757,N_12729,N_12638);
nand U12758 (N_12758,N_12634,N_12509);
or U12759 (N_12759,N_12665,N_12573);
and U12760 (N_12760,N_12678,N_12600);
nand U12761 (N_12761,N_12617,N_12535);
nor U12762 (N_12762,N_12717,N_12596);
nor U12763 (N_12763,N_12562,N_12609);
and U12764 (N_12764,N_12647,N_12570);
xor U12765 (N_12765,N_12740,N_12578);
and U12766 (N_12766,N_12523,N_12532);
or U12767 (N_12767,N_12704,N_12674);
and U12768 (N_12768,N_12676,N_12654);
or U12769 (N_12769,N_12736,N_12581);
xnor U12770 (N_12770,N_12594,N_12527);
or U12771 (N_12771,N_12555,N_12510);
and U12772 (N_12772,N_12521,N_12667);
nand U12773 (N_12773,N_12568,N_12544);
and U12774 (N_12774,N_12601,N_12681);
nor U12775 (N_12775,N_12648,N_12566);
nand U12776 (N_12776,N_12582,N_12520);
or U12777 (N_12777,N_12561,N_12675);
xnor U12778 (N_12778,N_12650,N_12627);
and U12779 (N_12779,N_12572,N_12529);
nand U12780 (N_12780,N_12735,N_12694);
nand U12781 (N_12781,N_12584,N_12557);
or U12782 (N_12782,N_12739,N_12628);
xor U12783 (N_12783,N_12715,N_12749);
nor U12784 (N_12784,N_12723,N_12525);
and U12785 (N_12785,N_12554,N_12513);
xor U12786 (N_12786,N_12642,N_12542);
or U12787 (N_12787,N_12574,N_12727);
or U12788 (N_12788,N_12560,N_12713);
nand U12789 (N_12789,N_12548,N_12579);
and U12790 (N_12790,N_12515,N_12576);
nand U12791 (N_12791,N_12631,N_12614);
nor U12792 (N_12792,N_12664,N_12517);
nand U12793 (N_12793,N_12508,N_12550);
or U12794 (N_12794,N_12666,N_12663);
or U12795 (N_12795,N_12575,N_12746);
or U12796 (N_12796,N_12538,N_12687);
nand U12797 (N_12797,N_12537,N_12690);
nor U12798 (N_12798,N_12545,N_12593);
or U12799 (N_12799,N_12553,N_12747);
xnor U12800 (N_12800,N_12571,N_12565);
and U12801 (N_12801,N_12526,N_12503);
xor U12802 (N_12802,N_12519,N_12688);
nand U12803 (N_12803,N_12697,N_12744);
nor U12804 (N_12804,N_12658,N_12522);
xnor U12805 (N_12805,N_12668,N_12705);
xor U12806 (N_12806,N_12543,N_12536);
nor U12807 (N_12807,N_12615,N_12602);
nor U12808 (N_12808,N_12656,N_12629);
nor U12809 (N_12809,N_12624,N_12604);
xor U12810 (N_12810,N_12748,N_12651);
xnor U12811 (N_12811,N_12673,N_12708);
or U12812 (N_12812,N_12618,N_12531);
xnor U12813 (N_12813,N_12707,N_12564);
nor U12814 (N_12814,N_12613,N_12605);
xor U12815 (N_12815,N_12590,N_12589);
nand U12816 (N_12816,N_12728,N_12696);
and U12817 (N_12817,N_12657,N_12702);
or U12818 (N_12818,N_12620,N_12644);
xnor U12819 (N_12819,N_12649,N_12541);
and U12820 (N_12820,N_12587,N_12655);
nand U12821 (N_12821,N_12731,N_12551);
nand U12822 (N_12822,N_12691,N_12712);
nor U12823 (N_12823,N_12661,N_12659);
nand U12824 (N_12824,N_12725,N_12559);
xnor U12825 (N_12825,N_12534,N_12684);
nor U12826 (N_12826,N_12586,N_12500);
and U12827 (N_12827,N_12563,N_12652);
and U12828 (N_12828,N_12645,N_12547);
xnor U12829 (N_12829,N_12507,N_12621);
nor U12830 (N_12830,N_12595,N_12518);
and U12831 (N_12831,N_12743,N_12679);
or U12832 (N_12832,N_12686,N_12730);
nor U12833 (N_12833,N_12610,N_12726);
nor U12834 (N_12834,N_12546,N_12626);
nor U12835 (N_12835,N_12672,N_12549);
nand U12836 (N_12836,N_12567,N_12682);
nand U12837 (N_12837,N_12716,N_12556);
nand U12838 (N_12838,N_12722,N_12701);
or U12839 (N_12839,N_12718,N_12700);
xor U12840 (N_12840,N_12552,N_12585);
xnor U12841 (N_12841,N_12512,N_12524);
nand U12842 (N_12842,N_12695,N_12693);
or U12843 (N_12843,N_12637,N_12737);
or U12844 (N_12844,N_12592,N_12703);
or U12845 (N_12845,N_12588,N_12641);
and U12846 (N_12846,N_12677,N_12643);
nand U12847 (N_12847,N_12741,N_12692);
nand U12848 (N_12848,N_12639,N_12714);
or U12849 (N_12849,N_12611,N_12612);
nor U12850 (N_12850,N_12516,N_12742);
xnor U12851 (N_12851,N_12683,N_12640);
nor U12852 (N_12852,N_12504,N_12734);
xnor U12853 (N_12853,N_12501,N_12528);
or U12854 (N_12854,N_12632,N_12671);
xnor U12855 (N_12855,N_12607,N_12623);
nor U12856 (N_12856,N_12502,N_12540);
or U12857 (N_12857,N_12558,N_12689);
or U12858 (N_12858,N_12598,N_12745);
and U12859 (N_12859,N_12706,N_12653);
and U12860 (N_12860,N_12580,N_12738);
nor U12861 (N_12861,N_12619,N_12599);
nand U12862 (N_12862,N_12630,N_12732);
nand U12863 (N_12863,N_12646,N_12662);
and U12864 (N_12864,N_12685,N_12711);
nor U12865 (N_12865,N_12698,N_12583);
nand U12866 (N_12866,N_12597,N_12533);
and U12867 (N_12867,N_12603,N_12616);
and U12868 (N_12868,N_12710,N_12719);
xor U12869 (N_12869,N_12625,N_12606);
nor U12870 (N_12870,N_12569,N_12608);
and U12871 (N_12871,N_12591,N_12724);
and U12872 (N_12872,N_12530,N_12506);
and U12873 (N_12873,N_12721,N_12636);
and U12874 (N_12874,N_12660,N_12669);
nor U12875 (N_12875,N_12523,N_12685);
and U12876 (N_12876,N_12538,N_12742);
nand U12877 (N_12877,N_12664,N_12627);
nor U12878 (N_12878,N_12625,N_12696);
or U12879 (N_12879,N_12571,N_12510);
nor U12880 (N_12880,N_12599,N_12500);
and U12881 (N_12881,N_12607,N_12696);
xnor U12882 (N_12882,N_12653,N_12605);
and U12883 (N_12883,N_12702,N_12653);
nand U12884 (N_12884,N_12630,N_12585);
nand U12885 (N_12885,N_12688,N_12629);
nand U12886 (N_12886,N_12619,N_12575);
nor U12887 (N_12887,N_12699,N_12647);
xor U12888 (N_12888,N_12567,N_12680);
xor U12889 (N_12889,N_12587,N_12515);
or U12890 (N_12890,N_12588,N_12502);
xnor U12891 (N_12891,N_12690,N_12554);
and U12892 (N_12892,N_12635,N_12504);
nor U12893 (N_12893,N_12687,N_12534);
nor U12894 (N_12894,N_12704,N_12590);
xnor U12895 (N_12895,N_12626,N_12602);
and U12896 (N_12896,N_12722,N_12725);
nor U12897 (N_12897,N_12595,N_12527);
xor U12898 (N_12898,N_12537,N_12743);
nand U12899 (N_12899,N_12628,N_12697);
xor U12900 (N_12900,N_12709,N_12696);
and U12901 (N_12901,N_12521,N_12612);
xnor U12902 (N_12902,N_12596,N_12549);
nand U12903 (N_12903,N_12666,N_12679);
or U12904 (N_12904,N_12621,N_12643);
nand U12905 (N_12905,N_12668,N_12687);
and U12906 (N_12906,N_12512,N_12700);
and U12907 (N_12907,N_12604,N_12642);
xor U12908 (N_12908,N_12517,N_12567);
nor U12909 (N_12909,N_12738,N_12658);
and U12910 (N_12910,N_12675,N_12625);
nand U12911 (N_12911,N_12669,N_12572);
nor U12912 (N_12912,N_12681,N_12518);
and U12913 (N_12913,N_12743,N_12651);
xnor U12914 (N_12914,N_12576,N_12569);
nand U12915 (N_12915,N_12661,N_12680);
xnor U12916 (N_12916,N_12598,N_12660);
xnor U12917 (N_12917,N_12624,N_12679);
or U12918 (N_12918,N_12534,N_12566);
nor U12919 (N_12919,N_12644,N_12509);
xnor U12920 (N_12920,N_12550,N_12669);
and U12921 (N_12921,N_12622,N_12587);
xor U12922 (N_12922,N_12599,N_12657);
nand U12923 (N_12923,N_12666,N_12561);
and U12924 (N_12924,N_12531,N_12572);
nand U12925 (N_12925,N_12664,N_12701);
and U12926 (N_12926,N_12692,N_12720);
nor U12927 (N_12927,N_12730,N_12603);
nor U12928 (N_12928,N_12556,N_12744);
nand U12929 (N_12929,N_12718,N_12595);
or U12930 (N_12930,N_12575,N_12552);
nor U12931 (N_12931,N_12602,N_12554);
nor U12932 (N_12932,N_12625,N_12502);
and U12933 (N_12933,N_12698,N_12637);
nand U12934 (N_12934,N_12525,N_12709);
xnor U12935 (N_12935,N_12576,N_12511);
and U12936 (N_12936,N_12640,N_12731);
xnor U12937 (N_12937,N_12687,N_12698);
nor U12938 (N_12938,N_12572,N_12549);
nand U12939 (N_12939,N_12522,N_12571);
xor U12940 (N_12940,N_12696,N_12536);
or U12941 (N_12941,N_12613,N_12618);
nor U12942 (N_12942,N_12513,N_12602);
and U12943 (N_12943,N_12703,N_12524);
and U12944 (N_12944,N_12748,N_12733);
and U12945 (N_12945,N_12537,N_12584);
and U12946 (N_12946,N_12556,N_12601);
or U12947 (N_12947,N_12518,N_12741);
or U12948 (N_12948,N_12738,N_12640);
or U12949 (N_12949,N_12579,N_12564);
and U12950 (N_12950,N_12508,N_12574);
or U12951 (N_12951,N_12600,N_12560);
and U12952 (N_12952,N_12516,N_12548);
or U12953 (N_12953,N_12663,N_12713);
and U12954 (N_12954,N_12662,N_12661);
or U12955 (N_12955,N_12720,N_12560);
nand U12956 (N_12956,N_12543,N_12566);
and U12957 (N_12957,N_12512,N_12608);
and U12958 (N_12958,N_12566,N_12711);
nor U12959 (N_12959,N_12541,N_12673);
xnor U12960 (N_12960,N_12680,N_12697);
nor U12961 (N_12961,N_12619,N_12678);
xnor U12962 (N_12962,N_12645,N_12512);
nor U12963 (N_12963,N_12699,N_12574);
xnor U12964 (N_12964,N_12607,N_12697);
nand U12965 (N_12965,N_12511,N_12711);
or U12966 (N_12966,N_12570,N_12663);
nand U12967 (N_12967,N_12546,N_12641);
nor U12968 (N_12968,N_12626,N_12687);
or U12969 (N_12969,N_12646,N_12722);
and U12970 (N_12970,N_12739,N_12615);
and U12971 (N_12971,N_12531,N_12581);
xnor U12972 (N_12972,N_12622,N_12670);
nand U12973 (N_12973,N_12744,N_12742);
nor U12974 (N_12974,N_12742,N_12571);
and U12975 (N_12975,N_12740,N_12695);
nor U12976 (N_12976,N_12542,N_12650);
xnor U12977 (N_12977,N_12736,N_12735);
nand U12978 (N_12978,N_12585,N_12606);
nand U12979 (N_12979,N_12515,N_12702);
nor U12980 (N_12980,N_12544,N_12597);
nor U12981 (N_12981,N_12504,N_12730);
xor U12982 (N_12982,N_12701,N_12535);
and U12983 (N_12983,N_12539,N_12653);
and U12984 (N_12984,N_12748,N_12641);
and U12985 (N_12985,N_12536,N_12745);
xnor U12986 (N_12986,N_12605,N_12524);
xor U12987 (N_12987,N_12580,N_12673);
xor U12988 (N_12988,N_12729,N_12633);
nor U12989 (N_12989,N_12636,N_12726);
nor U12990 (N_12990,N_12507,N_12744);
xnor U12991 (N_12991,N_12707,N_12517);
xnor U12992 (N_12992,N_12675,N_12576);
xor U12993 (N_12993,N_12591,N_12684);
or U12994 (N_12994,N_12656,N_12530);
nor U12995 (N_12995,N_12734,N_12500);
and U12996 (N_12996,N_12658,N_12746);
and U12997 (N_12997,N_12622,N_12573);
and U12998 (N_12998,N_12749,N_12546);
and U12999 (N_12999,N_12564,N_12528);
xnor U13000 (N_13000,N_12867,N_12994);
or U13001 (N_13001,N_12990,N_12848);
and U13002 (N_13002,N_12791,N_12775);
nand U13003 (N_13003,N_12750,N_12955);
nand U13004 (N_13004,N_12821,N_12871);
or U13005 (N_13005,N_12916,N_12830);
nor U13006 (N_13006,N_12999,N_12947);
xor U13007 (N_13007,N_12965,N_12964);
nand U13008 (N_13008,N_12929,N_12991);
nand U13009 (N_13009,N_12763,N_12900);
or U13010 (N_13010,N_12940,N_12767);
nor U13011 (N_13011,N_12813,N_12860);
nand U13012 (N_13012,N_12805,N_12910);
or U13013 (N_13013,N_12928,N_12981);
or U13014 (N_13014,N_12765,N_12825);
nor U13015 (N_13015,N_12943,N_12890);
and U13016 (N_13016,N_12762,N_12864);
xnor U13017 (N_13017,N_12812,N_12939);
and U13018 (N_13018,N_12970,N_12880);
nand U13019 (N_13019,N_12780,N_12945);
nor U13020 (N_13020,N_12996,N_12925);
nand U13021 (N_13021,N_12835,N_12893);
xnor U13022 (N_13022,N_12877,N_12870);
and U13023 (N_13023,N_12809,N_12901);
nand U13024 (N_13024,N_12799,N_12930);
or U13025 (N_13025,N_12972,N_12833);
xor U13026 (N_13026,N_12934,N_12841);
or U13027 (N_13027,N_12754,N_12752);
or U13028 (N_13028,N_12909,N_12976);
and U13029 (N_13029,N_12853,N_12951);
and U13030 (N_13030,N_12963,N_12790);
and U13031 (N_13031,N_12984,N_12923);
and U13032 (N_13032,N_12859,N_12985);
and U13033 (N_13033,N_12997,N_12768);
nand U13034 (N_13034,N_12779,N_12856);
or U13035 (N_13035,N_12800,N_12850);
nand U13036 (N_13036,N_12846,N_12926);
or U13037 (N_13037,N_12807,N_12832);
nand U13038 (N_13038,N_12865,N_12887);
xnor U13039 (N_13039,N_12814,N_12808);
or U13040 (N_13040,N_12952,N_12834);
nor U13041 (N_13041,N_12975,N_12840);
and U13042 (N_13042,N_12989,N_12785);
or U13043 (N_13043,N_12881,N_12849);
nand U13044 (N_13044,N_12914,N_12896);
or U13045 (N_13045,N_12897,N_12944);
nor U13046 (N_13046,N_12776,N_12879);
and U13047 (N_13047,N_12782,N_12756);
xnor U13048 (N_13048,N_12917,N_12953);
nand U13049 (N_13049,N_12918,N_12962);
and U13050 (N_13050,N_12804,N_12761);
nand U13051 (N_13051,N_12878,N_12995);
or U13052 (N_13052,N_12874,N_12854);
xnor U13053 (N_13053,N_12902,N_12772);
nand U13054 (N_13054,N_12827,N_12869);
nand U13055 (N_13055,N_12764,N_12933);
xnor U13056 (N_13056,N_12950,N_12771);
or U13057 (N_13057,N_12758,N_12942);
or U13058 (N_13058,N_12815,N_12801);
nor U13059 (N_13059,N_12967,N_12773);
nor U13060 (N_13060,N_12786,N_12937);
and U13061 (N_13061,N_12872,N_12898);
xor U13062 (N_13062,N_12993,N_12770);
nor U13063 (N_13063,N_12875,N_12863);
xor U13064 (N_13064,N_12883,N_12783);
and U13065 (N_13065,N_12988,N_12968);
xor U13066 (N_13066,N_12811,N_12847);
and U13067 (N_13067,N_12802,N_12982);
nand U13068 (N_13068,N_12857,N_12960);
xor U13069 (N_13069,N_12938,N_12803);
nand U13070 (N_13070,N_12983,N_12885);
or U13071 (N_13071,N_12904,N_12793);
nand U13072 (N_13072,N_12977,N_12816);
xnor U13073 (N_13073,N_12959,N_12873);
xor U13074 (N_13074,N_12819,N_12882);
xor U13075 (N_13075,N_12911,N_12852);
nand U13076 (N_13076,N_12753,N_12810);
or U13077 (N_13077,N_12927,N_12876);
and U13078 (N_13078,N_12855,N_12766);
or U13079 (N_13079,N_12843,N_12941);
or U13080 (N_13080,N_12913,N_12836);
nor U13081 (N_13081,N_12795,N_12755);
xnor U13082 (N_13082,N_12956,N_12922);
and U13083 (N_13083,N_12888,N_12792);
and U13084 (N_13084,N_12824,N_12978);
or U13085 (N_13085,N_12891,N_12778);
and U13086 (N_13086,N_12957,N_12806);
nor U13087 (N_13087,N_12759,N_12966);
and U13088 (N_13088,N_12895,N_12788);
nand U13089 (N_13089,N_12822,N_12920);
and U13090 (N_13090,N_12936,N_12931);
and U13091 (N_13091,N_12921,N_12915);
nor U13092 (N_13092,N_12907,N_12861);
xor U13093 (N_13093,N_12839,N_12906);
or U13094 (N_13094,N_12992,N_12796);
and U13095 (N_13095,N_12817,N_12889);
nand U13096 (N_13096,N_12862,N_12798);
or U13097 (N_13097,N_12844,N_12908);
and U13098 (N_13098,N_12829,N_12831);
and U13099 (N_13099,N_12971,N_12774);
or U13100 (N_13100,N_12884,N_12858);
nand U13101 (N_13101,N_12919,N_12946);
and U13102 (N_13102,N_12912,N_12818);
xnor U13103 (N_13103,N_12838,N_12837);
xnor U13104 (N_13104,N_12842,N_12826);
nand U13105 (N_13105,N_12892,N_12979);
nand U13106 (N_13106,N_12769,N_12899);
nand U13107 (N_13107,N_12935,N_12787);
or U13108 (N_13108,N_12998,N_12932);
nor U13109 (N_13109,N_12924,N_12948);
or U13110 (N_13110,N_12903,N_12797);
xnor U13111 (N_13111,N_12760,N_12777);
xnor U13112 (N_13112,N_12894,N_12784);
xnor U13113 (N_13113,N_12820,N_12828);
or U13114 (N_13114,N_12781,N_12751);
and U13115 (N_13115,N_12986,N_12969);
nor U13116 (N_13116,N_12866,N_12954);
nor U13117 (N_13117,N_12905,N_12868);
or U13118 (N_13118,N_12973,N_12794);
nor U13119 (N_13119,N_12789,N_12757);
nand U13120 (N_13120,N_12949,N_12987);
xnor U13121 (N_13121,N_12886,N_12961);
or U13122 (N_13122,N_12974,N_12851);
and U13123 (N_13123,N_12845,N_12980);
nor U13124 (N_13124,N_12823,N_12958);
nand U13125 (N_13125,N_12891,N_12987);
and U13126 (N_13126,N_12869,N_12953);
xor U13127 (N_13127,N_12831,N_12973);
and U13128 (N_13128,N_12824,N_12875);
or U13129 (N_13129,N_12836,N_12821);
nand U13130 (N_13130,N_12908,N_12903);
nand U13131 (N_13131,N_12830,N_12987);
xor U13132 (N_13132,N_12949,N_12843);
nand U13133 (N_13133,N_12783,N_12763);
nand U13134 (N_13134,N_12959,N_12757);
xor U13135 (N_13135,N_12814,N_12819);
xor U13136 (N_13136,N_12917,N_12915);
nand U13137 (N_13137,N_12753,N_12908);
and U13138 (N_13138,N_12792,N_12807);
or U13139 (N_13139,N_12816,N_12937);
and U13140 (N_13140,N_12850,N_12798);
and U13141 (N_13141,N_12780,N_12862);
or U13142 (N_13142,N_12800,N_12873);
or U13143 (N_13143,N_12890,N_12756);
nor U13144 (N_13144,N_12864,N_12882);
xor U13145 (N_13145,N_12806,N_12912);
nand U13146 (N_13146,N_12769,N_12836);
or U13147 (N_13147,N_12759,N_12807);
nor U13148 (N_13148,N_12840,N_12862);
and U13149 (N_13149,N_12943,N_12989);
nor U13150 (N_13150,N_12890,N_12764);
nand U13151 (N_13151,N_12780,N_12793);
or U13152 (N_13152,N_12910,N_12845);
nor U13153 (N_13153,N_12840,N_12878);
or U13154 (N_13154,N_12785,N_12964);
or U13155 (N_13155,N_12811,N_12922);
nand U13156 (N_13156,N_12884,N_12759);
nor U13157 (N_13157,N_12799,N_12820);
xor U13158 (N_13158,N_12808,N_12866);
nor U13159 (N_13159,N_12851,N_12867);
or U13160 (N_13160,N_12753,N_12987);
xnor U13161 (N_13161,N_12845,N_12904);
or U13162 (N_13162,N_12808,N_12974);
or U13163 (N_13163,N_12943,N_12753);
or U13164 (N_13164,N_12895,N_12830);
nor U13165 (N_13165,N_12991,N_12851);
or U13166 (N_13166,N_12785,N_12945);
and U13167 (N_13167,N_12896,N_12764);
nor U13168 (N_13168,N_12828,N_12885);
xor U13169 (N_13169,N_12784,N_12977);
or U13170 (N_13170,N_12767,N_12876);
xor U13171 (N_13171,N_12819,N_12772);
xnor U13172 (N_13172,N_12898,N_12808);
or U13173 (N_13173,N_12991,N_12804);
or U13174 (N_13174,N_12887,N_12772);
nand U13175 (N_13175,N_12934,N_12891);
and U13176 (N_13176,N_12825,N_12908);
xor U13177 (N_13177,N_12935,N_12828);
nor U13178 (N_13178,N_12852,N_12965);
and U13179 (N_13179,N_12970,N_12948);
or U13180 (N_13180,N_12770,N_12861);
or U13181 (N_13181,N_12766,N_12966);
or U13182 (N_13182,N_12816,N_12904);
xor U13183 (N_13183,N_12816,N_12783);
xnor U13184 (N_13184,N_12929,N_12898);
xor U13185 (N_13185,N_12769,N_12995);
or U13186 (N_13186,N_12805,N_12885);
nor U13187 (N_13187,N_12840,N_12845);
xnor U13188 (N_13188,N_12998,N_12801);
nand U13189 (N_13189,N_12904,N_12886);
xnor U13190 (N_13190,N_12837,N_12893);
nor U13191 (N_13191,N_12751,N_12948);
nor U13192 (N_13192,N_12804,N_12842);
and U13193 (N_13193,N_12909,N_12987);
nand U13194 (N_13194,N_12933,N_12760);
xor U13195 (N_13195,N_12932,N_12839);
nor U13196 (N_13196,N_12771,N_12784);
or U13197 (N_13197,N_12892,N_12964);
or U13198 (N_13198,N_12882,N_12797);
or U13199 (N_13199,N_12921,N_12950);
nand U13200 (N_13200,N_12864,N_12763);
or U13201 (N_13201,N_12930,N_12864);
nor U13202 (N_13202,N_12973,N_12770);
xnor U13203 (N_13203,N_12808,N_12764);
nor U13204 (N_13204,N_12883,N_12796);
nand U13205 (N_13205,N_12952,N_12900);
nor U13206 (N_13206,N_12829,N_12871);
xor U13207 (N_13207,N_12905,N_12931);
or U13208 (N_13208,N_12762,N_12954);
or U13209 (N_13209,N_12902,N_12966);
or U13210 (N_13210,N_12827,N_12995);
xor U13211 (N_13211,N_12965,N_12969);
and U13212 (N_13212,N_12868,N_12910);
and U13213 (N_13213,N_12784,N_12907);
or U13214 (N_13214,N_12851,N_12971);
nand U13215 (N_13215,N_12897,N_12866);
xnor U13216 (N_13216,N_12780,N_12893);
nand U13217 (N_13217,N_12876,N_12933);
and U13218 (N_13218,N_12890,N_12754);
nor U13219 (N_13219,N_12941,N_12833);
and U13220 (N_13220,N_12928,N_12889);
or U13221 (N_13221,N_12833,N_12860);
and U13222 (N_13222,N_12953,N_12761);
and U13223 (N_13223,N_12823,N_12999);
xnor U13224 (N_13224,N_12975,N_12953);
nor U13225 (N_13225,N_12992,N_12799);
and U13226 (N_13226,N_12766,N_12844);
nand U13227 (N_13227,N_12901,N_12880);
and U13228 (N_13228,N_12751,N_12970);
xnor U13229 (N_13229,N_12754,N_12894);
xnor U13230 (N_13230,N_12786,N_12750);
or U13231 (N_13231,N_12841,N_12875);
xor U13232 (N_13232,N_12929,N_12772);
and U13233 (N_13233,N_12962,N_12847);
nor U13234 (N_13234,N_12855,N_12944);
or U13235 (N_13235,N_12793,N_12851);
or U13236 (N_13236,N_12839,N_12847);
xnor U13237 (N_13237,N_12990,N_12946);
xor U13238 (N_13238,N_12920,N_12860);
xor U13239 (N_13239,N_12937,N_12861);
xor U13240 (N_13240,N_12753,N_12803);
nor U13241 (N_13241,N_12897,N_12819);
nor U13242 (N_13242,N_12880,N_12800);
nor U13243 (N_13243,N_12897,N_12769);
nor U13244 (N_13244,N_12986,N_12835);
or U13245 (N_13245,N_12851,N_12759);
nor U13246 (N_13246,N_12837,N_12865);
nor U13247 (N_13247,N_12814,N_12813);
nand U13248 (N_13248,N_12988,N_12822);
nor U13249 (N_13249,N_12950,N_12817);
xnor U13250 (N_13250,N_13228,N_13238);
nor U13251 (N_13251,N_13144,N_13055);
xor U13252 (N_13252,N_13075,N_13185);
nor U13253 (N_13253,N_13081,N_13007);
nor U13254 (N_13254,N_13219,N_13000);
nor U13255 (N_13255,N_13119,N_13134);
and U13256 (N_13256,N_13147,N_13194);
and U13257 (N_13257,N_13064,N_13243);
xnor U13258 (N_13258,N_13038,N_13042);
nor U13259 (N_13259,N_13120,N_13034);
and U13260 (N_13260,N_13188,N_13218);
nand U13261 (N_13261,N_13244,N_13186);
or U13262 (N_13262,N_13125,N_13065);
and U13263 (N_13263,N_13221,N_13091);
or U13264 (N_13264,N_13140,N_13019);
or U13265 (N_13265,N_13090,N_13168);
nor U13266 (N_13266,N_13138,N_13003);
or U13267 (N_13267,N_13180,N_13040);
and U13268 (N_13268,N_13234,N_13110);
nor U13269 (N_13269,N_13237,N_13107);
xnor U13270 (N_13270,N_13214,N_13208);
nand U13271 (N_13271,N_13156,N_13176);
nor U13272 (N_13272,N_13230,N_13009);
and U13273 (N_13273,N_13128,N_13210);
and U13274 (N_13274,N_13171,N_13068);
or U13275 (N_13275,N_13053,N_13002);
or U13276 (N_13276,N_13051,N_13056);
or U13277 (N_13277,N_13071,N_13044);
nand U13278 (N_13278,N_13101,N_13212);
nor U13279 (N_13279,N_13121,N_13111);
or U13280 (N_13280,N_13223,N_13058);
and U13281 (N_13281,N_13112,N_13173);
and U13282 (N_13282,N_13200,N_13132);
xor U13283 (N_13283,N_13116,N_13072);
and U13284 (N_13284,N_13103,N_13117);
nand U13285 (N_13285,N_13189,N_13216);
nand U13286 (N_13286,N_13215,N_13149);
nand U13287 (N_13287,N_13067,N_13073);
nand U13288 (N_13288,N_13145,N_13182);
and U13289 (N_13289,N_13164,N_13157);
xor U13290 (N_13290,N_13241,N_13197);
nor U13291 (N_13291,N_13059,N_13135);
nand U13292 (N_13292,N_13233,N_13008);
xnor U13293 (N_13293,N_13001,N_13232);
nor U13294 (N_13294,N_13082,N_13196);
xor U13295 (N_13295,N_13021,N_13027);
and U13296 (N_13296,N_13098,N_13158);
or U13297 (N_13297,N_13222,N_13187);
xnor U13298 (N_13298,N_13165,N_13026);
xnor U13299 (N_13299,N_13113,N_13122);
xnor U13300 (N_13300,N_13015,N_13025);
and U13301 (N_13301,N_13209,N_13195);
nor U13302 (N_13302,N_13037,N_13154);
nand U13303 (N_13303,N_13069,N_13052);
nand U13304 (N_13304,N_13050,N_13179);
xor U13305 (N_13305,N_13202,N_13220);
xnor U13306 (N_13306,N_13126,N_13192);
nor U13307 (N_13307,N_13018,N_13203);
nor U13308 (N_13308,N_13242,N_13246);
nor U13309 (N_13309,N_13004,N_13093);
nor U13310 (N_13310,N_13177,N_13161);
or U13311 (N_13311,N_13205,N_13136);
and U13312 (N_13312,N_13229,N_13178);
xor U13313 (N_13313,N_13118,N_13014);
nand U13314 (N_13314,N_13123,N_13077);
nand U13315 (N_13315,N_13028,N_13199);
nand U13316 (N_13316,N_13049,N_13029);
xnor U13317 (N_13317,N_13137,N_13170);
and U13318 (N_13318,N_13226,N_13247);
xnor U13319 (N_13319,N_13041,N_13109);
xor U13320 (N_13320,N_13204,N_13023);
and U13321 (N_13321,N_13240,N_13054);
nand U13322 (N_13322,N_13142,N_13013);
nor U13323 (N_13323,N_13146,N_13150);
xor U13324 (N_13324,N_13160,N_13236);
nor U13325 (N_13325,N_13063,N_13239);
xnor U13326 (N_13326,N_13087,N_13151);
nor U13327 (N_13327,N_13163,N_13048);
xnor U13328 (N_13328,N_13245,N_13094);
xnor U13329 (N_13329,N_13036,N_13005);
nor U13330 (N_13330,N_13035,N_13129);
nand U13331 (N_13331,N_13062,N_13190);
or U13332 (N_13332,N_13235,N_13224);
and U13333 (N_13333,N_13159,N_13102);
and U13334 (N_13334,N_13083,N_13088);
nor U13335 (N_13335,N_13078,N_13183);
and U13336 (N_13336,N_13012,N_13175);
or U13337 (N_13337,N_13057,N_13061);
nor U13338 (N_13338,N_13024,N_13174);
nor U13339 (N_13339,N_13089,N_13039);
nand U13340 (N_13340,N_13152,N_13079);
or U13341 (N_13341,N_13033,N_13086);
and U13342 (N_13342,N_13249,N_13045);
xor U13343 (N_13343,N_13172,N_13115);
or U13344 (N_13344,N_13031,N_13108);
and U13345 (N_13345,N_13106,N_13153);
or U13346 (N_13346,N_13084,N_13131);
nor U13347 (N_13347,N_13201,N_13043);
or U13348 (N_13348,N_13198,N_13162);
or U13349 (N_13349,N_13248,N_13030);
and U13350 (N_13350,N_13076,N_13207);
nor U13351 (N_13351,N_13020,N_13217);
or U13352 (N_13352,N_13085,N_13227);
nand U13353 (N_13353,N_13167,N_13010);
or U13354 (N_13354,N_13022,N_13127);
and U13355 (N_13355,N_13011,N_13006);
xnor U13356 (N_13356,N_13032,N_13046);
nor U13357 (N_13357,N_13193,N_13066);
xor U13358 (N_13358,N_13206,N_13096);
nor U13359 (N_13359,N_13092,N_13099);
or U13360 (N_13360,N_13017,N_13184);
or U13361 (N_13361,N_13141,N_13100);
and U13362 (N_13362,N_13225,N_13016);
and U13363 (N_13363,N_13080,N_13169);
nor U13364 (N_13364,N_13060,N_13191);
nand U13365 (N_13365,N_13105,N_13097);
nor U13366 (N_13366,N_13133,N_13231);
and U13367 (N_13367,N_13211,N_13070);
and U13368 (N_13368,N_13148,N_13074);
xor U13369 (N_13369,N_13124,N_13047);
xnor U13370 (N_13370,N_13104,N_13139);
xor U13371 (N_13371,N_13213,N_13155);
xor U13372 (N_13372,N_13181,N_13166);
and U13373 (N_13373,N_13095,N_13130);
nor U13374 (N_13374,N_13114,N_13143);
or U13375 (N_13375,N_13242,N_13194);
xnor U13376 (N_13376,N_13170,N_13210);
or U13377 (N_13377,N_13041,N_13143);
xor U13378 (N_13378,N_13084,N_13238);
nand U13379 (N_13379,N_13105,N_13089);
or U13380 (N_13380,N_13019,N_13054);
and U13381 (N_13381,N_13108,N_13221);
or U13382 (N_13382,N_13237,N_13240);
nand U13383 (N_13383,N_13166,N_13012);
nand U13384 (N_13384,N_13144,N_13122);
nand U13385 (N_13385,N_13068,N_13034);
or U13386 (N_13386,N_13083,N_13198);
nand U13387 (N_13387,N_13098,N_13054);
xor U13388 (N_13388,N_13026,N_13225);
nand U13389 (N_13389,N_13093,N_13230);
or U13390 (N_13390,N_13044,N_13042);
or U13391 (N_13391,N_13120,N_13020);
and U13392 (N_13392,N_13093,N_13135);
xnor U13393 (N_13393,N_13029,N_13146);
or U13394 (N_13394,N_13229,N_13246);
and U13395 (N_13395,N_13207,N_13090);
xnor U13396 (N_13396,N_13237,N_13096);
and U13397 (N_13397,N_13225,N_13129);
nor U13398 (N_13398,N_13052,N_13014);
or U13399 (N_13399,N_13188,N_13044);
nand U13400 (N_13400,N_13044,N_13118);
and U13401 (N_13401,N_13218,N_13132);
nor U13402 (N_13402,N_13189,N_13246);
nand U13403 (N_13403,N_13211,N_13217);
nor U13404 (N_13404,N_13174,N_13005);
nand U13405 (N_13405,N_13044,N_13242);
or U13406 (N_13406,N_13079,N_13024);
nand U13407 (N_13407,N_13041,N_13169);
nor U13408 (N_13408,N_13128,N_13075);
nand U13409 (N_13409,N_13157,N_13031);
and U13410 (N_13410,N_13243,N_13076);
or U13411 (N_13411,N_13029,N_13203);
xor U13412 (N_13412,N_13087,N_13023);
and U13413 (N_13413,N_13233,N_13220);
xnor U13414 (N_13414,N_13248,N_13060);
xnor U13415 (N_13415,N_13220,N_13194);
xor U13416 (N_13416,N_13101,N_13178);
nand U13417 (N_13417,N_13215,N_13130);
and U13418 (N_13418,N_13157,N_13104);
nor U13419 (N_13419,N_13191,N_13136);
and U13420 (N_13420,N_13195,N_13236);
and U13421 (N_13421,N_13242,N_13057);
xor U13422 (N_13422,N_13119,N_13044);
nor U13423 (N_13423,N_13084,N_13190);
xor U13424 (N_13424,N_13036,N_13223);
xor U13425 (N_13425,N_13116,N_13178);
xnor U13426 (N_13426,N_13081,N_13239);
nand U13427 (N_13427,N_13134,N_13230);
nor U13428 (N_13428,N_13015,N_13067);
nand U13429 (N_13429,N_13086,N_13213);
xnor U13430 (N_13430,N_13204,N_13025);
or U13431 (N_13431,N_13113,N_13175);
xor U13432 (N_13432,N_13205,N_13052);
or U13433 (N_13433,N_13225,N_13233);
xnor U13434 (N_13434,N_13224,N_13096);
and U13435 (N_13435,N_13196,N_13200);
or U13436 (N_13436,N_13166,N_13011);
or U13437 (N_13437,N_13013,N_13188);
or U13438 (N_13438,N_13068,N_13067);
nor U13439 (N_13439,N_13075,N_13245);
and U13440 (N_13440,N_13224,N_13142);
xnor U13441 (N_13441,N_13025,N_13049);
xnor U13442 (N_13442,N_13216,N_13147);
and U13443 (N_13443,N_13051,N_13093);
xor U13444 (N_13444,N_13210,N_13071);
or U13445 (N_13445,N_13160,N_13180);
or U13446 (N_13446,N_13144,N_13025);
nand U13447 (N_13447,N_13081,N_13140);
xor U13448 (N_13448,N_13148,N_13072);
nor U13449 (N_13449,N_13078,N_13162);
nor U13450 (N_13450,N_13174,N_13049);
xnor U13451 (N_13451,N_13068,N_13231);
or U13452 (N_13452,N_13144,N_13141);
nor U13453 (N_13453,N_13091,N_13054);
nor U13454 (N_13454,N_13200,N_13008);
and U13455 (N_13455,N_13173,N_13085);
and U13456 (N_13456,N_13232,N_13112);
xor U13457 (N_13457,N_13010,N_13140);
xor U13458 (N_13458,N_13163,N_13108);
or U13459 (N_13459,N_13110,N_13008);
or U13460 (N_13460,N_13136,N_13122);
xnor U13461 (N_13461,N_13078,N_13095);
nor U13462 (N_13462,N_13164,N_13201);
or U13463 (N_13463,N_13033,N_13196);
xnor U13464 (N_13464,N_13070,N_13170);
or U13465 (N_13465,N_13107,N_13119);
nand U13466 (N_13466,N_13046,N_13239);
xor U13467 (N_13467,N_13084,N_13023);
and U13468 (N_13468,N_13115,N_13240);
or U13469 (N_13469,N_13139,N_13230);
and U13470 (N_13470,N_13044,N_13007);
xnor U13471 (N_13471,N_13063,N_13112);
xnor U13472 (N_13472,N_13220,N_13002);
nor U13473 (N_13473,N_13069,N_13193);
xnor U13474 (N_13474,N_13084,N_13050);
nor U13475 (N_13475,N_13012,N_13213);
or U13476 (N_13476,N_13088,N_13015);
xor U13477 (N_13477,N_13223,N_13039);
nand U13478 (N_13478,N_13194,N_13232);
nand U13479 (N_13479,N_13185,N_13038);
or U13480 (N_13480,N_13196,N_13202);
nor U13481 (N_13481,N_13035,N_13181);
and U13482 (N_13482,N_13099,N_13161);
nand U13483 (N_13483,N_13117,N_13060);
and U13484 (N_13484,N_13248,N_13037);
or U13485 (N_13485,N_13165,N_13187);
xor U13486 (N_13486,N_13048,N_13157);
and U13487 (N_13487,N_13128,N_13177);
xnor U13488 (N_13488,N_13139,N_13093);
nor U13489 (N_13489,N_13211,N_13074);
and U13490 (N_13490,N_13173,N_13044);
nor U13491 (N_13491,N_13054,N_13238);
xor U13492 (N_13492,N_13185,N_13049);
nand U13493 (N_13493,N_13060,N_13241);
nand U13494 (N_13494,N_13198,N_13171);
nor U13495 (N_13495,N_13146,N_13028);
or U13496 (N_13496,N_13058,N_13161);
or U13497 (N_13497,N_13058,N_13104);
nand U13498 (N_13498,N_13043,N_13233);
xor U13499 (N_13499,N_13154,N_13093);
xnor U13500 (N_13500,N_13411,N_13442);
nand U13501 (N_13501,N_13317,N_13365);
nand U13502 (N_13502,N_13356,N_13284);
xnor U13503 (N_13503,N_13422,N_13483);
nor U13504 (N_13504,N_13450,N_13331);
xnor U13505 (N_13505,N_13440,N_13462);
xnor U13506 (N_13506,N_13354,N_13302);
nor U13507 (N_13507,N_13385,N_13330);
xnor U13508 (N_13508,N_13352,N_13324);
nand U13509 (N_13509,N_13339,N_13412);
nand U13510 (N_13510,N_13493,N_13466);
and U13511 (N_13511,N_13413,N_13437);
xor U13512 (N_13512,N_13328,N_13383);
xnor U13513 (N_13513,N_13272,N_13418);
xor U13514 (N_13514,N_13469,N_13311);
nor U13515 (N_13515,N_13260,N_13405);
xor U13516 (N_13516,N_13305,N_13306);
xor U13517 (N_13517,N_13435,N_13491);
and U13518 (N_13518,N_13485,N_13338);
xor U13519 (N_13519,N_13386,N_13291);
or U13520 (N_13520,N_13275,N_13427);
nor U13521 (N_13521,N_13467,N_13479);
nand U13522 (N_13522,N_13280,N_13313);
nand U13523 (N_13523,N_13406,N_13309);
nor U13524 (N_13524,N_13451,N_13375);
nor U13525 (N_13525,N_13267,N_13318);
nand U13526 (N_13526,N_13428,N_13400);
nand U13527 (N_13527,N_13464,N_13323);
and U13528 (N_13528,N_13351,N_13327);
xnor U13529 (N_13529,N_13399,N_13376);
nand U13530 (N_13530,N_13460,N_13395);
xnor U13531 (N_13531,N_13377,N_13388);
nand U13532 (N_13532,N_13310,N_13304);
xnor U13533 (N_13533,N_13307,N_13370);
xnor U13534 (N_13534,N_13256,N_13369);
nand U13535 (N_13535,N_13329,N_13264);
nor U13536 (N_13536,N_13495,N_13315);
nand U13537 (N_13537,N_13362,N_13490);
nand U13538 (N_13538,N_13484,N_13308);
or U13539 (N_13539,N_13340,N_13364);
xnor U13540 (N_13540,N_13251,N_13455);
and U13541 (N_13541,N_13278,N_13293);
nand U13542 (N_13542,N_13394,N_13259);
and U13543 (N_13543,N_13470,N_13367);
or U13544 (N_13544,N_13456,N_13414);
and U13545 (N_13545,N_13443,N_13453);
or U13546 (N_13546,N_13392,N_13343);
and U13547 (N_13547,N_13431,N_13445);
nor U13548 (N_13548,N_13446,N_13333);
and U13549 (N_13549,N_13289,N_13266);
xor U13550 (N_13550,N_13274,N_13444);
nor U13551 (N_13551,N_13316,N_13410);
and U13552 (N_13552,N_13268,N_13417);
or U13553 (N_13553,N_13403,N_13371);
xor U13554 (N_13554,N_13404,N_13421);
xnor U13555 (N_13555,N_13265,N_13285);
xor U13556 (N_13556,N_13252,N_13349);
xor U13557 (N_13557,N_13258,N_13429);
nand U13558 (N_13558,N_13345,N_13294);
or U13559 (N_13559,N_13496,N_13457);
nand U13560 (N_13560,N_13472,N_13374);
xor U13561 (N_13561,N_13459,N_13497);
and U13562 (N_13562,N_13312,N_13426);
and U13563 (N_13563,N_13334,N_13419);
or U13564 (N_13564,N_13290,N_13295);
nand U13565 (N_13565,N_13322,N_13487);
and U13566 (N_13566,N_13301,N_13270);
or U13567 (N_13567,N_13436,N_13281);
nand U13568 (N_13568,N_13441,N_13353);
xor U13569 (N_13569,N_13468,N_13432);
or U13570 (N_13570,N_13409,N_13366);
or U13571 (N_13571,N_13262,N_13297);
nor U13572 (N_13572,N_13398,N_13286);
xor U13573 (N_13573,N_13321,N_13299);
and U13574 (N_13574,N_13360,N_13424);
xnor U13575 (N_13575,N_13279,N_13300);
nor U13576 (N_13576,N_13430,N_13389);
and U13577 (N_13577,N_13402,N_13350);
nand U13578 (N_13578,N_13449,N_13499);
nand U13579 (N_13579,N_13282,N_13346);
and U13580 (N_13580,N_13434,N_13425);
or U13581 (N_13581,N_13271,N_13397);
or U13582 (N_13582,N_13373,N_13257);
or U13583 (N_13583,N_13255,N_13387);
xnor U13584 (N_13584,N_13348,N_13269);
and U13585 (N_13585,N_13382,N_13277);
nand U13586 (N_13586,N_13420,N_13361);
xor U13587 (N_13587,N_13452,N_13489);
nor U13588 (N_13588,N_13358,N_13498);
or U13589 (N_13589,N_13465,N_13481);
xnor U13590 (N_13590,N_13475,N_13474);
and U13591 (N_13591,N_13471,N_13378);
nand U13592 (N_13592,N_13433,N_13492);
and U13593 (N_13593,N_13261,N_13320);
and U13594 (N_13594,N_13407,N_13336);
xnor U13595 (N_13595,N_13296,N_13298);
and U13596 (N_13596,N_13253,N_13303);
nand U13597 (N_13597,N_13314,N_13494);
nor U13598 (N_13598,N_13273,N_13488);
xor U13599 (N_13599,N_13380,N_13393);
xor U13600 (N_13600,N_13391,N_13384);
xnor U13601 (N_13601,N_13372,N_13335);
nor U13602 (N_13602,N_13288,N_13416);
xor U13603 (N_13603,N_13423,N_13477);
or U13604 (N_13604,N_13381,N_13355);
nand U13605 (N_13605,N_13357,N_13458);
xnor U13606 (N_13606,N_13415,N_13454);
and U13607 (N_13607,N_13447,N_13448);
or U13608 (N_13608,N_13401,N_13254);
nor U13609 (N_13609,N_13359,N_13482);
xnor U13610 (N_13610,N_13463,N_13480);
and U13611 (N_13611,N_13473,N_13344);
or U13612 (N_13612,N_13363,N_13250);
nor U13613 (N_13613,N_13476,N_13379);
or U13614 (N_13614,N_13332,N_13287);
nor U13615 (N_13615,N_13337,N_13408);
and U13616 (N_13616,N_13292,N_13439);
and U13617 (N_13617,N_13438,N_13325);
and U13618 (N_13618,N_13368,N_13461);
nand U13619 (N_13619,N_13486,N_13283);
nor U13620 (N_13620,N_13276,N_13263);
nand U13621 (N_13621,N_13347,N_13319);
nand U13622 (N_13622,N_13390,N_13326);
nor U13623 (N_13623,N_13396,N_13341);
or U13624 (N_13624,N_13478,N_13342);
nor U13625 (N_13625,N_13250,N_13433);
and U13626 (N_13626,N_13469,N_13461);
xor U13627 (N_13627,N_13326,N_13275);
xor U13628 (N_13628,N_13377,N_13426);
nor U13629 (N_13629,N_13399,N_13252);
or U13630 (N_13630,N_13451,N_13340);
nand U13631 (N_13631,N_13346,N_13419);
nor U13632 (N_13632,N_13484,N_13257);
nor U13633 (N_13633,N_13375,N_13388);
nand U13634 (N_13634,N_13322,N_13411);
xor U13635 (N_13635,N_13376,N_13280);
nand U13636 (N_13636,N_13488,N_13382);
and U13637 (N_13637,N_13317,N_13453);
nor U13638 (N_13638,N_13316,N_13390);
or U13639 (N_13639,N_13318,N_13284);
nor U13640 (N_13640,N_13290,N_13338);
and U13641 (N_13641,N_13389,N_13473);
nand U13642 (N_13642,N_13261,N_13416);
or U13643 (N_13643,N_13337,N_13291);
nor U13644 (N_13644,N_13363,N_13417);
nor U13645 (N_13645,N_13468,N_13253);
xor U13646 (N_13646,N_13450,N_13357);
xor U13647 (N_13647,N_13375,N_13428);
nand U13648 (N_13648,N_13258,N_13361);
or U13649 (N_13649,N_13350,N_13290);
nor U13650 (N_13650,N_13437,N_13442);
nand U13651 (N_13651,N_13255,N_13340);
nand U13652 (N_13652,N_13451,N_13433);
nand U13653 (N_13653,N_13347,N_13413);
nand U13654 (N_13654,N_13266,N_13316);
or U13655 (N_13655,N_13486,N_13346);
nand U13656 (N_13656,N_13398,N_13297);
nand U13657 (N_13657,N_13284,N_13405);
nor U13658 (N_13658,N_13301,N_13337);
or U13659 (N_13659,N_13256,N_13465);
and U13660 (N_13660,N_13369,N_13310);
or U13661 (N_13661,N_13373,N_13446);
and U13662 (N_13662,N_13455,N_13254);
or U13663 (N_13663,N_13283,N_13250);
and U13664 (N_13664,N_13251,N_13313);
and U13665 (N_13665,N_13251,N_13486);
and U13666 (N_13666,N_13386,N_13493);
or U13667 (N_13667,N_13343,N_13453);
or U13668 (N_13668,N_13262,N_13400);
xnor U13669 (N_13669,N_13442,N_13499);
nand U13670 (N_13670,N_13352,N_13257);
and U13671 (N_13671,N_13471,N_13451);
xnor U13672 (N_13672,N_13292,N_13408);
xor U13673 (N_13673,N_13322,N_13346);
xor U13674 (N_13674,N_13349,N_13308);
nor U13675 (N_13675,N_13310,N_13273);
xnor U13676 (N_13676,N_13302,N_13399);
or U13677 (N_13677,N_13416,N_13324);
or U13678 (N_13678,N_13263,N_13271);
nor U13679 (N_13679,N_13393,N_13406);
and U13680 (N_13680,N_13354,N_13471);
xnor U13681 (N_13681,N_13492,N_13353);
or U13682 (N_13682,N_13324,N_13450);
xnor U13683 (N_13683,N_13320,N_13361);
and U13684 (N_13684,N_13390,N_13375);
and U13685 (N_13685,N_13454,N_13377);
nor U13686 (N_13686,N_13448,N_13432);
nand U13687 (N_13687,N_13410,N_13331);
xor U13688 (N_13688,N_13341,N_13491);
nor U13689 (N_13689,N_13460,N_13382);
xor U13690 (N_13690,N_13271,N_13434);
xnor U13691 (N_13691,N_13434,N_13469);
nand U13692 (N_13692,N_13326,N_13417);
xor U13693 (N_13693,N_13370,N_13393);
nor U13694 (N_13694,N_13387,N_13289);
nand U13695 (N_13695,N_13289,N_13320);
nor U13696 (N_13696,N_13274,N_13357);
nand U13697 (N_13697,N_13297,N_13411);
and U13698 (N_13698,N_13386,N_13256);
xor U13699 (N_13699,N_13475,N_13374);
nor U13700 (N_13700,N_13495,N_13386);
nor U13701 (N_13701,N_13382,N_13495);
nand U13702 (N_13702,N_13370,N_13347);
and U13703 (N_13703,N_13289,N_13443);
nand U13704 (N_13704,N_13469,N_13276);
and U13705 (N_13705,N_13258,N_13321);
nor U13706 (N_13706,N_13438,N_13328);
or U13707 (N_13707,N_13293,N_13396);
and U13708 (N_13708,N_13485,N_13397);
and U13709 (N_13709,N_13327,N_13407);
nor U13710 (N_13710,N_13412,N_13401);
or U13711 (N_13711,N_13323,N_13261);
and U13712 (N_13712,N_13298,N_13384);
nor U13713 (N_13713,N_13398,N_13373);
and U13714 (N_13714,N_13412,N_13314);
or U13715 (N_13715,N_13359,N_13250);
xor U13716 (N_13716,N_13254,N_13418);
and U13717 (N_13717,N_13456,N_13421);
nor U13718 (N_13718,N_13350,N_13399);
or U13719 (N_13719,N_13417,N_13328);
or U13720 (N_13720,N_13318,N_13477);
nand U13721 (N_13721,N_13438,N_13258);
nor U13722 (N_13722,N_13455,N_13307);
nand U13723 (N_13723,N_13262,N_13281);
or U13724 (N_13724,N_13304,N_13340);
xnor U13725 (N_13725,N_13445,N_13281);
xor U13726 (N_13726,N_13448,N_13387);
nand U13727 (N_13727,N_13367,N_13417);
nand U13728 (N_13728,N_13488,N_13431);
nand U13729 (N_13729,N_13397,N_13364);
or U13730 (N_13730,N_13383,N_13340);
nand U13731 (N_13731,N_13302,N_13364);
nand U13732 (N_13732,N_13252,N_13267);
and U13733 (N_13733,N_13477,N_13296);
or U13734 (N_13734,N_13335,N_13462);
and U13735 (N_13735,N_13448,N_13401);
or U13736 (N_13736,N_13279,N_13266);
nor U13737 (N_13737,N_13341,N_13404);
nand U13738 (N_13738,N_13311,N_13414);
nand U13739 (N_13739,N_13309,N_13319);
xor U13740 (N_13740,N_13400,N_13439);
and U13741 (N_13741,N_13301,N_13452);
xnor U13742 (N_13742,N_13320,N_13302);
and U13743 (N_13743,N_13349,N_13499);
nor U13744 (N_13744,N_13396,N_13308);
xor U13745 (N_13745,N_13364,N_13470);
xnor U13746 (N_13746,N_13294,N_13276);
nand U13747 (N_13747,N_13336,N_13477);
nand U13748 (N_13748,N_13351,N_13377);
nand U13749 (N_13749,N_13447,N_13302);
or U13750 (N_13750,N_13676,N_13681);
nand U13751 (N_13751,N_13634,N_13533);
nor U13752 (N_13752,N_13667,N_13637);
xor U13753 (N_13753,N_13625,N_13527);
nor U13754 (N_13754,N_13569,N_13671);
xor U13755 (N_13755,N_13571,N_13706);
or U13756 (N_13756,N_13629,N_13564);
xnor U13757 (N_13757,N_13538,N_13719);
and U13758 (N_13758,N_13574,N_13528);
and U13759 (N_13759,N_13611,N_13605);
or U13760 (N_13760,N_13501,N_13714);
or U13761 (N_13761,N_13516,N_13649);
and U13762 (N_13762,N_13641,N_13690);
nand U13763 (N_13763,N_13529,N_13664);
nor U13764 (N_13764,N_13536,N_13698);
nand U13765 (N_13765,N_13545,N_13615);
and U13766 (N_13766,N_13577,N_13651);
and U13767 (N_13767,N_13620,N_13591);
or U13768 (N_13768,N_13653,N_13713);
and U13769 (N_13769,N_13743,N_13601);
nand U13770 (N_13770,N_13708,N_13683);
and U13771 (N_13771,N_13630,N_13650);
xor U13772 (N_13772,N_13524,N_13745);
and U13773 (N_13773,N_13502,N_13525);
xnor U13774 (N_13774,N_13505,N_13703);
nor U13775 (N_13775,N_13731,N_13739);
xor U13776 (N_13776,N_13623,N_13685);
or U13777 (N_13777,N_13515,N_13672);
and U13778 (N_13778,N_13588,N_13663);
xnor U13779 (N_13779,N_13689,N_13619);
nor U13780 (N_13780,N_13682,N_13546);
nand U13781 (N_13781,N_13568,N_13677);
and U13782 (N_13782,N_13679,N_13539);
or U13783 (N_13783,N_13748,N_13554);
xnor U13784 (N_13784,N_13638,N_13707);
nor U13785 (N_13785,N_13666,N_13660);
nor U13786 (N_13786,N_13702,N_13716);
nor U13787 (N_13787,N_13590,N_13612);
and U13788 (N_13788,N_13610,N_13656);
or U13789 (N_13789,N_13730,N_13540);
or U13790 (N_13790,N_13506,N_13626);
or U13791 (N_13791,N_13604,N_13697);
xor U13792 (N_13792,N_13747,N_13556);
or U13793 (N_13793,N_13537,N_13578);
and U13794 (N_13794,N_13674,N_13544);
xnor U13795 (N_13795,N_13511,N_13632);
and U13796 (N_13796,N_13520,N_13737);
nor U13797 (N_13797,N_13652,N_13729);
xnor U13798 (N_13798,N_13642,N_13603);
nand U13799 (N_13799,N_13710,N_13721);
nor U13800 (N_13800,N_13686,N_13639);
nand U13801 (N_13801,N_13742,N_13732);
or U13802 (N_13802,N_13636,N_13648);
nor U13803 (N_13803,N_13513,N_13608);
or U13804 (N_13804,N_13573,N_13728);
or U13805 (N_13805,N_13535,N_13599);
nand U13806 (N_13806,N_13504,N_13635);
nor U13807 (N_13807,N_13675,N_13644);
and U13808 (N_13808,N_13643,N_13680);
xor U13809 (N_13809,N_13518,N_13640);
nor U13810 (N_13810,N_13543,N_13500);
and U13811 (N_13811,N_13662,N_13715);
nand U13812 (N_13812,N_13646,N_13584);
or U13813 (N_13813,N_13657,N_13627);
and U13814 (N_13814,N_13622,N_13665);
nand U13815 (N_13815,N_13744,N_13618);
xnor U13816 (N_13816,N_13613,N_13531);
nand U13817 (N_13817,N_13687,N_13526);
nor U13818 (N_13818,N_13562,N_13631);
or U13819 (N_13819,N_13580,N_13542);
or U13820 (N_13820,N_13594,N_13509);
and U13821 (N_13821,N_13596,N_13583);
nor U13822 (N_13822,N_13624,N_13684);
or U13823 (N_13823,N_13694,N_13550);
xnor U13824 (N_13824,N_13724,N_13733);
xor U13825 (N_13825,N_13517,N_13709);
nor U13826 (N_13826,N_13555,N_13600);
nand U13827 (N_13827,N_13659,N_13606);
or U13828 (N_13828,N_13575,N_13565);
and U13829 (N_13829,N_13589,N_13567);
or U13830 (N_13830,N_13602,N_13586);
nand U13831 (N_13831,N_13532,N_13551);
xor U13832 (N_13832,N_13582,N_13736);
nor U13833 (N_13833,N_13668,N_13616);
and U13834 (N_13834,N_13658,N_13558);
and U13835 (N_13835,N_13579,N_13712);
or U13836 (N_13836,N_13741,N_13701);
or U13837 (N_13837,N_13738,N_13711);
xnor U13838 (N_13838,N_13592,N_13559);
xnor U13839 (N_13839,N_13560,N_13678);
nand U13840 (N_13840,N_13566,N_13521);
or U13841 (N_13841,N_13522,N_13645);
or U13842 (N_13842,N_13749,N_13547);
nand U13843 (N_13843,N_13734,N_13699);
nor U13844 (N_13844,N_13740,N_13688);
and U13845 (N_13845,N_13727,N_13633);
xor U13846 (N_13846,N_13510,N_13726);
nand U13847 (N_13847,N_13507,N_13598);
or U13848 (N_13848,N_13593,N_13695);
nand U13849 (N_13849,N_13587,N_13549);
nor U13850 (N_13850,N_13523,N_13508);
nand U13851 (N_13851,N_13585,N_13735);
nor U13852 (N_13852,N_13621,N_13552);
nor U13853 (N_13853,N_13693,N_13553);
and U13854 (N_13854,N_13717,N_13557);
xnor U13855 (N_13855,N_13617,N_13576);
nor U13856 (N_13856,N_13692,N_13691);
nor U13857 (N_13857,N_13572,N_13595);
xnor U13858 (N_13858,N_13561,N_13581);
or U13859 (N_13859,N_13570,N_13661);
nand U13860 (N_13860,N_13700,N_13548);
nor U13861 (N_13861,N_13512,N_13746);
or U13862 (N_13862,N_13673,N_13530);
nor U13863 (N_13863,N_13514,N_13655);
nor U13864 (N_13864,N_13647,N_13704);
and U13865 (N_13865,N_13519,N_13628);
xor U13866 (N_13866,N_13718,N_13597);
and U13867 (N_13867,N_13541,N_13723);
and U13868 (N_13868,N_13563,N_13669);
nor U13869 (N_13869,N_13534,N_13720);
or U13870 (N_13870,N_13722,N_13725);
or U13871 (N_13871,N_13607,N_13614);
nand U13872 (N_13872,N_13705,N_13696);
and U13873 (N_13873,N_13609,N_13654);
nor U13874 (N_13874,N_13670,N_13503);
xor U13875 (N_13875,N_13639,N_13623);
nand U13876 (N_13876,N_13654,N_13601);
or U13877 (N_13877,N_13586,N_13745);
and U13878 (N_13878,N_13749,N_13551);
nand U13879 (N_13879,N_13709,N_13647);
and U13880 (N_13880,N_13533,N_13506);
or U13881 (N_13881,N_13562,N_13544);
nor U13882 (N_13882,N_13692,N_13602);
or U13883 (N_13883,N_13568,N_13599);
nand U13884 (N_13884,N_13651,N_13684);
or U13885 (N_13885,N_13647,N_13731);
xnor U13886 (N_13886,N_13537,N_13568);
xnor U13887 (N_13887,N_13743,N_13630);
nand U13888 (N_13888,N_13714,N_13674);
nor U13889 (N_13889,N_13595,N_13541);
or U13890 (N_13890,N_13651,N_13593);
and U13891 (N_13891,N_13632,N_13712);
nand U13892 (N_13892,N_13656,N_13620);
nor U13893 (N_13893,N_13522,N_13585);
xnor U13894 (N_13894,N_13620,N_13650);
xnor U13895 (N_13895,N_13738,N_13644);
nand U13896 (N_13896,N_13736,N_13738);
xor U13897 (N_13897,N_13677,N_13577);
nand U13898 (N_13898,N_13597,N_13660);
nand U13899 (N_13899,N_13568,N_13574);
and U13900 (N_13900,N_13681,N_13705);
or U13901 (N_13901,N_13524,N_13634);
and U13902 (N_13902,N_13626,N_13603);
nor U13903 (N_13903,N_13725,N_13521);
and U13904 (N_13904,N_13746,N_13619);
nand U13905 (N_13905,N_13683,N_13550);
or U13906 (N_13906,N_13741,N_13588);
xnor U13907 (N_13907,N_13549,N_13712);
xnor U13908 (N_13908,N_13729,N_13661);
nor U13909 (N_13909,N_13688,N_13731);
and U13910 (N_13910,N_13685,N_13733);
and U13911 (N_13911,N_13565,N_13627);
xnor U13912 (N_13912,N_13706,N_13708);
and U13913 (N_13913,N_13537,N_13540);
and U13914 (N_13914,N_13540,N_13635);
and U13915 (N_13915,N_13657,N_13720);
or U13916 (N_13916,N_13576,N_13742);
xnor U13917 (N_13917,N_13636,N_13719);
and U13918 (N_13918,N_13683,N_13692);
xor U13919 (N_13919,N_13550,N_13628);
xnor U13920 (N_13920,N_13505,N_13515);
or U13921 (N_13921,N_13533,N_13512);
and U13922 (N_13922,N_13652,N_13714);
and U13923 (N_13923,N_13559,N_13689);
nand U13924 (N_13924,N_13735,N_13667);
or U13925 (N_13925,N_13683,N_13535);
and U13926 (N_13926,N_13550,N_13546);
and U13927 (N_13927,N_13600,N_13711);
or U13928 (N_13928,N_13571,N_13529);
nor U13929 (N_13929,N_13646,N_13674);
or U13930 (N_13930,N_13710,N_13658);
or U13931 (N_13931,N_13636,N_13747);
and U13932 (N_13932,N_13613,N_13608);
xor U13933 (N_13933,N_13501,N_13587);
and U13934 (N_13934,N_13722,N_13519);
nand U13935 (N_13935,N_13620,N_13607);
or U13936 (N_13936,N_13557,N_13661);
nor U13937 (N_13937,N_13731,N_13704);
nand U13938 (N_13938,N_13651,N_13695);
nand U13939 (N_13939,N_13712,N_13556);
and U13940 (N_13940,N_13735,N_13611);
nor U13941 (N_13941,N_13508,N_13614);
and U13942 (N_13942,N_13696,N_13604);
nor U13943 (N_13943,N_13542,N_13623);
or U13944 (N_13944,N_13611,N_13543);
nand U13945 (N_13945,N_13569,N_13617);
nand U13946 (N_13946,N_13538,N_13558);
nor U13947 (N_13947,N_13686,N_13681);
xnor U13948 (N_13948,N_13724,N_13629);
xor U13949 (N_13949,N_13580,N_13746);
nor U13950 (N_13950,N_13575,N_13631);
and U13951 (N_13951,N_13574,N_13611);
nand U13952 (N_13952,N_13625,N_13733);
and U13953 (N_13953,N_13734,N_13595);
nor U13954 (N_13954,N_13696,N_13625);
and U13955 (N_13955,N_13707,N_13611);
and U13956 (N_13956,N_13502,N_13529);
nor U13957 (N_13957,N_13581,N_13652);
or U13958 (N_13958,N_13702,N_13672);
nor U13959 (N_13959,N_13676,N_13593);
and U13960 (N_13960,N_13538,N_13720);
xor U13961 (N_13961,N_13607,N_13691);
or U13962 (N_13962,N_13717,N_13502);
nor U13963 (N_13963,N_13706,N_13527);
nand U13964 (N_13964,N_13654,N_13556);
nand U13965 (N_13965,N_13514,N_13530);
and U13966 (N_13966,N_13619,N_13507);
xnor U13967 (N_13967,N_13569,N_13705);
xor U13968 (N_13968,N_13687,N_13678);
and U13969 (N_13969,N_13728,N_13632);
nand U13970 (N_13970,N_13589,N_13647);
and U13971 (N_13971,N_13699,N_13523);
or U13972 (N_13972,N_13691,N_13728);
xor U13973 (N_13973,N_13723,N_13613);
nor U13974 (N_13974,N_13587,N_13554);
nor U13975 (N_13975,N_13643,N_13679);
or U13976 (N_13976,N_13683,N_13548);
nor U13977 (N_13977,N_13510,N_13730);
or U13978 (N_13978,N_13539,N_13515);
and U13979 (N_13979,N_13527,N_13590);
and U13980 (N_13980,N_13666,N_13682);
nand U13981 (N_13981,N_13595,N_13547);
nor U13982 (N_13982,N_13597,N_13646);
and U13983 (N_13983,N_13554,N_13651);
and U13984 (N_13984,N_13561,N_13502);
and U13985 (N_13985,N_13547,N_13611);
nand U13986 (N_13986,N_13514,N_13526);
nand U13987 (N_13987,N_13518,N_13689);
and U13988 (N_13988,N_13546,N_13595);
nand U13989 (N_13989,N_13697,N_13647);
or U13990 (N_13990,N_13516,N_13622);
or U13991 (N_13991,N_13708,N_13550);
and U13992 (N_13992,N_13727,N_13604);
xor U13993 (N_13993,N_13723,N_13542);
or U13994 (N_13994,N_13551,N_13592);
nor U13995 (N_13995,N_13654,N_13575);
nor U13996 (N_13996,N_13536,N_13523);
and U13997 (N_13997,N_13748,N_13649);
and U13998 (N_13998,N_13742,N_13655);
nand U13999 (N_13999,N_13512,N_13737);
xor U14000 (N_14000,N_13908,N_13833);
or U14001 (N_14001,N_13896,N_13816);
nand U14002 (N_14002,N_13809,N_13890);
or U14003 (N_14003,N_13814,N_13933);
or U14004 (N_14004,N_13857,N_13870);
xor U14005 (N_14005,N_13980,N_13787);
xor U14006 (N_14006,N_13970,N_13851);
nor U14007 (N_14007,N_13947,N_13768);
and U14008 (N_14008,N_13967,N_13826);
xnor U14009 (N_14009,N_13957,N_13847);
nor U14010 (N_14010,N_13776,N_13966);
nand U14011 (N_14011,N_13825,N_13765);
and U14012 (N_14012,N_13859,N_13984);
or U14013 (N_14013,N_13839,N_13855);
nor U14014 (N_14014,N_13894,N_13937);
nand U14015 (N_14015,N_13779,N_13892);
xor U14016 (N_14016,N_13829,N_13899);
nor U14017 (N_14017,N_13963,N_13797);
or U14018 (N_14018,N_13864,N_13803);
and U14019 (N_14019,N_13844,N_13819);
nor U14020 (N_14020,N_13856,N_13930);
nand U14021 (N_14021,N_13869,N_13988);
nand U14022 (N_14022,N_13960,N_13999);
and U14023 (N_14023,N_13822,N_13961);
or U14024 (N_14024,N_13794,N_13753);
xor U14025 (N_14025,N_13882,N_13848);
nand U14026 (N_14026,N_13982,N_13951);
and U14027 (N_14027,N_13813,N_13811);
or U14028 (N_14028,N_13893,N_13981);
and U14029 (N_14029,N_13771,N_13830);
and U14030 (N_14030,N_13790,N_13846);
and U14031 (N_14031,N_13889,N_13751);
xor U14032 (N_14032,N_13940,N_13943);
nand U14033 (N_14033,N_13928,N_13777);
xnor U14034 (N_14034,N_13913,N_13840);
xnor U14035 (N_14035,N_13903,N_13979);
nand U14036 (N_14036,N_13885,N_13878);
or U14037 (N_14037,N_13824,N_13769);
nand U14038 (N_14038,N_13843,N_13959);
xor U14039 (N_14039,N_13998,N_13788);
nor U14040 (N_14040,N_13868,N_13918);
xor U14041 (N_14041,N_13949,N_13810);
and U14042 (N_14042,N_13860,N_13887);
xor U14043 (N_14043,N_13983,N_13879);
or U14044 (N_14044,N_13798,N_13997);
and U14045 (N_14045,N_13919,N_13770);
nor U14046 (N_14046,N_13883,N_13783);
nand U14047 (N_14047,N_13977,N_13911);
nand U14048 (N_14048,N_13954,N_13761);
or U14049 (N_14049,N_13898,N_13774);
nand U14050 (N_14050,N_13952,N_13762);
nand U14051 (N_14051,N_13827,N_13866);
nand U14052 (N_14052,N_13756,N_13752);
xor U14053 (N_14053,N_13853,N_13804);
nor U14054 (N_14054,N_13845,N_13796);
xnor U14055 (N_14055,N_13948,N_13755);
nand U14056 (N_14056,N_13793,N_13912);
or U14057 (N_14057,N_13985,N_13917);
nand U14058 (N_14058,N_13759,N_13852);
xnor U14059 (N_14059,N_13766,N_13950);
or U14060 (N_14060,N_13791,N_13897);
or U14061 (N_14061,N_13964,N_13925);
xor U14062 (N_14062,N_13750,N_13995);
xnor U14063 (N_14063,N_13993,N_13936);
nor U14064 (N_14064,N_13915,N_13962);
nand U14065 (N_14065,N_13781,N_13900);
nor U14066 (N_14066,N_13921,N_13895);
or U14067 (N_14067,N_13877,N_13975);
nor U14068 (N_14068,N_13976,N_13806);
xor U14069 (N_14069,N_13946,N_13764);
and U14070 (N_14070,N_13935,N_13812);
nand U14071 (N_14071,N_13758,N_13942);
nand U14072 (N_14072,N_13832,N_13801);
or U14073 (N_14073,N_13923,N_13994);
nor U14074 (N_14074,N_13974,N_13888);
nor U14075 (N_14075,N_13862,N_13969);
and U14076 (N_14076,N_13795,N_13958);
or U14077 (N_14077,N_13991,N_13775);
nand U14078 (N_14078,N_13865,N_13934);
nor U14079 (N_14079,N_13757,N_13876);
nor U14080 (N_14080,N_13867,N_13820);
nand U14081 (N_14081,N_13910,N_13973);
nand U14082 (N_14082,N_13754,N_13772);
xor U14083 (N_14083,N_13802,N_13807);
nand U14084 (N_14084,N_13786,N_13835);
and U14085 (N_14085,N_13834,N_13875);
xor U14086 (N_14086,N_13792,N_13861);
nor U14087 (N_14087,N_13858,N_13907);
nor U14088 (N_14088,N_13902,N_13837);
nand U14089 (N_14089,N_13996,N_13909);
or U14090 (N_14090,N_13784,N_13987);
xor U14091 (N_14091,N_13905,N_13941);
nor U14092 (N_14092,N_13955,N_13965);
xor U14093 (N_14093,N_13817,N_13799);
and U14094 (N_14094,N_13990,N_13939);
nor U14095 (N_14095,N_13916,N_13838);
and U14096 (N_14096,N_13818,N_13836);
or U14097 (N_14097,N_13849,N_13920);
or U14098 (N_14098,N_13821,N_13901);
and U14099 (N_14099,N_13926,N_13854);
nor U14100 (N_14100,N_13767,N_13914);
xnor U14101 (N_14101,N_13815,N_13789);
xnor U14102 (N_14102,N_13906,N_13904);
and U14103 (N_14103,N_13872,N_13881);
xor U14104 (N_14104,N_13932,N_13891);
or U14105 (N_14105,N_13808,N_13805);
or U14106 (N_14106,N_13831,N_13778);
or U14107 (N_14107,N_13863,N_13972);
nor U14108 (N_14108,N_13924,N_13968);
nor U14109 (N_14109,N_13823,N_13800);
and U14110 (N_14110,N_13938,N_13773);
nand U14111 (N_14111,N_13944,N_13956);
nand U14112 (N_14112,N_13927,N_13884);
or U14113 (N_14113,N_13841,N_13986);
and U14114 (N_14114,N_13953,N_13871);
or U14115 (N_14115,N_13931,N_13850);
xor U14116 (N_14116,N_13886,N_13978);
xor U14117 (N_14117,N_13873,N_13780);
and U14118 (N_14118,N_13989,N_13828);
xor U14119 (N_14119,N_13992,N_13971);
or U14120 (N_14120,N_13880,N_13929);
or U14121 (N_14121,N_13763,N_13760);
or U14122 (N_14122,N_13842,N_13922);
nor U14123 (N_14123,N_13945,N_13782);
or U14124 (N_14124,N_13785,N_13874);
xnor U14125 (N_14125,N_13968,N_13761);
xnor U14126 (N_14126,N_13889,N_13899);
xnor U14127 (N_14127,N_13772,N_13830);
xnor U14128 (N_14128,N_13859,N_13902);
nand U14129 (N_14129,N_13799,N_13838);
nand U14130 (N_14130,N_13813,N_13880);
and U14131 (N_14131,N_13760,N_13890);
and U14132 (N_14132,N_13773,N_13970);
nand U14133 (N_14133,N_13924,N_13943);
nor U14134 (N_14134,N_13833,N_13951);
and U14135 (N_14135,N_13850,N_13959);
and U14136 (N_14136,N_13801,N_13783);
xnor U14137 (N_14137,N_13888,N_13993);
and U14138 (N_14138,N_13914,N_13821);
and U14139 (N_14139,N_13753,N_13907);
xor U14140 (N_14140,N_13864,N_13939);
and U14141 (N_14141,N_13876,N_13768);
or U14142 (N_14142,N_13830,N_13785);
or U14143 (N_14143,N_13844,N_13969);
or U14144 (N_14144,N_13783,N_13788);
xor U14145 (N_14145,N_13809,N_13916);
nor U14146 (N_14146,N_13987,N_13861);
nand U14147 (N_14147,N_13905,N_13854);
xor U14148 (N_14148,N_13976,N_13907);
nand U14149 (N_14149,N_13984,N_13974);
or U14150 (N_14150,N_13803,N_13900);
nor U14151 (N_14151,N_13793,N_13990);
or U14152 (N_14152,N_13785,N_13764);
xor U14153 (N_14153,N_13756,N_13997);
or U14154 (N_14154,N_13993,N_13834);
or U14155 (N_14155,N_13992,N_13886);
and U14156 (N_14156,N_13891,N_13950);
xor U14157 (N_14157,N_13868,N_13782);
nand U14158 (N_14158,N_13867,N_13767);
xnor U14159 (N_14159,N_13796,N_13957);
and U14160 (N_14160,N_13800,N_13994);
and U14161 (N_14161,N_13897,N_13987);
nor U14162 (N_14162,N_13873,N_13834);
nand U14163 (N_14163,N_13917,N_13821);
xnor U14164 (N_14164,N_13949,N_13876);
nand U14165 (N_14165,N_13914,N_13864);
or U14166 (N_14166,N_13827,N_13831);
nor U14167 (N_14167,N_13834,N_13889);
or U14168 (N_14168,N_13774,N_13757);
nor U14169 (N_14169,N_13791,N_13920);
nand U14170 (N_14170,N_13819,N_13803);
or U14171 (N_14171,N_13962,N_13936);
or U14172 (N_14172,N_13850,N_13798);
and U14173 (N_14173,N_13889,N_13987);
nor U14174 (N_14174,N_13782,N_13760);
xor U14175 (N_14175,N_13883,N_13906);
and U14176 (N_14176,N_13796,N_13897);
xnor U14177 (N_14177,N_13928,N_13972);
nand U14178 (N_14178,N_13778,N_13817);
nor U14179 (N_14179,N_13918,N_13938);
nor U14180 (N_14180,N_13781,N_13858);
nand U14181 (N_14181,N_13967,N_13924);
nor U14182 (N_14182,N_13915,N_13908);
nor U14183 (N_14183,N_13803,N_13784);
and U14184 (N_14184,N_13869,N_13864);
nor U14185 (N_14185,N_13941,N_13807);
or U14186 (N_14186,N_13955,N_13768);
or U14187 (N_14187,N_13992,N_13972);
nor U14188 (N_14188,N_13935,N_13810);
nor U14189 (N_14189,N_13864,N_13855);
nor U14190 (N_14190,N_13825,N_13936);
and U14191 (N_14191,N_13944,N_13959);
nor U14192 (N_14192,N_13940,N_13835);
and U14193 (N_14193,N_13774,N_13900);
and U14194 (N_14194,N_13929,N_13987);
xnor U14195 (N_14195,N_13916,N_13792);
and U14196 (N_14196,N_13773,N_13933);
or U14197 (N_14197,N_13836,N_13817);
nor U14198 (N_14198,N_13915,N_13924);
nor U14199 (N_14199,N_13980,N_13772);
nand U14200 (N_14200,N_13917,N_13991);
nor U14201 (N_14201,N_13924,N_13963);
or U14202 (N_14202,N_13957,N_13868);
or U14203 (N_14203,N_13964,N_13896);
or U14204 (N_14204,N_13868,N_13916);
nor U14205 (N_14205,N_13979,N_13779);
xor U14206 (N_14206,N_13766,N_13917);
or U14207 (N_14207,N_13768,N_13851);
xor U14208 (N_14208,N_13948,N_13783);
or U14209 (N_14209,N_13973,N_13935);
or U14210 (N_14210,N_13891,N_13783);
nand U14211 (N_14211,N_13923,N_13840);
nand U14212 (N_14212,N_13780,N_13852);
nand U14213 (N_14213,N_13875,N_13924);
and U14214 (N_14214,N_13793,N_13816);
and U14215 (N_14215,N_13956,N_13911);
nand U14216 (N_14216,N_13946,N_13962);
and U14217 (N_14217,N_13763,N_13794);
or U14218 (N_14218,N_13870,N_13848);
nor U14219 (N_14219,N_13916,N_13835);
nor U14220 (N_14220,N_13925,N_13784);
xnor U14221 (N_14221,N_13847,N_13960);
xnor U14222 (N_14222,N_13790,N_13813);
or U14223 (N_14223,N_13839,N_13798);
xnor U14224 (N_14224,N_13961,N_13824);
nor U14225 (N_14225,N_13783,N_13833);
nor U14226 (N_14226,N_13932,N_13955);
xor U14227 (N_14227,N_13773,N_13824);
or U14228 (N_14228,N_13775,N_13835);
and U14229 (N_14229,N_13941,N_13792);
xor U14230 (N_14230,N_13799,N_13913);
xnor U14231 (N_14231,N_13948,N_13965);
xnor U14232 (N_14232,N_13838,N_13781);
or U14233 (N_14233,N_13776,N_13761);
nor U14234 (N_14234,N_13895,N_13754);
xnor U14235 (N_14235,N_13867,N_13976);
nor U14236 (N_14236,N_13926,N_13952);
nand U14237 (N_14237,N_13788,N_13982);
xor U14238 (N_14238,N_13878,N_13890);
xor U14239 (N_14239,N_13851,N_13869);
xnor U14240 (N_14240,N_13849,N_13976);
nor U14241 (N_14241,N_13817,N_13954);
nor U14242 (N_14242,N_13774,N_13986);
or U14243 (N_14243,N_13918,N_13904);
or U14244 (N_14244,N_13857,N_13935);
nor U14245 (N_14245,N_13843,N_13878);
or U14246 (N_14246,N_13998,N_13946);
or U14247 (N_14247,N_13764,N_13788);
and U14248 (N_14248,N_13807,N_13798);
and U14249 (N_14249,N_13812,N_13945);
or U14250 (N_14250,N_14137,N_14119);
and U14251 (N_14251,N_14231,N_14094);
nor U14252 (N_14252,N_14025,N_14178);
nand U14253 (N_14253,N_14187,N_14040);
nor U14254 (N_14254,N_14246,N_14076);
nor U14255 (N_14255,N_14073,N_14026);
or U14256 (N_14256,N_14120,N_14087);
and U14257 (N_14257,N_14111,N_14049);
or U14258 (N_14258,N_14156,N_14125);
and U14259 (N_14259,N_14192,N_14248);
xor U14260 (N_14260,N_14036,N_14038);
xnor U14261 (N_14261,N_14140,N_14199);
nand U14262 (N_14262,N_14244,N_14173);
and U14263 (N_14263,N_14210,N_14202);
nor U14264 (N_14264,N_14037,N_14032);
nor U14265 (N_14265,N_14136,N_14109);
nor U14266 (N_14266,N_14006,N_14091);
xor U14267 (N_14267,N_14127,N_14013);
nor U14268 (N_14268,N_14208,N_14090);
or U14269 (N_14269,N_14216,N_14180);
nor U14270 (N_14270,N_14072,N_14234);
nand U14271 (N_14271,N_14242,N_14001);
nor U14272 (N_14272,N_14068,N_14190);
nand U14273 (N_14273,N_14238,N_14078);
nand U14274 (N_14274,N_14205,N_14217);
nor U14275 (N_14275,N_14058,N_14245);
xor U14276 (N_14276,N_14074,N_14154);
xnor U14277 (N_14277,N_14128,N_14243);
nand U14278 (N_14278,N_14066,N_14077);
and U14279 (N_14279,N_14207,N_14130);
and U14280 (N_14280,N_14169,N_14027);
and U14281 (N_14281,N_14174,N_14124);
or U14282 (N_14282,N_14197,N_14041);
xor U14283 (N_14283,N_14166,N_14113);
xor U14284 (N_14284,N_14144,N_14224);
xor U14285 (N_14285,N_14200,N_14241);
and U14286 (N_14286,N_14053,N_14134);
nand U14287 (N_14287,N_14062,N_14050);
nor U14288 (N_14288,N_14171,N_14141);
or U14289 (N_14289,N_14160,N_14064);
xor U14290 (N_14290,N_14002,N_14017);
nand U14291 (N_14291,N_14034,N_14181);
and U14292 (N_14292,N_14143,N_14146);
xnor U14293 (N_14293,N_14220,N_14020);
nor U14294 (N_14294,N_14148,N_14235);
and U14295 (N_14295,N_14196,N_14188);
xor U14296 (N_14296,N_14043,N_14110);
and U14297 (N_14297,N_14047,N_14007);
nor U14298 (N_14298,N_14052,N_14195);
or U14299 (N_14299,N_14218,N_14240);
nor U14300 (N_14300,N_14162,N_14182);
or U14301 (N_14301,N_14067,N_14044);
and U14302 (N_14302,N_14211,N_14164);
and U14303 (N_14303,N_14232,N_14086);
nand U14304 (N_14304,N_14048,N_14168);
nor U14305 (N_14305,N_14114,N_14206);
or U14306 (N_14306,N_14215,N_14228);
xnor U14307 (N_14307,N_14029,N_14161);
xor U14308 (N_14308,N_14147,N_14219);
nor U14309 (N_14309,N_14225,N_14230);
nand U14310 (N_14310,N_14193,N_14236);
and U14311 (N_14311,N_14172,N_14088);
nand U14312 (N_14312,N_14028,N_14033);
xnor U14313 (N_14313,N_14183,N_14070);
or U14314 (N_14314,N_14203,N_14097);
nand U14315 (N_14315,N_14080,N_14159);
or U14316 (N_14316,N_14055,N_14079);
nand U14317 (N_14317,N_14155,N_14008);
nand U14318 (N_14318,N_14054,N_14084);
and U14319 (N_14319,N_14004,N_14065);
and U14320 (N_14320,N_14011,N_14118);
or U14321 (N_14321,N_14151,N_14158);
nor U14322 (N_14322,N_14117,N_14142);
and U14323 (N_14323,N_14209,N_14045);
or U14324 (N_14324,N_14022,N_14138);
or U14325 (N_14325,N_14247,N_14081);
or U14326 (N_14326,N_14061,N_14106);
and U14327 (N_14327,N_14249,N_14108);
or U14328 (N_14328,N_14176,N_14095);
and U14329 (N_14329,N_14018,N_14170);
or U14330 (N_14330,N_14129,N_14239);
or U14331 (N_14331,N_14194,N_14057);
xnor U14332 (N_14332,N_14213,N_14112);
nor U14333 (N_14333,N_14139,N_14093);
or U14334 (N_14334,N_14085,N_14191);
nand U14335 (N_14335,N_14101,N_14145);
or U14336 (N_14336,N_14123,N_14126);
or U14337 (N_14337,N_14009,N_14019);
and U14338 (N_14338,N_14131,N_14104);
or U14339 (N_14339,N_14082,N_14179);
and U14340 (N_14340,N_14184,N_14021);
and U14341 (N_14341,N_14000,N_14030);
nor U14342 (N_14342,N_14157,N_14115);
xnor U14343 (N_14343,N_14237,N_14003);
or U14344 (N_14344,N_14063,N_14185);
nor U14345 (N_14345,N_14233,N_14089);
xnor U14346 (N_14346,N_14177,N_14201);
and U14347 (N_14347,N_14102,N_14152);
or U14348 (N_14348,N_14149,N_14132);
nor U14349 (N_14349,N_14105,N_14024);
nand U14350 (N_14350,N_14098,N_14214);
nor U14351 (N_14351,N_14186,N_14229);
and U14352 (N_14352,N_14226,N_14103);
nor U14353 (N_14353,N_14167,N_14222);
nor U14354 (N_14354,N_14122,N_14204);
nand U14355 (N_14355,N_14056,N_14133);
or U14356 (N_14356,N_14012,N_14010);
and U14357 (N_14357,N_14060,N_14031);
nor U14358 (N_14358,N_14016,N_14121);
or U14359 (N_14359,N_14035,N_14083);
nor U14360 (N_14360,N_14189,N_14135);
or U14361 (N_14361,N_14165,N_14075);
or U14362 (N_14362,N_14071,N_14175);
or U14363 (N_14363,N_14092,N_14005);
nor U14364 (N_14364,N_14015,N_14051);
or U14365 (N_14365,N_14223,N_14163);
xor U14366 (N_14366,N_14059,N_14221);
xor U14367 (N_14367,N_14046,N_14014);
xnor U14368 (N_14368,N_14107,N_14212);
and U14369 (N_14369,N_14099,N_14227);
nor U14370 (N_14370,N_14069,N_14153);
nand U14371 (N_14371,N_14150,N_14116);
nand U14372 (N_14372,N_14039,N_14100);
nand U14373 (N_14373,N_14042,N_14096);
and U14374 (N_14374,N_14198,N_14023);
and U14375 (N_14375,N_14068,N_14049);
or U14376 (N_14376,N_14047,N_14091);
nand U14377 (N_14377,N_14242,N_14061);
and U14378 (N_14378,N_14068,N_14088);
or U14379 (N_14379,N_14001,N_14170);
xor U14380 (N_14380,N_14015,N_14171);
nor U14381 (N_14381,N_14028,N_14177);
xnor U14382 (N_14382,N_14215,N_14089);
xor U14383 (N_14383,N_14092,N_14001);
or U14384 (N_14384,N_14001,N_14237);
or U14385 (N_14385,N_14194,N_14222);
nor U14386 (N_14386,N_14016,N_14028);
nand U14387 (N_14387,N_14197,N_14232);
xnor U14388 (N_14388,N_14138,N_14136);
xnor U14389 (N_14389,N_14096,N_14072);
nand U14390 (N_14390,N_14222,N_14161);
and U14391 (N_14391,N_14235,N_14134);
nor U14392 (N_14392,N_14011,N_14184);
and U14393 (N_14393,N_14004,N_14165);
xnor U14394 (N_14394,N_14088,N_14222);
or U14395 (N_14395,N_14101,N_14015);
nand U14396 (N_14396,N_14173,N_14010);
or U14397 (N_14397,N_14115,N_14214);
nand U14398 (N_14398,N_14210,N_14058);
or U14399 (N_14399,N_14156,N_14131);
or U14400 (N_14400,N_14052,N_14147);
nor U14401 (N_14401,N_14071,N_14003);
or U14402 (N_14402,N_14056,N_14093);
nor U14403 (N_14403,N_14170,N_14233);
and U14404 (N_14404,N_14157,N_14215);
nor U14405 (N_14405,N_14076,N_14020);
nor U14406 (N_14406,N_14018,N_14171);
nor U14407 (N_14407,N_14161,N_14005);
xor U14408 (N_14408,N_14057,N_14154);
nand U14409 (N_14409,N_14069,N_14162);
and U14410 (N_14410,N_14132,N_14117);
xor U14411 (N_14411,N_14130,N_14223);
nand U14412 (N_14412,N_14160,N_14129);
or U14413 (N_14413,N_14227,N_14212);
nand U14414 (N_14414,N_14246,N_14227);
xor U14415 (N_14415,N_14215,N_14003);
nand U14416 (N_14416,N_14108,N_14101);
xnor U14417 (N_14417,N_14219,N_14029);
and U14418 (N_14418,N_14087,N_14243);
or U14419 (N_14419,N_14242,N_14238);
or U14420 (N_14420,N_14019,N_14068);
nand U14421 (N_14421,N_14106,N_14010);
nand U14422 (N_14422,N_14025,N_14120);
and U14423 (N_14423,N_14107,N_14169);
nand U14424 (N_14424,N_14078,N_14069);
xnor U14425 (N_14425,N_14003,N_14063);
nand U14426 (N_14426,N_14204,N_14032);
and U14427 (N_14427,N_14055,N_14108);
or U14428 (N_14428,N_14132,N_14180);
nor U14429 (N_14429,N_14111,N_14150);
xnor U14430 (N_14430,N_14195,N_14222);
nand U14431 (N_14431,N_14133,N_14184);
xnor U14432 (N_14432,N_14172,N_14241);
xnor U14433 (N_14433,N_14151,N_14111);
xor U14434 (N_14434,N_14026,N_14012);
nor U14435 (N_14435,N_14170,N_14210);
and U14436 (N_14436,N_14162,N_14220);
or U14437 (N_14437,N_14006,N_14123);
xor U14438 (N_14438,N_14086,N_14183);
xnor U14439 (N_14439,N_14096,N_14100);
nand U14440 (N_14440,N_14101,N_14234);
nor U14441 (N_14441,N_14008,N_14003);
xor U14442 (N_14442,N_14083,N_14185);
xnor U14443 (N_14443,N_14164,N_14223);
xnor U14444 (N_14444,N_14246,N_14078);
nor U14445 (N_14445,N_14098,N_14216);
nand U14446 (N_14446,N_14064,N_14050);
and U14447 (N_14447,N_14249,N_14098);
and U14448 (N_14448,N_14058,N_14157);
nor U14449 (N_14449,N_14210,N_14165);
nor U14450 (N_14450,N_14153,N_14015);
xnor U14451 (N_14451,N_14218,N_14169);
nor U14452 (N_14452,N_14225,N_14062);
nor U14453 (N_14453,N_14219,N_14092);
xor U14454 (N_14454,N_14102,N_14122);
xnor U14455 (N_14455,N_14180,N_14231);
and U14456 (N_14456,N_14188,N_14244);
or U14457 (N_14457,N_14234,N_14196);
or U14458 (N_14458,N_14046,N_14164);
nor U14459 (N_14459,N_14249,N_14095);
and U14460 (N_14460,N_14050,N_14216);
and U14461 (N_14461,N_14142,N_14122);
xnor U14462 (N_14462,N_14132,N_14115);
nor U14463 (N_14463,N_14175,N_14111);
xor U14464 (N_14464,N_14217,N_14082);
xnor U14465 (N_14465,N_14100,N_14193);
and U14466 (N_14466,N_14027,N_14064);
and U14467 (N_14467,N_14161,N_14247);
xor U14468 (N_14468,N_14204,N_14097);
and U14469 (N_14469,N_14061,N_14180);
xor U14470 (N_14470,N_14238,N_14140);
nand U14471 (N_14471,N_14228,N_14003);
nand U14472 (N_14472,N_14084,N_14201);
or U14473 (N_14473,N_14172,N_14099);
nand U14474 (N_14474,N_14174,N_14201);
xnor U14475 (N_14475,N_14229,N_14193);
nor U14476 (N_14476,N_14245,N_14225);
nor U14477 (N_14477,N_14027,N_14129);
nor U14478 (N_14478,N_14022,N_14160);
and U14479 (N_14479,N_14166,N_14199);
and U14480 (N_14480,N_14238,N_14209);
and U14481 (N_14481,N_14106,N_14189);
or U14482 (N_14482,N_14139,N_14228);
or U14483 (N_14483,N_14200,N_14234);
nand U14484 (N_14484,N_14228,N_14037);
or U14485 (N_14485,N_14132,N_14130);
and U14486 (N_14486,N_14129,N_14113);
nor U14487 (N_14487,N_14018,N_14130);
xnor U14488 (N_14488,N_14105,N_14041);
nand U14489 (N_14489,N_14059,N_14169);
nand U14490 (N_14490,N_14052,N_14108);
or U14491 (N_14491,N_14095,N_14089);
nand U14492 (N_14492,N_14101,N_14215);
nand U14493 (N_14493,N_14074,N_14009);
nor U14494 (N_14494,N_14012,N_14171);
nand U14495 (N_14495,N_14047,N_14055);
and U14496 (N_14496,N_14057,N_14216);
xor U14497 (N_14497,N_14249,N_14133);
nor U14498 (N_14498,N_14172,N_14131);
nor U14499 (N_14499,N_14170,N_14123);
nor U14500 (N_14500,N_14292,N_14414);
xnor U14501 (N_14501,N_14296,N_14473);
nand U14502 (N_14502,N_14453,N_14260);
or U14503 (N_14503,N_14488,N_14395);
or U14504 (N_14504,N_14428,N_14424);
nor U14505 (N_14505,N_14437,N_14382);
xor U14506 (N_14506,N_14407,N_14299);
or U14507 (N_14507,N_14376,N_14405);
nor U14508 (N_14508,N_14363,N_14494);
or U14509 (N_14509,N_14457,N_14496);
nor U14510 (N_14510,N_14479,N_14338);
nand U14511 (N_14511,N_14469,N_14259);
nor U14512 (N_14512,N_14321,N_14442);
or U14513 (N_14513,N_14410,N_14438);
and U14514 (N_14514,N_14358,N_14446);
and U14515 (N_14515,N_14398,N_14319);
nand U14516 (N_14516,N_14477,N_14250);
or U14517 (N_14517,N_14380,N_14465);
xnor U14518 (N_14518,N_14409,N_14336);
and U14519 (N_14519,N_14432,N_14288);
nor U14520 (N_14520,N_14289,N_14255);
nor U14521 (N_14521,N_14345,N_14396);
and U14522 (N_14522,N_14433,N_14331);
and U14523 (N_14523,N_14458,N_14316);
and U14524 (N_14524,N_14378,N_14417);
and U14525 (N_14525,N_14310,N_14328);
or U14526 (N_14526,N_14337,N_14371);
nand U14527 (N_14527,N_14252,N_14377);
xnor U14528 (N_14528,N_14273,N_14370);
xor U14529 (N_14529,N_14305,N_14295);
or U14530 (N_14530,N_14491,N_14450);
or U14531 (N_14531,N_14297,N_14468);
xor U14532 (N_14532,N_14434,N_14429);
or U14533 (N_14533,N_14350,N_14286);
or U14534 (N_14534,N_14493,N_14430);
nand U14535 (N_14535,N_14394,N_14412);
nand U14536 (N_14536,N_14352,N_14492);
or U14537 (N_14537,N_14304,N_14478);
nand U14538 (N_14538,N_14443,N_14413);
and U14539 (N_14539,N_14423,N_14283);
xor U14540 (N_14540,N_14384,N_14421);
nor U14541 (N_14541,N_14256,N_14268);
nor U14542 (N_14542,N_14324,N_14356);
nand U14543 (N_14543,N_14274,N_14373);
xnor U14544 (N_14544,N_14451,N_14386);
or U14545 (N_14545,N_14461,N_14426);
nand U14546 (N_14546,N_14422,N_14333);
xnor U14547 (N_14547,N_14475,N_14464);
and U14548 (N_14548,N_14339,N_14460);
and U14549 (N_14549,N_14416,N_14303);
xor U14550 (N_14550,N_14367,N_14311);
and U14551 (N_14551,N_14301,N_14397);
xnor U14552 (N_14552,N_14489,N_14449);
or U14553 (N_14553,N_14462,N_14399);
nand U14554 (N_14554,N_14309,N_14404);
nand U14555 (N_14555,N_14360,N_14271);
nand U14556 (N_14556,N_14452,N_14330);
and U14557 (N_14557,N_14466,N_14406);
or U14558 (N_14558,N_14480,N_14393);
nand U14559 (N_14559,N_14281,N_14392);
nor U14560 (N_14560,N_14359,N_14419);
and U14561 (N_14561,N_14364,N_14354);
nand U14562 (N_14562,N_14278,N_14298);
nand U14563 (N_14563,N_14342,N_14455);
and U14564 (N_14564,N_14253,N_14411);
nor U14565 (N_14565,N_14490,N_14314);
xor U14566 (N_14566,N_14318,N_14420);
nand U14567 (N_14567,N_14361,N_14302);
or U14568 (N_14568,N_14445,N_14385);
or U14569 (N_14569,N_14379,N_14300);
and U14570 (N_14570,N_14335,N_14389);
xor U14571 (N_14571,N_14467,N_14448);
nor U14572 (N_14572,N_14401,N_14463);
and U14573 (N_14573,N_14355,N_14357);
and U14574 (N_14574,N_14497,N_14456);
nand U14575 (N_14575,N_14258,N_14344);
nand U14576 (N_14576,N_14277,N_14280);
xnor U14577 (N_14577,N_14435,N_14307);
nand U14578 (N_14578,N_14366,N_14391);
xnor U14579 (N_14579,N_14263,N_14291);
xor U14580 (N_14580,N_14486,N_14425);
nor U14581 (N_14581,N_14276,N_14483);
and U14582 (N_14582,N_14346,N_14320);
or U14583 (N_14583,N_14322,N_14390);
or U14584 (N_14584,N_14326,N_14270);
nand U14585 (N_14585,N_14317,N_14427);
nor U14586 (N_14586,N_14372,N_14474);
and U14587 (N_14587,N_14343,N_14347);
or U14588 (N_14588,N_14471,N_14340);
or U14589 (N_14589,N_14472,N_14383);
nand U14590 (N_14590,N_14323,N_14264);
nor U14591 (N_14591,N_14334,N_14327);
or U14592 (N_14592,N_14315,N_14374);
and U14593 (N_14593,N_14341,N_14402);
xor U14594 (N_14594,N_14251,N_14369);
nor U14595 (N_14595,N_14431,N_14284);
or U14596 (N_14596,N_14387,N_14313);
nor U14597 (N_14597,N_14362,N_14293);
xor U14598 (N_14598,N_14470,N_14351);
nand U14599 (N_14599,N_14294,N_14499);
nand U14600 (N_14600,N_14487,N_14332);
and U14601 (N_14601,N_14272,N_14329);
nand U14602 (N_14602,N_14441,N_14481);
nor U14603 (N_14603,N_14290,N_14436);
and U14604 (N_14604,N_14482,N_14285);
and U14605 (N_14605,N_14365,N_14498);
or U14606 (N_14606,N_14349,N_14254);
nor U14607 (N_14607,N_14400,N_14262);
nor U14608 (N_14608,N_14485,N_14476);
and U14609 (N_14609,N_14375,N_14267);
and U14610 (N_14610,N_14459,N_14269);
or U14611 (N_14611,N_14495,N_14312);
or U14612 (N_14612,N_14368,N_14265);
or U14613 (N_14613,N_14348,N_14306);
xor U14614 (N_14614,N_14418,N_14408);
nand U14615 (N_14615,N_14261,N_14484);
nor U14616 (N_14616,N_14353,N_14266);
nor U14617 (N_14617,N_14444,N_14257);
nand U14618 (N_14618,N_14275,N_14325);
or U14619 (N_14619,N_14381,N_14439);
and U14620 (N_14620,N_14287,N_14440);
xor U14621 (N_14621,N_14403,N_14447);
xor U14622 (N_14622,N_14415,N_14454);
or U14623 (N_14623,N_14282,N_14308);
xnor U14624 (N_14624,N_14388,N_14279);
and U14625 (N_14625,N_14484,N_14303);
and U14626 (N_14626,N_14315,N_14456);
xnor U14627 (N_14627,N_14436,N_14489);
and U14628 (N_14628,N_14269,N_14387);
or U14629 (N_14629,N_14452,N_14364);
xor U14630 (N_14630,N_14411,N_14306);
and U14631 (N_14631,N_14341,N_14403);
nand U14632 (N_14632,N_14461,N_14475);
nand U14633 (N_14633,N_14450,N_14495);
nand U14634 (N_14634,N_14299,N_14279);
or U14635 (N_14635,N_14363,N_14484);
and U14636 (N_14636,N_14373,N_14343);
xor U14637 (N_14637,N_14489,N_14445);
nand U14638 (N_14638,N_14374,N_14339);
or U14639 (N_14639,N_14282,N_14292);
xnor U14640 (N_14640,N_14326,N_14305);
nor U14641 (N_14641,N_14303,N_14346);
or U14642 (N_14642,N_14279,N_14324);
nand U14643 (N_14643,N_14393,N_14296);
and U14644 (N_14644,N_14407,N_14493);
nand U14645 (N_14645,N_14472,N_14337);
nand U14646 (N_14646,N_14265,N_14484);
nor U14647 (N_14647,N_14258,N_14301);
nor U14648 (N_14648,N_14332,N_14342);
and U14649 (N_14649,N_14315,N_14491);
xor U14650 (N_14650,N_14343,N_14405);
nor U14651 (N_14651,N_14476,N_14292);
nand U14652 (N_14652,N_14335,N_14422);
xnor U14653 (N_14653,N_14355,N_14438);
nor U14654 (N_14654,N_14254,N_14458);
and U14655 (N_14655,N_14379,N_14450);
xnor U14656 (N_14656,N_14359,N_14274);
xnor U14657 (N_14657,N_14351,N_14490);
xor U14658 (N_14658,N_14287,N_14263);
nor U14659 (N_14659,N_14326,N_14477);
nor U14660 (N_14660,N_14272,N_14442);
or U14661 (N_14661,N_14471,N_14368);
or U14662 (N_14662,N_14383,N_14347);
xnor U14663 (N_14663,N_14305,N_14425);
xnor U14664 (N_14664,N_14451,N_14253);
or U14665 (N_14665,N_14324,N_14410);
nand U14666 (N_14666,N_14359,N_14302);
nand U14667 (N_14667,N_14461,N_14471);
or U14668 (N_14668,N_14486,N_14394);
or U14669 (N_14669,N_14361,N_14432);
nor U14670 (N_14670,N_14269,N_14365);
xnor U14671 (N_14671,N_14458,N_14436);
and U14672 (N_14672,N_14402,N_14356);
nand U14673 (N_14673,N_14400,N_14356);
xnor U14674 (N_14674,N_14343,N_14452);
xnor U14675 (N_14675,N_14287,N_14281);
or U14676 (N_14676,N_14374,N_14455);
and U14677 (N_14677,N_14428,N_14389);
nor U14678 (N_14678,N_14401,N_14492);
xor U14679 (N_14679,N_14386,N_14368);
and U14680 (N_14680,N_14405,N_14373);
nand U14681 (N_14681,N_14482,N_14449);
or U14682 (N_14682,N_14301,N_14316);
nand U14683 (N_14683,N_14351,N_14275);
or U14684 (N_14684,N_14285,N_14274);
nor U14685 (N_14685,N_14444,N_14495);
nor U14686 (N_14686,N_14389,N_14424);
xnor U14687 (N_14687,N_14356,N_14452);
and U14688 (N_14688,N_14412,N_14304);
or U14689 (N_14689,N_14346,N_14302);
nand U14690 (N_14690,N_14292,N_14488);
nand U14691 (N_14691,N_14402,N_14390);
and U14692 (N_14692,N_14325,N_14469);
xor U14693 (N_14693,N_14451,N_14287);
xnor U14694 (N_14694,N_14405,N_14445);
or U14695 (N_14695,N_14265,N_14365);
or U14696 (N_14696,N_14266,N_14330);
xnor U14697 (N_14697,N_14302,N_14299);
xor U14698 (N_14698,N_14417,N_14448);
xnor U14699 (N_14699,N_14314,N_14437);
nor U14700 (N_14700,N_14363,N_14490);
or U14701 (N_14701,N_14448,N_14304);
or U14702 (N_14702,N_14296,N_14377);
nand U14703 (N_14703,N_14438,N_14409);
and U14704 (N_14704,N_14411,N_14353);
xor U14705 (N_14705,N_14367,N_14324);
nand U14706 (N_14706,N_14288,N_14321);
and U14707 (N_14707,N_14448,N_14383);
and U14708 (N_14708,N_14351,N_14499);
nand U14709 (N_14709,N_14264,N_14267);
nor U14710 (N_14710,N_14273,N_14338);
nand U14711 (N_14711,N_14294,N_14435);
nor U14712 (N_14712,N_14429,N_14290);
and U14713 (N_14713,N_14331,N_14307);
nand U14714 (N_14714,N_14317,N_14365);
xnor U14715 (N_14715,N_14342,N_14381);
nand U14716 (N_14716,N_14297,N_14462);
xor U14717 (N_14717,N_14396,N_14293);
and U14718 (N_14718,N_14472,N_14477);
nand U14719 (N_14719,N_14390,N_14296);
nor U14720 (N_14720,N_14346,N_14432);
nor U14721 (N_14721,N_14255,N_14406);
xor U14722 (N_14722,N_14326,N_14483);
xor U14723 (N_14723,N_14361,N_14338);
nor U14724 (N_14724,N_14363,N_14334);
or U14725 (N_14725,N_14486,N_14403);
nand U14726 (N_14726,N_14378,N_14352);
and U14727 (N_14727,N_14441,N_14319);
nand U14728 (N_14728,N_14387,N_14293);
nor U14729 (N_14729,N_14273,N_14385);
nand U14730 (N_14730,N_14423,N_14280);
or U14731 (N_14731,N_14344,N_14475);
or U14732 (N_14732,N_14302,N_14432);
xor U14733 (N_14733,N_14477,N_14485);
or U14734 (N_14734,N_14488,N_14353);
nand U14735 (N_14735,N_14268,N_14266);
and U14736 (N_14736,N_14469,N_14260);
and U14737 (N_14737,N_14399,N_14354);
nor U14738 (N_14738,N_14319,N_14366);
nor U14739 (N_14739,N_14420,N_14356);
nand U14740 (N_14740,N_14445,N_14285);
xnor U14741 (N_14741,N_14339,N_14280);
nand U14742 (N_14742,N_14293,N_14486);
nand U14743 (N_14743,N_14472,N_14317);
or U14744 (N_14744,N_14384,N_14413);
or U14745 (N_14745,N_14339,N_14308);
nand U14746 (N_14746,N_14499,N_14318);
nand U14747 (N_14747,N_14346,N_14499);
nand U14748 (N_14748,N_14416,N_14309);
nand U14749 (N_14749,N_14415,N_14418);
xor U14750 (N_14750,N_14668,N_14510);
xor U14751 (N_14751,N_14582,N_14579);
nor U14752 (N_14752,N_14698,N_14734);
and U14753 (N_14753,N_14622,N_14521);
nor U14754 (N_14754,N_14740,N_14679);
nor U14755 (N_14755,N_14595,N_14617);
xnor U14756 (N_14756,N_14523,N_14706);
nand U14757 (N_14757,N_14688,N_14725);
or U14758 (N_14758,N_14596,N_14500);
or U14759 (N_14759,N_14558,N_14546);
xnor U14760 (N_14760,N_14549,N_14509);
or U14761 (N_14761,N_14570,N_14682);
nor U14762 (N_14762,N_14605,N_14749);
or U14763 (N_14763,N_14718,N_14665);
or U14764 (N_14764,N_14527,N_14606);
or U14765 (N_14765,N_14647,N_14735);
xnor U14766 (N_14766,N_14673,N_14723);
nor U14767 (N_14767,N_14631,N_14654);
nor U14768 (N_14768,N_14738,N_14638);
nor U14769 (N_14769,N_14678,N_14694);
xor U14770 (N_14770,N_14737,N_14575);
xor U14771 (N_14771,N_14552,N_14711);
nand U14772 (N_14772,N_14634,N_14710);
and U14773 (N_14773,N_14586,N_14534);
xnor U14774 (N_14774,N_14644,N_14610);
and U14775 (N_14775,N_14651,N_14732);
nor U14776 (N_14776,N_14699,N_14611);
nand U14777 (N_14777,N_14614,N_14529);
or U14778 (N_14778,N_14720,N_14506);
nor U14779 (N_14779,N_14539,N_14573);
nor U14780 (N_14780,N_14733,N_14553);
and U14781 (N_14781,N_14674,N_14703);
or U14782 (N_14782,N_14649,N_14724);
or U14783 (N_14783,N_14685,N_14667);
or U14784 (N_14784,N_14680,N_14512);
nor U14785 (N_14785,N_14692,N_14592);
xor U14786 (N_14786,N_14600,N_14658);
and U14787 (N_14787,N_14603,N_14587);
nand U14788 (N_14788,N_14618,N_14642);
and U14789 (N_14789,N_14623,N_14508);
xnor U14790 (N_14790,N_14686,N_14722);
and U14791 (N_14791,N_14639,N_14628);
nand U14792 (N_14792,N_14503,N_14609);
nand U14793 (N_14793,N_14591,N_14637);
or U14794 (N_14794,N_14536,N_14513);
and U14795 (N_14795,N_14540,N_14619);
and U14796 (N_14796,N_14728,N_14677);
nand U14797 (N_14797,N_14683,N_14571);
and U14798 (N_14798,N_14602,N_14613);
nor U14799 (N_14799,N_14577,N_14726);
xor U14800 (N_14800,N_14630,N_14716);
nand U14801 (N_14801,N_14578,N_14650);
nand U14802 (N_14802,N_14648,N_14567);
or U14803 (N_14803,N_14709,N_14607);
or U14804 (N_14804,N_14541,N_14538);
xor U14805 (N_14805,N_14676,N_14608);
nor U14806 (N_14806,N_14507,N_14675);
and U14807 (N_14807,N_14743,N_14544);
nor U14808 (N_14808,N_14612,N_14656);
nor U14809 (N_14809,N_14629,N_14568);
and U14810 (N_14810,N_14632,N_14700);
nand U14811 (N_14811,N_14559,N_14655);
and U14812 (N_14812,N_14712,N_14601);
nor U14813 (N_14813,N_14746,N_14528);
nand U14814 (N_14814,N_14621,N_14660);
xnor U14815 (N_14815,N_14585,N_14548);
nor U14816 (N_14816,N_14641,N_14670);
xor U14817 (N_14817,N_14652,N_14659);
and U14818 (N_14818,N_14542,N_14730);
and U14819 (N_14819,N_14616,N_14620);
nor U14820 (N_14820,N_14545,N_14727);
or U14821 (N_14821,N_14731,N_14531);
nand U14822 (N_14822,N_14717,N_14689);
xnor U14823 (N_14823,N_14627,N_14633);
xnor U14824 (N_14824,N_14705,N_14671);
nor U14825 (N_14825,N_14520,N_14533);
nor U14826 (N_14826,N_14526,N_14708);
nand U14827 (N_14827,N_14530,N_14625);
nand U14828 (N_14828,N_14624,N_14581);
or U14829 (N_14829,N_14547,N_14714);
nand U14830 (N_14830,N_14704,N_14560);
nand U14831 (N_14831,N_14604,N_14590);
xnor U14832 (N_14832,N_14646,N_14701);
xnor U14833 (N_14833,N_14669,N_14742);
xnor U14834 (N_14834,N_14696,N_14691);
nor U14835 (N_14835,N_14518,N_14713);
nand U14836 (N_14836,N_14672,N_14745);
xor U14837 (N_14837,N_14741,N_14511);
xnor U14838 (N_14838,N_14572,N_14597);
xor U14839 (N_14839,N_14556,N_14532);
xnor U14840 (N_14840,N_14588,N_14635);
xor U14841 (N_14841,N_14574,N_14519);
and U14842 (N_14842,N_14565,N_14643);
or U14843 (N_14843,N_14666,N_14525);
xnor U14844 (N_14844,N_14636,N_14517);
nand U14845 (N_14845,N_14557,N_14663);
and U14846 (N_14846,N_14748,N_14569);
nand U14847 (N_14847,N_14684,N_14583);
nor U14848 (N_14848,N_14576,N_14697);
nor U14849 (N_14849,N_14645,N_14593);
or U14850 (N_14850,N_14640,N_14555);
nor U14851 (N_14851,N_14739,N_14502);
nor U14852 (N_14852,N_14687,N_14580);
and U14853 (N_14853,N_14543,N_14661);
and U14854 (N_14854,N_14664,N_14615);
nor U14855 (N_14855,N_14515,N_14721);
xnor U14856 (N_14856,N_14504,N_14662);
nand U14857 (N_14857,N_14566,N_14522);
nand U14858 (N_14858,N_14693,N_14681);
xor U14859 (N_14859,N_14554,N_14653);
nor U14860 (N_14860,N_14564,N_14561);
or U14861 (N_14861,N_14736,N_14505);
and U14862 (N_14862,N_14562,N_14563);
nor U14863 (N_14863,N_14702,N_14514);
and U14864 (N_14864,N_14690,N_14537);
nand U14865 (N_14865,N_14626,N_14747);
nor U14866 (N_14866,N_14729,N_14719);
and U14867 (N_14867,N_14695,N_14594);
xnor U14868 (N_14868,N_14598,N_14516);
xnor U14869 (N_14869,N_14599,N_14744);
and U14870 (N_14870,N_14551,N_14584);
xnor U14871 (N_14871,N_14501,N_14524);
or U14872 (N_14872,N_14589,N_14715);
xnor U14873 (N_14873,N_14535,N_14707);
nor U14874 (N_14874,N_14657,N_14550);
nor U14875 (N_14875,N_14651,N_14697);
nand U14876 (N_14876,N_14510,N_14597);
or U14877 (N_14877,N_14649,N_14549);
or U14878 (N_14878,N_14593,N_14720);
or U14879 (N_14879,N_14686,N_14741);
or U14880 (N_14880,N_14523,N_14594);
nor U14881 (N_14881,N_14605,N_14655);
and U14882 (N_14882,N_14572,N_14629);
or U14883 (N_14883,N_14569,N_14534);
or U14884 (N_14884,N_14609,N_14739);
or U14885 (N_14885,N_14680,N_14665);
nor U14886 (N_14886,N_14649,N_14662);
and U14887 (N_14887,N_14553,N_14569);
xor U14888 (N_14888,N_14606,N_14626);
and U14889 (N_14889,N_14632,N_14548);
nor U14890 (N_14890,N_14684,N_14641);
or U14891 (N_14891,N_14728,N_14564);
nor U14892 (N_14892,N_14563,N_14722);
nor U14893 (N_14893,N_14619,N_14657);
and U14894 (N_14894,N_14726,N_14610);
nand U14895 (N_14895,N_14740,N_14690);
and U14896 (N_14896,N_14717,N_14653);
or U14897 (N_14897,N_14513,N_14509);
or U14898 (N_14898,N_14615,N_14551);
xnor U14899 (N_14899,N_14611,N_14686);
and U14900 (N_14900,N_14569,N_14540);
and U14901 (N_14901,N_14718,N_14739);
nor U14902 (N_14902,N_14619,N_14745);
nand U14903 (N_14903,N_14542,N_14509);
nor U14904 (N_14904,N_14560,N_14642);
xnor U14905 (N_14905,N_14613,N_14642);
nand U14906 (N_14906,N_14741,N_14705);
and U14907 (N_14907,N_14618,N_14603);
or U14908 (N_14908,N_14747,N_14537);
and U14909 (N_14909,N_14625,N_14501);
and U14910 (N_14910,N_14552,N_14737);
and U14911 (N_14911,N_14673,N_14679);
xor U14912 (N_14912,N_14616,N_14531);
xnor U14913 (N_14913,N_14683,N_14665);
nor U14914 (N_14914,N_14605,N_14746);
nor U14915 (N_14915,N_14529,N_14510);
or U14916 (N_14916,N_14749,N_14527);
nand U14917 (N_14917,N_14562,N_14631);
or U14918 (N_14918,N_14508,N_14525);
or U14919 (N_14919,N_14720,N_14501);
nand U14920 (N_14920,N_14746,N_14725);
xnor U14921 (N_14921,N_14741,N_14735);
nand U14922 (N_14922,N_14566,N_14592);
xnor U14923 (N_14923,N_14556,N_14526);
or U14924 (N_14924,N_14570,N_14662);
nor U14925 (N_14925,N_14555,N_14704);
and U14926 (N_14926,N_14695,N_14699);
nor U14927 (N_14927,N_14728,N_14725);
nand U14928 (N_14928,N_14559,N_14589);
xor U14929 (N_14929,N_14670,N_14669);
and U14930 (N_14930,N_14580,N_14645);
nand U14931 (N_14931,N_14571,N_14576);
nand U14932 (N_14932,N_14657,N_14681);
nor U14933 (N_14933,N_14745,N_14560);
or U14934 (N_14934,N_14743,N_14688);
nor U14935 (N_14935,N_14509,N_14669);
xor U14936 (N_14936,N_14748,N_14529);
nor U14937 (N_14937,N_14550,N_14621);
xor U14938 (N_14938,N_14559,N_14576);
xnor U14939 (N_14939,N_14673,N_14509);
or U14940 (N_14940,N_14565,N_14617);
nor U14941 (N_14941,N_14549,N_14680);
or U14942 (N_14942,N_14506,N_14726);
xor U14943 (N_14943,N_14549,N_14623);
xnor U14944 (N_14944,N_14718,N_14503);
nand U14945 (N_14945,N_14649,N_14616);
or U14946 (N_14946,N_14675,N_14715);
nand U14947 (N_14947,N_14687,N_14517);
nand U14948 (N_14948,N_14628,N_14687);
nand U14949 (N_14949,N_14591,N_14716);
and U14950 (N_14950,N_14668,N_14712);
xnor U14951 (N_14951,N_14741,N_14580);
and U14952 (N_14952,N_14671,N_14740);
and U14953 (N_14953,N_14721,N_14701);
nor U14954 (N_14954,N_14539,N_14583);
nor U14955 (N_14955,N_14643,N_14533);
and U14956 (N_14956,N_14730,N_14592);
xnor U14957 (N_14957,N_14528,N_14530);
and U14958 (N_14958,N_14556,N_14694);
nand U14959 (N_14959,N_14731,N_14596);
nand U14960 (N_14960,N_14667,N_14625);
nand U14961 (N_14961,N_14728,N_14693);
or U14962 (N_14962,N_14537,N_14624);
xor U14963 (N_14963,N_14652,N_14567);
and U14964 (N_14964,N_14666,N_14655);
nor U14965 (N_14965,N_14547,N_14671);
and U14966 (N_14966,N_14530,N_14731);
or U14967 (N_14967,N_14742,N_14578);
or U14968 (N_14968,N_14651,N_14546);
xnor U14969 (N_14969,N_14568,N_14513);
nand U14970 (N_14970,N_14720,N_14683);
nor U14971 (N_14971,N_14672,N_14505);
and U14972 (N_14972,N_14699,N_14595);
or U14973 (N_14973,N_14699,N_14552);
nand U14974 (N_14974,N_14705,N_14568);
nand U14975 (N_14975,N_14698,N_14697);
xor U14976 (N_14976,N_14671,N_14619);
xor U14977 (N_14977,N_14685,N_14666);
nand U14978 (N_14978,N_14535,N_14672);
or U14979 (N_14979,N_14653,N_14688);
nor U14980 (N_14980,N_14678,N_14741);
nor U14981 (N_14981,N_14620,N_14558);
nand U14982 (N_14982,N_14635,N_14678);
nand U14983 (N_14983,N_14733,N_14681);
or U14984 (N_14984,N_14744,N_14621);
nand U14985 (N_14985,N_14670,N_14672);
or U14986 (N_14986,N_14655,N_14699);
xor U14987 (N_14987,N_14507,N_14661);
and U14988 (N_14988,N_14509,N_14537);
nand U14989 (N_14989,N_14526,N_14643);
nand U14990 (N_14990,N_14540,N_14732);
or U14991 (N_14991,N_14730,N_14637);
nand U14992 (N_14992,N_14593,N_14649);
and U14993 (N_14993,N_14500,N_14573);
xor U14994 (N_14994,N_14704,N_14589);
and U14995 (N_14995,N_14546,N_14667);
nand U14996 (N_14996,N_14600,N_14704);
xnor U14997 (N_14997,N_14630,N_14598);
nand U14998 (N_14998,N_14698,N_14515);
and U14999 (N_14999,N_14581,N_14679);
xor U15000 (N_15000,N_14945,N_14764);
xnor U15001 (N_15001,N_14944,N_14954);
nand U15002 (N_15002,N_14780,N_14797);
nand U15003 (N_15003,N_14993,N_14960);
nand U15004 (N_15004,N_14817,N_14928);
nor U15005 (N_15005,N_14980,N_14950);
nor U15006 (N_15006,N_14885,N_14992);
nor U15007 (N_15007,N_14899,N_14752);
and U15008 (N_15008,N_14793,N_14852);
or U15009 (N_15009,N_14922,N_14761);
and U15010 (N_15010,N_14844,N_14925);
nor U15011 (N_15011,N_14838,N_14792);
xnor U15012 (N_15012,N_14995,N_14805);
xnor U15013 (N_15013,N_14896,N_14860);
and U15014 (N_15014,N_14831,N_14847);
and U15015 (N_15015,N_14964,N_14789);
xor U15016 (N_15016,N_14875,N_14753);
and U15017 (N_15017,N_14905,N_14946);
nor U15018 (N_15018,N_14943,N_14953);
nor U15019 (N_15019,N_14903,N_14756);
or U15020 (N_15020,N_14842,N_14877);
nor U15021 (N_15021,N_14982,N_14975);
xor U15022 (N_15022,N_14806,N_14812);
and U15023 (N_15023,N_14892,N_14799);
or U15024 (N_15024,N_14777,N_14942);
and U15025 (N_15025,N_14949,N_14791);
nand U15026 (N_15026,N_14986,N_14781);
or U15027 (N_15027,N_14801,N_14839);
or U15028 (N_15028,N_14814,N_14965);
nand U15029 (N_15029,N_14865,N_14935);
or U15030 (N_15030,N_14878,N_14873);
xor U15031 (N_15031,N_14917,N_14809);
nand U15032 (N_15032,N_14826,N_14768);
nor U15033 (N_15033,N_14807,N_14947);
or U15034 (N_15034,N_14895,N_14904);
nor U15035 (N_15035,N_14908,N_14759);
and U15036 (N_15036,N_14921,N_14835);
nand U15037 (N_15037,N_14959,N_14971);
and U15038 (N_15038,N_14923,N_14999);
nand U15039 (N_15039,N_14762,N_14914);
and U15040 (N_15040,N_14751,N_14910);
or U15041 (N_15041,N_14821,N_14803);
or U15042 (N_15042,N_14977,N_14888);
nor U15043 (N_15043,N_14936,N_14989);
nor U15044 (N_15044,N_14769,N_14798);
nand U15045 (N_15045,N_14871,N_14783);
nor U15046 (N_15046,N_14926,N_14802);
nor U15047 (N_15047,N_14952,N_14787);
nand U15048 (N_15048,N_14760,N_14755);
nand U15049 (N_15049,N_14879,N_14909);
nor U15050 (N_15050,N_14851,N_14939);
nor U15051 (N_15051,N_14984,N_14819);
and U15052 (N_15052,N_14786,N_14775);
xnor U15053 (N_15053,N_14828,N_14957);
nor U15054 (N_15054,N_14836,N_14985);
or U15055 (N_15055,N_14998,N_14815);
nand U15056 (N_15056,N_14973,N_14778);
and U15057 (N_15057,N_14902,N_14932);
or U15058 (N_15058,N_14848,N_14773);
xnor U15059 (N_15059,N_14988,N_14820);
and U15060 (N_15060,N_14987,N_14996);
nor U15061 (N_15061,N_14933,N_14808);
nand U15062 (N_15062,N_14884,N_14754);
and U15063 (N_15063,N_14767,N_14758);
nor U15064 (N_15064,N_14931,N_14859);
nand U15065 (N_15065,N_14800,N_14887);
or U15066 (N_15066,N_14834,N_14927);
nor U15067 (N_15067,N_14890,N_14765);
or U15068 (N_15068,N_14862,N_14850);
or U15069 (N_15069,N_14958,N_14937);
nor U15070 (N_15070,N_14855,N_14916);
xnor U15071 (N_15071,N_14963,N_14837);
or U15072 (N_15072,N_14840,N_14856);
or U15073 (N_15073,N_14804,N_14938);
nor U15074 (N_15074,N_14997,N_14981);
and U15075 (N_15075,N_14880,N_14853);
and U15076 (N_15076,N_14920,N_14881);
xnor U15077 (N_15077,N_14874,N_14849);
or U15078 (N_15078,N_14841,N_14962);
nor U15079 (N_15079,N_14955,N_14845);
nor U15080 (N_15080,N_14823,N_14915);
nor U15081 (N_15081,N_14824,N_14846);
and U15082 (N_15082,N_14951,N_14779);
and U15083 (N_15083,N_14940,N_14757);
nor U15084 (N_15084,N_14961,N_14968);
or U15085 (N_15085,N_14872,N_14766);
or U15086 (N_15086,N_14869,N_14970);
nor U15087 (N_15087,N_14919,N_14790);
nand U15088 (N_15088,N_14913,N_14911);
and U15089 (N_15089,N_14934,N_14900);
and U15090 (N_15090,N_14893,N_14827);
nor U15091 (N_15091,N_14948,N_14774);
nand U15092 (N_15092,N_14882,N_14924);
or U15093 (N_15093,N_14991,N_14784);
and U15094 (N_15094,N_14897,N_14941);
or U15095 (N_15095,N_14788,N_14969);
nor U15096 (N_15096,N_14883,N_14907);
and U15097 (N_15097,N_14843,N_14794);
or U15098 (N_15098,N_14857,N_14816);
nor U15099 (N_15099,N_14898,N_14864);
xor U15100 (N_15100,N_14876,N_14811);
and U15101 (N_15101,N_14912,N_14763);
xor U15102 (N_15102,N_14854,N_14863);
nor U15103 (N_15103,N_14796,N_14967);
nor U15104 (N_15104,N_14889,N_14906);
or U15105 (N_15105,N_14976,N_14858);
or U15106 (N_15106,N_14974,N_14825);
nor U15107 (N_15107,N_14866,N_14822);
nand U15108 (N_15108,N_14994,N_14829);
xor U15109 (N_15109,N_14979,N_14956);
nand U15110 (N_15110,N_14861,N_14813);
nor U15111 (N_15111,N_14810,N_14830);
or U15112 (N_15112,N_14918,N_14983);
nand U15113 (N_15113,N_14972,N_14870);
or U15114 (N_15114,N_14782,N_14832);
nor U15115 (N_15115,N_14886,N_14978);
nand U15116 (N_15116,N_14891,N_14772);
nor U15117 (N_15117,N_14894,N_14770);
xor U15118 (N_15118,N_14750,N_14901);
and U15119 (N_15119,N_14990,N_14867);
xnor U15120 (N_15120,N_14795,N_14771);
or U15121 (N_15121,N_14966,N_14785);
xor U15122 (N_15122,N_14929,N_14818);
nand U15123 (N_15123,N_14776,N_14868);
or U15124 (N_15124,N_14833,N_14930);
xnor U15125 (N_15125,N_14962,N_14788);
and U15126 (N_15126,N_14880,N_14995);
xor U15127 (N_15127,N_14870,N_14935);
or U15128 (N_15128,N_14996,N_14790);
or U15129 (N_15129,N_14892,N_14819);
xor U15130 (N_15130,N_14778,N_14980);
nor U15131 (N_15131,N_14755,N_14818);
nor U15132 (N_15132,N_14961,N_14942);
nor U15133 (N_15133,N_14772,N_14920);
nor U15134 (N_15134,N_14831,N_14855);
and U15135 (N_15135,N_14757,N_14896);
nor U15136 (N_15136,N_14962,N_14892);
xnor U15137 (N_15137,N_14983,N_14929);
nand U15138 (N_15138,N_14787,N_14762);
or U15139 (N_15139,N_14826,N_14857);
nand U15140 (N_15140,N_14839,N_14761);
or U15141 (N_15141,N_14768,N_14973);
nor U15142 (N_15142,N_14988,N_14901);
nand U15143 (N_15143,N_14949,N_14953);
xor U15144 (N_15144,N_14817,N_14753);
or U15145 (N_15145,N_14800,N_14858);
and U15146 (N_15146,N_14820,N_14836);
and U15147 (N_15147,N_14957,N_14857);
and U15148 (N_15148,N_14958,N_14897);
xor U15149 (N_15149,N_14858,N_14846);
nor U15150 (N_15150,N_14935,N_14802);
nand U15151 (N_15151,N_14784,N_14878);
xor U15152 (N_15152,N_14751,N_14758);
nor U15153 (N_15153,N_14762,N_14850);
nor U15154 (N_15154,N_14906,N_14961);
and U15155 (N_15155,N_14766,N_14861);
nand U15156 (N_15156,N_14867,N_14833);
nand U15157 (N_15157,N_14817,N_14812);
and U15158 (N_15158,N_14833,N_14807);
nor U15159 (N_15159,N_14930,N_14754);
xnor U15160 (N_15160,N_14850,N_14907);
nand U15161 (N_15161,N_14786,N_14845);
or U15162 (N_15162,N_14920,N_14784);
xor U15163 (N_15163,N_14924,N_14958);
and U15164 (N_15164,N_14854,N_14918);
and U15165 (N_15165,N_14958,N_14882);
nor U15166 (N_15166,N_14926,N_14940);
xor U15167 (N_15167,N_14828,N_14906);
nor U15168 (N_15168,N_14793,N_14931);
nor U15169 (N_15169,N_14881,N_14999);
nand U15170 (N_15170,N_14883,N_14790);
or U15171 (N_15171,N_14861,N_14844);
nand U15172 (N_15172,N_14984,N_14940);
xor U15173 (N_15173,N_14849,N_14952);
or U15174 (N_15174,N_14978,N_14961);
or U15175 (N_15175,N_14894,N_14873);
and U15176 (N_15176,N_14839,N_14987);
nor U15177 (N_15177,N_14990,N_14919);
and U15178 (N_15178,N_14762,N_14909);
nor U15179 (N_15179,N_14783,N_14842);
xnor U15180 (N_15180,N_14768,N_14992);
and U15181 (N_15181,N_14911,N_14779);
nor U15182 (N_15182,N_14805,N_14912);
or U15183 (N_15183,N_14816,N_14817);
and U15184 (N_15184,N_14975,N_14845);
xnor U15185 (N_15185,N_14979,N_14776);
and U15186 (N_15186,N_14854,N_14947);
xnor U15187 (N_15187,N_14896,N_14935);
nor U15188 (N_15188,N_14782,N_14762);
and U15189 (N_15189,N_14952,N_14751);
nor U15190 (N_15190,N_14860,N_14780);
or U15191 (N_15191,N_14932,N_14984);
xnor U15192 (N_15192,N_14917,N_14771);
or U15193 (N_15193,N_14948,N_14934);
nand U15194 (N_15194,N_14789,N_14906);
and U15195 (N_15195,N_14820,N_14928);
or U15196 (N_15196,N_14852,N_14836);
nand U15197 (N_15197,N_14863,N_14767);
xor U15198 (N_15198,N_14768,N_14774);
nor U15199 (N_15199,N_14885,N_14813);
nor U15200 (N_15200,N_14788,N_14935);
nor U15201 (N_15201,N_14816,N_14969);
nor U15202 (N_15202,N_14875,N_14985);
or U15203 (N_15203,N_14938,N_14997);
nor U15204 (N_15204,N_14971,N_14836);
nand U15205 (N_15205,N_14892,N_14766);
nand U15206 (N_15206,N_14768,N_14829);
xnor U15207 (N_15207,N_14862,N_14984);
xnor U15208 (N_15208,N_14904,N_14930);
nor U15209 (N_15209,N_14981,N_14978);
nand U15210 (N_15210,N_14759,N_14900);
nand U15211 (N_15211,N_14887,N_14929);
nand U15212 (N_15212,N_14880,N_14865);
xor U15213 (N_15213,N_14886,N_14996);
or U15214 (N_15214,N_14761,N_14860);
or U15215 (N_15215,N_14787,N_14931);
and U15216 (N_15216,N_14987,N_14837);
and U15217 (N_15217,N_14973,N_14793);
nor U15218 (N_15218,N_14792,N_14864);
and U15219 (N_15219,N_14955,N_14976);
xnor U15220 (N_15220,N_14786,N_14865);
and U15221 (N_15221,N_14789,N_14982);
and U15222 (N_15222,N_14795,N_14801);
xnor U15223 (N_15223,N_14846,N_14793);
nand U15224 (N_15224,N_14784,N_14886);
nand U15225 (N_15225,N_14765,N_14854);
or U15226 (N_15226,N_14822,N_14915);
and U15227 (N_15227,N_14802,N_14987);
or U15228 (N_15228,N_14823,N_14764);
and U15229 (N_15229,N_14777,N_14965);
xor U15230 (N_15230,N_14975,N_14913);
xor U15231 (N_15231,N_14900,N_14908);
xor U15232 (N_15232,N_14883,N_14934);
nor U15233 (N_15233,N_14966,N_14777);
xor U15234 (N_15234,N_14973,N_14846);
or U15235 (N_15235,N_14826,N_14840);
nand U15236 (N_15236,N_14869,N_14897);
nand U15237 (N_15237,N_14825,N_14797);
or U15238 (N_15238,N_14934,N_14952);
xor U15239 (N_15239,N_14751,N_14958);
and U15240 (N_15240,N_14808,N_14947);
nor U15241 (N_15241,N_14761,N_14756);
or U15242 (N_15242,N_14782,N_14909);
or U15243 (N_15243,N_14970,N_14998);
and U15244 (N_15244,N_14884,N_14966);
or U15245 (N_15245,N_14791,N_14753);
nor U15246 (N_15246,N_14932,N_14769);
nand U15247 (N_15247,N_14779,N_14936);
xor U15248 (N_15248,N_14842,N_14871);
nor U15249 (N_15249,N_14944,N_14862);
nand U15250 (N_15250,N_15114,N_15105);
or U15251 (N_15251,N_15241,N_15240);
or U15252 (N_15252,N_15090,N_15118);
nand U15253 (N_15253,N_15142,N_15186);
nor U15254 (N_15254,N_15139,N_15202);
nor U15255 (N_15255,N_15169,N_15013);
xnor U15256 (N_15256,N_15049,N_15191);
xnor U15257 (N_15257,N_15155,N_15144);
nor U15258 (N_15258,N_15089,N_15020);
nand U15259 (N_15259,N_15168,N_15182);
and U15260 (N_15260,N_15231,N_15172);
xor U15261 (N_15261,N_15236,N_15085);
or U15262 (N_15262,N_15154,N_15176);
nor U15263 (N_15263,N_15037,N_15216);
nor U15264 (N_15264,N_15164,N_15012);
and U15265 (N_15265,N_15221,N_15199);
or U15266 (N_15266,N_15131,N_15080);
and U15267 (N_15267,N_15094,N_15051);
nand U15268 (N_15268,N_15235,N_15219);
or U15269 (N_15269,N_15092,N_15067);
nand U15270 (N_15270,N_15185,N_15061);
or U15271 (N_15271,N_15224,N_15163);
nor U15272 (N_15272,N_15156,N_15056);
nor U15273 (N_15273,N_15147,N_15053);
or U15274 (N_15274,N_15245,N_15178);
xor U15275 (N_15275,N_15009,N_15135);
nand U15276 (N_15276,N_15032,N_15023);
and U15277 (N_15277,N_15208,N_15126);
xor U15278 (N_15278,N_15054,N_15174);
or U15279 (N_15279,N_15160,N_15116);
or U15280 (N_15280,N_15151,N_15138);
or U15281 (N_15281,N_15211,N_15152);
xor U15282 (N_15282,N_15048,N_15076);
xor U15283 (N_15283,N_15077,N_15022);
nand U15284 (N_15284,N_15088,N_15228);
or U15285 (N_15285,N_15084,N_15187);
nor U15286 (N_15286,N_15098,N_15002);
nand U15287 (N_15287,N_15119,N_15166);
nor U15288 (N_15288,N_15093,N_15081);
nor U15289 (N_15289,N_15167,N_15045);
or U15290 (N_15290,N_15181,N_15003);
nand U15291 (N_15291,N_15004,N_15043);
nand U15292 (N_15292,N_15158,N_15226);
nand U15293 (N_15293,N_15217,N_15177);
xnor U15294 (N_15294,N_15055,N_15001);
and U15295 (N_15295,N_15227,N_15150);
nor U15296 (N_15296,N_15014,N_15115);
xnor U15297 (N_15297,N_15060,N_15243);
and U15298 (N_15298,N_15042,N_15040);
and U15299 (N_15299,N_15058,N_15173);
xor U15300 (N_15300,N_15161,N_15196);
and U15301 (N_15301,N_15159,N_15036);
nand U15302 (N_15302,N_15021,N_15044);
xnor U15303 (N_15303,N_15179,N_15189);
or U15304 (N_15304,N_15145,N_15108);
xnor U15305 (N_15305,N_15071,N_15242);
or U15306 (N_15306,N_15033,N_15206);
xnor U15307 (N_15307,N_15097,N_15095);
xor U15308 (N_15308,N_15210,N_15008);
or U15309 (N_15309,N_15079,N_15006);
and U15310 (N_15310,N_15096,N_15019);
and U15311 (N_15311,N_15062,N_15148);
and U15312 (N_15312,N_15034,N_15130);
nor U15313 (N_15313,N_15101,N_15025);
and U15314 (N_15314,N_15068,N_15143);
and U15315 (N_15315,N_15165,N_15057);
and U15316 (N_15316,N_15074,N_15244);
xnor U15317 (N_15317,N_15229,N_15201);
nand U15318 (N_15318,N_15180,N_15117);
xor U15319 (N_15319,N_15247,N_15125);
and U15320 (N_15320,N_15220,N_15213);
and U15321 (N_15321,N_15141,N_15171);
xor U15322 (N_15322,N_15075,N_15027);
nand U15323 (N_15323,N_15234,N_15153);
and U15324 (N_15324,N_15207,N_15050);
nor U15325 (N_15325,N_15222,N_15212);
nand U15326 (N_15326,N_15183,N_15066);
nor U15327 (N_15327,N_15200,N_15188);
nor U15328 (N_15328,N_15112,N_15065);
nand U15329 (N_15329,N_15017,N_15195);
xor U15330 (N_15330,N_15007,N_15120);
nand U15331 (N_15331,N_15078,N_15010);
xor U15332 (N_15332,N_15133,N_15106);
or U15333 (N_15333,N_15215,N_15073);
xnor U15334 (N_15334,N_15030,N_15121);
xor U15335 (N_15335,N_15083,N_15104);
and U15336 (N_15336,N_15197,N_15005);
nor U15337 (N_15337,N_15099,N_15232);
xnor U15338 (N_15338,N_15136,N_15249);
xnor U15339 (N_15339,N_15122,N_15192);
nor U15340 (N_15340,N_15204,N_15132);
nor U15341 (N_15341,N_15052,N_15137);
nor U15342 (N_15342,N_15016,N_15233);
nand U15343 (N_15343,N_15248,N_15184);
nor U15344 (N_15344,N_15129,N_15011);
or U15345 (N_15345,N_15047,N_15072);
xor U15346 (N_15346,N_15087,N_15237);
and U15347 (N_15347,N_15123,N_15046);
and U15348 (N_15348,N_15026,N_15086);
or U15349 (N_15349,N_15162,N_15175);
xor U15350 (N_15350,N_15239,N_15103);
or U15351 (N_15351,N_15015,N_15024);
nor U15352 (N_15352,N_15134,N_15028);
nor U15353 (N_15353,N_15128,N_15107);
and U15354 (N_15354,N_15238,N_15100);
or U15355 (N_15355,N_15039,N_15069);
or U15356 (N_15356,N_15018,N_15140);
nor U15357 (N_15357,N_15198,N_15038);
nor U15358 (N_15358,N_15124,N_15246);
nor U15359 (N_15359,N_15063,N_15190);
nand U15360 (N_15360,N_15193,N_15091);
nand U15361 (N_15361,N_15209,N_15102);
nand U15362 (N_15362,N_15127,N_15064);
nor U15363 (N_15363,N_15109,N_15149);
nor U15364 (N_15364,N_15035,N_15230);
xnor U15365 (N_15365,N_15059,N_15029);
nand U15366 (N_15366,N_15225,N_15146);
or U15367 (N_15367,N_15223,N_15082);
and U15368 (N_15368,N_15110,N_15111);
nor U15369 (N_15369,N_15000,N_15194);
nor U15370 (N_15370,N_15205,N_15031);
nand U15371 (N_15371,N_15170,N_15070);
xor U15372 (N_15372,N_15041,N_15113);
and U15373 (N_15373,N_15214,N_15218);
nor U15374 (N_15374,N_15157,N_15203);
nor U15375 (N_15375,N_15101,N_15074);
xnor U15376 (N_15376,N_15165,N_15114);
or U15377 (N_15377,N_15232,N_15059);
and U15378 (N_15378,N_15137,N_15144);
and U15379 (N_15379,N_15110,N_15206);
xor U15380 (N_15380,N_15230,N_15203);
xor U15381 (N_15381,N_15087,N_15051);
and U15382 (N_15382,N_15023,N_15008);
nand U15383 (N_15383,N_15200,N_15119);
nand U15384 (N_15384,N_15002,N_15114);
nand U15385 (N_15385,N_15165,N_15164);
or U15386 (N_15386,N_15174,N_15105);
and U15387 (N_15387,N_15189,N_15015);
and U15388 (N_15388,N_15094,N_15025);
nor U15389 (N_15389,N_15123,N_15216);
nor U15390 (N_15390,N_15219,N_15071);
nand U15391 (N_15391,N_15233,N_15103);
nor U15392 (N_15392,N_15078,N_15247);
xor U15393 (N_15393,N_15128,N_15101);
nor U15394 (N_15394,N_15042,N_15097);
nand U15395 (N_15395,N_15192,N_15132);
and U15396 (N_15396,N_15213,N_15021);
nor U15397 (N_15397,N_15224,N_15084);
and U15398 (N_15398,N_15092,N_15143);
and U15399 (N_15399,N_15209,N_15190);
nor U15400 (N_15400,N_15067,N_15068);
xnor U15401 (N_15401,N_15094,N_15202);
xnor U15402 (N_15402,N_15075,N_15172);
xnor U15403 (N_15403,N_15119,N_15099);
nand U15404 (N_15404,N_15043,N_15020);
or U15405 (N_15405,N_15026,N_15203);
and U15406 (N_15406,N_15019,N_15028);
and U15407 (N_15407,N_15042,N_15110);
nand U15408 (N_15408,N_15109,N_15047);
nor U15409 (N_15409,N_15125,N_15084);
xor U15410 (N_15410,N_15159,N_15095);
nand U15411 (N_15411,N_15210,N_15133);
xor U15412 (N_15412,N_15023,N_15121);
or U15413 (N_15413,N_15174,N_15215);
nor U15414 (N_15414,N_15074,N_15051);
xor U15415 (N_15415,N_15164,N_15211);
xor U15416 (N_15416,N_15154,N_15100);
nand U15417 (N_15417,N_15035,N_15160);
xor U15418 (N_15418,N_15061,N_15121);
nor U15419 (N_15419,N_15137,N_15205);
xor U15420 (N_15420,N_15081,N_15144);
nand U15421 (N_15421,N_15011,N_15013);
nor U15422 (N_15422,N_15145,N_15139);
nor U15423 (N_15423,N_15063,N_15096);
nor U15424 (N_15424,N_15090,N_15044);
xnor U15425 (N_15425,N_15069,N_15127);
nor U15426 (N_15426,N_15039,N_15025);
xor U15427 (N_15427,N_15163,N_15032);
nor U15428 (N_15428,N_15034,N_15230);
xnor U15429 (N_15429,N_15178,N_15109);
xor U15430 (N_15430,N_15110,N_15092);
nor U15431 (N_15431,N_15169,N_15015);
nand U15432 (N_15432,N_15017,N_15071);
or U15433 (N_15433,N_15117,N_15191);
xor U15434 (N_15434,N_15101,N_15055);
and U15435 (N_15435,N_15015,N_15060);
nand U15436 (N_15436,N_15072,N_15208);
nor U15437 (N_15437,N_15163,N_15187);
and U15438 (N_15438,N_15134,N_15204);
nand U15439 (N_15439,N_15211,N_15117);
nand U15440 (N_15440,N_15210,N_15209);
nand U15441 (N_15441,N_15218,N_15234);
nor U15442 (N_15442,N_15067,N_15209);
nand U15443 (N_15443,N_15131,N_15017);
nand U15444 (N_15444,N_15129,N_15115);
nand U15445 (N_15445,N_15112,N_15154);
or U15446 (N_15446,N_15124,N_15101);
or U15447 (N_15447,N_15023,N_15117);
xnor U15448 (N_15448,N_15157,N_15097);
nor U15449 (N_15449,N_15144,N_15103);
nand U15450 (N_15450,N_15166,N_15164);
and U15451 (N_15451,N_15175,N_15135);
nand U15452 (N_15452,N_15084,N_15225);
nor U15453 (N_15453,N_15245,N_15077);
nor U15454 (N_15454,N_15159,N_15204);
and U15455 (N_15455,N_15124,N_15106);
xnor U15456 (N_15456,N_15038,N_15051);
and U15457 (N_15457,N_15208,N_15157);
nand U15458 (N_15458,N_15235,N_15052);
nor U15459 (N_15459,N_15020,N_15238);
nand U15460 (N_15460,N_15235,N_15020);
or U15461 (N_15461,N_15142,N_15043);
nand U15462 (N_15462,N_15109,N_15239);
nand U15463 (N_15463,N_15149,N_15010);
nor U15464 (N_15464,N_15022,N_15068);
or U15465 (N_15465,N_15227,N_15009);
nand U15466 (N_15466,N_15104,N_15243);
xnor U15467 (N_15467,N_15120,N_15221);
nand U15468 (N_15468,N_15023,N_15099);
or U15469 (N_15469,N_15188,N_15083);
nor U15470 (N_15470,N_15138,N_15186);
nor U15471 (N_15471,N_15076,N_15119);
nor U15472 (N_15472,N_15018,N_15181);
and U15473 (N_15473,N_15156,N_15074);
nand U15474 (N_15474,N_15069,N_15061);
and U15475 (N_15475,N_15063,N_15245);
xnor U15476 (N_15476,N_15020,N_15000);
or U15477 (N_15477,N_15081,N_15219);
or U15478 (N_15478,N_15056,N_15127);
or U15479 (N_15479,N_15134,N_15133);
xnor U15480 (N_15480,N_15060,N_15129);
or U15481 (N_15481,N_15117,N_15161);
or U15482 (N_15482,N_15160,N_15113);
nand U15483 (N_15483,N_15027,N_15121);
nand U15484 (N_15484,N_15214,N_15203);
nor U15485 (N_15485,N_15111,N_15010);
xnor U15486 (N_15486,N_15204,N_15133);
or U15487 (N_15487,N_15233,N_15122);
nor U15488 (N_15488,N_15115,N_15232);
nor U15489 (N_15489,N_15137,N_15092);
or U15490 (N_15490,N_15077,N_15200);
and U15491 (N_15491,N_15193,N_15114);
or U15492 (N_15492,N_15242,N_15093);
nor U15493 (N_15493,N_15146,N_15111);
nand U15494 (N_15494,N_15075,N_15179);
nand U15495 (N_15495,N_15149,N_15241);
xnor U15496 (N_15496,N_15233,N_15119);
or U15497 (N_15497,N_15168,N_15000);
and U15498 (N_15498,N_15124,N_15120);
nand U15499 (N_15499,N_15045,N_15124);
or U15500 (N_15500,N_15405,N_15395);
nor U15501 (N_15501,N_15415,N_15269);
nand U15502 (N_15502,N_15447,N_15327);
nand U15503 (N_15503,N_15452,N_15303);
nand U15504 (N_15504,N_15433,N_15279);
nor U15505 (N_15505,N_15349,N_15258);
nor U15506 (N_15506,N_15440,N_15419);
nor U15507 (N_15507,N_15470,N_15272);
nor U15508 (N_15508,N_15277,N_15453);
and U15509 (N_15509,N_15449,N_15265);
xor U15510 (N_15510,N_15488,N_15469);
nand U15511 (N_15511,N_15271,N_15289);
and U15512 (N_15512,N_15370,N_15474);
and U15513 (N_15513,N_15264,N_15344);
nor U15514 (N_15514,N_15443,N_15495);
nand U15515 (N_15515,N_15260,N_15274);
or U15516 (N_15516,N_15311,N_15493);
xnor U15517 (N_15517,N_15430,N_15448);
and U15518 (N_15518,N_15280,N_15255);
and U15519 (N_15519,N_15499,N_15396);
nand U15520 (N_15520,N_15489,N_15334);
nor U15521 (N_15521,N_15391,N_15438);
nor U15522 (N_15522,N_15298,N_15444);
xnor U15523 (N_15523,N_15252,N_15445);
nand U15524 (N_15524,N_15356,N_15475);
and U15525 (N_15525,N_15473,N_15299);
and U15526 (N_15526,N_15418,N_15262);
nand U15527 (N_15527,N_15461,N_15388);
xor U15528 (N_15528,N_15292,N_15486);
and U15529 (N_15529,N_15250,N_15284);
or U15530 (N_15530,N_15427,N_15342);
nor U15531 (N_15531,N_15256,N_15350);
and U15532 (N_15532,N_15273,N_15472);
and U15533 (N_15533,N_15457,N_15476);
nand U15534 (N_15534,N_15336,N_15425);
nand U15535 (N_15535,N_15317,N_15335);
and U15536 (N_15536,N_15385,N_15439);
nand U15537 (N_15537,N_15376,N_15330);
nand U15538 (N_15538,N_15384,N_15351);
xor U15539 (N_15539,N_15429,N_15463);
nor U15540 (N_15540,N_15333,N_15362);
and U15541 (N_15541,N_15485,N_15466);
nor U15542 (N_15542,N_15383,N_15341);
and U15543 (N_15543,N_15367,N_15426);
or U15544 (N_15544,N_15328,N_15352);
nor U15545 (N_15545,N_15455,N_15421);
and U15546 (N_15546,N_15302,N_15295);
or U15547 (N_15547,N_15268,N_15481);
xnor U15548 (N_15548,N_15320,N_15313);
and U15549 (N_15549,N_15484,N_15436);
and U15550 (N_15550,N_15358,N_15324);
and U15551 (N_15551,N_15435,N_15413);
and U15552 (N_15552,N_15431,N_15454);
or U15553 (N_15553,N_15306,N_15373);
or U15554 (N_15554,N_15267,N_15315);
xor U15555 (N_15555,N_15393,N_15378);
nand U15556 (N_15556,N_15403,N_15287);
xnor U15557 (N_15557,N_15340,N_15451);
nor U15558 (N_15558,N_15307,N_15364);
nand U15559 (N_15559,N_15397,N_15490);
and U15560 (N_15560,N_15404,N_15323);
nand U15561 (N_15561,N_15354,N_15257);
nand U15562 (N_15562,N_15355,N_15291);
and U15563 (N_15563,N_15253,N_15305);
xor U15564 (N_15564,N_15346,N_15316);
or U15565 (N_15565,N_15266,N_15437);
xnor U15566 (N_15566,N_15487,N_15331);
or U15567 (N_15567,N_15275,N_15337);
or U15568 (N_15568,N_15310,N_15251);
nor U15569 (N_15569,N_15392,N_15468);
or U15570 (N_15570,N_15412,N_15497);
xnor U15571 (N_15571,N_15319,N_15417);
nand U15572 (N_15572,N_15312,N_15399);
and U15573 (N_15573,N_15377,N_15278);
or U15574 (N_15574,N_15398,N_15290);
and U15575 (N_15575,N_15283,N_15477);
xnor U15576 (N_15576,N_15282,N_15343);
nor U15577 (N_15577,N_15353,N_15288);
nor U15578 (N_15578,N_15394,N_15498);
nand U15579 (N_15579,N_15380,N_15365);
or U15580 (N_15580,N_15270,N_15366);
nand U15581 (N_15581,N_15479,N_15363);
nand U15582 (N_15582,N_15308,N_15326);
or U15583 (N_15583,N_15450,N_15329);
nand U15584 (N_15584,N_15401,N_15471);
and U15585 (N_15585,N_15357,N_15423);
and U15586 (N_15586,N_15478,N_15332);
and U15587 (N_15587,N_15459,N_15318);
nor U15588 (N_15588,N_15491,N_15390);
or U15589 (N_15589,N_15259,N_15345);
and U15590 (N_15590,N_15381,N_15371);
xnor U15591 (N_15591,N_15347,N_15314);
or U15592 (N_15592,N_15360,N_15386);
nor U15593 (N_15593,N_15482,N_15387);
xor U15594 (N_15594,N_15480,N_15296);
nor U15595 (N_15595,N_15309,N_15494);
xnor U15596 (N_15596,N_15441,N_15408);
or U15597 (N_15597,N_15424,N_15322);
xnor U15598 (N_15598,N_15338,N_15467);
or U15599 (N_15599,N_15422,N_15446);
and U15600 (N_15600,N_15297,N_15432);
xor U15601 (N_15601,N_15414,N_15458);
and U15602 (N_15602,N_15382,N_15379);
nand U15603 (N_15603,N_15416,N_15389);
nor U15604 (N_15604,N_15281,N_15301);
nor U15605 (N_15605,N_15400,N_15361);
or U15606 (N_15606,N_15434,N_15304);
xor U15607 (N_15607,N_15372,N_15293);
and U15608 (N_15608,N_15285,N_15254);
nor U15609 (N_15609,N_15261,N_15374);
xnor U15610 (N_15610,N_15464,N_15465);
nor U15611 (N_15611,N_15420,N_15409);
nand U15612 (N_15612,N_15483,N_15410);
xor U15613 (N_15613,N_15321,N_15348);
xnor U15614 (N_15614,N_15460,N_15368);
or U15615 (N_15615,N_15294,N_15286);
xor U15616 (N_15616,N_15462,N_15369);
nor U15617 (N_15617,N_15496,N_15411);
nor U15618 (N_15618,N_15263,N_15325);
nor U15619 (N_15619,N_15442,N_15402);
xor U15620 (N_15620,N_15359,N_15456);
and U15621 (N_15621,N_15406,N_15428);
and U15622 (N_15622,N_15375,N_15492);
xnor U15623 (N_15623,N_15276,N_15407);
or U15624 (N_15624,N_15300,N_15339);
nand U15625 (N_15625,N_15286,N_15291);
and U15626 (N_15626,N_15482,N_15334);
xor U15627 (N_15627,N_15467,N_15351);
nor U15628 (N_15628,N_15302,N_15279);
and U15629 (N_15629,N_15469,N_15284);
nand U15630 (N_15630,N_15468,N_15404);
nor U15631 (N_15631,N_15419,N_15420);
xnor U15632 (N_15632,N_15440,N_15369);
nor U15633 (N_15633,N_15416,N_15480);
xnor U15634 (N_15634,N_15401,N_15274);
and U15635 (N_15635,N_15379,N_15459);
nor U15636 (N_15636,N_15322,N_15368);
or U15637 (N_15637,N_15300,N_15328);
nor U15638 (N_15638,N_15339,N_15345);
nand U15639 (N_15639,N_15422,N_15250);
xnor U15640 (N_15640,N_15497,N_15293);
or U15641 (N_15641,N_15454,N_15479);
nor U15642 (N_15642,N_15399,N_15281);
nand U15643 (N_15643,N_15454,N_15405);
or U15644 (N_15644,N_15447,N_15475);
nand U15645 (N_15645,N_15253,N_15407);
nor U15646 (N_15646,N_15445,N_15408);
xnor U15647 (N_15647,N_15400,N_15467);
or U15648 (N_15648,N_15303,N_15407);
nor U15649 (N_15649,N_15494,N_15482);
or U15650 (N_15650,N_15256,N_15385);
and U15651 (N_15651,N_15440,N_15299);
xnor U15652 (N_15652,N_15383,N_15407);
nor U15653 (N_15653,N_15346,N_15280);
and U15654 (N_15654,N_15404,N_15415);
xnor U15655 (N_15655,N_15287,N_15389);
and U15656 (N_15656,N_15385,N_15251);
and U15657 (N_15657,N_15423,N_15343);
or U15658 (N_15658,N_15254,N_15471);
or U15659 (N_15659,N_15453,N_15326);
xnor U15660 (N_15660,N_15437,N_15357);
or U15661 (N_15661,N_15301,N_15357);
and U15662 (N_15662,N_15316,N_15311);
and U15663 (N_15663,N_15474,N_15345);
nor U15664 (N_15664,N_15374,N_15298);
nand U15665 (N_15665,N_15389,N_15395);
nor U15666 (N_15666,N_15341,N_15296);
or U15667 (N_15667,N_15259,N_15377);
nor U15668 (N_15668,N_15334,N_15313);
or U15669 (N_15669,N_15323,N_15347);
xor U15670 (N_15670,N_15296,N_15376);
and U15671 (N_15671,N_15285,N_15451);
or U15672 (N_15672,N_15261,N_15473);
xor U15673 (N_15673,N_15315,N_15407);
or U15674 (N_15674,N_15487,N_15341);
nor U15675 (N_15675,N_15409,N_15324);
nor U15676 (N_15676,N_15353,N_15320);
nor U15677 (N_15677,N_15285,N_15419);
or U15678 (N_15678,N_15342,N_15393);
nor U15679 (N_15679,N_15324,N_15297);
or U15680 (N_15680,N_15264,N_15368);
nand U15681 (N_15681,N_15490,N_15370);
nand U15682 (N_15682,N_15307,N_15337);
or U15683 (N_15683,N_15491,N_15395);
nor U15684 (N_15684,N_15369,N_15311);
or U15685 (N_15685,N_15330,N_15373);
xor U15686 (N_15686,N_15252,N_15318);
nand U15687 (N_15687,N_15278,N_15472);
nor U15688 (N_15688,N_15348,N_15449);
nand U15689 (N_15689,N_15382,N_15475);
nor U15690 (N_15690,N_15399,N_15483);
nor U15691 (N_15691,N_15254,N_15296);
or U15692 (N_15692,N_15434,N_15480);
nor U15693 (N_15693,N_15457,N_15381);
and U15694 (N_15694,N_15430,N_15254);
or U15695 (N_15695,N_15278,N_15467);
nor U15696 (N_15696,N_15461,N_15409);
and U15697 (N_15697,N_15279,N_15267);
xor U15698 (N_15698,N_15263,N_15371);
and U15699 (N_15699,N_15354,N_15490);
or U15700 (N_15700,N_15393,N_15417);
nor U15701 (N_15701,N_15322,N_15450);
nor U15702 (N_15702,N_15413,N_15281);
xnor U15703 (N_15703,N_15434,N_15391);
or U15704 (N_15704,N_15257,N_15276);
xor U15705 (N_15705,N_15263,N_15485);
xor U15706 (N_15706,N_15420,N_15279);
nand U15707 (N_15707,N_15477,N_15450);
and U15708 (N_15708,N_15271,N_15490);
xnor U15709 (N_15709,N_15354,N_15391);
nor U15710 (N_15710,N_15364,N_15280);
nor U15711 (N_15711,N_15444,N_15313);
or U15712 (N_15712,N_15420,N_15432);
nand U15713 (N_15713,N_15261,N_15253);
and U15714 (N_15714,N_15373,N_15307);
or U15715 (N_15715,N_15413,N_15344);
or U15716 (N_15716,N_15393,N_15253);
or U15717 (N_15717,N_15330,N_15349);
or U15718 (N_15718,N_15271,N_15408);
and U15719 (N_15719,N_15472,N_15474);
and U15720 (N_15720,N_15433,N_15499);
nor U15721 (N_15721,N_15280,N_15286);
nor U15722 (N_15722,N_15270,N_15294);
nor U15723 (N_15723,N_15390,N_15472);
or U15724 (N_15724,N_15320,N_15444);
nor U15725 (N_15725,N_15434,N_15264);
nor U15726 (N_15726,N_15266,N_15277);
and U15727 (N_15727,N_15405,N_15341);
xor U15728 (N_15728,N_15446,N_15298);
nand U15729 (N_15729,N_15400,N_15279);
nand U15730 (N_15730,N_15289,N_15295);
and U15731 (N_15731,N_15380,N_15260);
nand U15732 (N_15732,N_15362,N_15432);
and U15733 (N_15733,N_15348,N_15446);
and U15734 (N_15734,N_15442,N_15322);
nor U15735 (N_15735,N_15366,N_15485);
nand U15736 (N_15736,N_15374,N_15442);
nor U15737 (N_15737,N_15460,N_15331);
or U15738 (N_15738,N_15416,N_15464);
or U15739 (N_15739,N_15341,N_15353);
or U15740 (N_15740,N_15334,N_15478);
nor U15741 (N_15741,N_15434,N_15449);
or U15742 (N_15742,N_15475,N_15319);
or U15743 (N_15743,N_15310,N_15457);
xnor U15744 (N_15744,N_15489,N_15475);
and U15745 (N_15745,N_15356,N_15486);
and U15746 (N_15746,N_15294,N_15253);
and U15747 (N_15747,N_15467,N_15406);
and U15748 (N_15748,N_15499,N_15274);
and U15749 (N_15749,N_15301,N_15294);
xnor U15750 (N_15750,N_15539,N_15736);
nand U15751 (N_15751,N_15708,N_15711);
xor U15752 (N_15752,N_15667,N_15635);
nor U15753 (N_15753,N_15664,N_15558);
nand U15754 (N_15754,N_15570,N_15716);
nand U15755 (N_15755,N_15593,N_15526);
and U15756 (N_15756,N_15617,N_15553);
xor U15757 (N_15757,N_15659,N_15724);
or U15758 (N_15758,N_15655,N_15612);
nand U15759 (N_15759,N_15505,N_15685);
xor U15760 (N_15760,N_15529,N_15639);
nand U15761 (N_15761,N_15517,N_15583);
xor U15762 (N_15762,N_15504,N_15695);
nand U15763 (N_15763,N_15707,N_15693);
xor U15764 (N_15764,N_15599,N_15706);
or U15765 (N_15765,N_15637,N_15531);
xor U15766 (N_15766,N_15748,N_15523);
or U15767 (N_15767,N_15646,N_15564);
or U15768 (N_15768,N_15611,N_15532);
xnor U15769 (N_15769,N_15502,N_15710);
or U15770 (N_15770,N_15568,N_15730);
nand U15771 (N_15771,N_15731,N_15616);
and U15772 (N_15772,N_15641,N_15687);
nor U15773 (N_15773,N_15729,N_15740);
nand U15774 (N_15774,N_15520,N_15511);
and U15775 (N_15775,N_15737,N_15661);
and U15776 (N_15776,N_15585,N_15521);
nor U15777 (N_15777,N_15565,N_15647);
nand U15778 (N_15778,N_15733,N_15645);
and U15779 (N_15779,N_15545,N_15668);
nor U15780 (N_15780,N_15572,N_15590);
and U15781 (N_15781,N_15522,N_15717);
nand U15782 (N_15782,N_15549,N_15606);
xor U15783 (N_15783,N_15671,N_15663);
or U15784 (N_15784,N_15614,N_15629);
and U15785 (N_15785,N_15584,N_15578);
nor U15786 (N_15786,N_15676,N_15747);
xor U15787 (N_15787,N_15556,N_15746);
or U15788 (N_15788,N_15686,N_15688);
nor U15789 (N_15789,N_15591,N_15588);
or U15790 (N_15790,N_15527,N_15550);
nor U15791 (N_15791,N_15613,N_15709);
and U15792 (N_15792,N_15609,N_15749);
nor U15793 (N_15793,N_15538,N_15597);
nand U15794 (N_15794,N_15742,N_15734);
and U15795 (N_15795,N_15623,N_15620);
xnor U15796 (N_15796,N_15683,N_15607);
nand U15797 (N_15797,N_15712,N_15579);
nor U15798 (N_15798,N_15547,N_15682);
or U15799 (N_15799,N_15662,N_15563);
nand U15800 (N_15800,N_15700,N_15721);
nand U15801 (N_15801,N_15500,N_15725);
or U15802 (N_15802,N_15560,N_15622);
and U15803 (N_15803,N_15626,N_15543);
nand U15804 (N_15804,N_15628,N_15503);
or U15805 (N_15805,N_15510,N_15632);
and U15806 (N_15806,N_15694,N_15670);
and U15807 (N_15807,N_15516,N_15648);
or U15808 (N_15808,N_15665,N_15720);
or U15809 (N_15809,N_15586,N_15743);
nand U15810 (N_15810,N_15652,N_15719);
nand U15811 (N_15811,N_15684,N_15644);
xnor U15812 (N_15812,N_15513,N_15714);
xor U15813 (N_15813,N_15643,N_15501);
or U15814 (N_15814,N_15675,N_15554);
or U15815 (N_15815,N_15696,N_15574);
xnor U15816 (N_15816,N_15669,N_15602);
nor U15817 (N_15817,N_15515,N_15530);
or U15818 (N_15818,N_15656,N_15638);
and U15819 (N_15819,N_15557,N_15608);
nor U15820 (N_15820,N_15519,N_15535);
or U15821 (N_15821,N_15533,N_15544);
and U15822 (N_15822,N_15571,N_15598);
xnor U15823 (N_15823,N_15534,N_15735);
and U15824 (N_15824,N_15744,N_15703);
and U15825 (N_15825,N_15698,N_15567);
and U15826 (N_15826,N_15536,N_15555);
xnor U15827 (N_15827,N_15601,N_15634);
nand U15828 (N_15828,N_15559,N_15651);
xnor U15829 (N_15829,N_15605,N_15594);
xnor U15830 (N_15830,N_15587,N_15576);
nor U15831 (N_15831,N_15658,N_15745);
xor U15832 (N_15832,N_15525,N_15580);
nor U15833 (N_15833,N_15689,N_15615);
nand U15834 (N_15834,N_15630,N_15723);
or U15835 (N_15835,N_15596,N_15577);
nor U15836 (N_15836,N_15581,N_15713);
and U15837 (N_15837,N_15618,N_15739);
or U15838 (N_15838,N_15702,N_15681);
nor U15839 (N_15839,N_15672,N_15528);
xor U15840 (N_15840,N_15573,N_15705);
and U15841 (N_15841,N_15624,N_15540);
xnor U15842 (N_15842,N_15506,N_15625);
or U15843 (N_15843,N_15569,N_15589);
nand U15844 (N_15844,N_15690,N_15582);
nand U15845 (N_15845,N_15562,N_15509);
nand U15846 (N_15846,N_15619,N_15657);
nand U15847 (N_15847,N_15701,N_15518);
xnor U15848 (N_15848,N_15697,N_15722);
nor U15849 (N_15849,N_15514,N_15603);
nand U15850 (N_15850,N_15566,N_15726);
xor U15851 (N_15851,N_15512,N_15537);
and U15852 (N_15852,N_15699,N_15649);
xor U15853 (N_15853,N_15674,N_15715);
nor U15854 (N_15854,N_15524,N_15631);
nand U15855 (N_15855,N_15633,N_15718);
xnor U15856 (N_15856,N_15621,N_15741);
nand U15857 (N_15857,N_15679,N_15610);
xnor U15858 (N_15858,N_15541,N_15738);
nand U15859 (N_15859,N_15592,N_15636);
xnor U15860 (N_15860,N_15650,N_15546);
nand U15861 (N_15861,N_15508,N_15666);
nand U15862 (N_15862,N_15728,N_15600);
or U15863 (N_15863,N_15542,N_15551);
nor U15864 (N_15864,N_15548,N_15552);
nor U15865 (N_15865,N_15654,N_15732);
nor U15866 (N_15866,N_15604,N_15640);
nor U15867 (N_15867,N_15627,N_15677);
nand U15868 (N_15868,N_15727,N_15595);
nand U15869 (N_15869,N_15673,N_15653);
nor U15870 (N_15870,N_15642,N_15575);
nand U15871 (N_15871,N_15660,N_15680);
and U15872 (N_15872,N_15561,N_15692);
nand U15873 (N_15873,N_15678,N_15507);
xnor U15874 (N_15874,N_15691,N_15704);
nor U15875 (N_15875,N_15727,N_15636);
nand U15876 (N_15876,N_15506,N_15621);
nor U15877 (N_15877,N_15582,N_15571);
nand U15878 (N_15878,N_15692,N_15568);
or U15879 (N_15879,N_15603,N_15709);
xnor U15880 (N_15880,N_15559,N_15568);
nand U15881 (N_15881,N_15520,N_15746);
nand U15882 (N_15882,N_15586,N_15645);
nand U15883 (N_15883,N_15584,N_15704);
xnor U15884 (N_15884,N_15713,N_15540);
or U15885 (N_15885,N_15618,N_15748);
nand U15886 (N_15886,N_15584,N_15732);
nor U15887 (N_15887,N_15611,N_15721);
nor U15888 (N_15888,N_15539,N_15510);
nor U15889 (N_15889,N_15706,N_15542);
and U15890 (N_15890,N_15692,N_15716);
nand U15891 (N_15891,N_15617,N_15527);
nor U15892 (N_15892,N_15509,N_15576);
or U15893 (N_15893,N_15713,N_15511);
nand U15894 (N_15894,N_15611,N_15561);
and U15895 (N_15895,N_15742,N_15518);
nand U15896 (N_15896,N_15747,N_15649);
and U15897 (N_15897,N_15547,N_15636);
nand U15898 (N_15898,N_15514,N_15600);
and U15899 (N_15899,N_15714,N_15641);
xor U15900 (N_15900,N_15698,N_15593);
xor U15901 (N_15901,N_15660,N_15612);
or U15902 (N_15902,N_15650,N_15561);
xnor U15903 (N_15903,N_15607,N_15568);
or U15904 (N_15904,N_15682,N_15734);
nor U15905 (N_15905,N_15722,N_15567);
and U15906 (N_15906,N_15721,N_15649);
xor U15907 (N_15907,N_15638,N_15725);
and U15908 (N_15908,N_15655,N_15553);
and U15909 (N_15909,N_15573,N_15517);
xor U15910 (N_15910,N_15689,N_15698);
and U15911 (N_15911,N_15530,N_15610);
nor U15912 (N_15912,N_15669,N_15605);
nand U15913 (N_15913,N_15568,N_15509);
nand U15914 (N_15914,N_15629,N_15579);
nand U15915 (N_15915,N_15668,N_15739);
xnor U15916 (N_15916,N_15595,N_15502);
xor U15917 (N_15917,N_15685,N_15524);
nand U15918 (N_15918,N_15647,N_15691);
nand U15919 (N_15919,N_15588,N_15681);
xor U15920 (N_15920,N_15519,N_15599);
nand U15921 (N_15921,N_15592,N_15660);
nand U15922 (N_15922,N_15620,N_15683);
or U15923 (N_15923,N_15746,N_15604);
and U15924 (N_15924,N_15621,N_15690);
or U15925 (N_15925,N_15538,N_15550);
and U15926 (N_15926,N_15576,N_15719);
nand U15927 (N_15927,N_15524,N_15689);
or U15928 (N_15928,N_15614,N_15579);
and U15929 (N_15929,N_15703,N_15528);
nor U15930 (N_15930,N_15638,N_15661);
nand U15931 (N_15931,N_15599,N_15674);
nor U15932 (N_15932,N_15675,N_15550);
nand U15933 (N_15933,N_15538,N_15594);
nor U15934 (N_15934,N_15672,N_15612);
and U15935 (N_15935,N_15606,N_15660);
and U15936 (N_15936,N_15565,N_15711);
nor U15937 (N_15937,N_15746,N_15614);
or U15938 (N_15938,N_15544,N_15517);
xor U15939 (N_15939,N_15649,N_15542);
xor U15940 (N_15940,N_15742,N_15515);
nor U15941 (N_15941,N_15682,N_15736);
xnor U15942 (N_15942,N_15748,N_15545);
nor U15943 (N_15943,N_15694,N_15681);
or U15944 (N_15944,N_15720,N_15639);
and U15945 (N_15945,N_15749,N_15583);
or U15946 (N_15946,N_15642,N_15606);
and U15947 (N_15947,N_15718,N_15667);
nand U15948 (N_15948,N_15711,N_15724);
or U15949 (N_15949,N_15746,N_15555);
nor U15950 (N_15950,N_15610,N_15519);
or U15951 (N_15951,N_15714,N_15741);
nor U15952 (N_15952,N_15640,N_15728);
and U15953 (N_15953,N_15708,N_15678);
xnor U15954 (N_15954,N_15641,N_15594);
xor U15955 (N_15955,N_15616,N_15570);
xor U15956 (N_15956,N_15580,N_15676);
and U15957 (N_15957,N_15731,N_15584);
nand U15958 (N_15958,N_15630,N_15600);
or U15959 (N_15959,N_15531,N_15599);
or U15960 (N_15960,N_15510,N_15687);
or U15961 (N_15961,N_15627,N_15516);
xnor U15962 (N_15962,N_15695,N_15714);
or U15963 (N_15963,N_15745,N_15563);
and U15964 (N_15964,N_15683,N_15616);
and U15965 (N_15965,N_15532,N_15615);
or U15966 (N_15966,N_15663,N_15652);
xnor U15967 (N_15967,N_15540,N_15737);
or U15968 (N_15968,N_15557,N_15628);
nand U15969 (N_15969,N_15724,N_15627);
xor U15970 (N_15970,N_15698,N_15635);
and U15971 (N_15971,N_15529,N_15667);
nor U15972 (N_15972,N_15587,N_15604);
or U15973 (N_15973,N_15531,N_15628);
and U15974 (N_15974,N_15657,N_15749);
nor U15975 (N_15975,N_15521,N_15563);
nor U15976 (N_15976,N_15542,N_15605);
nand U15977 (N_15977,N_15713,N_15634);
or U15978 (N_15978,N_15623,N_15527);
nand U15979 (N_15979,N_15688,N_15736);
nand U15980 (N_15980,N_15507,N_15502);
xnor U15981 (N_15981,N_15732,N_15592);
nor U15982 (N_15982,N_15631,N_15732);
nor U15983 (N_15983,N_15590,N_15681);
and U15984 (N_15984,N_15660,N_15582);
and U15985 (N_15985,N_15666,N_15512);
xor U15986 (N_15986,N_15650,N_15645);
xnor U15987 (N_15987,N_15500,N_15597);
nand U15988 (N_15988,N_15553,N_15741);
and U15989 (N_15989,N_15673,N_15524);
nor U15990 (N_15990,N_15564,N_15544);
nand U15991 (N_15991,N_15708,N_15516);
nor U15992 (N_15992,N_15528,N_15732);
or U15993 (N_15993,N_15714,N_15579);
and U15994 (N_15994,N_15649,N_15520);
and U15995 (N_15995,N_15675,N_15589);
nor U15996 (N_15996,N_15592,N_15524);
or U15997 (N_15997,N_15724,N_15658);
nand U15998 (N_15998,N_15572,N_15630);
and U15999 (N_15999,N_15612,N_15677);
and U16000 (N_16000,N_15966,N_15939);
and U16001 (N_16001,N_15963,N_15832);
nand U16002 (N_16002,N_15813,N_15975);
xor U16003 (N_16003,N_15753,N_15779);
nor U16004 (N_16004,N_15843,N_15822);
and U16005 (N_16005,N_15752,N_15994);
xnor U16006 (N_16006,N_15866,N_15848);
xor U16007 (N_16007,N_15911,N_15785);
xor U16008 (N_16008,N_15996,N_15930);
and U16009 (N_16009,N_15760,N_15825);
and U16010 (N_16010,N_15829,N_15772);
or U16011 (N_16011,N_15956,N_15949);
nor U16012 (N_16012,N_15835,N_15915);
and U16013 (N_16013,N_15921,N_15762);
or U16014 (N_16014,N_15984,N_15831);
or U16015 (N_16015,N_15877,N_15993);
xor U16016 (N_16016,N_15981,N_15796);
and U16017 (N_16017,N_15790,N_15937);
or U16018 (N_16018,N_15952,N_15839);
nor U16019 (N_16019,N_15973,N_15924);
nand U16020 (N_16020,N_15859,N_15869);
nor U16021 (N_16021,N_15820,N_15938);
xnor U16022 (N_16022,N_15857,N_15935);
nor U16023 (N_16023,N_15983,N_15929);
nor U16024 (N_16024,N_15936,N_15765);
and U16025 (N_16025,N_15844,N_15786);
xor U16026 (N_16026,N_15957,N_15814);
and U16027 (N_16027,N_15858,N_15971);
and U16028 (N_16028,N_15992,N_15799);
nor U16029 (N_16029,N_15985,N_15978);
nor U16030 (N_16030,N_15912,N_15826);
xnor U16031 (N_16031,N_15806,N_15932);
xor U16032 (N_16032,N_15933,N_15775);
xnor U16033 (N_16033,N_15898,N_15905);
or U16034 (N_16034,N_15886,N_15865);
nand U16035 (N_16035,N_15754,N_15809);
or U16036 (N_16036,N_15855,N_15900);
nor U16037 (N_16037,N_15884,N_15890);
nor U16038 (N_16038,N_15766,N_15888);
nand U16039 (N_16039,N_15876,N_15962);
xor U16040 (N_16040,N_15852,N_15879);
nor U16041 (N_16041,N_15934,N_15986);
nand U16042 (N_16042,N_15910,N_15816);
and U16043 (N_16043,N_15927,N_15802);
and U16044 (N_16044,N_15803,N_15953);
and U16045 (N_16045,N_15926,N_15794);
xor U16046 (N_16046,N_15868,N_15955);
nand U16047 (N_16047,N_15977,N_15842);
or U16048 (N_16048,N_15959,N_15928);
xnor U16049 (N_16049,N_15761,N_15811);
nor U16050 (N_16050,N_15787,N_15968);
nand U16051 (N_16051,N_15836,N_15894);
or U16052 (N_16052,N_15818,N_15960);
or U16053 (N_16053,N_15948,N_15906);
xor U16054 (N_16054,N_15770,N_15941);
xor U16055 (N_16055,N_15798,N_15828);
and U16056 (N_16056,N_15834,N_15807);
or U16057 (N_16057,N_15789,N_15970);
nand U16058 (N_16058,N_15768,N_15998);
and U16059 (N_16059,N_15864,N_15942);
nor U16060 (N_16060,N_15860,N_15874);
and U16061 (N_16061,N_15817,N_15819);
and U16062 (N_16062,N_15919,N_15950);
or U16063 (N_16063,N_15861,N_15883);
xnor U16064 (N_16064,N_15782,N_15997);
nand U16065 (N_16065,N_15792,N_15778);
nand U16066 (N_16066,N_15914,N_15922);
nor U16067 (N_16067,N_15751,N_15812);
nor U16068 (N_16068,N_15882,N_15870);
and U16069 (N_16069,N_15849,N_15947);
nand U16070 (N_16070,N_15943,N_15885);
or U16071 (N_16071,N_15946,N_15856);
xnor U16072 (N_16072,N_15989,N_15951);
nand U16073 (N_16073,N_15873,N_15773);
nand U16074 (N_16074,N_15815,N_15776);
xor U16075 (N_16075,N_15784,N_15824);
nand U16076 (N_16076,N_15783,N_15974);
xnor U16077 (N_16077,N_15777,N_15845);
and U16078 (N_16078,N_15801,N_15899);
or U16079 (N_16079,N_15823,N_15850);
nor U16080 (N_16080,N_15954,N_15780);
nor U16081 (N_16081,N_15895,N_15755);
nand U16082 (N_16082,N_15764,N_15756);
nor U16083 (N_16083,N_15918,N_15931);
nand U16084 (N_16084,N_15917,N_15995);
xnor U16085 (N_16085,N_15804,N_15800);
xor U16086 (N_16086,N_15797,N_15944);
xnor U16087 (N_16087,N_15774,N_15880);
nor U16088 (N_16088,N_15923,N_15907);
and U16089 (N_16089,N_15808,N_15972);
or U16090 (N_16090,N_15925,N_15990);
or U16091 (N_16091,N_15838,N_15988);
xnor U16092 (N_16092,N_15889,N_15969);
and U16093 (N_16093,N_15940,N_15961);
nor U16094 (N_16094,N_15976,N_15872);
nor U16095 (N_16095,N_15902,N_15891);
xor U16096 (N_16096,N_15805,N_15887);
nand U16097 (N_16097,N_15758,N_15833);
xnor U16098 (N_16098,N_15901,N_15987);
nor U16099 (N_16099,N_15965,N_15904);
nand U16100 (N_16100,N_15903,N_15771);
nand U16101 (N_16101,N_15863,N_15827);
and U16102 (N_16102,N_15875,N_15945);
and U16103 (N_16103,N_15908,N_15847);
and U16104 (N_16104,N_15913,N_15867);
nand U16105 (N_16105,N_15871,N_15896);
and U16106 (N_16106,N_15892,N_15759);
xnor U16107 (N_16107,N_15846,N_15881);
nor U16108 (N_16108,N_15893,N_15979);
nand U16109 (N_16109,N_15757,N_15878);
xor U16110 (N_16110,N_15810,N_15795);
or U16111 (N_16111,N_15853,N_15967);
nand U16112 (N_16112,N_15982,N_15763);
xnor U16113 (N_16113,N_15980,N_15999);
nor U16114 (N_16114,N_15821,N_15840);
nand U16115 (N_16115,N_15781,N_15837);
nand U16116 (N_16116,N_15851,N_15854);
and U16117 (N_16117,N_15767,N_15750);
or U16118 (N_16118,N_15958,N_15909);
xnor U16119 (N_16119,N_15964,N_15841);
and U16120 (N_16120,N_15791,N_15769);
nor U16121 (N_16121,N_15862,N_15793);
or U16122 (N_16122,N_15916,N_15788);
or U16123 (N_16123,N_15991,N_15920);
nand U16124 (N_16124,N_15830,N_15897);
nor U16125 (N_16125,N_15867,N_15791);
and U16126 (N_16126,N_15947,N_15959);
xor U16127 (N_16127,N_15993,N_15977);
nor U16128 (N_16128,N_15993,N_15869);
nor U16129 (N_16129,N_15806,N_15776);
and U16130 (N_16130,N_15857,N_15791);
or U16131 (N_16131,N_15988,N_15978);
and U16132 (N_16132,N_15932,N_15976);
and U16133 (N_16133,N_15858,N_15831);
nor U16134 (N_16134,N_15822,N_15891);
or U16135 (N_16135,N_15889,N_15809);
nor U16136 (N_16136,N_15947,N_15750);
and U16137 (N_16137,N_15964,N_15806);
and U16138 (N_16138,N_15965,N_15833);
xor U16139 (N_16139,N_15999,N_15900);
nand U16140 (N_16140,N_15971,N_15802);
and U16141 (N_16141,N_15871,N_15772);
and U16142 (N_16142,N_15799,N_15884);
nand U16143 (N_16143,N_15845,N_15832);
nand U16144 (N_16144,N_15960,N_15981);
and U16145 (N_16145,N_15825,N_15872);
or U16146 (N_16146,N_15836,N_15785);
nand U16147 (N_16147,N_15775,N_15783);
or U16148 (N_16148,N_15907,N_15788);
nor U16149 (N_16149,N_15878,N_15793);
and U16150 (N_16150,N_15990,N_15959);
nand U16151 (N_16151,N_15956,N_15878);
nor U16152 (N_16152,N_15950,N_15954);
or U16153 (N_16153,N_15927,N_15884);
and U16154 (N_16154,N_15815,N_15778);
or U16155 (N_16155,N_15867,N_15898);
or U16156 (N_16156,N_15801,N_15843);
or U16157 (N_16157,N_15932,N_15934);
nor U16158 (N_16158,N_15988,N_15756);
and U16159 (N_16159,N_15826,N_15899);
nor U16160 (N_16160,N_15934,N_15823);
nand U16161 (N_16161,N_15775,N_15921);
or U16162 (N_16162,N_15818,N_15999);
nor U16163 (N_16163,N_15908,N_15799);
xor U16164 (N_16164,N_15988,N_15982);
or U16165 (N_16165,N_15798,N_15961);
nor U16166 (N_16166,N_15872,N_15993);
nor U16167 (N_16167,N_15959,N_15783);
and U16168 (N_16168,N_15936,N_15872);
or U16169 (N_16169,N_15817,N_15935);
or U16170 (N_16170,N_15975,N_15765);
nand U16171 (N_16171,N_15840,N_15778);
nand U16172 (N_16172,N_15865,N_15968);
xor U16173 (N_16173,N_15997,N_15905);
nand U16174 (N_16174,N_15922,N_15754);
and U16175 (N_16175,N_15954,N_15751);
nand U16176 (N_16176,N_15899,N_15882);
or U16177 (N_16177,N_15883,N_15782);
and U16178 (N_16178,N_15977,N_15902);
or U16179 (N_16179,N_15767,N_15818);
nor U16180 (N_16180,N_15804,N_15939);
or U16181 (N_16181,N_15921,N_15848);
nand U16182 (N_16182,N_15963,N_15851);
nand U16183 (N_16183,N_15785,N_15879);
and U16184 (N_16184,N_15956,N_15928);
xor U16185 (N_16185,N_15782,N_15780);
or U16186 (N_16186,N_15789,N_15784);
and U16187 (N_16187,N_15805,N_15837);
xor U16188 (N_16188,N_15886,N_15842);
or U16189 (N_16189,N_15830,N_15790);
and U16190 (N_16190,N_15915,N_15845);
and U16191 (N_16191,N_15952,N_15940);
nand U16192 (N_16192,N_15793,N_15775);
nor U16193 (N_16193,N_15983,N_15951);
and U16194 (N_16194,N_15754,N_15762);
nand U16195 (N_16195,N_15776,N_15886);
nor U16196 (N_16196,N_15865,N_15970);
nand U16197 (N_16197,N_15987,N_15895);
nor U16198 (N_16198,N_15769,N_15792);
nor U16199 (N_16199,N_15898,N_15841);
and U16200 (N_16200,N_15975,N_15893);
and U16201 (N_16201,N_15925,N_15943);
or U16202 (N_16202,N_15857,N_15940);
nor U16203 (N_16203,N_15785,N_15799);
nor U16204 (N_16204,N_15998,N_15798);
nor U16205 (N_16205,N_15762,N_15827);
or U16206 (N_16206,N_15832,N_15755);
nand U16207 (N_16207,N_15935,N_15932);
nand U16208 (N_16208,N_15937,N_15752);
xnor U16209 (N_16209,N_15884,N_15839);
xor U16210 (N_16210,N_15957,N_15938);
and U16211 (N_16211,N_15819,N_15911);
nor U16212 (N_16212,N_15811,N_15870);
or U16213 (N_16213,N_15947,N_15916);
nand U16214 (N_16214,N_15995,N_15993);
or U16215 (N_16215,N_15774,N_15781);
nand U16216 (N_16216,N_15961,N_15973);
and U16217 (N_16217,N_15765,N_15850);
and U16218 (N_16218,N_15892,N_15978);
nand U16219 (N_16219,N_15975,N_15929);
and U16220 (N_16220,N_15901,N_15945);
xor U16221 (N_16221,N_15852,N_15976);
nor U16222 (N_16222,N_15871,N_15913);
nand U16223 (N_16223,N_15778,N_15952);
nand U16224 (N_16224,N_15929,N_15985);
xor U16225 (N_16225,N_15955,N_15789);
xnor U16226 (N_16226,N_15896,N_15884);
nor U16227 (N_16227,N_15816,N_15817);
nor U16228 (N_16228,N_15919,N_15968);
xor U16229 (N_16229,N_15857,N_15821);
xor U16230 (N_16230,N_15962,N_15890);
nor U16231 (N_16231,N_15817,N_15881);
nand U16232 (N_16232,N_15825,N_15895);
or U16233 (N_16233,N_15760,N_15919);
or U16234 (N_16234,N_15834,N_15963);
nand U16235 (N_16235,N_15755,N_15961);
or U16236 (N_16236,N_15780,N_15795);
and U16237 (N_16237,N_15825,N_15898);
xor U16238 (N_16238,N_15803,N_15756);
xor U16239 (N_16239,N_15913,N_15805);
nand U16240 (N_16240,N_15963,N_15844);
xor U16241 (N_16241,N_15933,N_15987);
xnor U16242 (N_16242,N_15868,N_15750);
nor U16243 (N_16243,N_15839,N_15984);
and U16244 (N_16244,N_15918,N_15920);
xor U16245 (N_16245,N_15913,N_15986);
or U16246 (N_16246,N_15783,N_15976);
and U16247 (N_16247,N_15820,N_15826);
nor U16248 (N_16248,N_15803,N_15847);
nand U16249 (N_16249,N_15886,N_15940);
and U16250 (N_16250,N_16073,N_16154);
xor U16251 (N_16251,N_16080,N_16146);
and U16252 (N_16252,N_16204,N_16035);
nor U16253 (N_16253,N_16195,N_16147);
and U16254 (N_16254,N_16017,N_16007);
xnor U16255 (N_16255,N_16177,N_16236);
or U16256 (N_16256,N_16166,N_16156);
nor U16257 (N_16257,N_16019,N_16002);
or U16258 (N_16258,N_16003,N_16091);
nand U16259 (N_16259,N_16135,N_16041);
xor U16260 (N_16260,N_16130,N_16153);
nor U16261 (N_16261,N_16123,N_16067);
nand U16262 (N_16262,N_16132,N_16056);
and U16263 (N_16263,N_16125,N_16114);
or U16264 (N_16264,N_16223,N_16097);
or U16265 (N_16265,N_16072,N_16136);
nor U16266 (N_16266,N_16093,N_16060);
and U16267 (N_16267,N_16138,N_16043);
nor U16268 (N_16268,N_16233,N_16157);
and U16269 (N_16269,N_16065,N_16026);
xor U16270 (N_16270,N_16165,N_16163);
xnor U16271 (N_16271,N_16249,N_16189);
xor U16272 (N_16272,N_16109,N_16052);
or U16273 (N_16273,N_16042,N_16243);
or U16274 (N_16274,N_16103,N_16063);
nor U16275 (N_16275,N_16004,N_16092);
nor U16276 (N_16276,N_16222,N_16010);
or U16277 (N_16277,N_16182,N_16173);
or U16278 (N_16278,N_16142,N_16078);
nor U16279 (N_16279,N_16225,N_16240);
nor U16280 (N_16280,N_16082,N_16169);
nor U16281 (N_16281,N_16047,N_16158);
or U16282 (N_16282,N_16176,N_16029);
xnor U16283 (N_16283,N_16190,N_16014);
or U16284 (N_16284,N_16149,N_16016);
nor U16285 (N_16285,N_16025,N_16087);
or U16286 (N_16286,N_16127,N_16085);
nor U16287 (N_16287,N_16232,N_16167);
and U16288 (N_16288,N_16077,N_16148);
or U16289 (N_16289,N_16234,N_16124);
nand U16290 (N_16290,N_16180,N_16044);
nor U16291 (N_16291,N_16074,N_16079);
nand U16292 (N_16292,N_16113,N_16241);
xor U16293 (N_16293,N_16219,N_16096);
nor U16294 (N_16294,N_16160,N_16203);
and U16295 (N_16295,N_16140,N_16066);
nand U16296 (N_16296,N_16213,N_16058);
or U16297 (N_16297,N_16128,N_16107);
or U16298 (N_16298,N_16202,N_16133);
xnor U16299 (N_16299,N_16245,N_16178);
nor U16300 (N_16300,N_16118,N_16229);
and U16301 (N_16301,N_16030,N_16231);
xor U16302 (N_16302,N_16089,N_16151);
xor U16303 (N_16303,N_16012,N_16199);
nor U16304 (N_16304,N_16183,N_16120);
or U16305 (N_16305,N_16221,N_16186);
nand U16306 (N_16306,N_16001,N_16244);
and U16307 (N_16307,N_16020,N_16101);
nand U16308 (N_16308,N_16045,N_16054);
or U16309 (N_16309,N_16239,N_16179);
nand U16310 (N_16310,N_16242,N_16110);
or U16311 (N_16311,N_16216,N_16106);
nand U16312 (N_16312,N_16238,N_16137);
nor U16313 (N_16313,N_16129,N_16039);
xnor U16314 (N_16314,N_16011,N_16055);
xor U16315 (N_16315,N_16100,N_16064);
nand U16316 (N_16316,N_16168,N_16036);
xnor U16317 (N_16317,N_16134,N_16115);
and U16318 (N_16318,N_16246,N_16040);
nand U16319 (N_16319,N_16224,N_16227);
nand U16320 (N_16320,N_16145,N_16088);
nor U16321 (N_16321,N_16230,N_16150);
xor U16322 (N_16322,N_16068,N_16126);
and U16323 (N_16323,N_16211,N_16018);
and U16324 (N_16324,N_16198,N_16009);
or U16325 (N_16325,N_16184,N_16038);
nor U16326 (N_16326,N_16164,N_16000);
xor U16327 (N_16327,N_16141,N_16108);
nor U16328 (N_16328,N_16059,N_16116);
and U16329 (N_16329,N_16021,N_16215);
or U16330 (N_16330,N_16105,N_16152);
or U16331 (N_16331,N_16122,N_16139);
and U16332 (N_16332,N_16049,N_16005);
and U16333 (N_16333,N_16172,N_16194);
nand U16334 (N_16334,N_16237,N_16181);
and U16335 (N_16335,N_16171,N_16174);
and U16336 (N_16336,N_16062,N_16048);
or U16337 (N_16337,N_16095,N_16143);
xor U16338 (N_16338,N_16117,N_16193);
nand U16339 (N_16339,N_16031,N_16013);
or U16340 (N_16340,N_16015,N_16144);
xor U16341 (N_16341,N_16188,N_16076);
nor U16342 (N_16342,N_16191,N_16070);
and U16343 (N_16343,N_16061,N_16083);
nor U16344 (N_16344,N_16104,N_16081);
nor U16345 (N_16345,N_16196,N_16170);
and U16346 (N_16346,N_16159,N_16205);
or U16347 (N_16347,N_16226,N_16023);
xnor U16348 (N_16348,N_16155,N_16034);
xnor U16349 (N_16349,N_16094,N_16084);
nor U16350 (N_16350,N_16008,N_16247);
or U16351 (N_16351,N_16071,N_16112);
nand U16352 (N_16352,N_16032,N_16098);
and U16353 (N_16353,N_16027,N_16185);
nor U16354 (N_16354,N_16046,N_16050);
and U16355 (N_16355,N_16228,N_16053);
nor U16356 (N_16356,N_16131,N_16197);
xor U16357 (N_16357,N_16192,N_16121);
or U16358 (N_16358,N_16006,N_16209);
nand U16359 (N_16359,N_16162,N_16111);
or U16360 (N_16360,N_16075,N_16037);
nand U16361 (N_16361,N_16201,N_16069);
nand U16362 (N_16362,N_16086,N_16033);
or U16363 (N_16363,N_16200,N_16022);
xor U16364 (N_16364,N_16220,N_16161);
xnor U16365 (N_16365,N_16207,N_16051);
xnor U16366 (N_16366,N_16090,N_16206);
xor U16367 (N_16367,N_16218,N_16212);
or U16368 (N_16368,N_16187,N_16217);
or U16369 (N_16369,N_16214,N_16057);
nand U16370 (N_16370,N_16028,N_16102);
or U16371 (N_16371,N_16208,N_16210);
and U16372 (N_16372,N_16235,N_16024);
xnor U16373 (N_16373,N_16119,N_16175);
nand U16374 (N_16374,N_16099,N_16248);
or U16375 (N_16375,N_16097,N_16166);
xor U16376 (N_16376,N_16138,N_16102);
nor U16377 (N_16377,N_16006,N_16135);
nand U16378 (N_16378,N_16021,N_16111);
xor U16379 (N_16379,N_16188,N_16240);
nand U16380 (N_16380,N_16036,N_16046);
xnor U16381 (N_16381,N_16158,N_16235);
nor U16382 (N_16382,N_16193,N_16115);
and U16383 (N_16383,N_16047,N_16078);
and U16384 (N_16384,N_16048,N_16241);
or U16385 (N_16385,N_16043,N_16180);
nor U16386 (N_16386,N_16158,N_16187);
and U16387 (N_16387,N_16091,N_16217);
nor U16388 (N_16388,N_16101,N_16102);
or U16389 (N_16389,N_16069,N_16247);
nor U16390 (N_16390,N_16132,N_16110);
nor U16391 (N_16391,N_16106,N_16247);
or U16392 (N_16392,N_16084,N_16141);
nand U16393 (N_16393,N_16237,N_16183);
and U16394 (N_16394,N_16174,N_16014);
nand U16395 (N_16395,N_16249,N_16143);
nor U16396 (N_16396,N_16212,N_16055);
nand U16397 (N_16397,N_16239,N_16204);
or U16398 (N_16398,N_16166,N_16019);
or U16399 (N_16399,N_16096,N_16105);
or U16400 (N_16400,N_16092,N_16188);
nand U16401 (N_16401,N_16130,N_16161);
nand U16402 (N_16402,N_16019,N_16160);
and U16403 (N_16403,N_16213,N_16174);
nand U16404 (N_16404,N_16157,N_16187);
xnor U16405 (N_16405,N_16188,N_16033);
and U16406 (N_16406,N_16237,N_16005);
or U16407 (N_16407,N_16094,N_16093);
nor U16408 (N_16408,N_16103,N_16219);
nand U16409 (N_16409,N_16015,N_16042);
nand U16410 (N_16410,N_16155,N_16218);
and U16411 (N_16411,N_16210,N_16178);
and U16412 (N_16412,N_16044,N_16002);
xnor U16413 (N_16413,N_16223,N_16166);
or U16414 (N_16414,N_16143,N_16110);
or U16415 (N_16415,N_16065,N_16138);
nor U16416 (N_16416,N_16028,N_16040);
xor U16417 (N_16417,N_16243,N_16241);
xnor U16418 (N_16418,N_16031,N_16138);
xnor U16419 (N_16419,N_16005,N_16016);
xnor U16420 (N_16420,N_16040,N_16124);
nor U16421 (N_16421,N_16038,N_16144);
nand U16422 (N_16422,N_16033,N_16193);
nor U16423 (N_16423,N_16192,N_16181);
nand U16424 (N_16424,N_16149,N_16227);
and U16425 (N_16425,N_16085,N_16169);
or U16426 (N_16426,N_16020,N_16211);
or U16427 (N_16427,N_16247,N_16093);
nor U16428 (N_16428,N_16112,N_16057);
nor U16429 (N_16429,N_16110,N_16170);
nand U16430 (N_16430,N_16011,N_16203);
or U16431 (N_16431,N_16081,N_16145);
nor U16432 (N_16432,N_16132,N_16219);
nor U16433 (N_16433,N_16153,N_16232);
nor U16434 (N_16434,N_16084,N_16128);
xor U16435 (N_16435,N_16043,N_16183);
and U16436 (N_16436,N_16164,N_16092);
nor U16437 (N_16437,N_16006,N_16093);
nor U16438 (N_16438,N_16003,N_16248);
xor U16439 (N_16439,N_16220,N_16065);
nor U16440 (N_16440,N_16134,N_16249);
xor U16441 (N_16441,N_16146,N_16088);
or U16442 (N_16442,N_16081,N_16149);
nand U16443 (N_16443,N_16034,N_16071);
and U16444 (N_16444,N_16092,N_16078);
or U16445 (N_16445,N_16142,N_16023);
and U16446 (N_16446,N_16189,N_16030);
or U16447 (N_16447,N_16088,N_16218);
nand U16448 (N_16448,N_16041,N_16188);
and U16449 (N_16449,N_16069,N_16080);
or U16450 (N_16450,N_16130,N_16098);
and U16451 (N_16451,N_16066,N_16204);
xor U16452 (N_16452,N_16012,N_16011);
nor U16453 (N_16453,N_16072,N_16012);
nor U16454 (N_16454,N_16225,N_16227);
nand U16455 (N_16455,N_16044,N_16177);
or U16456 (N_16456,N_16139,N_16034);
nor U16457 (N_16457,N_16092,N_16006);
or U16458 (N_16458,N_16238,N_16003);
xor U16459 (N_16459,N_16206,N_16226);
and U16460 (N_16460,N_16091,N_16245);
xnor U16461 (N_16461,N_16034,N_16194);
xnor U16462 (N_16462,N_16215,N_16127);
nor U16463 (N_16463,N_16225,N_16209);
nor U16464 (N_16464,N_16014,N_16124);
or U16465 (N_16465,N_16025,N_16210);
nand U16466 (N_16466,N_16044,N_16010);
or U16467 (N_16467,N_16102,N_16199);
or U16468 (N_16468,N_16218,N_16085);
nand U16469 (N_16469,N_16021,N_16189);
nor U16470 (N_16470,N_16044,N_16117);
or U16471 (N_16471,N_16204,N_16201);
nor U16472 (N_16472,N_16123,N_16241);
xor U16473 (N_16473,N_16065,N_16015);
or U16474 (N_16474,N_16018,N_16135);
nor U16475 (N_16475,N_16148,N_16206);
nand U16476 (N_16476,N_16161,N_16218);
nand U16477 (N_16477,N_16122,N_16136);
nor U16478 (N_16478,N_16014,N_16144);
or U16479 (N_16479,N_16204,N_16048);
nor U16480 (N_16480,N_16182,N_16069);
or U16481 (N_16481,N_16161,N_16164);
and U16482 (N_16482,N_16036,N_16122);
nor U16483 (N_16483,N_16042,N_16019);
nor U16484 (N_16484,N_16136,N_16127);
or U16485 (N_16485,N_16135,N_16245);
nor U16486 (N_16486,N_16097,N_16024);
and U16487 (N_16487,N_16044,N_16025);
and U16488 (N_16488,N_16118,N_16060);
or U16489 (N_16489,N_16205,N_16161);
nand U16490 (N_16490,N_16231,N_16238);
and U16491 (N_16491,N_16181,N_16034);
nor U16492 (N_16492,N_16183,N_16094);
and U16493 (N_16493,N_16249,N_16185);
xor U16494 (N_16494,N_16125,N_16097);
nand U16495 (N_16495,N_16208,N_16134);
xor U16496 (N_16496,N_16101,N_16119);
xor U16497 (N_16497,N_16045,N_16006);
or U16498 (N_16498,N_16184,N_16056);
nor U16499 (N_16499,N_16099,N_16202);
or U16500 (N_16500,N_16441,N_16460);
xnor U16501 (N_16501,N_16341,N_16428);
nor U16502 (N_16502,N_16371,N_16389);
and U16503 (N_16503,N_16340,N_16259);
or U16504 (N_16504,N_16321,N_16402);
nor U16505 (N_16505,N_16462,N_16427);
nand U16506 (N_16506,N_16457,N_16374);
xnor U16507 (N_16507,N_16294,N_16337);
and U16508 (N_16508,N_16264,N_16476);
xor U16509 (N_16509,N_16478,N_16342);
nor U16510 (N_16510,N_16388,N_16253);
nor U16511 (N_16511,N_16417,N_16404);
nand U16512 (N_16512,N_16318,N_16414);
and U16513 (N_16513,N_16263,N_16411);
nand U16514 (N_16514,N_16379,N_16310);
xor U16515 (N_16515,N_16490,N_16426);
nor U16516 (N_16516,N_16488,N_16421);
and U16517 (N_16517,N_16416,N_16383);
xnor U16518 (N_16518,N_16333,N_16398);
and U16519 (N_16519,N_16312,N_16307);
or U16520 (N_16520,N_16257,N_16328);
nand U16521 (N_16521,N_16255,N_16293);
nor U16522 (N_16522,N_16471,N_16297);
and U16523 (N_16523,N_16407,N_16267);
and U16524 (N_16524,N_16309,N_16439);
nor U16525 (N_16525,N_16399,N_16452);
nand U16526 (N_16526,N_16258,N_16372);
xor U16527 (N_16527,N_16466,N_16287);
and U16528 (N_16528,N_16378,N_16285);
nand U16529 (N_16529,N_16306,N_16283);
xor U16530 (N_16530,N_16477,N_16420);
nand U16531 (N_16531,N_16376,N_16296);
and U16532 (N_16532,N_16268,N_16410);
nor U16533 (N_16533,N_16424,N_16369);
and U16534 (N_16534,N_16415,N_16348);
xnor U16535 (N_16535,N_16338,N_16298);
nand U16536 (N_16536,N_16300,N_16386);
xor U16537 (N_16537,N_16269,N_16373);
nor U16538 (N_16538,N_16412,N_16270);
xnor U16539 (N_16539,N_16302,N_16380);
and U16540 (N_16540,N_16438,N_16375);
xnor U16541 (N_16541,N_16409,N_16482);
nand U16542 (N_16542,N_16350,N_16450);
or U16543 (N_16543,N_16358,N_16262);
or U16544 (N_16544,N_16317,N_16431);
and U16545 (N_16545,N_16394,N_16304);
and U16546 (N_16546,N_16495,N_16481);
and U16547 (N_16547,N_16390,N_16385);
xnor U16548 (N_16548,N_16278,N_16282);
or U16549 (N_16549,N_16251,N_16393);
or U16550 (N_16550,N_16479,N_16382);
and U16551 (N_16551,N_16280,N_16423);
and U16552 (N_16552,N_16354,N_16408);
or U16553 (N_16553,N_16316,N_16273);
nand U16554 (N_16554,N_16433,N_16305);
or U16555 (N_16555,N_16472,N_16281);
and U16556 (N_16556,N_16397,N_16435);
xnor U16557 (N_16557,N_16492,N_16497);
nand U16558 (N_16558,N_16365,N_16325);
nor U16559 (N_16559,N_16455,N_16319);
and U16560 (N_16560,N_16436,N_16361);
nand U16561 (N_16561,N_16413,N_16367);
and U16562 (N_16562,N_16437,N_16467);
nand U16563 (N_16563,N_16326,N_16334);
xor U16564 (N_16564,N_16391,N_16336);
or U16565 (N_16565,N_16443,N_16403);
nand U16566 (N_16566,N_16475,N_16445);
nor U16567 (N_16567,N_16366,N_16483);
nor U16568 (N_16568,N_16276,N_16453);
and U16569 (N_16569,N_16355,N_16352);
and U16570 (N_16570,N_16335,N_16396);
nor U16571 (N_16571,N_16464,N_16480);
and U16572 (N_16572,N_16362,N_16486);
and U16573 (N_16573,N_16311,N_16401);
and U16574 (N_16574,N_16370,N_16346);
and U16575 (N_16575,N_16286,N_16384);
and U16576 (N_16576,N_16459,N_16498);
xnor U16577 (N_16577,N_16430,N_16252);
and U16578 (N_16578,N_16301,N_16451);
or U16579 (N_16579,N_16324,N_16491);
nand U16580 (N_16580,N_16327,N_16499);
xor U16581 (N_16581,N_16320,N_16465);
and U16582 (N_16582,N_16406,N_16496);
nor U16583 (N_16583,N_16377,N_16494);
and U16584 (N_16584,N_16425,N_16400);
or U16585 (N_16585,N_16351,N_16359);
or U16586 (N_16586,N_16434,N_16456);
and U16587 (N_16587,N_16313,N_16299);
or U16588 (N_16588,N_16418,N_16329);
or U16589 (N_16589,N_16363,N_16469);
nor U16590 (N_16590,N_16332,N_16353);
nor U16591 (N_16591,N_16303,N_16289);
xor U16592 (N_16592,N_16260,N_16470);
nand U16593 (N_16593,N_16315,N_16458);
nor U16594 (N_16594,N_16485,N_16291);
nand U16595 (N_16595,N_16256,N_16487);
nor U16596 (N_16596,N_16489,N_16274);
nand U16597 (N_16597,N_16473,N_16288);
nor U16598 (N_16598,N_16345,N_16349);
nand U16599 (N_16599,N_16429,N_16261);
xnor U16600 (N_16600,N_16339,N_16308);
and U16601 (N_16601,N_16265,N_16484);
nor U16602 (N_16602,N_16254,N_16347);
xnor U16603 (N_16603,N_16272,N_16284);
xnor U16604 (N_16604,N_16405,N_16446);
xnor U16605 (N_16605,N_16440,N_16279);
and U16606 (N_16606,N_16368,N_16295);
and U16607 (N_16607,N_16277,N_16442);
and U16608 (N_16608,N_16357,N_16419);
and U16609 (N_16609,N_16356,N_16292);
and U16610 (N_16610,N_16343,N_16422);
xnor U16611 (N_16611,N_16447,N_16449);
and U16612 (N_16612,N_16461,N_16364);
xnor U16613 (N_16613,N_16454,N_16271);
xnor U16614 (N_16614,N_16314,N_16474);
nor U16615 (N_16615,N_16387,N_16322);
or U16616 (N_16616,N_16448,N_16331);
and U16617 (N_16617,N_16275,N_16323);
nor U16618 (N_16618,N_16360,N_16330);
nor U16619 (N_16619,N_16344,N_16463);
xor U16620 (N_16620,N_16493,N_16266);
nand U16621 (N_16621,N_16432,N_16444);
xnor U16622 (N_16622,N_16290,N_16381);
nand U16623 (N_16623,N_16395,N_16468);
nand U16624 (N_16624,N_16392,N_16250);
or U16625 (N_16625,N_16485,N_16427);
nor U16626 (N_16626,N_16390,N_16297);
or U16627 (N_16627,N_16297,N_16307);
nand U16628 (N_16628,N_16488,N_16419);
or U16629 (N_16629,N_16409,N_16476);
or U16630 (N_16630,N_16328,N_16334);
and U16631 (N_16631,N_16253,N_16497);
and U16632 (N_16632,N_16369,N_16326);
and U16633 (N_16633,N_16254,N_16332);
and U16634 (N_16634,N_16355,N_16291);
or U16635 (N_16635,N_16254,N_16410);
nand U16636 (N_16636,N_16498,N_16382);
and U16637 (N_16637,N_16365,N_16302);
xnor U16638 (N_16638,N_16269,N_16285);
nand U16639 (N_16639,N_16269,N_16315);
or U16640 (N_16640,N_16470,N_16255);
nor U16641 (N_16641,N_16477,N_16318);
nor U16642 (N_16642,N_16467,N_16363);
or U16643 (N_16643,N_16273,N_16360);
or U16644 (N_16644,N_16337,N_16290);
and U16645 (N_16645,N_16451,N_16485);
nor U16646 (N_16646,N_16338,N_16416);
and U16647 (N_16647,N_16340,N_16452);
nand U16648 (N_16648,N_16276,N_16422);
nor U16649 (N_16649,N_16272,N_16345);
xnor U16650 (N_16650,N_16325,N_16274);
and U16651 (N_16651,N_16266,N_16322);
xnor U16652 (N_16652,N_16269,N_16415);
nor U16653 (N_16653,N_16440,N_16432);
xnor U16654 (N_16654,N_16287,N_16336);
and U16655 (N_16655,N_16380,N_16372);
or U16656 (N_16656,N_16275,N_16356);
xnor U16657 (N_16657,N_16448,N_16461);
nor U16658 (N_16658,N_16254,N_16330);
or U16659 (N_16659,N_16422,N_16287);
nor U16660 (N_16660,N_16262,N_16311);
nand U16661 (N_16661,N_16461,N_16483);
nand U16662 (N_16662,N_16270,N_16427);
and U16663 (N_16663,N_16336,N_16467);
nand U16664 (N_16664,N_16432,N_16471);
and U16665 (N_16665,N_16270,N_16350);
nor U16666 (N_16666,N_16488,N_16352);
or U16667 (N_16667,N_16482,N_16481);
and U16668 (N_16668,N_16347,N_16278);
and U16669 (N_16669,N_16308,N_16291);
or U16670 (N_16670,N_16410,N_16424);
nor U16671 (N_16671,N_16462,N_16278);
nand U16672 (N_16672,N_16357,N_16284);
nand U16673 (N_16673,N_16415,N_16391);
or U16674 (N_16674,N_16390,N_16469);
and U16675 (N_16675,N_16322,N_16482);
or U16676 (N_16676,N_16364,N_16422);
and U16677 (N_16677,N_16284,N_16441);
xor U16678 (N_16678,N_16264,N_16345);
or U16679 (N_16679,N_16266,N_16499);
nand U16680 (N_16680,N_16319,N_16348);
nor U16681 (N_16681,N_16416,N_16299);
xor U16682 (N_16682,N_16387,N_16338);
nand U16683 (N_16683,N_16398,N_16395);
nand U16684 (N_16684,N_16367,N_16330);
xor U16685 (N_16685,N_16274,N_16433);
and U16686 (N_16686,N_16435,N_16373);
nand U16687 (N_16687,N_16374,N_16293);
or U16688 (N_16688,N_16293,N_16291);
nand U16689 (N_16689,N_16464,N_16403);
nand U16690 (N_16690,N_16364,N_16272);
nand U16691 (N_16691,N_16270,N_16353);
and U16692 (N_16692,N_16293,N_16295);
or U16693 (N_16693,N_16276,N_16346);
nand U16694 (N_16694,N_16417,N_16302);
nand U16695 (N_16695,N_16363,N_16452);
and U16696 (N_16696,N_16390,N_16352);
nand U16697 (N_16697,N_16394,N_16467);
nor U16698 (N_16698,N_16471,N_16475);
nor U16699 (N_16699,N_16368,N_16454);
or U16700 (N_16700,N_16353,N_16421);
and U16701 (N_16701,N_16430,N_16327);
and U16702 (N_16702,N_16368,N_16290);
nand U16703 (N_16703,N_16336,N_16395);
nand U16704 (N_16704,N_16430,N_16478);
and U16705 (N_16705,N_16409,N_16410);
and U16706 (N_16706,N_16398,N_16337);
and U16707 (N_16707,N_16378,N_16310);
nand U16708 (N_16708,N_16457,N_16257);
or U16709 (N_16709,N_16311,N_16484);
xnor U16710 (N_16710,N_16414,N_16465);
nor U16711 (N_16711,N_16372,N_16412);
or U16712 (N_16712,N_16268,N_16359);
xnor U16713 (N_16713,N_16250,N_16337);
xnor U16714 (N_16714,N_16329,N_16331);
nand U16715 (N_16715,N_16285,N_16442);
and U16716 (N_16716,N_16253,N_16333);
nor U16717 (N_16717,N_16376,N_16385);
xnor U16718 (N_16718,N_16438,N_16367);
nand U16719 (N_16719,N_16318,N_16267);
or U16720 (N_16720,N_16360,N_16359);
nor U16721 (N_16721,N_16379,N_16449);
and U16722 (N_16722,N_16457,N_16357);
nand U16723 (N_16723,N_16326,N_16405);
and U16724 (N_16724,N_16344,N_16389);
xor U16725 (N_16725,N_16472,N_16397);
or U16726 (N_16726,N_16482,N_16484);
and U16727 (N_16727,N_16276,N_16477);
and U16728 (N_16728,N_16368,N_16273);
xnor U16729 (N_16729,N_16452,N_16334);
or U16730 (N_16730,N_16260,N_16497);
and U16731 (N_16731,N_16392,N_16281);
nor U16732 (N_16732,N_16451,N_16359);
and U16733 (N_16733,N_16318,N_16394);
nor U16734 (N_16734,N_16456,N_16291);
or U16735 (N_16735,N_16389,N_16478);
xor U16736 (N_16736,N_16380,N_16288);
and U16737 (N_16737,N_16400,N_16402);
and U16738 (N_16738,N_16458,N_16454);
xnor U16739 (N_16739,N_16444,N_16462);
and U16740 (N_16740,N_16368,N_16282);
and U16741 (N_16741,N_16453,N_16469);
nand U16742 (N_16742,N_16380,N_16357);
xor U16743 (N_16743,N_16476,N_16482);
or U16744 (N_16744,N_16320,N_16255);
xnor U16745 (N_16745,N_16489,N_16329);
nand U16746 (N_16746,N_16320,N_16254);
or U16747 (N_16747,N_16476,N_16425);
nand U16748 (N_16748,N_16490,N_16286);
and U16749 (N_16749,N_16355,N_16379);
nand U16750 (N_16750,N_16662,N_16658);
nor U16751 (N_16751,N_16522,N_16721);
xor U16752 (N_16752,N_16666,N_16697);
and U16753 (N_16753,N_16618,N_16733);
and U16754 (N_16754,N_16531,N_16535);
xnor U16755 (N_16755,N_16626,N_16639);
nor U16756 (N_16756,N_16627,N_16582);
nor U16757 (N_16757,N_16716,N_16726);
xor U16758 (N_16758,N_16576,N_16525);
or U16759 (N_16759,N_16654,N_16581);
or U16760 (N_16760,N_16507,N_16688);
and U16761 (N_16761,N_16536,N_16604);
nand U16762 (N_16762,N_16743,N_16622);
or U16763 (N_16763,N_16571,N_16564);
or U16764 (N_16764,N_16676,N_16583);
xor U16765 (N_16765,N_16601,N_16606);
and U16766 (N_16766,N_16738,N_16749);
nor U16767 (N_16767,N_16737,N_16506);
and U16768 (N_16768,N_16603,N_16530);
and U16769 (N_16769,N_16691,N_16669);
nand U16770 (N_16770,N_16569,N_16673);
nand U16771 (N_16771,N_16647,N_16500);
or U16772 (N_16772,N_16698,N_16596);
and U16773 (N_16773,N_16515,N_16709);
nor U16774 (N_16774,N_16529,N_16703);
and U16775 (N_16775,N_16527,N_16693);
nand U16776 (N_16776,N_16549,N_16600);
or U16777 (N_16777,N_16517,N_16731);
or U16778 (N_16778,N_16577,N_16505);
xnor U16779 (N_16779,N_16521,N_16718);
xor U16780 (N_16780,N_16740,N_16663);
nor U16781 (N_16781,N_16635,N_16748);
nor U16782 (N_16782,N_16539,N_16623);
and U16783 (N_16783,N_16540,N_16580);
and U16784 (N_16784,N_16545,N_16561);
nor U16785 (N_16785,N_16547,N_16584);
nor U16786 (N_16786,N_16645,N_16516);
or U16787 (N_16787,N_16544,N_16675);
nor U16788 (N_16788,N_16509,N_16724);
nor U16789 (N_16789,N_16620,N_16548);
nand U16790 (N_16790,N_16586,N_16652);
nor U16791 (N_16791,N_16538,N_16742);
and U16792 (N_16792,N_16661,N_16612);
xor U16793 (N_16793,N_16690,N_16682);
xnor U16794 (N_16794,N_16741,N_16653);
nor U16795 (N_16795,N_16725,N_16573);
or U16796 (N_16796,N_16602,N_16723);
nor U16797 (N_16797,N_16649,N_16686);
and U16798 (N_16798,N_16514,N_16651);
nor U16799 (N_16799,N_16713,N_16615);
nor U16800 (N_16800,N_16665,N_16629);
and U16801 (N_16801,N_16502,N_16542);
and U16802 (N_16802,N_16519,N_16613);
and U16803 (N_16803,N_16533,N_16575);
xor U16804 (N_16804,N_16554,N_16659);
nand U16805 (N_16805,N_16719,N_16558);
nand U16806 (N_16806,N_16624,N_16736);
nand U16807 (N_16807,N_16727,N_16672);
and U16808 (N_16808,N_16707,N_16714);
nand U16809 (N_16809,N_16543,N_16734);
nand U16810 (N_16810,N_16578,N_16617);
nand U16811 (N_16811,N_16699,N_16568);
or U16812 (N_16812,N_16504,N_16608);
and U16813 (N_16813,N_16598,N_16656);
or U16814 (N_16814,N_16503,N_16550);
xor U16815 (N_16815,N_16594,N_16557);
and U16816 (N_16816,N_16694,N_16735);
xnor U16817 (N_16817,N_16619,N_16621);
and U16818 (N_16818,N_16706,N_16609);
nand U16819 (N_16819,N_16689,N_16563);
xnor U16820 (N_16820,N_16587,N_16732);
nand U16821 (N_16821,N_16674,N_16566);
or U16822 (N_16822,N_16556,N_16715);
nor U16823 (N_16823,N_16570,N_16729);
nor U16824 (N_16824,N_16643,N_16705);
nor U16825 (N_16825,N_16560,N_16501);
nand U16826 (N_16826,N_16526,N_16524);
or U16827 (N_16827,N_16546,N_16746);
nand U16828 (N_16828,N_16523,N_16593);
xor U16829 (N_16829,N_16508,N_16589);
nand U16830 (N_16830,N_16616,N_16660);
xnor U16831 (N_16831,N_16520,N_16551);
nand U16832 (N_16832,N_16534,N_16687);
nand U16833 (N_16833,N_16711,N_16671);
nor U16834 (N_16834,N_16552,N_16646);
xor U16835 (N_16835,N_16704,N_16605);
nand U16836 (N_16836,N_16744,N_16510);
nor U16837 (N_16837,N_16712,N_16730);
xnor U16838 (N_16838,N_16597,N_16630);
and U16839 (N_16839,N_16684,N_16528);
or U16840 (N_16840,N_16681,N_16678);
or U16841 (N_16841,N_16553,N_16632);
or U16842 (N_16842,N_16592,N_16512);
nand U16843 (N_16843,N_16679,N_16591);
and U16844 (N_16844,N_16631,N_16588);
and U16845 (N_16845,N_16638,N_16722);
nor U16846 (N_16846,N_16511,N_16633);
or U16847 (N_16847,N_16642,N_16701);
nor U16848 (N_16848,N_16650,N_16692);
nand U16849 (N_16849,N_16648,N_16565);
xor U16850 (N_16850,N_16667,N_16668);
xnor U16851 (N_16851,N_16541,N_16590);
and U16852 (N_16852,N_16717,N_16610);
and U16853 (N_16853,N_16657,N_16685);
nand U16854 (N_16854,N_16641,N_16555);
and U16855 (N_16855,N_16567,N_16728);
or U16856 (N_16856,N_16572,N_16655);
nand U16857 (N_16857,N_16747,N_16513);
nand U16858 (N_16858,N_16628,N_16574);
or U16859 (N_16859,N_16696,N_16710);
nand U16860 (N_16860,N_16702,N_16677);
xor U16861 (N_16861,N_16670,N_16695);
and U16862 (N_16862,N_16700,N_16637);
or U16863 (N_16863,N_16636,N_16537);
nor U16864 (N_16864,N_16683,N_16634);
xnor U16865 (N_16865,N_16518,N_16599);
nor U16866 (N_16866,N_16680,N_16708);
xnor U16867 (N_16867,N_16611,N_16532);
xnor U16868 (N_16868,N_16579,N_16625);
and U16869 (N_16869,N_16644,N_16664);
xor U16870 (N_16870,N_16720,N_16585);
xnor U16871 (N_16871,N_16559,N_16745);
nand U16872 (N_16872,N_16739,N_16640);
nor U16873 (N_16873,N_16614,N_16607);
nand U16874 (N_16874,N_16595,N_16562);
nor U16875 (N_16875,N_16593,N_16742);
nor U16876 (N_16876,N_16668,N_16511);
nand U16877 (N_16877,N_16657,N_16591);
nor U16878 (N_16878,N_16689,N_16693);
xnor U16879 (N_16879,N_16597,N_16523);
nand U16880 (N_16880,N_16502,N_16656);
and U16881 (N_16881,N_16692,N_16505);
xnor U16882 (N_16882,N_16708,N_16696);
nand U16883 (N_16883,N_16519,N_16624);
or U16884 (N_16884,N_16734,N_16516);
or U16885 (N_16885,N_16594,N_16644);
xor U16886 (N_16886,N_16648,N_16513);
nand U16887 (N_16887,N_16615,N_16660);
nand U16888 (N_16888,N_16550,N_16743);
nand U16889 (N_16889,N_16711,N_16714);
nand U16890 (N_16890,N_16725,N_16553);
nand U16891 (N_16891,N_16527,N_16584);
xor U16892 (N_16892,N_16736,N_16653);
or U16893 (N_16893,N_16645,N_16603);
and U16894 (N_16894,N_16548,N_16516);
nor U16895 (N_16895,N_16744,N_16656);
nor U16896 (N_16896,N_16638,N_16699);
and U16897 (N_16897,N_16511,N_16541);
xnor U16898 (N_16898,N_16573,N_16662);
xnor U16899 (N_16899,N_16575,N_16673);
or U16900 (N_16900,N_16507,N_16726);
and U16901 (N_16901,N_16597,N_16547);
nand U16902 (N_16902,N_16727,N_16557);
nor U16903 (N_16903,N_16681,N_16559);
or U16904 (N_16904,N_16557,N_16596);
nor U16905 (N_16905,N_16563,N_16627);
xnor U16906 (N_16906,N_16629,N_16641);
or U16907 (N_16907,N_16539,N_16556);
nor U16908 (N_16908,N_16732,N_16502);
or U16909 (N_16909,N_16739,N_16567);
nand U16910 (N_16910,N_16611,N_16530);
nor U16911 (N_16911,N_16504,N_16650);
nand U16912 (N_16912,N_16650,N_16631);
nor U16913 (N_16913,N_16673,N_16538);
nor U16914 (N_16914,N_16748,N_16555);
nand U16915 (N_16915,N_16669,N_16582);
or U16916 (N_16916,N_16585,N_16711);
xor U16917 (N_16917,N_16513,N_16525);
nand U16918 (N_16918,N_16552,N_16514);
nor U16919 (N_16919,N_16524,N_16535);
or U16920 (N_16920,N_16507,N_16675);
or U16921 (N_16921,N_16555,N_16679);
nand U16922 (N_16922,N_16704,N_16510);
nand U16923 (N_16923,N_16541,N_16695);
and U16924 (N_16924,N_16548,N_16744);
and U16925 (N_16925,N_16648,N_16518);
or U16926 (N_16926,N_16545,N_16696);
nand U16927 (N_16927,N_16640,N_16655);
nand U16928 (N_16928,N_16724,N_16594);
nor U16929 (N_16929,N_16574,N_16718);
and U16930 (N_16930,N_16688,N_16533);
xnor U16931 (N_16931,N_16546,N_16587);
xnor U16932 (N_16932,N_16715,N_16546);
or U16933 (N_16933,N_16580,N_16585);
or U16934 (N_16934,N_16692,N_16604);
xnor U16935 (N_16935,N_16746,N_16656);
nor U16936 (N_16936,N_16630,N_16702);
or U16937 (N_16937,N_16576,N_16580);
nand U16938 (N_16938,N_16611,N_16679);
nor U16939 (N_16939,N_16563,N_16739);
and U16940 (N_16940,N_16639,N_16586);
and U16941 (N_16941,N_16670,N_16693);
or U16942 (N_16942,N_16670,N_16525);
and U16943 (N_16943,N_16650,N_16663);
nand U16944 (N_16944,N_16632,N_16611);
nand U16945 (N_16945,N_16708,N_16623);
nor U16946 (N_16946,N_16531,N_16697);
or U16947 (N_16947,N_16642,N_16722);
and U16948 (N_16948,N_16601,N_16747);
nor U16949 (N_16949,N_16616,N_16566);
xnor U16950 (N_16950,N_16703,N_16626);
or U16951 (N_16951,N_16503,N_16525);
nor U16952 (N_16952,N_16656,N_16626);
xor U16953 (N_16953,N_16653,N_16592);
or U16954 (N_16954,N_16630,N_16583);
or U16955 (N_16955,N_16534,N_16575);
nand U16956 (N_16956,N_16614,N_16731);
xnor U16957 (N_16957,N_16698,N_16524);
nor U16958 (N_16958,N_16707,N_16551);
nand U16959 (N_16959,N_16635,N_16529);
nor U16960 (N_16960,N_16500,N_16746);
nand U16961 (N_16961,N_16655,N_16624);
or U16962 (N_16962,N_16666,N_16578);
or U16963 (N_16963,N_16558,N_16593);
or U16964 (N_16964,N_16505,N_16528);
or U16965 (N_16965,N_16562,N_16565);
or U16966 (N_16966,N_16734,N_16534);
or U16967 (N_16967,N_16513,N_16588);
nor U16968 (N_16968,N_16585,N_16698);
or U16969 (N_16969,N_16564,N_16521);
nor U16970 (N_16970,N_16546,N_16513);
xor U16971 (N_16971,N_16679,N_16525);
nor U16972 (N_16972,N_16728,N_16681);
nand U16973 (N_16973,N_16700,N_16670);
xor U16974 (N_16974,N_16517,N_16748);
or U16975 (N_16975,N_16506,N_16607);
and U16976 (N_16976,N_16694,N_16704);
and U16977 (N_16977,N_16560,N_16712);
xnor U16978 (N_16978,N_16537,N_16617);
nand U16979 (N_16979,N_16737,N_16664);
and U16980 (N_16980,N_16631,N_16617);
and U16981 (N_16981,N_16609,N_16616);
xnor U16982 (N_16982,N_16506,N_16719);
nand U16983 (N_16983,N_16732,N_16683);
xor U16984 (N_16984,N_16561,N_16664);
and U16985 (N_16985,N_16737,N_16690);
and U16986 (N_16986,N_16703,N_16620);
or U16987 (N_16987,N_16571,N_16511);
or U16988 (N_16988,N_16676,N_16715);
nand U16989 (N_16989,N_16598,N_16621);
nor U16990 (N_16990,N_16580,N_16608);
and U16991 (N_16991,N_16531,N_16686);
and U16992 (N_16992,N_16748,N_16525);
or U16993 (N_16993,N_16543,N_16649);
nor U16994 (N_16994,N_16739,N_16630);
or U16995 (N_16995,N_16511,N_16561);
and U16996 (N_16996,N_16620,N_16736);
xnor U16997 (N_16997,N_16644,N_16646);
xnor U16998 (N_16998,N_16685,N_16729);
xnor U16999 (N_16999,N_16643,N_16629);
nand U17000 (N_17000,N_16991,N_16992);
nand U17001 (N_17001,N_16855,N_16989);
nor U17002 (N_17002,N_16924,N_16854);
or U17003 (N_17003,N_16884,N_16877);
and U17004 (N_17004,N_16885,N_16865);
nor U17005 (N_17005,N_16775,N_16914);
or U17006 (N_17006,N_16882,N_16873);
xnor U17007 (N_17007,N_16892,N_16838);
xnor U17008 (N_17008,N_16891,N_16994);
nand U17009 (N_17009,N_16782,N_16887);
or U17010 (N_17010,N_16979,N_16922);
nor U17011 (N_17011,N_16793,N_16988);
nor U17012 (N_17012,N_16751,N_16795);
or U17013 (N_17013,N_16761,N_16964);
xor U17014 (N_17014,N_16801,N_16978);
or U17015 (N_17015,N_16764,N_16916);
xor U17016 (N_17016,N_16990,N_16813);
or U17017 (N_17017,N_16796,N_16966);
or U17018 (N_17018,N_16819,N_16844);
or U17019 (N_17019,N_16980,N_16934);
nor U17020 (N_17020,N_16859,N_16953);
nor U17021 (N_17021,N_16845,N_16785);
and U17022 (N_17022,N_16802,N_16757);
and U17023 (N_17023,N_16883,N_16961);
or U17024 (N_17024,N_16791,N_16901);
nor U17025 (N_17025,N_16833,N_16843);
xor U17026 (N_17026,N_16940,N_16875);
and U17027 (N_17027,N_16888,N_16907);
or U17028 (N_17028,N_16759,N_16899);
nand U17029 (N_17029,N_16913,N_16918);
and U17030 (N_17030,N_16783,N_16823);
xor U17031 (N_17031,N_16937,N_16968);
nor U17032 (N_17032,N_16935,N_16822);
xnor U17033 (N_17033,N_16930,N_16815);
nor U17034 (N_17034,N_16837,N_16977);
xnor U17035 (N_17035,N_16772,N_16849);
nand U17036 (N_17036,N_16932,N_16797);
and U17037 (N_17037,N_16763,N_16829);
nor U17038 (N_17038,N_16834,N_16963);
or U17039 (N_17039,N_16766,N_16920);
nand U17040 (N_17040,N_16773,N_16794);
or U17041 (N_17041,N_16906,N_16821);
xor U17042 (N_17042,N_16771,N_16840);
nor U17043 (N_17043,N_16809,N_16879);
nand U17044 (N_17044,N_16959,N_16832);
nor U17045 (N_17045,N_16758,N_16826);
xor U17046 (N_17046,N_16956,N_16902);
nand U17047 (N_17047,N_16944,N_16921);
nand U17048 (N_17048,N_16862,N_16933);
nor U17049 (N_17049,N_16972,N_16811);
nor U17050 (N_17050,N_16805,N_16919);
xnor U17051 (N_17051,N_16965,N_16752);
nor U17052 (N_17052,N_16903,N_16756);
and U17053 (N_17053,N_16828,N_16860);
and U17054 (N_17054,N_16905,N_16942);
nand U17055 (N_17055,N_16886,N_16911);
xor U17056 (N_17056,N_16957,N_16871);
or U17057 (N_17057,N_16850,N_16841);
or U17058 (N_17058,N_16970,N_16869);
nand U17059 (N_17059,N_16820,N_16835);
xor U17060 (N_17060,N_16998,N_16857);
or U17061 (N_17061,N_16825,N_16951);
or U17062 (N_17062,N_16769,N_16755);
and U17063 (N_17063,N_16868,N_16867);
nor U17064 (N_17064,N_16852,N_16804);
and U17065 (N_17065,N_16952,N_16962);
nand U17066 (N_17066,N_16798,N_16760);
and U17067 (N_17067,N_16807,N_16851);
nand U17068 (N_17068,N_16974,N_16925);
nand U17069 (N_17069,N_16982,N_16910);
and U17070 (N_17070,N_16799,N_16864);
xnor U17071 (N_17071,N_16770,N_16839);
nand U17072 (N_17072,N_16790,N_16872);
or U17073 (N_17073,N_16858,N_16950);
and U17074 (N_17074,N_16817,N_16784);
and U17075 (N_17075,N_16881,N_16776);
nor U17076 (N_17076,N_16993,N_16768);
nor U17077 (N_17077,N_16848,N_16904);
or U17078 (N_17078,N_16927,N_16917);
xor U17079 (N_17079,N_16774,N_16975);
xnor U17080 (N_17080,N_16971,N_16827);
or U17081 (N_17081,N_16831,N_16787);
or U17082 (N_17082,N_16778,N_16870);
nor U17083 (N_17083,N_16847,N_16792);
xnor U17084 (N_17084,N_16846,N_16810);
or U17085 (N_17085,N_16987,N_16830);
nor U17086 (N_17086,N_16836,N_16929);
nand U17087 (N_17087,N_16945,N_16954);
or U17088 (N_17088,N_16861,N_16786);
xnor U17089 (N_17089,N_16880,N_16876);
or U17090 (N_17090,N_16788,N_16936);
nand U17091 (N_17091,N_16941,N_16908);
nand U17092 (N_17092,N_16949,N_16824);
and U17093 (N_17093,N_16863,N_16983);
xor U17094 (N_17094,N_16814,N_16750);
and U17095 (N_17095,N_16931,N_16874);
xor U17096 (N_17096,N_16789,N_16897);
nor U17097 (N_17097,N_16909,N_16939);
nor U17098 (N_17098,N_16866,N_16753);
or U17099 (N_17099,N_16985,N_16893);
nand U17100 (N_17100,N_16878,N_16856);
nand U17101 (N_17101,N_16960,N_16955);
nand U17102 (N_17102,N_16762,N_16812);
and U17103 (N_17103,N_16754,N_16842);
nand U17104 (N_17104,N_16943,N_16894);
and U17105 (N_17105,N_16896,N_16926);
nor U17106 (N_17106,N_16976,N_16803);
and U17107 (N_17107,N_16946,N_16947);
nor U17108 (N_17108,N_16958,N_16765);
nand U17109 (N_17109,N_16973,N_16915);
nand U17110 (N_17110,N_16808,N_16767);
xnor U17111 (N_17111,N_16800,N_16999);
nor U17112 (N_17112,N_16816,N_16969);
nand U17113 (N_17113,N_16984,N_16806);
nand U17114 (N_17114,N_16781,N_16780);
xnor U17115 (N_17115,N_16938,N_16997);
xnor U17116 (N_17116,N_16853,N_16996);
and U17117 (N_17117,N_16928,N_16948);
nor U17118 (N_17118,N_16889,N_16779);
and U17119 (N_17119,N_16900,N_16912);
nand U17120 (N_17120,N_16967,N_16986);
xor U17121 (N_17121,N_16890,N_16923);
nand U17122 (N_17122,N_16777,N_16818);
nor U17123 (N_17123,N_16898,N_16895);
xor U17124 (N_17124,N_16995,N_16981);
nand U17125 (N_17125,N_16910,N_16816);
nand U17126 (N_17126,N_16809,N_16805);
xnor U17127 (N_17127,N_16952,N_16959);
and U17128 (N_17128,N_16834,N_16785);
nand U17129 (N_17129,N_16810,N_16911);
nor U17130 (N_17130,N_16809,N_16812);
xor U17131 (N_17131,N_16923,N_16949);
and U17132 (N_17132,N_16864,N_16772);
nor U17133 (N_17133,N_16750,N_16861);
or U17134 (N_17134,N_16928,N_16767);
nand U17135 (N_17135,N_16769,N_16966);
nand U17136 (N_17136,N_16934,N_16846);
nand U17137 (N_17137,N_16981,N_16810);
or U17138 (N_17138,N_16929,N_16915);
nor U17139 (N_17139,N_16766,N_16979);
nor U17140 (N_17140,N_16878,N_16922);
nor U17141 (N_17141,N_16852,N_16885);
or U17142 (N_17142,N_16783,N_16778);
and U17143 (N_17143,N_16761,N_16911);
and U17144 (N_17144,N_16850,N_16967);
and U17145 (N_17145,N_16886,N_16974);
or U17146 (N_17146,N_16911,N_16937);
xnor U17147 (N_17147,N_16836,N_16789);
and U17148 (N_17148,N_16829,N_16793);
xnor U17149 (N_17149,N_16901,N_16814);
or U17150 (N_17150,N_16924,N_16900);
nand U17151 (N_17151,N_16968,N_16766);
xor U17152 (N_17152,N_16913,N_16962);
or U17153 (N_17153,N_16957,N_16873);
nand U17154 (N_17154,N_16766,N_16997);
and U17155 (N_17155,N_16817,N_16819);
nand U17156 (N_17156,N_16769,N_16921);
nand U17157 (N_17157,N_16835,N_16887);
nor U17158 (N_17158,N_16877,N_16975);
or U17159 (N_17159,N_16828,N_16856);
nand U17160 (N_17160,N_16789,N_16902);
xor U17161 (N_17161,N_16951,N_16963);
nor U17162 (N_17162,N_16961,N_16828);
nand U17163 (N_17163,N_16924,N_16757);
or U17164 (N_17164,N_16887,N_16839);
xor U17165 (N_17165,N_16796,N_16781);
or U17166 (N_17166,N_16970,N_16973);
nand U17167 (N_17167,N_16977,N_16906);
or U17168 (N_17168,N_16958,N_16978);
xnor U17169 (N_17169,N_16979,N_16812);
nor U17170 (N_17170,N_16786,N_16770);
nor U17171 (N_17171,N_16856,N_16976);
nand U17172 (N_17172,N_16848,N_16797);
nand U17173 (N_17173,N_16902,N_16986);
xor U17174 (N_17174,N_16901,N_16876);
nand U17175 (N_17175,N_16929,N_16850);
nand U17176 (N_17176,N_16943,N_16806);
nor U17177 (N_17177,N_16870,N_16836);
nor U17178 (N_17178,N_16975,N_16907);
xor U17179 (N_17179,N_16839,N_16960);
nand U17180 (N_17180,N_16978,N_16953);
and U17181 (N_17181,N_16919,N_16908);
xnor U17182 (N_17182,N_16971,N_16829);
nor U17183 (N_17183,N_16973,N_16917);
and U17184 (N_17184,N_16832,N_16780);
nor U17185 (N_17185,N_16859,N_16757);
nand U17186 (N_17186,N_16858,N_16898);
nor U17187 (N_17187,N_16909,N_16921);
nand U17188 (N_17188,N_16868,N_16772);
or U17189 (N_17189,N_16908,N_16786);
nand U17190 (N_17190,N_16848,N_16954);
nand U17191 (N_17191,N_16875,N_16895);
xnor U17192 (N_17192,N_16982,N_16859);
and U17193 (N_17193,N_16828,N_16776);
or U17194 (N_17194,N_16854,N_16792);
nor U17195 (N_17195,N_16851,N_16872);
nor U17196 (N_17196,N_16955,N_16825);
xnor U17197 (N_17197,N_16763,N_16945);
and U17198 (N_17198,N_16756,N_16799);
or U17199 (N_17199,N_16754,N_16990);
nor U17200 (N_17200,N_16917,N_16987);
nor U17201 (N_17201,N_16895,N_16764);
or U17202 (N_17202,N_16907,N_16901);
nor U17203 (N_17203,N_16819,N_16815);
and U17204 (N_17204,N_16790,N_16995);
and U17205 (N_17205,N_16785,N_16861);
nand U17206 (N_17206,N_16773,N_16767);
xnor U17207 (N_17207,N_16842,N_16983);
nand U17208 (N_17208,N_16908,N_16805);
nor U17209 (N_17209,N_16817,N_16884);
nand U17210 (N_17210,N_16853,N_16902);
xor U17211 (N_17211,N_16975,N_16894);
nor U17212 (N_17212,N_16922,N_16754);
xnor U17213 (N_17213,N_16759,N_16978);
nand U17214 (N_17214,N_16955,N_16939);
nor U17215 (N_17215,N_16855,N_16751);
nor U17216 (N_17216,N_16848,N_16981);
or U17217 (N_17217,N_16802,N_16837);
or U17218 (N_17218,N_16839,N_16838);
nor U17219 (N_17219,N_16914,N_16847);
nand U17220 (N_17220,N_16754,N_16967);
and U17221 (N_17221,N_16767,N_16869);
and U17222 (N_17222,N_16778,N_16943);
and U17223 (N_17223,N_16853,N_16931);
xnor U17224 (N_17224,N_16750,N_16818);
or U17225 (N_17225,N_16764,N_16800);
nor U17226 (N_17226,N_16878,N_16979);
nand U17227 (N_17227,N_16973,N_16909);
nor U17228 (N_17228,N_16954,N_16760);
and U17229 (N_17229,N_16764,N_16864);
xnor U17230 (N_17230,N_16826,N_16760);
and U17231 (N_17231,N_16933,N_16942);
nand U17232 (N_17232,N_16781,N_16930);
and U17233 (N_17233,N_16820,N_16919);
and U17234 (N_17234,N_16771,N_16797);
and U17235 (N_17235,N_16845,N_16843);
nor U17236 (N_17236,N_16958,N_16955);
nand U17237 (N_17237,N_16910,N_16824);
and U17238 (N_17238,N_16875,N_16943);
nor U17239 (N_17239,N_16859,N_16758);
nor U17240 (N_17240,N_16787,N_16845);
or U17241 (N_17241,N_16988,N_16966);
xnor U17242 (N_17242,N_16852,N_16884);
nor U17243 (N_17243,N_16926,N_16935);
xnor U17244 (N_17244,N_16996,N_16948);
xor U17245 (N_17245,N_16911,N_16965);
nor U17246 (N_17246,N_16825,N_16756);
and U17247 (N_17247,N_16901,N_16952);
and U17248 (N_17248,N_16873,N_16859);
nor U17249 (N_17249,N_16916,N_16896);
and U17250 (N_17250,N_17022,N_17210);
or U17251 (N_17251,N_17014,N_17104);
nor U17252 (N_17252,N_17085,N_17156);
xor U17253 (N_17253,N_17109,N_17000);
nor U17254 (N_17254,N_17007,N_17149);
nand U17255 (N_17255,N_17028,N_17064);
and U17256 (N_17256,N_17213,N_17114);
nand U17257 (N_17257,N_17170,N_17133);
and U17258 (N_17258,N_17055,N_17226);
xnor U17259 (N_17259,N_17079,N_17101);
nor U17260 (N_17260,N_17186,N_17177);
and U17261 (N_17261,N_17225,N_17152);
nand U17262 (N_17262,N_17023,N_17172);
and U17263 (N_17263,N_17042,N_17142);
nor U17264 (N_17264,N_17088,N_17120);
nor U17265 (N_17265,N_17159,N_17129);
nor U17266 (N_17266,N_17036,N_17082);
nand U17267 (N_17267,N_17232,N_17209);
nor U17268 (N_17268,N_17113,N_17005);
nand U17269 (N_17269,N_17092,N_17026);
nand U17270 (N_17270,N_17160,N_17017);
nand U17271 (N_17271,N_17110,N_17157);
nand U17272 (N_17272,N_17094,N_17090);
xor U17273 (N_17273,N_17001,N_17033);
or U17274 (N_17274,N_17009,N_17121);
nand U17275 (N_17275,N_17103,N_17089);
and U17276 (N_17276,N_17173,N_17068);
nor U17277 (N_17277,N_17027,N_17218);
xor U17278 (N_17278,N_17185,N_17011);
or U17279 (N_17279,N_17201,N_17025);
nand U17280 (N_17280,N_17097,N_17031);
xnor U17281 (N_17281,N_17056,N_17204);
nand U17282 (N_17282,N_17207,N_17229);
nor U17283 (N_17283,N_17248,N_17205);
and U17284 (N_17284,N_17029,N_17118);
xnor U17285 (N_17285,N_17153,N_17061);
or U17286 (N_17286,N_17182,N_17168);
and U17287 (N_17287,N_17234,N_17143);
nor U17288 (N_17288,N_17141,N_17069);
xor U17289 (N_17289,N_17112,N_17034);
or U17290 (N_17290,N_17239,N_17048);
or U17291 (N_17291,N_17083,N_17193);
xnor U17292 (N_17292,N_17087,N_17190);
nor U17293 (N_17293,N_17035,N_17191);
nor U17294 (N_17294,N_17108,N_17115);
or U17295 (N_17295,N_17222,N_17006);
or U17296 (N_17296,N_17155,N_17164);
xnor U17297 (N_17297,N_17166,N_17214);
or U17298 (N_17298,N_17139,N_17242);
or U17299 (N_17299,N_17039,N_17163);
or U17300 (N_17300,N_17077,N_17111);
nor U17301 (N_17301,N_17008,N_17013);
nor U17302 (N_17302,N_17203,N_17236);
and U17303 (N_17303,N_17073,N_17070);
and U17304 (N_17304,N_17054,N_17223);
or U17305 (N_17305,N_17158,N_17187);
nor U17306 (N_17306,N_17053,N_17198);
nand U17307 (N_17307,N_17049,N_17220);
and U17308 (N_17308,N_17067,N_17117);
nor U17309 (N_17309,N_17241,N_17043);
and U17310 (N_17310,N_17125,N_17199);
nor U17311 (N_17311,N_17084,N_17154);
xnor U17312 (N_17312,N_17127,N_17058);
and U17313 (N_17313,N_17194,N_17136);
and U17314 (N_17314,N_17140,N_17135);
nand U17315 (N_17315,N_17217,N_17010);
and U17316 (N_17316,N_17192,N_17231);
nand U17317 (N_17317,N_17196,N_17063);
and U17318 (N_17318,N_17004,N_17151);
or U17319 (N_17319,N_17030,N_17024);
or U17320 (N_17320,N_17128,N_17044);
and U17321 (N_17321,N_17012,N_17122);
nor U17322 (N_17322,N_17002,N_17057);
and U17323 (N_17323,N_17091,N_17208);
and U17324 (N_17324,N_17072,N_17216);
nand U17325 (N_17325,N_17219,N_17075);
nand U17326 (N_17326,N_17184,N_17145);
and U17327 (N_17327,N_17037,N_17124);
nand U17328 (N_17328,N_17071,N_17020);
xor U17329 (N_17329,N_17211,N_17221);
nand U17330 (N_17330,N_17246,N_17243);
and U17331 (N_17331,N_17137,N_17181);
nand U17332 (N_17332,N_17147,N_17224);
xor U17333 (N_17333,N_17233,N_17126);
nor U17334 (N_17334,N_17095,N_17046);
and U17335 (N_17335,N_17021,N_17244);
and U17336 (N_17336,N_17227,N_17116);
xnor U17337 (N_17337,N_17228,N_17189);
xnor U17338 (N_17338,N_17179,N_17123);
nor U17339 (N_17339,N_17107,N_17134);
nand U17340 (N_17340,N_17144,N_17045);
xnor U17341 (N_17341,N_17235,N_17098);
and U17342 (N_17342,N_17080,N_17176);
nor U17343 (N_17343,N_17169,N_17059);
nor U17344 (N_17344,N_17060,N_17200);
nand U17345 (N_17345,N_17138,N_17047);
nor U17346 (N_17346,N_17212,N_17018);
and U17347 (N_17347,N_17041,N_17171);
nand U17348 (N_17348,N_17238,N_17131);
xor U17349 (N_17349,N_17245,N_17230);
and U17350 (N_17350,N_17050,N_17081);
xnor U17351 (N_17351,N_17052,N_17078);
or U17352 (N_17352,N_17093,N_17240);
or U17353 (N_17353,N_17180,N_17202);
or U17354 (N_17354,N_17040,N_17032);
nand U17355 (N_17355,N_17119,N_17086);
nor U17356 (N_17356,N_17247,N_17099);
xnor U17357 (N_17357,N_17132,N_17174);
nand U17358 (N_17358,N_17016,N_17096);
nor U17359 (N_17359,N_17206,N_17146);
nand U17360 (N_17360,N_17249,N_17161);
nand U17361 (N_17361,N_17165,N_17066);
nor U17362 (N_17362,N_17074,N_17076);
or U17363 (N_17363,N_17197,N_17003);
nand U17364 (N_17364,N_17215,N_17051);
or U17365 (N_17365,N_17105,N_17188);
and U17366 (N_17366,N_17065,N_17162);
nand U17367 (N_17367,N_17167,N_17183);
or U17368 (N_17368,N_17130,N_17100);
and U17369 (N_17369,N_17102,N_17175);
nor U17370 (N_17370,N_17150,N_17178);
nand U17371 (N_17371,N_17106,N_17195);
and U17372 (N_17372,N_17237,N_17019);
or U17373 (N_17373,N_17062,N_17148);
xnor U17374 (N_17374,N_17038,N_17015);
nor U17375 (N_17375,N_17037,N_17062);
or U17376 (N_17376,N_17045,N_17111);
nor U17377 (N_17377,N_17097,N_17192);
or U17378 (N_17378,N_17215,N_17241);
and U17379 (N_17379,N_17050,N_17142);
nand U17380 (N_17380,N_17075,N_17077);
nand U17381 (N_17381,N_17120,N_17177);
nand U17382 (N_17382,N_17119,N_17129);
nor U17383 (N_17383,N_17061,N_17075);
nand U17384 (N_17384,N_17104,N_17105);
nor U17385 (N_17385,N_17071,N_17047);
xnor U17386 (N_17386,N_17092,N_17091);
and U17387 (N_17387,N_17095,N_17243);
nor U17388 (N_17388,N_17197,N_17216);
and U17389 (N_17389,N_17215,N_17072);
nand U17390 (N_17390,N_17050,N_17159);
xnor U17391 (N_17391,N_17214,N_17144);
nand U17392 (N_17392,N_17221,N_17124);
xor U17393 (N_17393,N_17013,N_17183);
nand U17394 (N_17394,N_17022,N_17223);
xnor U17395 (N_17395,N_17189,N_17004);
nand U17396 (N_17396,N_17221,N_17038);
nor U17397 (N_17397,N_17178,N_17127);
or U17398 (N_17398,N_17137,N_17082);
and U17399 (N_17399,N_17214,N_17178);
or U17400 (N_17400,N_17068,N_17246);
or U17401 (N_17401,N_17158,N_17023);
nand U17402 (N_17402,N_17239,N_17126);
or U17403 (N_17403,N_17144,N_17149);
or U17404 (N_17404,N_17018,N_17114);
and U17405 (N_17405,N_17087,N_17186);
nor U17406 (N_17406,N_17080,N_17051);
and U17407 (N_17407,N_17095,N_17192);
or U17408 (N_17408,N_17009,N_17010);
xor U17409 (N_17409,N_17148,N_17185);
nand U17410 (N_17410,N_17142,N_17000);
nor U17411 (N_17411,N_17144,N_17118);
and U17412 (N_17412,N_17093,N_17111);
and U17413 (N_17413,N_17076,N_17233);
xor U17414 (N_17414,N_17093,N_17211);
xnor U17415 (N_17415,N_17229,N_17197);
or U17416 (N_17416,N_17166,N_17025);
or U17417 (N_17417,N_17007,N_17173);
or U17418 (N_17418,N_17184,N_17062);
or U17419 (N_17419,N_17195,N_17146);
and U17420 (N_17420,N_17171,N_17090);
nor U17421 (N_17421,N_17191,N_17108);
nand U17422 (N_17422,N_17219,N_17085);
nand U17423 (N_17423,N_17013,N_17195);
and U17424 (N_17424,N_17213,N_17173);
nand U17425 (N_17425,N_17070,N_17161);
nor U17426 (N_17426,N_17161,N_17219);
nor U17427 (N_17427,N_17154,N_17168);
nand U17428 (N_17428,N_17144,N_17016);
nand U17429 (N_17429,N_17031,N_17043);
nand U17430 (N_17430,N_17102,N_17200);
xnor U17431 (N_17431,N_17204,N_17160);
nor U17432 (N_17432,N_17242,N_17208);
or U17433 (N_17433,N_17028,N_17090);
nand U17434 (N_17434,N_17234,N_17108);
and U17435 (N_17435,N_17102,N_17203);
nor U17436 (N_17436,N_17014,N_17101);
xnor U17437 (N_17437,N_17075,N_17221);
or U17438 (N_17438,N_17195,N_17022);
xor U17439 (N_17439,N_17179,N_17012);
or U17440 (N_17440,N_17195,N_17154);
nor U17441 (N_17441,N_17115,N_17239);
xor U17442 (N_17442,N_17143,N_17247);
or U17443 (N_17443,N_17201,N_17115);
or U17444 (N_17444,N_17236,N_17004);
nor U17445 (N_17445,N_17089,N_17163);
nand U17446 (N_17446,N_17207,N_17010);
or U17447 (N_17447,N_17157,N_17049);
nand U17448 (N_17448,N_17230,N_17208);
or U17449 (N_17449,N_17173,N_17113);
or U17450 (N_17450,N_17000,N_17031);
nor U17451 (N_17451,N_17093,N_17183);
and U17452 (N_17452,N_17043,N_17216);
xor U17453 (N_17453,N_17015,N_17152);
xor U17454 (N_17454,N_17210,N_17064);
nand U17455 (N_17455,N_17203,N_17178);
nor U17456 (N_17456,N_17176,N_17221);
or U17457 (N_17457,N_17162,N_17231);
and U17458 (N_17458,N_17120,N_17116);
or U17459 (N_17459,N_17063,N_17213);
nand U17460 (N_17460,N_17134,N_17102);
and U17461 (N_17461,N_17144,N_17164);
or U17462 (N_17462,N_17230,N_17249);
nand U17463 (N_17463,N_17226,N_17184);
or U17464 (N_17464,N_17077,N_17058);
nor U17465 (N_17465,N_17203,N_17148);
or U17466 (N_17466,N_17054,N_17247);
xor U17467 (N_17467,N_17115,N_17221);
nand U17468 (N_17468,N_17128,N_17065);
or U17469 (N_17469,N_17119,N_17019);
nand U17470 (N_17470,N_17006,N_17143);
xnor U17471 (N_17471,N_17058,N_17200);
and U17472 (N_17472,N_17230,N_17039);
nor U17473 (N_17473,N_17176,N_17140);
and U17474 (N_17474,N_17201,N_17178);
and U17475 (N_17475,N_17167,N_17192);
or U17476 (N_17476,N_17101,N_17055);
or U17477 (N_17477,N_17075,N_17047);
and U17478 (N_17478,N_17029,N_17177);
nand U17479 (N_17479,N_17010,N_17042);
and U17480 (N_17480,N_17030,N_17022);
xor U17481 (N_17481,N_17091,N_17244);
and U17482 (N_17482,N_17045,N_17159);
nand U17483 (N_17483,N_17164,N_17191);
xor U17484 (N_17484,N_17002,N_17026);
xnor U17485 (N_17485,N_17209,N_17040);
xor U17486 (N_17486,N_17122,N_17206);
nand U17487 (N_17487,N_17167,N_17153);
nor U17488 (N_17488,N_17106,N_17086);
xnor U17489 (N_17489,N_17198,N_17142);
nor U17490 (N_17490,N_17077,N_17117);
xor U17491 (N_17491,N_17124,N_17123);
and U17492 (N_17492,N_17060,N_17000);
and U17493 (N_17493,N_17217,N_17162);
xor U17494 (N_17494,N_17051,N_17057);
xnor U17495 (N_17495,N_17198,N_17021);
or U17496 (N_17496,N_17027,N_17097);
and U17497 (N_17497,N_17225,N_17014);
nor U17498 (N_17498,N_17059,N_17016);
and U17499 (N_17499,N_17150,N_17129);
nand U17500 (N_17500,N_17385,N_17361);
nand U17501 (N_17501,N_17390,N_17287);
xor U17502 (N_17502,N_17270,N_17376);
nor U17503 (N_17503,N_17372,N_17290);
and U17504 (N_17504,N_17331,N_17264);
nor U17505 (N_17505,N_17320,N_17425);
nand U17506 (N_17506,N_17424,N_17415);
nor U17507 (N_17507,N_17493,N_17429);
and U17508 (N_17508,N_17260,N_17349);
xor U17509 (N_17509,N_17363,N_17337);
xor U17510 (N_17510,N_17457,N_17325);
nand U17511 (N_17511,N_17346,N_17366);
or U17512 (N_17512,N_17449,N_17381);
and U17513 (N_17513,N_17427,N_17255);
nand U17514 (N_17514,N_17259,N_17477);
nor U17515 (N_17515,N_17471,N_17265);
and U17516 (N_17516,N_17404,N_17402);
nor U17517 (N_17517,N_17343,N_17479);
xnor U17518 (N_17518,N_17269,N_17340);
xor U17519 (N_17519,N_17447,N_17304);
xor U17520 (N_17520,N_17485,N_17250);
nand U17521 (N_17521,N_17487,N_17309);
and U17522 (N_17522,N_17375,N_17461);
nor U17523 (N_17523,N_17489,N_17262);
xnor U17524 (N_17524,N_17319,N_17384);
nor U17525 (N_17525,N_17322,N_17383);
nor U17526 (N_17526,N_17444,N_17432);
nand U17527 (N_17527,N_17279,N_17339);
nor U17528 (N_17528,N_17408,N_17327);
nand U17529 (N_17529,N_17344,N_17464);
or U17530 (N_17530,N_17295,N_17365);
nand U17531 (N_17531,N_17296,N_17283);
nor U17532 (N_17532,N_17347,N_17379);
nand U17533 (N_17533,N_17303,N_17282);
and U17534 (N_17534,N_17266,N_17275);
nor U17535 (N_17535,N_17450,N_17488);
or U17536 (N_17536,N_17498,N_17333);
nand U17537 (N_17537,N_17434,N_17360);
nand U17538 (N_17538,N_17353,N_17435);
and U17539 (N_17539,N_17417,N_17418);
xor U17540 (N_17540,N_17368,N_17317);
nand U17541 (N_17541,N_17297,N_17356);
nand U17542 (N_17542,N_17367,N_17463);
nand U17543 (N_17543,N_17268,N_17336);
nor U17544 (N_17544,N_17284,N_17338);
nand U17545 (N_17545,N_17438,N_17314);
nand U17546 (N_17546,N_17332,N_17423);
xor U17547 (N_17547,N_17410,N_17403);
nor U17548 (N_17548,N_17495,N_17351);
nor U17549 (N_17549,N_17496,N_17451);
xnor U17550 (N_17550,N_17326,N_17292);
or U17551 (N_17551,N_17389,N_17380);
nand U17552 (N_17552,N_17345,N_17422);
xor U17553 (N_17553,N_17305,N_17302);
xor U17554 (N_17554,N_17378,N_17306);
and U17555 (N_17555,N_17342,N_17310);
nand U17556 (N_17556,N_17293,N_17377);
nor U17557 (N_17557,N_17452,N_17473);
or U17558 (N_17558,N_17370,N_17359);
and U17559 (N_17559,N_17459,N_17430);
xor U17560 (N_17560,N_17276,N_17469);
xor U17561 (N_17561,N_17362,N_17416);
and U17562 (N_17562,N_17455,N_17286);
and U17563 (N_17563,N_17396,N_17480);
and U17564 (N_17564,N_17492,N_17399);
nand U17565 (N_17565,N_17257,N_17474);
nand U17566 (N_17566,N_17273,N_17354);
xnor U17567 (N_17567,N_17288,N_17355);
nor U17568 (N_17568,N_17433,N_17482);
and U17569 (N_17569,N_17406,N_17407);
nor U17570 (N_17570,N_17400,N_17294);
nor U17571 (N_17571,N_17437,N_17419);
or U17572 (N_17572,N_17258,N_17280);
xor U17573 (N_17573,N_17312,N_17401);
and U17574 (N_17574,N_17478,N_17315);
nor U17575 (N_17575,N_17490,N_17484);
or U17576 (N_17576,N_17440,N_17335);
or U17577 (N_17577,N_17466,N_17373);
and U17578 (N_17578,N_17278,N_17443);
or U17579 (N_17579,N_17261,N_17470);
or U17580 (N_17580,N_17387,N_17454);
xnor U17581 (N_17581,N_17291,N_17420);
xor U17582 (N_17582,N_17300,N_17299);
or U17583 (N_17583,N_17395,N_17456);
nand U17584 (N_17584,N_17393,N_17446);
xnor U17585 (N_17585,N_17491,N_17431);
nand U17586 (N_17586,N_17272,N_17374);
and U17587 (N_17587,N_17394,N_17426);
or U17588 (N_17588,N_17442,N_17324);
xor U17589 (N_17589,N_17285,N_17298);
or U17590 (N_17590,N_17313,N_17301);
nand U17591 (N_17591,N_17369,N_17328);
and U17592 (N_17592,N_17357,N_17436);
xnor U17593 (N_17593,N_17318,N_17467);
xor U17594 (N_17594,N_17350,N_17392);
nor U17595 (N_17595,N_17271,N_17476);
xnor U17596 (N_17596,N_17251,N_17468);
nor U17597 (N_17597,N_17316,N_17254);
xor U17598 (N_17598,N_17475,N_17499);
or U17599 (N_17599,N_17462,N_17321);
nand U17600 (N_17600,N_17371,N_17307);
xnor U17601 (N_17601,N_17445,N_17414);
nand U17602 (N_17602,N_17364,N_17441);
or U17603 (N_17603,N_17323,N_17330);
nand U17604 (N_17604,N_17391,N_17409);
or U17605 (N_17605,N_17458,N_17334);
xnor U17606 (N_17606,N_17352,N_17281);
nor U17607 (N_17607,N_17494,N_17252);
xnor U17608 (N_17608,N_17439,N_17329);
and U17609 (N_17609,N_17358,N_17388);
xnor U17610 (N_17610,N_17460,N_17428);
and U17611 (N_17611,N_17472,N_17483);
or U17612 (N_17612,N_17308,N_17448);
nand U17613 (N_17613,N_17386,N_17411);
nand U17614 (N_17614,N_17348,N_17253);
nor U17615 (N_17615,N_17465,N_17497);
xor U17616 (N_17616,N_17398,N_17421);
and U17617 (N_17617,N_17413,N_17341);
and U17618 (N_17618,N_17289,N_17481);
nor U17619 (N_17619,N_17267,N_17382);
nor U17620 (N_17620,N_17486,N_17311);
nor U17621 (N_17621,N_17274,N_17412);
xor U17622 (N_17622,N_17277,N_17397);
and U17623 (N_17623,N_17256,N_17405);
nor U17624 (N_17624,N_17263,N_17453);
xor U17625 (N_17625,N_17359,N_17474);
and U17626 (N_17626,N_17256,N_17418);
nor U17627 (N_17627,N_17350,N_17493);
nor U17628 (N_17628,N_17293,N_17469);
nand U17629 (N_17629,N_17284,N_17354);
nand U17630 (N_17630,N_17311,N_17408);
or U17631 (N_17631,N_17294,N_17439);
nor U17632 (N_17632,N_17407,N_17378);
or U17633 (N_17633,N_17496,N_17399);
nand U17634 (N_17634,N_17476,N_17300);
or U17635 (N_17635,N_17435,N_17367);
or U17636 (N_17636,N_17472,N_17476);
and U17637 (N_17637,N_17444,N_17413);
xor U17638 (N_17638,N_17429,N_17284);
xnor U17639 (N_17639,N_17341,N_17284);
and U17640 (N_17640,N_17363,N_17472);
nor U17641 (N_17641,N_17271,N_17332);
nor U17642 (N_17642,N_17365,N_17492);
and U17643 (N_17643,N_17347,N_17384);
or U17644 (N_17644,N_17422,N_17421);
nor U17645 (N_17645,N_17429,N_17470);
xor U17646 (N_17646,N_17349,N_17338);
nor U17647 (N_17647,N_17471,N_17479);
xnor U17648 (N_17648,N_17419,N_17366);
or U17649 (N_17649,N_17423,N_17441);
nand U17650 (N_17650,N_17366,N_17458);
nor U17651 (N_17651,N_17286,N_17274);
nand U17652 (N_17652,N_17259,N_17257);
nand U17653 (N_17653,N_17333,N_17476);
or U17654 (N_17654,N_17312,N_17332);
and U17655 (N_17655,N_17493,N_17262);
nand U17656 (N_17656,N_17455,N_17260);
nand U17657 (N_17657,N_17378,N_17453);
xnor U17658 (N_17658,N_17431,N_17436);
nand U17659 (N_17659,N_17479,N_17484);
xor U17660 (N_17660,N_17396,N_17279);
nand U17661 (N_17661,N_17342,N_17433);
and U17662 (N_17662,N_17276,N_17279);
nor U17663 (N_17663,N_17453,N_17338);
nand U17664 (N_17664,N_17287,N_17486);
xor U17665 (N_17665,N_17317,N_17274);
xor U17666 (N_17666,N_17299,N_17394);
xnor U17667 (N_17667,N_17263,N_17288);
xnor U17668 (N_17668,N_17342,N_17455);
or U17669 (N_17669,N_17461,N_17441);
xor U17670 (N_17670,N_17343,N_17354);
nor U17671 (N_17671,N_17254,N_17412);
and U17672 (N_17672,N_17435,N_17375);
and U17673 (N_17673,N_17478,N_17338);
xnor U17674 (N_17674,N_17408,N_17334);
or U17675 (N_17675,N_17260,N_17470);
nor U17676 (N_17676,N_17261,N_17250);
and U17677 (N_17677,N_17357,N_17490);
nor U17678 (N_17678,N_17309,N_17340);
xnor U17679 (N_17679,N_17269,N_17464);
or U17680 (N_17680,N_17433,N_17462);
and U17681 (N_17681,N_17338,N_17446);
nand U17682 (N_17682,N_17279,N_17284);
xnor U17683 (N_17683,N_17364,N_17389);
and U17684 (N_17684,N_17278,N_17480);
and U17685 (N_17685,N_17301,N_17322);
nand U17686 (N_17686,N_17269,N_17421);
nor U17687 (N_17687,N_17395,N_17442);
xor U17688 (N_17688,N_17289,N_17297);
or U17689 (N_17689,N_17447,N_17289);
nand U17690 (N_17690,N_17355,N_17349);
nor U17691 (N_17691,N_17481,N_17342);
or U17692 (N_17692,N_17402,N_17337);
xor U17693 (N_17693,N_17445,N_17425);
and U17694 (N_17694,N_17255,N_17302);
and U17695 (N_17695,N_17499,N_17340);
and U17696 (N_17696,N_17298,N_17459);
or U17697 (N_17697,N_17341,N_17326);
and U17698 (N_17698,N_17331,N_17454);
xnor U17699 (N_17699,N_17482,N_17497);
or U17700 (N_17700,N_17455,N_17449);
nor U17701 (N_17701,N_17282,N_17487);
or U17702 (N_17702,N_17253,N_17441);
nand U17703 (N_17703,N_17341,N_17376);
xnor U17704 (N_17704,N_17268,N_17304);
or U17705 (N_17705,N_17269,N_17293);
nand U17706 (N_17706,N_17430,N_17432);
xnor U17707 (N_17707,N_17384,N_17340);
xnor U17708 (N_17708,N_17314,N_17268);
and U17709 (N_17709,N_17304,N_17497);
or U17710 (N_17710,N_17448,N_17257);
nand U17711 (N_17711,N_17283,N_17483);
nand U17712 (N_17712,N_17412,N_17260);
nor U17713 (N_17713,N_17359,N_17493);
xor U17714 (N_17714,N_17482,N_17284);
or U17715 (N_17715,N_17493,N_17377);
nand U17716 (N_17716,N_17283,N_17282);
xnor U17717 (N_17717,N_17274,N_17259);
nand U17718 (N_17718,N_17298,N_17386);
and U17719 (N_17719,N_17443,N_17305);
nor U17720 (N_17720,N_17321,N_17434);
nor U17721 (N_17721,N_17304,N_17342);
and U17722 (N_17722,N_17460,N_17380);
xnor U17723 (N_17723,N_17490,N_17251);
or U17724 (N_17724,N_17375,N_17296);
nand U17725 (N_17725,N_17372,N_17473);
xnor U17726 (N_17726,N_17480,N_17348);
and U17727 (N_17727,N_17264,N_17397);
xor U17728 (N_17728,N_17298,N_17266);
xor U17729 (N_17729,N_17367,N_17416);
nand U17730 (N_17730,N_17294,N_17265);
and U17731 (N_17731,N_17295,N_17279);
xnor U17732 (N_17732,N_17294,N_17260);
xor U17733 (N_17733,N_17427,N_17463);
nand U17734 (N_17734,N_17357,N_17440);
xnor U17735 (N_17735,N_17282,N_17333);
and U17736 (N_17736,N_17449,N_17395);
or U17737 (N_17737,N_17341,N_17307);
nor U17738 (N_17738,N_17291,N_17274);
nor U17739 (N_17739,N_17278,N_17498);
xor U17740 (N_17740,N_17459,N_17350);
and U17741 (N_17741,N_17433,N_17466);
nand U17742 (N_17742,N_17400,N_17302);
nand U17743 (N_17743,N_17404,N_17445);
nand U17744 (N_17744,N_17420,N_17276);
and U17745 (N_17745,N_17287,N_17355);
nand U17746 (N_17746,N_17480,N_17287);
nor U17747 (N_17747,N_17321,N_17373);
or U17748 (N_17748,N_17251,N_17375);
or U17749 (N_17749,N_17385,N_17271);
nor U17750 (N_17750,N_17749,N_17591);
and U17751 (N_17751,N_17583,N_17532);
and U17752 (N_17752,N_17562,N_17659);
nand U17753 (N_17753,N_17622,N_17740);
nor U17754 (N_17754,N_17597,N_17525);
nand U17755 (N_17755,N_17539,N_17556);
xor U17756 (N_17756,N_17601,N_17733);
nor U17757 (N_17757,N_17743,N_17720);
or U17758 (N_17758,N_17676,N_17746);
and U17759 (N_17759,N_17508,N_17538);
nor U17760 (N_17760,N_17579,N_17585);
nand U17761 (N_17761,N_17633,N_17594);
nand U17762 (N_17762,N_17645,N_17501);
nand U17763 (N_17763,N_17542,N_17576);
nor U17764 (N_17764,N_17515,N_17714);
and U17765 (N_17765,N_17735,N_17516);
xor U17766 (N_17766,N_17521,N_17653);
nor U17767 (N_17767,N_17624,N_17702);
and U17768 (N_17768,N_17552,N_17719);
and U17769 (N_17769,N_17565,N_17745);
and U17770 (N_17770,N_17514,N_17674);
xor U17771 (N_17771,N_17736,N_17707);
nand U17772 (N_17772,N_17685,N_17711);
nand U17773 (N_17773,N_17600,N_17741);
nand U17774 (N_17774,N_17681,N_17502);
xnor U17775 (N_17775,N_17587,N_17662);
nand U17776 (N_17776,N_17527,N_17713);
and U17777 (N_17777,N_17543,N_17620);
nand U17778 (N_17778,N_17715,N_17709);
or U17779 (N_17779,N_17545,N_17544);
and U17780 (N_17780,N_17573,N_17505);
nor U17781 (N_17781,N_17560,N_17548);
and U17782 (N_17782,N_17522,N_17626);
and U17783 (N_17783,N_17574,N_17533);
and U17784 (N_17784,N_17666,N_17649);
nor U17785 (N_17785,N_17553,N_17596);
or U17786 (N_17786,N_17535,N_17717);
xnor U17787 (N_17787,N_17716,N_17647);
nand U17788 (N_17788,N_17689,N_17684);
xor U17789 (N_17789,N_17584,N_17517);
and U17790 (N_17790,N_17621,N_17593);
xnor U17791 (N_17791,N_17657,N_17555);
nand U17792 (N_17792,N_17729,N_17737);
nand U17793 (N_17793,N_17682,N_17531);
or U17794 (N_17794,N_17726,N_17605);
nor U17795 (N_17795,N_17558,N_17683);
nand U17796 (N_17796,N_17500,N_17569);
and U17797 (N_17797,N_17698,N_17612);
nor U17798 (N_17798,N_17547,N_17615);
nand U17799 (N_17799,N_17526,N_17665);
xor U17800 (N_17800,N_17701,N_17744);
nor U17801 (N_17801,N_17634,N_17732);
and U17802 (N_17802,N_17642,N_17678);
xnor U17803 (N_17803,N_17534,N_17655);
nand U17804 (N_17804,N_17567,N_17673);
xor U17805 (N_17805,N_17710,N_17667);
nand U17806 (N_17806,N_17523,N_17725);
nor U17807 (N_17807,N_17581,N_17616);
xnor U17808 (N_17808,N_17513,N_17672);
or U17809 (N_17809,N_17690,N_17618);
and U17810 (N_17810,N_17561,N_17656);
xnor U17811 (N_17811,N_17648,N_17660);
and U17812 (N_17812,N_17510,N_17602);
nor U17813 (N_17813,N_17646,N_17727);
and U17814 (N_17814,N_17632,N_17731);
and U17815 (N_17815,N_17705,N_17747);
or U17816 (N_17816,N_17704,N_17703);
and U17817 (N_17817,N_17628,N_17699);
nor U17818 (N_17818,N_17603,N_17636);
nand U17819 (N_17819,N_17688,N_17519);
and U17820 (N_17820,N_17518,N_17650);
and U17821 (N_17821,N_17693,N_17595);
and U17822 (N_17822,N_17658,N_17619);
or U17823 (N_17823,N_17564,N_17611);
xor U17824 (N_17824,N_17580,N_17638);
or U17825 (N_17825,N_17609,N_17586);
nand U17826 (N_17826,N_17694,N_17623);
and U17827 (N_17827,N_17604,N_17568);
nand U17828 (N_17828,N_17520,N_17550);
or U17829 (N_17829,N_17570,N_17546);
nor U17830 (N_17830,N_17738,N_17697);
xor U17831 (N_17831,N_17509,N_17652);
nor U17832 (N_17832,N_17669,N_17617);
and U17833 (N_17833,N_17629,N_17578);
and U17834 (N_17834,N_17692,N_17577);
and U17835 (N_17835,N_17563,N_17696);
nand U17836 (N_17836,N_17507,N_17748);
nor U17837 (N_17837,N_17549,N_17721);
or U17838 (N_17838,N_17512,N_17686);
or U17839 (N_17839,N_17588,N_17599);
or U17840 (N_17840,N_17530,N_17575);
and U17841 (N_17841,N_17559,N_17613);
or U17842 (N_17842,N_17635,N_17722);
nand U17843 (N_17843,N_17718,N_17610);
nor U17844 (N_17844,N_17644,N_17506);
nand U17845 (N_17845,N_17708,N_17592);
xnor U17846 (N_17846,N_17503,N_17723);
nor U17847 (N_17847,N_17641,N_17691);
or U17848 (N_17848,N_17557,N_17566);
or U17849 (N_17849,N_17728,N_17631);
and U17850 (N_17850,N_17571,N_17554);
nand U17851 (N_17851,N_17541,N_17661);
xor U17852 (N_17852,N_17643,N_17677);
nand U17853 (N_17853,N_17536,N_17630);
or U17854 (N_17854,N_17606,N_17695);
nor U17855 (N_17855,N_17734,N_17529);
or U17856 (N_17856,N_17687,N_17664);
nor U17857 (N_17857,N_17675,N_17504);
or U17858 (N_17858,N_17654,N_17551);
or U17859 (N_17859,N_17625,N_17589);
nor U17860 (N_17860,N_17679,N_17608);
nand U17861 (N_17861,N_17670,N_17671);
nor U17862 (N_17862,N_17524,N_17739);
or U17863 (N_17863,N_17639,N_17706);
nand U17864 (N_17864,N_17742,N_17651);
xnor U17865 (N_17865,N_17663,N_17712);
or U17866 (N_17866,N_17540,N_17640);
and U17867 (N_17867,N_17637,N_17614);
and U17868 (N_17868,N_17582,N_17607);
and U17869 (N_17869,N_17724,N_17590);
and U17870 (N_17870,N_17598,N_17700);
nor U17871 (N_17871,N_17528,N_17730);
and U17872 (N_17872,N_17537,N_17511);
nand U17873 (N_17873,N_17668,N_17572);
or U17874 (N_17874,N_17627,N_17680);
or U17875 (N_17875,N_17572,N_17705);
or U17876 (N_17876,N_17618,N_17686);
xnor U17877 (N_17877,N_17557,N_17626);
nand U17878 (N_17878,N_17679,N_17552);
xor U17879 (N_17879,N_17705,N_17679);
and U17880 (N_17880,N_17713,N_17534);
xnor U17881 (N_17881,N_17671,N_17572);
nor U17882 (N_17882,N_17605,N_17636);
or U17883 (N_17883,N_17649,N_17567);
xnor U17884 (N_17884,N_17728,N_17632);
nand U17885 (N_17885,N_17743,N_17614);
and U17886 (N_17886,N_17742,N_17511);
nand U17887 (N_17887,N_17512,N_17714);
nand U17888 (N_17888,N_17719,N_17712);
xor U17889 (N_17889,N_17724,N_17653);
nand U17890 (N_17890,N_17637,N_17699);
xor U17891 (N_17891,N_17559,N_17525);
nand U17892 (N_17892,N_17619,N_17690);
nand U17893 (N_17893,N_17596,N_17602);
and U17894 (N_17894,N_17564,N_17664);
nand U17895 (N_17895,N_17730,N_17603);
or U17896 (N_17896,N_17500,N_17572);
nor U17897 (N_17897,N_17527,N_17586);
nand U17898 (N_17898,N_17619,N_17566);
xnor U17899 (N_17899,N_17694,N_17717);
nor U17900 (N_17900,N_17504,N_17679);
nor U17901 (N_17901,N_17735,N_17636);
and U17902 (N_17902,N_17585,N_17565);
xor U17903 (N_17903,N_17659,N_17709);
nand U17904 (N_17904,N_17507,N_17554);
and U17905 (N_17905,N_17615,N_17710);
and U17906 (N_17906,N_17600,N_17594);
nor U17907 (N_17907,N_17539,N_17746);
nor U17908 (N_17908,N_17552,N_17676);
nor U17909 (N_17909,N_17719,N_17662);
and U17910 (N_17910,N_17575,N_17520);
nor U17911 (N_17911,N_17588,N_17511);
or U17912 (N_17912,N_17713,N_17577);
xnor U17913 (N_17913,N_17627,N_17746);
nor U17914 (N_17914,N_17540,N_17546);
xor U17915 (N_17915,N_17502,N_17748);
nor U17916 (N_17916,N_17627,N_17607);
or U17917 (N_17917,N_17728,N_17738);
nand U17918 (N_17918,N_17724,N_17726);
and U17919 (N_17919,N_17590,N_17744);
xor U17920 (N_17920,N_17572,N_17686);
nand U17921 (N_17921,N_17561,N_17558);
or U17922 (N_17922,N_17688,N_17549);
nand U17923 (N_17923,N_17532,N_17721);
nor U17924 (N_17924,N_17547,N_17677);
and U17925 (N_17925,N_17517,N_17641);
nand U17926 (N_17926,N_17598,N_17717);
nor U17927 (N_17927,N_17644,N_17730);
nor U17928 (N_17928,N_17697,N_17634);
or U17929 (N_17929,N_17585,N_17718);
or U17930 (N_17930,N_17602,N_17627);
and U17931 (N_17931,N_17565,N_17550);
or U17932 (N_17932,N_17652,N_17583);
and U17933 (N_17933,N_17670,N_17741);
nor U17934 (N_17934,N_17505,N_17658);
nor U17935 (N_17935,N_17572,N_17667);
and U17936 (N_17936,N_17501,N_17582);
nand U17937 (N_17937,N_17629,N_17545);
nand U17938 (N_17938,N_17614,N_17671);
xor U17939 (N_17939,N_17604,N_17534);
or U17940 (N_17940,N_17659,N_17657);
or U17941 (N_17941,N_17662,N_17532);
xnor U17942 (N_17942,N_17702,N_17623);
nor U17943 (N_17943,N_17680,N_17602);
nand U17944 (N_17944,N_17704,N_17533);
nand U17945 (N_17945,N_17693,N_17533);
and U17946 (N_17946,N_17544,N_17672);
nand U17947 (N_17947,N_17501,N_17638);
nor U17948 (N_17948,N_17581,N_17590);
and U17949 (N_17949,N_17732,N_17573);
and U17950 (N_17950,N_17700,N_17577);
xor U17951 (N_17951,N_17603,N_17605);
or U17952 (N_17952,N_17663,N_17535);
or U17953 (N_17953,N_17610,N_17708);
and U17954 (N_17954,N_17637,N_17573);
xor U17955 (N_17955,N_17632,N_17553);
nand U17956 (N_17956,N_17557,N_17558);
and U17957 (N_17957,N_17667,N_17577);
nand U17958 (N_17958,N_17702,N_17606);
xnor U17959 (N_17959,N_17545,N_17619);
nand U17960 (N_17960,N_17670,N_17594);
nand U17961 (N_17961,N_17576,N_17604);
and U17962 (N_17962,N_17566,N_17598);
nor U17963 (N_17963,N_17639,N_17556);
or U17964 (N_17964,N_17675,N_17559);
or U17965 (N_17965,N_17712,N_17540);
and U17966 (N_17966,N_17724,N_17528);
and U17967 (N_17967,N_17605,N_17567);
and U17968 (N_17968,N_17749,N_17728);
xnor U17969 (N_17969,N_17572,N_17719);
and U17970 (N_17970,N_17699,N_17688);
nor U17971 (N_17971,N_17727,N_17654);
nor U17972 (N_17972,N_17685,N_17581);
or U17973 (N_17973,N_17633,N_17644);
and U17974 (N_17974,N_17735,N_17597);
nor U17975 (N_17975,N_17509,N_17545);
or U17976 (N_17976,N_17574,N_17597);
nand U17977 (N_17977,N_17641,N_17532);
nor U17978 (N_17978,N_17734,N_17630);
xor U17979 (N_17979,N_17517,N_17725);
and U17980 (N_17980,N_17521,N_17635);
nor U17981 (N_17981,N_17741,N_17651);
nor U17982 (N_17982,N_17605,N_17660);
nor U17983 (N_17983,N_17716,N_17541);
or U17984 (N_17984,N_17706,N_17561);
and U17985 (N_17985,N_17599,N_17671);
xnor U17986 (N_17986,N_17725,N_17616);
nor U17987 (N_17987,N_17600,N_17521);
or U17988 (N_17988,N_17612,N_17682);
nor U17989 (N_17989,N_17545,N_17521);
xnor U17990 (N_17990,N_17650,N_17605);
nand U17991 (N_17991,N_17505,N_17659);
nand U17992 (N_17992,N_17598,N_17719);
or U17993 (N_17993,N_17681,N_17735);
and U17994 (N_17994,N_17748,N_17711);
nand U17995 (N_17995,N_17673,N_17542);
nand U17996 (N_17996,N_17627,N_17679);
or U17997 (N_17997,N_17511,N_17523);
nor U17998 (N_17998,N_17590,N_17532);
or U17999 (N_17999,N_17723,N_17583);
and U18000 (N_18000,N_17845,N_17842);
nor U18001 (N_18001,N_17753,N_17999);
nand U18002 (N_18002,N_17987,N_17764);
nor U18003 (N_18003,N_17866,N_17936);
nor U18004 (N_18004,N_17826,N_17769);
nor U18005 (N_18005,N_17966,N_17953);
or U18006 (N_18006,N_17807,N_17766);
xnor U18007 (N_18007,N_17939,N_17955);
or U18008 (N_18008,N_17831,N_17924);
or U18009 (N_18009,N_17948,N_17872);
or U18010 (N_18010,N_17762,N_17930);
and U18011 (N_18011,N_17781,N_17993);
xor U18012 (N_18012,N_17771,N_17963);
xnor U18013 (N_18013,N_17787,N_17756);
xnor U18014 (N_18014,N_17919,N_17829);
nand U18015 (N_18015,N_17864,N_17871);
nor U18016 (N_18016,N_17933,N_17915);
nor U18017 (N_18017,N_17759,N_17757);
nand U18018 (N_18018,N_17921,N_17954);
nor U18019 (N_18019,N_17931,N_17946);
xnor U18020 (N_18020,N_17980,N_17902);
nand U18021 (N_18021,N_17794,N_17814);
nand U18022 (N_18022,N_17976,N_17777);
and U18023 (N_18023,N_17832,N_17834);
nand U18024 (N_18024,N_17882,N_17891);
nand U18025 (N_18025,N_17887,N_17994);
and U18026 (N_18026,N_17860,N_17925);
xnor U18027 (N_18027,N_17827,N_17808);
nor U18028 (N_18028,N_17984,N_17959);
and U18029 (N_18029,N_17960,N_17815);
or U18030 (N_18030,N_17935,N_17788);
nand U18031 (N_18031,N_17750,N_17928);
xnor U18032 (N_18032,N_17922,N_17792);
nand U18033 (N_18033,N_17983,N_17811);
nor U18034 (N_18034,N_17947,N_17877);
or U18035 (N_18035,N_17818,N_17893);
nor U18036 (N_18036,N_17982,N_17810);
xor U18037 (N_18037,N_17837,N_17909);
xor U18038 (N_18038,N_17790,N_17995);
or U18039 (N_18039,N_17956,N_17835);
or U18040 (N_18040,N_17853,N_17758);
and U18041 (N_18041,N_17836,N_17906);
nor U18042 (N_18042,N_17961,N_17817);
and U18043 (N_18043,N_17772,N_17949);
xor U18044 (N_18044,N_17791,N_17876);
xor U18045 (N_18045,N_17868,N_17912);
nand U18046 (N_18046,N_17997,N_17800);
nand U18047 (N_18047,N_17819,N_17805);
nor U18048 (N_18048,N_17934,N_17768);
or U18049 (N_18049,N_17784,N_17825);
nor U18050 (N_18050,N_17973,N_17820);
xnor U18051 (N_18051,N_17850,N_17920);
nand U18052 (N_18052,N_17904,N_17867);
or U18053 (N_18053,N_17978,N_17824);
nor U18054 (N_18054,N_17856,N_17752);
nor U18055 (N_18055,N_17918,N_17884);
and U18056 (N_18056,N_17962,N_17754);
xnor U18057 (N_18057,N_17943,N_17965);
or U18058 (N_18058,N_17843,N_17861);
or U18059 (N_18059,N_17958,N_17970);
nor U18060 (N_18060,N_17760,N_17951);
or U18061 (N_18061,N_17763,N_17900);
nor U18062 (N_18062,N_17917,N_17989);
nand U18063 (N_18063,N_17780,N_17879);
nand U18064 (N_18064,N_17975,N_17940);
and U18065 (N_18065,N_17991,N_17941);
nor U18066 (N_18066,N_17896,N_17926);
or U18067 (N_18067,N_17968,N_17767);
and U18068 (N_18068,N_17981,N_17778);
nor U18069 (N_18069,N_17913,N_17839);
nor U18070 (N_18070,N_17992,N_17775);
nor U18071 (N_18071,N_17770,N_17806);
xor U18072 (N_18072,N_17899,N_17849);
xnor U18073 (N_18073,N_17971,N_17952);
and U18074 (N_18074,N_17886,N_17932);
or U18075 (N_18075,N_17789,N_17785);
nor U18076 (N_18076,N_17841,N_17793);
nor U18077 (N_18077,N_17897,N_17911);
and U18078 (N_18078,N_17802,N_17916);
nand U18079 (N_18079,N_17964,N_17873);
nand U18080 (N_18080,N_17822,N_17799);
nor U18081 (N_18081,N_17852,N_17828);
nor U18082 (N_18082,N_17874,N_17990);
nor U18083 (N_18083,N_17977,N_17858);
xnor U18084 (N_18084,N_17972,N_17796);
or U18085 (N_18085,N_17844,N_17988);
and U18086 (N_18086,N_17929,N_17797);
and U18087 (N_18087,N_17945,N_17863);
nor U18088 (N_18088,N_17798,N_17821);
or U18089 (N_18089,N_17927,N_17950);
or U18090 (N_18090,N_17782,N_17998);
and U18091 (N_18091,N_17881,N_17908);
or U18092 (N_18092,N_17880,N_17944);
nor U18093 (N_18093,N_17795,N_17986);
nor U18094 (N_18094,N_17903,N_17967);
nand U18095 (N_18095,N_17761,N_17783);
nand U18096 (N_18096,N_17957,N_17830);
nand U18097 (N_18097,N_17895,N_17854);
or U18098 (N_18098,N_17883,N_17996);
or U18099 (N_18099,N_17812,N_17801);
and U18100 (N_18100,N_17985,N_17969);
nand U18101 (N_18101,N_17938,N_17755);
nor U18102 (N_18102,N_17823,N_17846);
nand U18103 (N_18103,N_17776,N_17765);
or U18104 (N_18104,N_17905,N_17859);
xnor U18105 (N_18105,N_17898,N_17833);
and U18106 (N_18106,N_17979,N_17890);
or U18107 (N_18107,N_17809,N_17894);
nand U18108 (N_18108,N_17875,N_17914);
xor U18109 (N_18109,N_17774,N_17847);
nand U18110 (N_18110,N_17974,N_17813);
or U18111 (N_18111,N_17942,N_17869);
or U18112 (N_18112,N_17803,N_17816);
nor U18113 (N_18113,N_17910,N_17892);
xor U18114 (N_18114,N_17751,N_17889);
and U18115 (N_18115,N_17870,N_17840);
and U18116 (N_18116,N_17865,N_17773);
xor U18117 (N_18117,N_17878,N_17786);
xor U18118 (N_18118,N_17779,N_17804);
and U18119 (N_18119,N_17888,N_17848);
xor U18120 (N_18120,N_17907,N_17851);
nor U18121 (N_18121,N_17838,N_17855);
xnor U18122 (N_18122,N_17901,N_17862);
nand U18123 (N_18123,N_17937,N_17885);
nand U18124 (N_18124,N_17923,N_17857);
nor U18125 (N_18125,N_17929,N_17763);
or U18126 (N_18126,N_17922,N_17818);
nor U18127 (N_18127,N_17896,N_17766);
nor U18128 (N_18128,N_17767,N_17948);
nand U18129 (N_18129,N_17816,N_17751);
or U18130 (N_18130,N_17931,N_17894);
nand U18131 (N_18131,N_17775,N_17805);
or U18132 (N_18132,N_17850,N_17796);
nor U18133 (N_18133,N_17846,N_17955);
and U18134 (N_18134,N_17918,N_17797);
nand U18135 (N_18135,N_17765,N_17971);
nor U18136 (N_18136,N_17768,N_17805);
nor U18137 (N_18137,N_17859,N_17834);
xnor U18138 (N_18138,N_17920,N_17941);
nor U18139 (N_18139,N_17969,N_17807);
nand U18140 (N_18140,N_17886,N_17950);
nor U18141 (N_18141,N_17767,N_17840);
or U18142 (N_18142,N_17966,N_17786);
nand U18143 (N_18143,N_17841,N_17809);
or U18144 (N_18144,N_17909,N_17817);
or U18145 (N_18145,N_17961,N_17844);
nand U18146 (N_18146,N_17966,N_17895);
or U18147 (N_18147,N_17933,N_17753);
nor U18148 (N_18148,N_17773,N_17821);
and U18149 (N_18149,N_17890,N_17962);
xnor U18150 (N_18150,N_17900,N_17813);
or U18151 (N_18151,N_17822,N_17827);
and U18152 (N_18152,N_17825,N_17947);
nor U18153 (N_18153,N_17979,N_17907);
or U18154 (N_18154,N_17925,N_17868);
nand U18155 (N_18155,N_17977,N_17979);
and U18156 (N_18156,N_17963,N_17809);
nand U18157 (N_18157,N_17984,N_17927);
or U18158 (N_18158,N_17896,N_17936);
nand U18159 (N_18159,N_17769,N_17968);
xnor U18160 (N_18160,N_17766,N_17921);
and U18161 (N_18161,N_17936,N_17874);
or U18162 (N_18162,N_17959,N_17901);
and U18163 (N_18163,N_17998,N_17901);
and U18164 (N_18164,N_17929,N_17838);
or U18165 (N_18165,N_17823,N_17930);
or U18166 (N_18166,N_17891,N_17938);
nand U18167 (N_18167,N_17867,N_17944);
nand U18168 (N_18168,N_17963,N_17871);
or U18169 (N_18169,N_17929,N_17988);
and U18170 (N_18170,N_17883,N_17974);
nand U18171 (N_18171,N_17919,N_17962);
nand U18172 (N_18172,N_17987,N_17962);
nor U18173 (N_18173,N_17954,N_17925);
and U18174 (N_18174,N_17817,N_17887);
or U18175 (N_18175,N_17786,N_17936);
nor U18176 (N_18176,N_17773,N_17973);
nor U18177 (N_18177,N_17825,N_17853);
nand U18178 (N_18178,N_17807,N_17765);
nor U18179 (N_18179,N_17952,N_17947);
nand U18180 (N_18180,N_17820,N_17986);
nor U18181 (N_18181,N_17919,N_17800);
or U18182 (N_18182,N_17958,N_17803);
or U18183 (N_18183,N_17868,N_17776);
nand U18184 (N_18184,N_17926,N_17786);
nor U18185 (N_18185,N_17879,N_17947);
nand U18186 (N_18186,N_17912,N_17903);
or U18187 (N_18187,N_17949,N_17877);
nand U18188 (N_18188,N_17986,N_17840);
or U18189 (N_18189,N_17809,N_17967);
or U18190 (N_18190,N_17929,N_17912);
and U18191 (N_18191,N_17938,N_17825);
nand U18192 (N_18192,N_17750,N_17895);
nand U18193 (N_18193,N_17994,N_17842);
xnor U18194 (N_18194,N_17927,N_17754);
xnor U18195 (N_18195,N_17890,N_17867);
xor U18196 (N_18196,N_17846,N_17924);
nor U18197 (N_18197,N_17865,N_17939);
nand U18198 (N_18198,N_17932,N_17984);
and U18199 (N_18199,N_17982,N_17913);
nand U18200 (N_18200,N_17855,N_17963);
nor U18201 (N_18201,N_17782,N_17996);
and U18202 (N_18202,N_17884,N_17972);
and U18203 (N_18203,N_17998,N_17978);
nand U18204 (N_18204,N_17918,N_17988);
nand U18205 (N_18205,N_17888,N_17882);
xor U18206 (N_18206,N_17827,N_17897);
and U18207 (N_18207,N_17883,N_17871);
or U18208 (N_18208,N_17882,N_17908);
or U18209 (N_18209,N_17761,N_17932);
nand U18210 (N_18210,N_17979,N_17778);
or U18211 (N_18211,N_17776,N_17999);
nand U18212 (N_18212,N_17754,N_17961);
nand U18213 (N_18213,N_17860,N_17958);
nor U18214 (N_18214,N_17995,N_17834);
nor U18215 (N_18215,N_17955,N_17913);
nand U18216 (N_18216,N_17772,N_17777);
or U18217 (N_18217,N_17770,N_17754);
nand U18218 (N_18218,N_17871,N_17913);
xnor U18219 (N_18219,N_17904,N_17851);
or U18220 (N_18220,N_17769,N_17791);
xor U18221 (N_18221,N_17870,N_17805);
nor U18222 (N_18222,N_17884,N_17883);
nor U18223 (N_18223,N_17851,N_17996);
nor U18224 (N_18224,N_17862,N_17910);
xnor U18225 (N_18225,N_17798,N_17764);
nor U18226 (N_18226,N_17755,N_17945);
and U18227 (N_18227,N_17891,N_17775);
xor U18228 (N_18228,N_17846,N_17803);
nand U18229 (N_18229,N_17885,N_17820);
nor U18230 (N_18230,N_17798,N_17951);
xnor U18231 (N_18231,N_17981,N_17953);
or U18232 (N_18232,N_17760,N_17778);
nand U18233 (N_18233,N_17805,N_17838);
and U18234 (N_18234,N_17765,N_17988);
and U18235 (N_18235,N_17811,N_17992);
nand U18236 (N_18236,N_17754,N_17970);
nand U18237 (N_18237,N_17796,N_17867);
and U18238 (N_18238,N_17847,N_17975);
and U18239 (N_18239,N_17760,N_17923);
or U18240 (N_18240,N_17816,N_17989);
nand U18241 (N_18241,N_17826,N_17810);
and U18242 (N_18242,N_17772,N_17801);
and U18243 (N_18243,N_17815,N_17810);
or U18244 (N_18244,N_17786,N_17834);
and U18245 (N_18245,N_17775,N_17993);
nand U18246 (N_18246,N_17920,N_17767);
xnor U18247 (N_18247,N_17871,N_17912);
nand U18248 (N_18248,N_17948,N_17907);
or U18249 (N_18249,N_17960,N_17862);
nor U18250 (N_18250,N_18057,N_18034);
xor U18251 (N_18251,N_18113,N_18180);
nand U18252 (N_18252,N_18004,N_18242);
and U18253 (N_18253,N_18212,N_18111);
and U18254 (N_18254,N_18229,N_18020);
or U18255 (N_18255,N_18134,N_18064);
and U18256 (N_18256,N_18219,N_18037);
xnor U18257 (N_18257,N_18070,N_18237);
nand U18258 (N_18258,N_18213,N_18231);
nor U18259 (N_18259,N_18179,N_18077);
nor U18260 (N_18260,N_18071,N_18010);
and U18261 (N_18261,N_18118,N_18066);
nand U18262 (N_18262,N_18052,N_18218);
and U18263 (N_18263,N_18008,N_18209);
or U18264 (N_18264,N_18076,N_18097);
and U18265 (N_18265,N_18226,N_18177);
or U18266 (N_18266,N_18173,N_18043);
nor U18267 (N_18267,N_18027,N_18083);
xnor U18268 (N_18268,N_18195,N_18090);
xor U18269 (N_18269,N_18046,N_18061);
nor U18270 (N_18270,N_18028,N_18187);
and U18271 (N_18271,N_18102,N_18155);
and U18272 (N_18272,N_18072,N_18192);
and U18273 (N_18273,N_18031,N_18082);
and U18274 (N_18274,N_18205,N_18060);
xor U18275 (N_18275,N_18156,N_18148);
nor U18276 (N_18276,N_18200,N_18087);
and U18277 (N_18277,N_18021,N_18171);
or U18278 (N_18278,N_18005,N_18119);
xor U18279 (N_18279,N_18085,N_18048);
nor U18280 (N_18280,N_18032,N_18074);
nor U18281 (N_18281,N_18249,N_18240);
nor U18282 (N_18282,N_18128,N_18065);
nand U18283 (N_18283,N_18232,N_18116);
nand U18284 (N_18284,N_18172,N_18185);
or U18285 (N_18285,N_18035,N_18112);
or U18286 (N_18286,N_18132,N_18103);
nor U18287 (N_18287,N_18024,N_18106);
nor U18288 (N_18288,N_18091,N_18135);
nor U18289 (N_18289,N_18093,N_18176);
nor U18290 (N_18290,N_18063,N_18001);
nand U18291 (N_18291,N_18053,N_18007);
nor U18292 (N_18292,N_18150,N_18041);
or U18293 (N_18293,N_18207,N_18055);
xor U18294 (N_18294,N_18015,N_18158);
and U18295 (N_18295,N_18220,N_18095);
or U18296 (N_18296,N_18023,N_18164);
or U18297 (N_18297,N_18030,N_18166);
nor U18298 (N_18298,N_18012,N_18115);
or U18299 (N_18299,N_18243,N_18058);
nand U18300 (N_18300,N_18040,N_18157);
and U18301 (N_18301,N_18216,N_18109);
and U18302 (N_18302,N_18126,N_18182);
nor U18303 (N_18303,N_18038,N_18107);
xor U18304 (N_18304,N_18086,N_18002);
nand U18305 (N_18305,N_18227,N_18017);
nor U18306 (N_18306,N_18245,N_18140);
and U18307 (N_18307,N_18047,N_18141);
and U18308 (N_18308,N_18153,N_18121);
nand U18309 (N_18309,N_18014,N_18206);
or U18310 (N_18310,N_18248,N_18143);
nand U18311 (N_18311,N_18122,N_18186);
or U18312 (N_18312,N_18105,N_18241);
xnor U18313 (N_18313,N_18168,N_18025);
nand U18314 (N_18314,N_18050,N_18049);
nand U18315 (N_18315,N_18127,N_18099);
xnor U18316 (N_18316,N_18003,N_18018);
xnor U18317 (N_18317,N_18051,N_18224);
and U18318 (N_18318,N_18045,N_18145);
xor U18319 (N_18319,N_18190,N_18165);
or U18320 (N_18320,N_18221,N_18006);
and U18321 (N_18321,N_18081,N_18144);
or U18322 (N_18322,N_18230,N_18170);
and U18323 (N_18323,N_18191,N_18120);
nand U18324 (N_18324,N_18042,N_18110);
nor U18325 (N_18325,N_18100,N_18247);
xor U18326 (N_18326,N_18246,N_18201);
nand U18327 (N_18327,N_18033,N_18183);
or U18328 (N_18328,N_18142,N_18210);
or U18329 (N_18329,N_18022,N_18215);
or U18330 (N_18330,N_18084,N_18181);
and U18331 (N_18331,N_18124,N_18096);
xor U18332 (N_18332,N_18234,N_18197);
or U18333 (N_18333,N_18152,N_18235);
nor U18334 (N_18334,N_18089,N_18189);
nor U18335 (N_18335,N_18188,N_18238);
xor U18336 (N_18336,N_18092,N_18088);
xor U18337 (N_18337,N_18009,N_18178);
and U18338 (N_18338,N_18069,N_18101);
xor U18339 (N_18339,N_18067,N_18167);
nor U18340 (N_18340,N_18075,N_18016);
or U18341 (N_18341,N_18214,N_18094);
nand U18342 (N_18342,N_18223,N_18013);
and U18343 (N_18343,N_18133,N_18117);
or U18344 (N_18344,N_18217,N_18211);
nand U18345 (N_18345,N_18199,N_18080);
xor U18346 (N_18346,N_18062,N_18149);
and U18347 (N_18347,N_18138,N_18203);
nand U18348 (N_18348,N_18114,N_18159);
or U18349 (N_18349,N_18125,N_18160);
nand U18350 (N_18350,N_18073,N_18151);
or U18351 (N_18351,N_18054,N_18161);
and U18352 (N_18352,N_18225,N_18162);
nand U18353 (N_18353,N_18233,N_18154);
or U18354 (N_18354,N_18194,N_18131);
nand U18355 (N_18355,N_18000,N_18036);
or U18356 (N_18356,N_18239,N_18222);
xor U18357 (N_18357,N_18026,N_18130);
or U18358 (N_18358,N_18011,N_18068);
or U18359 (N_18359,N_18136,N_18202);
nand U18360 (N_18360,N_18196,N_18098);
nand U18361 (N_18361,N_18146,N_18056);
xor U18362 (N_18362,N_18059,N_18078);
nand U18363 (N_18363,N_18108,N_18236);
xor U18364 (N_18364,N_18147,N_18193);
xor U18365 (N_18365,N_18198,N_18228);
nor U18366 (N_18366,N_18184,N_18174);
and U18367 (N_18367,N_18019,N_18169);
nand U18368 (N_18368,N_18029,N_18129);
xnor U18369 (N_18369,N_18208,N_18204);
nor U18370 (N_18370,N_18079,N_18137);
and U18371 (N_18371,N_18123,N_18039);
nor U18372 (N_18372,N_18244,N_18163);
or U18373 (N_18373,N_18044,N_18139);
or U18374 (N_18374,N_18104,N_18175);
or U18375 (N_18375,N_18247,N_18190);
nand U18376 (N_18376,N_18030,N_18120);
xnor U18377 (N_18377,N_18020,N_18027);
xnor U18378 (N_18378,N_18129,N_18229);
or U18379 (N_18379,N_18168,N_18169);
and U18380 (N_18380,N_18044,N_18209);
xor U18381 (N_18381,N_18221,N_18112);
nor U18382 (N_18382,N_18215,N_18109);
nand U18383 (N_18383,N_18179,N_18248);
or U18384 (N_18384,N_18227,N_18230);
nand U18385 (N_18385,N_18213,N_18235);
nor U18386 (N_18386,N_18096,N_18195);
nand U18387 (N_18387,N_18197,N_18225);
xnor U18388 (N_18388,N_18126,N_18221);
nor U18389 (N_18389,N_18066,N_18236);
or U18390 (N_18390,N_18000,N_18132);
nor U18391 (N_18391,N_18076,N_18029);
nor U18392 (N_18392,N_18189,N_18244);
nand U18393 (N_18393,N_18179,N_18132);
and U18394 (N_18394,N_18043,N_18154);
and U18395 (N_18395,N_18158,N_18102);
nand U18396 (N_18396,N_18020,N_18158);
and U18397 (N_18397,N_18056,N_18090);
and U18398 (N_18398,N_18066,N_18100);
or U18399 (N_18399,N_18039,N_18240);
or U18400 (N_18400,N_18003,N_18223);
or U18401 (N_18401,N_18156,N_18189);
and U18402 (N_18402,N_18125,N_18083);
nand U18403 (N_18403,N_18193,N_18125);
xnor U18404 (N_18404,N_18249,N_18027);
nand U18405 (N_18405,N_18138,N_18135);
and U18406 (N_18406,N_18193,N_18223);
xor U18407 (N_18407,N_18025,N_18238);
or U18408 (N_18408,N_18010,N_18134);
nor U18409 (N_18409,N_18109,N_18088);
xnor U18410 (N_18410,N_18228,N_18142);
or U18411 (N_18411,N_18081,N_18077);
nor U18412 (N_18412,N_18195,N_18065);
nor U18413 (N_18413,N_18023,N_18199);
nand U18414 (N_18414,N_18114,N_18007);
or U18415 (N_18415,N_18130,N_18033);
or U18416 (N_18416,N_18118,N_18194);
xor U18417 (N_18417,N_18169,N_18186);
or U18418 (N_18418,N_18207,N_18099);
nand U18419 (N_18419,N_18247,N_18032);
or U18420 (N_18420,N_18109,N_18122);
nand U18421 (N_18421,N_18033,N_18155);
and U18422 (N_18422,N_18092,N_18074);
nor U18423 (N_18423,N_18071,N_18229);
nor U18424 (N_18424,N_18193,N_18124);
xor U18425 (N_18425,N_18021,N_18249);
nand U18426 (N_18426,N_18040,N_18241);
xnor U18427 (N_18427,N_18051,N_18101);
nor U18428 (N_18428,N_18128,N_18159);
and U18429 (N_18429,N_18184,N_18005);
or U18430 (N_18430,N_18209,N_18061);
nand U18431 (N_18431,N_18079,N_18089);
xor U18432 (N_18432,N_18110,N_18031);
or U18433 (N_18433,N_18207,N_18242);
or U18434 (N_18434,N_18218,N_18129);
and U18435 (N_18435,N_18172,N_18110);
nand U18436 (N_18436,N_18072,N_18048);
nand U18437 (N_18437,N_18011,N_18240);
nand U18438 (N_18438,N_18153,N_18170);
nor U18439 (N_18439,N_18004,N_18154);
and U18440 (N_18440,N_18249,N_18204);
or U18441 (N_18441,N_18227,N_18062);
and U18442 (N_18442,N_18131,N_18152);
nand U18443 (N_18443,N_18044,N_18039);
or U18444 (N_18444,N_18196,N_18026);
or U18445 (N_18445,N_18111,N_18185);
nor U18446 (N_18446,N_18012,N_18185);
xor U18447 (N_18447,N_18105,N_18028);
nor U18448 (N_18448,N_18060,N_18122);
or U18449 (N_18449,N_18124,N_18089);
xnor U18450 (N_18450,N_18098,N_18085);
nand U18451 (N_18451,N_18120,N_18160);
and U18452 (N_18452,N_18066,N_18109);
nand U18453 (N_18453,N_18236,N_18150);
or U18454 (N_18454,N_18105,N_18222);
nor U18455 (N_18455,N_18011,N_18010);
xor U18456 (N_18456,N_18149,N_18076);
and U18457 (N_18457,N_18158,N_18038);
nor U18458 (N_18458,N_18129,N_18130);
nand U18459 (N_18459,N_18009,N_18023);
and U18460 (N_18460,N_18193,N_18120);
or U18461 (N_18461,N_18060,N_18226);
xnor U18462 (N_18462,N_18171,N_18000);
nor U18463 (N_18463,N_18042,N_18149);
xnor U18464 (N_18464,N_18129,N_18233);
or U18465 (N_18465,N_18191,N_18230);
xor U18466 (N_18466,N_18146,N_18015);
nor U18467 (N_18467,N_18238,N_18012);
xor U18468 (N_18468,N_18107,N_18100);
xnor U18469 (N_18469,N_18086,N_18143);
xnor U18470 (N_18470,N_18141,N_18244);
nand U18471 (N_18471,N_18235,N_18013);
nor U18472 (N_18472,N_18020,N_18090);
or U18473 (N_18473,N_18089,N_18114);
and U18474 (N_18474,N_18140,N_18056);
nand U18475 (N_18475,N_18236,N_18095);
xor U18476 (N_18476,N_18191,N_18056);
nor U18477 (N_18477,N_18180,N_18136);
xnor U18478 (N_18478,N_18097,N_18031);
xor U18479 (N_18479,N_18235,N_18214);
nand U18480 (N_18480,N_18202,N_18090);
and U18481 (N_18481,N_18217,N_18215);
or U18482 (N_18482,N_18150,N_18081);
or U18483 (N_18483,N_18040,N_18085);
xnor U18484 (N_18484,N_18087,N_18014);
nand U18485 (N_18485,N_18239,N_18243);
nand U18486 (N_18486,N_18037,N_18108);
nor U18487 (N_18487,N_18075,N_18200);
and U18488 (N_18488,N_18073,N_18135);
xor U18489 (N_18489,N_18064,N_18171);
nor U18490 (N_18490,N_18181,N_18195);
nand U18491 (N_18491,N_18056,N_18100);
nand U18492 (N_18492,N_18027,N_18214);
nand U18493 (N_18493,N_18122,N_18081);
nor U18494 (N_18494,N_18069,N_18184);
nand U18495 (N_18495,N_18000,N_18223);
nand U18496 (N_18496,N_18034,N_18222);
and U18497 (N_18497,N_18219,N_18217);
and U18498 (N_18498,N_18130,N_18225);
or U18499 (N_18499,N_18079,N_18225);
and U18500 (N_18500,N_18437,N_18399);
or U18501 (N_18501,N_18270,N_18291);
nand U18502 (N_18502,N_18441,N_18366);
xor U18503 (N_18503,N_18489,N_18252);
nor U18504 (N_18504,N_18496,N_18331);
xnor U18505 (N_18505,N_18316,N_18384);
xnor U18506 (N_18506,N_18268,N_18376);
nor U18507 (N_18507,N_18417,N_18289);
or U18508 (N_18508,N_18320,N_18344);
nor U18509 (N_18509,N_18345,N_18348);
and U18510 (N_18510,N_18303,N_18492);
nand U18511 (N_18511,N_18449,N_18335);
and U18512 (N_18512,N_18420,N_18283);
nand U18513 (N_18513,N_18455,N_18482);
nor U18514 (N_18514,N_18256,N_18319);
nand U18515 (N_18515,N_18394,N_18397);
and U18516 (N_18516,N_18300,N_18360);
xnor U18517 (N_18517,N_18263,N_18462);
nand U18518 (N_18518,N_18266,N_18454);
nand U18519 (N_18519,N_18448,N_18471);
xor U18520 (N_18520,N_18307,N_18429);
nor U18521 (N_18521,N_18431,N_18378);
and U18522 (N_18522,N_18313,N_18416);
and U18523 (N_18523,N_18410,N_18355);
or U18524 (N_18524,N_18330,N_18432);
or U18525 (N_18525,N_18272,N_18282);
and U18526 (N_18526,N_18324,N_18364);
nand U18527 (N_18527,N_18499,N_18293);
xnor U18528 (N_18528,N_18327,N_18259);
nand U18529 (N_18529,N_18288,N_18491);
and U18530 (N_18530,N_18265,N_18373);
or U18531 (N_18531,N_18301,N_18434);
nand U18532 (N_18532,N_18474,N_18447);
or U18533 (N_18533,N_18356,N_18445);
nor U18534 (N_18534,N_18306,N_18275);
nand U18535 (N_18535,N_18285,N_18343);
nand U18536 (N_18536,N_18284,N_18273);
or U18537 (N_18537,N_18359,N_18374);
nand U18538 (N_18538,N_18279,N_18483);
xnor U18539 (N_18539,N_18261,N_18281);
or U18540 (N_18540,N_18457,N_18446);
xnor U18541 (N_18541,N_18458,N_18372);
xor U18542 (N_18542,N_18310,N_18287);
nand U18543 (N_18543,N_18329,N_18338);
nor U18544 (N_18544,N_18456,N_18383);
xnor U18545 (N_18545,N_18251,N_18321);
xor U18546 (N_18546,N_18426,N_18428);
nand U18547 (N_18547,N_18309,N_18361);
nand U18548 (N_18548,N_18485,N_18297);
nand U18549 (N_18549,N_18299,N_18495);
nor U18550 (N_18550,N_18402,N_18476);
nand U18551 (N_18551,N_18332,N_18400);
or U18552 (N_18552,N_18341,N_18296);
or U18553 (N_18553,N_18258,N_18371);
and U18554 (N_18554,N_18409,N_18422);
nor U18555 (N_18555,N_18326,N_18484);
xnor U18556 (N_18556,N_18468,N_18322);
nand U18557 (N_18557,N_18470,N_18488);
nor U18558 (N_18558,N_18487,N_18421);
nor U18559 (N_18559,N_18401,N_18435);
xnor U18560 (N_18560,N_18405,N_18423);
nor U18561 (N_18561,N_18369,N_18486);
nand U18562 (N_18562,N_18377,N_18357);
and U18563 (N_18563,N_18392,N_18302);
xor U18564 (N_18564,N_18419,N_18413);
nor U18565 (N_18565,N_18398,N_18418);
and U18566 (N_18566,N_18480,N_18467);
and U18567 (N_18567,N_18430,N_18255);
nand U18568 (N_18568,N_18336,N_18305);
nand U18569 (N_18569,N_18267,N_18498);
or U18570 (N_18570,N_18466,N_18439);
nand U18571 (N_18571,N_18393,N_18494);
xor U18572 (N_18572,N_18271,N_18342);
xnor U18573 (N_18573,N_18365,N_18478);
nor U18574 (N_18574,N_18274,N_18325);
nand U18575 (N_18575,N_18396,N_18451);
nor U18576 (N_18576,N_18286,N_18481);
nor U18577 (N_18577,N_18280,N_18452);
or U18578 (N_18578,N_18334,N_18351);
and U18579 (N_18579,N_18388,N_18386);
or U18580 (N_18580,N_18442,N_18278);
xor U18581 (N_18581,N_18407,N_18403);
nand U18582 (N_18582,N_18349,N_18363);
and U18583 (N_18583,N_18312,N_18277);
or U18584 (N_18584,N_18262,N_18444);
or U18585 (N_18585,N_18264,N_18414);
nor U18586 (N_18586,N_18391,N_18412);
nand U18587 (N_18587,N_18254,N_18440);
nand U18588 (N_18588,N_18380,N_18362);
or U18589 (N_18589,N_18333,N_18269);
or U18590 (N_18590,N_18415,N_18315);
or U18591 (N_18591,N_18337,N_18339);
and U18592 (N_18592,N_18276,N_18425);
nor U18593 (N_18593,N_18385,N_18472);
nand U18594 (N_18594,N_18475,N_18260);
or U18595 (N_18595,N_18479,N_18461);
or U18596 (N_18596,N_18370,N_18382);
xnor U18597 (N_18597,N_18469,N_18453);
or U18598 (N_18598,N_18477,N_18443);
nand U18599 (N_18599,N_18350,N_18404);
and U18600 (N_18600,N_18408,N_18358);
xnor U18601 (N_18601,N_18395,N_18389);
nand U18602 (N_18602,N_18311,N_18367);
or U18603 (N_18603,N_18438,N_18381);
or U18604 (N_18604,N_18298,N_18294);
xnor U18605 (N_18605,N_18353,N_18314);
nor U18606 (N_18606,N_18424,N_18368);
and U18607 (N_18607,N_18292,N_18295);
xor U18608 (N_18608,N_18465,N_18406);
nand U18609 (N_18609,N_18493,N_18411);
and U18610 (N_18610,N_18346,N_18490);
nand U18611 (N_18611,N_18257,N_18463);
or U18612 (N_18612,N_18497,N_18328);
and U18613 (N_18613,N_18340,N_18387);
or U18614 (N_18614,N_18379,N_18318);
nand U18615 (N_18615,N_18459,N_18304);
and U18616 (N_18616,N_18473,N_18354);
and U18617 (N_18617,N_18427,N_18375);
or U18618 (N_18618,N_18250,N_18460);
or U18619 (N_18619,N_18317,N_18347);
nand U18620 (N_18620,N_18450,N_18433);
nand U18621 (N_18621,N_18308,N_18436);
nor U18622 (N_18622,N_18253,N_18323);
or U18623 (N_18623,N_18290,N_18352);
and U18624 (N_18624,N_18390,N_18464);
nor U18625 (N_18625,N_18490,N_18336);
or U18626 (N_18626,N_18448,N_18470);
nand U18627 (N_18627,N_18311,N_18424);
nor U18628 (N_18628,N_18379,N_18380);
xor U18629 (N_18629,N_18280,N_18453);
nor U18630 (N_18630,N_18397,N_18283);
nor U18631 (N_18631,N_18368,N_18340);
nor U18632 (N_18632,N_18274,N_18470);
and U18633 (N_18633,N_18443,N_18468);
nor U18634 (N_18634,N_18438,N_18370);
or U18635 (N_18635,N_18296,N_18340);
nor U18636 (N_18636,N_18283,N_18321);
nand U18637 (N_18637,N_18354,N_18391);
xor U18638 (N_18638,N_18485,N_18338);
xnor U18639 (N_18639,N_18357,N_18385);
or U18640 (N_18640,N_18438,N_18424);
nor U18641 (N_18641,N_18439,N_18487);
and U18642 (N_18642,N_18416,N_18294);
xnor U18643 (N_18643,N_18282,N_18341);
xnor U18644 (N_18644,N_18381,N_18267);
xnor U18645 (N_18645,N_18353,N_18490);
xnor U18646 (N_18646,N_18268,N_18296);
xor U18647 (N_18647,N_18494,N_18360);
nand U18648 (N_18648,N_18416,N_18316);
xnor U18649 (N_18649,N_18487,N_18405);
xor U18650 (N_18650,N_18272,N_18425);
nor U18651 (N_18651,N_18461,N_18415);
nor U18652 (N_18652,N_18454,N_18411);
or U18653 (N_18653,N_18450,N_18352);
or U18654 (N_18654,N_18420,N_18303);
and U18655 (N_18655,N_18317,N_18480);
and U18656 (N_18656,N_18313,N_18308);
xor U18657 (N_18657,N_18458,N_18266);
nor U18658 (N_18658,N_18295,N_18345);
or U18659 (N_18659,N_18250,N_18428);
nor U18660 (N_18660,N_18278,N_18410);
xor U18661 (N_18661,N_18347,N_18416);
and U18662 (N_18662,N_18292,N_18268);
and U18663 (N_18663,N_18343,N_18258);
or U18664 (N_18664,N_18371,N_18323);
nor U18665 (N_18665,N_18391,N_18326);
or U18666 (N_18666,N_18340,N_18409);
and U18667 (N_18667,N_18304,N_18265);
or U18668 (N_18668,N_18471,N_18459);
nand U18669 (N_18669,N_18356,N_18348);
and U18670 (N_18670,N_18307,N_18337);
or U18671 (N_18671,N_18438,N_18290);
or U18672 (N_18672,N_18371,N_18384);
xnor U18673 (N_18673,N_18331,N_18281);
nand U18674 (N_18674,N_18322,N_18460);
nor U18675 (N_18675,N_18438,N_18295);
or U18676 (N_18676,N_18346,N_18426);
and U18677 (N_18677,N_18372,N_18274);
and U18678 (N_18678,N_18402,N_18260);
and U18679 (N_18679,N_18366,N_18393);
or U18680 (N_18680,N_18318,N_18469);
or U18681 (N_18681,N_18397,N_18476);
and U18682 (N_18682,N_18409,N_18452);
or U18683 (N_18683,N_18429,N_18499);
xor U18684 (N_18684,N_18431,N_18299);
and U18685 (N_18685,N_18364,N_18263);
xnor U18686 (N_18686,N_18313,N_18492);
and U18687 (N_18687,N_18363,N_18366);
xor U18688 (N_18688,N_18484,N_18366);
nand U18689 (N_18689,N_18408,N_18417);
nor U18690 (N_18690,N_18286,N_18322);
or U18691 (N_18691,N_18263,N_18283);
xnor U18692 (N_18692,N_18349,N_18458);
nand U18693 (N_18693,N_18386,N_18404);
xnor U18694 (N_18694,N_18447,N_18440);
nand U18695 (N_18695,N_18258,N_18470);
xor U18696 (N_18696,N_18361,N_18459);
nor U18697 (N_18697,N_18413,N_18270);
nand U18698 (N_18698,N_18397,N_18441);
and U18699 (N_18699,N_18491,N_18303);
nor U18700 (N_18700,N_18499,N_18355);
nand U18701 (N_18701,N_18318,N_18269);
or U18702 (N_18702,N_18486,N_18378);
or U18703 (N_18703,N_18412,N_18320);
or U18704 (N_18704,N_18398,N_18286);
and U18705 (N_18705,N_18494,N_18297);
or U18706 (N_18706,N_18494,N_18309);
nor U18707 (N_18707,N_18387,N_18439);
or U18708 (N_18708,N_18332,N_18410);
nor U18709 (N_18709,N_18337,N_18376);
and U18710 (N_18710,N_18338,N_18408);
nor U18711 (N_18711,N_18287,N_18395);
nand U18712 (N_18712,N_18483,N_18471);
nor U18713 (N_18713,N_18417,N_18372);
and U18714 (N_18714,N_18275,N_18469);
xor U18715 (N_18715,N_18491,N_18329);
nor U18716 (N_18716,N_18313,N_18334);
and U18717 (N_18717,N_18442,N_18401);
or U18718 (N_18718,N_18450,N_18364);
nor U18719 (N_18719,N_18336,N_18355);
xor U18720 (N_18720,N_18445,N_18289);
xor U18721 (N_18721,N_18368,N_18377);
nor U18722 (N_18722,N_18341,N_18316);
and U18723 (N_18723,N_18275,N_18355);
nand U18724 (N_18724,N_18400,N_18410);
or U18725 (N_18725,N_18388,N_18307);
or U18726 (N_18726,N_18254,N_18401);
nor U18727 (N_18727,N_18395,N_18478);
or U18728 (N_18728,N_18430,N_18319);
and U18729 (N_18729,N_18392,N_18425);
nand U18730 (N_18730,N_18410,N_18474);
and U18731 (N_18731,N_18476,N_18257);
or U18732 (N_18732,N_18266,N_18408);
xor U18733 (N_18733,N_18316,N_18379);
nand U18734 (N_18734,N_18427,N_18267);
or U18735 (N_18735,N_18323,N_18252);
nor U18736 (N_18736,N_18408,N_18488);
nand U18737 (N_18737,N_18384,N_18349);
nand U18738 (N_18738,N_18431,N_18309);
and U18739 (N_18739,N_18343,N_18378);
nor U18740 (N_18740,N_18339,N_18284);
nor U18741 (N_18741,N_18419,N_18485);
xnor U18742 (N_18742,N_18483,N_18423);
or U18743 (N_18743,N_18494,N_18430);
and U18744 (N_18744,N_18260,N_18399);
or U18745 (N_18745,N_18415,N_18422);
and U18746 (N_18746,N_18429,N_18392);
xor U18747 (N_18747,N_18440,N_18328);
nand U18748 (N_18748,N_18269,N_18284);
xor U18749 (N_18749,N_18299,N_18324);
or U18750 (N_18750,N_18563,N_18610);
nand U18751 (N_18751,N_18598,N_18537);
xnor U18752 (N_18752,N_18680,N_18597);
or U18753 (N_18753,N_18615,N_18717);
and U18754 (N_18754,N_18518,N_18504);
xnor U18755 (N_18755,N_18629,N_18679);
nand U18756 (N_18756,N_18650,N_18628);
nor U18757 (N_18757,N_18574,N_18667);
xor U18758 (N_18758,N_18626,N_18612);
and U18759 (N_18759,N_18607,N_18665);
and U18760 (N_18760,N_18546,N_18586);
and U18761 (N_18761,N_18535,N_18543);
nand U18762 (N_18762,N_18689,N_18572);
and U18763 (N_18763,N_18560,N_18506);
xor U18764 (N_18764,N_18538,N_18643);
or U18765 (N_18765,N_18663,N_18625);
nand U18766 (N_18766,N_18729,N_18556);
or U18767 (N_18767,N_18647,N_18743);
and U18768 (N_18768,N_18609,N_18671);
nor U18769 (N_18769,N_18527,N_18631);
nand U18770 (N_18770,N_18737,N_18588);
nand U18771 (N_18771,N_18664,N_18508);
nand U18772 (N_18772,N_18744,N_18569);
xor U18773 (N_18773,N_18548,N_18520);
or U18774 (N_18774,N_18703,N_18713);
and U18775 (N_18775,N_18693,N_18608);
xnor U18776 (N_18776,N_18551,N_18748);
or U18777 (N_18777,N_18512,N_18723);
or U18778 (N_18778,N_18639,N_18677);
nor U18779 (N_18779,N_18571,N_18613);
and U18780 (N_18780,N_18515,N_18657);
nand U18781 (N_18781,N_18594,N_18674);
xnor U18782 (N_18782,N_18519,N_18620);
xor U18783 (N_18783,N_18542,N_18500);
xnor U18784 (N_18784,N_18524,N_18636);
or U18785 (N_18785,N_18682,N_18559);
and U18786 (N_18786,N_18721,N_18553);
xnor U18787 (N_18787,N_18694,N_18521);
nor U18788 (N_18788,N_18741,N_18529);
or U18789 (N_18789,N_18644,N_18545);
and U18790 (N_18790,N_18745,N_18525);
xor U18791 (N_18791,N_18509,N_18699);
or U18792 (N_18792,N_18728,N_18532);
or U18793 (N_18793,N_18573,N_18730);
nand U18794 (N_18794,N_18541,N_18530);
or U18795 (N_18795,N_18687,N_18704);
and U18796 (N_18796,N_18513,N_18738);
nor U18797 (N_18797,N_18549,N_18690);
xor U18798 (N_18798,N_18547,N_18675);
xnor U18799 (N_18799,N_18581,N_18627);
nor U18800 (N_18800,N_18742,N_18714);
xnor U18801 (N_18801,N_18708,N_18531);
nor U18802 (N_18802,N_18692,N_18749);
xor U18803 (N_18803,N_18660,N_18735);
nand U18804 (N_18804,N_18661,N_18698);
nand U18805 (N_18805,N_18645,N_18510);
and U18806 (N_18806,N_18584,N_18653);
xor U18807 (N_18807,N_18666,N_18640);
nand U18808 (N_18808,N_18570,N_18649);
nand U18809 (N_18809,N_18678,N_18722);
or U18810 (N_18810,N_18720,N_18684);
nor U18811 (N_18811,N_18599,N_18540);
or U18812 (N_18812,N_18668,N_18582);
and U18813 (N_18813,N_18691,N_18732);
or U18814 (N_18814,N_18706,N_18623);
or U18815 (N_18815,N_18596,N_18580);
and U18816 (N_18816,N_18575,N_18734);
or U18817 (N_18817,N_18651,N_18696);
and U18818 (N_18818,N_18616,N_18746);
and U18819 (N_18819,N_18711,N_18605);
nand U18820 (N_18820,N_18731,N_18705);
and U18821 (N_18821,N_18523,N_18576);
xor U18822 (N_18822,N_18554,N_18740);
and U18823 (N_18823,N_18635,N_18726);
or U18824 (N_18824,N_18659,N_18579);
or U18825 (N_18825,N_18614,N_18514);
nand U18826 (N_18826,N_18590,N_18564);
xnor U18827 (N_18827,N_18503,N_18733);
or U18828 (N_18828,N_18585,N_18592);
xnor U18829 (N_18829,N_18621,N_18526);
xor U18830 (N_18830,N_18522,N_18646);
nand U18831 (N_18831,N_18648,N_18658);
nor U18832 (N_18832,N_18709,N_18539);
nor U18833 (N_18833,N_18662,N_18568);
nor U18834 (N_18834,N_18550,N_18565);
and U18835 (N_18835,N_18724,N_18669);
and U18836 (N_18836,N_18715,N_18618);
or U18837 (N_18837,N_18683,N_18686);
and U18838 (N_18838,N_18566,N_18601);
nor U18839 (N_18839,N_18511,N_18600);
and U18840 (N_18840,N_18656,N_18534);
nor U18841 (N_18841,N_18707,N_18517);
xnor U18842 (N_18842,N_18611,N_18670);
and U18843 (N_18843,N_18558,N_18700);
and U18844 (N_18844,N_18603,N_18617);
xor U18845 (N_18845,N_18697,N_18633);
nor U18846 (N_18846,N_18727,N_18712);
xor U18847 (N_18847,N_18604,N_18606);
nor U18848 (N_18848,N_18501,N_18718);
nand U18849 (N_18849,N_18739,N_18681);
nor U18850 (N_18850,N_18638,N_18637);
or U18851 (N_18851,N_18719,N_18641);
xnor U18852 (N_18852,N_18747,N_18630);
and U18853 (N_18853,N_18577,N_18642);
xor U18854 (N_18854,N_18716,N_18516);
nor U18855 (N_18855,N_18655,N_18676);
nor U18856 (N_18856,N_18502,N_18634);
nor U18857 (N_18857,N_18622,N_18505);
xnor U18858 (N_18858,N_18528,N_18533);
nor U18859 (N_18859,N_18552,N_18725);
or U18860 (N_18860,N_18702,N_18544);
xnor U18861 (N_18861,N_18578,N_18652);
and U18862 (N_18862,N_18619,N_18561);
xor U18863 (N_18863,N_18562,N_18602);
nor U18864 (N_18864,N_18688,N_18673);
nand U18865 (N_18865,N_18672,N_18567);
nand U18866 (N_18866,N_18654,N_18555);
nand U18867 (N_18867,N_18593,N_18685);
or U18868 (N_18868,N_18589,N_18632);
nor U18869 (N_18869,N_18701,N_18591);
nand U18870 (N_18870,N_18557,N_18507);
or U18871 (N_18871,N_18710,N_18624);
xor U18872 (N_18872,N_18587,N_18536);
nand U18873 (N_18873,N_18736,N_18695);
nor U18874 (N_18874,N_18583,N_18595);
xnor U18875 (N_18875,N_18734,N_18678);
xor U18876 (N_18876,N_18604,N_18724);
xnor U18877 (N_18877,N_18582,N_18503);
nor U18878 (N_18878,N_18605,N_18633);
nor U18879 (N_18879,N_18703,N_18581);
or U18880 (N_18880,N_18732,N_18718);
nand U18881 (N_18881,N_18646,N_18713);
nand U18882 (N_18882,N_18582,N_18639);
nor U18883 (N_18883,N_18597,N_18664);
xor U18884 (N_18884,N_18544,N_18570);
nor U18885 (N_18885,N_18605,N_18710);
or U18886 (N_18886,N_18594,N_18565);
nand U18887 (N_18887,N_18570,N_18533);
and U18888 (N_18888,N_18515,N_18610);
xnor U18889 (N_18889,N_18545,N_18543);
and U18890 (N_18890,N_18574,N_18625);
nand U18891 (N_18891,N_18652,N_18587);
xnor U18892 (N_18892,N_18722,N_18614);
or U18893 (N_18893,N_18671,N_18725);
or U18894 (N_18894,N_18729,N_18547);
nand U18895 (N_18895,N_18635,N_18748);
nor U18896 (N_18896,N_18658,N_18569);
nor U18897 (N_18897,N_18567,N_18516);
nor U18898 (N_18898,N_18615,N_18696);
nor U18899 (N_18899,N_18621,N_18636);
xnor U18900 (N_18900,N_18527,N_18546);
nor U18901 (N_18901,N_18640,N_18627);
or U18902 (N_18902,N_18708,N_18578);
nand U18903 (N_18903,N_18714,N_18740);
or U18904 (N_18904,N_18731,N_18566);
nand U18905 (N_18905,N_18600,N_18618);
nor U18906 (N_18906,N_18634,N_18705);
xor U18907 (N_18907,N_18747,N_18618);
or U18908 (N_18908,N_18746,N_18535);
nor U18909 (N_18909,N_18569,N_18574);
and U18910 (N_18910,N_18745,N_18697);
or U18911 (N_18911,N_18694,N_18565);
or U18912 (N_18912,N_18691,N_18671);
or U18913 (N_18913,N_18555,N_18582);
nand U18914 (N_18914,N_18610,N_18712);
nand U18915 (N_18915,N_18577,N_18630);
or U18916 (N_18916,N_18671,N_18628);
and U18917 (N_18917,N_18645,N_18562);
or U18918 (N_18918,N_18607,N_18731);
nor U18919 (N_18919,N_18505,N_18529);
and U18920 (N_18920,N_18516,N_18607);
or U18921 (N_18921,N_18676,N_18648);
nand U18922 (N_18922,N_18601,N_18744);
and U18923 (N_18923,N_18676,N_18689);
xnor U18924 (N_18924,N_18672,N_18594);
and U18925 (N_18925,N_18509,N_18506);
nor U18926 (N_18926,N_18670,N_18537);
nand U18927 (N_18927,N_18659,N_18596);
nor U18928 (N_18928,N_18705,N_18649);
nor U18929 (N_18929,N_18563,N_18746);
or U18930 (N_18930,N_18731,N_18662);
nand U18931 (N_18931,N_18524,N_18634);
and U18932 (N_18932,N_18573,N_18681);
xnor U18933 (N_18933,N_18736,N_18538);
and U18934 (N_18934,N_18539,N_18694);
nor U18935 (N_18935,N_18742,N_18568);
nor U18936 (N_18936,N_18586,N_18674);
nor U18937 (N_18937,N_18686,N_18574);
or U18938 (N_18938,N_18614,N_18730);
nand U18939 (N_18939,N_18533,N_18507);
or U18940 (N_18940,N_18593,N_18545);
or U18941 (N_18941,N_18661,N_18738);
xnor U18942 (N_18942,N_18617,N_18646);
nand U18943 (N_18943,N_18641,N_18683);
nor U18944 (N_18944,N_18651,N_18715);
nor U18945 (N_18945,N_18561,N_18610);
or U18946 (N_18946,N_18510,N_18501);
and U18947 (N_18947,N_18564,N_18708);
or U18948 (N_18948,N_18681,N_18517);
and U18949 (N_18949,N_18510,N_18686);
xnor U18950 (N_18950,N_18599,N_18533);
nand U18951 (N_18951,N_18622,N_18543);
and U18952 (N_18952,N_18615,N_18513);
and U18953 (N_18953,N_18585,N_18623);
nand U18954 (N_18954,N_18624,N_18617);
or U18955 (N_18955,N_18721,N_18580);
and U18956 (N_18956,N_18556,N_18515);
and U18957 (N_18957,N_18508,N_18639);
nand U18958 (N_18958,N_18535,N_18613);
and U18959 (N_18959,N_18566,N_18578);
or U18960 (N_18960,N_18700,N_18512);
or U18961 (N_18961,N_18571,N_18508);
nor U18962 (N_18962,N_18625,N_18746);
xor U18963 (N_18963,N_18631,N_18570);
nor U18964 (N_18964,N_18666,N_18620);
nand U18965 (N_18965,N_18519,N_18586);
nor U18966 (N_18966,N_18724,N_18657);
or U18967 (N_18967,N_18542,N_18539);
or U18968 (N_18968,N_18664,N_18707);
xnor U18969 (N_18969,N_18604,N_18664);
nand U18970 (N_18970,N_18691,N_18543);
or U18971 (N_18971,N_18540,N_18596);
nor U18972 (N_18972,N_18647,N_18734);
and U18973 (N_18973,N_18667,N_18542);
nand U18974 (N_18974,N_18504,N_18717);
nand U18975 (N_18975,N_18502,N_18505);
nor U18976 (N_18976,N_18570,N_18663);
nor U18977 (N_18977,N_18706,N_18524);
xor U18978 (N_18978,N_18548,N_18721);
xnor U18979 (N_18979,N_18506,N_18646);
xor U18980 (N_18980,N_18609,N_18640);
nor U18981 (N_18981,N_18695,N_18526);
nand U18982 (N_18982,N_18622,N_18581);
xor U18983 (N_18983,N_18578,N_18670);
or U18984 (N_18984,N_18648,N_18594);
nor U18985 (N_18985,N_18592,N_18707);
xnor U18986 (N_18986,N_18565,N_18679);
xnor U18987 (N_18987,N_18653,N_18585);
and U18988 (N_18988,N_18652,N_18616);
nand U18989 (N_18989,N_18711,N_18651);
nand U18990 (N_18990,N_18555,N_18580);
or U18991 (N_18991,N_18510,N_18657);
nor U18992 (N_18992,N_18736,N_18663);
nand U18993 (N_18993,N_18529,N_18600);
nor U18994 (N_18994,N_18662,N_18623);
and U18995 (N_18995,N_18538,N_18580);
xor U18996 (N_18996,N_18630,N_18641);
xnor U18997 (N_18997,N_18698,N_18687);
xnor U18998 (N_18998,N_18577,N_18511);
xnor U18999 (N_18999,N_18685,N_18709);
nand U19000 (N_19000,N_18944,N_18770);
xnor U19001 (N_19001,N_18791,N_18925);
nor U19002 (N_19002,N_18974,N_18834);
xnor U19003 (N_19003,N_18750,N_18863);
xor U19004 (N_19004,N_18828,N_18924);
or U19005 (N_19005,N_18775,N_18996);
nand U19006 (N_19006,N_18890,N_18782);
xnor U19007 (N_19007,N_18803,N_18835);
nand U19008 (N_19008,N_18966,N_18855);
nor U19009 (N_19009,N_18839,N_18850);
xor U19010 (N_19010,N_18942,N_18883);
nand U19011 (N_19011,N_18956,N_18906);
nor U19012 (N_19012,N_18773,N_18967);
or U19013 (N_19013,N_18948,N_18777);
and U19014 (N_19014,N_18827,N_18756);
and U19015 (N_19015,N_18911,N_18814);
nor U19016 (N_19016,N_18951,N_18862);
nor U19017 (N_19017,N_18846,N_18832);
and U19018 (N_19018,N_18810,N_18926);
xor U19019 (N_19019,N_18845,N_18757);
nand U19020 (N_19020,N_18772,N_18927);
nor U19021 (N_19021,N_18954,N_18792);
xor U19022 (N_19022,N_18797,N_18997);
nand U19023 (N_19023,N_18935,N_18795);
xor U19024 (N_19024,N_18752,N_18811);
or U19025 (N_19025,N_18858,N_18889);
and U19026 (N_19026,N_18960,N_18824);
nand U19027 (N_19027,N_18872,N_18887);
nand U19028 (N_19028,N_18952,N_18866);
xnor U19029 (N_19029,N_18784,N_18842);
nand U19030 (N_19030,N_18976,N_18809);
or U19031 (N_19031,N_18953,N_18776);
nor U19032 (N_19032,N_18787,N_18841);
nor U19033 (N_19033,N_18760,N_18875);
and U19034 (N_19034,N_18922,N_18965);
nor U19035 (N_19035,N_18767,N_18980);
xor U19036 (N_19036,N_18892,N_18915);
or U19037 (N_19037,N_18794,N_18812);
and U19038 (N_19038,N_18946,N_18877);
nand U19039 (N_19039,N_18920,N_18985);
xnor U19040 (N_19040,N_18848,N_18938);
nand U19041 (N_19041,N_18964,N_18999);
or U19042 (N_19042,N_18774,N_18755);
nor U19043 (N_19043,N_18816,N_18878);
xor U19044 (N_19044,N_18901,N_18837);
nor U19045 (N_19045,N_18753,N_18793);
xor U19046 (N_19046,N_18916,N_18761);
and U19047 (N_19047,N_18765,N_18836);
xnor U19048 (N_19048,N_18886,N_18778);
or U19049 (N_19049,N_18898,N_18766);
xnor U19050 (N_19050,N_18940,N_18936);
nand U19051 (N_19051,N_18779,N_18959);
xnor U19052 (N_19052,N_18994,N_18785);
nor U19053 (N_19053,N_18970,N_18847);
nand U19054 (N_19054,N_18822,N_18993);
or U19055 (N_19055,N_18808,N_18815);
nand U19056 (N_19056,N_18977,N_18879);
or U19057 (N_19057,N_18800,N_18790);
and U19058 (N_19058,N_18860,N_18813);
nor U19059 (N_19059,N_18851,N_18831);
nor U19060 (N_19060,N_18918,N_18806);
and U19061 (N_19061,N_18897,N_18998);
xor U19062 (N_19062,N_18789,N_18932);
xnor U19063 (N_19063,N_18856,N_18949);
xor U19064 (N_19064,N_18871,N_18868);
or U19065 (N_19065,N_18958,N_18941);
or U19066 (N_19066,N_18933,N_18764);
and U19067 (N_19067,N_18961,N_18909);
or U19068 (N_19068,N_18963,N_18874);
xnor U19069 (N_19069,N_18882,N_18881);
nand U19070 (N_19070,N_18904,N_18894);
or U19071 (N_19071,N_18931,N_18838);
or U19072 (N_19072,N_18913,N_18751);
nand U19073 (N_19073,N_18972,N_18989);
xor U19074 (N_19074,N_18759,N_18919);
or U19075 (N_19075,N_18857,N_18910);
and U19076 (N_19076,N_18947,N_18902);
or U19077 (N_19077,N_18992,N_18786);
or U19078 (N_19078,N_18939,N_18903);
and U19079 (N_19079,N_18950,N_18833);
nor U19080 (N_19080,N_18869,N_18973);
nand U19081 (N_19081,N_18807,N_18979);
xnor U19082 (N_19082,N_18804,N_18829);
or U19083 (N_19083,N_18771,N_18895);
or U19084 (N_19084,N_18955,N_18820);
nand U19085 (N_19085,N_18930,N_18984);
nand U19086 (N_19086,N_18943,N_18830);
and U19087 (N_19087,N_18991,N_18802);
nand U19088 (N_19088,N_18957,N_18962);
xnor U19089 (N_19089,N_18880,N_18884);
xor U19090 (N_19090,N_18891,N_18928);
and U19091 (N_19091,N_18818,N_18798);
nor U19092 (N_19092,N_18921,N_18817);
nor U19093 (N_19093,N_18995,N_18865);
nand U19094 (N_19094,N_18988,N_18893);
nand U19095 (N_19095,N_18796,N_18873);
nor U19096 (N_19096,N_18969,N_18826);
and U19097 (N_19097,N_18912,N_18754);
and U19098 (N_19098,N_18768,N_18870);
and U19099 (N_19099,N_18853,N_18885);
nand U19100 (N_19100,N_18934,N_18981);
xor U19101 (N_19101,N_18888,N_18914);
nor U19102 (N_19102,N_18843,N_18799);
and U19103 (N_19103,N_18900,N_18908);
xor U19104 (N_19104,N_18945,N_18876);
nand U19105 (N_19105,N_18840,N_18971);
nor U19106 (N_19106,N_18859,N_18864);
nand U19107 (N_19107,N_18896,N_18899);
xor U19108 (N_19108,N_18907,N_18975);
or U19109 (N_19109,N_18849,N_18937);
nand U19110 (N_19110,N_18780,N_18990);
nand U19111 (N_19111,N_18861,N_18923);
nor U19112 (N_19112,N_18781,N_18905);
xor U19113 (N_19113,N_18852,N_18823);
nor U19114 (N_19114,N_18982,N_18968);
nand U19115 (N_19115,N_18769,N_18983);
nor U19116 (N_19116,N_18801,N_18867);
xor U19117 (N_19117,N_18978,N_18929);
nor U19118 (N_19118,N_18986,N_18917);
xor U19119 (N_19119,N_18819,N_18821);
and U19120 (N_19120,N_18758,N_18783);
and U19121 (N_19121,N_18825,N_18762);
xor U19122 (N_19122,N_18987,N_18763);
xnor U19123 (N_19123,N_18788,N_18805);
xnor U19124 (N_19124,N_18854,N_18844);
or U19125 (N_19125,N_18782,N_18774);
and U19126 (N_19126,N_18814,N_18857);
xor U19127 (N_19127,N_18793,N_18774);
nor U19128 (N_19128,N_18833,N_18881);
xor U19129 (N_19129,N_18887,N_18979);
nand U19130 (N_19130,N_18951,N_18930);
xnor U19131 (N_19131,N_18926,N_18955);
or U19132 (N_19132,N_18898,N_18864);
or U19133 (N_19133,N_18807,N_18801);
and U19134 (N_19134,N_18971,N_18980);
and U19135 (N_19135,N_18989,N_18923);
xnor U19136 (N_19136,N_18965,N_18929);
or U19137 (N_19137,N_18947,N_18834);
nand U19138 (N_19138,N_18894,N_18907);
and U19139 (N_19139,N_18836,N_18938);
nor U19140 (N_19140,N_18806,N_18998);
nor U19141 (N_19141,N_18804,N_18992);
xnor U19142 (N_19142,N_18914,N_18870);
xnor U19143 (N_19143,N_18845,N_18965);
nor U19144 (N_19144,N_18967,N_18990);
nand U19145 (N_19145,N_18782,N_18771);
or U19146 (N_19146,N_18927,N_18785);
or U19147 (N_19147,N_18934,N_18942);
nor U19148 (N_19148,N_18906,N_18895);
xor U19149 (N_19149,N_18777,N_18873);
nor U19150 (N_19150,N_18961,N_18833);
or U19151 (N_19151,N_18915,N_18785);
xor U19152 (N_19152,N_18889,N_18941);
nor U19153 (N_19153,N_18847,N_18926);
nor U19154 (N_19154,N_18992,N_18919);
or U19155 (N_19155,N_18897,N_18770);
or U19156 (N_19156,N_18923,N_18849);
xnor U19157 (N_19157,N_18902,N_18805);
nand U19158 (N_19158,N_18999,N_18787);
nor U19159 (N_19159,N_18810,N_18767);
nor U19160 (N_19160,N_18935,N_18918);
nor U19161 (N_19161,N_18799,N_18906);
xor U19162 (N_19162,N_18764,N_18945);
nand U19163 (N_19163,N_18821,N_18779);
nor U19164 (N_19164,N_18938,N_18881);
and U19165 (N_19165,N_18841,N_18811);
xor U19166 (N_19166,N_18751,N_18966);
and U19167 (N_19167,N_18994,N_18959);
and U19168 (N_19168,N_18882,N_18964);
xnor U19169 (N_19169,N_18882,N_18993);
and U19170 (N_19170,N_18807,N_18793);
or U19171 (N_19171,N_18981,N_18855);
xnor U19172 (N_19172,N_18899,N_18942);
nand U19173 (N_19173,N_18829,N_18858);
and U19174 (N_19174,N_18970,N_18843);
nand U19175 (N_19175,N_18965,N_18761);
or U19176 (N_19176,N_18920,N_18885);
nor U19177 (N_19177,N_18907,N_18985);
or U19178 (N_19178,N_18790,N_18919);
and U19179 (N_19179,N_18796,N_18751);
or U19180 (N_19180,N_18991,N_18768);
or U19181 (N_19181,N_18890,N_18885);
and U19182 (N_19182,N_18976,N_18988);
and U19183 (N_19183,N_18789,N_18957);
xnor U19184 (N_19184,N_18985,N_18754);
nand U19185 (N_19185,N_18956,N_18970);
nor U19186 (N_19186,N_18758,N_18962);
nor U19187 (N_19187,N_18845,N_18952);
xor U19188 (N_19188,N_18786,N_18801);
nor U19189 (N_19189,N_18772,N_18919);
nand U19190 (N_19190,N_18928,N_18799);
and U19191 (N_19191,N_18835,N_18943);
nand U19192 (N_19192,N_18843,N_18992);
or U19193 (N_19193,N_18917,N_18981);
nor U19194 (N_19194,N_18771,N_18979);
nor U19195 (N_19195,N_18925,N_18866);
or U19196 (N_19196,N_18939,N_18839);
nor U19197 (N_19197,N_18895,N_18966);
xnor U19198 (N_19198,N_18957,N_18787);
or U19199 (N_19199,N_18796,N_18889);
nor U19200 (N_19200,N_18976,N_18909);
xor U19201 (N_19201,N_18843,N_18872);
or U19202 (N_19202,N_18904,N_18921);
or U19203 (N_19203,N_18758,N_18769);
nor U19204 (N_19204,N_18816,N_18776);
xor U19205 (N_19205,N_18944,N_18923);
or U19206 (N_19206,N_18883,N_18935);
or U19207 (N_19207,N_18833,N_18812);
nor U19208 (N_19208,N_18865,N_18834);
nor U19209 (N_19209,N_18773,N_18815);
xor U19210 (N_19210,N_18835,N_18815);
xor U19211 (N_19211,N_18760,N_18985);
nand U19212 (N_19212,N_18969,N_18959);
or U19213 (N_19213,N_18826,N_18810);
nor U19214 (N_19214,N_18837,N_18806);
nand U19215 (N_19215,N_18899,N_18928);
nand U19216 (N_19216,N_18788,N_18750);
xnor U19217 (N_19217,N_18986,N_18898);
or U19218 (N_19218,N_18780,N_18850);
xor U19219 (N_19219,N_18787,N_18946);
nor U19220 (N_19220,N_18776,N_18925);
nor U19221 (N_19221,N_18895,N_18931);
nor U19222 (N_19222,N_18842,N_18840);
nor U19223 (N_19223,N_18979,N_18791);
xnor U19224 (N_19224,N_18959,N_18967);
xnor U19225 (N_19225,N_18917,N_18755);
or U19226 (N_19226,N_18902,N_18807);
xnor U19227 (N_19227,N_18774,N_18960);
nand U19228 (N_19228,N_18805,N_18757);
nor U19229 (N_19229,N_18921,N_18863);
and U19230 (N_19230,N_18994,N_18853);
nor U19231 (N_19231,N_18779,N_18947);
or U19232 (N_19232,N_18957,N_18783);
and U19233 (N_19233,N_18971,N_18957);
and U19234 (N_19234,N_18779,N_18993);
xnor U19235 (N_19235,N_18848,N_18916);
and U19236 (N_19236,N_18879,N_18778);
and U19237 (N_19237,N_18818,N_18922);
nor U19238 (N_19238,N_18925,N_18977);
xor U19239 (N_19239,N_18896,N_18761);
and U19240 (N_19240,N_18920,N_18900);
nor U19241 (N_19241,N_18991,N_18995);
xor U19242 (N_19242,N_18831,N_18939);
nand U19243 (N_19243,N_18789,N_18912);
and U19244 (N_19244,N_18826,N_18984);
xnor U19245 (N_19245,N_18932,N_18800);
or U19246 (N_19246,N_18855,N_18791);
nand U19247 (N_19247,N_18993,N_18772);
xor U19248 (N_19248,N_18850,N_18978);
xor U19249 (N_19249,N_18859,N_18880);
or U19250 (N_19250,N_19049,N_19057);
or U19251 (N_19251,N_19224,N_19127);
xnor U19252 (N_19252,N_19037,N_19137);
or U19253 (N_19253,N_19084,N_19218);
nor U19254 (N_19254,N_19202,N_19028);
or U19255 (N_19255,N_19228,N_19227);
nor U19256 (N_19256,N_19158,N_19038);
and U19257 (N_19257,N_19087,N_19030);
xnor U19258 (N_19258,N_19237,N_19231);
and U19259 (N_19259,N_19021,N_19067);
xnor U19260 (N_19260,N_19174,N_19195);
nor U19261 (N_19261,N_19175,N_19076);
and U19262 (N_19262,N_19153,N_19016);
xnor U19263 (N_19263,N_19064,N_19181);
xnor U19264 (N_19264,N_19155,N_19099);
nor U19265 (N_19265,N_19140,N_19012);
or U19266 (N_19266,N_19185,N_19241);
or U19267 (N_19267,N_19098,N_19033);
and U19268 (N_19268,N_19234,N_19050);
or U19269 (N_19269,N_19133,N_19215);
and U19270 (N_19270,N_19168,N_19197);
or U19271 (N_19271,N_19122,N_19022);
nor U19272 (N_19272,N_19120,N_19062);
or U19273 (N_19273,N_19232,N_19123);
or U19274 (N_19274,N_19208,N_19249);
nor U19275 (N_19275,N_19220,N_19005);
nand U19276 (N_19276,N_19119,N_19248);
or U19277 (N_19277,N_19214,N_19097);
nand U19278 (N_19278,N_19014,N_19040);
nand U19279 (N_19279,N_19013,N_19141);
xor U19280 (N_19280,N_19089,N_19129);
xnor U19281 (N_19281,N_19128,N_19245);
nand U19282 (N_19282,N_19102,N_19166);
nand U19283 (N_19283,N_19118,N_19217);
and U19284 (N_19284,N_19145,N_19044);
nor U19285 (N_19285,N_19052,N_19211);
nand U19286 (N_19286,N_19088,N_19080);
and U19287 (N_19287,N_19045,N_19199);
xnor U19288 (N_19288,N_19075,N_19172);
xnor U19289 (N_19289,N_19068,N_19223);
nand U19290 (N_19290,N_19077,N_19190);
or U19291 (N_19291,N_19156,N_19072);
and U19292 (N_19292,N_19161,N_19207);
and U19293 (N_19293,N_19143,N_19047);
xor U19294 (N_19294,N_19154,N_19108);
or U19295 (N_19295,N_19183,N_19186);
or U19296 (N_19296,N_19191,N_19126);
xor U19297 (N_19297,N_19230,N_19204);
and U19298 (N_19298,N_19056,N_19018);
nor U19299 (N_19299,N_19082,N_19023);
xnor U19300 (N_19300,N_19019,N_19200);
nor U19301 (N_19301,N_19124,N_19229);
and U19302 (N_19302,N_19216,N_19169);
nor U19303 (N_19303,N_19003,N_19006);
xor U19304 (N_19304,N_19065,N_19144);
and U19305 (N_19305,N_19074,N_19173);
nand U19306 (N_19306,N_19073,N_19225);
and U19307 (N_19307,N_19162,N_19150);
xor U19308 (N_19308,N_19247,N_19210);
or U19309 (N_19309,N_19004,N_19095);
xor U19310 (N_19310,N_19032,N_19063);
or U19311 (N_19311,N_19196,N_19152);
xnor U19312 (N_19312,N_19219,N_19139);
and U19313 (N_19313,N_19055,N_19130);
or U19314 (N_19314,N_19193,N_19066);
or U19315 (N_19315,N_19239,N_19201);
and U19316 (N_19316,N_19081,N_19236);
nor U19317 (N_19317,N_19036,N_19165);
nor U19318 (N_19318,N_19131,N_19093);
nor U19319 (N_19319,N_19100,N_19048);
nor U19320 (N_19320,N_19206,N_19242);
xor U19321 (N_19321,N_19112,N_19105);
nor U19322 (N_19322,N_19035,N_19017);
or U19323 (N_19323,N_19205,N_19009);
xnor U19324 (N_19324,N_19148,N_19104);
nand U19325 (N_19325,N_19061,N_19147);
xnor U19326 (N_19326,N_19085,N_19146);
xor U19327 (N_19327,N_19110,N_19034);
xnor U19328 (N_19328,N_19078,N_19015);
nand U19329 (N_19329,N_19060,N_19000);
xnor U19330 (N_19330,N_19086,N_19167);
or U19331 (N_19331,N_19069,N_19222);
xor U19332 (N_19332,N_19058,N_19192);
xnor U19333 (N_19333,N_19233,N_19024);
or U19334 (N_19334,N_19180,N_19071);
and U19335 (N_19335,N_19092,N_19083);
xor U19336 (N_19336,N_19025,N_19001);
nand U19337 (N_19337,N_19116,N_19209);
nor U19338 (N_19338,N_19179,N_19113);
xnor U19339 (N_19339,N_19135,N_19054);
xor U19340 (N_19340,N_19151,N_19125);
nand U19341 (N_19341,N_19238,N_19157);
nand U19342 (N_19342,N_19111,N_19164);
xnor U19343 (N_19343,N_19031,N_19243);
xnor U19344 (N_19344,N_19246,N_19043);
nand U19345 (N_19345,N_19240,N_19042);
nor U19346 (N_19346,N_19117,N_19226);
nor U19347 (N_19347,N_19138,N_19090);
or U19348 (N_19348,N_19203,N_19115);
or U19349 (N_19349,N_19103,N_19149);
and U19350 (N_19350,N_19187,N_19059);
nand U19351 (N_19351,N_19027,N_19020);
or U19352 (N_19352,N_19094,N_19039);
nand U19353 (N_19353,N_19184,N_19221);
or U19354 (N_19354,N_19163,N_19096);
nand U19355 (N_19355,N_19159,N_19107);
xnor U19356 (N_19356,N_19008,N_19053);
or U19357 (N_19357,N_19132,N_19007);
or U19358 (N_19358,N_19244,N_19079);
nand U19359 (N_19359,N_19091,N_19070);
nand U19360 (N_19360,N_19026,N_19121);
and U19361 (N_19361,N_19046,N_19101);
nor U19362 (N_19362,N_19177,N_19029);
xnor U19363 (N_19363,N_19106,N_19182);
nor U19364 (N_19364,N_19002,N_19213);
xnor U19365 (N_19365,N_19142,N_19198);
or U19366 (N_19366,N_19109,N_19114);
xor U19367 (N_19367,N_19010,N_19041);
xnor U19368 (N_19368,N_19176,N_19011);
and U19369 (N_19369,N_19170,N_19212);
or U19370 (N_19370,N_19178,N_19051);
and U19371 (N_19371,N_19188,N_19171);
xnor U19372 (N_19372,N_19235,N_19136);
xnor U19373 (N_19373,N_19189,N_19134);
nand U19374 (N_19374,N_19160,N_19194);
xnor U19375 (N_19375,N_19161,N_19131);
or U19376 (N_19376,N_19080,N_19179);
or U19377 (N_19377,N_19162,N_19065);
xor U19378 (N_19378,N_19051,N_19137);
nor U19379 (N_19379,N_19142,N_19131);
nor U19380 (N_19380,N_19056,N_19119);
nand U19381 (N_19381,N_19083,N_19098);
nand U19382 (N_19382,N_19095,N_19225);
or U19383 (N_19383,N_19129,N_19013);
xor U19384 (N_19384,N_19005,N_19100);
or U19385 (N_19385,N_19029,N_19022);
and U19386 (N_19386,N_19071,N_19116);
and U19387 (N_19387,N_19020,N_19111);
or U19388 (N_19388,N_19116,N_19184);
nand U19389 (N_19389,N_19155,N_19072);
or U19390 (N_19390,N_19052,N_19044);
or U19391 (N_19391,N_19188,N_19216);
and U19392 (N_19392,N_19246,N_19102);
nand U19393 (N_19393,N_19162,N_19246);
nand U19394 (N_19394,N_19072,N_19057);
nor U19395 (N_19395,N_19237,N_19106);
nor U19396 (N_19396,N_19136,N_19033);
nor U19397 (N_19397,N_19140,N_19136);
nand U19398 (N_19398,N_19024,N_19232);
xor U19399 (N_19399,N_19186,N_19144);
and U19400 (N_19400,N_19139,N_19119);
nand U19401 (N_19401,N_19077,N_19045);
nand U19402 (N_19402,N_19222,N_19216);
nor U19403 (N_19403,N_19173,N_19183);
or U19404 (N_19404,N_19009,N_19217);
nand U19405 (N_19405,N_19093,N_19071);
nand U19406 (N_19406,N_19108,N_19195);
nand U19407 (N_19407,N_19246,N_19007);
xor U19408 (N_19408,N_19090,N_19071);
and U19409 (N_19409,N_19096,N_19013);
and U19410 (N_19410,N_19241,N_19229);
xnor U19411 (N_19411,N_19164,N_19097);
nor U19412 (N_19412,N_19050,N_19240);
nand U19413 (N_19413,N_19224,N_19073);
and U19414 (N_19414,N_19132,N_19066);
and U19415 (N_19415,N_19123,N_19016);
xor U19416 (N_19416,N_19120,N_19219);
xnor U19417 (N_19417,N_19152,N_19014);
or U19418 (N_19418,N_19064,N_19177);
xor U19419 (N_19419,N_19137,N_19024);
nor U19420 (N_19420,N_19243,N_19057);
and U19421 (N_19421,N_19119,N_19214);
and U19422 (N_19422,N_19226,N_19073);
nand U19423 (N_19423,N_19034,N_19245);
or U19424 (N_19424,N_19032,N_19079);
and U19425 (N_19425,N_19063,N_19191);
xnor U19426 (N_19426,N_19037,N_19042);
or U19427 (N_19427,N_19194,N_19000);
xor U19428 (N_19428,N_19063,N_19209);
or U19429 (N_19429,N_19011,N_19053);
nor U19430 (N_19430,N_19164,N_19177);
nand U19431 (N_19431,N_19244,N_19080);
and U19432 (N_19432,N_19093,N_19176);
nor U19433 (N_19433,N_19073,N_19219);
nand U19434 (N_19434,N_19197,N_19125);
or U19435 (N_19435,N_19069,N_19215);
or U19436 (N_19436,N_19046,N_19171);
or U19437 (N_19437,N_19067,N_19069);
xor U19438 (N_19438,N_19038,N_19207);
nor U19439 (N_19439,N_19160,N_19115);
nand U19440 (N_19440,N_19139,N_19132);
xnor U19441 (N_19441,N_19134,N_19052);
nor U19442 (N_19442,N_19039,N_19014);
or U19443 (N_19443,N_19041,N_19019);
nand U19444 (N_19444,N_19101,N_19133);
or U19445 (N_19445,N_19050,N_19002);
or U19446 (N_19446,N_19085,N_19058);
nand U19447 (N_19447,N_19142,N_19138);
or U19448 (N_19448,N_19230,N_19023);
nor U19449 (N_19449,N_19205,N_19069);
xor U19450 (N_19450,N_19161,N_19197);
and U19451 (N_19451,N_19201,N_19213);
xor U19452 (N_19452,N_19174,N_19011);
nor U19453 (N_19453,N_19188,N_19017);
and U19454 (N_19454,N_19050,N_19165);
and U19455 (N_19455,N_19110,N_19074);
xnor U19456 (N_19456,N_19154,N_19133);
or U19457 (N_19457,N_19204,N_19148);
xor U19458 (N_19458,N_19207,N_19119);
nand U19459 (N_19459,N_19010,N_19022);
and U19460 (N_19460,N_19156,N_19043);
nand U19461 (N_19461,N_19129,N_19208);
xor U19462 (N_19462,N_19010,N_19244);
or U19463 (N_19463,N_19183,N_19157);
xnor U19464 (N_19464,N_19127,N_19011);
and U19465 (N_19465,N_19026,N_19221);
or U19466 (N_19466,N_19217,N_19196);
or U19467 (N_19467,N_19164,N_19016);
or U19468 (N_19468,N_19108,N_19005);
xnor U19469 (N_19469,N_19135,N_19150);
nand U19470 (N_19470,N_19205,N_19130);
or U19471 (N_19471,N_19050,N_19249);
nand U19472 (N_19472,N_19051,N_19143);
nand U19473 (N_19473,N_19128,N_19180);
or U19474 (N_19474,N_19183,N_19002);
xnor U19475 (N_19475,N_19120,N_19025);
and U19476 (N_19476,N_19132,N_19232);
xor U19477 (N_19477,N_19089,N_19067);
xnor U19478 (N_19478,N_19022,N_19239);
nand U19479 (N_19479,N_19240,N_19168);
and U19480 (N_19480,N_19139,N_19057);
xnor U19481 (N_19481,N_19014,N_19164);
xnor U19482 (N_19482,N_19229,N_19199);
nor U19483 (N_19483,N_19035,N_19043);
and U19484 (N_19484,N_19028,N_19035);
nor U19485 (N_19485,N_19076,N_19230);
xor U19486 (N_19486,N_19069,N_19091);
nand U19487 (N_19487,N_19166,N_19044);
and U19488 (N_19488,N_19068,N_19051);
nor U19489 (N_19489,N_19184,N_19031);
and U19490 (N_19490,N_19175,N_19145);
xnor U19491 (N_19491,N_19062,N_19158);
or U19492 (N_19492,N_19139,N_19191);
nor U19493 (N_19493,N_19005,N_19127);
xnor U19494 (N_19494,N_19132,N_19120);
nor U19495 (N_19495,N_19013,N_19107);
or U19496 (N_19496,N_19054,N_19145);
and U19497 (N_19497,N_19137,N_19062);
or U19498 (N_19498,N_19135,N_19204);
nor U19499 (N_19499,N_19110,N_19022);
nand U19500 (N_19500,N_19434,N_19430);
nor U19501 (N_19501,N_19309,N_19490);
and U19502 (N_19502,N_19433,N_19453);
nand U19503 (N_19503,N_19318,N_19258);
xnor U19504 (N_19504,N_19428,N_19385);
xor U19505 (N_19505,N_19404,N_19380);
or U19506 (N_19506,N_19470,N_19423);
and U19507 (N_19507,N_19276,N_19375);
nor U19508 (N_19508,N_19278,N_19326);
or U19509 (N_19509,N_19383,N_19341);
nor U19510 (N_19510,N_19371,N_19499);
nand U19511 (N_19511,N_19292,N_19286);
and U19512 (N_19512,N_19424,N_19478);
or U19513 (N_19513,N_19367,N_19361);
nor U19514 (N_19514,N_19355,N_19397);
xnor U19515 (N_19515,N_19356,N_19271);
xnor U19516 (N_19516,N_19415,N_19317);
nor U19517 (N_19517,N_19483,N_19265);
nor U19518 (N_19518,N_19401,N_19270);
and U19519 (N_19519,N_19310,N_19273);
nand U19520 (N_19520,N_19488,N_19370);
and U19521 (N_19521,N_19438,N_19458);
xnor U19522 (N_19522,N_19452,N_19336);
xnor U19523 (N_19523,N_19477,N_19342);
nor U19524 (N_19524,N_19426,N_19295);
and U19525 (N_19525,N_19436,N_19285);
xor U19526 (N_19526,N_19338,N_19456);
or U19527 (N_19527,N_19260,N_19298);
and U19528 (N_19528,N_19354,N_19360);
xnor U19529 (N_19529,N_19303,N_19384);
nand U19530 (N_19530,N_19254,N_19305);
nand U19531 (N_19531,N_19293,N_19274);
nand U19532 (N_19532,N_19410,N_19474);
nand U19533 (N_19533,N_19297,N_19381);
and U19534 (N_19534,N_19429,N_19431);
xor U19535 (N_19535,N_19376,N_19358);
nor U19536 (N_19536,N_19389,N_19498);
or U19537 (N_19537,N_19422,N_19406);
or U19538 (N_19538,N_19465,N_19302);
nand U19539 (N_19539,N_19301,N_19394);
nor U19540 (N_19540,N_19388,N_19387);
and U19541 (N_19541,N_19340,N_19345);
xnor U19542 (N_19542,N_19497,N_19441);
or U19543 (N_19543,N_19259,N_19476);
nand U19544 (N_19544,N_19275,N_19282);
or U19545 (N_19545,N_19250,N_19251);
and U19546 (N_19546,N_19485,N_19390);
or U19547 (N_19547,N_19427,N_19311);
or U19548 (N_19548,N_19418,N_19405);
or U19549 (N_19549,N_19480,N_19277);
xor U19550 (N_19550,N_19495,N_19432);
nor U19551 (N_19551,N_19268,N_19403);
nand U19552 (N_19552,N_19449,N_19439);
nand U19553 (N_19553,N_19447,N_19473);
xor U19554 (N_19554,N_19409,N_19289);
xor U19555 (N_19555,N_19307,N_19333);
xor U19556 (N_19556,N_19475,N_19442);
nor U19557 (N_19557,N_19471,N_19369);
nand U19558 (N_19558,N_19382,N_19420);
or U19559 (N_19559,N_19462,N_19255);
or U19560 (N_19560,N_19294,N_19283);
or U19561 (N_19561,N_19451,N_19407);
nand U19562 (N_19562,N_19339,N_19335);
or U19563 (N_19563,N_19264,N_19316);
or U19564 (N_19564,N_19445,N_19416);
nand U19565 (N_19565,N_19343,N_19372);
and U19566 (N_19566,N_19398,N_19486);
nor U19567 (N_19567,N_19267,N_19402);
and U19568 (N_19568,N_19469,N_19417);
nor U19569 (N_19569,N_19392,N_19327);
or U19570 (N_19570,N_19257,N_19411);
nand U19571 (N_19571,N_19279,N_19378);
or U19572 (N_19572,N_19466,N_19413);
nor U19573 (N_19573,N_19365,N_19350);
or U19574 (N_19574,N_19314,N_19290);
nor U19575 (N_19575,N_19435,N_19331);
nand U19576 (N_19576,N_19472,N_19368);
and U19577 (N_19577,N_19252,N_19308);
nand U19578 (N_19578,N_19332,N_19287);
xor U19579 (N_19579,N_19379,N_19306);
xor U19580 (N_19580,N_19324,N_19304);
or U19581 (N_19581,N_19443,N_19359);
and U19582 (N_19582,N_19344,N_19351);
nand U19583 (N_19583,N_19347,N_19364);
and U19584 (N_19584,N_19496,N_19353);
nor U19585 (N_19585,N_19377,N_19269);
or U19586 (N_19586,N_19312,N_19349);
xor U19587 (N_19587,N_19446,N_19395);
xnor U19588 (N_19588,N_19479,N_19284);
nor U19589 (N_19589,N_19459,N_19357);
nor U19590 (N_19590,N_19337,N_19440);
xor U19591 (N_19591,N_19280,N_19281);
xnor U19592 (N_19592,N_19363,N_19300);
nand U19593 (N_19593,N_19487,N_19322);
xnor U19594 (N_19594,N_19492,N_19455);
nand U19595 (N_19595,N_19464,N_19315);
or U19596 (N_19596,N_19329,N_19493);
and U19597 (N_19597,N_19334,N_19467);
and U19598 (N_19598,N_19412,N_19450);
and U19599 (N_19599,N_19468,N_19373);
nor U19600 (N_19600,N_19481,N_19419);
and U19601 (N_19601,N_19484,N_19457);
and U19602 (N_19602,N_19346,N_19393);
and U19603 (N_19603,N_19319,N_19253);
and U19604 (N_19604,N_19425,N_19272);
or U19605 (N_19605,N_19256,N_19461);
and U19606 (N_19606,N_19321,N_19299);
nor U19607 (N_19607,N_19261,N_19352);
or U19608 (N_19608,N_19494,N_19266);
or U19609 (N_19609,N_19328,N_19291);
or U19610 (N_19610,N_19399,N_19391);
nor U19611 (N_19611,N_19288,N_19320);
nor U19612 (N_19612,N_19482,N_19323);
or U19613 (N_19613,N_19491,N_19374);
and U19614 (N_19614,N_19448,N_19348);
nor U19615 (N_19615,N_19386,N_19366);
nor U19616 (N_19616,N_19444,N_19463);
or U19617 (N_19617,N_19489,N_19414);
or U19618 (N_19618,N_19454,N_19460);
or U19619 (N_19619,N_19263,N_19362);
or U19620 (N_19620,N_19396,N_19262);
nor U19621 (N_19621,N_19437,N_19421);
nor U19622 (N_19622,N_19330,N_19313);
nor U19623 (N_19623,N_19325,N_19296);
nor U19624 (N_19624,N_19400,N_19408);
nor U19625 (N_19625,N_19310,N_19281);
xor U19626 (N_19626,N_19364,N_19487);
xnor U19627 (N_19627,N_19345,N_19436);
nand U19628 (N_19628,N_19470,N_19427);
or U19629 (N_19629,N_19492,N_19497);
or U19630 (N_19630,N_19451,N_19401);
and U19631 (N_19631,N_19289,N_19399);
and U19632 (N_19632,N_19319,N_19460);
and U19633 (N_19633,N_19429,N_19407);
nand U19634 (N_19634,N_19349,N_19292);
and U19635 (N_19635,N_19317,N_19329);
and U19636 (N_19636,N_19428,N_19347);
xor U19637 (N_19637,N_19284,N_19312);
nand U19638 (N_19638,N_19305,N_19436);
nor U19639 (N_19639,N_19333,N_19383);
and U19640 (N_19640,N_19363,N_19258);
nand U19641 (N_19641,N_19323,N_19396);
nor U19642 (N_19642,N_19337,N_19482);
and U19643 (N_19643,N_19498,N_19420);
and U19644 (N_19644,N_19344,N_19368);
nor U19645 (N_19645,N_19449,N_19261);
nand U19646 (N_19646,N_19281,N_19282);
nand U19647 (N_19647,N_19493,N_19294);
and U19648 (N_19648,N_19442,N_19477);
nand U19649 (N_19649,N_19492,N_19277);
or U19650 (N_19650,N_19262,N_19432);
xnor U19651 (N_19651,N_19372,N_19281);
or U19652 (N_19652,N_19416,N_19328);
xnor U19653 (N_19653,N_19320,N_19452);
and U19654 (N_19654,N_19278,N_19461);
or U19655 (N_19655,N_19495,N_19429);
nor U19656 (N_19656,N_19419,N_19316);
nor U19657 (N_19657,N_19424,N_19275);
and U19658 (N_19658,N_19250,N_19341);
and U19659 (N_19659,N_19257,N_19394);
nand U19660 (N_19660,N_19309,N_19470);
xnor U19661 (N_19661,N_19434,N_19444);
and U19662 (N_19662,N_19405,N_19278);
nand U19663 (N_19663,N_19448,N_19409);
and U19664 (N_19664,N_19444,N_19426);
nand U19665 (N_19665,N_19390,N_19445);
nand U19666 (N_19666,N_19487,N_19338);
nor U19667 (N_19667,N_19493,N_19425);
and U19668 (N_19668,N_19490,N_19467);
xor U19669 (N_19669,N_19429,N_19365);
nor U19670 (N_19670,N_19329,N_19281);
nor U19671 (N_19671,N_19352,N_19469);
nor U19672 (N_19672,N_19462,N_19429);
nor U19673 (N_19673,N_19326,N_19293);
or U19674 (N_19674,N_19363,N_19296);
nor U19675 (N_19675,N_19269,N_19429);
nand U19676 (N_19676,N_19346,N_19252);
and U19677 (N_19677,N_19458,N_19268);
or U19678 (N_19678,N_19393,N_19381);
or U19679 (N_19679,N_19370,N_19297);
or U19680 (N_19680,N_19250,N_19432);
nor U19681 (N_19681,N_19423,N_19321);
xnor U19682 (N_19682,N_19369,N_19308);
and U19683 (N_19683,N_19321,N_19344);
or U19684 (N_19684,N_19253,N_19286);
xnor U19685 (N_19685,N_19337,N_19443);
nor U19686 (N_19686,N_19359,N_19413);
and U19687 (N_19687,N_19473,N_19331);
or U19688 (N_19688,N_19356,N_19474);
nand U19689 (N_19689,N_19330,N_19431);
and U19690 (N_19690,N_19286,N_19256);
nand U19691 (N_19691,N_19256,N_19372);
nand U19692 (N_19692,N_19376,N_19396);
or U19693 (N_19693,N_19471,N_19265);
and U19694 (N_19694,N_19433,N_19334);
nor U19695 (N_19695,N_19379,N_19464);
nand U19696 (N_19696,N_19271,N_19464);
or U19697 (N_19697,N_19269,N_19471);
or U19698 (N_19698,N_19371,N_19412);
and U19699 (N_19699,N_19406,N_19360);
or U19700 (N_19700,N_19271,N_19466);
nor U19701 (N_19701,N_19446,N_19287);
nand U19702 (N_19702,N_19371,N_19263);
xnor U19703 (N_19703,N_19425,N_19461);
nand U19704 (N_19704,N_19338,N_19477);
nand U19705 (N_19705,N_19251,N_19322);
or U19706 (N_19706,N_19422,N_19381);
or U19707 (N_19707,N_19462,N_19370);
and U19708 (N_19708,N_19295,N_19469);
and U19709 (N_19709,N_19462,N_19400);
nor U19710 (N_19710,N_19293,N_19433);
nand U19711 (N_19711,N_19348,N_19440);
xor U19712 (N_19712,N_19396,N_19258);
and U19713 (N_19713,N_19477,N_19317);
nor U19714 (N_19714,N_19471,N_19281);
or U19715 (N_19715,N_19474,N_19466);
nor U19716 (N_19716,N_19420,N_19418);
nand U19717 (N_19717,N_19309,N_19357);
xnor U19718 (N_19718,N_19367,N_19289);
or U19719 (N_19719,N_19443,N_19492);
or U19720 (N_19720,N_19255,N_19317);
nor U19721 (N_19721,N_19424,N_19406);
or U19722 (N_19722,N_19402,N_19325);
and U19723 (N_19723,N_19494,N_19299);
xnor U19724 (N_19724,N_19363,N_19265);
nor U19725 (N_19725,N_19358,N_19313);
nand U19726 (N_19726,N_19470,N_19328);
xnor U19727 (N_19727,N_19484,N_19345);
nor U19728 (N_19728,N_19325,N_19496);
and U19729 (N_19729,N_19489,N_19336);
or U19730 (N_19730,N_19432,N_19465);
xor U19731 (N_19731,N_19404,N_19409);
and U19732 (N_19732,N_19406,N_19303);
xor U19733 (N_19733,N_19334,N_19300);
nand U19734 (N_19734,N_19413,N_19351);
nor U19735 (N_19735,N_19406,N_19353);
and U19736 (N_19736,N_19439,N_19307);
nor U19737 (N_19737,N_19397,N_19437);
nor U19738 (N_19738,N_19362,N_19282);
xnor U19739 (N_19739,N_19475,N_19431);
or U19740 (N_19740,N_19265,N_19254);
and U19741 (N_19741,N_19433,N_19280);
and U19742 (N_19742,N_19341,N_19284);
xnor U19743 (N_19743,N_19377,N_19288);
nand U19744 (N_19744,N_19435,N_19361);
and U19745 (N_19745,N_19381,N_19432);
nor U19746 (N_19746,N_19468,N_19430);
nand U19747 (N_19747,N_19453,N_19324);
and U19748 (N_19748,N_19382,N_19443);
nor U19749 (N_19749,N_19399,N_19495);
nor U19750 (N_19750,N_19610,N_19569);
and U19751 (N_19751,N_19727,N_19740);
nand U19752 (N_19752,N_19628,N_19514);
and U19753 (N_19753,N_19599,N_19724);
xnor U19754 (N_19754,N_19605,N_19548);
or U19755 (N_19755,N_19613,N_19539);
nor U19756 (N_19756,N_19572,N_19729);
and U19757 (N_19757,N_19525,N_19591);
nor U19758 (N_19758,N_19711,N_19732);
nand U19759 (N_19759,N_19547,N_19576);
nand U19760 (N_19760,N_19618,N_19719);
and U19761 (N_19761,N_19556,N_19667);
nand U19762 (N_19762,N_19688,N_19554);
nor U19763 (N_19763,N_19635,N_19701);
nor U19764 (N_19764,N_19694,N_19677);
or U19765 (N_19765,N_19606,N_19670);
and U19766 (N_19766,N_19654,N_19617);
and U19767 (N_19767,N_19717,N_19524);
nand U19768 (N_19768,N_19523,N_19515);
nand U19769 (N_19769,N_19693,N_19546);
or U19770 (N_19770,N_19535,N_19520);
and U19771 (N_19771,N_19638,N_19622);
nor U19772 (N_19772,N_19623,N_19682);
nor U19773 (N_19773,N_19699,N_19544);
and U19774 (N_19774,N_19681,N_19716);
or U19775 (N_19775,N_19709,N_19584);
nor U19776 (N_19776,N_19646,N_19602);
nand U19777 (N_19777,N_19692,N_19721);
xor U19778 (N_19778,N_19660,N_19714);
and U19779 (N_19779,N_19537,N_19615);
and U19780 (N_19780,N_19695,N_19550);
nand U19781 (N_19781,N_19552,N_19668);
xor U19782 (N_19782,N_19737,N_19634);
xnor U19783 (N_19783,N_19558,N_19508);
and U19784 (N_19784,N_19565,N_19577);
xnor U19785 (N_19785,N_19506,N_19704);
xor U19786 (N_19786,N_19531,N_19590);
nand U19787 (N_19787,N_19560,N_19522);
xnor U19788 (N_19788,N_19671,N_19648);
nor U19789 (N_19789,N_19609,N_19553);
or U19790 (N_19790,N_19647,N_19627);
or U19791 (N_19791,N_19629,N_19510);
or U19792 (N_19792,N_19662,N_19595);
nand U19793 (N_19793,N_19529,N_19509);
nand U19794 (N_19794,N_19549,N_19641);
nor U19795 (N_19795,N_19561,N_19749);
nor U19796 (N_19796,N_19645,N_19663);
or U19797 (N_19797,N_19652,N_19518);
xor U19798 (N_19798,N_19715,N_19587);
and U19799 (N_19799,N_19567,N_19642);
xor U19800 (N_19800,N_19726,N_19744);
and U19801 (N_19801,N_19574,N_19538);
or U19802 (N_19802,N_19702,N_19637);
nor U19803 (N_19803,N_19707,N_19748);
and U19804 (N_19804,N_19739,N_19517);
xor U19805 (N_19805,N_19728,N_19666);
nand U19806 (N_19806,N_19564,N_19706);
and U19807 (N_19807,N_19683,N_19588);
nor U19808 (N_19808,N_19612,N_19579);
and U19809 (N_19809,N_19733,N_19516);
nand U19810 (N_19810,N_19700,N_19734);
nand U19811 (N_19811,N_19527,N_19689);
nor U19812 (N_19812,N_19691,N_19745);
xnor U19813 (N_19813,N_19686,N_19665);
nor U19814 (N_19814,N_19586,N_19644);
or U19815 (N_19815,N_19601,N_19608);
nand U19816 (N_19816,N_19626,N_19532);
and U19817 (N_19817,N_19673,N_19543);
or U19818 (N_19818,N_19541,N_19607);
and U19819 (N_19819,N_19675,N_19680);
or U19820 (N_19820,N_19621,N_19712);
nand U19821 (N_19821,N_19685,N_19659);
nand U19822 (N_19822,N_19743,N_19513);
nor U19823 (N_19823,N_19710,N_19722);
xor U19824 (N_19824,N_19505,N_19697);
xnor U19825 (N_19825,N_19557,N_19708);
nor U19826 (N_19826,N_19585,N_19746);
xnor U19827 (N_19827,N_19578,N_19600);
and U19828 (N_19828,N_19519,N_19649);
nand U19829 (N_19829,N_19718,N_19619);
nand U19830 (N_19830,N_19632,N_19583);
nand U19831 (N_19831,N_19720,N_19503);
or U19832 (N_19832,N_19723,N_19611);
or U19833 (N_19833,N_19542,N_19575);
nand U19834 (N_19834,N_19676,N_19528);
nand U19835 (N_19835,N_19551,N_19526);
and U19836 (N_19836,N_19684,N_19616);
and U19837 (N_19837,N_19533,N_19713);
nand U19838 (N_19838,N_19568,N_19573);
and U19839 (N_19839,N_19580,N_19566);
and U19840 (N_19840,N_19594,N_19636);
and U19841 (N_19841,N_19731,N_19624);
and U19842 (N_19842,N_19614,N_19512);
nor U19843 (N_19843,N_19678,N_19511);
nor U19844 (N_19844,N_19559,N_19598);
and U19845 (N_19845,N_19501,N_19653);
or U19846 (N_19846,N_19603,N_19639);
xor U19847 (N_19847,N_19597,N_19521);
and U19848 (N_19848,N_19742,N_19650);
and U19849 (N_19849,N_19536,N_19655);
nand U19850 (N_19850,N_19725,N_19589);
nor U19851 (N_19851,N_19570,N_19705);
nor U19852 (N_19852,N_19504,N_19730);
nor U19853 (N_19853,N_19596,N_19620);
and U19854 (N_19854,N_19604,N_19738);
nor U19855 (N_19855,N_19657,N_19679);
or U19856 (N_19856,N_19690,N_19656);
or U19857 (N_19857,N_19582,N_19640);
nor U19858 (N_19858,N_19631,N_19563);
nand U19859 (N_19859,N_19661,N_19530);
and U19860 (N_19860,N_19633,N_19674);
nand U19861 (N_19861,N_19555,N_19672);
xor U19862 (N_19862,N_19545,N_19625);
or U19863 (N_19863,N_19540,N_19736);
or U19864 (N_19864,N_19534,N_19502);
or U19865 (N_19865,N_19562,N_19571);
or U19866 (N_19866,N_19630,N_19643);
nor U19867 (N_19867,N_19592,N_19703);
xor U19868 (N_19868,N_19651,N_19664);
nand U19869 (N_19869,N_19687,N_19500);
xor U19870 (N_19870,N_19669,N_19507);
xor U19871 (N_19871,N_19735,N_19696);
nor U19872 (N_19872,N_19698,N_19658);
nor U19873 (N_19873,N_19747,N_19741);
nor U19874 (N_19874,N_19593,N_19581);
and U19875 (N_19875,N_19634,N_19743);
nor U19876 (N_19876,N_19561,N_19606);
xnor U19877 (N_19877,N_19606,N_19728);
nor U19878 (N_19878,N_19559,N_19731);
nor U19879 (N_19879,N_19611,N_19633);
or U19880 (N_19880,N_19720,N_19709);
nand U19881 (N_19881,N_19576,N_19584);
xor U19882 (N_19882,N_19557,N_19707);
nor U19883 (N_19883,N_19602,N_19508);
xnor U19884 (N_19884,N_19563,N_19572);
and U19885 (N_19885,N_19565,N_19621);
xor U19886 (N_19886,N_19542,N_19697);
nor U19887 (N_19887,N_19674,N_19592);
and U19888 (N_19888,N_19502,N_19596);
nand U19889 (N_19889,N_19730,N_19720);
nor U19890 (N_19890,N_19602,N_19679);
nor U19891 (N_19891,N_19679,N_19715);
nor U19892 (N_19892,N_19631,N_19539);
or U19893 (N_19893,N_19690,N_19541);
nand U19894 (N_19894,N_19654,N_19567);
nand U19895 (N_19895,N_19697,N_19722);
nor U19896 (N_19896,N_19726,N_19634);
or U19897 (N_19897,N_19561,N_19627);
nand U19898 (N_19898,N_19500,N_19606);
or U19899 (N_19899,N_19630,N_19728);
xor U19900 (N_19900,N_19501,N_19595);
xnor U19901 (N_19901,N_19505,N_19604);
or U19902 (N_19902,N_19537,N_19504);
nor U19903 (N_19903,N_19577,N_19548);
nor U19904 (N_19904,N_19746,N_19524);
nand U19905 (N_19905,N_19629,N_19728);
nor U19906 (N_19906,N_19625,N_19718);
nand U19907 (N_19907,N_19641,N_19711);
and U19908 (N_19908,N_19679,N_19640);
and U19909 (N_19909,N_19646,N_19655);
nand U19910 (N_19910,N_19509,N_19658);
and U19911 (N_19911,N_19571,N_19715);
and U19912 (N_19912,N_19703,N_19643);
nor U19913 (N_19913,N_19500,N_19559);
xnor U19914 (N_19914,N_19691,N_19614);
nand U19915 (N_19915,N_19639,N_19516);
xor U19916 (N_19916,N_19676,N_19707);
and U19917 (N_19917,N_19519,N_19667);
nor U19918 (N_19918,N_19732,N_19741);
nand U19919 (N_19919,N_19504,N_19502);
xor U19920 (N_19920,N_19512,N_19717);
nor U19921 (N_19921,N_19728,N_19586);
and U19922 (N_19922,N_19741,N_19700);
nor U19923 (N_19923,N_19624,N_19674);
and U19924 (N_19924,N_19719,N_19624);
xor U19925 (N_19925,N_19691,N_19595);
or U19926 (N_19926,N_19532,N_19647);
xor U19927 (N_19927,N_19629,N_19674);
nor U19928 (N_19928,N_19639,N_19545);
or U19929 (N_19929,N_19518,N_19660);
nand U19930 (N_19930,N_19720,N_19510);
nand U19931 (N_19931,N_19714,N_19713);
and U19932 (N_19932,N_19570,N_19590);
and U19933 (N_19933,N_19585,N_19602);
nor U19934 (N_19934,N_19523,N_19572);
nand U19935 (N_19935,N_19506,N_19622);
xor U19936 (N_19936,N_19696,N_19515);
or U19937 (N_19937,N_19714,N_19611);
nor U19938 (N_19938,N_19714,N_19598);
xor U19939 (N_19939,N_19724,N_19690);
nor U19940 (N_19940,N_19528,N_19585);
or U19941 (N_19941,N_19623,N_19588);
or U19942 (N_19942,N_19608,N_19645);
xor U19943 (N_19943,N_19630,N_19740);
nor U19944 (N_19944,N_19700,N_19718);
nor U19945 (N_19945,N_19633,N_19520);
and U19946 (N_19946,N_19535,N_19532);
xor U19947 (N_19947,N_19651,N_19649);
and U19948 (N_19948,N_19663,N_19622);
nand U19949 (N_19949,N_19747,N_19711);
or U19950 (N_19950,N_19506,N_19691);
nand U19951 (N_19951,N_19740,N_19645);
nand U19952 (N_19952,N_19684,N_19724);
nor U19953 (N_19953,N_19680,N_19518);
and U19954 (N_19954,N_19679,N_19555);
nand U19955 (N_19955,N_19746,N_19535);
nand U19956 (N_19956,N_19622,N_19702);
xnor U19957 (N_19957,N_19511,N_19542);
or U19958 (N_19958,N_19666,N_19693);
nor U19959 (N_19959,N_19671,N_19734);
xnor U19960 (N_19960,N_19575,N_19645);
nor U19961 (N_19961,N_19593,N_19699);
xor U19962 (N_19962,N_19554,N_19615);
xor U19963 (N_19963,N_19742,N_19612);
or U19964 (N_19964,N_19591,N_19599);
xor U19965 (N_19965,N_19640,N_19513);
xnor U19966 (N_19966,N_19621,N_19557);
xnor U19967 (N_19967,N_19612,N_19704);
xnor U19968 (N_19968,N_19636,N_19668);
and U19969 (N_19969,N_19551,N_19646);
xnor U19970 (N_19970,N_19607,N_19673);
or U19971 (N_19971,N_19568,N_19628);
and U19972 (N_19972,N_19546,N_19655);
or U19973 (N_19973,N_19613,N_19522);
nor U19974 (N_19974,N_19695,N_19740);
nor U19975 (N_19975,N_19521,N_19693);
or U19976 (N_19976,N_19624,N_19557);
nor U19977 (N_19977,N_19540,N_19600);
nor U19978 (N_19978,N_19507,N_19599);
or U19979 (N_19979,N_19506,N_19535);
nand U19980 (N_19980,N_19631,N_19667);
xor U19981 (N_19981,N_19692,N_19704);
nor U19982 (N_19982,N_19692,N_19625);
nor U19983 (N_19983,N_19718,N_19507);
xor U19984 (N_19984,N_19626,N_19545);
nor U19985 (N_19985,N_19668,N_19603);
nand U19986 (N_19986,N_19579,N_19738);
nor U19987 (N_19987,N_19706,N_19613);
xor U19988 (N_19988,N_19731,N_19712);
or U19989 (N_19989,N_19598,N_19698);
nand U19990 (N_19990,N_19625,N_19515);
and U19991 (N_19991,N_19602,N_19658);
and U19992 (N_19992,N_19541,N_19657);
or U19993 (N_19993,N_19571,N_19691);
and U19994 (N_19994,N_19637,N_19609);
xor U19995 (N_19995,N_19696,N_19521);
xor U19996 (N_19996,N_19572,N_19676);
xnor U19997 (N_19997,N_19574,N_19627);
or U19998 (N_19998,N_19659,N_19582);
xnor U19999 (N_19999,N_19542,N_19717);
or U20000 (N_20000,N_19848,N_19956);
xnor U20001 (N_20001,N_19852,N_19867);
and U20002 (N_20002,N_19997,N_19819);
nand U20003 (N_20003,N_19826,N_19978);
xnor U20004 (N_20004,N_19966,N_19797);
and U20005 (N_20005,N_19962,N_19950);
nor U20006 (N_20006,N_19992,N_19839);
or U20007 (N_20007,N_19779,N_19930);
nor U20008 (N_20008,N_19921,N_19878);
or U20009 (N_20009,N_19975,N_19995);
or U20010 (N_20010,N_19874,N_19943);
nand U20011 (N_20011,N_19769,N_19977);
nand U20012 (N_20012,N_19803,N_19946);
nand U20013 (N_20013,N_19861,N_19855);
nand U20014 (N_20014,N_19818,N_19792);
and U20015 (N_20015,N_19845,N_19881);
and U20016 (N_20016,N_19775,N_19888);
or U20017 (N_20017,N_19873,N_19938);
and U20018 (N_20018,N_19784,N_19964);
xor U20019 (N_20019,N_19804,N_19916);
or U20020 (N_20020,N_19915,N_19924);
xnor U20021 (N_20021,N_19970,N_19751);
and U20022 (N_20022,N_19833,N_19863);
nand U20023 (N_20023,N_19788,N_19894);
nand U20024 (N_20024,N_19778,N_19822);
and U20025 (N_20025,N_19882,N_19942);
nor U20026 (N_20026,N_19851,N_19911);
nor U20027 (N_20027,N_19860,N_19947);
xnor U20028 (N_20028,N_19890,N_19896);
nor U20029 (N_20029,N_19759,N_19862);
nor U20030 (N_20030,N_19794,N_19866);
or U20031 (N_20031,N_19774,N_19982);
nand U20032 (N_20032,N_19892,N_19791);
nand U20033 (N_20033,N_19996,N_19815);
nand U20034 (N_20034,N_19941,N_19891);
xnor U20035 (N_20035,N_19802,N_19805);
xnor U20036 (N_20036,N_19953,N_19770);
or U20037 (N_20037,N_19944,N_19918);
or U20038 (N_20038,N_19875,N_19776);
nor U20039 (N_20039,N_19868,N_19999);
or U20040 (N_20040,N_19903,N_19793);
nor U20041 (N_20041,N_19898,N_19799);
nand U20042 (N_20042,N_19893,N_19780);
and U20043 (N_20043,N_19787,N_19974);
and U20044 (N_20044,N_19902,N_19828);
nor U20045 (N_20045,N_19883,N_19807);
or U20046 (N_20046,N_19773,N_19800);
and U20047 (N_20047,N_19831,N_19785);
or U20048 (N_20048,N_19864,N_19857);
nand U20049 (N_20049,N_19981,N_19765);
xor U20050 (N_20050,N_19917,N_19935);
nand U20051 (N_20051,N_19920,N_19912);
nor U20052 (N_20052,N_19909,N_19789);
or U20053 (N_20053,N_19990,N_19919);
nor U20054 (N_20054,N_19786,N_19980);
or U20055 (N_20055,N_19767,N_19993);
or U20056 (N_20056,N_19931,N_19754);
and U20057 (N_20057,N_19764,N_19832);
nor U20058 (N_20058,N_19936,N_19923);
nor U20059 (N_20059,N_19844,N_19985);
nor U20060 (N_20060,N_19817,N_19922);
xor U20061 (N_20061,N_19809,N_19963);
nor U20062 (N_20062,N_19979,N_19972);
nand U20063 (N_20063,N_19820,N_19823);
xnor U20064 (N_20064,N_19856,N_19932);
nor U20065 (N_20065,N_19762,N_19782);
nand U20066 (N_20066,N_19959,N_19954);
and U20067 (N_20067,N_19795,N_19937);
nand U20068 (N_20068,N_19879,N_19991);
nand U20069 (N_20069,N_19854,N_19830);
or U20070 (N_20070,N_19814,N_19900);
nor U20071 (N_20071,N_19812,N_19842);
or U20072 (N_20072,N_19834,N_19934);
xor U20073 (N_20073,N_19870,N_19836);
or U20074 (N_20074,N_19756,N_19885);
and U20075 (N_20075,N_19984,N_19927);
xnor U20076 (N_20076,N_19808,N_19824);
xnor U20077 (N_20077,N_19829,N_19772);
xnor U20078 (N_20078,N_19987,N_19886);
or U20079 (N_20079,N_19955,N_19929);
nor U20080 (N_20080,N_19957,N_19761);
xnor U20081 (N_20081,N_19968,N_19766);
or U20082 (N_20082,N_19887,N_19847);
nand U20083 (N_20083,N_19880,N_19849);
nand U20084 (N_20084,N_19825,N_19869);
nand U20085 (N_20085,N_19960,N_19948);
nor U20086 (N_20086,N_19925,N_19877);
nor U20087 (N_20087,N_19910,N_19904);
nand U20088 (N_20088,N_19965,N_19850);
xnor U20089 (N_20089,N_19895,N_19913);
and U20090 (N_20090,N_19926,N_19958);
xnor U20091 (N_20091,N_19859,N_19945);
nor U20092 (N_20092,N_19889,N_19906);
and U20093 (N_20093,N_19901,N_19988);
nor U20094 (N_20094,N_19755,N_19994);
xor U20095 (N_20095,N_19949,N_19908);
nand U20096 (N_20096,N_19837,N_19760);
and U20097 (N_20097,N_19976,N_19752);
or U20098 (N_20098,N_19983,N_19853);
nand U20099 (N_20099,N_19781,N_19810);
or U20100 (N_20100,N_19928,N_19969);
nand U20101 (N_20101,N_19806,N_19757);
nor U20102 (N_20102,N_19940,N_19865);
or U20103 (N_20103,N_19884,N_19967);
nand U20104 (N_20104,N_19858,N_19872);
xor U20105 (N_20105,N_19798,N_19783);
nor U20106 (N_20106,N_19939,N_19827);
nand U20107 (N_20107,N_19986,N_19811);
nor U20108 (N_20108,N_19971,N_19907);
and U20109 (N_20109,N_19841,N_19871);
nand U20110 (N_20110,N_19801,N_19768);
and U20111 (N_20111,N_19840,N_19821);
nor U20112 (N_20112,N_19843,N_19989);
nand U20113 (N_20113,N_19973,N_19914);
xnor U20114 (N_20114,N_19846,N_19753);
nor U20115 (N_20115,N_19899,N_19777);
nor U20116 (N_20116,N_19813,N_19758);
xnor U20117 (N_20117,N_19951,N_19816);
and U20118 (N_20118,N_19961,N_19905);
nand U20119 (N_20119,N_19998,N_19838);
or U20120 (N_20120,N_19771,N_19952);
xnor U20121 (N_20121,N_19790,N_19750);
nor U20122 (N_20122,N_19835,N_19897);
and U20123 (N_20123,N_19796,N_19876);
xor U20124 (N_20124,N_19933,N_19763);
or U20125 (N_20125,N_19946,N_19828);
and U20126 (N_20126,N_19935,N_19883);
or U20127 (N_20127,N_19911,N_19771);
nor U20128 (N_20128,N_19934,N_19825);
or U20129 (N_20129,N_19961,N_19858);
nor U20130 (N_20130,N_19819,N_19906);
or U20131 (N_20131,N_19982,N_19928);
nand U20132 (N_20132,N_19961,N_19808);
nand U20133 (N_20133,N_19850,N_19838);
and U20134 (N_20134,N_19991,N_19840);
xor U20135 (N_20135,N_19808,N_19797);
xnor U20136 (N_20136,N_19938,N_19850);
and U20137 (N_20137,N_19851,N_19865);
or U20138 (N_20138,N_19981,N_19885);
and U20139 (N_20139,N_19815,N_19932);
and U20140 (N_20140,N_19999,N_19845);
or U20141 (N_20141,N_19904,N_19924);
and U20142 (N_20142,N_19882,N_19808);
nand U20143 (N_20143,N_19784,N_19891);
and U20144 (N_20144,N_19865,N_19870);
and U20145 (N_20145,N_19789,N_19771);
or U20146 (N_20146,N_19791,N_19905);
nand U20147 (N_20147,N_19882,N_19912);
xnor U20148 (N_20148,N_19984,N_19801);
nand U20149 (N_20149,N_19765,N_19842);
or U20150 (N_20150,N_19835,N_19991);
nand U20151 (N_20151,N_19817,N_19982);
nor U20152 (N_20152,N_19962,N_19764);
xor U20153 (N_20153,N_19863,N_19981);
nand U20154 (N_20154,N_19893,N_19765);
or U20155 (N_20155,N_19876,N_19859);
and U20156 (N_20156,N_19986,N_19965);
nand U20157 (N_20157,N_19797,N_19918);
and U20158 (N_20158,N_19838,N_19889);
nor U20159 (N_20159,N_19893,N_19926);
and U20160 (N_20160,N_19808,N_19807);
nor U20161 (N_20161,N_19886,N_19758);
nor U20162 (N_20162,N_19898,N_19911);
xor U20163 (N_20163,N_19902,N_19787);
or U20164 (N_20164,N_19812,N_19920);
nor U20165 (N_20165,N_19775,N_19970);
and U20166 (N_20166,N_19883,N_19789);
xor U20167 (N_20167,N_19839,N_19780);
and U20168 (N_20168,N_19941,N_19944);
nand U20169 (N_20169,N_19805,N_19875);
and U20170 (N_20170,N_19862,N_19777);
nand U20171 (N_20171,N_19972,N_19866);
and U20172 (N_20172,N_19893,N_19868);
nand U20173 (N_20173,N_19866,N_19863);
or U20174 (N_20174,N_19904,N_19845);
nor U20175 (N_20175,N_19835,N_19753);
and U20176 (N_20176,N_19770,N_19834);
and U20177 (N_20177,N_19853,N_19879);
nor U20178 (N_20178,N_19901,N_19968);
and U20179 (N_20179,N_19761,N_19843);
xor U20180 (N_20180,N_19941,N_19853);
and U20181 (N_20181,N_19893,N_19930);
xnor U20182 (N_20182,N_19754,N_19820);
and U20183 (N_20183,N_19765,N_19958);
and U20184 (N_20184,N_19917,N_19971);
nor U20185 (N_20185,N_19959,N_19869);
or U20186 (N_20186,N_19896,N_19933);
or U20187 (N_20187,N_19974,N_19888);
xor U20188 (N_20188,N_19978,N_19885);
xor U20189 (N_20189,N_19827,N_19945);
or U20190 (N_20190,N_19818,N_19957);
or U20191 (N_20191,N_19862,N_19860);
nand U20192 (N_20192,N_19777,N_19839);
xnor U20193 (N_20193,N_19982,N_19925);
or U20194 (N_20194,N_19935,N_19979);
and U20195 (N_20195,N_19846,N_19965);
and U20196 (N_20196,N_19842,N_19793);
xor U20197 (N_20197,N_19830,N_19866);
and U20198 (N_20198,N_19997,N_19833);
xor U20199 (N_20199,N_19869,N_19890);
xor U20200 (N_20200,N_19779,N_19878);
xor U20201 (N_20201,N_19907,N_19856);
nand U20202 (N_20202,N_19906,N_19752);
and U20203 (N_20203,N_19796,N_19851);
xnor U20204 (N_20204,N_19772,N_19891);
nand U20205 (N_20205,N_19863,N_19955);
or U20206 (N_20206,N_19896,N_19864);
or U20207 (N_20207,N_19939,N_19805);
nor U20208 (N_20208,N_19839,N_19873);
and U20209 (N_20209,N_19828,N_19751);
and U20210 (N_20210,N_19830,N_19933);
and U20211 (N_20211,N_19939,N_19849);
xor U20212 (N_20212,N_19817,N_19990);
nor U20213 (N_20213,N_19869,N_19996);
or U20214 (N_20214,N_19909,N_19868);
and U20215 (N_20215,N_19931,N_19906);
nor U20216 (N_20216,N_19963,N_19974);
nor U20217 (N_20217,N_19876,N_19752);
or U20218 (N_20218,N_19895,N_19808);
xor U20219 (N_20219,N_19880,N_19754);
nor U20220 (N_20220,N_19965,N_19980);
nand U20221 (N_20221,N_19946,N_19860);
nor U20222 (N_20222,N_19984,N_19916);
nand U20223 (N_20223,N_19765,N_19829);
nor U20224 (N_20224,N_19960,N_19900);
nand U20225 (N_20225,N_19868,N_19947);
and U20226 (N_20226,N_19988,N_19995);
and U20227 (N_20227,N_19829,N_19898);
and U20228 (N_20228,N_19997,N_19856);
nand U20229 (N_20229,N_19807,N_19968);
or U20230 (N_20230,N_19869,N_19902);
nand U20231 (N_20231,N_19974,N_19764);
or U20232 (N_20232,N_19942,N_19938);
and U20233 (N_20233,N_19957,N_19940);
nor U20234 (N_20234,N_19864,N_19898);
nand U20235 (N_20235,N_19760,N_19783);
nor U20236 (N_20236,N_19786,N_19802);
nand U20237 (N_20237,N_19840,N_19787);
or U20238 (N_20238,N_19849,N_19851);
nand U20239 (N_20239,N_19936,N_19909);
nand U20240 (N_20240,N_19845,N_19847);
nand U20241 (N_20241,N_19804,N_19957);
nand U20242 (N_20242,N_19947,N_19960);
nand U20243 (N_20243,N_19828,N_19933);
or U20244 (N_20244,N_19802,N_19956);
nand U20245 (N_20245,N_19903,N_19998);
and U20246 (N_20246,N_19878,N_19867);
nand U20247 (N_20247,N_19919,N_19784);
nand U20248 (N_20248,N_19864,N_19881);
nor U20249 (N_20249,N_19856,N_19794);
nor U20250 (N_20250,N_20190,N_20101);
xor U20251 (N_20251,N_20108,N_20112);
xnor U20252 (N_20252,N_20110,N_20193);
and U20253 (N_20253,N_20118,N_20143);
or U20254 (N_20254,N_20185,N_20123);
nor U20255 (N_20255,N_20030,N_20078);
nand U20256 (N_20256,N_20107,N_20121);
nor U20257 (N_20257,N_20095,N_20046);
xor U20258 (N_20258,N_20072,N_20081);
nand U20259 (N_20259,N_20167,N_20200);
xor U20260 (N_20260,N_20234,N_20160);
and U20261 (N_20261,N_20214,N_20127);
xor U20262 (N_20262,N_20189,N_20005);
and U20263 (N_20263,N_20013,N_20048);
nand U20264 (N_20264,N_20082,N_20119);
or U20265 (N_20265,N_20087,N_20028);
xnor U20266 (N_20266,N_20057,N_20139);
and U20267 (N_20267,N_20241,N_20128);
and U20268 (N_20268,N_20137,N_20243);
or U20269 (N_20269,N_20052,N_20187);
nand U20270 (N_20270,N_20237,N_20212);
nor U20271 (N_20271,N_20098,N_20058);
nor U20272 (N_20272,N_20073,N_20181);
or U20273 (N_20273,N_20135,N_20033);
nand U20274 (N_20274,N_20104,N_20047);
nor U20275 (N_20275,N_20061,N_20197);
and U20276 (N_20276,N_20019,N_20036);
xnor U20277 (N_20277,N_20111,N_20147);
xor U20278 (N_20278,N_20201,N_20177);
xnor U20279 (N_20279,N_20029,N_20122);
or U20280 (N_20280,N_20242,N_20062);
and U20281 (N_20281,N_20230,N_20192);
nor U20282 (N_20282,N_20218,N_20238);
nand U20283 (N_20283,N_20198,N_20209);
nor U20284 (N_20284,N_20141,N_20161);
and U20285 (N_20285,N_20159,N_20231);
and U20286 (N_20286,N_20207,N_20051);
nor U20287 (N_20287,N_20109,N_20210);
or U20288 (N_20288,N_20102,N_20085);
xor U20289 (N_20289,N_20050,N_20220);
xor U20290 (N_20290,N_20076,N_20232);
or U20291 (N_20291,N_20038,N_20186);
nand U20292 (N_20292,N_20031,N_20064);
nor U20293 (N_20293,N_20136,N_20114);
and U20294 (N_20294,N_20016,N_20074);
xor U20295 (N_20295,N_20023,N_20024);
nor U20296 (N_20296,N_20096,N_20115);
nand U20297 (N_20297,N_20091,N_20065);
or U20298 (N_20298,N_20228,N_20166);
xor U20299 (N_20299,N_20199,N_20157);
nor U20300 (N_20300,N_20203,N_20168);
and U20301 (N_20301,N_20195,N_20227);
xor U20302 (N_20302,N_20066,N_20131);
or U20303 (N_20303,N_20151,N_20054);
and U20304 (N_20304,N_20240,N_20133);
nor U20305 (N_20305,N_20215,N_20229);
and U20306 (N_20306,N_20248,N_20010);
or U20307 (N_20307,N_20097,N_20247);
or U20308 (N_20308,N_20043,N_20080);
nor U20309 (N_20309,N_20090,N_20044);
and U20310 (N_20310,N_20027,N_20129);
xor U20311 (N_20311,N_20079,N_20134);
xnor U20312 (N_20312,N_20003,N_20130);
or U20313 (N_20313,N_20146,N_20035);
or U20314 (N_20314,N_20142,N_20236);
xnor U20315 (N_20315,N_20086,N_20083);
nor U20316 (N_20316,N_20056,N_20100);
nand U20317 (N_20317,N_20249,N_20158);
nand U20318 (N_20318,N_20042,N_20165);
and U20319 (N_20319,N_20103,N_20155);
nand U20320 (N_20320,N_20017,N_20049);
nand U20321 (N_20321,N_20001,N_20032);
or U20322 (N_20322,N_20223,N_20244);
or U20323 (N_20323,N_20002,N_20009);
nor U20324 (N_20324,N_20026,N_20060);
and U20325 (N_20325,N_20020,N_20055);
and U20326 (N_20326,N_20180,N_20117);
or U20327 (N_20327,N_20039,N_20217);
nor U20328 (N_20328,N_20233,N_20040);
or U20329 (N_20329,N_20124,N_20171);
xnor U20330 (N_20330,N_20182,N_20106);
nor U20331 (N_20331,N_20041,N_20053);
nand U20332 (N_20332,N_20144,N_20089);
or U20333 (N_20333,N_20093,N_20196);
and U20334 (N_20334,N_20116,N_20145);
xor U20335 (N_20335,N_20148,N_20125);
nand U20336 (N_20336,N_20173,N_20140);
xnor U20337 (N_20337,N_20191,N_20163);
nand U20338 (N_20338,N_20170,N_20169);
nor U20339 (N_20339,N_20034,N_20211);
and U20340 (N_20340,N_20164,N_20092);
xor U20341 (N_20341,N_20172,N_20045);
or U20342 (N_20342,N_20011,N_20178);
nor U20343 (N_20343,N_20088,N_20126);
nor U20344 (N_20344,N_20183,N_20179);
or U20345 (N_20345,N_20099,N_20120);
nand U20346 (N_20346,N_20012,N_20156);
or U20347 (N_20347,N_20007,N_20004);
xor U20348 (N_20348,N_20015,N_20077);
and U20349 (N_20349,N_20239,N_20037);
and U20350 (N_20350,N_20213,N_20174);
nand U20351 (N_20351,N_20084,N_20067);
and U20352 (N_20352,N_20021,N_20245);
and U20353 (N_20353,N_20224,N_20188);
xor U20354 (N_20354,N_20000,N_20132);
nand U20355 (N_20355,N_20226,N_20205);
xor U20356 (N_20356,N_20194,N_20216);
and U20357 (N_20357,N_20008,N_20105);
xnor U20358 (N_20358,N_20221,N_20113);
nand U20359 (N_20359,N_20063,N_20153);
and U20360 (N_20360,N_20075,N_20025);
and U20361 (N_20361,N_20235,N_20149);
xor U20362 (N_20362,N_20152,N_20225);
nand U20363 (N_20363,N_20246,N_20059);
or U20364 (N_20364,N_20094,N_20138);
or U20365 (N_20365,N_20069,N_20006);
xor U20366 (N_20366,N_20070,N_20202);
and U20367 (N_20367,N_20071,N_20014);
xnor U20368 (N_20368,N_20154,N_20204);
xor U20369 (N_20369,N_20162,N_20222);
or U20370 (N_20370,N_20184,N_20150);
xnor U20371 (N_20371,N_20208,N_20206);
xor U20372 (N_20372,N_20175,N_20022);
nand U20373 (N_20373,N_20219,N_20018);
and U20374 (N_20374,N_20176,N_20068);
nand U20375 (N_20375,N_20169,N_20124);
or U20376 (N_20376,N_20002,N_20087);
nand U20377 (N_20377,N_20113,N_20076);
xnor U20378 (N_20378,N_20182,N_20058);
nor U20379 (N_20379,N_20240,N_20039);
or U20380 (N_20380,N_20079,N_20210);
xor U20381 (N_20381,N_20096,N_20243);
nor U20382 (N_20382,N_20146,N_20118);
xnor U20383 (N_20383,N_20150,N_20231);
and U20384 (N_20384,N_20117,N_20034);
or U20385 (N_20385,N_20113,N_20093);
xor U20386 (N_20386,N_20009,N_20078);
nand U20387 (N_20387,N_20192,N_20166);
and U20388 (N_20388,N_20035,N_20137);
nand U20389 (N_20389,N_20003,N_20197);
nor U20390 (N_20390,N_20184,N_20050);
or U20391 (N_20391,N_20065,N_20202);
xnor U20392 (N_20392,N_20056,N_20081);
xnor U20393 (N_20393,N_20050,N_20130);
nor U20394 (N_20394,N_20014,N_20183);
xor U20395 (N_20395,N_20197,N_20052);
nand U20396 (N_20396,N_20111,N_20184);
nand U20397 (N_20397,N_20099,N_20174);
nor U20398 (N_20398,N_20155,N_20064);
xor U20399 (N_20399,N_20050,N_20213);
xor U20400 (N_20400,N_20041,N_20167);
nor U20401 (N_20401,N_20112,N_20002);
xor U20402 (N_20402,N_20168,N_20143);
xnor U20403 (N_20403,N_20006,N_20191);
xnor U20404 (N_20404,N_20059,N_20014);
nor U20405 (N_20405,N_20241,N_20082);
nand U20406 (N_20406,N_20167,N_20168);
and U20407 (N_20407,N_20043,N_20175);
nor U20408 (N_20408,N_20191,N_20112);
and U20409 (N_20409,N_20084,N_20093);
nor U20410 (N_20410,N_20157,N_20129);
and U20411 (N_20411,N_20035,N_20015);
xnor U20412 (N_20412,N_20018,N_20013);
xnor U20413 (N_20413,N_20231,N_20126);
xor U20414 (N_20414,N_20249,N_20128);
and U20415 (N_20415,N_20130,N_20024);
nand U20416 (N_20416,N_20013,N_20215);
xor U20417 (N_20417,N_20072,N_20019);
nand U20418 (N_20418,N_20131,N_20107);
or U20419 (N_20419,N_20129,N_20140);
nor U20420 (N_20420,N_20204,N_20110);
nor U20421 (N_20421,N_20081,N_20058);
or U20422 (N_20422,N_20232,N_20067);
nor U20423 (N_20423,N_20117,N_20244);
xor U20424 (N_20424,N_20142,N_20226);
or U20425 (N_20425,N_20141,N_20055);
xor U20426 (N_20426,N_20237,N_20102);
nand U20427 (N_20427,N_20118,N_20026);
nand U20428 (N_20428,N_20046,N_20003);
nor U20429 (N_20429,N_20036,N_20067);
xor U20430 (N_20430,N_20186,N_20168);
nor U20431 (N_20431,N_20171,N_20017);
nand U20432 (N_20432,N_20176,N_20134);
nor U20433 (N_20433,N_20128,N_20005);
nor U20434 (N_20434,N_20029,N_20012);
nand U20435 (N_20435,N_20244,N_20022);
xor U20436 (N_20436,N_20073,N_20041);
xnor U20437 (N_20437,N_20229,N_20015);
nor U20438 (N_20438,N_20219,N_20061);
and U20439 (N_20439,N_20101,N_20044);
xnor U20440 (N_20440,N_20062,N_20041);
nand U20441 (N_20441,N_20063,N_20060);
and U20442 (N_20442,N_20238,N_20058);
nor U20443 (N_20443,N_20137,N_20177);
or U20444 (N_20444,N_20054,N_20069);
xor U20445 (N_20445,N_20241,N_20103);
and U20446 (N_20446,N_20023,N_20053);
nor U20447 (N_20447,N_20168,N_20099);
nand U20448 (N_20448,N_20041,N_20028);
nor U20449 (N_20449,N_20122,N_20200);
and U20450 (N_20450,N_20097,N_20241);
nand U20451 (N_20451,N_20181,N_20071);
and U20452 (N_20452,N_20223,N_20130);
and U20453 (N_20453,N_20190,N_20025);
nor U20454 (N_20454,N_20071,N_20150);
and U20455 (N_20455,N_20032,N_20179);
nand U20456 (N_20456,N_20039,N_20106);
and U20457 (N_20457,N_20040,N_20061);
or U20458 (N_20458,N_20045,N_20052);
nand U20459 (N_20459,N_20146,N_20202);
and U20460 (N_20460,N_20063,N_20140);
xnor U20461 (N_20461,N_20061,N_20160);
nor U20462 (N_20462,N_20044,N_20174);
and U20463 (N_20463,N_20019,N_20224);
nand U20464 (N_20464,N_20197,N_20178);
or U20465 (N_20465,N_20224,N_20067);
or U20466 (N_20466,N_20023,N_20225);
nor U20467 (N_20467,N_20108,N_20145);
or U20468 (N_20468,N_20010,N_20071);
and U20469 (N_20469,N_20078,N_20019);
nand U20470 (N_20470,N_20133,N_20244);
xnor U20471 (N_20471,N_20077,N_20031);
or U20472 (N_20472,N_20133,N_20017);
and U20473 (N_20473,N_20007,N_20208);
or U20474 (N_20474,N_20095,N_20111);
nor U20475 (N_20475,N_20074,N_20237);
nor U20476 (N_20476,N_20176,N_20168);
and U20477 (N_20477,N_20135,N_20220);
or U20478 (N_20478,N_20145,N_20156);
or U20479 (N_20479,N_20203,N_20211);
or U20480 (N_20480,N_20043,N_20161);
and U20481 (N_20481,N_20203,N_20183);
nand U20482 (N_20482,N_20135,N_20090);
or U20483 (N_20483,N_20229,N_20186);
xor U20484 (N_20484,N_20125,N_20026);
xnor U20485 (N_20485,N_20039,N_20139);
or U20486 (N_20486,N_20035,N_20028);
xor U20487 (N_20487,N_20048,N_20219);
xor U20488 (N_20488,N_20163,N_20182);
nor U20489 (N_20489,N_20058,N_20078);
xnor U20490 (N_20490,N_20088,N_20080);
nor U20491 (N_20491,N_20120,N_20187);
nor U20492 (N_20492,N_20138,N_20190);
nand U20493 (N_20493,N_20110,N_20059);
and U20494 (N_20494,N_20052,N_20162);
or U20495 (N_20495,N_20245,N_20200);
or U20496 (N_20496,N_20157,N_20118);
nand U20497 (N_20497,N_20162,N_20205);
or U20498 (N_20498,N_20124,N_20095);
xor U20499 (N_20499,N_20002,N_20076);
or U20500 (N_20500,N_20370,N_20382);
and U20501 (N_20501,N_20415,N_20300);
and U20502 (N_20502,N_20290,N_20354);
nor U20503 (N_20503,N_20473,N_20389);
and U20504 (N_20504,N_20417,N_20289);
nand U20505 (N_20505,N_20455,N_20485);
and U20506 (N_20506,N_20264,N_20279);
nor U20507 (N_20507,N_20378,N_20282);
xor U20508 (N_20508,N_20348,N_20428);
or U20509 (N_20509,N_20498,N_20325);
or U20510 (N_20510,N_20291,N_20489);
nand U20511 (N_20511,N_20438,N_20288);
xor U20512 (N_20512,N_20269,N_20471);
xor U20513 (N_20513,N_20345,N_20446);
or U20514 (N_20514,N_20475,N_20443);
nand U20515 (N_20515,N_20301,N_20297);
nor U20516 (N_20516,N_20349,N_20412);
nand U20517 (N_20517,N_20459,N_20369);
nor U20518 (N_20518,N_20283,N_20402);
nor U20519 (N_20519,N_20319,N_20356);
and U20520 (N_20520,N_20333,N_20299);
or U20521 (N_20521,N_20364,N_20405);
and U20522 (N_20522,N_20421,N_20419);
or U20523 (N_20523,N_20451,N_20445);
and U20524 (N_20524,N_20447,N_20263);
and U20525 (N_20525,N_20461,N_20329);
and U20526 (N_20526,N_20454,N_20314);
and U20527 (N_20527,N_20499,N_20380);
xnor U20528 (N_20528,N_20358,N_20462);
xor U20529 (N_20529,N_20448,N_20432);
and U20530 (N_20530,N_20406,N_20334);
nand U20531 (N_20531,N_20361,N_20425);
nand U20532 (N_20532,N_20388,N_20366);
nor U20533 (N_20533,N_20497,N_20395);
and U20534 (N_20534,N_20278,N_20324);
nor U20535 (N_20535,N_20496,N_20396);
and U20536 (N_20536,N_20467,N_20427);
xor U20537 (N_20537,N_20352,N_20465);
xnor U20538 (N_20538,N_20260,N_20373);
and U20539 (N_20539,N_20304,N_20483);
and U20540 (N_20540,N_20296,N_20371);
nor U20541 (N_20541,N_20478,N_20423);
xnor U20542 (N_20542,N_20433,N_20346);
nand U20543 (N_20543,N_20275,N_20408);
nor U20544 (N_20544,N_20397,N_20258);
nand U20545 (N_20545,N_20326,N_20318);
xor U20546 (N_20546,N_20259,N_20399);
and U20547 (N_20547,N_20312,N_20424);
and U20548 (N_20548,N_20426,N_20359);
nor U20549 (N_20549,N_20456,N_20468);
nand U20550 (N_20550,N_20305,N_20458);
xnor U20551 (N_20551,N_20347,N_20390);
nand U20552 (N_20552,N_20479,N_20482);
nor U20553 (N_20553,N_20442,N_20310);
or U20554 (N_20554,N_20295,N_20376);
or U20555 (N_20555,N_20480,N_20267);
xor U20556 (N_20556,N_20268,N_20493);
xor U20557 (N_20557,N_20253,N_20271);
nand U20558 (N_20558,N_20315,N_20306);
or U20559 (N_20559,N_20252,N_20327);
nor U20560 (N_20560,N_20463,N_20335);
nor U20561 (N_20561,N_20464,N_20392);
and U20562 (N_20562,N_20466,N_20407);
xnor U20563 (N_20563,N_20339,N_20449);
xor U20564 (N_20564,N_20416,N_20492);
and U20565 (N_20565,N_20411,N_20435);
nand U20566 (N_20566,N_20377,N_20383);
and U20567 (N_20567,N_20313,N_20284);
nor U20568 (N_20568,N_20418,N_20307);
nand U20569 (N_20569,N_20453,N_20470);
nand U20570 (N_20570,N_20460,N_20484);
and U20571 (N_20571,N_20394,N_20273);
nand U20572 (N_20572,N_20431,N_20270);
nand U20573 (N_20573,N_20337,N_20422);
nor U20574 (N_20574,N_20420,N_20342);
xor U20575 (N_20575,N_20262,N_20294);
xor U20576 (N_20576,N_20266,N_20401);
nand U20577 (N_20577,N_20477,N_20495);
nor U20578 (N_20578,N_20277,N_20320);
or U20579 (N_20579,N_20298,N_20437);
and U20580 (N_20580,N_20257,N_20341);
xor U20581 (N_20581,N_20374,N_20434);
xnor U20582 (N_20582,N_20350,N_20436);
nand U20583 (N_20583,N_20343,N_20398);
nand U20584 (N_20584,N_20487,N_20311);
nand U20585 (N_20585,N_20292,N_20410);
or U20586 (N_20586,N_20256,N_20250);
xnor U20587 (N_20587,N_20365,N_20452);
xor U20588 (N_20588,N_20323,N_20387);
xor U20589 (N_20589,N_20385,N_20280);
or U20590 (N_20590,N_20251,N_20386);
nand U20591 (N_20591,N_20363,N_20486);
nor U20592 (N_20592,N_20276,N_20285);
xnor U20593 (N_20593,N_20391,N_20302);
or U20594 (N_20594,N_20322,N_20360);
xnor U20595 (N_20595,N_20265,N_20404);
xor U20596 (N_20596,N_20254,N_20481);
nand U20597 (N_20597,N_20472,N_20457);
or U20598 (N_20598,N_20393,N_20440);
and U20599 (N_20599,N_20286,N_20336);
nand U20600 (N_20600,N_20309,N_20272);
nor U20601 (N_20601,N_20429,N_20317);
and U20602 (N_20602,N_20450,N_20355);
nand U20603 (N_20603,N_20274,N_20403);
nand U20604 (N_20604,N_20439,N_20344);
xnor U20605 (N_20605,N_20375,N_20474);
and U20606 (N_20606,N_20281,N_20353);
or U20607 (N_20607,N_20357,N_20321);
xor U20608 (N_20608,N_20367,N_20381);
nor U20609 (N_20609,N_20490,N_20351);
xnor U20610 (N_20610,N_20316,N_20441);
and U20611 (N_20611,N_20413,N_20409);
xor U20612 (N_20612,N_20414,N_20400);
xor U20613 (N_20613,N_20255,N_20379);
nand U20614 (N_20614,N_20384,N_20330);
nor U20615 (N_20615,N_20340,N_20372);
nor U20616 (N_20616,N_20368,N_20328);
xnor U20617 (N_20617,N_20331,N_20308);
or U20618 (N_20618,N_20332,N_20287);
or U20619 (N_20619,N_20261,N_20430);
or U20620 (N_20620,N_20476,N_20303);
or U20621 (N_20621,N_20469,N_20444);
xnor U20622 (N_20622,N_20488,N_20338);
and U20623 (N_20623,N_20293,N_20491);
nand U20624 (N_20624,N_20362,N_20494);
xnor U20625 (N_20625,N_20365,N_20305);
or U20626 (N_20626,N_20326,N_20467);
xor U20627 (N_20627,N_20429,N_20444);
or U20628 (N_20628,N_20489,N_20464);
or U20629 (N_20629,N_20346,N_20372);
and U20630 (N_20630,N_20487,N_20454);
and U20631 (N_20631,N_20381,N_20346);
xnor U20632 (N_20632,N_20357,N_20367);
or U20633 (N_20633,N_20440,N_20288);
and U20634 (N_20634,N_20481,N_20349);
and U20635 (N_20635,N_20422,N_20312);
or U20636 (N_20636,N_20356,N_20496);
or U20637 (N_20637,N_20492,N_20428);
and U20638 (N_20638,N_20318,N_20483);
xor U20639 (N_20639,N_20296,N_20492);
or U20640 (N_20640,N_20296,N_20281);
nand U20641 (N_20641,N_20426,N_20441);
nor U20642 (N_20642,N_20391,N_20329);
and U20643 (N_20643,N_20260,N_20345);
nand U20644 (N_20644,N_20473,N_20308);
nand U20645 (N_20645,N_20338,N_20329);
or U20646 (N_20646,N_20294,N_20442);
xor U20647 (N_20647,N_20372,N_20308);
nor U20648 (N_20648,N_20492,N_20381);
xor U20649 (N_20649,N_20275,N_20480);
xor U20650 (N_20650,N_20456,N_20408);
nand U20651 (N_20651,N_20388,N_20424);
xnor U20652 (N_20652,N_20283,N_20446);
or U20653 (N_20653,N_20402,N_20270);
and U20654 (N_20654,N_20364,N_20338);
and U20655 (N_20655,N_20329,N_20353);
and U20656 (N_20656,N_20488,N_20353);
xor U20657 (N_20657,N_20453,N_20495);
or U20658 (N_20658,N_20340,N_20414);
or U20659 (N_20659,N_20398,N_20366);
and U20660 (N_20660,N_20350,N_20467);
nand U20661 (N_20661,N_20309,N_20409);
xnor U20662 (N_20662,N_20456,N_20294);
xor U20663 (N_20663,N_20466,N_20271);
nor U20664 (N_20664,N_20295,N_20438);
or U20665 (N_20665,N_20409,N_20391);
or U20666 (N_20666,N_20463,N_20445);
nor U20667 (N_20667,N_20377,N_20360);
and U20668 (N_20668,N_20389,N_20290);
nand U20669 (N_20669,N_20429,N_20376);
and U20670 (N_20670,N_20425,N_20496);
or U20671 (N_20671,N_20314,N_20436);
nor U20672 (N_20672,N_20480,N_20498);
nor U20673 (N_20673,N_20481,N_20407);
and U20674 (N_20674,N_20378,N_20310);
nand U20675 (N_20675,N_20409,N_20456);
and U20676 (N_20676,N_20464,N_20290);
or U20677 (N_20677,N_20329,N_20497);
and U20678 (N_20678,N_20290,N_20498);
and U20679 (N_20679,N_20296,N_20372);
and U20680 (N_20680,N_20252,N_20496);
nand U20681 (N_20681,N_20310,N_20451);
xnor U20682 (N_20682,N_20471,N_20330);
xor U20683 (N_20683,N_20351,N_20318);
nor U20684 (N_20684,N_20278,N_20496);
and U20685 (N_20685,N_20472,N_20470);
nor U20686 (N_20686,N_20392,N_20260);
nand U20687 (N_20687,N_20493,N_20255);
nor U20688 (N_20688,N_20313,N_20250);
and U20689 (N_20689,N_20301,N_20296);
nand U20690 (N_20690,N_20396,N_20495);
xor U20691 (N_20691,N_20275,N_20499);
nand U20692 (N_20692,N_20480,N_20325);
or U20693 (N_20693,N_20382,N_20440);
or U20694 (N_20694,N_20333,N_20443);
xor U20695 (N_20695,N_20485,N_20374);
nor U20696 (N_20696,N_20354,N_20357);
xor U20697 (N_20697,N_20412,N_20450);
nor U20698 (N_20698,N_20295,N_20469);
nand U20699 (N_20699,N_20300,N_20465);
nor U20700 (N_20700,N_20276,N_20310);
xnor U20701 (N_20701,N_20451,N_20304);
or U20702 (N_20702,N_20461,N_20456);
or U20703 (N_20703,N_20352,N_20321);
xor U20704 (N_20704,N_20404,N_20375);
and U20705 (N_20705,N_20280,N_20381);
xnor U20706 (N_20706,N_20255,N_20495);
and U20707 (N_20707,N_20432,N_20431);
and U20708 (N_20708,N_20264,N_20453);
and U20709 (N_20709,N_20281,N_20264);
xnor U20710 (N_20710,N_20493,N_20318);
and U20711 (N_20711,N_20329,N_20487);
and U20712 (N_20712,N_20269,N_20480);
and U20713 (N_20713,N_20259,N_20302);
xor U20714 (N_20714,N_20309,N_20485);
or U20715 (N_20715,N_20477,N_20273);
nand U20716 (N_20716,N_20400,N_20434);
nand U20717 (N_20717,N_20409,N_20269);
nor U20718 (N_20718,N_20271,N_20377);
nand U20719 (N_20719,N_20458,N_20389);
or U20720 (N_20720,N_20254,N_20329);
xor U20721 (N_20721,N_20489,N_20258);
xnor U20722 (N_20722,N_20362,N_20283);
nand U20723 (N_20723,N_20263,N_20349);
xor U20724 (N_20724,N_20363,N_20258);
nand U20725 (N_20725,N_20426,N_20389);
xor U20726 (N_20726,N_20472,N_20256);
or U20727 (N_20727,N_20395,N_20375);
nand U20728 (N_20728,N_20265,N_20253);
xnor U20729 (N_20729,N_20436,N_20419);
nor U20730 (N_20730,N_20471,N_20336);
xnor U20731 (N_20731,N_20300,N_20279);
nand U20732 (N_20732,N_20432,N_20323);
and U20733 (N_20733,N_20427,N_20375);
and U20734 (N_20734,N_20293,N_20396);
or U20735 (N_20735,N_20321,N_20379);
xor U20736 (N_20736,N_20324,N_20413);
and U20737 (N_20737,N_20344,N_20270);
nand U20738 (N_20738,N_20360,N_20253);
or U20739 (N_20739,N_20265,N_20382);
xnor U20740 (N_20740,N_20278,N_20266);
or U20741 (N_20741,N_20321,N_20351);
nor U20742 (N_20742,N_20462,N_20383);
nor U20743 (N_20743,N_20337,N_20276);
nor U20744 (N_20744,N_20322,N_20484);
nand U20745 (N_20745,N_20332,N_20293);
nand U20746 (N_20746,N_20417,N_20374);
nor U20747 (N_20747,N_20426,N_20386);
nand U20748 (N_20748,N_20296,N_20345);
nand U20749 (N_20749,N_20265,N_20424);
nand U20750 (N_20750,N_20613,N_20599);
nand U20751 (N_20751,N_20509,N_20527);
and U20752 (N_20752,N_20739,N_20589);
xnor U20753 (N_20753,N_20683,N_20504);
nand U20754 (N_20754,N_20520,N_20611);
xnor U20755 (N_20755,N_20673,N_20670);
nor U20756 (N_20756,N_20582,N_20692);
nand U20757 (N_20757,N_20579,N_20648);
nand U20758 (N_20758,N_20603,N_20587);
and U20759 (N_20759,N_20634,N_20747);
nand U20760 (N_20760,N_20702,N_20627);
and U20761 (N_20761,N_20662,N_20538);
and U20762 (N_20762,N_20618,N_20568);
nand U20763 (N_20763,N_20560,N_20617);
xnor U20764 (N_20764,N_20506,N_20633);
nor U20765 (N_20765,N_20734,N_20635);
xnor U20766 (N_20766,N_20594,N_20588);
and U20767 (N_20767,N_20686,N_20596);
nor U20768 (N_20768,N_20566,N_20614);
xor U20769 (N_20769,N_20745,N_20525);
and U20770 (N_20770,N_20555,N_20671);
or U20771 (N_20771,N_20748,N_20646);
and U20772 (N_20772,N_20665,N_20743);
or U20773 (N_20773,N_20553,N_20619);
xor U20774 (N_20774,N_20605,N_20681);
nand U20775 (N_20775,N_20580,N_20517);
nand U20776 (N_20776,N_20700,N_20721);
nor U20777 (N_20777,N_20616,N_20650);
or U20778 (N_20778,N_20740,N_20667);
nand U20779 (N_20779,N_20602,N_20659);
and U20780 (N_20780,N_20562,N_20699);
and U20781 (N_20781,N_20717,N_20746);
and U20782 (N_20782,N_20511,N_20530);
and U20783 (N_20783,N_20724,N_20624);
or U20784 (N_20784,N_20676,N_20674);
xnor U20785 (N_20785,N_20607,N_20679);
or U20786 (N_20786,N_20719,N_20507);
xnor U20787 (N_20787,N_20685,N_20675);
xnor U20788 (N_20788,N_20666,N_20708);
xor U20789 (N_20789,N_20711,N_20501);
nand U20790 (N_20790,N_20541,N_20533);
nor U20791 (N_20791,N_20696,N_20690);
and U20792 (N_20792,N_20678,N_20658);
nor U20793 (N_20793,N_20653,N_20652);
nand U20794 (N_20794,N_20697,N_20581);
and U20795 (N_20795,N_20592,N_20590);
or U20796 (N_20796,N_20638,N_20502);
or U20797 (N_20797,N_20691,N_20632);
and U20798 (N_20798,N_20548,N_20707);
and U20799 (N_20799,N_20519,N_20521);
and U20800 (N_20800,N_20625,N_20636);
nor U20801 (N_20801,N_20537,N_20500);
xnor U20802 (N_20802,N_20585,N_20578);
nor U20803 (N_20803,N_20583,N_20641);
or U20804 (N_20804,N_20556,N_20606);
nor U20805 (N_20805,N_20680,N_20749);
xor U20806 (N_20806,N_20565,N_20733);
nor U20807 (N_20807,N_20515,N_20698);
nand U20808 (N_20808,N_20570,N_20727);
nor U20809 (N_20809,N_20516,N_20712);
nor U20810 (N_20810,N_20723,N_20647);
and U20811 (N_20811,N_20549,N_20532);
nor U20812 (N_20812,N_20584,N_20572);
nand U20813 (N_20813,N_20522,N_20535);
nor U20814 (N_20814,N_20701,N_20639);
or U20815 (N_20815,N_20654,N_20561);
xor U20816 (N_20816,N_20615,N_20689);
or U20817 (N_20817,N_20655,N_20669);
nor U20818 (N_20818,N_20503,N_20524);
and U20819 (N_20819,N_20718,N_20593);
xnor U20820 (N_20820,N_20597,N_20640);
nand U20821 (N_20821,N_20591,N_20598);
nand U20822 (N_20822,N_20694,N_20629);
nand U20823 (N_20823,N_20609,N_20608);
and U20824 (N_20824,N_20687,N_20513);
xnor U20825 (N_20825,N_20703,N_20672);
xor U20826 (N_20826,N_20728,N_20643);
nor U20827 (N_20827,N_20656,N_20558);
nor U20828 (N_20828,N_20577,N_20518);
and U20829 (N_20829,N_20628,N_20545);
nand U20830 (N_20830,N_20738,N_20631);
and U20831 (N_20831,N_20661,N_20512);
nor U20832 (N_20832,N_20709,N_20531);
and U20833 (N_20833,N_20729,N_20612);
and U20834 (N_20834,N_20663,N_20651);
xor U20835 (N_20835,N_20576,N_20715);
nand U20836 (N_20836,N_20564,N_20610);
xor U20837 (N_20837,N_20540,N_20505);
and U20838 (N_20838,N_20604,N_20668);
nand U20839 (N_20839,N_20664,N_20621);
nor U20840 (N_20840,N_20704,N_20737);
and U20841 (N_20841,N_20574,N_20657);
xor U20842 (N_20842,N_20725,N_20735);
xnor U20843 (N_20843,N_20526,N_20626);
or U20844 (N_20844,N_20573,N_20623);
or U20845 (N_20845,N_20543,N_20550);
and U20846 (N_20846,N_20741,N_20534);
xnor U20847 (N_20847,N_20529,N_20544);
and U20848 (N_20848,N_20567,N_20677);
xor U20849 (N_20849,N_20714,N_20551);
xnor U20850 (N_20850,N_20559,N_20706);
nor U20851 (N_20851,N_20528,N_20688);
or U20852 (N_20852,N_20736,N_20637);
nor U20853 (N_20853,N_20682,N_20547);
xnor U20854 (N_20854,N_20710,N_20552);
or U20855 (N_20855,N_20620,N_20630);
and U20856 (N_20856,N_20649,N_20595);
xnor U20857 (N_20857,N_20726,N_20622);
nand U20858 (N_20858,N_20684,N_20536);
nor U20859 (N_20859,N_20732,N_20705);
or U20860 (N_20860,N_20716,N_20563);
xor U20861 (N_20861,N_20660,N_20644);
nor U20862 (N_20862,N_20693,N_20523);
nand U20863 (N_20863,N_20730,N_20557);
nor U20864 (N_20864,N_20510,N_20695);
or U20865 (N_20865,N_20546,N_20742);
xnor U20866 (N_20866,N_20586,N_20539);
nand U20867 (N_20867,N_20514,N_20575);
nand U20868 (N_20868,N_20720,N_20722);
xnor U20869 (N_20869,N_20645,N_20554);
nor U20870 (N_20870,N_20571,N_20600);
nand U20871 (N_20871,N_20642,N_20731);
xnor U20872 (N_20872,N_20542,N_20744);
nor U20873 (N_20873,N_20713,N_20508);
nor U20874 (N_20874,N_20569,N_20601);
and U20875 (N_20875,N_20514,N_20650);
or U20876 (N_20876,N_20687,N_20500);
and U20877 (N_20877,N_20649,N_20535);
and U20878 (N_20878,N_20560,N_20641);
nor U20879 (N_20879,N_20617,N_20537);
xnor U20880 (N_20880,N_20717,N_20608);
nor U20881 (N_20881,N_20541,N_20642);
or U20882 (N_20882,N_20708,N_20576);
xnor U20883 (N_20883,N_20723,N_20725);
and U20884 (N_20884,N_20671,N_20678);
or U20885 (N_20885,N_20506,N_20704);
xnor U20886 (N_20886,N_20737,N_20582);
nand U20887 (N_20887,N_20562,N_20511);
nand U20888 (N_20888,N_20631,N_20616);
nand U20889 (N_20889,N_20682,N_20624);
and U20890 (N_20890,N_20722,N_20639);
nand U20891 (N_20891,N_20694,N_20729);
and U20892 (N_20892,N_20613,N_20619);
and U20893 (N_20893,N_20732,N_20591);
nand U20894 (N_20894,N_20704,N_20708);
nand U20895 (N_20895,N_20534,N_20587);
and U20896 (N_20896,N_20538,N_20507);
nor U20897 (N_20897,N_20568,N_20738);
and U20898 (N_20898,N_20718,N_20681);
nor U20899 (N_20899,N_20745,N_20567);
and U20900 (N_20900,N_20681,N_20648);
or U20901 (N_20901,N_20576,N_20609);
nor U20902 (N_20902,N_20674,N_20733);
or U20903 (N_20903,N_20680,N_20705);
or U20904 (N_20904,N_20578,N_20579);
nand U20905 (N_20905,N_20518,N_20741);
nor U20906 (N_20906,N_20610,N_20667);
and U20907 (N_20907,N_20533,N_20554);
and U20908 (N_20908,N_20648,N_20526);
and U20909 (N_20909,N_20600,N_20513);
xor U20910 (N_20910,N_20562,N_20596);
nor U20911 (N_20911,N_20525,N_20609);
nor U20912 (N_20912,N_20733,N_20668);
nand U20913 (N_20913,N_20501,N_20559);
or U20914 (N_20914,N_20595,N_20611);
nand U20915 (N_20915,N_20634,N_20609);
nor U20916 (N_20916,N_20716,N_20589);
or U20917 (N_20917,N_20733,N_20594);
nand U20918 (N_20918,N_20709,N_20626);
or U20919 (N_20919,N_20632,N_20701);
nand U20920 (N_20920,N_20573,N_20612);
nor U20921 (N_20921,N_20741,N_20717);
nand U20922 (N_20922,N_20545,N_20745);
or U20923 (N_20923,N_20588,N_20631);
nor U20924 (N_20924,N_20503,N_20570);
or U20925 (N_20925,N_20653,N_20590);
or U20926 (N_20926,N_20716,N_20641);
nor U20927 (N_20927,N_20677,N_20613);
nand U20928 (N_20928,N_20594,N_20586);
xnor U20929 (N_20929,N_20537,N_20561);
or U20930 (N_20930,N_20674,N_20522);
xnor U20931 (N_20931,N_20701,N_20531);
or U20932 (N_20932,N_20737,N_20547);
and U20933 (N_20933,N_20501,N_20624);
nand U20934 (N_20934,N_20595,N_20520);
nor U20935 (N_20935,N_20550,N_20687);
or U20936 (N_20936,N_20668,N_20545);
or U20937 (N_20937,N_20733,N_20642);
xnor U20938 (N_20938,N_20686,N_20703);
nor U20939 (N_20939,N_20615,N_20737);
and U20940 (N_20940,N_20674,N_20545);
nand U20941 (N_20941,N_20631,N_20578);
and U20942 (N_20942,N_20577,N_20708);
nand U20943 (N_20943,N_20710,N_20590);
and U20944 (N_20944,N_20554,N_20604);
or U20945 (N_20945,N_20543,N_20747);
or U20946 (N_20946,N_20722,N_20636);
or U20947 (N_20947,N_20700,N_20631);
or U20948 (N_20948,N_20620,N_20733);
or U20949 (N_20949,N_20542,N_20736);
xnor U20950 (N_20950,N_20696,N_20638);
nand U20951 (N_20951,N_20708,N_20723);
nor U20952 (N_20952,N_20555,N_20684);
xnor U20953 (N_20953,N_20516,N_20710);
or U20954 (N_20954,N_20641,N_20594);
nand U20955 (N_20955,N_20531,N_20577);
and U20956 (N_20956,N_20564,N_20648);
nor U20957 (N_20957,N_20578,N_20648);
xnor U20958 (N_20958,N_20639,N_20640);
and U20959 (N_20959,N_20687,N_20545);
and U20960 (N_20960,N_20625,N_20715);
xor U20961 (N_20961,N_20663,N_20549);
or U20962 (N_20962,N_20609,N_20642);
xnor U20963 (N_20963,N_20620,N_20553);
nand U20964 (N_20964,N_20502,N_20706);
or U20965 (N_20965,N_20538,N_20542);
or U20966 (N_20966,N_20657,N_20511);
and U20967 (N_20967,N_20513,N_20675);
xor U20968 (N_20968,N_20558,N_20702);
xor U20969 (N_20969,N_20574,N_20670);
nor U20970 (N_20970,N_20684,N_20622);
nor U20971 (N_20971,N_20667,N_20513);
nor U20972 (N_20972,N_20687,N_20625);
and U20973 (N_20973,N_20742,N_20551);
xor U20974 (N_20974,N_20530,N_20651);
and U20975 (N_20975,N_20573,N_20657);
or U20976 (N_20976,N_20722,N_20716);
nand U20977 (N_20977,N_20748,N_20731);
xnor U20978 (N_20978,N_20693,N_20697);
xor U20979 (N_20979,N_20642,N_20680);
nand U20980 (N_20980,N_20701,N_20608);
nor U20981 (N_20981,N_20626,N_20573);
and U20982 (N_20982,N_20747,N_20650);
xor U20983 (N_20983,N_20619,N_20555);
or U20984 (N_20984,N_20747,N_20737);
or U20985 (N_20985,N_20694,N_20547);
and U20986 (N_20986,N_20511,N_20672);
xor U20987 (N_20987,N_20640,N_20625);
or U20988 (N_20988,N_20552,N_20718);
or U20989 (N_20989,N_20532,N_20653);
and U20990 (N_20990,N_20562,N_20666);
or U20991 (N_20991,N_20571,N_20525);
and U20992 (N_20992,N_20524,N_20526);
xor U20993 (N_20993,N_20530,N_20508);
or U20994 (N_20994,N_20593,N_20676);
nor U20995 (N_20995,N_20597,N_20694);
xor U20996 (N_20996,N_20720,N_20506);
or U20997 (N_20997,N_20595,N_20686);
xnor U20998 (N_20998,N_20593,N_20566);
nor U20999 (N_20999,N_20508,N_20522);
and U21000 (N_21000,N_20805,N_20915);
nor U21001 (N_21001,N_20770,N_20870);
nor U21002 (N_21002,N_20971,N_20950);
xnor U21003 (N_21003,N_20964,N_20850);
nor U21004 (N_21004,N_20859,N_20757);
or U21005 (N_21005,N_20990,N_20780);
or U21006 (N_21006,N_20823,N_20980);
nand U21007 (N_21007,N_20777,N_20932);
nand U21008 (N_21008,N_20945,N_20752);
xor U21009 (N_21009,N_20843,N_20935);
nand U21010 (N_21010,N_20802,N_20769);
nand U21011 (N_21011,N_20953,N_20986);
or U21012 (N_21012,N_20985,N_20783);
nor U21013 (N_21013,N_20812,N_20886);
nor U21014 (N_21014,N_20889,N_20919);
and U21015 (N_21015,N_20988,N_20982);
xor U21016 (N_21016,N_20934,N_20911);
nor U21017 (N_21017,N_20961,N_20778);
xnor U21018 (N_21018,N_20775,N_20981);
nor U21019 (N_21019,N_20841,N_20910);
nor U21020 (N_21020,N_20872,N_20907);
xor U21021 (N_21021,N_20926,N_20967);
and U21022 (N_21022,N_20858,N_20943);
xnor U21023 (N_21023,N_20898,N_20972);
nor U21024 (N_21024,N_20913,N_20947);
xor U21025 (N_21025,N_20903,N_20811);
and U21026 (N_21026,N_20931,N_20874);
xnor U21027 (N_21027,N_20813,N_20867);
nand U21028 (N_21028,N_20974,N_20968);
nor U21029 (N_21029,N_20786,N_20925);
xor U21030 (N_21030,N_20834,N_20809);
or U21031 (N_21031,N_20948,N_20869);
and U21032 (N_21032,N_20938,N_20900);
xnor U21033 (N_21033,N_20865,N_20836);
nand U21034 (N_21034,N_20860,N_20999);
xnor U21035 (N_21035,N_20791,N_20766);
nor U21036 (N_21036,N_20877,N_20863);
or U21037 (N_21037,N_20929,N_20979);
or U21038 (N_21038,N_20973,N_20893);
nor U21039 (N_21039,N_20774,N_20866);
nor U21040 (N_21040,N_20820,N_20760);
xor U21041 (N_21041,N_20857,N_20958);
and U21042 (N_21042,N_20887,N_20906);
and U21043 (N_21043,N_20751,N_20914);
nand U21044 (N_21044,N_20785,N_20896);
or U21045 (N_21045,N_20796,N_20816);
and U21046 (N_21046,N_20789,N_20918);
nand U21047 (N_21047,N_20772,N_20917);
or U21048 (N_21048,N_20846,N_20838);
and U21049 (N_21049,N_20810,N_20835);
or U21050 (N_21050,N_20868,N_20821);
nor U21051 (N_21051,N_20797,N_20951);
nor U21052 (N_21052,N_20983,N_20801);
nor U21053 (N_21053,N_20781,N_20997);
xnor U21054 (N_21054,N_20878,N_20765);
xnor U21055 (N_21055,N_20849,N_20880);
and U21056 (N_21056,N_20848,N_20761);
xor U21057 (N_21057,N_20895,N_20794);
and U21058 (N_21058,N_20828,N_20939);
and U21059 (N_21059,N_20759,N_20976);
xnor U21060 (N_21060,N_20944,N_20930);
or U21061 (N_21061,N_20881,N_20936);
nand U21062 (N_21062,N_20842,N_20806);
and U21063 (N_21063,N_20832,N_20890);
nand U21064 (N_21064,N_20864,N_20755);
and U21065 (N_21065,N_20884,N_20819);
nand U21066 (N_21066,N_20800,N_20984);
nor U21067 (N_21067,N_20901,N_20963);
nand U21068 (N_21068,N_20764,N_20771);
and U21069 (N_21069,N_20818,N_20782);
and U21070 (N_21070,N_20827,N_20792);
nand U21071 (N_21071,N_20768,N_20798);
nand U21072 (N_21072,N_20891,N_20933);
nor U21073 (N_21073,N_20753,N_20856);
or U21074 (N_21074,N_20970,N_20804);
or U21075 (N_21075,N_20885,N_20949);
nand U21076 (N_21076,N_20837,N_20991);
xor U21077 (N_21077,N_20815,N_20839);
nand U21078 (N_21078,N_20784,N_20965);
and U21079 (N_21079,N_20787,N_20975);
xor U21080 (N_21080,N_20894,N_20923);
and U21081 (N_21081,N_20873,N_20799);
xor U21082 (N_21082,N_20960,N_20969);
nand U21083 (N_21083,N_20847,N_20854);
nand U21084 (N_21084,N_20904,N_20831);
xnor U21085 (N_21085,N_20956,N_20978);
and U21086 (N_21086,N_20952,N_20996);
nand U21087 (N_21087,N_20922,N_20807);
xnor U21088 (N_21088,N_20822,N_20845);
nor U21089 (N_21089,N_20920,N_20954);
nor U21090 (N_21090,N_20897,N_20927);
or U21091 (N_21091,N_20773,N_20962);
xor U21092 (N_21092,N_20908,N_20892);
and U21093 (N_21093,N_20795,N_20758);
and U21094 (N_21094,N_20957,N_20879);
or U21095 (N_21095,N_20928,N_20862);
and U21096 (N_21096,N_20750,N_20987);
nand U21097 (N_21097,N_20763,N_20829);
nand U21098 (N_21098,N_20909,N_20912);
and U21099 (N_21099,N_20808,N_20788);
and U21100 (N_21100,N_20994,N_20940);
nor U21101 (N_21101,N_20942,N_20756);
and U21102 (N_21102,N_20882,N_20883);
and U21103 (N_21103,N_20833,N_20955);
or U21104 (N_21104,N_20825,N_20851);
nand U21105 (N_21105,N_20817,N_20966);
xor U21106 (N_21106,N_20875,N_20992);
nor U21107 (N_21107,N_20853,N_20762);
and U21108 (N_21108,N_20824,N_20861);
and U21109 (N_21109,N_20754,N_20855);
nand U21110 (N_21110,N_20941,N_20767);
or U21111 (N_21111,N_20921,N_20840);
xor U21112 (N_21112,N_20779,N_20995);
xnor U21113 (N_21113,N_20902,N_20998);
nor U21114 (N_21114,N_20993,N_20790);
and U21115 (N_21115,N_20830,N_20871);
and U21116 (N_21116,N_20826,N_20899);
and U21117 (N_21117,N_20905,N_20793);
or U21118 (N_21118,N_20924,N_20989);
and U21119 (N_21119,N_20916,N_20876);
or U21120 (N_21120,N_20803,N_20946);
or U21121 (N_21121,N_20814,N_20977);
nor U21122 (N_21122,N_20776,N_20959);
nor U21123 (N_21123,N_20852,N_20937);
or U21124 (N_21124,N_20844,N_20888);
or U21125 (N_21125,N_20946,N_20899);
xor U21126 (N_21126,N_20853,N_20759);
nor U21127 (N_21127,N_20778,N_20868);
xor U21128 (N_21128,N_20786,N_20941);
xor U21129 (N_21129,N_20921,N_20862);
or U21130 (N_21130,N_20951,N_20814);
xor U21131 (N_21131,N_20834,N_20835);
or U21132 (N_21132,N_20823,N_20840);
nor U21133 (N_21133,N_20803,N_20756);
xor U21134 (N_21134,N_20943,N_20794);
xnor U21135 (N_21135,N_20991,N_20894);
and U21136 (N_21136,N_20759,N_20918);
or U21137 (N_21137,N_20911,N_20759);
or U21138 (N_21138,N_20883,N_20908);
xnor U21139 (N_21139,N_20960,N_20761);
or U21140 (N_21140,N_20969,N_20911);
xnor U21141 (N_21141,N_20957,N_20831);
xnor U21142 (N_21142,N_20917,N_20895);
xor U21143 (N_21143,N_20774,N_20906);
or U21144 (N_21144,N_20873,N_20839);
or U21145 (N_21145,N_20814,N_20842);
and U21146 (N_21146,N_20782,N_20963);
and U21147 (N_21147,N_20767,N_20763);
xor U21148 (N_21148,N_20772,N_20765);
nor U21149 (N_21149,N_20985,N_20999);
and U21150 (N_21150,N_20892,N_20929);
or U21151 (N_21151,N_20861,N_20963);
nor U21152 (N_21152,N_20920,N_20930);
nor U21153 (N_21153,N_20943,N_20962);
or U21154 (N_21154,N_20904,N_20826);
and U21155 (N_21155,N_20874,N_20762);
nor U21156 (N_21156,N_20754,N_20920);
and U21157 (N_21157,N_20833,N_20940);
nand U21158 (N_21158,N_20908,N_20957);
xnor U21159 (N_21159,N_20839,N_20798);
xor U21160 (N_21160,N_20900,N_20857);
nand U21161 (N_21161,N_20863,N_20848);
or U21162 (N_21162,N_20983,N_20818);
nand U21163 (N_21163,N_20972,N_20986);
and U21164 (N_21164,N_20841,N_20808);
nor U21165 (N_21165,N_20860,N_20784);
nand U21166 (N_21166,N_20751,N_20869);
xor U21167 (N_21167,N_20923,N_20790);
nor U21168 (N_21168,N_20900,N_20947);
nor U21169 (N_21169,N_20990,N_20993);
and U21170 (N_21170,N_20796,N_20856);
nor U21171 (N_21171,N_20779,N_20973);
nor U21172 (N_21172,N_20796,N_20903);
nand U21173 (N_21173,N_20926,N_20874);
and U21174 (N_21174,N_20870,N_20755);
and U21175 (N_21175,N_20828,N_20891);
nor U21176 (N_21176,N_20812,N_20935);
or U21177 (N_21177,N_20826,N_20979);
or U21178 (N_21178,N_20757,N_20831);
and U21179 (N_21179,N_20859,N_20944);
and U21180 (N_21180,N_20853,N_20754);
nand U21181 (N_21181,N_20930,N_20767);
xnor U21182 (N_21182,N_20774,N_20957);
xnor U21183 (N_21183,N_20822,N_20994);
nand U21184 (N_21184,N_20762,N_20834);
nand U21185 (N_21185,N_20978,N_20840);
or U21186 (N_21186,N_20891,N_20864);
xnor U21187 (N_21187,N_20914,N_20843);
nor U21188 (N_21188,N_20993,N_20984);
or U21189 (N_21189,N_20754,N_20973);
nor U21190 (N_21190,N_20783,N_20773);
nand U21191 (N_21191,N_20841,N_20882);
nand U21192 (N_21192,N_20917,N_20792);
nor U21193 (N_21193,N_20940,N_20846);
and U21194 (N_21194,N_20753,N_20751);
nand U21195 (N_21195,N_20769,N_20944);
nor U21196 (N_21196,N_20869,N_20930);
xor U21197 (N_21197,N_20971,N_20967);
or U21198 (N_21198,N_20990,N_20991);
xnor U21199 (N_21199,N_20896,N_20969);
and U21200 (N_21200,N_20963,N_20920);
or U21201 (N_21201,N_20902,N_20804);
xor U21202 (N_21202,N_20843,N_20857);
nor U21203 (N_21203,N_20866,N_20797);
nor U21204 (N_21204,N_20823,N_20847);
or U21205 (N_21205,N_20995,N_20880);
or U21206 (N_21206,N_20974,N_20845);
or U21207 (N_21207,N_20912,N_20757);
nor U21208 (N_21208,N_20763,N_20802);
nand U21209 (N_21209,N_20836,N_20881);
or U21210 (N_21210,N_20761,N_20825);
nor U21211 (N_21211,N_20763,N_20931);
and U21212 (N_21212,N_20889,N_20887);
or U21213 (N_21213,N_20784,N_20961);
nand U21214 (N_21214,N_20757,N_20901);
nand U21215 (N_21215,N_20930,N_20859);
and U21216 (N_21216,N_20815,N_20878);
xor U21217 (N_21217,N_20830,N_20915);
nor U21218 (N_21218,N_20938,N_20876);
xor U21219 (N_21219,N_20808,N_20843);
and U21220 (N_21220,N_20832,N_20860);
nor U21221 (N_21221,N_20858,N_20904);
xnor U21222 (N_21222,N_20846,N_20904);
or U21223 (N_21223,N_20985,N_20812);
and U21224 (N_21224,N_20916,N_20859);
xnor U21225 (N_21225,N_20824,N_20920);
and U21226 (N_21226,N_20930,N_20905);
and U21227 (N_21227,N_20822,N_20913);
nor U21228 (N_21228,N_20993,N_20877);
nand U21229 (N_21229,N_20941,N_20918);
nand U21230 (N_21230,N_20980,N_20754);
nor U21231 (N_21231,N_20923,N_20844);
xnor U21232 (N_21232,N_20842,N_20929);
and U21233 (N_21233,N_20907,N_20945);
nand U21234 (N_21234,N_20801,N_20762);
nor U21235 (N_21235,N_20867,N_20761);
nor U21236 (N_21236,N_20961,N_20791);
or U21237 (N_21237,N_20965,N_20842);
nand U21238 (N_21238,N_20933,N_20787);
or U21239 (N_21239,N_20761,N_20968);
xnor U21240 (N_21240,N_20977,N_20780);
xor U21241 (N_21241,N_20853,N_20780);
xor U21242 (N_21242,N_20954,N_20800);
nor U21243 (N_21243,N_20989,N_20855);
and U21244 (N_21244,N_20829,N_20824);
xor U21245 (N_21245,N_20896,N_20946);
xor U21246 (N_21246,N_20770,N_20764);
and U21247 (N_21247,N_20992,N_20782);
nor U21248 (N_21248,N_20965,N_20851);
xor U21249 (N_21249,N_20814,N_20762);
nor U21250 (N_21250,N_21104,N_21010);
nor U21251 (N_21251,N_21147,N_21075);
nor U21252 (N_21252,N_21043,N_21016);
or U21253 (N_21253,N_21093,N_21209);
or U21254 (N_21254,N_21241,N_21187);
and U21255 (N_21255,N_21127,N_21157);
or U21256 (N_21256,N_21155,N_21196);
or U21257 (N_21257,N_21109,N_21161);
nor U21258 (N_21258,N_21151,N_21116);
nand U21259 (N_21259,N_21235,N_21015);
or U21260 (N_21260,N_21133,N_21124);
and U21261 (N_21261,N_21059,N_21185);
or U21262 (N_21262,N_21199,N_21006);
nand U21263 (N_21263,N_21020,N_21173);
and U21264 (N_21264,N_21156,N_21142);
or U21265 (N_21265,N_21094,N_21089);
nand U21266 (N_21266,N_21129,N_21174);
xor U21267 (N_21267,N_21179,N_21125);
or U21268 (N_21268,N_21122,N_21097);
nor U21269 (N_21269,N_21188,N_21216);
nand U21270 (N_21270,N_21211,N_21207);
xor U21271 (N_21271,N_21165,N_21240);
nor U21272 (N_21272,N_21138,N_21163);
or U21273 (N_21273,N_21052,N_21014);
or U21274 (N_21274,N_21086,N_21153);
and U21275 (N_21275,N_21120,N_21001);
and U21276 (N_21276,N_21139,N_21198);
xor U21277 (N_21277,N_21191,N_21132);
and U21278 (N_21278,N_21072,N_21065);
xor U21279 (N_21279,N_21044,N_21041);
nand U21280 (N_21280,N_21146,N_21180);
and U21281 (N_21281,N_21242,N_21067);
nand U21282 (N_21282,N_21085,N_21215);
xnor U21283 (N_21283,N_21051,N_21115);
xor U21284 (N_21284,N_21219,N_21084);
and U21285 (N_21285,N_21239,N_21070);
nand U21286 (N_21286,N_21246,N_21225);
xor U21287 (N_21287,N_21024,N_21222);
or U21288 (N_21288,N_21193,N_21164);
or U21289 (N_21289,N_21099,N_21181);
xor U21290 (N_21290,N_21066,N_21111);
xor U21291 (N_21291,N_21077,N_21103);
nor U21292 (N_21292,N_21083,N_21100);
xnor U21293 (N_21293,N_21244,N_21134);
nor U21294 (N_21294,N_21035,N_21121);
nand U21295 (N_21295,N_21055,N_21080);
xnor U21296 (N_21296,N_21069,N_21057);
or U21297 (N_21297,N_21201,N_21012);
xnor U21298 (N_21298,N_21123,N_21208);
or U21299 (N_21299,N_21171,N_21137);
nand U21300 (N_21300,N_21169,N_21063);
nor U21301 (N_21301,N_21042,N_21149);
nand U21302 (N_21302,N_21140,N_21249);
xor U21303 (N_21303,N_21136,N_21029);
nor U21304 (N_21304,N_21056,N_21025);
and U21305 (N_21305,N_21054,N_21177);
nor U21306 (N_21306,N_21194,N_21036);
xor U21307 (N_21307,N_21095,N_21224);
xnor U21308 (N_21308,N_21243,N_21189);
and U21309 (N_21309,N_21232,N_21234);
nand U21310 (N_21310,N_21184,N_21212);
or U21311 (N_21311,N_21226,N_21106);
nand U21312 (N_21312,N_21018,N_21039);
or U21313 (N_21313,N_21028,N_21108);
xor U21314 (N_21314,N_21168,N_21105);
and U21315 (N_21315,N_21118,N_21202);
nand U21316 (N_21316,N_21166,N_21131);
and U21317 (N_21317,N_21186,N_21087);
or U21318 (N_21318,N_21195,N_21079);
and U21319 (N_21319,N_21013,N_21101);
xor U21320 (N_21320,N_21159,N_21228);
nand U21321 (N_21321,N_21230,N_21114);
or U21322 (N_21322,N_21183,N_21062);
nor U21323 (N_21323,N_21007,N_21221);
nor U21324 (N_21324,N_21218,N_21229);
nor U21325 (N_21325,N_21049,N_21068);
and U21326 (N_21326,N_21026,N_21037);
xor U21327 (N_21327,N_21197,N_21182);
or U21328 (N_21328,N_21081,N_21210);
nor U21329 (N_21329,N_21203,N_21048);
or U21330 (N_21330,N_21027,N_21002);
or U21331 (N_21331,N_21091,N_21061);
nor U21332 (N_21332,N_21032,N_21078);
and U21333 (N_21333,N_21017,N_21172);
and U21334 (N_21334,N_21150,N_21170);
or U21335 (N_21335,N_21217,N_21128);
nand U21336 (N_21336,N_21088,N_21021);
nand U21337 (N_21337,N_21064,N_21030);
nor U21338 (N_21338,N_21058,N_21213);
nor U21339 (N_21339,N_21248,N_21205);
and U21340 (N_21340,N_21190,N_21141);
nand U21341 (N_21341,N_21019,N_21033);
and U21342 (N_21342,N_21098,N_21011);
and U21343 (N_21343,N_21192,N_21231);
and U21344 (N_21344,N_21023,N_21220);
and U21345 (N_21345,N_21126,N_21238);
nand U21346 (N_21346,N_21008,N_21076);
nand U21347 (N_21347,N_21247,N_21223);
nand U21348 (N_21348,N_21175,N_21162);
xnor U21349 (N_21349,N_21090,N_21047);
nand U21350 (N_21350,N_21071,N_21152);
and U21351 (N_21351,N_21092,N_21214);
nand U21352 (N_21352,N_21046,N_21119);
or U21353 (N_21353,N_21096,N_21113);
or U21354 (N_21354,N_21206,N_21073);
or U21355 (N_21355,N_21130,N_21009);
or U21356 (N_21356,N_21236,N_21148);
and U21357 (N_21357,N_21038,N_21154);
nand U21358 (N_21358,N_21107,N_21167);
nand U21359 (N_21359,N_21227,N_21178);
nand U21360 (N_21360,N_21237,N_21022);
or U21361 (N_21361,N_21003,N_21000);
and U21362 (N_21362,N_21117,N_21060);
and U21363 (N_21363,N_21200,N_21045);
or U21364 (N_21364,N_21082,N_21050);
nand U21365 (N_21365,N_21053,N_21135);
and U21366 (N_21366,N_21160,N_21040);
nor U21367 (N_21367,N_21158,N_21110);
or U21368 (N_21368,N_21245,N_21176);
xnor U21369 (N_21369,N_21031,N_21204);
nor U21370 (N_21370,N_21102,N_21143);
xor U21371 (N_21371,N_21233,N_21074);
and U21372 (N_21372,N_21005,N_21144);
nand U21373 (N_21373,N_21034,N_21112);
nand U21374 (N_21374,N_21145,N_21004);
nand U21375 (N_21375,N_21063,N_21164);
or U21376 (N_21376,N_21198,N_21171);
or U21377 (N_21377,N_21011,N_21092);
nand U21378 (N_21378,N_21077,N_21113);
and U21379 (N_21379,N_21047,N_21232);
and U21380 (N_21380,N_21137,N_21048);
xor U21381 (N_21381,N_21010,N_21133);
xor U21382 (N_21382,N_21153,N_21125);
xor U21383 (N_21383,N_21078,N_21111);
nor U21384 (N_21384,N_21144,N_21243);
or U21385 (N_21385,N_21135,N_21132);
nor U21386 (N_21386,N_21155,N_21208);
or U21387 (N_21387,N_21176,N_21235);
nand U21388 (N_21388,N_21005,N_21173);
or U21389 (N_21389,N_21148,N_21066);
nand U21390 (N_21390,N_21010,N_21181);
or U21391 (N_21391,N_21243,N_21208);
xor U21392 (N_21392,N_21112,N_21234);
nand U21393 (N_21393,N_21159,N_21082);
nor U21394 (N_21394,N_21006,N_21170);
nand U21395 (N_21395,N_21036,N_21239);
nand U21396 (N_21396,N_21208,N_21152);
xor U21397 (N_21397,N_21070,N_21157);
or U21398 (N_21398,N_21015,N_21127);
nand U21399 (N_21399,N_21030,N_21185);
or U21400 (N_21400,N_21079,N_21031);
nor U21401 (N_21401,N_21171,N_21176);
and U21402 (N_21402,N_21249,N_21072);
nor U21403 (N_21403,N_21087,N_21106);
nor U21404 (N_21404,N_21205,N_21207);
nand U21405 (N_21405,N_21007,N_21084);
nor U21406 (N_21406,N_21206,N_21195);
and U21407 (N_21407,N_21067,N_21214);
nand U21408 (N_21408,N_21054,N_21144);
or U21409 (N_21409,N_21056,N_21222);
nand U21410 (N_21410,N_21168,N_21200);
nor U21411 (N_21411,N_21156,N_21186);
and U21412 (N_21412,N_21208,N_21204);
and U21413 (N_21413,N_21025,N_21175);
xnor U21414 (N_21414,N_21162,N_21025);
xnor U21415 (N_21415,N_21005,N_21187);
and U21416 (N_21416,N_21067,N_21211);
nand U21417 (N_21417,N_21132,N_21129);
or U21418 (N_21418,N_21066,N_21183);
nor U21419 (N_21419,N_21008,N_21078);
or U21420 (N_21420,N_21174,N_21077);
xnor U21421 (N_21421,N_21021,N_21005);
nor U21422 (N_21422,N_21216,N_21228);
xnor U21423 (N_21423,N_21242,N_21216);
nand U21424 (N_21424,N_21089,N_21166);
and U21425 (N_21425,N_21099,N_21092);
nor U21426 (N_21426,N_21090,N_21042);
nand U21427 (N_21427,N_21018,N_21132);
or U21428 (N_21428,N_21178,N_21038);
xor U21429 (N_21429,N_21193,N_21215);
nor U21430 (N_21430,N_21115,N_21210);
or U21431 (N_21431,N_21073,N_21185);
and U21432 (N_21432,N_21062,N_21147);
xnor U21433 (N_21433,N_21077,N_21241);
and U21434 (N_21434,N_21004,N_21241);
xor U21435 (N_21435,N_21018,N_21194);
nand U21436 (N_21436,N_21210,N_21223);
and U21437 (N_21437,N_21220,N_21149);
and U21438 (N_21438,N_21058,N_21004);
nand U21439 (N_21439,N_21142,N_21076);
nand U21440 (N_21440,N_21001,N_21082);
xor U21441 (N_21441,N_21090,N_21213);
or U21442 (N_21442,N_21140,N_21148);
nand U21443 (N_21443,N_21118,N_21072);
xor U21444 (N_21444,N_21012,N_21049);
or U21445 (N_21445,N_21143,N_21093);
and U21446 (N_21446,N_21233,N_21070);
xor U21447 (N_21447,N_21125,N_21010);
xor U21448 (N_21448,N_21162,N_21123);
or U21449 (N_21449,N_21211,N_21052);
nand U21450 (N_21450,N_21034,N_21140);
and U21451 (N_21451,N_21164,N_21064);
nor U21452 (N_21452,N_21108,N_21235);
or U21453 (N_21453,N_21215,N_21197);
xnor U21454 (N_21454,N_21089,N_21194);
xnor U21455 (N_21455,N_21016,N_21025);
nor U21456 (N_21456,N_21226,N_21157);
or U21457 (N_21457,N_21240,N_21022);
nand U21458 (N_21458,N_21195,N_21189);
nor U21459 (N_21459,N_21173,N_21095);
and U21460 (N_21460,N_21195,N_21153);
nor U21461 (N_21461,N_21037,N_21039);
or U21462 (N_21462,N_21224,N_21096);
and U21463 (N_21463,N_21155,N_21246);
nor U21464 (N_21464,N_21057,N_21070);
xnor U21465 (N_21465,N_21246,N_21065);
and U21466 (N_21466,N_21243,N_21222);
nor U21467 (N_21467,N_21156,N_21150);
xnor U21468 (N_21468,N_21020,N_21212);
and U21469 (N_21469,N_21065,N_21090);
xor U21470 (N_21470,N_21095,N_21174);
nand U21471 (N_21471,N_21113,N_21051);
and U21472 (N_21472,N_21089,N_21029);
nor U21473 (N_21473,N_21248,N_21196);
nor U21474 (N_21474,N_21026,N_21153);
nor U21475 (N_21475,N_21206,N_21137);
nor U21476 (N_21476,N_21156,N_21181);
nor U21477 (N_21477,N_21064,N_21085);
xor U21478 (N_21478,N_21188,N_21061);
nand U21479 (N_21479,N_21042,N_21073);
or U21480 (N_21480,N_21219,N_21013);
xnor U21481 (N_21481,N_21233,N_21058);
and U21482 (N_21482,N_21040,N_21199);
nand U21483 (N_21483,N_21046,N_21006);
and U21484 (N_21484,N_21106,N_21246);
and U21485 (N_21485,N_21123,N_21098);
nand U21486 (N_21486,N_21109,N_21208);
and U21487 (N_21487,N_21238,N_21076);
or U21488 (N_21488,N_21100,N_21164);
or U21489 (N_21489,N_21152,N_21065);
xnor U21490 (N_21490,N_21194,N_21105);
nand U21491 (N_21491,N_21010,N_21177);
and U21492 (N_21492,N_21243,N_21058);
nor U21493 (N_21493,N_21191,N_21030);
or U21494 (N_21494,N_21240,N_21097);
nand U21495 (N_21495,N_21099,N_21168);
nand U21496 (N_21496,N_21068,N_21100);
nand U21497 (N_21497,N_21115,N_21097);
xor U21498 (N_21498,N_21030,N_21205);
nand U21499 (N_21499,N_21154,N_21202);
nor U21500 (N_21500,N_21472,N_21282);
or U21501 (N_21501,N_21445,N_21372);
or U21502 (N_21502,N_21278,N_21464);
nor U21503 (N_21503,N_21476,N_21325);
and U21504 (N_21504,N_21438,N_21390);
xor U21505 (N_21505,N_21406,N_21331);
nor U21506 (N_21506,N_21320,N_21279);
nor U21507 (N_21507,N_21419,N_21414);
xnor U21508 (N_21508,N_21388,N_21403);
nor U21509 (N_21509,N_21352,N_21417);
nor U21510 (N_21510,N_21357,N_21275);
xor U21511 (N_21511,N_21374,N_21281);
or U21512 (N_21512,N_21466,N_21497);
and U21513 (N_21513,N_21470,N_21335);
nand U21514 (N_21514,N_21340,N_21465);
xnor U21515 (N_21515,N_21260,N_21328);
and U21516 (N_21516,N_21333,N_21385);
and U21517 (N_21517,N_21400,N_21319);
nand U21518 (N_21518,N_21410,N_21270);
xnor U21519 (N_21519,N_21444,N_21484);
nand U21520 (N_21520,N_21477,N_21268);
or U21521 (N_21521,N_21493,N_21392);
nand U21522 (N_21522,N_21269,N_21342);
xor U21523 (N_21523,N_21277,N_21349);
and U21524 (N_21524,N_21286,N_21394);
xnor U21525 (N_21525,N_21361,N_21381);
and U21526 (N_21526,N_21450,N_21370);
or U21527 (N_21527,N_21266,N_21364);
nand U21528 (N_21528,N_21274,N_21489);
and U21529 (N_21529,N_21495,N_21480);
xnor U21530 (N_21530,N_21289,N_21262);
nor U21531 (N_21531,N_21413,N_21276);
or U21532 (N_21532,N_21359,N_21448);
nor U21533 (N_21533,N_21300,N_21442);
nor U21534 (N_21534,N_21367,N_21330);
xnor U21535 (N_21535,N_21411,N_21308);
and U21536 (N_21536,N_21272,N_21421);
xor U21537 (N_21537,N_21261,N_21306);
and U21538 (N_21538,N_21440,N_21360);
nor U21539 (N_21539,N_21327,N_21259);
or U21540 (N_21540,N_21354,N_21312);
nor U21541 (N_21541,N_21280,N_21407);
xnor U21542 (N_21542,N_21290,N_21473);
nand U21543 (N_21543,N_21323,N_21437);
nand U21544 (N_21544,N_21492,N_21334);
or U21545 (N_21545,N_21426,N_21479);
nor U21546 (N_21546,N_21251,N_21378);
nand U21547 (N_21547,N_21474,N_21355);
nor U21548 (N_21548,N_21399,N_21256);
or U21549 (N_21549,N_21324,N_21386);
or U21550 (N_21550,N_21412,N_21366);
nand U21551 (N_21551,N_21391,N_21310);
nor U21552 (N_21552,N_21343,N_21432);
or U21553 (N_21553,N_21405,N_21384);
xor U21554 (N_21554,N_21318,N_21346);
nand U21555 (N_21555,N_21396,N_21255);
or U21556 (N_21556,N_21283,N_21429);
nor U21557 (N_21557,N_21447,N_21253);
nand U21558 (N_21558,N_21458,N_21423);
nand U21559 (N_21559,N_21404,N_21436);
nor U21560 (N_21560,N_21365,N_21402);
xor U21561 (N_21561,N_21299,N_21467);
nand U21562 (N_21562,N_21433,N_21428);
and U21563 (N_21563,N_21254,N_21463);
or U21564 (N_21564,N_21379,N_21491);
xor U21565 (N_21565,N_21475,N_21311);
xnor U21566 (N_21566,N_21338,N_21398);
xor U21567 (N_21567,N_21315,N_21337);
or U21568 (N_21568,N_21336,N_21303);
nand U21569 (N_21569,N_21409,N_21356);
xor U21570 (N_21570,N_21264,N_21258);
nand U21571 (N_21571,N_21288,N_21257);
xor U21572 (N_21572,N_21462,N_21457);
and U21573 (N_21573,N_21449,N_21375);
xor U21574 (N_21574,N_21295,N_21482);
xnor U21575 (N_21575,N_21353,N_21397);
nor U21576 (N_21576,N_21427,N_21494);
and U21577 (N_21577,N_21485,N_21393);
nor U21578 (N_21578,N_21309,N_21304);
and U21579 (N_21579,N_21368,N_21496);
nand U21580 (N_21580,N_21297,N_21362);
nor U21581 (N_21581,N_21294,N_21345);
xnor U21582 (N_21582,N_21291,N_21273);
xor U21583 (N_21583,N_21487,N_21443);
and U21584 (N_21584,N_21369,N_21424);
xor U21585 (N_21585,N_21305,N_21382);
and U21586 (N_21586,N_21296,N_21452);
and U21587 (N_21587,N_21321,N_21313);
nand U21588 (N_21588,N_21358,N_21326);
nand U21589 (N_21589,N_21418,N_21351);
xor U21590 (N_21590,N_21483,N_21332);
or U21591 (N_21591,N_21471,N_21329);
nand U21592 (N_21592,N_21395,N_21347);
nor U21593 (N_21593,N_21441,N_21344);
nand U21594 (N_21594,N_21389,N_21287);
nand U21595 (N_21595,N_21285,N_21387);
nor U21596 (N_21596,N_21339,N_21435);
nor U21597 (N_21597,N_21298,N_21454);
xor U21598 (N_21598,N_21314,N_21265);
nor U21599 (N_21599,N_21460,N_21446);
and U21600 (N_21600,N_21383,N_21499);
nand U21601 (N_21601,N_21431,N_21416);
or U21602 (N_21602,N_21348,N_21434);
or U21603 (N_21603,N_21373,N_21293);
and U21604 (N_21604,N_21498,N_21451);
and U21605 (N_21605,N_21267,N_21422);
nand U21606 (N_21606,N_21363,N_21486);
nor U21607 (N_21607,N_21317,N_21302);
and U21608 (N_21608,N_21488,N_21469);
or U21609 (N_21609,N_21292,N_21307);
or U21610 (N_21610,N_21456,N_21341);
nor U21611 (N_21611,N_21453,N_21439);
nor U21612 (N_21612,N_21490,N_21481);
xor U21613 (N_21613,N_21284,N_21271);
xor U21614 (N_21614,N_21468,N_21263);
xor U21615 (N_21615,N_21376,N_21371);
and U21616 (N_21616,N_21408,N_21415);
or U21617 (N_21617,N_21380,N_21322);
xnor U21618 (N_21618,N_21250,N_21420);
nand U21619 (N_21619,N_21478,N_21377);
or U21620 (N_21620,N_21252,N_21459);
or U21621 (N_21621,N_21401,N_21301);
nor U21622 (N_21622,N_21430,N_21461);
nor U21623 (N_21623,N_21316,N_21425);
xnor U21624 (N_21624,N_21455,N_21350);
or U21625 (N_21625,N_21473,N_21259);
xor U21626 (N_21626,N_21269,N_21453);
and U21627 (N_21627,N_21329,N_21454);
xnor U21628 (N_21628,N_21312,N_21393);
or U21629 (N_21629,N_21392,N_21422);
xnor U21630 (N_21630,N_21406,N_21271);
and U21631 (N_21631,N_21445,N_21333);
and U21632 (N_21632,N_21401,N_21398);
nand U21633 (N_21633,N_21290,N_21417);
xor U21634 (N_21634,N_21377,N_21352);
or U21635 (N_21635,N_21251,N_21439);
nor U21636 (N_21636,N_21443,N_21303);
and U21637 (N_21637,N_21277,N_21289);
and U21638 (N_21638,N_21354,N_21350);
nand U21639 (N_21639,N_21393,N_21488);
and U21640 (N_21640,N_21480,N_21353);
or U21641 (N_21641,N_21287,N_21382);
nand U21642 (N_21642,N_21411,N_21439);
nor U21643 (N_21643,N_21265,N_21340);
and U21644 (N_21644,N_21288,N_21450);
and U21645 (N_21645,N_21336,N_21483);
xnor U21646 (N_21646,N_21343,N_21465);
xnor U21647 (N_21647,N_21428,N_21336);
nor U21648 (N_21648,N_21434,N_21476);
xor U21649 (N_21649,N_21465,N_21277);
or U21650 (N_21650,N_21317,N_21428);
nand U21651 (N_21651,N_21359,N_21361);
and U21652 (N_21652,N_21367,N_21268);
nor U21653 (N_21653,N_21383,N_21376);
or U21654 (N_21654,N_21297,N_21422);
nor U21655 (N_21655,N_21391,N_21250);
nand U21656 (N_21656,N_21455,N_21499);
nor U21657 (N_21657,N_21389,N_21336);
nand U21658 (N_21658,N_21466,N_21291);
and U21659 (N_21659,N_21305,N_21343);
nor U21660 (N_21660,N_21272,N_21402);
nor U21661 (N_21661,N_21365,N_21253);
or U21662 (N_21662,N_21475,N_21499);
and U21663 (N_21663,N_21408,N_21414);
or U21664 (N_21664,N_21497,N_21268);
and U21665 (N_21665,N_21322,N_21341);
nor U21666 (N_21666,N_21273,N_21365);
or U21667 (N_21667,N_21328,N_21383);
nor U21668 (N_21668,N_21331,N_21271);
nor U21669 (N_21669,N_21374,N_21461);
or U21670 (N_21670,N_21344,N_21276);
nor U21671 (N_21671,N_21466,N_21325);
nand U21672 (N_21672,N_21366,N_21475);
or U21673 (N_21673,N_21253,N_21476);
nor U21674 (N_21674,N_21492,N_21387);
xor U21675 (N_21675,N_21264,N_21250);
nand U21676 (N_21676,N_21400,N_21377);
nand U21677 (N_21677,N_21476,N_21355);
nor U21678 (N_21678,N_21442,N_21356);
nand U21679 (N_21679,N_21464,N_21377);
nand U21680 (N_21680,N_21479,N_21382);
or U21681 (N_21681,N_21457,N_21429);
nand U21682 (N_21682,N_21439,N_21270);
and U21683 (N_21683,N_21464,N_21401);
or U21684 (N_21684,N_21302,N_21429);
xnor U21685 (N_21685,N_21340,N_21405);
nor U21686 (N_21686,N_21433,N_21323);
and U21687 (N_21687,N_21342,N_21489);
xnor U21688 (N_21688,N_21478,N_21362);
and U21689 (N_21689,N_21499,N_21329);
and U21690 (N_21690,N_21466,N_21393);
or U21691 (N_21691,N_21383,N_21347);
or U21692 (N_21692,N_21375,N_21392);
nand U21693 (N_21693,N_21283,N_21439);
nand U21694 (N_21694,N_21340,N_21468);
xor U21695 (N_21695,N_21283,N_21338);
and U21696 (N_21696,N_21470,N_21486);
and U21697 (N_21697,N_21261,N_21469);
nand U21698 (N_21698,N_21441,N_21498);
nor U21699 (N_21699,N_21355,N_21477);
or U21700 (N_21700,N_21377,N_21270);
and U21701 (N_21701,N_21280,N_21448);
nand U21702 (N_21702,N_21260,N_21355);
or U21703 (N_21703,N_21395,N_21353);
xor U21704 (N_21704,N_21475,N_21291);
xnor U21705 (N_21705,N_21376,N_21414);
nand U21706 (N_21706,N_21363,N_21268);
or U21707 (N_21707,N_21289,N_21329);
xnor U21708 (N_21708,N_21436,N_21335);
xor U21709 (N_21709,N_21458,N_21337);
nand U21710 (N_21710,N_21309,N_21382);
xnor U21711 (N_21711,N_21377,N_21406);
xnor U21712 (N_21712,N_21398,N_21383);
xor U21713 (N_21713,N_21287,N_21433);
nand U21714 (N_21714,N_21257,N_21492);
nor U21715 (N_21715,N_21250,N_21300);
nand U21716 (N_21716,N_21337,N_21344);
and U21717 (N_21717,N_21275,N_21297);
or U21718 (N_21718,N_21371,N_21292);
and U21719 (N_21719,N_21372,N_21331);
xor U21720 (N_21720,N_21343,N_21477);
nor U21721 (N_21721,N_21307,N_21462);
and U21722 (N_21722,N_21327,N_21293);
nor U21723 (N_21723,N_21326,N_21295);
or U21724 (N_21724,N_21321,N_21459);
xnor U21725 (N_21725,N_21395,N_21373);
xnor U21726 (N_21726,N_21384,N_21303);
or U21727 (N_21727,N_21410,N_21316);
nor U21728 (N_21728,N_21490,N_21467);
nand U21729 (N_21729,N_21374,N_21291);
xor U21730 (N_21730,N_21495,N_21481);
and U21731 (N_21731,N_21450,N_21471);
or U21732 (N_21732,N_21499,N_21285);
xor U21733 (N_21733,N_21426,N_21251);
nand U21734 (N_21734,N_21274,N_21273);
and U21735 (N_21735,N_21256,N_21408);
xnor U21736 (N_21736,N_21373,N_21324);
nor U21737 (N_21737,N_21417,N_21268);
and U21738 (N_21738,N_21348,N_21398);
nor U21739 (N_21739,N_21467,N_21477);
or U21740 (N_21740,N_21292,N_21317);
nor U21741 (N_21741,N_21376,N_21294);
nor U21742 (N_21742,N_21318,N_21493);
and U21743 (N_21743,N_21496,N_21370);
and U21744 (N_21744,N_21322,N_21339);
or U21745 (N_21745,N_21435,N_21395);
or U21746 (N_21746,N_21397,N_21324);
or U21747 (N_21747,N_21363,N_21309);
and U21748 (N_21748,N_21254,N_21442);
nand U21749 (N_21749,N_21316,N_21385);
xor U21750 (N_21750,N_21644,N_21536);
xnor U21751 (N_21751,N_21709,N_21605);
nor U21752 (N_21752,N_21560,N_21542);
nor U21753 (N_21753,N_21587,N_21656);
xnor U21754 (N_21754,N_21505,N_21686);
and U21755 (N_21755,N_21527,N_21654);
nor U21756 (N_21756,N_21699,N_21609);
xnor U21757 (N_21757,N_21626,N_21611);
and U21758 (N_21758,N_21503,N_21738);
nor U21759 (N_21759,N_21680,N_21578);
and U21760 (N_21760,N_21546,N_21511);
xnor U21761 (N_21761,N_21566,N_21531);
xor U21762 (N_21762,N_21691,N_21675);
xnor U21763 (N_21763,N_21603,N_21621);
nand U21764 (N_21764,N_21519,N_21634);
and U21765 (N_21765,N_21633,N_21647);
nand U21766 (N_21766,N_21722,N_21522);
or U21767 (N_21767,N_21517,N_21668);
or U21768 (N_21768,N_21562,N_21665);
and U21769 (N_21769,N_21606,N_21617);
and U21770 (N_21770,N_21741,N_21518);
xnor U21771 (N_21771,N_21627,N_21748);
nand U21772 (N_21772,N_21506,N_21586);
xnor U21773 (N_21773,N_21544,N_21698);
nor U21774 (N_21774,N_21583,N_21704);
and U21775 (N_21775,N_21701,N_21613);
nor U21776 (N_21776,N_21660,N_21574);
nand U21777 (N_21777,N_21657,N_21702);
and U21778 (N_21778,N_21658,N_21715);
or U21779 (N_21779,N_21696,N_21508);
nand U21780 (N_21780,N_21557,N_21664);
xor U21781 (N_21781,N_21735,N_21661);
nor U21782 (N_21782,N_21565,N_21520);
nor U21783 (N_21783,N_21650,N_21620);
or U21784 (N_21784,N_21512,N_21602);
xnor U21785 (N_21785,N_21729,N_21711);
or U21786 (N_21786,N_21618,N_21734);
xor U21787 (N_21787,N_21585,N_21721);
nand U21788 (N_21788,N_21552,N_21526);
and U21789 (N_21789,N_21539,N_21676);
xor U21790 (N_21790,N_21513,N_21652);
nand U21791 (N_21791,N_21684,N_21577);
or U21792 (N_21792,N_21662,N_21563);
nor U21793 (N_21793,N_21730,N_21608);
and U21794 (N_21794,N_21706,N_21538);
or U21795 (N_21795,N_21573,N_21708);
nor U21796 (N_21796,N_21590,N_21718);
and U21797 (N_21797,N_21631,N_21612);
nor U21798 (N_21798,N_21543,N_21619);
nand U21799 (N_21799,N_21521,N_21582);
nand U21800 (N_21800,N_21659,N_21670);
xnor U21801 (N_21801,N_21651,N_21584);
nand U21802 (N_21802,N_21549,N_21713);
and U21803 (N_21803,N_21726,N_21710);
and U21804 (N_21804,N_21632,N_21604);
or U21805 (N_21805,N_21559,N_21690);
or U21806 (N_21806,N_21623,N_21558);
nor U21807 (N_21807,N_21591,N_21588);
xor U21808 (N_21808,N_21622,N_21693);
nand U21809 (N_21809,N_21534,N_21733);
nor U21810 (N_21810,N_21616,N_21663);
nor U21811 (N_21811,N_21674,N_21695);
or U21812 (N_21812,N_21745,N_21714);
nand U21813 (N_21813,N_21598,N_21571);
and U21814 (N_21814,N_21524,N_21599);
or U21815 (N_21815,N_21553,N_21689);
nor U21816 (N_21816,N_21731,N_21640);
nor U21817 (N_21817,N_21725,N_21610);
xnor U21818 (N_21818,N_21672,N_21700);
nand U21819 (N_21819,N_21593,N_21507);
and U21820 (N_21820,N_21717,N_21548);
or U21821 (N_21821,N_21705,N_21597);
nand U21822 (N_21822,N_21724,N_21596);
or U21823 (N_21823,N_21692,N_21648);
nor U21824 (N_21824,N_21638,N_21561);
nor U21825 (N_21825,N_21630,N_21643);
xor U21826 (N_21826,N_21592,N_21607);
nor U21827 (N_21827,N_21637,N_21569);
or U21828 (N_21828,N_21579,N_21635);
nand U21829 (N_21829,N_21697,N_21510);
xnor U21830 (N_21830,N_21550,N_21625);
xor U21831 (N_21831,N_21589,N_21515);
xor U21832 (N_21832,N_21501,N_21514);
nand U21833 (N_21833,N_21739,N_21547);
xor U21834 (N_21834,N_21594,N_21545);
nor U21835 (N_21835,N_21564,N_21737);
or U21836 (N_21836,N_21649,N_21740);
nand U21837 (N_21837,N_21677,N_21567);
xnor U21838 (N_21838,N_21646,N_21727);
nor U21839 (N_21839,N_21723,N_21642);
or U21840 (N_21840,N_21694,N_21673);
nor U21841 (N_21841,N_21535,N_21749);
or U21842 (N_21842,N_21614,N_21525);
and U21843 (N_21843,N_21533,N_21502);
and U21844 (N_21844,N_21682,N_21728);
and U21845 (N_21845,N_21595,N_21707);
nand U21846 (N_21846,N_21576,N_21720);
nand U21847 (N_21847,N_21555,N_21580);
nor U21848 (N_21848,N_21703,N_21655);
xor U21849 (N_21849,N_21575,N_21509);
nand U21850 (N_21850,N_21645,N_21541);
nand U21851 (N_21851,N_21570,N_21744);
xor U21852 (N_21852,N_21601,N_21639);
or U21853 (N_21853,N_21581,N_21681);
or U21854 (N_21854,N_21732,N_21529);
xnor U21855 (N_21855,N_21712,N_21500);
or U21856 (N_21856,N_21683,N_21551);
nand U21857 (N_21857,N_21516,N_21600);
and U21858 (N_21858,N_21678,N_21688);
nor U21859 (N_21859,N_21685,N_21679);
xnor U21860 (N_21860,N_21669,N_21504);
nand U21861 (N_21861,N_21641,N_21736);
and U21862 (N_21862,N_21540,N_21687);
and U21863 (N_21863,N_21572,N_21537);
xor U21864 (N_21864,N_21671,N_21636);
nand U21865 (N_21865,N_21742,N_21615);
and U21866 (N_21866,N_21568,N_21666);
nand U21867 (N_21867,N_21554,N_21719);
or U21868 (N_21868,N_21629,N_21716);
and U21869 (N_21869,N_21667,N_21532);
nor U21870 (N_21870,N_21743,N_21628);
nand U21871 (N_21871,N_21747,N_21556);
xnor U21872 (N_21872,N_21530,N_21528);
nor U21873 (N_21873,N_21746,N_21624);
or U21874 (N_21874,N_21523,N_21653);
nor U21875 (N_21875,N_21740,N_21691);
and U21876 (N_21876,N_21532,N_21656);
or U21877 (N_21877,N_21538,N_21718);
xor U21878 (N_21878,N_21745,N_21749);
and U21879 (N_21879,N_21698,N_21719);
nand U21880 (N_21880,N_21714,N_21502);
or U21881 (N_21881,N_21579,N_21595);
nand U21882 (N_21882,N_21667,N_21605);
and U21883 (N_21883,N_21745,N_21681);
xor U21884 (N_21884,N_21642,N_21634);
xnor U21885 (N_21885,N_21611,N_21508);
and U21886 (N_21886,N_21713,N_21603);
and U21887 (N_21887,N_21649,N_21644);
nor U21888 (N_21888,N_21642,N_21691);
or U21889 (N_21889,N_21544,N_21528);
nand U21890 (N_21890,N_21512,N_21697);
or U21891 (N_21891,N_21528,N_21504);
and U21892 (N_21892,N_21739,N_21749);
nor U21893 (N_21893,N_21594,N_21505);
nand U21894 (N_21894,N_21637,N_21519);
nand U21895 (N_21895,N_21664,N_21737);
xnor U21896 (N_21896,N_21612,N_21531);
nor U21897 (N_21897,N_21719,N_21659);
nand U21898 (N_21898,N_21502,N_21740);
nor U21899 (N_21899,N_21503,N_21641);
nor U21900 (N_21900,N_21746,N_21595);
or U21901 (N_21901,N_21676,N_21730);
xor U21902 (N_21902,N_21501,N_21747);
nand U21903 (N_21903,N_21578,N_21695);
xor U21904 (N_21904,N_21577,N_21547);
or U21905 (N_21905,N_21625,N_21646);
nand U21906 (N_21906,N_21591,N_21633);
or U21907 (N_21907,N_21623,N_21686);
nand U21908 (N_21908,N_21668,N_21690);
or U21909 (N_21909,N_21561,N_21662);
nand U21910 (N_21910,N_21542,N_21543);
nor U21911 (N_21911,N_21554,N_21727);
or U21912 (N_21912,N_21657,N_21612);
nor U21913 (N_21913,N_21572,N_21610);
xor U21914 (N_21914,N_21500,N_21601);
nand U21915 (N_21915,N_21533,N_21681);
nand U21916 (N_21916,N_21582,N_21522);
xnor U21917 (N_21917,N_21613,N_21671);
nor U21918 (N_21918,N_21642,N_21557);
or U21919 (N_21919,N_21539,N_21629);
or U21920 (N_21920,N_21646,N_21557);
or U21921 (N_21921,N_21575,N_21691);
nand U21922 (N_21922,N_21537,N_21720);
or U21923 (N_21923,N_21678,N_21748);
nor U21924 (N_21924,N_21577,N_21575);
nor U21925 (N_21925,N_21737,N_21531);
nor U21926 (N_21926,N_21647,N_21571);
nand U21927 (N_21927,N_21646,N_21601);
nand U21928 (N_21928,N_21529,N_21664);
nand U21929 (N_21929,N_21686,N_21507);
or U21930 (N_21930,N_21681,N_21631);
and U21931 (N_21931,N_21615,N_21596);
nor U21932 (N_21932,N_21597,N_21710);
xnor U21933 (N_21933,N_21704,N_21510);
or U21934 (N_21934,N_21577,N_21742);
or U21935 (N_21935,N_21603,N_21531);
and U21936 (N_21936,N_21541,N_21654);
xor U21937 (N_21937,N_21722,N_21708);
xnor U21938 (N_21938,N_21701,N_21592);
nand U21939 (N_21939,N_21601,N_21552);
nand U21940 (N_21940,N_21521,N_21630);
xnor U21941 (N_21941,N_21551,N_21742);
or U21942 (N_21942,N_21715,N_21707);
nand U21943 (N_21943,N_21585,N_21695);
or U21944 (N_21944,N_21534,N_21582);
nor U21945 (N_21945,N_21599,N_21627);
or U21946 (N_21946,N_21564,N_21574);
or U21947 (N_21947,N_21694,N_21593);
and U21948 (N_21948,N_21686,N_21643);
and U21949 (N_21949,N_21731,N_21570);
nand U21950 (N_21950,N_21582,N_21729);
or U21951 (N_21951,N_21560,N_21677);
nand U21952 (N_21952,N_21691,N_21555);
nand U21953 (N_21953,N_21526,N_21742);
xor U21954 (N_21954,N_21714,N_21721);
nand U21955 (N_21955,N_21549,N_21502);
and U21956 (N_21956,N_21665,N_21604);
nand U21957 (N_21957,N_21643,N_21724);
nor U21958 (N_21958,N_21545,N_21555);
or U21959 (N_21959,N_21717,N_21529);
and U21960 (N_21960,N_21611,N_21613);
or U21961 (N_21961,N_21598,N_21668);
and U21962 (N_21962,N_21580,N_21724);
xor U21963 (N_21963,N_21694,N_21625);
xor U21964 (N_21964,N_21710,N_21631);
and U21965 (N_21965,N_21588,N_21716);
nor U21966 (N_21966,N_21528,N_21666);
xnor U21967 (N_21967,N_21718,N_21530);
and U21968 (N_21968,N_21691,N_21641);
xor U21969 (N_21969,N_21747,N_21554);
nand U21970 (N_21970,N_21540,N_21611);
nand U21971 (N_21971,N_21677,N_21632);
and U21972 (N_21972,N_21682,N_21537);
and U21973 (N_21973,N_21661,N_21747);
xor U21974 (N_21974,N_21575,N_21512);
xor U21975 (N_21975,N_21618,N_21665);
nand U21976 (N_21976,N_21687,N_21524);
or U21977 (N_21977,N_21628,N_21717);
or U21978 (N_21978,N_21707,N_21710);
or U21979 (N_21979,N_21602,N_21533);
xor U21980 (N_21980,N_21698,N_21713);
nor U21981 (N_21981,N_21523,N_21732);
nand U21982 (N_21982,N_21745,N_21666);
nor U21983 (N_21983,N_21685,N_21716);
nor U21984 (N_21984,N_21553,N_21709);
and U21985 (N_21985,N_21681,N_21522);
and U21986 (N_21986,N_21557,N_21702);
and U21987 (N_21987,N_21604,N_21549);
nor U21988 (N_21988,N_21600,N_21736);
xor U21989 (N_21989,N_21734,N_21673);
and U21990 (N_21990,N_21520,N_21569);
xor U21991 (N_21991,N_21693,N_21617);
or U21992 (N_21992,N_21672,N_21641);
xor U21993 (N_21993,N_21628,N_21736);
and U21994 (N_21994,N_21600,N_21656);
xnor U21995 (N_21995,N_21694,N_21747);
or U21996 (N_21996,N_21582,N_21567);
or U21997 (N_21997,N_21594,N_21700);
nand U21998 (N_21998,N_21520,N_21749);
nand U21999 (N_21999,N_21728,N_21611);
or U22000 (N_22000,N_21835,N_21775);
or U22001 (N_22001,N_21999,N_21855);
nand U22002 (N_22002,N_21811,N_21988);
nand U22003 (N_22003,N_21843,N_21960);
nor U22004 (N_22004,N_21758,N_21910);
nand U22005 (N_22005,N_21787,N_21878);
xor U22006 (N_22006,N_21861,N_21957);
xor U22007 (N_22007,N_21992,N_21981);
xor U22008 (N_22008,N_21929,N_21970);
and U22009 (N_22009,N_21871,N_21862);
or U22010 (N_22010,N_21978,N_21954);
nor U22011 (N_22011,N_21967,N_21905);
xor U22012 (N_22012,N_21779,N_21808);
or U22013 (N_22013,N_21942,N_21868);
and U22014 (N_22014,N_21955,N_21791);
nor U22015 (N_22015,N_21993,N_21977);
and U22016 (N_22016,N_21937,N_21824);
and U22017 (N_22017,N_21872,N_21854);
nor U22018 (N_22018,N_21925,N_21947);
and U22019 (N_22019,N_21839,N_21900);
and U22020 (N_22020,N_21965,N_21917);
or U22021 (N_22021,N_21897,N_21788);
nor U22022 (N_22022,N_21891,N_21783);
xor U22023 (N_22023,N_21934,N_21903);
nor U22024 (N_22024,N_21928,N_21939);
xnor U22025 (N_22025,N_21781,N_21936);
nand U22026 (N_22026,N_21828,N_21831);
xnor U22027 (N_22027,N_21819,N_21794);
nor U22028 (N_22028,N_21909,N_21969);
or U22029 (N_22029,N_21818,N_21989);
and U22030 (N_22030,N_21906,N_21885);
and U22031 (N_22031,N_21904,N_21948);
or U22032 (N_22032,N_21887,N_21964);
and U22033 (N_22033,N_21777,N_21851);
nand U22034 (N_22034,N_21813,N_21973);
xnor U22035 (N_22035,N_21852,N_21884);
nand U22036 (N_22036,N_21952,N_21867);
or U22037 (N_22037,N_21963,N_21821);
nor U22038 (N_22038,N_21816,N_21807);
nor U22039 (N_22039,N_21796,N_21982);
and U22040 (N_22040,N_21950,N_21888);
or U22041 (N_22041,N_21853,N_21763);
or U22042 (N_22042,N_21890,N_21784);
or U22043 (N_22043,N_21926,N_21859);
nor U22044 (N_22044,N_21953,N_21951);
nand U22045 (N_22045,N_21832,N_21765);
or U22046 (N_22046,N_21924,N_21901);
xor U22047 (N_22047,N_21930,N_21764);
nor U22048 (N_22048,N_21801,N_21927);
xnor U22049 (N_22049,N_21789,N_21911);
xor U22050 (N_22050,N_21792,N_21983);
xnor U22051 (N_22051,N_21908,N_21753);
nand U22052 (N_22052,N_21771,N_21817);
nand U22053 (N_22053,N_21757,N_21938);
xor U22054 (N_22054,N_21756,N_21877);
or U22055 (N_22055,N_21804,N_21769);
nand U22056 (N_22056,N_21920,N_21760);
nor U22057 (N_22057,N_21889,N_21844);
nand U22058 (N_22058,N_21914,N_21767);
xor U22059 (N_22059,N_21991,N_21799);
or U22060 (N_22060,N_21795,N_21902);
and U22061 (N_22061,N_21976,N_21880);
nand U22062 (N_22062,N_21933,N_21815);
and U22063 (N_22063,N_21941,N_21840);
nor U22064 (N_22064,N_21921,N_21766);
or U22065 (N_22065,N_21860,N_21834);
xor U22066 (N_22066,N_21800,N_21845);
nor U22067 (N_22067,N_21864,N_21886);
and U22068 (N_22068,N_21797,N_21874);
nor U22069 (N_22069,N_21847,N_21959);
or U22070 (N_22070,N_21849,N_21833);
nor U22071 (N_22071,N_21785,N_21896);
and U22072 (N_22072,N_21987,N_21912);
and U22073 (N_22073,N_21883,N_21949);
nand U22074 (N_22074,N_21966,N_21761);
xnor U22075 (N_22075,N_21944,N_21858);
xnor U22076 (N_22076,N_21986,N_21857);
nand U22077 (N_22077,N_21958,N_21923);
and U22078 (N_22078,N_21997,N_21984);
or U22079 (N_22079,N_21946,N_21809);
nor U22080 (N_22080,N_21995,N_21848);
or U22081 (N_22081,N_21956,N_21894);
and U22082 (N_22082,N_21968,N_21772);
xnor U22083 (N_22083,N_21759,N_21866);
nand U22084 (N_22084,N_21931,N_21842);
or U22085 (N_22085,N_21856,N_21962);
or U22086 (N_22086,N_21980,N_21822);
nor U22087 (N_22087,N_21899,N_21971);
and U22088 (N_22088,N_21943,N_21907);
or U22089 (N_22089,N_21895,N_21836);
xor U22090 (N_22090,N_21774,N_21935);
nor U22091 (N_22091,N_21922,N_21994);
nand U22092 (N_22092,N_21841,N_21870);
or U22093 (N_22093,N_21780,N_21812);
and U22094 (N_22094,N_21916,N_21919);
xor U22095 (N_22095,N_21873,N_21881);
nor U22096 (N_22096,N_21974,N_21837);
and U22097 (N_22097,N_21893,N_21750);
xnor U22098 (N_22098,N_21826,N_21770);
or U22099 (N_22099,N_21790,N_21802);
or U22100 (N_22100,N_21829,N_21918);
xor U22101 (N_22101,N_21869,N_21782);
and U22102 (N_22102,N_21972,N_21755);
and U22103 (N_22103,N_21882,N_21798);
xnor U22104 (N_22104,N_21892,N_21786);
nand U22105 (N_22105,N_21751,N_21876);
nor U22106 (N_22106,N_21979,N_21915);
xnor U22107 (N_22107,N_21996,N_21754);
xnor U22108 (N_22108,N_21823,N_21810);
nand U22109 (N_22109,N_21850,N_21803);
nand U22110 (N_22110,N_21879,N_21865);
nand U22111 (N_22111,N_21961,N_21820);
and U22112 (N_22112,N_21985,N_21762);
and U22113 (N_22113,N_21863,N_21805);
nor U22114 (N_22114,N_21814,N_21975);
nor U22115 (N_22115,N_21846,N_21932);
and U22116 (N_22116,N_21998,N_21793);
nor U22117 (N_22117,N_21913,N_21990);
nand U22118 (N_22118,N_21806,N_21830);
and U22119 (N_22119,N_21827,N_21776);
and U22120 (N_22120,N_21945,N_21940);
and U22121 (N_22121,N_21768,N_21838);
and U22122 (N_22122,N_21875,N_21773);
and U22123 (N_22123,N_21825,N_21752);
and U22124 (N_22124,N_21778,N_21898);
and U22125 (N_22125,N_21958,N_21914);
nor U22126 (N_22126,N_21797,N_21910);
xor U22127 (N_22127,N_21754,N_21894);
nand U22128 (N_22128,N_21768,N_21875);
and U22129 (N_22129,N_21930,N_21961);
xnor U22130 (N_22130,N_21964,N_21880);
xor U22131 (N_22131,N_21830,N_21991);
xor U22132 (N_22132,N_21916,N_21926);
nor U22133 (N_22133,N_21995,N_21877);
nor U22134 (N_22134,N_21806,N_21856);
nand U22135 (N_22135,N_21992,N_21767);
nor U22136 (N_22136,N_21778,N_21848);
or U22137 (N_22137,N_21807,N_21804);
and U22138 (N_22138,N_21758,N_21870);
xor U22139 (N_22139,N_21777,N_21948);
xor U22140 (N_22140,N_21767,N_21753);
nor U22141 (N_22141,N_21760,N_21848);
xnor U22142 (N_22142,N_21757,N_21761);
xor U22143 (N_22143,N_21966,N_21837);
xor U22144 (N_22144,N_21801,N_21849);
nand U22145 (N_22145,N_21989,N_21938);
and U22146 (N_22146,N_21817,N_21779);
nand U22147 (N_22147,N_21806,N_21815);
nand U22148 (N_22148,N_21817,N_21781);
nand U22149 (N_22149,N_21858,N_21769);
or U22150 (N_22150,N_21878,N_21930);
and U22151 (N_22151,N_21918,N_21853);
or U22152 (N_22152,N_21888,N_21858);
and U22153 (N_22153,N_21881,N_21951);
xnor U22154 (N_22154,N_21996,N_21963);
or U22155 (N_22155,N_21943,N_21992);
nor U22156 (N_22156,N_21850,N_21792);
and U22157 (N_22157,N_21963,N_21990);
and U22158 (N_22158,N_21761,N_21755);
xnor U22159 (N_22159,N_21960,N_21913);
xnor U22160 (N_22160,N_21958,N_21916);
or U22161 (N_22161,N_21791,N_21809);
or U22162 (N_22162,N_21882,N_21898);
nor U22163 (N_22163,N_21772,N_21859);
nor U22164 (N_22164,N_21910,N_21977);
nand U22165 (N_22165,N_21892,N_21912);
nor U22166 (N_22166,N_21786,N_21805);
or U22167 (N_22167,N_21790,N_21825);
nor U22168 (N_22168,N_21989,N_21905);
and U22169 (N_22169,N_21825,N_21826);
xnor U22170 (N_22170,N_21840,N_21925);
nor U22171 (N_22171,N_21778,N_21900);
nand U22172 (N_22172,N_21968,N_21978);
nor U22173 (N_22173,N_21965,N_21890);
or U22174 (N_22174,N_21909,N_21807);
or U22175 (N_22175,N_21897,N_21909);
xnor U22176 (N_22176,N_21803,N_21848);
or U22177 (N_22177,N_21768,N_21821);
and U22178 (N_22178,N_21894,N_21796);
or U22179 (N_22179,N_21839,N_21979);
and U22180 (N_22180,N_21808,N_21883);
and U22181 (N_22181,N_21774,N_21788);
and U22182 (N_22182,N_21969,N_21946);
or U22183 (N_22183,N_21846,N_21789);
xnor U22184 (N_22184,N_21977,N_21799);
nand U22185 (N_22185,N_21973,N_21898);
and U22186 (N_22186,N_21794,N_21855);
and U22187 (N_22187,N_21878,N_21858);
xnor U22188 (N_22188,N_21875,N_21837);
nand U22189 (N_22189,N_21795,N_21750);
and U22190 (N_22190,N_21859,N_21836);
and U22191 (N_22191,N_21780,N_21854);
xor U22192 (N_22192,N_21827,N_21950);
or U22193 (N_22193,N_21902,N_21756);
nor U22194 (N_22194,N_21998,N_21884);
nand U22195 (N_22195,N_21800,N_21760);
nor U22196 (N_22196,N_21855,N_21758);
nand U22197 (N_22197,N_21763,N_21799);
nor U22198 (N_22198,N_21785,N_21889);
xnor U22199 (N_22199,N_21937,N_21828);
and U22200 (N_22200,N_21772,N_21864);
nor U22201 (N_22201,N_21925,N_21911);
xor U22202 (N_22202,N_21982,N_21823);
or U22203 (N_22203,N_21966,N_21879);
or U22204 (N_22204,N_21851,N_21885);
nand U22205 (N_22205,N_21777,N_21968);
and U22206 (N_22206,N_21977,N_21843);
or U22207 (N_22207,N_21970,N_21887);
and U22208 (N_22208,N_21906,N_21863);
nand U22209 (N_22209,N_21791,N_21835);
nand U22210 (N_22210,N_21904,N_21991);
or U22211 (N_22211,N_21924,N_21951);
and U22212 (N_22212,N_21979,N_21783);
or U22213 (N_22213,N_21869,N_21910);
nor U22214 (N_22214,N_21820,N_21881);
and U22215 (N_22215,N_21938,N_21800);
and U22216 (N_22216,N_21958,N_21826);
nor U22217 (N_22217,N_21986,N_21855);
and U22218 (N_22218,N_21795,N_21880);
or U22219 (N_22219,N_21770,N_21885);
xor U22220 (N_22220,N_21915,N_21948);
nand U22221 (N_22221,N_21807,N_21958);
nand U22222 (N_22222,N_21766,N_21977);
nor U22223 (N_22223,N_21831,N_21884);
nand U22224 (N_22224,N_21761,N_21963);
and U22225 (N_22225,N_21844,N_21843);
nor U22226 (N_22226,N_21861,N_21859);
or U22227 (N_22227,N_21877,N_21980);
or U22228 (N_22228,N_21843,N_21856);
xor U22229 (N_22229,N_21925,N_21774);
nor U22230 (N_22230,N_21785,N_21844);
nand U22231 (N_22231,N_21887,N_21833);
xor U22232 (N_22232,N_21849,N_21840);
or U22233 (N_22233,N_21929,N_21998);
or U22234 (N_22234,N_21969,N_21756);
nor U22235 (N_22235,N_21966,N_21927);
or U22236 (N_22236,N_21906,N_21841);
nand U22237 (N_22237,N_21903,N_21925);
and U22238 (N_22238,N_21983,N_21928);
xnor U22239 (N_22239,N_21851,N_21927);
or U22240 (N_22240,N_21799,N_21888);
nor U22241 (N_22241,N_21838,N_21779);
and U22242 (N_22242,N_21913,N_21857);
xnor U22243 (N_22243,N_21788,N_21953);
xnor U22244 (N_22244,N_21910,N_21777);
xnor U22245 (N_22245,N_21766,N_21853);
nand U22246 (N_22246,N_21976,N_21987);
and U22247 (N_22247,N_21886,N_21778);
nand U22248 (N_22248,N_21897,N_21791);
xnor U22249 (N_22249,N_21855,N_21839);
nand U22250 (N_22250,N_22212,N_22089);
or U22251 (N_22251,N_22101,N_22069);
and U22252 (N_22252,N_22008,N_22058);
xor U22253 (N_22253,N_22004,N_22220);
nor U22254 (N_22254,N_22156,N_22093);
and U22255 (N_22255,N_22150,N_22000);
nand U22256 (N_22256,N_22096,N_22038);
nand U22257 (N_22257,N_22181,N_22182);
and U22258 (N_22258,N_22064,N_22235);
nand U22259 (N_22259,N_22194,N_22110);
and U22260 (N_22260,N_22134,N_22129);
nand U22261 (N_22261,N_22246,N_22189);
and U22262 (N_22262,N_22006,N_22188);
and U22263 (N_22263,N_22198,N_22208);
nand U22264 (N_22264,N_22226,N_22245);
nor U22265 (N_22265,N_22161,N_22046);
xor U22266 (N_22266,N_22209,N_22190);
or U22267 (N_22267,N_22137,N_22071);
and U22268 (N_22268,N_22185,N_22230);
nand U22269 (N_22269,N_22221,N_22196);
or U22270 (N_22270,N_22128,N_22169);
xnor U22271 (N_22271,N_22041,N_22079);
or U22272 (N_22272,N_22073,N_22139);
xnor U22273 (N_22273,N_22030,N_22216);
xor U22274 (N_22274,N_22201,N_22075);
or U22275 (N_22275,N_22233,N_22056);
or U22276 (N_22276,N_22237,N_22033);
nor U22277 (N_22277,N_22215,N_22088);
xor U22278 (N_22278,N_22214,N_22067);
xnor U22279 (N_22279,N_22010,N_22239);
and U22280 (N_22280,N_22231,N_22159);
or U22281 (N_22281,N_22107,N_22116);
or U22282 (N_22282,N_22082,N_22118);
nor U22283 (N_22283,N_22044,N_22153);
xnor U22284 (N_22284,N_22115,N_22094);
or U22285 (N_22285,N_22105,N_22070);
nand U22286 (N_22286,N_22242,N_22244);
or U22287 (N_22287,N_22057,N_22184);
or U22288 (N_22288,N_22229,N_22234);
xnor U22289 (N_22289,N_22095,N_22236);
xnor U22290 (N_22290,N_22133,N_22136);
and U22291 (N_22291,N_22204,N_22016);
or U22292 (N_22292,N_22199,N_22213);
xor U22293 (N_22293,N_22218,N_22002);
and U22294 (N_22294,N_22238,N_22164);
and U22295 (N_22295,N_22060,N_22009);
and U22296 (N_22296,N_22167,N_22225);
or U22297 (N_22297,N_22012,N_22114);
and U22298 (N_22298,N_22232,N_22059);
nor U22299 (N_22299,N_22126,N_22195);
and U22300 (N_22300,N_22011,N_22022);
nand U22301 (N_22301,N_22145,N_22162);
xnor U22302 (N_22302,N_22035,N_22158);
xor U22303 (N_22303,N_22020,N_22018);
xor U22304 (N_22304,N_22055,N_22178);
xor U22305 (N_22305,N_22005,N_22243);
nand U22306 (N_22306,N_22074,N_22138);
nand U22307 (N_22307,N_22048,N_22027);
and U22308 (N_22308,N_22183,N_22121);
nand U22309 (N_22309,N_22191,N_22100);
nor U22310 (N_22310,N_22200,N_22175);
nor U22311 (N_22311,N_22036,N_22142);
nand U22312 (N_22312,N_22052,N_22154);
xnor U22313 (N_22313,N_22104,N_22098);
and U22314 (N_22314,N_22143,N_22090);
or U22315 (N_22315,N_22034,N_22102);
or U22316 (N_22316,N_22039,N_22028);
xor U22317 (N_22317,N_22174,N_22014);
nand U22318 (N_22318,N_22109,N_22023);
and U22319 (N_22319,N_22155,N_22179);
and U22320 (N_22320,N_22108,N_22206);
and U22321 (N_22321,N_22049,N_22224);
and U22322 (N_22322,N_22054,N_22066);
nor U22323 (N_22323,N_22122,N_22147);
nor U22324 (N_22324,N_22219,N_22127);
or U22325 (N_22325,N_22021,N_22026);
nand U22326 (N_22326,N_22037,N_22111);
nand U22327 (N_22327,N_22050,N_22097);
xor U22328 (N_22328,N_22144,N_22125);
or U22329 (N_22329,N_22103,N_22141);
nand U22330 (N_22330,N_22007,N_22076);
or U22331 (N_22331,N_22083,N_22077);
nor U22332 (N_22332,N_22157,N_22180);
and U22333 (N_22333,N_22013,N_22140);
or U22334 (N_22334,N_22032,N_22047);
xor U22335 (N_22335,N_22241,N_22163);
nor U22336 (N_22336,N_22119,N_22227);
and U22337 (N_22337,N_22065,N_22160);
xor U22338 (N_22338,N_22078,N_22132);
or U22339 (N_22339,N_22130,N_22113);
or U22340 (N_22340,N_22063,N_22168);
nand U22341 (N_22341,N_22176,N_22084);
and U22342 (N_22342,N_22172,N_22015);
xnor U22343 (N_22343,N_22166,N_22203);
and U22344 (N_22344,N_22053,N_22186);
nand U22345 (N_22345,N_22085,N_22120);
nand U22346 (N_22346,N_22086,N_22040);
or U22347 (N_22347,N_22081,N_22062);
nand U22348 (N_22348,N_22131,N_22051);
and U22349 (N_22349,N_22197,N_22123);
or U22350 (N_22350,N_22222,N_22117);
xnor U22351 (N_22351,N_22217,N_22149);
nor U22352 (N_22352,N_22249,N_22072);
nand U22353 (N_22353,N_22202,N_22207);
nor U22354 (N_22354,N_22106,N_22001);
and U22355 (N_22355,N_22043,N_22124);
nor U22356 (N_22356,N_22152,N_22177);
or U22357 (N_22357,N_22171,N_22017);
or U22358 (N_22358,N_22092,N_22193);
or U22359 (N_22359,N_22151,N_22112);
nor U22360 (N_22360,N_22146,N_22187);
nor U22361 (N_22361,N_22061,N_22211);
nor U22362 (N_22362,N_22029,N_22228);
nor U22363 (N_22363,N_22248,N_22003);
or U22364 (N_22364,N_22170,N_22042);
or U22365 (N_22365,N_22165,N_22045);
and U22366 (N_22366,N_22247,N_22031);
or U22367 (N_22367,N_22024,N_22205);
and U22368 (N_22368,N_22087,N_22173);
nor U22369 (N_22369,N_22223,N_22091);
xor U22370 (N_22370,N_22192,N_22019);
nor U22371 (N_22371,N_22210,N_22099);
nand U22372 (N_22372,N_22068,N_22025);
xor U22373 (N_22373,N_22148,N_22240);
nor U22374 (N_22374,N_22080,N_22135);
xor U22375 (N_22375,N_22209,N_22247);
nand U22376 (N_22376,N_22111,N_22114);
nor U22377 (N_22377,N_22060,N_22242);
and U22378 (N_22378,N_22168,N_22237);
and U22379 (N_22379,N_22164,N_22117);
nor U22380 (N_22380,N_22057,N_22072);
and U22381 (N_22381,N_22125,N_22197);
nand U22382 (N_22382,N_22201,N_22064);
nand U22383 (N_22383,N_22007,N_22004);
or U22384 (N_22384,N_22080,N_22106);
nor U22385 (N_22385,N_22242,N_22206);
nand U22386 (N_22386,N_22245,N_22199);
nor U22387 (N_22387,N_22201,N_22142);
nor U22388 (N_22388,N_22247,N_22213);
nand U22389 (N_22389,N_22086,N_22178);
xnor U22390 (N_22390,N_22175,N_22223);
xnor U22391 (N_22391,N_22070,N_22201);
and U22392 (N_22392,N_22022,N_22058);
nor U22393 (N_22393,N_22004,N_22225);
nand U22394 (N_22394,N_22249,N_22094);
nor U22395 (N_22395,N_22128,N_22003);
xnor U22396 (N_22396,N_22062,N_22108);
and U22397 (N_22397,N_22222,N_22178);
nor U22398 (N_22398,N_22209,N_22139);
or U22399 (N_22399,N_22215,N_22181);
nand U22400 (N_22400,N_22196,N_22053);
and U22401 (N_22401,N_22221,N_22029);
xor U22402 (N_22402,N_22071,N_22156);
nor U22403 (N_22403,N_22190,N_22204);
nor U22404 (N_22404,N_22036,N_22019);
nand U22405 (N_22405,N_22188,N_22040);
nand U22406 (N_22406,N_22101,N_22214);
or U22407 (N_22407,N_22059,N_22111);
nor U22408 (N_22408,N_22207,N_22100);
or U22409 (N_22409,N_22182,N_22093);
and U22410 (N_22410,N_22000,N_22127);
and U22411 (N_22411,N_22037,N_22242);
xnor U22412 (N_22412,N_22221,N_22210);
and U22413 (N_22413,N_22138,N_22197);
nand U22414 (N_22414,N_22224,N_22029);
xnor U22415 (N_22415,N_22101,N_22173);
nor U22416 (N_22416,N_22196,N_22120);
nor U22417 (N_22417,N_22046,N_22234);
nand U22418 (N_22418,N_22173,N_22150);
xor U22419 (N_22419,N_22235,N_22071);
and U22420 (N_22420,N_22234,N_22043);
and U22421 (N_22421,N_22197,N_22060);
nand U22422 (N_22422,N_22030,N_22045);
or U22423 (N_22423,N_22247,N_22052);
nand U22424 (N_22424,N_22195,N_22037);
or U22425 (N_22425,N_22132,N_22041);
or U22426 (N_22426,N_22085,N_22050);
nand U22427 (N_22427,N_22224,N_22167);
nand U22428 (N_22428,N_22210,N_22230);
nor U22429 (N_22429,N_22237,N_22204);
xor U22430 (N_22430,N_22065,N_22151);
nand U22431 (N_22431,N_22105,N_22060);
and U22432 (N_22432,N_22141,N_22034);
nor U22433 (N_22433,N_22074,N_22226);
nor U22434 (N_22434,N_22154,N_22193);
nand U22435 (N_22435,N_22097,N_22072);
or U22436 (N_22436,N_22134,N_22142);
nor U22437 (N_22437,N_22208,N_22102);
nor U22438 (N_22438,N_22117,N_22198);
nor U22439 (N_22439,N_22225,N_22234);
nor U22440 (N_22440,N_22016,N_22103);
nor U22441 (N_22441,N_22120,N_22122);
and U22442 (N_22442,N_22006,N_22033);
nor U22443 (N_22443,N_22209,N_22074);
and U22444 (N_22444,N_22248,N_22208);
xnor U22445 (N_22445,N_22057,N_22167);
xnor U22446 (N_22446,N_22173,N_22056);
nor U22447 (N_22447,N_22053,N_22241);
nor U22448 (N_22448,N_22189,N_22127);
nor U22449 (N_22449,N_22122,N_22201);
and U22450 (N_22450,N_22156,N_22005);
nor U22451 (N_22451,N_22111,N_22014);
nor U22452 (N_22452,N_22201,N_22014);
or U22453 (N_22453,N_22014,N_22044);
and U22454 (N_22454,N_22006,N_22236);
or U22455 (N_22455,N_22040,N_22105);
nand U22456 (N_22456,N_22091,N_22248);
xnor U22457 (N_22457,N_22236,N_22007);
nand U22458 (N_22458,N_22116,N_22190);
xor U22459 (N_22459,N_22031,N_22231);
and U22460 (N_22460,N_22169,N_22148);
xor U22461 (N_22461,N_22238,N_22186);
and U22462 (N_22462,N_22158,N_22248);
nand U22463 (N_22463,N_22002,N_22140);
nor U22464 (N_22464,N_22070,N_22159);
and U22465 (N_22465,N_22137,N_22157);
or U22466 (N_22466,N_22210,N_22156);
xor U22467 (N_22467,N_22187,N_22082);
nor U22468 (N_22468,N_22229,N_22174);
and U22469 (N_22469,N_22149,N_22209);
or U22470 (N_22470,N_22056,N_22092);
nor U22471 (N_22471,N_22151,N_22084);
and U22472 (N_22472,N_22054,N_22069);
xor U22473 (N_22473,N_22019,N_22043);
nand U22474 (N_22474,N_22124,N_22085);
nor U22475 (N_22475,N_22078,N_22125);
xor U22476 (N_22476,N_22081,N_22002);
xor U22477 (N_22477,N_22118,N_22175);
nor U22478 (N_22478,N_22209,N_22193);
and U22479 (N_22479,N_22115,N_22216);
xor U22480 (N_22480,N_22090,N_22220);
and U22481 (N_22481,N_22076,N_22210);
nor U22482 (N_22482,N_22085,N_22220);
nand U22483 (N_22483,N_22090,N_22080);
or U22484 (N_22484,N_22151,N_22005);
and U22485 (N_22485,N_22124,N_22062);
nand U22486 (N_22486,N_22166,N_22122);
xnor U22487 (N_22487,N_22100,N_22184);
xor U22488 (N_22488,N_22020,N_22241);
nand U22489 (N_22489,N_22083,N_22148);
or U22490 (N_22490,N_22071,N_22237);
or U22491 (N_22491,N_22148,N_22087);
or U22492 (N_22492,N_22235,N_22047);
nand U22493 (N_22493,N_22126,N_22059);
xnor U22494 (N_22494,N_22050,N_22227);
or U22495 (N_22495,N_22079,N_22170);
xnor U22496 (N_22496,N_22208,N_22204);
nand U22497 (N_22497,N_22222,N_22106);
nand U22498 (N_22498,N_22128,N_22135);
and U22499 (N_22499,N_22139,N_22071);
or U22500 (N_22500,N_22283,N_22335);
nor U22501 (N_22501,N_22311,N_22350);
nor U22502 (N_22502,N_22323,N_22264);
and U22503 (N_22503,N_22392,N_22442);
nand U22504 (N_22504,N_22255,N_22312);
and U22505 (N_22505,N_22358,N_22262);
nor U22506 (N_22506,N_22489,N_22338);
and U22507 (N_22507,N_22415,N_22368);
or U22508 (N_22508,N_22417,N_22495);
nor U22509 (N_22509,N_22393,N_22270);
or U22510 (N_22510,N_22397,N_22492);
xor U22511 (N_22511,N_22276,N_22253);
xor U22512 (N_22512,N_22403,N_22294);
or U22513 (N_22513,N_22362,N_22346);
nor U22514 (N_22514,N_22325,N_22268);
nand U22515 (N_22515,N_22469,N_22260);
xor U22516 (N_22516,N_22376,N_22271);
and U22517 (N_22517,N_22466,N_22386);
nor U22518 (N_22518,N_22378,N_22394);
nand U22519 (N_22519,N_22465,N_22257);
nor U22520 (N_22520,N_22296,N_22360);
or U22521 (N_22521,N_22331,N_22491);
nor U22522 (N_22522,N_22425,N_22298);
and U22523 (N_22523,N_22412,N_22457);
nor U22524 (N_22524,N_22423,N_22478);
and U22525 (N_22525,N_22309,N_22313);
nand U22526 (N_22526,N_22322,N_22290);
nor U22527 (N_22527,N_22250,N_22314);
xnor U22528 (N_22528,N_22432,N_22259);
or U22529 (N_22529,N_22382,N_22407);
or U22530 (N_22530,N_22494,N_22333);
nor U22531 (N_22531,N_22419,N_22327);
nor U22532 (N_22532,N_22473,N_22299);
and U22533 (N_22533,N_22266,N_22414);
and U22534 (N_22534,N_22352,N_22275);
xor U22535 (N_22535,N_22440,N_22406);
xor U22536 (N_22536,N_22361,N_22474);
nand U22537 (N_22537,N_22453,N_22458);
nor U22538 (N_22538,N_22301,N_22287);
or U22539 (N_22539,N_22450,N_22499);
xnor U22540 (N_22540,N_22345,N_22355);
nand U22541 (N_22541,N_22344,N_22289);
nor U22542 (N_22542,N_22436,N_22349);
nor U22543 (N_22543,N_22404,N_22421);
nand U22544 (N_22544,N_22405,N_22359);
or U22545 (N_22545,N_22459,N_22303);
nand U22546 (N_22546,N_22334,N_22449);
nor U22547 (N_22547,N_22348,N_22429);
nand U22548 (N_22548,N_22461,N_22373);
xor U22549 (N_22549,N_22263,N_22278);
and U22550 (N_22550,N_22326,N_22497);
nor U22551 (N_22551,N_22291,N_22252);
xnor U22552 (N_22552,N_22488,N_22402);
nor U22553 (N_22553,N_22433,N_22475);
nand U22554 (N_22554,N_22487,N_22439);
or U22555 (N_22555,N_22413,N_22267);
nor U22556 (N_22556,N_22293,N_22330);
or U22557 (N_22557,N_22416,N_22424);
and U22558 (N_22558,N_22265,N_22353);
nand U22559 (N_22559,N_22365,N_22445);
xnor U22560 (N_22560,N_22482,N_22347);
xnor U22561 (N_22561,N_22396,N_22258);
or U22562 (N_22562,N_22277,N_22329);
nand U22563 (N_22563,N_22464,N_22448);
or U22564 (N_22564,N_22357,N_22336);
and U22565 (N_22565,N_22374,N_22462);
nand U22566 (N_22566,N_22295,N_22320);
nor U22567 (N_22567,N_22444,N_22454);
nor U22568 (N_22568,N_22384,N_22390);
nor U22569 (N_22569,N_22381,N_22281);
nor U22570 (N_22570,N_22480,N_22292);
nor U22571 (N_22571,N_22446,N_22471);
nor U22572 (N_22572,N_22460,N_22430);
xnor U22573 (N_22573,N_22318,N_22304);
nand U22574 (N_22574,N_22317,N_22443);
nor U22575 (N_22575,N_22274,N_22387);
and U22576 (N_22576,N_22498,N_22251);
nor U22577 (N_22577,N_22485,N_22256);
or U22578 (N_22578,N_22308,N_22410);
or U22579 (N_22579,N_22305,N_22385);
xnor U22580 (N_22580,N_22426,N_22339);
xor U22581 (N_22581,N_22422,N_22437);
or U22582 (N_22582,N_22310,N_22493);
xor U22583 (N_22583,N_22370,N_22435);
xor U22584 (N_22584,N_22332,N_22398);
xnor U22585 (N_22585,N_22254,N_22395);
or U22586 (N_22586,N_22328,N_22476);
or U22587 (N_22587,N_22284,N_22288);
xnor U22588 (N_22588,N_22315,N_22383);
nand U22589 (N_22589,N_22316,N_22452);
nor U22590 (N_22590,N_22297,N_22367);
nand U22591 (N_22591,N_22377,N_22472);
xnor U22592 (N_22592,N_22371,N_22486);
and U22593 (N_22593,N_22428,N_22272);
nand U22594 (N_22594,N_22434,N_22490);
or U22595 (N_22595,N_22427,N_22441);
nand U22596 (N_22596,N_22401,N_22399);
nor U22597 (N_22597,N_22282,N_22463);
nand U22598 (N_22598,N_22340,N_22468);
nand U22599 (N_22599,N_22341,N_22455);
and U22600 (N_22600,N_22389,N_22481);
xor U22601 (N_22601,N_22321,N_22369);
nor U22602 (N_22602,N_22456,N_22380);
or U22603 (N_22603,N_22363,N_22375);
nor U22604 (N_22604,N_22409,N_22496);
and U22605 (N_22605,N_22342,N_22319);
xnor U22606 (N_22606,N_22354,N_22470);
xor U22607 (N_22607,N_22351,N_22286);
or U22608 (N_22608,N_22408,N_22261);
and U22609 (N_22609,N_22479,N_22477);
and U22610 (N_22610,N_22356,N_22431);
nand U22611 (N_22611,N_22366,N_22343);
nor U22612 (N_22612,N_22438,N_22400);
xor U22613 (N_22613,N_22300,N_22273);
nor U22614 (N_22614,N_22484,N_22467);
and U22615 (N_22615,N_22324,N_22420);
or U22616 (N_22616,N_22447,N_22418);
and U22617 (N_22617,N_22451,N_22306);
nor U22618 (N_22618,N_22364,N_22302);
and U22619 (N_22619,N_22269,N_22285);
or U22620 (N_22620,N_22379,N_22483);
nand U22621 (N_22621,N_22391,N_22279);
xor U22622 (N_22622,N_22411,N_22372);
nor U22623 (N_22623,N_22307,N_22388);
nor U22624 (N_22624,N_22280,N_22337);
and U22625 (N_22625,N_22263,N_22250);
xor U22626 (N_22626,N_22396,N_22278);
xnor U22627 (N_22627,N_22311,N_22353);
nand U22628 (N_22628,N_22376,N_22465);
or U22629 (N_22629,N_22430,N_22269);
and U22630 (N_22630,N_22265,N_22362);
or U22631 (N_22631,N_22305,N_22328);
nor U22632 (N_22632,N_22377,N_22445);
xnor U22633 (N_22633,N_22386,N_22298);
xnor U22634 (N_22634,N_22407,N_22400);
nand U22635 (N_22635,N_22481,N_22327);
xnor U22636 (N_22636,N_22252,N_22484);
or U22637 (N_22637,N_22432,N_22433);
xnor U22638 (N_22638,N_22477,N_22490);
xnor U22639 (N_22639,N_22404,N_22437);
or U22640 (N_22640,N_22361,N_22425);
nand U22641 (N_22641,N_22336,N_22447);
or U22642 (N_22642,N_22265,N_22447);
xor U22643 (N_22643,N_22293,N_22351);
nand U22644 (N_22644,N_22357,N_22416);
nor U22645 (N_22645,N_22295,N_22372);
or U22646 (N_22646,N_22362,N_22259);
and U22647 (N_22647,N_22358,N_22368);
or U22648 (N_22648,N_22455,N_22499);
nand U22649 (N_22649,N_22273,N_22252);
nor U22650 (N_22650,N_22302,N_22440);
or U22651 (N_22651,N_22298,N_22390);
or U22652 (N_22652,N_22400,N_22395);
nor U22653 (N_22653,N_22393,N_22312);
xor U22654 (N_22654,N_22442,N_22255);
nor U22655 (N_22655,N_22417,N_22361);
or U22656 (N_22656,N_22464,N_22316);
nor U22657 (N_22657,N_22386,N_22258);
or U22658 (N_22658,N_22409,N_22435);
or U22659 (N_22659,N_22461,N_22420);
xor U22660 (N_22660,N_22348,N_22320);
nor U22661 (N_22661,N_22262,N_22455);
or U22662 (N_22662,N_22496,N_22323);
nand U22663 (N_22663,N_22389,N_22499);
nor U22664 (N_22664,N_22313,N_22461);
and U22665 (N_22665,N_22397,N_22289);
xnor U22666 (N_22666,N_22291,N_22267);
xnor U22667 (N_22667,N_22495,N_22344);
and U22668 (N_22668,N_22414,N_22442);
nand U22669 (N_22669,N_22415,N_22443);
nand U22670 (N_22670,N_22484,N_22381);
or U22671 (N_22671,N_22263,N_22406);
nor U22672 (N_22672,N_22348,N_22321);
and U22673 (N_22673,N_22368,N_22319);
xor U22674 (N_22674,N_22433,N_22290);
nor U22675 (N_22675,N_22449,N_22405);
xnor U22676 (N_22676,N_22310,N_22250);
or U22677 (N_22677,N_22350,N_22457);
xnor U22678 (N_22678,N_22462,N_22322);
nor U22679 (N_22679,N_22375,N_22301);
and U22680 (N_22680,N_22410,N_22258);
xor U22681 (N_22681,N_22335,N_22324);
nor U22682 (N_22682,N_22306,N_22313);
xor U22683 (N_22683,N_22276,N_22273);
xor U22684 (N_22684,N_22458,N_22311);
xnor U22685 (N_22685,N_22367,N_22364);
nand U22686 (N_22686,N_22432,N_22423);
and U22687 (N_22687,N_22357,N_22319);
and U22688 (N_22688,N_22313,N_22459);
xor U22689 (N_22689,N_22373,N_22290);
nor U22690 (N_22690,N_22380,N_22275);
or U22691 (N_22691,N_22281,N_22444);
nor U22692 (N_22692,N_22300,N_22354);
nor U22693 (N_22693,N_22315,N_22380);
xor U22694 (N_22694,N_22321,N_22316);
xor U22695 (N_22695,N_22426,N_22370);
xor U22696 (N_22696,N_22486,N_22488);
or U22697 (N_22697,N_22478,N_22376);
xnor U22698 (N_22698,N_22404,N_22411);
or U22699 (N_22699,N_22257,N_22484);
nor U22700 (N_22700,N_22367,N_22342);
nand U22701 (N_22701,N_22368,N_22442);
xor U22702 (N_22702,N_22462,N_22415);
xor U22703 (N_22703,N_22462,N_22297);
and U22704 (N_22704,N_22490,N_22254);
and U22705 (N_22705,N_22440,N_22493);
xnor U22706 (N_22706,N_22333,N_22374);
and U22707 (N_22707,N_22386,N_22446);
and U22708 (N_22708,N_22478,N_22278);
nand U22709 (N_22709,N_22259,N_22439);
nand U22710 (N_22710,N_22444,N_22374);
nand U22711 (N_22711,N_22270,N_22390);
nor U22712 (N_22712,N_22450,N_22455);
and U22713 (N_22713,N_22421,N_22496);
xnor U22714 (N_22714,N_22366,N_22348);
nor U22715 (N_22715,N_22316,N_22338);
and U22716 (N_22716,N_22275,N_22357);
nor U22717 (N_22717,N_22368,N_22265);
nand U22718 (N_22718,N_22262,N_22438);
xnor U22719 (N_22719,N_22426,N_22329);
nand U22720 (N_22720,N_22266,N_22321);
and U22721 (N_22721,N_22481,N_22414);
and U22722 (N_22722,N_22478,N_22389);
and U22723 (N_22723,N_22256,N_22334);
nor U22724 (N_22724,N_22499,N_22315);
and U22725 (N_22725,N_22420,N_22292);
and U22726 (N_22726,N_22320,N_22466);
nand U22727 (N_22727,N_22309,N_22451);
and U22728 (N_22728,N_22376,N_22370);
and U22729 (N_22729,N_22376,N_22461);
nand U22730 (N_22730,N_22415,N_22414);
nor U22731 (N_22731,N_22320,N_22451);
nand U22732 (N_22732,N_22336,N_22463);
and U22733 (N_22733,N_22319,N_22376);
nor U22734 (N_22734,N_22266,N_22412);
and U22735 (N_22735,N_22485,N_22331);
and U22736 (N_22736,N_22364,N_22359);
xor U22737 (N_22737,N_22400,N_22455);
nor U22738 (N_22738,N_22287,N_22352);
and U22739 (N_22739,N_22342,N_22315);
xor U22740 (N_22740,N_22349,N_22378);
nor U22741 (N_22741,N_22397,N_22272);
nor U22742 (N_22742,N_22266,N_22455);
and U22743 (N_22743,N_22343,N_22315);
and U22744 (N_22744,N_22421,N_22499);
and U22745 (N_22745,N_22274,N_22467);
nand U22746 (N_22746,N_22298,N_22474);
nor U22747 (N_22747,N_22456,N_22266);
and U22748 (N_22748,N_22260,N_22303);
nand U22749 (N_22749,N_22353,N_22451);
and U22750 (N_22750,N_22677,N_22623);
xor U22751 (N_22751,N_22566,N_22564);
or U22752 (N_22752,N_22545,N_22698);
nand U22753 (N_22753,N_22611,N_22636);
and U22754 (N_22754,N_22620,N_22655);
xnor U22755 (N_22755,N_22509,N_22678);
xnor U22756 (N_22756,N_22514,N_22745);
xor U22757 (N_22757,N_22653,N_22553);
nand U22758 (N_22758,N_22634,N_22574);
and U22759 (N_22759,N_22664,N_22739);
nand U22760 (N_22760,N_22712,N_22546);
xor U22761 (N_22761,N_22530,N_22560);
or U22762 (N_22762,N_22749,N_22585);
and U22763 (N_22763,N_22502,N_22697);
xnor U22764 (N_22764,N_22531,N_22676);
or U22765 (N_22765,N_22688,N_22729);
and U22766 (N_22766,N_22621,N_22744);
nand U22767 (N_22767,N_22507,N_22670);
and U22768 (N_22768,N_22733,N_22635);
and U22769 (N_22769,N_22607,N_22715);
xor U22770 (N_22770,N_22646,N_22569);
nand U22771 (N_22771,N_22647,N_22624);
or U22772 (N_22772,N_22660,N_22556);
nor U22773 (N_22773,N_22552,N_22680);
or U22774 (N_22774,N_22673,N_22510);
xor U22775 (N_22775,N_22605,N_22734);
or U22776 (N_22776,N_22652,N_22631);
or U22777 (N_22777,N_22604,N_22747);
nand U22778 (N_22778,N_22666,N_22533);
and U22779 (N_22779,N_22736,N_22645);
xnor U22780 (N_22780,N_22682,N_22668);
xnor U22781 (N_22781,N_22633,N_22591);
or U22782 (N_22782,N_22526,N_22637);
and U22783 (N_22783,N_22724,N_22542);
or U22784 (N_22784,N_22656,N_22743);
nor U22785 (N_22785,N_22639,N_22681);
and U22786 (N_22786,N_22588,N_22707);
nor U22787 (N_22787,N_22568,N_22628);
nor U22788 (N_22788,N_22713,N_22551);
and U22789 (N_22789,N_22596,N_22741);
nand U22790 (N_22790,N_22732,N_22549);
nand U22791 (N_22791,N_22695,N_22609);
nor U22792 (N_22792,N_22521,N_22717);
nand U22793 (N_22793,N_22738,N_22718);
xnor U22794 (N_22794,N_22706,N_22561);
and U22795 (N_22795,N_22559,N_22650);
and U22796 (N_22796,N_22524,N_22513);
xnor U22797 (N_22797,N_22506,N_22601);
nor U22798 (N_22798,N_22685,N_22599);
or U22799 (N_22799,N_22689,N_22534);
xor U22800 (N_22800,N_22548,N_22555);
nand U22801 (N_22801,N_22711,N_22722);
and U22802 (N_22802,N_22539,N_22577);
nor U22803 (N_22803,N_22583,N_22716);
nand U22804 (N_22804,N_22598,N_22723);
xnor U22805 (N_22805,N_22538,N_22541);
and U22806 (N_22806,N_22587,N_22504);
or U22807 (N_22807,N_22579,N_22576);
xnor U22808 (N_22808,N_22573,N_22675);
nand U22809 (N_22809,N_22616,N_22694);
and U22810 (N_22810,N_22626,N_22501);
nand U22811 (N_22811,N_22575,N_22699);
and U22812 (N_22812,N_22567,N_22649);
xor U22813 (N_22813,N_22589,N_22705);
nand U22814 (N_22814,N_22525,N_22667);
xor U22815 (N_22815,N_22684,N_22565);
and U22816 (N_22816,N_22544,N_22529);
xor U22817 (N_22817,N_22537,N_22594);
or U22818 (N_22818,N_22570,N_22704);
nand U22819 (N_22819,N_22610,N_22580);
nor U22820 (N_22820,N_22586,N_22557);
nor U22821 (N_22821,N_22571,N_22679);
nor U22822 (N_22822,N_22550,N_22721);
and U22823 (N_22823,N_22687,N_22593);
nor U22824 (N_22824,N_22674,N_22701);
nor U22825 (N_22825,N_22516,N_22627);
nand U22826 (N_22826,N_22630,N_22662);
xor U22827 (N_22827,N_22584,N_22746);
nor U22828 (N_22828,N_22617,N_22527);
nor U22829 (N_22829,N_22505,N_22597);
nor U22830 (N_22830,N_22719,N_22671);
nor U22831 (N_22831,N_22508,N_22519);
nor U22832 (N_22832,N_22562,N_22641);
or U22833 (N_22833,N_22517,N_22731);
nor U22834 (N_22834,N_22710,N_22727);
and U22835 (N_22835,N_22692,N_22737);
or U22836 (N_22836,N_22500,N_22512);
nand U22837 (N_22837,N_22700,N_22686);
xnor U22838 (N_22838,N_22658,N_22726);
nor U22839 (N_22839,N_22563,N_22643);
or U22840 (N_22840,N_22742,N_22654);
nor U22841 (N_22841,N_22618,N_22523);
and U22842 (N_22842,N_22522,N_22572);
xnor U22843 (N_22843,N_22615,N_22638);
nor U22844 (N_22844,N_22582,N_22690);
or U22845 (N_22845,N_22740,N_22536);
or U22846 (N_22846,N_22613,N_22600);
or U22847 (N_22847,N_22648,N_22590);
and U22848 (N_22848,N_22532,N_22728);
and U22849 (N_22849,N_22625,N_22503);
nor U22850 (N_22850,N_22543,N_22693);
nand U22851 (N_22851,N_22720,N_22603);
xor U22852 (N_22852,N_22657,N_22554);
and U22853 (N_22853,N_22709,N_22608);
xnor U22854 (N_22854,N_22629,N_22661);
and U22855 (N_22855,N_22592,N_22602);
nor U22856 (N_22856,N_22702,N_22595);
xnor U22857 (N_22857,N_22578,N_22606);
nand U22858 (N_22858,N_22651,N_22683);
nor U22859 (N_22859,N_22528,N_22640);
xor U22860 (N_22860,N_22665,N_22691);
or U22861 (N_22861,N_22511,N_22540);
nor U22862 (N_22862,N_22714,N_22725);
or U22863 (N_22863,N_22558,N_22735);
nor U22864 (N_22864,N_22644,N_22581);
nand U22865 (N_22865,N_22730,N_22619);
xnor U22866 (N_22866,N_22703,N_22708);
nor U22867 (N_22867,N_22632,N_22663);
xnor U22868 (N_22868,N_22547,N_22642);
or U22869 (N_22869,N_22515,N_22669);
nand U22870 (N_22870,N_22622,N_22748);
nor U22871 (N_22871,N_22672,N_22535);
and U22872 (N_22872,N_22696,N_22614);
nor U22873 (N_22873,N_22518,N_22612);
and U22874 (N_22874,N_22659,N_22520);
nand U22875 (N_22875,N_22643,N_22693);
nor U22876 (N_22876,N_22500,N_22585);
nand U22877 (N_22877,N_22734,N_22620);
nand U22878 (N_22878,N_22656,N_22645);
or U22879 (N_22879,N_22632,N_22575);
and U22880 (N_22880,N_22664,N_22681);
xnor U22881 (N_22881,N_22624,N_22728);
or U22882 (N_22882,N_22679,N_22637);
or U22883 (N_22883,N_22652,N_22594);
xor U22884 (N_22884,N_22614,N_22506);
and U22885 (N_22885,N_22508,N_22674);
and U22886 (N_22886,N_22561,N_22522);
xor U22887 (N_22887,N_22563,N_22713);
nor U22888 (N_22888,N_22554,N_22542);
and U22889 (N_22889,N_22531,N_22714);
and U22890 (N_22890,N_22531,N_22524);
nor U22891 (N_22891,N_22694,N_22641);
nor U22892 (N_22892,N_22747,N_22628);
nor U22893 (N_22893,N_22629,N_22719);
nor U22894 (N_22894,N_22669,N_22641);
nor U22895 (N_22895,N_22537,N_22540);
nor U22896 (N_22896,N_22702,N_22693);
xor U22897 (N_22897,N_22599,N_22547);
or U22898 (N_22898,N_22602,N_22619);
nor U22899 (N_22899,N_22532,N_22517);
and U22900 (N_22900,N_22717,N_22577);
nand U22901 (N_22901,N_22716,N_22549);
nand U22902 (N_22902,N_22511,N_22679);
and U22903 (N_22903,N_22588,N_22730);
and U22904 (N_22904,N_22704,N_22723);
nor U22905 (N_22905,N_22679,N_22715);
xnor U22906 (N_22906,N_22592,N_22528);
or U22907 (N_22907,N_22626,N_22630);
and U22908 (N_22908,N_22668,N_22632);
and U22909 (N_22909,N_22547,N_22654);
nand U22910 (N_22910,N_22629,N_22567);
nand U22911 (N_22911,N_22650,N_22652);
nor U22912 (N_22912,N_22731,N_22543);
or U22913 (N_22913,N_22540,N_22722);
nand U22914 (N_22914,N_22612,N_22580);
nor U22915 (N_22915,N_22632,N_22694);
xor U22916 (N_22916,N_22625,N_22694);
xnor U22917 (N_22917,N_22747,N_22637);
nand U22918 (N_22918,N_22575,N_22709);
and U22919 (N_22919,N_22710,N_22620);
or U22920 (N_22920,N_22563,N_22700);
nand U22921 (N_22921,N_22505,N_22683);
nand U22922 (N_22922,N_22574,N_22589);
and U22923 (N_22923,N_22550,N_22525);
and U22924 (N_22924,N_22685,N_22673);
nor U22925 (N_22925,N_22607,N_22588);
or U22926 (N_22926,N_22545,N_22550);
xnor U22927 (N_22927,N_22540,N_22703);
and U22928 (N_22928,N_22677,N_22663);
xor U22929 (N_22929,N_22565,N_22528);
and U22930 (N_22930,N_22628,N_22715);
or U22931 (N_22931,N_22544,N_22714);
xor U22932 (N_22932,N_22552,N_22695);
nor U22933 (N_22933,N_22520,N_22516);
nor U22934 (N_22934,N_22612,N_22620);
nand U22935 (N_22935,N_22661,N_22704);
or U22936 (N_22936,N_22616,N_22515);
nand U22937 (N_22937,N_22610,N_22547);
nand U22938 (N_22938,N_22622,N_22658);
nor U22939 (N_22939,N_22620,N_22745);
xor U22940 (N_22940,N_22696,N_22535);
nor U22941 (N_22941,N_22681,N_22561);
nor U22942 (N_22942,N_22599,N_22502);
nor U22943 (N_22943,N_22667,N_22572);
or U22944 (N_22944,N_22511,N_22618);
nand U22945 (N_22945,N_22559,N_22686);
nand U22946 (N_22946,N_22628,N_22668);
nor U22947 (N_22947,N_22715,N_22504);
nand U22948 (N_22948,N_22544,N_22538);
or U22949 (N_22949,N_22542,N_22670);
and U22950 (N_22950,N_22511,N_22663);
xor U22951 (N_22951,N_22553,N_22538);
and U22952 (N_22952,N_22740,N_22696);
xnor U22953 (N_22953,N_22532,N_22715);
nor U22954 (N_22954,N_22539,N_22509);
xor U22955 (N_22955,N_22589,N_22596);
and U22956 (N_22956,N_22742,N_22730);
nand U22957 (N_22957,N_22501,N_22519);
nor U22958 (N_22958,N_22618,N_22509);
nand U22959 (N_22959,N_22732,N_22617);
and U22960 (N_22960,N_22580,N_22684);
or U22961 (N_22961,N_22501,N_22609);
nand U22962 (N_22962,N_22645,N_22717);
xnor U22963 (N_22963,N_22651,N_22706);
nand U22964 (N_22964,N_22692,N_22733);
nor U22965 (N_22965,N_22724,N_22689);
and U22966 (N_22966,N_22507,N_22608);
nor U22967 (N_22967,N_22738,N_22522);
nand U22968 (N_22968,N_22724,N_22723);
nand U22969 (N_22969,N_22567,N_22579);
nor U22970 (N_22970,N_22700,N_22642);
nand U22971 (N_22971,N_22598,N_22576);
nand U22972 (N_22972,N_22679,N_22561);
xnor U22973 (N_22973,N_22522,N_22585);
xnor U22974 (N_22974,N_22636,N_22666);
or U22975 (N_22975,N_22610,N_22618);
nor U22976 (N_22976,N_22559,N_22548);
and U22977 (N_22977,N_22611,N_22728);
and U22978 (N_22978,N_22663,N_22713);
or U22979 (N_22979,N_22579,N_22666);
or U22980 (N_22980,N_22562,N_22521);
nand U22981 (N_22981,N_22594,N_22581);
or U22982 (N_22982,N_22684,N_22682);
and U22983 (N_22983,N_22505,N_22682);
nand U22984 (N_22984,N_22615,N_22544);
nor U22985 (N_22985,N_22745,N_22649);
or U22986 (N_22986,N_22711,N_22526);
or U22987 (N_22987,N_22503,N_22601);
xnor U22988 (N_22988,N_22538,N_22649);
xor U22989 (N_22989,N_22540,N_22748);
nand U22990 (N_22990,N_22655,N_22549);
nor U22991 (N_22991,N_22708,N_22637);
and U22992 (N_22992,N_22661,N_22715);
and U22993 (N_22993,N_22672,N_22606);
or U22994 (N_22994,N_22545,N_22603);
or U22995 (N_22995,N_22734,N_22603);
nor U22996 (N_22996,N_22657,N_22524);
nand U22997 (N_22997,N_22578,N_22733);
nor U22998 (N_22998,N_22681,N_22716);
xor U22999 (N_22999,N_22677,N_22619);
nor U23000 (N_23000,N_22757,N_22946);
xnor U23001 (N_23001,N_22927,N_22920);
or U23002 (N_23002,N_22949,N_22984);
nand U23003 (N_23003,N_22762,N_22846);
xnor U23004 (N_23004,N_22780,N_22853);
or U23005 (N_23005,N_22855,N_22849);
nor U23006 (N_23006,N_22941,N_22923);
nand U23007 (N_23007,N_22957,N_22843);
nor U23008 (N_23008,N_22773,N_22886);
and U23009 (N_23009,N_22814,N_22758);
nor U23010 (N_23010,N_22820,N_22863);
nand U23011 (N_23011,N_22996,N_22935);
nor U23012 (N_23012,N_22854,N_22896);
and U23013 (N_23013,N_22959,N_22830);
and U23014 (N_23014,N_22789,N_22982);
xnor U23015 (N_23015,N_22848,N_22791);
xor U23016 (N_23016,N_22983,N_22822);
nand U23017 (N_23017,N_22939,N_22966);
xor U23018 (N_23018,N_22777,N_22951);
and U23019 (N_23019,N_22812,N_22911);
nand U23020 (N_23020,N_22771,N_22769);
nand U23021 (N_23021,N_22772,N_22973);
nand U23022 (N_23022,N_22766,N_22844);
or U23023 (N_23023,N_22907,N_22754);
or U23024 (N_23024,N_22816,N_22835);
nor U23025 (N_23025,N_22796,N_22914);
nand U23026 (N_23026,N_22997,N_22962);
xor U23027 (N_23027,N_22753,N_22936);
nor U23028 (N_23028,N_22770,N_22767);
nor U23029 (N_23029,N_22870,N_22768);
nor U23030 (N_23030,N_22874,N_22906);
nor U23031 (N_23031,N_22808,N_22943);
nor U23032 (N_23032,N_22991,N_22954);
and U23033 (N_23033,N_22919,N_22892);
or U23034 (N_23034,N_22894,N_22832);
xor U23035 (N_23035,N_22977,N_22929);
xor U23036 (N_23036,N_22995,N_22819);
nor U23037 (N_23037,N_22937,N_22931);
nor U23038 (N_23038,N_22987,N_22850);
nor U23039 (N_23039,N_22761,N_22904);
or U23040 (N_23040,N_22999,N_22828);
nor U23041 (N_23041,N_22833,N_22925);
nor U23042 (N_23042,N_22990,N_22787);
or U23043 (N_23043,N_22998,N_22905);
xnor U23044 (N_23044,N_22751,N_22889);
xor U23045 (N_23045,N_22798,N_22841);
and U23046 (N_23046,N_22775,N_22921);
nand U23047 (N_23047,N_22975,N_22953);
or U23048 (N_23048,N_22805,N_22809);
or U23049 (N_23049,N_22869,N_22898);
nor U23050 (N_23050,N_22944,N_22928);
nor U23051 (N_23051,N_22960,N_22945);
nor U23052 (N_23052,N_22794,N_22915);
nand U23053 (N_23053,N_22806,N_22795);
xnor U23054 (N_23054,N_22810,N_22948);
and U23055 (N_23055,N_22895,N_22888);
and U23056 (N_23056,N_22964,N_22778);
nor U23057 (N_23057,N_22913,N_22976);
or U23058 (N_23058,N_22799,N_22824);
nor U23059 (N_23059,N_22852,N_22882);
nor U23060 (N_23060,N_22823,N_22912);
and U23061 (N_23061,N_22755,N_22947);
nand U23062 (N_23062,N_22909,N_22858);
nor U23063 (N_23063,N_22837,N_22897);
nand U23064 (N_23064,N_22872,N_22900);
and U23065 (N_23065,N_22847,N_22986);
nand U23066 (N_23066,N_22908,N_22988);
or U23067 (N_23067,N_22783,N_22811);
or U23068 (N_23068,N_22926,N_22857);
nor U23069 (N_23069,N_22880,N_22800);
or U23070 (N_23070,N_22871,N_22968);
xor U23071 (N_23071,N_22774,N_22978);
nor U23072 (N_23072,N_22891,N_22933);
or U23073 (N_23073,N_22879,N_22902);
nand U23074 (N_23074,N_22938,N_22981);
nor U23075 (N_23075,N_22802,N_22916);
nand U23076 (N_23076,N_22950,N_22825);
nor U23077 (N_23077,N_22763,N_22776);
nor U23078 (N_23078,N_22932,N_22876);
or U23079 (N_23079,N_22952,N_22887);
nor U23080 (N_23080,N_22989,N_22890);
nor U23081 (N_23081,N_22961,N_22836);
nand U23082 (N_23082,N_22942,N_22972);
nand U23083 (N_23083,N_22985,N_22971);
and U23084 (N_23084,N_22865,N_22893);
or U23085 (N_23085,N_22862,N_22788);
nand U23086 (N_23086,N_22765,N_22881);
nor U23087 (N_23087,N_22804,N_22786);
xor U23088 (N_23088,N_22917,N_22801);
and U23089 (N_23089,N_22750,N_22845);
nand U23090 (N_23090,N_22873,N_22980);
xnor U23091 (N_23091,N_22860,N_22883);
nand U23092 (N_23092,N_22793,N_22784);
xor U23093 (N_23093,N_22979,N_22807);
nor U23094 (N_23094,N_22965,N_22930);
and U23095 (N_23095,N_22878,N_22839);
or U23096 (N_23096,N_22859,N_22956);
nor U23097 (N_23097,N_22831,N_22851);
xor U23098 (N_23098,N_22910,N_22877);
xor U23099 (N_23099,N_22970,N_22818);
and U23100 (N_23100,N_22866,N_22967);
or U23101 (N_23101,N_22992,N_22885);
nor U23102 (N_23102,N_22813,N_22759);
nor U23103 (N_23103,N_22815,N_22792);
or U23104 (N_23104,N_22868,N_22760);
and U23105 (N_23105,N_22785,N_22903);
or U23106 (N_23106,N_22834,N_22840);
and U23107 (N_23107,N_22918,N_22867);
nand U23108 (N_23108,N_22782,N_22856);
and U23109 (N_23109,N_22958,N_22817);
nor U23110 (N_23110,N_22899,N_22827);
nor U23111 (N_23111,N_22829,N_22994);
and U23112 (N_23112,N_22993,N_22790);
and U23113 (N_23113,N_22803,N_22797);
and U23114 (N_23114,N_22875,N_22969);
and U23115 (N_23115,N_22752,N_22861);
xnor U23116 (N_23116,N_22756,N_22826);
and U23117 (N_23117,N_22963,N_22821);
or U23118 (N_23118,N_22922,N_22974);
and U23119 (N_23119,N_22838,N_22781);
xor U23120 (N_23120,N_22864,N_22884);
xor U23121 (N_23121,N_22842,N_22764);
nor U23122 (N_23122,N_22924,N_22779);
xor U23123 (N_23123,N_22955,N_22940);
nor U23124 (N_23124,N_22934,N_22901);
or U23125 (N_23125,N_22774,N_22833);
or U23126 (N_23126,N_22763,N_22777);
nand U23127 (N_23127,N_22992,N_22937);
or U23128 (N_23128,N_22986,N_22966);
and U23129 (N_23129,N_22819,N_22918);
nor U23130 (N_23130,N_22875,N_22887);
xor U23131 (N_23131,N_22982,N_22936);
nor U23132 (N_23132,N_22923,N_22772);
xor U23133 (N_23133,N_22929,N_22806);
nor U23134 (N_23134,N_22787,N_22815);
xnor U23135 (N_23135,N_22790,N_22873);
xor U23136 (N_23136,N_22787,N_22998);
nand U23137 (N_23137,N_22985,N_22816);
nand U23138 (N_23138,N_22924,N_22968);
and U23139 (N_23139,N_22926,N_22789);
or U23140 (N_23140,N_22872,N_22870);
or U23141 (N_23141,N_22767,N_22986);
nand U23142 (N_23142,N_22908,N_22877);
nor U23143 (N_23143,N_22819,N_22854);
or U23144 (N_23144,N_22853,N_22877);
or U23145 (N_23145,N_22840,N_22943);
and U23146 (N_23146,N_22762,N_22912);
and U23147 (N_23147,N_22778,N_22977);
xnor U23148 (N_23148,N_22797,N_22864);
or U23149 (N_23149,N_22924,N_22950);
or U23150 (N_23150,N_22889,N_22920);
and U23151 (N_23151,N_22858,N_22870);
and U23152 (N_23152,N_22901,N_22974);
xnor U23153 (N_23153,N_22943,N_22959);
xnor U23154 (N_23154,N_22841,N_22752);
and U23155 (N_23155,N_22877,N_22925);
nand U23156 (N_23156,N_22875,N_22983);
or U23157 (N_23157,N_22801,N_22820);
or U23158 (N_23158,N_22945,N_22932);
nand U23159 (N_23159,N_22796,N_22872);
nor U23160 (N_23160,N_22797,N_22986);
or U23161 (N_23161,N_22881,N_22987);
nand U23162 (N_23162,N_22840,N_22872);
or U23163 (N_23163,N_22908,N_22831);
or U23164 (N_23164,N_22811,N_22918);
nand U23165 (N_23165,N_22991,N_22896);
or U23166 (N_23166,N_22977,N_22911);
and U23167 (N_23167,N_22823,N_22826);
nand U23168 (N_23168,N_22906,N_22825);
xor U23169 (N_23169,N_22898,N_22829);
and U23170 (N_23170,N_22928,N_22924);
nand U23171 (N_23171,N_22962,N_22936);
and U23172 (N_23172,N_22842,N_22937);
and U23173 (N_23173,N_22881,N_22785);
nand U23174 (N_23174,N_22802,N_22958);
or U23175 (N_23175,N_22835,N_22813);
or U23176 (N_23176,N_22766,N_22877);
nor U23177 (N_23177,N_22780,N_22812);
nand U23178 (N_23178,N_22945,N_22845);
nor U23179 (N_23179,N_22939,N_22921);
nor U23180 (N_23180,N_22839,N_22931);
or U23181 (N_23181,N_22896,N_22848);
xor U23182 (N_23182,N_22844,N_22775);
nand U23183 (N_23183,N_22985,N_22881);
xnor U23184 (N_23184,N_22879,N_22767);
or U23185 (N_23185,N_22768,N_22894);
nor U23186 (N_23186,N_22969,N_22775);
or U23187 (N_23187,N_22897,N_22931);
nand U23188 (N_23188,N_22822,N_22922);
or U23189 (N_23189,N_22853,N_22764);
xor U23190 (N_23190,N_22889,N_22907);
nor U23191 (N_23191,N_22821,N_22951);
xnor U23192 (N_23192,N_22922,N_22854);
or U23193 (N_23193,N_22799,N_22752);
and U23194 (N_23194,N_22977,N_22819);
nor U23195 (N_23195,N_22964,N_22956);
or U23196 (N_23196,N_22758,N_22991);
nand U23197 (N_23197,N_22862,N_22847);
nand U23198 (N_23198,N_22850,N_22832);
and U23199 (N_23199,N_22835,N_22858);
nor U23200 (N_23200,N_22930,N_22843);
xor U23201 (N_23201,N_22750,N_22869);
and U23202 (N_23202,N_22932,N_22760);
and U23203 (N_23203,N_22937,N_22954);
nand U23204 (N_23204,N_22955,N_22783);
and U23205 (N_23205,N_22880,N_22897);
xor U23206 (N_23206,N_22789,N_22823);
and U23207 (N_23207,N_22950,N_22804);
xor U23208 (N_23208,N_22890,N_22794);
and U23209 (N_23209,N_22928,N_22973);
nand U23210 (N_23210,N_22921,N_22797);
and U23211 (N_23211,N_22863,N_22996);
or U23212 (N_23212,N_22751,N_22847);
and U23213 (N_23213,N_22879,N_22972);
or U23214 (N_23214,N_22874,N_22967);
and U23215 (N_23215,N_22976,N_22933);
or U23216 (N_23216,N_22805,N_22905);
or U23217 (N_23217,N_22837,N_22925);
nand U23218 (N_23218,N_22925,N_22859);
and U23219 (N_23219,N_22758,N_22848);
nand U23220 (N_23220,N_22853,N_22940);
and U23221 (N_23221,N_22858,N_22902);
and U23222 (N_23222,N_22931,N_22915);
nor U23223 (N_23223,N_22923,N_22806);
or U23224 (N_23224,N_22933,N_22894);
and U23225 (N_23225,N_22804,N_22780);
nor U23226 (N_23226,N_22787,N_22966);
nand U23227 (N_23227,N_22770,N_22778);
nor U23228 (N_23228,N_22946,N_22802);
and U23229 (N_23229,N_22783,N_22842);
nor U23230 (N_23230,N_22915,N_22805);
nor U23231 (N_23231,N_22959,N_22920);
nand U23232 (N_23232,N_22968,N_22976);
or U23233 (N_23233,N_22836,N_22922);
and U23234 (N_23234,N_22763,N_22973);
xor U23235 (N_23235,N_22877,N_22980);
or U23236 (N_23236,N_22919,N_22950);
xnor U23237 (N_23237,N_22819,N_22889);
nor U23238 (N_23238,N_22880,N_22826);
xor U23239 (N_23239,N_22869,N_22787);
nand U23240 (N_23240,N_22906,N_22998);
and U23241 (N_23241,N_22866,N_22958);
nand U23242 (N_23242,N_22889,N_22881);
xor U23243 (N_23243,N_22800,N_22839);
nand U23244 (N_23244,N_22905,N_22973);
nand U23245 (N_23245,N_22941,N_22994);
or U23246 (N_23246,N_22881,N_22845);
xor U23247 (N_23247,N_22755,N_22929);
nand U23248 (N_23248,N_22802,N_22923);
nor U23249 (N_23249,N_22978,N_22768);
and U23250 (N_23250,N_23160,N_23162);
or U23251 (N_23251,N_23038,N_23222);
nand U23252 (N_23252,N_23243,N_23204);
or U23253 (N_23253,N_23029,N_23045);
nand U23254 (N_23254,N_23017,N_23197);
xnor U23255 (N_23255,N_23092,N_23249);
and U23256 (N_23256,N_23082,N_23156);
and U23257 (N_23257,N_23100,N_23050);
and U23258 (N_23258,N_23086,N_23219);
nand U23259 (N_23259,N_23033,N_23003);
or U23260 (N_23260,N_23142,N_23203);
and U23261 (N_23261,N_23132,N_23067);
nor U23262 (N_23262,N_23131,N_23211);
or U23263 (N_23263,N_23059,N_23168);
or U23264 (N_23264,N_23200,N_23087);
nor U23265 (N_23265,N_23034,N_23114);
and U23266 (N_23266,N_23137,N_23013);
and U23267 (N_23267,N_23036,N_23152);
nand U23268 (N_23268,N_23148,N_23216);
and U23269 (N_23269,N_23239,N_23210);
nand U23270 (N_23270,N_23058,N_23220);
nor U23271 (N_23271,N_23021,N_23169);
xor U23272 (N_23272,N_23218,N_23101);
xor U23273 (N_23273,N_23155,N_23193);
or U23274 (N_23274,N_23174,N_23069);
or U23275 (N_23275,N_23075,N_23229);
xor U23276 (N_23276,N_23042,N_23043);
and U23277 (N_23277,N_23099,N_23158);
and U23278 (N_23278,N_23238,N_23190);
nand U23279 (N_23279,N_23103,N_23061);
nor U23280 (N_23280,N_23111,N_23020);
or U23281 (N_23281,N_23235,N_23063);
and U23282 (N_23282,N_23151,N_23081);
and U23283 (N_23283,N_23171,N_23163);
or U23284 (N_23284,N_23141,N_23192);
or U23285 (N_23285,N_23157,N_23109);
nor U23286 (N_23286,N_23232,N_23196);
and U23287 (N_23287,N_23194,N_23121);
or U23288 (N_23288,N_23126,N_23140);
nor U23289 (N_23289,N_23173,N_23124);
nor U23290 (N_23290,N_23096,N_23053);
xnor U23291 (N_23291,N_23009,N_23221);
and U23292 (N_23292,N_23106,N_23236);
xnor U23293 (N_23293,N_23083,N_23031);
and U23294 (N_23294,N_23060,N_23015);
xnor U23295 (N_23295,N_23107,N_23001);
nand U23296 (N_23296,N_23000,N_23205);
nand U23297 (N_23297,N_23227,N_23198);
nor U23298 (N_23298,N_23127,N_23228);
nand U23299 (N_23299,N_23230,N_23037);
xnor U23300 (N_23300,N_23128,N_23223);
or U23301 (N_23301,N_23189,N_23165);
nor U23302 (N_23302,N_23102,N_23122);
or U23303 (N_23303,N_23054,N_23153);
and U23304 (N_23304,N_23016,N_23180);
xnor U23305 (N_23305,N_23008,N_23125);
nor U23306 (N_23306,N_23244,N_23150);
xnor U23307 (N_23307,N_23046,N_23166);
nor U23308 (N_23308,N_23185,N_23098);
or U23309 (N_23309,N_23178,N_23119);
and U23310 (N_23310,N_23242,N_23202);
xor U23311 (N_23311,N_23047,N_23110);
and U23312 (N_23312,N_23005,N_23032);
or U23313 (N_23313,N_23097,N_23146);
nor U23314 (N_23314,N_23091,N_23212);
or U23315 (N_23315,N_23245,N_23231);
and U23316 (N_23316,N_23093,N_23068);
nor U23317 (N_23317,N_23176,N_23186);
xnor U23318 (N_23318,N_23149,N_23177);
nor U23319 (N_23319,N_23187,N_23018);
and U23320 (N_23320,N_23246,N_23027);
nand U23321 (N_23321,N_23080,N_23070);
nand U23322 (N_23322,N_23088,N_23039);
nor U23323 (N_23323,N_23248,N_23049);
nor U23324 (N_23324,N_23057,N_23147);
and U23325 (N_23325,N_23072,N_23006);
xnor U23326 (N_23326,N_23184,N_23164);
xor U23327 (N_23327,N_23172,N_23112);
nand U23328 (N_23328,N_23175,N_23143);
nand U23329 (N_23329,N_23135,N_23133);
nand U23330 (N_23330,N_23108,N_23066);
xor U23331 (N_23331,N_23095,N_23048);
nand U23332 (N_23332,N_23226,N_23064);
nand U23333 (N_23333,N_23026,N_23134);
nand U23334 (N_23334,N_23145,N_23051);
nor U23335 (N_23335,N_23115,N_23209);
or U23336 (N_23336,N_23241,N_23028);
and U23337 (N_23337,N_23024,N_23188);
and U23338 (N_23338,N_23195,N_23056);
nor U23339 (N_23339,N_23170,N_23139);
nand U23340 (N_23340,N_23161,N_23213);
and U23341 (N_23341,N_23085,N_23182);
nor U23342 (N_23342,N_23215,N_23002);
nand U23343 (N_23343,N_23117,N_23074);
nand U23344 (N_23344,N_23201,N_23071);
xnor U23345 (N_23345,N_23073,N_23154);
or U23346 (N_23346,N_23240,N_23234);
nand U23347 (N_23347,N_23144,N_23052);
or U23348 (N_23348,N_23004,N_23167);
nor U23349 (N_23349,N_23214,N_23247);
nand U23350 (N_23350,N_23094,N_23207);
nand U23351 (N_23351,N_23076,N_23237);
nor U23352 (N_23352,N_23089,N_23118);
xor U23353 (N_23353,N_23116,N_23138);
or U23354 (N_23354,N_23030,N_23084);
xnor U23355 (N_23355,N_23105,N_23035);
and U23356 (N_23356,N_23136,N_23022);
xor U23357 (N_23357,N_23041,N_23007);
xnor U23358 (N_23358,N_23159,N_23011);
and U23359 (N_23359,N_23012,N_23104);
nor U23360 (N_23360,N_23065,N_23010);
and U23361 (N_23361,N_23014,N_23233);
nor U23362 (N_23362,N_23199,N_23181);
nor U23363 (N_23363,N_23062,N_23023);
xor U23364 (N_23364,N_23055,N_23183);
nand U23365 (N_23365,N_23225,N_23078);
and U23366 (N_23366,N_23179,N_23044);
nand U23367 (N_23367,N_23079,N_23123);
or U23368 (N_23368,N_23217,N_23113);
or U23369 (N_23369,N_23206,N_23224);
nand U23370 (N_23370,N_23040,N_23077);
and U23371 (N_23371,N_23019,N_23025);
nor U23372 (N_23372,N_23120,N_23130);
or U23373 (N_23373,N_23129,N_23191);
and U23374 (N_23374,N_23090,N_23208);
and U23375 (N_23375,N_23227,N_23005);
and U23376 (N_23376,N_23191,N_23145);
nor U23377 (N_23377,N_23105,N_23075);
nand U23378 (N_23378,N_23133,N_23110);
xor U23379 (N_23379,N_23036,N_23161);
xnor U23380 (N_23380,N_23177,N_23185);
nand U23381 (N_23381,N_23087,N_23092);
xnor U23382 (N_23382,N_23046,N_23090);
and U23383 (N_23383,N_23008,N_23241);
and U23384 (N_23384,N_23075,N_23074);
nand U23385 (N_23385,N_23027,N_23213);
xor U23386 (N_23386,N_23079,N_23032);
and U23387 (N_23387,N_23037,N_23000);
nand U23388 (N_23388,N_23071,N_23018);
nand U23389 (N_23389,N_23240,N_23029);
or U23390 (N_23390,N_23241,N_23150);
and U23391 (N_23391,N_23171,N_23120);
nor U23392 (N_23392,N_23147,N_23017);
nand U23393 (N_23393,N_23011,N_23132);
nor U23394 (N_23394,N_23166,N_23132);
or U23395 (N_23395,N_23182,N_23098);
and U23396 (N_23396,N_23004,N_23200);
xor U23397 (N_23397,N_23080,N_23048);
nand U23398 (N_23398,N_23065,N_23013);
nand U23399 (N_23399,N_23021,N_23245);
nor U23400 (N_23400,N_23057,N_23246);
nand U23401 (N_23401,N_23099,N_23013);
nand U23402 (N_23402,N_23128,N_23168);
or U23403 (N_23403,N_23174,N_23014);
nor U23404 (N_23404,N_23047,N_23130);
nand U23405 (N_23405,N_23016,N_23137);
xor U23406 (N_23406,N_23078,N_23029);
or U23407 (N_23407,N_23249,N_23066);
nor U23408 (N_23408,N_23157,N_23223);
nor U23409 (N_23409,N_23031,N_23064);
nand U23410 (N_23410,N_23199,N_23146);
xor U23411 (N_23411,N_23249,N_23146);
and U23412 (N_23412,N_23085,N_23100);
and U23413 (N_23413,N_23124,N_23092);
nand U23414 (N_23414,N_23131,N_23178);
xor U23415 (N_23415,N_23010,N_23067);
and U23416 (N_23416,N_23034,N_23065);
or U23417 (N_23417,N_23021,N_23213);
nand U23418 (N_23418,N_23182,N_23059);
xnor U23419 (N_23419,N_23032,N_23247);
and U23420 (N_23420,N_23215,N_23056);
and U23421 (N_23421,N_23233,N_23130);
and U23422 (N_23422,N_23088,N_23171);
nand U23423 (N_23423,N_23126,N_23207);
nand U23424 (N_23424,N_23228,N_23009);
nand U23425 (N_23425,N_23191,N_23131);
or U23426 (N_23426,N_23200,N_23088);
and U23427 (N_23427,N_23040,N_23218);
nand U23428 (N_23428,N_23168,N_23083);
or U23429 (N_23429,N_23117,N_23021);
nor U23430 (N_23430,N_23017,N_23237);
nor U23431 (N_23431,N_23205,N_23089);
xor U23432 (N_23432,N_23099,N_23136);
or U23433 (N_23433,N_23154,N_23018);
nor U23434 (N_23434,N_23076,N_23071);
or U23435 (N_23435,N_23146,N_23215);
nand U23436 (N_23436,N_23077,N_23062);
xor U23437 (N_23437,N_23077,N_23204);
and U23438 (N_23438,N_23182,N_23081);
nand U23439 (N_23439,N_23241,N_23228);
or U23440 (N_23440,N_23127,N_23143);
or U23441 (N_23441,N_23123,N_23103);
xnor U23442 (N_23442,N_23139,N_23012);
nor U23443 (N_23443,N_23068,N_23016);
and U23444 (N_23444,N_23096,N_23091);
or U23445 (N_23445,N_23093,N_23227);
and U23446 (N_23446,N_23187,N_23122);
nand U23447 (N_23447,N_23127,N_23087);
or U23448 (N_23448,N_23089,N_23082);
xnor U23449 (N_23449,N_23033,N_23144);
nor U23450 (N_23450,N_23083,N_23213);
and U23451 (N_23451,N_23000,N_23154);
nor U23452 (N_23452,N_23205,N_23196);
and U23453 (N_23453,N_23123,N_23142);
or U23454 (N_23454,N_23031,N_23209);
nor U23455 (N_23455,N_23084,N_23241);
nor U23456 (N_23456,N_23066,N_23084);
or U23457 (N_23457,N_23104,N_23135);
and U23458 (N_23458,N_23094,N_23235);
and U23459 (N_23459,N_23024,N_23108);
or U23460 (N_23460,N_23220,N_23033);
and U23461 (N_23461,N_23187,N_23234);
xor U23462 (N_23462,N_23150,N_23030);
nor U23463 (N_23463,N_23140,N_23232);
nand U23464 (N_23464,N_23021,N_23026);
nand U23465 (N_23465,N_23139,N_23245);
xnor U23466 (N_23466,N_23187,N_23189);
or U23467 (N_23467,N_23232,N_23048);
or U23468 (N_23468,N_23195,N_23113);
nor U23469 (N_23469,N_23231,N_23211);
nor U23470 (N_23470,N_23008,N_23081);
and U23471 (N_23471,N_23061,N_23026);
and U23472 (N_23472,N_23165,N_23138);
nor U23473 (N_23473,N_23144,N_23027);
nand U23474 (N_23474,N_23180,N_23013);
nand U23475 (N_23475,N_23141,N_23061);
and U23476 (N_23476,N_23156,N_23014);
nor U23477 (N_23477,N_23023,N_23159);
and U23478 (N_23478,N_23231,N_23015);
and U23479 (N_23479,N_23035,N_23162);
nand U23480 (N_23480,N_23055,N_23025);
xnor U23481 (N_23481,N_23224,N_23156);
xnor U23482 (N_23482,N_23015,N_23232);
or U23483 (N_23483,N_23205,N_23153);
and U23484 (N_23484,N_23146,N_23162);
and U23485 (N_23485,N_23090,N_23194);
or U23486 (N_23486,N_23150,N_23180);
and U23487 (N_23487,N_23007,N_23139);
or U23488 (N_23488,N_23163,N_23202);
and U23489 (N_23489,N_23160,N_23105);
and U23490 (N_23490,N_23246,N_23094);
or U23491 (N_23491,N_23124,N_23226);
and U23492 (N_23492,N_23071,N_23110);
and U23493 (N_23493,N_23219,N_23070);
nand U23494 (N_23494,N_23115,N_23128);
and U23495 (N_23495,N_23083,N_23230);
xnor U23496 (N_23496,N_23060,N_23213);
xnor U23497 (N_23497,N_23071,N_23221);
nor U23498 (N_23498,N_23207,N_23004);
xnor U23499 (N_23499,N_23073,N_23113);
and U23500 (N_23500,N_23331,N_23320);
xnor U23501 (N_23501,N_23336,N_23356);
nor U23502 (N_23502,N_23344,N_23406);
nor U23503 (N_23503,N_23474,N_23374);
xnor U23504 (N_23504,N_23273,N_23340);
nand U23505 (N_23505,N_23359,N_23268);
nor U23506 (N_23506,N_23452,N_23437);
and U23507 (N_23507,N_23477,N_23254);
and U23508 (N_23508,N_23305,N_23461);
nand U23509 (N_23509,N_23269,N_23416);
or U23510 (N_23510,N_23421,N_23289);
or U23511 (N_23511,N_23319,N_23330);
nor U23512 (N_23512,N_23353,N_23450);
xor U23513 (N_23513,N_23283,N_23458);
and U23514 (N_23514,N_23365,N_23424);
or U23515 (N_23515,N_23482,N_23386);
nor U23516 (N_23516,N_23311,N_23495);
xnor U23517 (N_23517,N_23298,N_23418);
nand U23518 (N_23518,N_23481,N_23489);
or U23519 (N_23519,N_23494,N_23264);
nor U23520 (N_23520,N_23380,N_23310);
xor U23521 (N_23521,N_23277,N_23355);
or U23522 (N_23522,N_23251,N_23397);
nand U23523 (N_23523,N_23366,N_23262);
nor U23524 (N_23524,N_23297,N_23413);
nand U23525 (N_23525,N_23449,N_23425);
nand U23526 (N_23526,N_23307,N_23472);
or U23527 (N_23527,N_23493,N_23480);
and U23528 (N_23528,N_23275,N_23479);
or U23529 (N_23529,N_23498,N_23491);
or U23530 (N_23530,N_23490,N_23326);
or U23531 (N_23531,N_23408,N_23306);
and U23532 (N_23532,N_23304,N_23260);
or U23533 (N_23533,N_23463,N_23272);
or U23534 (N_23534,N_23325,N_23476);
and U23535 (N_23535,N_23293,N_23339);
and U23536 (N_23536,N_23372,N_23379);
or U23537 (N_23537,N_23405,N_23337);
xor U23538 (N_23538,N_23459,N_23335);
nor U23539 (N_23539,N_23422,N_23362);
nor U23540 (N_23540,N_23485,N_23396);
nor U23541 (N_23541,N_23303,N_23391);
xnor U23542 (N_23542,N_23377,N_23456);
nand U23543 (N_23543,N_23350,N_23327);
xnor U23544 (N_23544,N_23341,N_23441);
or U23545 (N_23545,N_23387,N_23438);
or U23546 (N_23546,N_23381,N_23345);
or U23547 (N_23547,N_23445,N_23294);
or U23548 (N_23548,N_23488,N_23270);
and U23549 (N_23549,N_23499,N_23486);
xor U23550 (N_23550,N_23442,N_23349);
nor U23551 (N_23551,N_23258,N_23423);
nor U23552 (N_23552,N_23384,N_23357);
xnor U23553 (N_23553,N_23292,N_23440);
xor U23554 (N_23554,N_23465,N_23402);
nor U23555 (N_23555,N_23411,N_23360);
or U23556 (N_23556,N_23370,N_23271);
and U23557 (N_23557,N_23466,N_23316);
nand U23558 (N_23558,N_23315,N_23317);
and U23559 (N_23559,N_23288,N_23473);
and U23560 (N_23560,N_23388,N_23484);
or U23561 (N_23561,N_23407,N_23382);
or U23562 (N_23562,N_23256,N_23265);
nor U23563 (N_23563,N_23351,N_23492);
nor U23564 (N_23564,N_23389,N_23393);
xnor U23565 (N_23565,N_23276,N_23285);
or U23566 (N_23566,N_23253,N_23280);
or U23567 (N_23567,N_23301,N_23401);
xor U23568 (N_23568,N_23446,N_23410);
and U23569 (N_23569,N_23299,N_23329);
nand U23570 (N_23570,N_23312,N_23313);
nand U23571 (N_23571,N_23453,N_23274);
or U23572 (N_23572,N_23496,N_23309);
nand U23573 (N_23573,N_23390,N_23435);
and U23574 (N_23574,N_23318,N_23400);
nand U23575 (N_23575,N_23295,N_23469);
and U23576 (N_23576,N_23385,N_23475);
and U23577 (N_23577,N_23334,N_23281);
and U23578 (N_23578,N_23279,N_23375);
or U23579 (N_23579,N_23427,N_23428);
nand U23580 (N_23580,N_23347,N_23267);
and U23581 (N_23581,N_23324,N_23308);
nand U23582 (N_23582,N_23403,N_23348);
nor U23583 (N_23583,N_23426,N_23364);
nor U23584 (N_23584,N_23328,N_23420);
or U23585 (N_23585,N_23278,N_23286);
or U23586 (N_23586,N_23436,N_23468);
xor U23587 (N_23587,N_23399,N_23368);
nor U23588 (N_23588,N_23352,N_23419);
and U23589 (N_23589,N_23394,N_23415);
nor U23590 (N_23590,N_23263,N_23284);
xnor U23591 (N_23591,N_23338,N_23363);
nand U23592 (N_23592,N_23409,N_23395);
nor U23593 (N_23593,N_23323,N_23432);
nor U23594 (N_23594,N_23462,N_23257);
nor U23595 (N_23595,N_23342,N_23346);
xor U23596 (N_23596,N_23457,N_23255);
and U23597 (N_23597,N_23439,N_23464);
xor U23598 (N_23598,N_23414,N_23371);
nor U23599 (N_23599,N_23314,N_23404);
or U23600 (N_23600,N_23332,N_23290);
nand U23601 (N_23601,N_23296,N_23467);
or U23602 (N_23602,N_23321,N_23448);
nor U23603 (N_23603,N_23343,N_23398);
or U23604 (N_23604,N_23483,N_23333);
nand U23605 (N_23605,N_23478,N_23376);
or U23606 (N_23606,N_23447,N_23392);
xor U23607 (N_23607,N_23361,N_23300);
nand U23608 (N_23608,N_23431,N_23367);
or U23609 (N_23609,N_23434,N_23358);
nor U23610 (N_23610,N_23291,N_23250);
xnor U23611 (N_23611,N_23383,N_23454);
and U23612 (N_23612,N_23433,N_23417);
and U23613 (N_23613,N_23497,N_23369);
or U23614 (N_23614,N_23287,N_23259);
nand U23615 (N_23615,N_23443,N_23470);
and U23616 (N_23616,N_23471,N_23302);
and U23617 (N_23617,N_23261,N_23429);
xnor U23618 (N_23618,N_23487,N_23455);
xor U23619 (N_23619,N_23322,N_23460);
and U23620 (N_23620,N_23266,N_23354);
nand U23621 (N_23621,N_23282,N_23430);
nor U23622 (N_23622,N_23412,N_23373);
or U23623 (N_23623,N_23252,N_23378);
and U23624 (N_23624,N_23444,N_23451);
xor U23625 (N_23625,N_23304,N_23341);
and U23626 (N_23626,N_23320,N_23434);
nand U23627 (N_23627,N_23286,N_23470);
nor U23628 (N_23628,N_23262,N_23363);
nand U23629 (N_23629,N_23409,N_23255);
or U23630 (N_23630,N_23251,N_23378);
nor U23631 (N_23631,N_23356,N_23471);
xnor U23632 (N_23632,N_23384,N_23343);
and U23633 (N_23633,N_23435,N_23322);
xnor U23634 (N_23634,N_23409,N_23420);
or U23635 (N_23635,N_23469,N_23354);
xor U23636 (N_23636,N_23395,N_23332);
or U23637 (N_23637,N_23467,N_23411);
nand U23638 (N_23638,N_23309,N_23337);
xnor U23639 (N_23639,N_23329,N_23408);
or U23640 (N_23640,N_23395,N_23315);
and U23641 (N_23641,N_23466,N_23364);
or U23642 (N_23642,N_23254,N_23298);
nor U23643 (N_23643,N_23318,N_23315);
and U23644 (N_23644,N_23320,N_23382);
or U23645 (N_23645,N_23266,N_23292);
xnor U23646 (N_23646,N_23309,N_23498);
nand U23647 (N_23647,N_23270,N_23434);
xor U23648 (N_23648,N_23346,N_23309);
or U23649 (N_23649,N_23453,N_23258);
xnor U23650 (N_23650,N_23472,N_23381);
nor U23651 (N_23651,N_23267,N_23365);
and U23652 (N_23652,N_23487,N_23472);
and U23653 (N_23653,N_23260,N_23412);
or U23654 (N_23654,N_23334,N_23417);
or U23655 (N_23655,N_23297,N_23395);
or U23656 (N_23656,N_23404,N_23408);
xnor U23657 (N_23657,N_23424,N_23280);
or U23658 (N_23658,N_23487,N_23481);
xor U23659 (N_23659,N_23394,N_23424);
or U23660 (N_23660,N_23474,N_23354);
nor U23661 (N_23661,N_23250,N_23382);
or U23662 (N_23662,N_23464,N_23390);
or U23663 (N_23663,N_23311,N_23484);
xnor U23664 (N_23664,N_23482,N_23297);
nor U23665 (N_23665,N_23303,N_23280);
nand U23666 (N_23666,N_23325,N_23271);
nor U23667 (N_23667,N_23380,N_23379);
and U23668 (N_23668,N_23446,N_23434);
xnor U23669 (N_23669,N_23413,N_23437);
or U23670 (N_23670,N_23433,N_23338);
nand U23671 (N_23671,N_23318,N_23270);
nand U23672 (N_23672,N_23274,N_23363);
xor U23673 (N_23673,N_23285,N_23357);
nand U23674 (N_23674,N_23424,N_23475);
or U23675 (N_23675,N_23285,N_23272);
nand U23676 (N_23676,N_23257,N_23492);
xnor U23677 (N_23677,N_23323,N_23266);
and U23678 (N_23678,N_23389,N_23307);
xor U23679 (N_23679,N_23392,N_23270);
xor U23680 (N_23680,N_23322,N_23395);
nand U23681 (N_23681,N_23496,N_23373);
nand U23682 (N_23682,N_23480,N_23341);
nand U23683 (N_23683,N_23334,N_23344);
or U23684 (N_23684,N_23447,N_23266);
nor U23685 (N_23685,N_23467,N_23314);
nand U23686 (N_23686,N_23429,N_23394);
or U23687 (N_23687,N_23417,N_23465);
nand U23688 (N_23688,N_23475,N_23408);
and U23689 (N_23689,N_23334,N_23450);
nor U23690 (N_23690,N_23323,N_23305);
nor U23691 (N_23691,N_23362,N_23396);
nand U23692 (N_23692,N_23462,N_23253);
xnor U23693 (N_23693,N_23299,N_23370);
xor U23694 (N_23694,N_23369,N_23479);
xnor U23695 (N_23695,N_23391,N_23266);
or U23696 (N_23696,N_23373,N_23431);
xor U23697 (N_23697,N_23440,N_23379);
xor U23698 (N_23698,N_23364,N_23275);
or U23699 (N_23699,N_23331,N_23352);
or U23700 (N_23700,N_23290,N_23437);
nor U23701 (N_23701,N_23440,N_23356);
nand U23702 (N_23702,N_23455,N_23380);
nor U23703 (N_23703,N_23489,N_23279);
nand U23704 (N_23704,N_23314,N_23349);
and U23705 (N_23705,N_23413,N_23468);
nor U23706 (N_23706,N_23477,N_23301);
and U23707 (N_23707,N_23276,N_23415);
or U23708 (N_23708,N_23330,N_23283);
xor U23709 (N_23709,N_23480,N_23360);
or U23710 (N_23710,N_23304,N_23371);
nand U23711 (N_23711,N_23375,N_23271);
xnor U23712 (N_23712,N_23478,N_23339);
or U23713 (N_23713,N_23339,N_23457);
nor U23714 (N_23714,N_23390,N_23378);
xor U23715 (N_23715,N_23435,N_23463);
nor U23716 (N_23716,N_23411,N_23319);
xor U23717 (N_23717,N_23377,N_23457);
xnor U23718 (N_23718,N_23324,N_23441);
xnor U23719 (N_23719,N_23442,N_23319);
xor U23720 (N_23720,N_23298,N_23366);
and U23721 (N_23721,N_23378,N_23288);
and U23722 (N_23722,N_23373,N_23265);
or U23723 (N_23723,N_23261,N_23250);
xor U23724 (N_23724,N_23276,N_23457);
nor U23725 (N_23725,N_23445,N_23446);
nand U23726 (N_23726,N_23344,N_23304);
nor U23727 (N_23727,N_23409,N_23371);
xor U23728 (N_23728,N_23340,N_23291);
xnor U23729 (N_23729,N_23369,N_23404);
or U23730 (N_23730,N_23354,N_23320);
xnor U23731 (N_23731,N_23457,N_23383);
nand U23732 (N_23732,N_23264,N_23258);
or U23733 (N_23733,N_23456,N_23281);
xnor U23734 (N_23734,N_23311,N_23355);
nor U23735 (N_23735,N_23350,N_23378);
nor U23736 (N_23736,N_23304,N_23305);
or U23737 (N_23737,N_23450,N_23472);
nand U23738 (N_23738,N_23400,N_23438);
or U23739 (N_23739,N_23435,N_23471);
nor U23740 (N_23740,N_23368,N_23392);
xor U23741 (N_23741,N_23451,N_23377);
nand U23742 (N_23742,N_23377,N_23321);
and U23743 (N_23743,N_23477,N_23307);
nor U23744 (N_23744,N_23254,N_23323);
nor U23745 (N_23745,N_23481,N_23429);
nand U23746 (N_23746,N_23388,N_23275);
xnor U23747 (N_23747,N_23328,N_23251);
nor U23748 (N_23748,N_23386,N_23287);
nor U23749 (N_23749,N_23308,N_23382);
xnor U23750 (N_23750,N_23651,N_23735);
nor U23751 (N_23751,N_23567,N_23596);
nor U23752 (N_23752,N_23727,N_23539);
or U23753 (N_23753,N_23610,N_23646);
nand U23754 (N_23754,N_23599,N_23699);
or U23755 (N_23755,N_23739,N_23736);
and U23756 (N_23756,N_23561,N_23548);
nand U23757 (N_23757,N_23513,N_23505);
nor U23758 (N_23758,N_23632,N_23652);
xor U23759 (N_23759,N_23509,N_23745);
nor U23760 (N_23760,N_23722,N_23524);
nand U23761 (N_23761,N_23617,N_23729);
nor U23762 (N_23762,N_23525,N_23695);
xnor U23763 (N_23763,N_23517,N_23710);
xnor U23764 (N_23764,N_23607,N_23728);
and U23765 (N_23765,N_23580,N_23589);
nand U23766 (N_23766,N_23511,N_23721);
nor U23767 (N_23767,N_23566,N_23590);
nand U23768 (N_23768,N_23604,N_23606);
or U23769 (N_23769,N_23692,N_23522);
xnor U23770 (N_23770,N_23689,N_23623);
or U23771 (N_23771,N_23701,N_23719);
and U23772 (N_23772,N_23747,N_23593);
nor U23773 (N_23773,N_23663,N_23504);
or U23774 (N_23774,N_23621,N_23559);
nand U23775 (N_23775,N_23510,N_23746);
xnor U23776 (N_23776,N_23564,N_23698);
and U23777 (N_23777,N_23731,N_23565);
and U23778 (N_23778,N_23515,N_23712);
and U23779 (N_23779,N_23612,N_23666);
or U23780 (N_23780,N_23740,N_23609);
nand U23781 (N_23781,N_23625,N_23681);
and U23782 (N_23782,N_23616,N_23532);
or U23783 (N_23783,N_23624,N_23603);
xor U23784 (N_23784,N_23702,N_23647);
nand U23785 (N_23785,N_23634,N_23562);
xor U23786 (N_23786,N_23748,N_23709);
nand U23787 (N_23787,N_23725,N_23633);
or U23788 (N_23788,N_23742,N_23551);
nand U23789 (N_23789,N_23585,N_23635);
or U23790 (N_23790,N_23568,N_23584);
and U23791 (N_23791,N_23619,N_23643);
and U23792 (N_23792,N_23527,N_23713);
nor U23793 (N_23793,N_23654,N_23605);
nand U23794 (N_23794,N_23672,N_23690);
nand U23795 (N_23795,N_23639,N_23648);
or U23796 (N_23796,N_23547,N_23531);
and U23797 (N_23797,N_23519,N_23573);
and U23798 (N_23798,N_23611,N_23744);
xnor U23799 (N_23799,N_23536,N_23688);
and U23800 (N_23800,N_23583,N_23705);
nand U23801 (N_23801,N_23658,N_23732);
xor U23802 (N_23802,N_23544,N_23655);
xnor U23803 (N_23803,N_23708,N_23668);
or U23804 (N_23804,N_23540,N_23577);
and U23805 (N_23805,N_23726,N_23597);
nor U23806 (N_23806,N_23613,N_23506);
nand U23807 (N_23807,N_23626,N_23718);
nand U23808 (N_23808,N_23685,N_23642);
and U23809 (N_23809,N_23512,N_23669);
and U23810 (N_23810,N_23529,N_23707);
nor U23811 (N_23811,N_23697,N_23600);
xor U23812 (N_23812,N_23700,N_23683);
or U23813 (N_23813,N_23538,N_23737);
and U23814 (N_23814,N_23576,N_23704);
xor U23815 (N_23815,N_23514,N_23582);
or U23816 (N_23816,N_23686,N_23557);
and U23817 (N_23817,N_23591,N_23546);
nand U23818 (N_23818,N_23570,N_23595);
xor U23819 (N_23819,N_23684,N_23574);
and U23820 (N_23820,N_23649,N_23743);
nand U23821 (N_23821,N_23520,N_23622);
nor U23822 (N_23822,N_23716,N_23549);
nand U23823 (N_23823,N_23656,N_23521);
or U23824 (N_23824,N_23734,N_23670);
xnor U23825 (N_23825,N_23659,N_23667);
xor U23826 (N_23826,N_23543,N_23749);
or U23827 (N_23827,N_23638,N_23674);
xor U23828 (N_23828,N_23637,N_23545);
and U23829 (N_23829,N_23594,N_23660);
nand U23830 (N_23830,N_23693,N_23662);
nor U23831 (N_23831,N_23644,N_23508);
nand U23832 (N_23832,N_23550,N_23738);
nand U23833 (N_23833,N_23502,N_23664);
nor U23834 (N_23834,N_23552,N_23587);
and U23835 (N_23835,N_23586,N_23620);
nor U23836 (N_23836,N_23665,N_23653);
or U23837 (N_23837,N_23571,N_23630);
or U23838 (N_23838,N_23541,N_23680);
and U23839 (N_23839,N_23723,N_23501);
nand U23840 (N_23840,N_23650,N_23602);
and U23841 (N_23841,N_23628,N_23694);
and U23842 (N_23842,N_23588,N_23636);
xnor U23843 (N_23843,N_23592,N_23657);
or U23844 (N_23844,N_23556,N_23614);
nand U23845 (N_23845,N_23572,N_23631);
or U23846 (N_23846,N_23715,N_23645);
nor U23847 (N_23847,N_23711,N_23730);
nor U23848 (N_23848,N_23661,N_23555);
nor U23849 (N_23849,N_23569,N_23554);
or U23850 (N_23850,N_23640,N_23598);
or U23851 (N_23851,N_23741,N_23578);
xnor U23852 (N_23852,N_23675,N_23618);
nand U23853 (N_23853,N_23601,N_23575);
nand U23854 (N_23854,N_23720,N_23523);
nor U23855 (N_23855,N_23608,N_23563);
and U23856 (N_23856,N_23500,N_23534);
nor U23857 (N_23857,N_23673,N_23703);
and U23858 (N_23858,N_23679,N_23676);
or U23859 (N_23859,N_23503,N_23537);
or U23860 (N_23860,N_23533,N_23687);
nor U23861 (N_23861,N_23717,N_23706);
nor U23862 (N_23862,N_23518,N_23691);
or U23863 (N_23863,N_23724,N_23535);
nor U23864 (N_23864,N_23581,N_23526);
or U23865 (N_23865,N_23553,N_23671);
nor U23866 (N_23866,N_23677,N_23558);
or U23867 (N_23867,N_23641,N_23627);
or U23868 (N_23868,N_23516,N_23733);
and U23869 (N_23869,N_23528,N_23560);
or U23870 (N_23870,N_23579,N_23714);
and U23871 (N_23871,N_23629,N_23615);
xnor U23872 (N_23872,N_23507,N_23530);
xnor U23873 (N_23873,N_23678,N_23696);
nor U23874 (N_23874,N_23682,N_23542);
nor U23875 (N_23875,N_23660,N_23656);
xor U23876 (N_23876,N_23533,N_23693);
or U23877 (N_23877,N_23617,N_23710);
nor U23878 (N_23878,N_23677,N_23587);
nand U23879 (N_23879,N_23656,N_23598);
or U23880 (N_23880,N_23709,N_23609);
nor U23881 (N_23881,N_23563,N_23642);
xor U23882 (N_23882,N_23597,N_23558);
or U23883 (N_23883,N_23510,N_23527);
nand U23884 (N_23884,N_23517,N_23569);
nor U23885 (N_23885,N_23678,N_23685);
xnor U23886 (N_23886,N_23665,N_23589);
nand U23887 (N_23887,N_23716,N_23537);
xor U23888 (N_23888,N_23654,N_23533);
nor U23889 (N_23889,N_23505,N_23559);
or U23890 (N_23890,N_23590,N_23689);
and U23891 (N_23891,N_23550,N_23636);
xnor U23892 (N_23892,N_23582,N_23648);
nand U23893 (N_23893,N_23676,N_23642);
or U23894 (N_23894,N_23680,N_23528);
nor U23895 (N_23895,N_23528,N_23583);
nor U23896 (N_23896,N_23562,N_23670);
nand U23897 (N_23897,N_23589,N_23730);
nand U23898 (N_23898,N_23640,N_23671);
xor U23899 (N_23899,N_23611,N_23686);
nand U23900 (N_23900,N_23527,N_23540);
xnor U23901 (N_23901,N_23733,N_23645);
nor U23902 (N_23902,N_23698,N_23514);
and U23903 (N_23903,N_23605,N_23594);
nor U23904 (N_23904,N_23601,N_23510);
nor U23905 (N_23905,N_23598,N_23524);
or U23906 (N_23906,N_23561,N_23664);
or U23907 (N_23907,N_23666,N_23585);
nand U23908 (N_23908,N_23575,N_23622);
and U23909 (N_23909,N_23639,N_23695);
xnor U23910 (N_23910,N_23592,N_23599);
nor U23911 (N_23911,N_23658,N_23601);
nor U23912 (N_23912,N_23700,N_23644);
or U23913 (N_23913,N_23617,N_23570);
nand U23914 (N_23914,N_23588,N_23715);
and U23915 (N_23915,N_23631,N_23567);
nand U23916 (N_23916,N_23514,N_23672);
nand U23917 (N_23917,N_23696,N_23650);
nand U23918 (N_23918,N_23530,N_23538);
or U23919 (N_23919,N_23571,N_23565);
or U23920 (N_23920,N_23564,N_23560);
nand U23921 (N_23921,N_23658,N_23541);
nand U23922 (N_23922,N_23729,N_23719);
and U23923 (N_23923,N_23555,N_23715);
xor U23924 (N_23924,N_23543,N_23558);
nor U23925 (N_23925,N_23663,N_23627);
and U23926 (N_23926,N_23615,N_23527);
and U23927 (N_23927,N_23727,N_23551);
nor U23928 (N_23928,N_23658,N_23621);
nor U23929 (N_23929,N_23671,N_23614);
or U23930 (N_23930,N_23711,N_23557);
or U23931 (N_23931,N_23591,N_23652);
nor U23932 (N_23932,N_23747,N_23719);
or U23933 (N_23933,N_23636,N_23568);
nor U23934 (N_23934,N_23660,N_23735);
or U23935 (N_23935,N_23588,N_23556);
and U23936 (N_23936,N_23713,N_23570);
and U23937 (N_23937,N_23641,N_23726);
or U23938 (N_23938,N_23739,N_23643);
nor U23939 (N_23939,N_23563,N_23526);
nand U23940 (N_23940,N_23535,N_23603);
nor U23941 (N_23941,N_23591,N_23651);
and U23942 (N_23942,N_23525,N_23521);
and U23943 (N_23943,N_23547,N_23636);
nor U23944 (N_23944,N_23564,N_23690);
nor U23945 (N_23945,N_23708,N_23625);
xor U23946 (N_23946,N_23721,N_23547);
xor U23947 (N_23947,N_23614,N_23586);
nand U23948 (N_23948,N_23575,N_23534);
xnor U23949 (N_23949,N_23541,N_23684);
and U23950 (N_23950,N_23578,N_23637);
nor U23951 (N_23951,N_23618,N_23582);
and U23952 (N_23952,N_23631,N_23734);
nand U23953 (N_23953,N_23603,N_23630);
or U23954 (N_23954,N_23732,N_23598);
nand U23955 (N_23955,N_23538,N_23616);
or U23956 (N_23956,N_23663,N_23511);
and U23957 (N_23957,N_23521,N_23698);
nor U23958 (N_23958,N_23734,N_23714);
or U23959 (N_23959,N_23728,N_23689);
nand U23960 (N_23960,N_23595,N_23715);
nand U23961 (N_23961,N_23677,N_23708);
or U23962 (N_23962,N_23509,N_23656);
or U23963 (N_23963,N_23737,N_23588);
and U23964 (N_23964,N_23601,N_23635);
nor U23965 (N_23965,N_23533,N_23529);
or U23966 (N_23966,N_23648,N_23745);
xnor U23967 (N_23967,N_23561,N_23724);
and U23968 (N_23968,N_23547,N_23652);
or U23969 (N_23969,N_23744,N_23521);
or U23970 (N_23970,N_23574,N_23507);
xnor U23971 (N_23971,N_23741,N_23676);
nand U23972 (N_23972,N_23547,N_23736);
nor U23973 (N_23973,N_23601,N_23649);
and U23974 (N_23974,N_23562,N_23736);
or U23975 (N_23975,N_23563,N_23596);
nor U23976 (N_23976,N_23685,N_23552);
nor U23977 (N_23977,N_23573,N_23657);
xnor U23978 (N_23978,N_23506,N_23571);
xor U23979 (N_23979,N_23645,N_23545);
nor U23980 (N_23980,N_23713,N_23653);
and U23981 (N_23981,N_23534,N_23548);
nor U23982 (N_23982,N_23691,N_23519);
nor U23983 (N_23983,N_23504,N_23622);
nor U23984 (N_23984,N_23517,N_23674);
xnor U23985 (N_23985,N_23610,N_23693);
and U23986 (N_23986,N_23564,N_23599);
xnor U23987 (N_23987,N_23683,N_23531);
and U23988 (N_23988,N_23634,N_23681);
or U23989 (N_23989,N_23630,N_23559);
and U23990 (N_23990,N_23625,N_23716);
nand U23991 (N_23991,N_23592,N_23594);
xnor U23992 (N_23992,N_23740,N_23723);
and U23993 (N_23993,N_23731,N_23745);
and U23994 (N_23994,N_23692,N_23645);
or U23995 (N_23995,N_23657,N_23717);
and U23996 (N_23996,N_23518,N_23685);
and U23997 (N_23997,N_23534,N_23579);
nor U23998 (N_23998,N_23694,N_23592);
and U23999 (N_23999,N_23656,N_23588);
xor U24000 (N_24000,N_23799,N_23816);
nand U24001 (N_24001,N_23948,N_23950);
or U24002 (N_24002,N_23851,N_23904);
and U24003 (N_24003,N_23831,N_23787);
nor U24004 (N_24004,N_23918,N_23891);
and U24005 (N_24005,N_23941,N_23863);
and U24006 (N_24006,N_23761,N_23887);
nand U24007 (N_24007,N_23923,N_23846);
nand U24008 (N_24008,N_23955,N_23835);
and U24009 (N_24009,N_23814,N_23876);
nand U24010 (N_24010,N_23951,N_23884);
nand U24011 (N_24011,N_23866,N_23803);
xnor U24012 (N_24012,N_23764,N_23898);
nor U24013 (N_24013,N_23800,N_23882);
nor U24014 (N_24014,N_23822,N_23850);
xor U24015 (N_24015,N_23897,N_23855);
xor U24016 (N_24016,N_23989,N_23962);
nor U24017 (N_24017,N_23862,N_23965);
or U24018 (N_24018,N_23973,N_23790);
xnor U24019 (N_24019,N_23817,N_23769);
and U24020 (N_24020,N_23754,N_23883);
xnor U24021 (N_24021,N_23886,N_23881);
nand U24022 (N_24022,N_23992,N_23774);
and U24023 (N_24023,N_23802,N_23902);
and U24024 (N_24024,N_23762,N_23957);
or U24025 (N_24025,N_23808,N_23793);
nand U24026 (N_24026,N_23848,N_23836);
or U24027 (N_24027,N_23860,N_23924);
and U24028 (N_24028,N_23879,N_23824);
nor U24029 (N_24029,N_23781,N_23840);
xnor U24030 (N_24030,N_23777,N_23776);
xnor U24031 (N_24031,N_23966,N_23907);
xnor U24032 (N_24032,N_23757,N_23798);
xor U24033 (N_24033,N_23819,N_23751);
nor U24034 (N_24034,N_23784,N_23901);
nand U24035 (N_24035,N_23928,N_23826);
nand U24036 (N_24036,N_23919,N_23772);
xor U24037 (N_24037,N_23892,N_23982);
and U24038 (N_24038,N_23801,N_23981);
nand U24039 (N_24039,N_23807,N_23818);
xnor U24040 (N_24040,N_23976,N_23968);
and U24041 (N_24041,N_23760,N_23984);
and U24042 (N_24042,N_23841,N_23830);
nor U24043 (N_24043,N_23942,N_23820);
or U24044 (N_24044,N_23980,N_23806);
and U24045 (N_24045,N_23970,N_23933);
or U24046 (N_24046,N_23839,N_23837);
nand U24047 (N_24047,N_23921,N_23988);
xor U24048 (N_24048,N_23779,N_23927);
nand U24049 (N_24049,N_23880,N_23997);
nor U24050 (N_24050,N_23783,N_23995);
and U24051 (N_24051,N_23999,N_23952);
and U24052 (N_24052,N_23930,N_23805);
nor U24053 (N_24053,N_23785,N_23847);
xor U24054 (N_24054,N_23874,N_23797);
or U24055 (N_24055,N_23912,N_23963);
or U24056 (N_24056,N_23811,N_23867);
nand U24057 (N_24057,N_23983,N_23878);
xnor U24058 (N_24058,N_23870,N_23810);
xnor U24059 (N_24059,N_23939,N_23972);
nand U24060 (N_24060,N_23809,N_23961);
and U24061 (N_24061,N_23926,N_23825);
and U24062 (N_24062,N_23975,N_23922);
nor U24063 (N_24063,N_23789,N_23991);
or U24064 (N_24064,N_23813,N_23844);
and U24065 (N_24065,N_23873,N_23823);
or U24066 (N_24066,N_23895,N_23900);
or U24067 (N_24067,N_23959,N_23905);
and U24068 (N_24068,N_23944,N_23770);
and U24069 (N_24069,N_23849,N_23979);
nand U24070 (N_24070,N_23821,N_23894);
nand U24071 (N_24071,N_23788,N_23868);
nand U24072 (N_24072,N_23947,N_23750);
and U24073 (N_24073,N_23977,N_23865);
or U24074 (N_24074,N_23827,N_23791);
nand U24075 (N_24075,N_23937,N_23759);
nor U24076 (N_24076,N_23829,N_23974);
nor U24077 (N_24077,N_23856,N_23843);
and U24078 (N_24078,N_23889,N_23877);
or U24079 (N_24079,N_23990,N_23815);
and U24080 (N_24080,N_23916,N_23853);
xnor U24081 (N_24081,N_23940,N_23896);
xor U24082 (N_24082,N_23778,N_23775);
or U24083 (N_24083,N_23861,N_23932);
and U24084 (N_24084,N_23872,N_23890);
or U24085 (N_24085,N_23864,N_23804);
or U24086 (N_24086,N_23795,N_23756);
nor U24087 (N_24087,N_23986,N_23766);
or U24088 (N_24088,N_23845,N_23796);
nand U24089 (N_24089,N_23969,N_23929);
xor U24090 (N_24090,N_23925,N_23838);
xnor U24091 (N_24091,N_23953,N_23909);
and U24092 (N_24092,N_23958,N_23967);
xor U24093 (N_24093,N_23931,N_23934);
xor U24094 (N_24094,N_23935,N_23913);
nand U24095 (N_24095,N_23875,N_23888);
nor U24096 (N_24096,N_23782,N_23833);
nor U24097 (N_24097,N_23920,N_23964);
and U24098 (N_24098,N_23752,N_23885);
and U24099 (N_24099,N_23985,N_23945);
nor U24100 (N_24100,N_23938,N_23910);
and U24101 (N_24101,N_23768,N_23763);
nand U24102 (N_24102,N_23812,N_23871);
xor U24103 (N_24103,N_23903,N_23780);
xnor U24104 (N_24104,N_23773,N_23946);
or U24105 (N_24105,N_23978,N_23993);
xnor U24106 (N_24106,N_23869,N_23834);
or U24107 (N_24107,N_23915,N_23771);
nand U24108 (N_24108,N_23971,N_23954);
nor U24109 (N_24109,N_23794,N_23832);
nor U24110 (N_24110,N_23828,N_23852);
nand U24111 (N_24111,N_23854,N_23998);
and U24112 (N_24112,N_23960,N_23893);
or U24113 (N_24113,N_23996,N_23943);
nand U24114 (N_24114,N_23755,N_23767);
and U24115 (N_24115,N_23899,N_23956);
or U24116 (N_24116,N_23917,N_23994);
xor U24117 (N_24117,N_23949,N_23765);
nor U24118 (N_24118,N_23758,N_23842);
or U24119 (N_24119,N_23936,N_23859);
nand U24120 (N_24120,N_23857,N_23914);
nand U24121 (N_24121,N_23987,N_23786);
xnor U24122 (N_24122,N_23792,N_23753);
xnor U24123 (N_24123,N_23858,N_23908);
or U24124 (N_24124,N_23911,N_23906);
or U24125 (N_24125,N_23848,N_23969);
nor U24126 (N_24126,N_23945,N_23942);
nand U24127 (N_24127,N_23880,N_23996);
and U24128 (N_24128,N_23773,N_23754);
or U24129 (N_24129,N_23782,N_23915);
nand U24130 (N_24130,N_23992,N_23840);
xor U24131 (N_24131,N_23883,N_23899);
and U24132 (N_24132,N_23778,N_23883);
xnor U24133 (N_24133,N_23995,N_23982);
nand U24134 (N_24134,N_23776,N_23751);
xor U24135 (N_24135,N_23842,N_23961);
xor U24136 (N_24136,N_23930,N_23809);
xnor U24137 (N_24137,N_23988,N_23812);
nor U24138 (N_24138,N_23944,N_23810);
and U24139 (N_24139,N_23976,N_23889);
and U24140 (N_24140,N_23754,N_23963);
xnor U24141 (N_24141,N_23793,N_23973);
nor U24142 (N_24142,N_23982,N_23948);
and U24143 (N_24143,N_23804,N_23843);
or U24144 (N_24144,N_23774,N_23873);
nor U24145 (N_24145,N_23753,N_23750);
and U24146 (N_24146,N_23980,N_23921);
nor U24147 (N_24147,N_23798,N_23812);
nor U24148 (N_24148,N_23883,N_23851);
nand U24149 (N_24149,N_23836,N_23771);
or U24150 (N_24150,N_23823,N_23896);
nand U24151 (N_24151,N_23788,N_23925);
and U24152 (N_24152,N_23939,N_23997);
or U24153 (N_24153,N_23931,N_23945);
nor U24154 (N_24154,N_23760,N_23944);
nand U24155 (N_24155,N_23994,N_23890);
and U24156 (N_24156,N_23914,N_23795);
and U24157 (N_24157,N_23921,N_23795);
nand U24158 (N_24158,N_23810,N_23851);
and U24159 (N_24159,N_23842,N_23913);
xor U24160 (N_24160,N_23864,N_23998);
xor U24161 (N_24161,N_23848,N_23799);
nand U24162 (N_24162,N_23881,N_23949);
or U24163 (N_24163,N_23769,N_23937);
and U24164 (N_24164,N_23944,N_23956);
nor U24165 (N_24165,N_23794,N_23863);
nor U24166 (N_24166,N_23951,N_23776);
nor U24167 (N_24167,N_23833,N_23838);
xnor U24168 (N_24168,N_23826,N_23803);
or U24169 (N_24169,N_23807,N_23997);
nand U24170 (N_24170,N_23915,N_23904);
nor U24171 (N_24171,N_23774,N_23976);
and U24172 (N_24172,N_23757,N_23874);
and U24173 (N_24173,N_23856,N_23784);
nand U24174 (N_24174,N_23830,N_23763);
xor U24175 (N_24175,N_23975,N_23977);
xnor U24176 (N_24176,N_23883,N_23784);
and U24177 (N_24177,N_23803,N_23953);
xnor U24178 (N_24178,N_23843,N_23761);
and U24179 (N_24179,N_23976,N_23923);
and U24180 (N_24180,N_23806,N_23760);
or U24181 (N_24181,N_23810,N_23949);
and U24182 (N_24182,N_23882,N_23904);
and U24183 (N_24183,N_23809,N_23831);
nand U24184 (N_24184,N_23786,N_23859);
or U24185 (N_24185,N_23825,N_23973);
and U24186 (N_24186,N_23796,N_23966);
nor U24187 (N_24187,N_23816,N_23997);
nand U24188 (N_24188,N_23830,N_23761);
nor U24189 (N_24189,N_23925,N_23877);
or U24190 (N_24190,N_23954,N_23824);
or U24191 (N_24191,N_23923,N_23866);
or U24192 (N_24192,N_23915,N_23842);
xnor U24193 (N_24193,N_23981,N_23888);
or U24194 (N_24194,N_23801,N_23879);
and U24195 (N_24195,N_23768,N_23815);
xor U24196 (N_24196,N_23819,N_23846);
or U24197 (N_24197,N_23905,N_23832);
and U24198 (N_24198,N_23776,N_23894);
and U24199 (N_24199,N_23878,N_23803);
nor U24200 (N_24200,N_23978,N_23768);
and U24201 (N_24201,N_23939,N_23859);
and U24202 (N_24202,N_23948,N_23932);
xnor U24203 (N_24203,N_23961,N_23797);
nand U24204 (N_24204,N_23924,N_23911);
xor U24205 (N_24205,N_23909,N_23935);
nor U24206 (N_24206,N_23965,N_23856);
or U24207 (N_24207,N_23812,N_23813);
nand U24208 (N_24208,N_23969,N_23838);
and U24209 (N_24209,N_23860,N_23903);
or U24210 (N_24210,N_23785,N_23805);
or U24211 (N_24211,N_23807,N_23861);
or U24212 (N_24212,N_23987,N_23824);
nand U24213 (N_24213,N_23983,N_23841);
nand U24214 (N_24214,N_23843,N_23763);
and U24215 (N_24215,N_23991,N_23905);
or U24216 (N_24216,N_23787,N_23789);
xor U24217 (N_24217,N_23887,N_23803);
nor U24218 (N_24218,N_23927,N_23816);
nand U24219 (N_24219,N_23951,N_23943);
nand U24220 (N_24220,N_23991,N_23876);
nand U24221 (N_24221,N_23798,N_23944);
and U24222 (N_24222,N_23874,N_23831);
xor U24223 (N_24223,N_23990,N_23859);
nand U24224 (N_24224,N_23958,N_23873);
nor U24225 (N_24225,N_23861,N_23912);
or U24226 (N_24226,N_23811,N_23841);
xnor U24227 (N_24227,N_23954,N_23858);
nand U24228 (N_24228,N_23840,N_23880);
nand U24229 (N_24229,N_23871,N_23972);
and U24230 (N_24230,N_23756,N_23897);
nand U24231 (N_24231,N_23867,N_23972);
and U24232 (N_24232,N_23828,N_23970);
xnor U24233 (N_24233,N_23904,N_23820);
or U24234 (N_24234,N_23830,N_23773);
nor U24235 (N_24235,N_23962,N_23776);
nor U24236 (N_24236,N_23793,N_23882);
nor U24237 (N_24237,N_23940,N_23976);
nor U24238 (N_24238,N_23903,N_23754);
nor U24239 (N_24239,N_23911,N_23810);
or U24240 (N_24240,N_23929,N_23960);
or U24241 (N_24241,N_23947,N_23924);
or U24242 (N_24242,N_23938,N_23998);
and U24243 (N_24243,N_23764,N_23975);
nand U24244 (N_24244,N_23893,N_23975);
xor U24245 (N_24245,N_23781,N_23816);
xor U24246 (N_24246,N_23773,N_23928);
xor U24247 (N_24247,N_23915,N_23861);
and U24248 (N_24248,N_23772,N_23964);
and U24249 (N_24249,N_23927,N_23908);
xor U24250 (N_24250,N_24033,N_24103);
xor U24251 (N_24251,N_24092,N_24229);
or U24252 (N_24252,N_24179,N_24111);
xor U24253 (N_24253,N_24086,N_24160);
nand U24254 (N_24254,N_24048,N_24023);
nor U24255 (N_24255,N_24000,N_24047);
xor U24256 (N_24256,N_24110,N_24227);
xor U24257 (N_24257,N_24097,N_24083);
nand U24258 (N_24258,N_24054,N_24236);
or U24259 (N_24259,N_24031,N_24007);
xnor U24260 (N_24260,N_24099,N_24162);
or U24261 (N_24261,N_24043,N_24008);
or U24262 (N_24262,N_24188,N_24025);
nor U24263 (N_24263,N_24061,N_24030);
xnor U24264 (N_24264,N_24168,N_24208);
nor U24265 (N_24265,N_24034,N_24101);
and U24266 (N_24266,N_24203,N_24002);
and U24267 (N_24267,N_24196,N_24209);
and U24268 (N_24268,N_24166,N_24181);
or U24269 (N_24269,N_24214,N_24073);
nor U24270 (N_24270,N_24234,N_24184);
nor U24271 (N_24271,N_24036,N_24138);
xor U24272 (N_24272,N_24186,N_24137);
nand U24273 (N_24273,N_24165,N_24076);
nand U24274 (N_24274,N_24192,N_24230);
nor U24275 (N_24275,N_24156,N_24027);
nand U24276 (N_24276,N_24022,N_24131);
nand U24277 (N_24277,N_24206,N_24112);
xor U24278 (N_24278,N_24080,N_24109);
xnor U24279 (N_24279,N_24012,N_24224);
nor U24280 (N_24280,N_24220,N_24155);
xor U24281 (N_24281,N_24056,N_24177);
nand U24282 (N_24282,N_24248,N_24020);
nor U24283 (N_24283,N_24035,N_24094);
xor U24284 (N_24284,N_24215,N_24151);
or U24285 (N_24285,N_24051,N_24144);
nor U24286 (N_24286,N_24201,N_24090);
xor U24287 (N_24287,N_24010,N_24057);
or U24288 (N_24288,N_24242,N_24091);
or U24289 (N_24289,N_24211,N_24154);
nor U24290 (N_24290,N_24197,N_24009);
xor U24291 (N_24291,N_24149,N_24053);
nor U24292 (N_24292,N_24233,N_24107);
or U24293 (N_24293,N_24223,N_24077);
and U24294 (N_24294,N_24130,N_24241);
xnor U24295 (N_24295,N_24021,N_24128);
xor U24296 (N_24296,N_24147,N_24070);
nand U24297 (N_24297,N_24139,N_24032);
nor U24298 (N_24298,N_24153,N_24205);
xnor U24299 (N_24299,N_24175,N_24152);
xnor U24300 (N_24300,N_24018,N_24195);
nor U24301 (N_24301,N_24182,N_24060);
nand U24302 (N_24302,N_24169,N_24222);
nand U24303 (N_24303,N_24052,N_24158);
and U24304 (N_24304,N_24011,N_24124);
nor U24305 (N_24305,N_24055,N_24029);
or U24306 (N_24306,N_24243,N_24202);
nor U24307 (N_24307,N_24078,N_24232);
nand U24308 (N_24308,N_24063,N_24019);
nor U24309 (N_24309,N_24016,N_24095);
nand U24310 (N_24310,N_24150,N_24219);
and U24311 (N_24311,N_24038,N_24167);
nor U24312 (N_24312,N_24134,N_24189);
xnor U24313 (N_24313,N_24075,N_24100);
or U24314 (N_24314,N_24132,N_24164);
nor U24315 (N_24315,N_24216,N_24163);
or U24316 (N_24316,N_24239,N_24096);
or U24317 (N_24317,N_24004,N_24085);
nor U24318 (N_24318,N_24194,N_24140);
and U24319 (N_24319,N_24116,N_24244);
and U24320 (N_24320,N_24120,N_24171);
and U24321 (N_24321,N_24013,N_24074);
and U24322 (N_24322,N_24087,N_24231);
nor U24323 (N_24323,N_24245,N_24088);
nor U24324 (N_24324,N_24104,N_24026);
and U24325 (N_24325,N_24106,N_24246);
nand U24326 (N_24326,N_24121,N_24058);
or U24327 (N_24327,N_24142,N_24143);
xnor U24328 (N_24328,N_24235,N_24024);
and U24329 (N_24329,N_24176,N_24204);
or U24330 (N_24330,N_24113,N_24098);
and U24331 (N_24331,N_24122,N_24199);
and U24332 (N_24332,N_24062,N_24228);
nand U24333 (N_24333,N_24066,N_24159);
xor U24334 (N_24334,N_24041,N_24081);
xnor U24335 (N_24335,N_24017,N_24133);
xor U24336 (N_24336,N_24183,N_24079);
xor U24337 (N_24337,N_24003,N_24240);
and U24338 (N_24338,N_24072,N_24059);
nor U24339 (N_24339,N_24117,N_24200);
xor U24340 (N_24340,N_24119,N_24141);
or U24341 (N_24341,N_24042,N_24102);
nor U24342 (N_24342,N_24118,N_24185);
or U24343 (N_24343,N_24028,N_24174);
nand U24344 (N_24344,N_24191,N_24136);
or U24345 (N_24345,N_24040,N_24145);
and U24346 (N_24346,N_24225,N_24084);
nor U24347 (N_24347,N_24198,N_24238);
nor U24348 (N_24348,N_24014,N_24005);
or U24349 (N_24349,N_24046,N_24127);
and U24350 (N_24350,N_24114,N_24157);
or U24351 (N_24351,N_24126,N_24190);
nand U24352 (N_24352,N_24125,N_24180);
nand U24353 (N_24353,N_24193,N_24069);
nand U24354 (N_24354,N_24050,N_24247);
xnor U24355 (N_24355,N_24001,N_24217);
nor U24356 (N_24356,N_24146,N_24161);
and U24357 (N_24357,N_24221,N_24006);
xnor U24358 (N_24358,N_24173,N_24170);
and U24359 (N_24359,N_24226,N_24049);
xnor U24360 (N_24360,N_24064,N_24207);
and U24361 (N_24361,N_24045,N_24212);
and U24362 (N_24362,N_24082,N_24108);
xor U24363 (N_24363,N_24237,N_24039);
nor U24364 (N_24364,N_24015,N_24129);
and U24365 (N_24365,N_24213,N_24210);
and U24366 (N_24366,N_24218,N_24178);
xor U24367 (N_24367,N_24089,N_24105);
xnor U24368 (N_24368,N_24065,N_24148);
or U24369 (N_24369,N_24068,N_24115);
and U24370 (N_24370,N_24249,N_24123);
xnor U24371 (N_24371,N_24172,N_24071);
and U24372 (N_24372,N_24135,N_24187);
and U24373 (N_24373,N_24037,N_24067);
nand U24374 (N_24374,N_24093,N_24044);
nand U24375 (N_24375,N_24232,N_24166);
or U24376 (N_24376,N_24195,N_24140);
and U24377 (N_24377,N_24178,N_24165);
nor U24378 (N_24378,N_24119,N_24224);
or U24379 (N_24379,N_24199,N_24197);
and U24380 (N_24380,N_24241,N_24146);
and U24381 (N_24381,N_24184,N_24121);
nor U24382 (N_24382,N_24220,N_24010);
and U24383 (N_24383,N_24148,N_24037);
xor U24384 (N_24384,N_24168,N_24191);
nand U24385 (N_24385,N_24164,N_24161);
xor U24386 (N_24386,N_24012,N_24163);
nand U24387 (N_24387,N_24046,N_24105);
nand U24388 (N_24388,N_24148,N_24249);
nor U24389 (N_24389,N_24230,N_24102);
or U24390 (N_24390,N_24166,N_24139);
or U24391 (N_24391,N_24032,N_24167);
nand U24392 (N_24392,N_24110,N_24029);
and U24393 (N_24393,N_24119,N_24083);
and U24394 (N_24394,N_24099,N_24240);
nand U24395 (N_24395,N_24034,N_24157);
nor U24396 (N_24396,N_24200,N_24087);
or U24397 (N_24397,N_24181,N_24012);
or U24398 (N_24398,N_24112,N_24028);
nor U24399 (N_24399,N_24108,N_24206);
nor U24400 (N_24400,N_24174,N_24229);
xor U24401 (N_24401,N_24147,N_24182);
or U24402 (N_24402,N_24168,N_24042);
nor U24403 (N_24403,N_24170,N_24161);
nand U24404 (N_24404,N_24171,N_24142);
xor U24405 (N_24405,N_24149,N_24066);
and U24406 (N_24406,N_24137,N_24149);
nand U24407 (N_24407,N_24034,N_24243);
nor U24408 (N_24408,N_24154,N_24226);
or U24409 (N_24409,N_24224,N_24120);
or U24410 (N_24410,N_24180,N_24162);
and U24411 (N_24411,N_24155,N_24234);
nand U24412 (N_24412,N_24169,N_24132);
and U24413 (N_24413,N_24072,N_24214);
and U24414 (N_24414,N_24215,N_24175);
xor U24415 (N_24415,N_24063,N_24172);
nand U24416 (N_24416,N_24193,N_24043);
nor U24417 (N_24417,N_24023,N_24137);
and U24418 (N_24418,N_24019,N_24159);
or U24419 (N_24419,N_24049,N_24191);
or U24420 (N_24420,N_24153,N_24160);
and U24421 (N_24421,N_24017,N_24156);
and U24422 (N_24422,N_24117,N_24100);
and U24423 (N_24423,N_24085,N_24236);
or U24424 (N_24424,N_24190,N_24079);
nand U24425 (N_24425,N_24194,N_24138);
or U24426 (N_24426,N_24084,N_24176);
nand U24427 (N_24427,N_24199,N_24176);
or U24428 (N_24428,N_24082,N_24160);
and U24429 (N_24429,N_24172,N_24110);
or U24430 (N_24430,N_24121,N_24079);
nand U24431 (N_24431,N_24054,N_24075);
nand U24432 (N_24432,N_24036,N_24006);
nor U24433 (N_24433,N_24043,N_24208);
nand U24434 (N_24434,N_24185,N_24187);
and U24435 (N_24435,N_24087,N_24068);
and U24436 (N_24436,N_24220,N_24097);
nor U24437 (N_24437,N_24099,N_24176);
xor U24438 (N_24438,N_24192,N_24117);
nor U24439 (N_24439,N_24149,N_24023);
nor U24440 (N_24440,N_24221,N_24241);
or U24441 (N_24441,N_24003,N_24148);
and U24442 (N_24442,N_24243,N_24121);
and U24443 (N_24443,N_24171,N_24209);
xnor U24444 (N_24444,N_24026,N_24168);
nor U24445 (N_24445,N_24131,N_24115);
nor U24446 (N_24446,N_24044,N_24123);
or U24447 (N_24447,N_24248,N_24039);
xor U24448 (N_24448,N_24105,N_24097);
or U24449 (N_24449,N_24068,N_24030);
xor U24450 (N_24450,N_24099,N_24059);
nand U24451 (N_24451,N_24088,N_24208);
nor U24452 (N_24452,N_24014,N_24163);
nor U24453 (N_24453,N_24245,N_24105);
nand U24454 (N_24454,N_24083,N_24020);
xor U24455 (N_24455,N_24249,N_24104);
xor U24456 (N_24456,N_24011,N_24049);
xnor U24457 (N_24457,N_24003,N_24020);
nand U24458 (N_24458,N_24186,N_24031);
nor U24459 (N_24459,N_24070,N_24066);
nor U24460 (N_24460,N_24099,N_24236);
xnor U24461 (N_24461,N_24182,N_24169);
or U24462 (N_24462,N_24003,N_24084);
or U24463 (N_24463,N_24038,N_24066);
or U24464 (N_24464,N_24249,N_24032);
xnor U24465 (N_24465,N_24123,N_24211);
nor U24466 (N_24466,N_24244,N_24194);
xnor U24467 (N_24467,N_24174,N_24113);
or U24468 (N_24468,N_24119,N_24007);
nand U24469 (N_24469,N_24058,N_24110);
nor U24470 (N_24470,N_24081,N_24188);
nand U24471 (N_24471,N_24147,N_24030);
xor U24472 (N_24472,N_24017,N_24055);
nor U24473 (N_24473,N_24014,N_24012);
xnor U24474 (N_24474,N_24087,N_24187);
nor U24475 (N_24475,N_24080,N_24083);
or U24476 (N_24476,N_24120,N_24032);
nand U24477 (N_24477,N_24222,N_24120);
nand U24478 (N_24478,N_24205,N_24130);
xor U24479 (N_24479,N_24062,N_24143);
nor U24480 (N_24480,N_24103,N_24012);
xnor U24481 (N_24481,N_24103,N_24069);
or U24482 (N_24482,N_24038,N_24021);
and U24483 (N_24483,N_24178,N_24029);
and U24484 (N_24484,N_24003,N_24144);
nand U24485 (N_24485,N_24074,N_24016);
or U24486 (N_24486,N_24241,N_24192);
nand U24487 (N_24487,N_24091,N_24238);
nand U24488 (N_24488,N_24052,N_24210);
or U24489 (N_24489,N_24097,N_24022);
xnor U24490 (N_24490,N_24194,N_24190);
or U24491 (N_24491,N_24072,N_24069);
nand U24492 (N_24492,N_24137,N_24037);
nor U24493 (N_24493,N_24165,N_24158);
nor U24494 (N_24494,N_24108,N_24023);
xor U24495 (N_24495,N_24238,N_24077);
nor U24496 (N_24496,N_24199,N_24126);
xnor U24497 (N_24497,N_24170,N_24171);
and U24498 (N_24498,N_24048,N_24100);
and U24499 (N_24499,N_24013,N_24219);
nor U24500 (N_24500,N_24350,N_24439);
xor U24501 (N_24501,N_24344,N_24267);
nand U24502 (N_24502,N_24391,N_24404);
xnor U24503 (N_24503,N_24322,N_24318);
nor U24504 (N_24504,N_24284,N_24354);
and U24505 (N_24505,N_24272,N_24296);
and U24506 (N_24506,N_24371,N_24312);
nor U24507 (N_24507,N_24308,N_24377);
and U24508 (N_24508,N_24451,N_24429);
xor U24509 (N_24509,N_24300,N_24442);
nand U24510 (N_24510,N_24266,N_24328);
nor U24511 (N_24511,N_24368,N_24337);
xor U24512 (N_24512,N_24409,N_24254);
or U24513 (N_24513,N_24260,N_24352);
or U24514 (N_24514,N_24420,N_24405);
nor U24515 (N_24515,N_24473,N_24317);
nand U24516 (N_24516,N_24287,N_24295);
nor U24517 (N_24517,N_24392,N_24250);
nand U24518 (N_24518,N_24423,N_24252);
nand U24519 (N_24519,N_24433,N_24443);
and U24520 (N_24520,N_24324,N_24330);
nor U24521 (N_24521,N_24299,N_24407);
nor U24522 (N_24522,N_24410,N_24497);
nand U24523 (N_24523,N_24341,N_24380);
nor U24524 (N_24524,N_24251,N_24343);
and U24525 (N_24525,N_24413,N_24327);
or U24526 (N_24526,N_24477,N_24454);
and U24527 (N_24527,N_24446,N_24427);
nand U24528 (N_24528,N_24336,N_24282);
nor U24529 (N_24529,N_24263,N_24363);
or U24530 (N_24530,N_24349,N_24383);
nor U24531 (N_24531,N_24412,N_24387);
xor U24532 (N_24532,N_24453,N_24286);
xnor U24533 (N_24533,N_24458,N_24310);
xor U24534 (N_24534,N_24365,N_24345);
nand U24535 (N_24535,N_24273,N_24469);
or U24536 (N_24536,N_24465,N_24449);
and U24537 (N_24537,N_24393,N_24428);
nand U24538 (N_24538,N_24306,N_24478);
or U24539 (N_24539,N_24403,N_24361);
or U24540 (N_24540,N_24262,N_24493);
nand U24541 (N_24541,N_24321,N_24373);
nand U24542 (N_24542,N_24460,N_24489);
nor U24543 (N_24543,N_24358,N_24390);
xor U24544 (N_24544,N_24397,N_24258);
and U24545 (N_24545,N_24305,N_24325);
nand U24546 (N_24546,N_24357,N_24372);
nand U24547 (N_24547,N_24293,N_24483);
nor U24548 (N_24548,N_24471,N_24419);
and U24549 (N_24549,N_24370,N_24356);
nor U24550 (N_24550,N_24342,N_24333);
nor U24551 (N_24551,N_24276,N_24470);
nor U24552 (N_24552,N_24329,N_24472);
or U24553 (N_24553,N_24402,N_24285);
and U24554 (N_24554,N_24292,N_24386);
and U24555 (N_24555,N_24406,N_24467);
and U24556 (N_24556,N_24389,N_24416);
and U24557 (N_24557,N_24398,N_24332);
nor U24558 (N_24558,N_24297,N_24435);
nor U24559 (N_24559,N_24265,N_24264);
and U24560 (N_24560,N_24338,N_24290);
or U24561 (N_24561,N_24486,N_24440);
and U24562 (N_24562,N_24279,N_24311);
nand U24563 (N_24563,N_24418,N_24445);
nor U24564 (N_24564,N_24253,N_24426);
or U24565 (N_24565,N_24364,N_24359);
nand U24566 (N_24566,N_24268,N_24375);
and U24567 (N_24567,N_24360,N_24280);
xnor U24568 (N_24568,N_24259,N_24309);
xor U24569 (N_24569,N_24314,N_24274);
nor U24570 (N_24570,N_24436,N_24459);
and U24571 (N_24571,N_24256,N_24424);
nor U24572 (N_24572,N_24487,N_24421);
and U24573 (N_24573,N_24396,N_24385);
nand U24574 (N_24574,N_24294,N_24450);
xnor U24575 (N_24575,N_24485,N_24347);
nor U24576 (N_24576,N_24408,N_24269);
xor U24577 (N_24577,N_24366,N_24425);
and U24578 (N_24578,N_24320,N_24382);
or U24579 (N_24579,N_24304,N_24261);
xor U24580 (N_24580,N_24395,N_24491);
or U24581 (N_24581,N_24275,N_24379);
nand U24582 (N_24582,N_24351,N_24283);
nand U24583 (N_24583,N_24496,N_24464);
nor U24584 (N_24584,N_24326,N_24334);
xnor U24585 (N_24585,N_24301,N_24388);
xor U24586 (N_24586,N_24400,N_24481);
or U24587 (N_24587,N_24457,N_24495);
nand U24588 (N_24588,N_24476,N_24498);
xnor U24589 (N_24589,N_24432,N_24461);
or U24590 (N_24590,N_24434,N_24281);
and U24591 (N_24591,N_24289,N_24288);
nand U24592 (N_24592,N_24339,N_24319);
and U24593 (N_24593,N_24415,N_24499);
nand U24594 (N_24594,N_24422,N_24455);
nor U24595 (N_24595,N_24494,N_24255);
nor U24596 (N_24596,N_24374,N_24348);
xnor U24597 (N_24597,N_24401,N_24444);
xor U24598 (N_24598,N_24384,N_24456);
xnor U24599 (N_24599,N_24484,N_24466);
or U24600 (N_24600,N_24479,N_24315);
nand U24601 (N_24601,N_24303,N_24331);
and U24602 (N_24602,N_24316,N_24302);
xor U24603 (N_24603,N_24482,N_24452);
nand U24604 (N_24604,N_24313,N_24490);
nor U24605 (N_24605,N_24462,N_24411);
and U24606 (N_24606,N_24277,N_24367);
nor U24607 (N_24607,N_24335,N_24447);
nor U24608 (N_24608,N_24441,N_24376);
or U24609 (N_24609,N_24278,N_24369);
and U24610 (N_24610,N_24355,N_24430);
xnor U24611 (N_24611,N_24270,N_24257);
xor U24612 (N_24612,N_24291,N_24381);
nand U24613 (N_24613,N_24431,N_24298);
and U24614 (N_24614,N_24417,N_24414);
nand U24615 (N_24615,N_24271,N_24488);
or U24616 (N_24616,N_24474,N_24353);
and U24617 (N_24617,N_24394,N_24480);
nand U24618 (N_24618,N_24448,N_24340);
or U24619 (N_24619,N_24438,N_24463);
and U24620 (N_24620,N_24323,N_24399);
nand U24621 (N_24621,N_24437,N_24468);
nor U24622 (N_24622,N_24307,N_24492);
nand U24623 (N_24623,N_24346,N_24362);
nor U24624 (N_24624,N_24475,N_24378);
nand U24625 (N_24625,N_24461,N_24305);
nor U24626 (N_24626,N_24486,N_24326);
or U24627 (N_24627,N_24250,N_24478);
nor U24628 (N_24628,N_24361,N_24322);
and U24629 (N_24629,N_24417,N_24259);
or U24630 (N_24630,N_24411,N_24334);
xor U24631 (N_24631,N_24440,N_24429);
and U24632 (N_24632,N_24419,N_24351);
nor U24633 (N_24633,N_24348,N_24294);
nor U24634 (N_24634,N_24359,N_24401);
nand U24635 (N_24635,N_24333,N_24345);
nor U24636 (N_24636,N_24391,N_24364);
nor U24637 (N_24637,N_24483,N_24472);
nor U24638 (N_24638,N_24421,N_24370);
or U24639 (N_24639,N_24400,N_24478);
or U24640 (N_24640,N_24437,N_24369);
or U24641 (N_24641,N_24374,N_24494);
and U24642 (N_24642,N_24298,N_24344);
xor U24643 (N_24643,N_24460,N_24480);
nor U24644 (N_24644,N_24279,N_24350);
and U24645 (N_24645,N_24353,N_24499);
or U24646 (N_24646,N_24389,N_24376);
xor U24647 (N_24647,N_24420,N_24391);
nand U24648 (N_24648,N_24399,N_24359);
nor U24649 (N_24649,N_24335,N_24425);
xnor U24650 (N_24650,N_24301,N_24286);
or U24651 (N_24651,N_24426,N_24482);
nand U24652 (N_24652,N_24384,N_24286);
xor U24653 (N_24653,N_24433,N_24482);
and U24654 (N_24654,N_24292,N_24332);
xor U24655 (N_24655,N_24473,N_24419);
or U24656 (N_24656,N_24457,N_24402);
or U24657 (N_24657,N_24363,N_24388);
xnor U24658 (N_24658,N_24272,N_24251);
and U24659 (N_24659,N_24338,N_24409);
nor U24660 (N_24660,N_24388,N_24321);
nor U24661 (N_24661,N_24318,N_24360);
nor U24662 (N_24662,N_24470,N_24428);
nor U24663 (N_24663,N_24301,N_24497);
and U24664 (N_24664,N_24315,N_24337);
nor U24665 (N_24665,N_24297,N_24394);
and U24666 (N_24666,N_24438,N_24418);
or U24667 (N_24667,N_24493,N_24404);
and U24668 (N_24668,N_24287,N_24469);
nor U24669 (N_24669,N_24251,N_24349);
xnor U24670 (N_24670,N_24349,N_24411);
and U24671 (N_24671,N_24410,N_24334);
xnor U24672 (N_24672,N_24473,N_24347);
xnor U24673 (N_24673,N_24426,N_24361);
nor U24674 (N_24674,N_24252,N_24329);
and U24675 (N_24675,N_24260,N_24317);
and U24676 (N_24676,N_24392,N_24309);
or U24677 (N_24677,N_24351,N_24403);
nor U24678 (N_24678,N_24404,N_24319);
and U24679 (N_24679,N_24339,N_24366);
nand U24680 (N_24680,N_24496,N_24399);
xnor U24681 (N_24681,N_24396,N_24461);
and U24682 (N_24682,N_24381,N_24464);
or U24683 (N_24683,N_24407,N_24314);
xor U24684 (N_24684,N_24319,N_24423);
nor U24685 (N_24685,N_24257,N_24250);
or U24686 (N_24686,N_24381,N_24307);
nor U24687 (N_24687,N_24345,N_24383);
nand U24688 (N_24688,N_24288,N_24264);
nor U24689 (N_24689,N_24406,N_24275);
or U24690 (N_24690,N_24442,N_24456);
and U24691 (N_24691,N_24279,N_24410);
nand U24692 (N_24692,N_24448,N_24470);
and U24693 (N_24693,N_24283,N_24306);
and U24694 (N_24694,N_24385,N_24402);
or U24695 (N_24695,N_24391,N_24338);
nand U24696 (N_24696,N_24291,N_24262);
nand U24697 (N_24697,N_24342,N_24282);
nor U24698 (N_24698,N_24408,N_24255);
and U24699 (N_24699,N_24407,N_24415);
nor U24700 (N_24700,N_24449,N_24347);
nand U24701 (N_24701,N_24267,N_24372);
nand U24702 (N_24702,N_24317,N_24422);
nand U24703 (N_24703,N_24381,N_24300);
and U24704 (N_24704,N_24379,N_24463);
or U24705 (N_24705,N_24447,N_24359);
xor U24706 (N_24706,N_24465,N_24460);
nor U24707 (N_24707,N_24335,N_24250);
nand U24708 (N_24708,N_24408,N_24297);
nand U24709 (N_24709,N_24398,N_24383);
nand U24710 (N_24710,N_24398,N_24483);
nor U24711 (N_24711,N_24433,N_24478);
or U24712 (N_24712,N_24362,N_24378);
or U24713 (N_24713,N_24379,N_24280);
nor U24714 (N_24714,N_24429,N_24329);
nor U24715 (N_24715,N_24357,N_24256);
nor U24716 (N_24716,N_24307,N_24278);
xor U24717 (N_24717,N_24483,N_24485);
and U24718 (N_24718,N_24417,N_24436);
nand U24719 (N_24719,N_24312,N_24485);
or U24720 (N_24720,N_24493,N_24335);
and U24721 (N_24721,N_24345,N_24493);
or U24722 (N_24722,N_24278,N_24277);
xnor U24723 (N_24723,N_24435,N_24326);
or U24724 (N_24724,N_24321,N_24252);
or U24725 (N_24725,N_24265,N_24429);
xnor U24726 (N_24726,N_24385,N_24287);
xor U24727 (N_24727,N_24391,N_24311);
nand U24728 (N_24728,N_24433,N_24489);
or U24729 (N_24729,N_24435,N_24323);
nand U24730 (N_24730,N_24461,N_24486);
nand U24731 (N_24731,N_24437,N_24262);
xnor U24732 (N_24732,N_24272,N_24335);
or U24733 (N_24733,N_24297,N_24363);
xor U24734 (N_24734,N_24382,N_24492);
or U24735 (N_24735,N_24355,N_24348);
nand U24736 (N_24736,N_24358,N_24355);
xor U24737 (N_24737,N_24480,N_24359);
xor U24738 (N_24738,N_24357,N_24304);
or U24739 (N_24739,N_24309,N_24251);
nor U24740 (N_24740,N_24410,N_24480);
and U24741 (N_24741,N_24465,N_24411);
xnor U24742 (N_24742,N_24311,N_24361);
nor U24743 (N_24743,N_24496,N_24290);
xnor U24744 (N_24744,N_24267,N_24453);
nor U24745 (N_24745,N_24278,N_24440);
nor U24746 (N_24746,N_24393,N_24463);
or U24747 (N_24747,N_24397,N_24473);
nor U24748 (N_24748,N_24320,N_24329);
nand U24749 (N_24749,N_24307,N_24298);
nor U24750 (N_24750,N_24654,N_24684);
or U24751 (N_24751,N_24500,N_24720);
nand U24752 (N_24752,N_24659,N_24623);
nor U24753 (N_24753,N_24522,N_24545);
or U24754 (N_24754,N_24749,N_24657);
nor U24755 (N_24755,N_24591,N_24520);
and U24756 (N_24756,N_24601,N_24706);
nor U24757 (N_24757,N_24559,N_24595);
or U24758 (N_24758,N_24702,N_24586);
xor U24759 (N_24759,N_24596,N_24671);
nand U24760 (N_24760,N_24611,N_24570);
or U24761 (N_24761,N_24742,N_24538);
nor U24762 (N_24762,N_24650,N_24698);
nand U24763 (N_24763,N_24567,N_24539);
nor U24764 (N_24764,N_24518,N_24614);
and U24765 (N_24765,N_24687,N_24676);
nor U24766 (N_24766,N_24708,N_24587);
nor U24767 (N_24767,N_24686,N_24564);
xnor U24768 (N_24768,N_24747,N_24583);
nor U24769 (N_24769,N_24628,N_24725);
nand U24770 (N_24770,N_24662,N_24675);
nand U24771 (N_24771,N_24631,N_24673);
or U24772 (N_24772,N_24722,N_24584);
nor U24773 (N_24773,N_24593,N_24515);
or U24774 (N_24774,N_24592,N_24639);
or U24775 (N_24775,N_24705,N_24534);
or U24776 (N_24776,N_24716,N_24741);
xor U24777 (N_24777,N_24680,N_24560);
or U24778 (N_24778,N_24508,N_24691);
nand U24779 (N_24779,N_24597,N_24555);
nand U24780 (N_24780,N_24613,N_24565);
and U24781 (N_24781,N_24646,N_24590);
and U24782 (N_24782,N_24552,N_24575);
and U24783 (N_24783,N_24571,N_24600);
xor U24784 (N_24784,N_24636,N_24501);
and U24785 (N_24785,N_24503,N_24664);
nor U24786 (N_24786,N_24553,N_24549);
xnor U24787 (N_24787,N_24712,N_24670);
or U24788 (N_24788,N_24667,N_24707);
nor U24789 (N_24789,N_24577,N_24643);
nor U24790 (N_24790,N_24730,N_24732);
nor U24791 (N_24791,N_24609,N_24693);
xor U24792 (N_24792,N_24685,N_24502);
nor U24793 (N_24793,N_24551,N_24713);
or U24794 (N_24794,N_24731,N_24599);
nor U24795 (N_24795,N_24525,N_24535);
nor U24796 (N_24796,N_24633,N_24621);
nand U24797 (N_24797,N_24715,N_24516);
and U24798 (N_24798,N_24607,N_24701);
nor U24799 (N_24799,N_24729,N_24554);
or U24800 (N_24800,N_24724,N_24572);
and U24801 (N_24801,N_24620,N_24672);
xor U24802 (N_24802,N_24737,N_24576);
nand U24803 (N_24803,N_24524,N_24531);
or U24804 (N_24804,N_24589,N_24566);
nand U24805 (N_24805,N_24648,N_24637);
xnor U24806 (N_24806,N_24656,N_24626);
and U24807 (N_24807,N_24528,N_24542);
and U24808 (N_24808,N_24661,N_24649);
and U24809 (N_24809,N_24562,N_24641);
nor U24810 (N_24810,N_24588,N_24748);
and U24811 (N_24811,N_24507,N_24709);
and U24812 (N_24812,N_24666,N_24738);
or U24813 (N_24813,N_24678,N_24697);
and U24814 (N_24814,N_24580,N_24736);
nand U24815 (N_24815,N_24579,N_24728);
nor U24816 (N_24816,N_24504,N_24608);
nor U24817 (N_24817,N_24511,N_24585);
nor U24818 (N_24818,N_24546,N_24710);
or U24819 (N_24819,N_24533,N_24509);
or U24820 (N_24820,N_24735,N_24632);
or U24821 (N_24821,N_24548,N_24652);
nand U24822 (N_24822,N_24594,N_24658);
nand U24823 (N_24823,N_24746,N_24510);
xor U24824 (N_24824,N_24581,N_24618);
and U24825 (N_24825,N_24723,N_24521);
or U24826 (N_24826,N_24653,N_24512);
and U24827 (N_24827,N_24543,N_24714);
xor U24828 (N_24828,N_24660,N_24700);
xnor U24829 (N_24829,N_24561,N_24642);
or U24830 (N_24830,N_24612,N_24668);
nand U24831 (N_24831,N_24645,N_24734);
nand U24832 (N_24832,N_24556,N_24634);
nand U24833 (N_24833,N_24699,N_24743);
or U24834 (N_24834,N_24550,N_24695);
or U24835 (N_24835,N_24674,N_24616);
and U24836 (N_24836,N_24513,N_24692);
xor U24837 (N_24837,N_24630,N_24647);
nor U24838 (N_24838,N_24733,N_24617);
nand U24839 (N_24839,N_24703,N_24619);
and U24840 (N_24840,N_24665,N_24727);
nand U24841 (N_24841,N_24557,N_24719);
nor U24842 (N_24842,N_24615,N_24726);
and U24843 (N_24843,N_24544,N_24717);
and U24844 (N_24844,N_24547,N_24603);
nand U24845 (N_24845,N_24704,N_24625);
nand U24846 (N_24846,N_24573,N_24627);
or U24847 (N_24847,N_24505,N_24530);
xnor U24848 (N_24848,N_24651,N_24629);
nand U24849 (N_24849,N_24669,N_24606);
nor U24850 (N_24850,N_24679,N_24740);
nand U24851 (N_24851,N_24624,N_24519);
or U24852 (N_24852,N_24635,N_24523);
or U24853 (N_24853,N_24711,N_24537);
xor U24854 (N_24854,N_24578,N_24677);
nand U24855 (N_24855,N_24568,N_24640);
and U24856 (N_24856,N_24526,N_24529);
nand U24857 (N_24857,N_24541,N_24718);
nor U24858 (N_24858,N_24558,N_24598);
nor U24859 (N_24859,N_24682,N_24582);
nand U24860 (N_24860,N_24506,N_24602);
and U24861 (N_24861,N_24540,N_24604);
nor U24862 (N_24862,N_24605,N_24690);
or U24863 (N_24863,N_24688,N_24689);
nor U24864 (N_24864,N_24721,N_24739);
xor U24865 (N_24865,N_24683,N_24569);
or U24866 (N_24866,N_24745,N_24696);
xnor U24867 (N_24867,N_24563,N_24610);
nand U24868 (N_24868,N_24517,N_24532);
nor U24869 (N_24869,N_24644,N_24514);
nand U24870 (N_24870,N_24638,N_24663);
or U24871 (N_24871,N_24681,N_24574);
xor U24872 (N_24872,N_24744,N_24622);
nand U24873 (N_24873,N_24655,N_24536);
nor U24874 (N_24874,N_24527,N_24694);
nor U24875 (N_24875,N_24628,N_24573);
or U24876 (N_24876,N_24540,N_24586);
nand U24877 (N_24877,N_24730,N_24632);
nor U24878 (N_24878,N_24629,N_24722);
xnor U24879 (N_24879,N_24553,N_24691);
xnor U24880 (N_24880,N_24616,N_24555);
and U24881 (N_24881,N_24600,N_24627);
and U24882 (N_24882,N_24561,N_24686);
or U24883 (N_24883,N_24541,N_24733);
and U24884 (N_24884,N_24524,N_24618);
nor U24885 (N_24885,N_24583,N_24647);
xor U24886 (N_24886,N_24702,N_24604);
nor U24887 (N_24887,N_24653,N_24631);
nand U24888 (N_24888,N_24718,N_24616);
nand U24889 (N_24889,N_24737,N_24525);
and U24890 (N_24890,N_24531,N_24559);
nand U24891 (N_24891,N_24686,N_24622);
nor U24892 (N_24892,N_24581,N_24690);
and U24893 (N_24893,N_24647,N_24506);
xnor U24894 (N_24894,N_24524,N_24563);
nor U24895 (N_24895,N_24669,N_24566);
and U24896 (N_24896,N_24749,N_24586);
xnor U24897 (N_24897,N_24728,N_24646);
xor U24898 (N_24898,N_24554,N_24512);
and U24899 (N_24899,N_24690,N_24533);
and U24900 (N_24900,N_24626,N_24637);
nor U24901 (N_24901,N_24550,N_24682);
or U24902 (N_24902,N_24607,N_24525);
and U24903 (N_24903,N_24568,N_24604);
nor U24904 (N_24904,N_24553,N_24568);
nor U24905 (N_24905,N_24523,N_24656);
nand U24906 (N_24906,N_24585,N_24601);
and U24907 (N_24907,N_24667,N_24532);
nor U24908 (N_24908,N_24514,N_24606);
xnor U24909 (N_24909,N_24667,N_24515);
nand U24910 (N_24910,N_24733,N_24511);
xnor U24911 (N_24911,N_24651,N_24563);
nand U24912 (N_24912,N_24699,N_24573);
xor U24913 (N_24913,N_24504,N_24575);
and U24914 (N_24914,N_24576,N_24651);
xor U24915 (N_24915,N_24573,N_24567);
or U24916 (N_24916,N_24652,N_24698);
and U24917 (N_24917,N_24602,N_24505);
and U24918 (N_24918,N_24560,N_24593);
or U24919 (N_24919,N_24626,N_24663);
nor U24920 (N_24920,N_24542,N_24734);
xor U24921 (N_24921,N_24743,N_24581);
and U24922 (N_24922,N_24687,N_24508);
xnor U24923 (N_24923,N_24617,N_24590);
or U24924 (N_24924,N_24540,N_24579);
nor U24925 (N_24925,N_24731,N_24697);
nor U24926 (N_24926,N_24578,N_24685);
xnor U24927 (N_24927,N_24623,N_24711);
nand U24928 (N_24928,N_24521,N_24548);
xnor U24929 (N_24929,N_24529,N_24519);
nor U24930 (N_24930,N_24588,N_24529);
or U24931 (N_24931,N_24588,N_24630);
nand U24932 (N_24932,N_24659,N_24718);
or U24933 (N_24933,N_24585,N_24527);
and U24934 (N_24934,N_24700,N_24505);
or U24935 (N_24935,N_24550,N_24726);
nand U24936 (N_24936,N_24663,N_24540);
nor U24937 (N_24937,N_24669,N_24660);
and U24938 (N_24938,N_24546,N_24688);
nand U24939 (N_24939,N_24581,N_24534);
xnor U24940 (N_24940,N_24681,N_24607);
xor U24941 (N_24941,N_24542,N_24609);
or U24942 (N_24942,N_24528,N_24737);
or U24943 (N_24943,N_24639,N_24602);
and U24944 (N_24944,N_24702,N_24681);
nor U24945 (N_24945,N_24683,N_24637);
nor U24946 (N_24946,N_24513,N_24543);
nand U24947 (N_24947,N_24630,N_24575);
and U24948 (N_24948,N_24643,N_24541);
nor U24949 (N_24949,N_24612,N_24534);
and U24950 (N_24950,N_24652,N_24710);
nand U24951 (N_24951,N_24636,N_24590);
xor U24952 (N_24952,N_24694,N_24698);
nand U24953 (N_24953,N_24693,N_24570);
xnor U24954 (N_24954,N_24747,N_24566);
nand U24955 (N_24955,N_24723,N_24506);
or U24956 (N_24956,N_24733,N_24597);
or U24957 (N_24957,N_24636,N_24561);
and U24958 (N_24958,N_24608,N_24581);
xnor U24959 (N_24959,N_24620,N_24648);
nor U24960 (N_24960,N_24625,N_24708);
nor U24961 (N_24961,N_24692,N_24661);
nand U24962 (N_24962,N_24724,N_24706);
xor U24963 (N_24963,N_24588,N_24604);
nor U24964 (N_24964,N_24520,N_24563);
nor U24965 (N_24965,N_24680,N_24638);
nor U24966 (N_24966,N_24549,N_24534);
or U24967 (N_24967,N_24640,N_24663);
nor U24968 (N_24968,N_24732,N_24527);
or U24969 (N_24969,N_24592,N_24723);
nor U24970 (N_24970,N_24520,N_24707);
nand U24971 (N_24971,N_24559,N_24688);
nor U24972 (N_24972,N_24509,N_24551);
or U24973 (N_24973,N_24666,N_24741);
and U24974 (N_24974,N_24548,N_24534);
and U24975 (N_24975,N_24703,N_24642);
xor U24976 (N_24976,N_24691,N_24700);
nor U24977 (N_24977,N_24531,N_24523);
and U24978 (N_24978,N_24544,N_24500);
and U24979 (N_24979,N_24705,N_24686);
nor U24980 (N_24980,N_24579,N_24734);
nor U24981 (N_24981,N_24561,N_24511);
nand U24982 (N_24982,N_24700,N_24655);
or U24983 (N_24983,N_24635,N_24563);
nor U24984 (N_24984,N_24724,N_24642);
or U24985 (N_24985,N_24631,N_24583);
xnor U24986 (N_24986,N_24561,N_24739);
xor U24987 (N_24987,N_24700,N_24686);
nor U24988 (N_24988,N_24658,N_24747);
xor U24989 (N_24989,N_24558,N_24533);
or U24990 (N_24990,N_24565,N_24656);
or U24991 (N_24991,N_24708,N_24503);
nor U24992 (N_24992,N_24554,N_24607);
nor U24993 (N_24993,N_24743,N_24528);
nor U24994 (N_24994,N_24644,N_24719);
nand U24995 (N_24995,N_24540,N_24605);
nor U24996 (N_24996,N_24621,N_24608);
nand U24997 (N_24997,N_24569,N_24738);
xor U24998 (N_24998,N_24581,N_24706);
nor U24999 (N_24999,N_24650,N_24591);
xor UO_0 (O_0,N_24803,N_24827);
nor UO_1 (O_1,N_24882,N_24946);
and UO_2 (O_2,N_24865,N_24980);
nand UO_3 (O_3,N_24780,N_24752);
xnor UO_4 (O_4,N_24817,N_24923);
nor UO_5 (O_5,N_24836,N_24996);
xor UO_6 (O_6,N_24816,N_24958);
xnor UO_7 (O_7,N_24810,N_24928);
and UO_8 (O_8,N_24790,N_24753);
nand UO_9 (O_9,N_24763,N_24758);
nor UO_10 (O_10,N_24990,N_24921);
nand UO_11 (O_11,N_24801,N_24786);
nand UO_12 (O_12,N_24789,N_24968);
xnor UO_13 (O_13,N_24830,N_24911);
or UO_14 (O_14,N_24840,N_24893);
nor UO_15 (O_15,N_24945,N_24976);
nand UO_16 (O_16,N_24957,N_24807);
or UO_17 (O_17,N_24760,N_24851);
and UO_18 (O_18,N_24767,N_24906);
and UO_19 (O_19,N_24795,N_24787);
xor UO_20 (O_20,N_24779,N_24883);
xor UO_21 (O_21,N_24991,N_24890);
xnor UO_22 (O_22,N_24954,N_24940);
and UO_23 (O_23,N_24860,N_24988);
and UO_24 (O_24,N_24878,N_24839);
nand UO_25 (O_25,N_24873,N_24853);
nor UO_26 (O_26,N_24794,N_24825);
nand UO_27 (O_27,N_24821,N_24927);
and UO_28 (O_28,N_24899,N_24918);
nand UO_29 (O_29,N_24777,N_24887);
nor UO_30 (O_30,N_24997,N_24838);
nor UO_31 (O_31,N_24956,N_24811);
and UO_32 (O_32,N_24897,N_24755);
nand UO_33 (O_33,N_24778,N_24872);
or UO_34 (O_34,N_24953,N_24986);
nand UO_35 (O_35,N_24805,N_24866);
xor UO_36 (O_36,N_24796,N_24765);
xnor UO_37 (O_37,N_24961,N_24885);
and UO_38 (O_38,N_24857,N_24892);
nor UO_39 (O_39,N_24869,N_24971);
nor UO_40 (O_40,N_24783,N_24861);
and UO_41 (O_41,N_24868,N_24867);
or UO_42 (O_42,N_24877,N_24774);
or UO_43 (O_43,N_24973,N_24802);
or UO_44 (O_44,N_24907,N_24960);
nand UO_45 (O_45,N_24925,N_24913);
xor UO_46 (O_46,N_24999,N_24814);
nor UO_47 (O_47,N_24818,N_24766);
nor UO_48 (O_48,N_24895,N_24750);
or UO_49 (O_49,N_24959,N_24870);
xor UO_50 (O_50,N_24875,N_24813);
xor UO_51 (O_51,N_24942,N_24962);
nand UO_52 (O_52,N_24965,N_24936);
and UO_53 (O_53,N_24770,N_24823);
nor UO_54 (O_54,N_24975,N_24979);
and UO_55 (O_55,N_24987,N_24995);
xor UO_56 (O_56,N_24947,N_24854);
or UO_57 (O_57,N_24948,N_24841);
or UO_58 (O_58,N_24985,N_24799);
or UO_59 (O_59,N_24792,N_24993);
or UO_60 (O_60,N_24879,N_24800);
nor UO_61 (O_61,N_24884,N_24915);
or UO_62 (O_62,N_24889,N_24939);
xnor UO_63 (O_63,N_24924,N_24917);
nand UO_64 (O_64,N_24908,N_24919);
or UO_65 (O_65,N_24797,N_24930);
and UO_66 (O_66,N_24769,N_24757);
or UO_67 (O_67,N_24819,N_24754);
and UO_68 (O_68,N_24829,N_24863);
nand UO_69 (O_69,N_24934,N_24798);
nand UO_70 (O_70,N_24762,N_24859);
xor UO_71 (O_71,N_24929,N_24989);
or UO_72 (O_72,N_24828,N_24933);
and UO_73 (O_73,N_24848,N_24970);
or UO_74 (O_74,N_24808,N_24773);
xnor UO_75 (O_75,N_24864,N_24951);
nand UO_76 (O_76,N_24984,N_24888);
and UO_77 (O_77,N_24983,N_24920);
nor UO_78 (O_78,N_24922,N_24941);
or UO_79 (O_79,N_24806,N_24782);
xnor UO_80 (O_80,N_24912,N_24855);
xor UO_81 (O_81,N_24943,N_24771);
xor UO_82 (O_82,N_24931,N_24966);
nand UO_83 (O_83,N_24880,N_24998);
nand UO_84 (O_84,N_24916,N_24972);
or UO_85 (O_85,N_24764,N_24926);
nor UO_86 (O_86,N_24932,N_24756);
and UO_87 (O_87,N_24849,N_24898);
or UO_88 (O_88,N_24905,N_24886);
nor UO_89 (O_89,N_24751,N_24793);
or UO_90 (O_90,N_24791,N_24775);
and UO_91 (O_91,N_24852,N_24910);
nor UO_92 (O_92,N_24812,N_24901);
or UO_93 (O_93,N_24759,N_24978);
nor UO_94 (O_94,N_24761,N_24781);
xor UO_95 (O_95,N_24967,N_24862);
and UO_96 (O_96,N_24833,N_24955);
nand UO_97 (O_97,N_24842,N_24772);
nand UO_98 (O_98,N_24937,N_24831);
and UO_99 (O_99,N_24820,N_24850);
nor UO_100 (O_100,N_24824,N_24834);
or UO_101 (O_101,N_24856,N_24949);
or UO_102 (O_102,N_24904,N_24969);
xor UO_103 (O_103,N_24964,N_24843);
xnor UO_104 (O_104,N_24891,N_24871);
or UO_105 (O_105,N_24952,N_24981);
xnor UO_106 (O_106,N_24845,N_24896);
nor UO_107 (O_107,N_24902,N_24788);
xnor UO_108 (O_108,N_24900,N_24914);
or UO_109 (O_109,N_24903,N_24963);
and UO_110 (O_110,N_24858,N_24992);
or UO_111 (O_111,N_24822,N_24909);
nand UO_112 (O_112,N_24768,N_24935);
nor UO_113 (O_113,N_24844,N_24826);
xnor UO_114 (O_114,N_24881,N_24846);
nand UO_115 (O_115,N_24950,N_24837);
xor UO_116 (O_116,N_24994,N_24785);
or UO_117 (O_117,N_24944,N_24809);
nor UO_118 (O_118,N_24776,N_24938);
or UO_119 (O_119,N_24982,N_24974);
nand UO_120 (O_120,N_24977,N_24894);
or UO_121 (O_121,N_24847,N_24815);
and UO_122 (O_122,N_24874,N_24835);
and UO_123 (O_123,N_24876,N_24784);
xnor UO_124 (O_124,N_24804,N_24832);
nand UO_125 (O_125,N_24889,N_24787);
xor UO_126 (O_126,N_24837,N_24806);
and UO_127 (O_127,N_24924,N_24936);
and UO_128 (O_128,N_24829,N_24905);
and UO_129 (O_129,N_24884,N_24879);
and UO_130 (O_130,N_24879,N_24871);
and UO_131 (O_131,N_24760,N_24770);
nor UO_132 (O_132,N_24912,N_24931);
nand UO_133 (O_133,N_24900,N_24759);
xor UO_134 (O_134,N_24909,N_24809);
or UO_135 (O_135,N_24916,N_24759);
nand UO_136 (O_136,N_24771,N_24758);
nand UO_137 (O_137,N_24837,N_24845);
nor UO_138 (O_138,N_24911,N_24939);
xnor UO_139 (O_139,N_24853,N_24828);
and UO_140 (O_140,N_24881,N_24787);
nor UO_141 (O_141,N_24881,N_24920);
xor UO_142 (O_142,N_24905,N_24968);
or UO_143 (O_143,N_24782,N_24944);
nand UO_144 (O_144,N_24850,N_24848);
and UO_145 (O_145,N_24953,N_24854);
nor UO_146 (O_146,N_24781,N_24914);
and UO_147 (O_147,N_24829,N_24847);
and UO_148 (O_148,N_24940,N_24989);
or UO_149 (O_149,N_24991,N_24864);
nor UO_150 (O_150,N_24881,N_24759);
and UO_151 (O_151,N_24979,N_24767);
or UO_152 (O_152,N_24940,N_24864);
or UO_153 (O_153,N_24992,N_24925);
nand UO_154 (O_154,N_24810,N_24945);
nor UO_155 (O_155,N_24976,N_24815);
or UO_156 (O_156,N_24772,N_24811);
nand UO_157 (O_157,N_24930,N_24897);
nor UO_158 (O_158,N_24810,N_24762);
nand UO_159 (O_159,N_24840,N_24997);
nor UO_160 (O_160,N_24921,N_24784);
nand UO_161 (O_161,N_24798,N_24956);
nor UO_162 (O_162,N_24961,N_24787);
nor UO_163 (O_163,N_24964,N_24968);
xor UO_164 (O_164,N_24778,N_24896);
xnor UO_165 (O_165,N_24862,N_24979);
nand UO_166 (O_166,N_24908,N_24890);
xor UO_167 (O_167,N_24866,N_24841);
nor UO_168 (O_168,N_24837,N_24750);
xor UO_169 (O_169,N_24925,N_24838);
nor UO_170 (O_170,N_24822,N_24854);
and UO_171 (O_171,N_24961,N_24834);
nor UO_172 (O_172,N_24911,N_24750);
xor UO_173 (O_173,N_24847,N_24761);
xnor UO_174 (O_174,N_24822,N_24933);
nand UO_175 (O_175,N_24778,N_24933);
nor UO_176 (O_176,N_24804,N_24940);
xnor UO_177 (O_177,N_24794,N_24833);
nor UO_178 (O_178,N_24938,N_24753);
nand UO_179 (O_179,N_24867,N_24964);
or UO_180 (O_180,N_24945,N_24792);
nand UO_181 (O_181,N_24985,N_24978);
nand UO_182 (O_182,N_24864,N_24804);
nor UO_183 (O_183,N_24854,N_24792);
nand UO_184 (O_184,N_24803,N_24901);
and UO_185 (O_185,N_24819,N_24924);
and UO_186 (O_186,N_24777,N_24766);
or UO_187 (O_187,N_24761,N_24952);
and UO_188 (O_188,N_24768,N_24885);
or UO_189 (O_189,N_24906,N_24761);
nand UO_190 (O_190,N_24825,N_24850);
and UO_191 (O_191,N_24997,N_24992);
nand UO_192 (O_192,N_24818,N_24830);
or UO_193 (O_193,N_24842,N_24852);
and UO_194 (O_194,N_24859,N_24805);
nor UO_195 (O_195,N_24771,N_24857);
nand UO_196 (O_196,N_24906,N_24957);
nand UO_197 (O_197,N_24889,N_24995);
or UO_198 (O_198,N_24806,N_24948);
and UO_199 (O_199,N_24895,N_24813);
or UO_200 (O_200,N_24998,N_24785);
nand UO_201 (O_201,N_24777,N_24769);
xor UO_202 (O_202,N_24952,N_24965);
nor UO_203 (O_203,N_24816,N_24957);
nor UO_204 (O_204,N_24986,N_24876);
nand UO_205 (O_205,N_24812,N_24784);
nor UO_206 (O_206,N_24918,N_24796);
nand UO_207 (O_207,N_24897,N_24807);
nor UO_208 (O_208,N_24949,N_24756);
and UO_209 (O_209,N_24967,N_24917);
xnor UO_210 (O_210,N_24863,N_24932);
and UO_211 (O_211,N_24956,N_24792);
and UO_212 (O_212,N_24836,N_24966);
nand UO_213 (O_213,N_24801,N_24861);
nand UO_214 (O_214,N_24945,N_24956);
nand UO_215 (O_215,N_24867,N_24783);
and UO_216 (O_216,N_24897,N_24945);
nand UO_217 (O_217,N_24875,N_24867);
nand UO_218 (O_218,N_24806,N_24794);
nor UO_219 (O_219,N_24982,N_24795);
xnor UO_220 (O_220,N_24766,N_24888);
nor UO_221 (O_221,N_24929,N_24882);
xor UO_222 (O_222,N_24843,N_24869);
xnor UO_223 (O_223,N_24898,N_24907);
xor UO_224 (O_224,N_24815,N_24929);
nand UO_225 (O_225,N_24823,N_24934);
xnor UO_226 (O_226,N_24987,N_24932);
or UO_227 (O_227,N_24836,N_24907);
and UO_228 (O_228,N_24919,N_24787);
nor UO_229 (O_229,N_24798,N_24921);
and UO_230 (O_230,N_24900,N_24938);
xor UO_231 (O_231,N_24987,N_24847);
xnor UO_232 (O_232,N_24791,N_24804);
xnor UO_233 (O_233,N_24767,N_24904);
and UO_234 (O_234,N_24822,N_24752);
xnor UO_235 (O_235,N_24886,N_24866);
nor UO_236 (O_236,N_24791,N_24849);
and UO_237 (O_237,N_24959,N_24905);
xnor UO_238 (O_238,N_24906,N_24844);
or UO_239 (O_239,N_24843,N_24805);
xor UO_240 (O_240,N_24794,N_24815);
and UO_241 (O_241,N_24752,N_24784);
and UO_242 (O_242,N_24818,N_24973);
xnor UO_243 (O_243,N_24937,N_24874);
nand UO_244 (O_244,N_24911,N_24759);
or UO_245 (O_245,N_24835,N_24975);
xnor UO_246 (O_246,N_24754,N_24921);
nor UO_247 (O_247,N_24882,N_24907);
and UO_248 (O_248,N_24832,N_24989);
xnor UO_249 (O_249,N_24952,N_24883);
and UO_250 (O_250,N_24767,N_24756);
or UO_251 (O_251,N_24945,N_24841);
or UO_252 (O_252,N_24940,N_24772);
and UO_253 (O_253,N_24787,N_24772);
and UO_254 (O_254,N_24771,N_24814);
nor UO_255 (O_255,N_24814,N_24760);
or UO_256 (O_256,N_24886,N_24891);
nand UO_257 (O_257,N_24753,N_24964);
nand UO_258 (O_258,N_24818,N_24993);
nor UO_259 (O_259,N_24914,N_24986);
nor UO_260 (O_260,N_24760,N_24929);
xor UO_261 (O_261,N_24846,N_24987);
and UO_262 (O_262,N_24923,N_24994);
and UO_263 (O_263,N_24872,N_24791);
and UO_264 (O_264,N_24895,N_24851);
nor UO_265 (O_265,N_24875,N_24926);
nor UO_266 (O_266,N_24959,N_24963);
xor UO_267 (O_267,N_24975,N_24964);
and UO_268 (O_268,N_24951,N_24922);
nand UO_269 (O_269,N_24971,N_24922);
and UO_270 (O_270,N_24933,N_24947);
and UO_271 (O_271,N_24913,N_24982);
nor UO_272 (O_272,N_24832,N_24766);
and UO_273 (O_273,N_24915,N_24961);
and UO_274 (O_274,N_24782,N_24970);
or UO_275 (O_275,N_24878,N_24939);
and UO_276 (O_276,N_24996,N_24804);
or UO_277 (O_277,N_24985,N_24792);
nand UO_278 (O_278,N_24941,N_24844);
xor UO_279 (O_279,N_24990,N_24927);
and UO_280 (O_280,N_24777,N_24860);
xnor UO_281 (O_281,N_24913,N_24877);
or UO_282 (O_282,N_24811,N_24832);
nor UO_283 (O_283,N_24834,N_24889);
nand UO_284 (O_284,N_24996,N_24806);
nand UO_285 (O_285,N_24930,N_24970);
xor UO_286 (O_286,N_24853,N_24914);
or UO_287 (O_287,N_24988,N_24953);
and UO_288 (O_288,N_24842,N_24897);
or UO_289 (O_289,N_24756,N_24912);
and UO_290 (O_290,N_24826,N_24759);
nor UO_291 (O_291,N_24865,N_24797);
nand UO_292 (O_292,N_24862,N_24879);
and UO_293 (O_293,N_24931,N_24948);
xor UO_294 (O_294,N_24874,N_24903);
nor UO_295 (O_295,N_24946,N_24943);
nor UO_296 (O_296,N_24951,N_24846);
or UO_297 (O_297,N_24874,N_24770);
nand UO_298 (O_298,N_24899,N_24932);
and UO_299 (O_299,N_24801,N_24930);
or UO_300 (O_300,N_24957,N_24909);
xnor UO_301 (O_301,N_24929,N_24824);
xnor UO_302 (O_302,N_24866,N_24839);
nand UO_303 (O_303,N_24987,N_24994);
xor UO_304 (O_304,N_24756,N_24974);
or UO_305 (O_305,N_24750,N_24922);
xnor UO_306 (O_306,N_24755,N_24907);
xor UO_307 (O_307,N_24900,N_24758);
and UO_308 (O_308,N_24908,N_24937);
or UO_309 (O_309,N_24983,N_24914);
xnor UO_310 (O_310,N_24809,N_24777);
or UO_311 (O_311,N_24926,N_24765);
and UO_312 (O_312,N_24913,N_24804);
nand UO_313 (O_313,N_24918,N_24815);
nand UO_314 (O_314,N_24995,N_24779);
nand UO_315 (O_315,N_24951,N_24935);
and UO_316 (O_316,N_24973,N_24901);
or UO_317 (O_317,N_24810,N_24877);
and UO_318 (O_318,N_24796,N_24848);
nand UO_319 (O_319,N_24966,N_24801);
nor UO_320 (O_320,N_24908,N_24968);
or UO_321 (O_321,N_24937,N_24797);
or UO_322 (O_322,N_24873,N_24970);
nand UO_323 (O_323,N_24784,N_24875);
or UO_324 (O_324,N_24970,N_24812);
nand UO_325 (O_325,N_24765,N_24916);
nand UO_326 (O_326,N_24894,N_24906);
or UO_327 (O_327,N_24892,N_24932);
nor UO_328 (O_328,N_24762,N_24990);
nor UO_329 (O_329,N_24782,N_24754);
nor UO_330 (O_330,N_24884,N_24971);
and UO_331 (O_331,N_24980,N_24844);
or UO_332 (O_332,N_24910,N_24751);
and UO_333 (O_333,N_24913,N_24809);
or UO_334 (O_334,N_24770,N_24752);
nand UO_335 (O_335,N_24936,N_24805);
nor UO_336 (O_336,N_24981,N_24780);
nand UO_337 (O_337,N_24798,N_24960);
or UO_338 (O_338,N_24946,N_24824);
xor UO_339 (O_339,N_24903,N_24851);
xnor UO_340 (O_340,N_24805,N_24795);
and UO_341 (O_341,N_24950,N_24873);
xor UO_342 (O_342,N_24788,N_24852);
nor UO_343 (O_343,N_24988,N_24875);
nand UO_344 (O_344,N_24887,N_24795);
nand UO_345 (O_345,N_24768,N_24868);
and UO_346 (O_346,N_24971,N_24750);
nor UO_347 (O_347,N_24897,N_24770);
or UO_348 (O_348,N_24958,N_24912);
and UO_349 (O_349,N_24890,N_24975);
nand UO_350 (O_350,N_24996,N_24884);
xor UO_351 (O_351,N_24798,N_24915);
xnor UO_352 (O_352,N_24773,N_24882);
and UO_353 (O_353,N_24771,N_24767);
nand UO_354 (O_354,N_24835,N_24812);
or UO_355 (O_355,N_24922,N_24897);
or UO_356 (O_356,N_24855,N_24979);
or UO_357 (O_357,N_24854,N_24798);
or UO_358 (O_358,N_24780,N_24889);
or UO_359 (O_359,N_24759,N_24898);
nand UO_360 (O_360,N_24868,N_24946);
xor UO_361 (O_361,N_24952,N_24896);
nor UO_362 (O_362,N_24974,N_24876);
nor UO_363 (O_363,N_24828,N_24799);
or UO_364 (O_364,N_24807,N_24845);
nor UO_365 (O_365,N_24820,N_24952);
nand UO_366 (O_366,N_24770,N_24851);
or UO_367 (O_367,N_24981,N_24831);
and UO_368 (O_368,N_24817,N_24770);
xnor UO_369 (O_369,N_24940,N_24803);
xor UO_370 (O_370,N_24884,N_24811);
xnor UO_371 (O_371,N_24935,N_24958);
nor UO_372 (O_372,N_24846,N_24790);
and UO_373 (O_373,N_24873,N_24886);
nand UO_374 (O_374,N_24996,N_24833);
nand UO_375 (O_375,N_24798,N_24932);
nor UO_376 (O_376,N_24780,N_24944);
nor UO_377 (O_377,N_24757,N_24833);
and UO_378 (O_378,N_24970,N_24960);
nor UO_379 (O_379,N_24803,N_24788);
nand UO_380 (O_380,N_24950,N_24921);
or UO_381 (O_381,N_24825,N_24881);
nor UO_382 (O_382,N_24815,N_24779);
nor UO_383 (O_383,N_24884,N_24921);
nand UO_384 (O_384,N_24990,N_24865);
nand UO_385 (O_385,N_24960,N_24989);
nor UO_386 (O_386,N_24939,N_24885);
nand UO_387 (O_387,N_24961,N_24896);
nor UO_388 (O_388,N_24780,N_24922);
nand UO_389 (O_389,N_24945,N_24836);
xnor UO_390 (O_390,N_24859,N_24763);
nand UO_391 (O_391,N_24916,N_24982);
or UO_392 (O_392,N_24952,N_24865);
nand UO_393 (O_393,N_24758,N_24767);
nor UO_394 (O_394,N_24830,N_24974);
or UO_395 (O_395,N_24908,N_24857);
nor UO_396 (O_396,N_24928,N_24831);
nor UO_397 (O_397,N_24879,N_24986);
and UO_398 (O_398,N_24990,N_24884);
nor UO_399 (O_399,N_24962,N_24883);
xor UO_400 (O_400,N_24765,N_24831);
xnor UO_401 (O_401,N_24846,N_24974);
xnor UO_402 (O_402,N_24976,N_24812);
nor UO_403 (O_403,N_24887,N_24947);
nor UO_404 (O_404,N_24954,N_24925);
and UO_405 (O_405,N_24915,N_24797);
xor UO_406 (O_406,N_24837,N_24846);
and UO_407 (O_407,N_24851,N_24972);
or UO_408 (O_408,N_24899,N_24875);
nand UO_409 (O_409,N_24950,N_24751);
nand UO_410 (O_410,N_24808,N_24888);
or UO_411 (O_411,N_24873,N_24770);
xnor UO_412 (O_412,N_24828,N_24870);
or UO_413 (O_413,N_24988,N_24905);
nand UO_414 (O_414,N_24952,N_24829);
and UO_415 (O_415,N_24901,N_24873);
xnor UO_416 (O_416,N_24843,N_24770);
nand UO_417 (O_417,N_24966,N_24807);
nor UO_418 (O_418,N_24764,N_24884);
and UO_419 (O_419,N_24992,N_24921);
nand UO_420 (O_420,N_24875,N_24915);
xnor UO_421 (O_421,N_24835,N_24960);
xor UO_422 (O_422,N_24762,N_24802);
nor UO_423 (O_423,N_24926,N_24854);
nand UO_424 (O_424,N_24792,N_24927);
xnor UO_425 (O_425,N_24903,N_24987);
nand UO_426 (O_426,N_24974,N_24986);
xor UO_427 (O_427,N_24970,N_24906);
xnor UO_428 (O_428,N_24857,N_24936);
and UO_429 (O_429,N_24825,N_24883);
nor UO_430 (O_430,N_24964,N_24798);
nand UO_431 (O_431,N_24990,N_24883);
nand UO_432 (O_432,N_24962,N_24956);
and UO_433 (O_433,N_24752,N_24958);
or UO_434 (O_434,N_24836,N_24872);
and UO_435 (O_435,N_24841,N_24981);
nand UO_436 (O_436,N_24766,N_24885);
nand UO_437 (O_437,N_24813,N_24814);
or UO_438 (O_438,N_24885,N_24860);
or UO_439 (O_439,N_24772,N_24849);
nor UO_440 (O_440,N_24776,N_24787);
nor UO_441 (O_441,N_24800,N_24991);
nor UO_442 (O_442,N_24758,N_24815);
nor UO_443 (O_443,N_24767,N_24968);
nor UO_444 (O_444,N_24870,N_24940);
nand UO_445 (O_445,N_24841,N_24894);
nor UO_446 (O_446,N_24764,N_24971);
nor UO_447 (O_447,N_24993,N_24765);
or UO_448 (O_448,N_24837,N_24824);
or UO_449 (O_449,N_24961,N_24963);
or UO_450 (O_450,N_24772,N_24835);
nand UO_451 (O_451,N_24993,N_24801);
xnor UO_452 (O_452,N_24780,N_24928);
nand UO_453 (O_453,N_24853,N_24885);
and UO_454 (O_454,N_24900,N_24999);
xnor UO_455 (O_455,N_24841,N_24773);
xor UO_456 (O_456,N_24998,N_24853);
nor UO_457 (O_457,N_24960,N_24875);
xnor UO_458 (O_458,N_24826,N_24885);
or UO_459 (O_459,N_24891,N_24986);
and UO_460 (O_460,N_24869,N_24769);
nor UO_461 (O_461,N_24820,N_24944);
xor UO_462 (O_462,N_24864,N_24993);
or UO_463 (O_463,N_24858,N_24831);
nand UO_464 (O_464,N_24915,N_24983);
and UO_465 (O_465,N_24826,N_24754);
and UO_466 (O_466,N_24773,N_24750);
or UO_467 (O_467,N_24849,N_24753);
and UO_468 (O_468,N_24869,N_24988);
and UO_469 (O_469,N_24768,N_24919);
and UO_470 (O_470,N_24936,N_24766);
nand UO_471 (O_471,N_24792,N_24791);
and UO_472 (O_472,N_24864,N_24985);
nor UO_473 (O_473,N_24961,N_24843);
nand UO_474 (O_474,N_24889,N_24959);
or UO_475 (O_475,N_24871,N_24967);
nand UO_476 (O_476,N_24819,N_24946);
xnor UO_477 (O_477,N_24834,N_24926);
and UO_478 (O_478,N_24943,N_24760);
and UO_479 (O_479,N_24814,N_24929);
xor UO_480 (O_480,N_24966,N_24850);
or UO_481 (O_481,N_24844,N_24815);
and UO_482 (O_482,N_24829,N_24796);
nand UO_483 (O_483,N_24823,N_24828);
or UO_484 (O_484,N_24952,N_24780);
and UO_485 (O_485,N_24968,N_24979);
xnor UO_486 (O_486,N_24974,N_24814);
or UO_487 (O_487,N_24817,N_24823);
nand UO_488 (O_488,N_24821,N_24915);
nor UO_489 (O_489,N_24793,N_24769);
nand UO_490 (O_490,N_24886,N_24942);
nand UO_491 (O_491,N_24990,N_24773);
nor UO_492 (O_492,N_24812,N_24881);
xor UO_493 (O_493,N_24804,N_24838);
or UO_494 (O_494,N_24965,N_24979);
and UO_495 (O_495,N_24858,N_24891);
and UO_496 (O_496,N_24892,N_24996);
xor UO_497 (O_497,N_24887,N_24755);
xnor UO_498 (O_498,N_24789,N_24941);
xor UO_499 (O_499,N_24800,N_24790);
nand UO_500 (O_500,N_24809,N_24986);
nand UO_501 (O_501,N_24757,N_24795);
or UO_502 (O_502,N_24998,N_24807);
and UO_503 (O_503,N_24890,N_24902);
and UO_504 (O_504,N_24870,N_24805);
nor UO_505 (O_505,N_24915,N_24870);
or UO_506 (O_506,N_24795,N_24908);
and UO_507 (O_507,N_24970,N_24775);
and UO_508 (O_508,N_24887,N_24939);
nand UO_509 (O_509,N_24926,N_24802);
and UO_510 (O_510,N_24787,N_24761);
or UO_511 (O_511,N_24755,N_24758);
nor UO_512 (O_512,N_24803,N_24889);
xor UO_513 (O_513,N_24780,N_24987);
nor UO_514 (O_514,N_24800,N_24920);
and UO_515 (O_515,N_24886,N_24926);
xnor UO_516 (O_516,N_24964,N_24862);
xnor UO_517 (O_517,N_24839,N_24894);
xnor UO_518 (O_518,N_24906,N_24859);
or UO_519 (O_519,N_24815,N_24891);
nand UO_520 (O_520,N_24822,N_24857);
or UO_521 (O_521,N_24793,N_24858);
and UO_522 (O_522,N_24809,N_24984);
and UO_523 (O_523,N_24889,N_24852);
nor UO_524 (O_524,N_24901,N_24869);
and UO_525 (O_525,N_24871,N_24945);
or UO_526 (O_526,N_24985,N_24822);
nand UO_527 (O_527,N_24994,N_24997);
nor UO_528 (O_528,N_24796,N_24777);
nor UO_529 (O_529,N_24911,N_24984);
or UO_530 (O_530,N_24919,N_24999);
xnor UO_531 (O_531,N_24910,N_24819);
nand UO_532 (O_532,N_24918,N_24765);
nand UO_533 (O_533,N_24780,N_24878);
xnor UO_534 (O_534,N_24787,N_24918);
nor UO_535 (O_535,N_24965,N_24939);
nor UO_536 (O_536,N_24825,N_24870);
xor UO_537 (O_537,N_24771,N_24855);
and UO_538 (O_538,N_24842,N_24783);
nand UO_539 (O_539,N_24997,N_24822);
or UO_540 (O_540,N_24987,N_24839);
nor UO_541 (O_541,N_24839,N_24854);
nand UO_542 (O_542,N_24985,N_24923);
nand UO_543 (O_543,N_24814,N_24886);
or UO_544 (O_544,N_24776,N_24998);
xnor UO_545 (O_545,N_24816,N_24913);
nor UO_546 (O_546,N_24993,N_24914);
nor UO_547 (O_547,N_24761,N_24928);
and UO_548 (O_548,N_24982,N_24900);
or UO_549 (O_549,N_24914,N_24997);
or UO_550 (O_550,N_24920,N_24998);
nor UO_551 (O_551,N_24887,N_24997);
xnor UO_552 (O_552,N_24962,N_24826);
nor UO_553 (O_553,N_24961,N_24856);
and UO_554 (O_554,N_24918,N_24925);
or UO_555 (O_555,N_24998,N_24944);
nor UO_556 (O_556,N_24903,N_24997);
nand UO_557 (O_557,N_24868,N_24765);
or UO_558 (O_558,N_24943,N_24796);
xnor UO_559 (O_559,N_24762,N_24929);
xor UO_560 (O_560,N_24943,N_24994);
nand UO_561 (O_561,N_24991,N_24873);
or UO_562 (O_562,N_24881,N_24949);
nand UO_563 (O_563,N_24958,N_24959);
nor UO_564 (O_564,N_24888,N_24753);
and UO_565 (O_565,N_24918,N_24954);
xor UO_566 (O_566,N_24814,N_24769);
nor UO_567 (O_567,N_24927,N_24855);
xor UO_568 (O_568,N_24868,N_24752);
nand UO_569 (O_569,N_24781,N_24812);
and UO_570 (O_570,N_24895,N_24785);
nand UO_571 (O_571,N_24819,N_24874);
and UO_572 (O_572,N_24929,N_24887);
nand UO_573 (O_573,N_24906,N_24924);
or UO_574 (O_574,N_24993,N_24989);
xnor UO_575 (O_575,N_24931,N_24954);
nand UO_576 (O_576,N_24996,N_24890);
or UO_577 (O_577,N_24981,N_24799);
or UO_578 (O_578,N_24939,N_24907);
nand UO_579 (O_579,N_24894,N_24761);
xnor UO_580 (O_580,N_24856,N_24777);
nor UO_581 (O_581,N_24957,N_24849);
or UO_582 (O_582,N_24941,N_24924);
or UO_583 (O_583,N_24814,N_24866);
and UO_584 (O_584,N_24927,N_24790);
nor UO_585 (O_585,N_24750,N_24942);
or UO_586 (O_586,N_24906,N_24979);
nand UO_587 (O_587,N_24972,N_24885);
xnor UO_588 (O_588,N_24780,N_24848);
and UO_589 (O_589,N_24858,N_24785);
nor UO_590 (O_590,N_24831,N_24814);
and UO_591 (O_591,N_24985,N_24991);
xor UO_592 (O_592,N_24805,N_24903);
nand UO_593 (O_593,N_24869,N_24814);
or UO_594 (O_594,N_24808,N_24781);
xnor UO_595 (O_595,N_24920,N_24986);
nand UO_596 (O_596,N_24776,N_24921);
or UO_597 (O_597,N_24988,N_24787);
and UO_598 (O_598,N_24782,N_24798);
nor UO_599 (O_599,N_24852,N_24933);
nand UO_600 (O_600,N_24924,N_24930);
nor UO_601 (O_601,N_24847,N_24827);
or UO_602 (O_602,N_24828,N_24941);
nor UO_603 (O_603,N_24907,N_24881);
and UO_604 (O_604,N_24965,N_24911);
or UO_605 (O_605,N_24857,N_24850);
xor UO_606 (O_606,N_24949,N_24761);
nand UO_607 (O_607,N_24847,N_24916);
nand UO_608 (O_608,N_24853,N_24947);
nand UO_609 (O_609,N_24942,N_24865);
and UO_610 (O_610,N_24952,N_24890);
nor UO_611 (O_611,N_24816,N_24936);
nand UO_612 (O_612,N_24778,N_24787);
or UO_613 (O_613,N_24807,N_24850);
nand UO_614 (O_614,N_24766,N_24980);
or UO_615 (O_615,N_24793,N_24986);
nor UO_616 (O_616,N_24790,N_24993);
and UO_617 (O_617,N_24836,N_24913);
or UO_618 (O_618,N_24789,N_24869);
xnor UO_619 (O_619,N_24857,N_24905);
and UO_620 (O_620,N_24893,N_24880);
or UO_621 (O_621,N_24877,N_24916);
or UO_622 (O_622,N_24768,N_24982);
nor UO_623 (O_623,N_24862,N_24958);
nor UO_624 (O_624,N_24825,N_24793);
or UO_625 (O_625,N_24914,N_24963);
xnor UO_626 (O_626,N_24760,N_24830);
or UO_627 (O_627,N_24960,N_24756);
or UO_628 (O_628,N_24935,N_24913);
and UO_629 (O_629,N_24815,N_24934);
and UO_630 (O_630,N_24769,N_24987);
xnor UO_631 (O_631,N_24922,N_24807);
and UO_632 (O_632,N_24969,N_24892);
nand UO_633 (O_633,N_24906,N_24774);
xor UO_634 (O_634,N_24952,N_24972);
and UO_635 (O_635,N_24959,N_24972);
nand UO_636 (O_636,N_24980,N_24900);
and UO_637 (O_637,N_24943,N_24801);
nand UO_638 (O_638,N_24774,N_24953);
nor UO_639 (O_639,N_24854,N_24914);
nand UO_640 (O_640,N_24869,N_24937);
and UO_641 (O_641,N_24952,N_24821);
nand UO_642 (O_642,N_24991,N_24779);
nor UO_643 (O_643,N_24884,N_24986);
and UO_644 (O_644,N_24863,N_24972);
nand UO_645 (O_645,N_24883,N_24874);
and UO_646 (O_646,N_24794,N_24813);
nor UO_647 (O_647,N_24970,N_24820);
xnor UO_648 (O_648,N_24863,N_24894);
xnor UO_649 (O_649,N_24961,N_24855);
nor UO_650 (O_650,N_24799,N_24991);
nor UO_651 (O_651,N_24754,N_24803);
nand UO_652 (O_652,N_24956,N_24936);
and UO_653 (O_653,N_24831,N_24862);
xnor UO_654 (O_654,N_24761,N_24992);
or UO_655 (O_655,N_24842,N_24934);
or UO_656 (O_656,N_24904,N_24773);
xnor UO_657 (O_657,N_24795,N_24910);
nor UO_658 (O_658,N_24912,N_24885);
or UO_659 (O_659,N_24911,N_24812);
xnor UO_660 (O_660,N_24864,N_24798);
and UO_661 (O_661,N_24964,N_24850);
and UO_662 (O_662,N_24902,N_24767);
nand UO_663 (O_663,N_24879,N_24822);
xnor UO_664 (O_664,N_24781,N_24966);
xnor UO_665 (O_665,N_24931,N_24950);
xnor UO_666 (O_666,N_24837,N_24803);
and UO_667 (O_667,N_24995,N_24797);
and UO_668 (O_668,N_24898,N_24942);
nand UO_669 (O_669,N_24942,N_24916);
nand UO_670 (O_670,N_24892,N_24910);
or UO_671 (O_671,N_24750,N_24979);
nor UO_672 (O_672,N_24832,N_24834);
xnor UO_673 (O_673,N_24962,N_24911);
and UO_674 (O_674,N_24864,N_24982);
and UO_675 (O_675,N_24769,N_24914);
nand UO_676 (O_676,N_24779,N_24882);
nand UO_677 (O_677,N_24969,N_24975);
nor UO_678 (O_678,N_24758,N_24869);
nand UO_679 (O_679,N_24757,N_24827);
and UO_680 (O_680,N_24820,N_24772);
or UO_681 (O_681,N_24792,N_24807);
nor UO_682 (O_682,N_24936,N_24831);
or UO_683 (O_683,N_24773,N_24949);
nor UO_684 (O_684,N_24978,N_24993);
xor UO_685 (O_685,N_24760,N_24940);
nand UO_686 (O_686,N_24901,N_24896);
and UO_687 (O_687,N_24826,N_24827);
or UO_688 (O_688,N_24957,N_24894);
nor UO_689 (O_689,N_24867,N_24762);
nor UO_690 (O_690,N_24794,N_24899);
nor UO_691 (O_691,N_24776,N_24980);
or UO_692 (O_692,N_24811,N_24890);
nor UO_693 (O_693,N_24875,N_24762);
or UO_694 (O_694,N_24773,N_24963);
nor UO_695 (O_695,N_24825,N_24897);
nor UO_696 (O_696,N_24907,N_24969);
or UO_697 (O_697,N_24780,N_24894);
nor UO_698 (O_698,N_24820,N_24764);
nor UO_699 (O_699,N_24878,N_24819);
nor UO_700 (O_700,N_24975,N_24836);
xor UO_701 (O_701,N_24954,N_24834);
or UO_702 (O_702,N_24936,N_24898);
nand UO_703 (O_703,N_24780,N_24982);
or UO_704 (O_704,N_24888,N_24823);
and UO_705 (O_705,N_24894,N_24996);
and UO_706 (O_706,N_24835,N_24796);
nor UO_707 (O_707,N_24939,N_24843);
nand UO_708 (O_708,N_24990,N_24862);
and UO_709 (O_709,N_24963,N_24759);
and UO_710 (O_710,N_24864,N_24850);
nor UO_711 (O_711,N_24778,N_24965);
xnor UO_712 (O_712,N_24973,N_24821);
or UO_713 (O_713,N_24846,N_24986);
nand UO_714 (O_714,N_24919,N_24831);
and UO_715 (O_715,N_24804,N_24892);
xnor UO_716 (O_716,N_24783,N_24761);
xnor UO_717 (O_717,N_24803,N_24820);
and UO_718 (O_718,N_24993,N_24998);
xnor UO_719 (O_719,N_24961,N_24810);
and UO_720 (O_720,N_24937,N_24840);
or UO_721 (O_721,N_24807,N_24761);
xor UO_722 (O_722,N_24896,N_24948);
and UO_723 (O_723,N_24838,N_24883);
xnor UO_724 (O_724,N_24858,N_24927);
nand UO_725 (O_725,N_24781,N_24799);
xnor UO_726 (O_726,N_24969,N_24817);
nor UO_727 (O_727,N_24813,N_24896);
nor UO_728 (O_728,N_24771,N_24866);
or UO_729 (O_729,N_24854,N_24916);
xor UO_730 (O_730,N_24837,N_24891);
nand UO_731 (O_731,N_24875,N_24815);
nand UO_732 (O_732,N_24852,N_24832);
and UO_733 (O_733,N_24757,N_24936);
xor UO_734 (O_734,N_24796,N_24793);
xnor UO_735 (O_735,N_24956,N_24807);
nand UO_736 (O_736,N_24784,N_24979);
nand UO_737 (O_737,N_24945,N_24867);
nor UO_738 (O_738,N_24849,N_24971);
nand UO_739 (O_739,N_24929,N_24886);
or UO_740 (O_740,N_24788,N_24795);
nand UO_741 (O_741,N_24857,N_24765);
nor UO_742 (O_742,N_24961,N_24773);
nor UO_743 (O_743,N_24993,N_24940);
or UO_744 (O_744,N_24886,N_24806);
xor UO_745 (O_745,N_24996,N_24758);
nor UO_746 (O_746,N_24863,N_24989);
and UO_747 (O_747,N_24752,N_24979);
and UO_748 (O_748,N_24775,N_24953);
nor UO_749 (O_749,N_24903,N_24920);
xnor UO_750 (O_750,N_24875,N_24877);
nor UO_751 (O_751,N_24866,N_24857);
or UO_752 (O_752,N_24885,N_24888);
xor UO_753 (O_753,N_24802,N_24961);
nand UO_754 (O_754,N_24881,N_24767);
nor UO_755 (O_755,N_24774,N_24882);
xnor UO_756 (O_756,N_24768,N_24930);
and UO_757 (O_757,N_24906,N_24878);
and UO_758 (O_758,N_24858,N_24917);
or UO_759 (O_759,N_24779,N_24894);
nor UO_760 (O_760,N_24777,N_24952);
or UO_761 (O_761,N_24898,N_24997);
nor UO_762 (O_762,N_24876,N_24861);
nor UO_763 (O_763,N_24820,N_24971);
nor UO_764 (O_764,N_24785,N_24853);
nor UO_765 (O_765,N_24974,N_24968);
nor UO_766 (O_766,N_24818,N_24813);
nor UO_767 (O_767,N_24963,N_24919);
nor UO_768 (O_768,N_24947,N_24955);
and UO_769 (O_769,N_24872,N_24780);
or UO_770 (O_770,N_24942,N_24893);
xnor UO_771 (O_771,N_24969,N_24775);
xnor UO_772 (O_772,N_24876,N_24796);
nand UO_773 (O_773,N_24842,N_24940);
xor UO_774 (O_774,N_24758,N_24800);
and UO_775 (O_775,N_24917,N_24897);
and UO_776 (O_776,N_24905,N_24877);
nand UO_777 (O_777,N_24760,N_24823);
or UO_778 (O_778,N_24840,N_24887);
nand UO_779 (O_779,N_24998,N_24764);
nand UO_780 (O_780,N_24846,N_24778);
xor UO_781 (O_781,N_24827,N_24758);
nand UO_782 (O_782,N_24755,N_24857);
nor UO_783 (O_783,N_24862,N_24912);
xnor UO_784 (O_784,N_24946,N_24922);
nand UO_785 (O_785,N_24909,N_24988);
nand UO_786 (O_786,N_24940,N_24784);
xor UO_787 (O_787,N_24821,N_24759);
xnor UO_788 (O_788,N_24835,N_24961);
xnor UO_789 (O_789,N_24981,N_24938);
nor UO_790 (O_790,N_24865,N_24982);
nor UO_791 (O_791,N_24758,N_24899);
nor UO_792 (O_792,N_24853,N_24789);
or UO_793 (O_793,N_24889,N_24757);
or UO_794 (O_794,N_24830,N_24900);
or UO_795 (O_795,N_24808,N_24775);
and UO_796 (O_796,N_24886,N_24969);
and UO_797 (O_797,N_24762,N_24975);
and UO_798 (O_798,N_24826,N_24857);
nor UO_799 (O_799,N_24765,N_24944);
xor UO_800 (O_800,N_24847,N_24854);
nand UO_801 (O_801,N_24874,N_24975);
nand UO_802 (O_802,N_24814,N_24912);
and UO_803 (O_803,N_24899,N_24821);
nand UO_804 (O_804,N_24870,N_24806);
nor UO_805 (O_805,N_24961,N_24976);
nor UO_806 (O_806,N_24900,N_24896);
xnor UO_807 (O_807,N_24885,N_24862);
nand UO_808 (O_808,N_24864,N_24972);
and UO_809 (O_809,N_24951,N_24967);
and UO_810 (O_810,N_24797,N_24889);
and UO_811 (O_811,N_24788,N_24824);
xor UO_812 (O_812,N_24781,N_24904);
xor UO_813 (O_813,N_24832,N_24997);
nor UO_814 (O_814,N_24884,N_24770);
nor UO_815 (O_815,N_24861,N_24893);
nor UO_816 (O_816,N_24871,N_24920);
xnor UO_817 (O_817,N_24963,N_24922);
or UO_818 (O_818,N_24771,N_24877);
nor UO_819 (O_819,N_24994,N_24787);
xor UO_820 (O_820,N_24803,N_24792);
and UO_821 (O_821,N_24754,N_24812);
xnor UO_822 (O_822,N_24916,N_24980);
or UO_823 (O_823,N_24972,N_24935);
or UO_824 (O_824,N_24830,N_24901);
nand UO_825 (O_825,N_24798,N_24787);
xnor UO_826 (O_826,N_24916,N_24796);
nor UO_827 (O_827,N_24971,N_24937);
or UO_828 (O_828,N_24837,N_24969);
xnor UO_829 (O_829,N_24847,N_24985);
and UO_830 (O_830,N_24962,N_24866);
and UO_831 (O_831,N_24927,N_24758);
nand UO_832 (O_832,N_24907,N_24957);
and UO_833 (O_833,N_24830,N_24869);
xor UO_834 (O_834,N_24828,N_24829);
nand UO_835 (O_835,N_24986,N_24991);
and UO_836 (O_836,N_24881,N_24886);
nand UO_837 (O_837,N_24860,N_24815);
or UO_838 (O_838,N_24966,N_24753);
nor UO_839 (O_839,N_24991,N_24974);
or UO_840 (O_840,N_24878,N_24934);
xor UO_841 (O_841,N_24939,N_24948);
nand UO_842 (O_842,N_24990,N_24834);
nand UO_843 (O_843,N_24933,N_24905);
and UO_844 (O_844,N_24942,N_24838);
nand UO_845 (O_845,N_24777,N_24995);
or UO_846 (O_846,N_24757,N_24806);
and UO_847 (O_847,N_24814,N_24966);
and UO_848 (O_848,N_24846,N_24833);
nand UO_849 (O_849,N_24792,N_24785);
and UO_850 (O_850,N_24816,N_24900);
xor UO_851 (O_851,N_24885,N_24874);
xor UO_852 (O_852,N_24898,N_24905);
or UO_853 (O_853,N_24934,N_24912);
or UO_854 (O_854,N_24820,N_24980);
xnor UO_855 (O_855,N_24996,N_24985);
xnor UO_856 (O_856,N_24995,N_24950);
nand UO_857 (O_857,N_24776,N_24920);
nor UO_858 (O_858,N_24954,N_24783);
xnor UO_859 (O_859,N_24809,N_24773);
xnor UO_860 (O_860,N_24805,N_24893);
or UO_861 (O_861,N_24837,N_24908);
nor UO_862 (O_862,N_24840,N_24950);
xor UO_863 (O_863,N_24875,N_24851);
nor UO_864 (O_864,N_24858,N_24808);
or UO_865 (O_865,N_24761,N_24779);
or UO_866 (O_866,N_24871,N_24761);
nand UO_867 (O_867,N_24955,N_24795);
nand UO_868 (O_868,N_24930,N_24816);
and UO_869 (O_869,N_24826,N_24941);
nand UO_870 (O_870,N_24895,N_24795);
xor UO_871 (O_871,N_24876,N_24920);
xor UO_872 (O_872,N_24766,N_24982);
nand UO_873 (O_873,N_24832,N_24753);
nand UO_874 (O_874,N_24994,N_24949);
and UO_875 (O_875,N_24869,N_24812);
nand UO_876 (O_876,N_24794,N_24776);
xor UO_877 (O_877,N_24960,N_24973);
nor UO_878 (O_878,N_24938,N_24844);
nor UO_879 (O_879,N_24994,N_24758);
and UO_880 (O_880,N_24788,N_24829);
or UO_881 (O_881,N_24949,N_24918);
xor UO_882 (O_882,N_24953,N_24910);
nor UO_883 (O_883,N_24750,N_24996);
or UO_884 (O_884,N_24878,N_24872);
nand UO_885 (O_885,N_24822,N_24815);
xor UO_886 (O_886,N_24872,N_24979);
or UO_887 (O_887,N_24852,N_24892);
or UO_888 (O_888,N_24785,N_24886);
nand UO_889 (O_889,N_24944,N_24785);
nor UO_890 (O_890,N_24971,N_24805);
nand UO_891 (O_891,N_24899,N_24765);
xnor UO_892 (O_892,N_24817,N_24811);
nand UO_893 (O_893,N_24998,N_24873);
and UO_894 (O_894,N_24880,N_24869);
nor UO_895 (O_895,N_24757,N_24986);
and UO_896 (O_896,N_24872,N_24977);
nor UO_897 (O_897,N_24784,N_24980);
xor UO_898 (O_898,N_24770,N_24796);
and UO_899 (O_899,N_24967,N_24826);
xnor UO_900 (O_900,N_24959,N_24975);
nand UO_901 (O_901,N_24942,N_24906);
or UO_902 (O_902,N_24788,N_24760);
xnor UO_903 (O_903,N_24897,N_24958);
nor UO_904 (O_904,N_24783,N_24754);
or UO_905 (O_905,N_24940,N_24758);
nor UO_906 (O_906,N_24917,N_24765);
or UO_907 (O_907,N_24776,N_24770);
nor UO_908 (O_908,N_24929,N_24884);
and UO_909 (O_909,N_24766,N_24855);
nand UO_910 (O_910,N_24783,N_24901);
nand UO_911 (O_911,N_24804,N_24938);
xor UO_912 (O_912,N_24909,N_24754);
nand UO_913 (O_913,N_24948,N_24928);
or UO_914 (O_914,N_24829,N_24979);
and UO_915 (O_915,N_24823,N_24845);
nand UO_916 (O_916,N_24962,N_24991);
nand UO_917 (O_917,N_24841,N_24938);
and UO_918 (O_918,N_24931,N_24900);
or UO_919 (O_919,N_24860,N_24766);
nor UO_920 (O_920,N_24945,N_24916);
and UO_921 (O_921,N_24770,N_24927);
or UO_922 (O_922,N_24813,N_24874);
nor UO_923 (O_923,N_24851,N_24870);
nor UO_924 (O_924,N_24988,N_24757);
nor UO_925 (O_925,N_24786,N_24982);
and UO_926 (O_926,N_24900,N_24942);
or UO_927 (O_927,N_24758,N_24820);
nand UO_928 (O_928,N_24757,N_24879);
nor UO_929 (O_929,N_24807,N_24963);
or UO_930 (O_930,N_24901,N_24820);
or UO_931 (O_931,N_24823,N_24822);
nor UO_932 (O_932,N_24806,N_24990);
or UO_933 (O_933,N_24784,N_24964);
nor UO_934 (O_934,N_24910,N_24814);
nand UO_935 (O_935,N_24863,N_24798);
nand UO_936 (O_936,N_24948,N_24886);
nand UO_937 (O_937,N_24817,N_24971);
nand UO_938 (O_938,N_24821,N_24966);
nand UO_939 (O_939,N_24973,N_24899);
nor UO_940 (O_940,N_24927,N_24948);
nand UO_941 (O_941,N_24949,N_24830);
or UO_942 (O_942,N_24850,N_24994);
nor UO_943 (O_943,N_24824,N_24937);
and UO_944 (O_944,N_24816,N_24844);
and UO_945 (O_945,N_24888,N_24906);
and UO_946 (O_946,N_24956,N_24875);
xor UO_947 (O_947,N_24916,N_24965);
or UO_948 (O_948,N_24921,N_24880);
nand UO_949 (O_949,N_24814,N_24840);
or UO_950 (O_950,N_24917,N_24928);
nand UO_951 (O_951,N_24861,N_24997);
nor UO_952 (O_952,N_24991,N_24945);
and UO_953 (O_953,N_24928,N_24916);
or UO_954 (O_954,N_24773,N_24967);
and UO_955 (O_955,N_24829,N_24780);
or UO_956 (O_956,N_24992,N_24976);
or UO_957 (O_957,N_24878,N_24822);
nand UO_958 (O_958,N_24866,N_24769);
nand UO_959 (O_959,N_24888,N_24847);
or UO_960 (O_960,N_24983,N_24892);
or UO_961 (O_961,N_24875,N_24840);
xor UO_962 (O_962,N_24888,N_24918);
nand UO_963 (O_963,N_24832,N_24831);
xnor UO_964 (O_964,N_24752,N_24832);
nor UO_965 (O_965,N_24802,N_24893);
xnor UO_966 (O_966,N_24831,N_24813);
nor UO_967 (O_967,N_24990,N_24943);
xnor UO_968 (O_968,N_24790,N_24793);
and UO_969 (O_969,N_24854,N_24796);
nand UO_970 (O_970,N_24992,N_24873);
or UO_971 (O_971,N_24900,N_24894);
xor UO_972 (O_972,N_24939,N_24776);
or UO_973 (O_973,N_24837,N_24961);
nor UO_974 (O_974,N_24983,N_24842);
nand UO_975 (O_975,N_24880,N_24792);
nand UO_976 (O_976,N_24937,N_24781);
or UO_977 (O_977,N_24845,N_24929);
or UO_978 (O_978,N_24946,N_24813);
and UO_979 (O_979,N_24849,N_24817);
or UO_980 (O_980,N_24900,N_24828);
and UO_981 (O_981,N_24852,N_24993);
and UO_982 (O_982,N_24894,N_24917);
or UO_983 (O_983,N_24876,N_24977);
xor UO_984 (O_984,N_24973,N_24930);
or UO_985 (O_985,N_24790,N_24789);
nor UO_986 (O_986,N_24885,N_24866);
and UO_987 (O_987,N_24835,N_24831);
and UO_988 (O_988,N_24848,N_24847);
and UO_989 (O_989,N_24996,N_24930);
nor UO_990 (O_990,N_24983,N_24999);
nor UO_991 (O_991,N_24760,N_24810);
nand UO_992 (O_992,N_24816,N_24935);
or UO_993 (O_993,N_24840,N_24804);
nand UO_994 (O_994,N_24958,N_24992);
nand UO_995 (O_995,N_24757,N_24864);
nor UO_996 (O_996,N_24911,N_24929);
and UO_997 (O_997,N_24980,N_24894);
xnor UO_998 (O_998,N_24775,N_24852);
or UO_999 (O_999,N_24809,N_24759);
nand UO_1000 (O_1000,N_24759,N_24766);
or UO_1001 (O_1001,N_24916,N_24885);
or UO_1002 (O_1002,N_24998,N_24798);
and UO_1003 (O_1003,N_24888,N_24921);
or UO_1004 (O_1004,N_24792,N_24821);
nand UO_1005 (O_1005,N_24965,N_24830);
or UO_1006 (O_1006,N_24978,N_24783);
or UO_1007 (O_1007,N_24778,N_24963);
and UO_1008 (O_1008,N_24839,N_24857);
or UO_1009 (O_1009,N_24997,N_24760);
nand UO_1010 (O_1010,N_24920,N_24796);
nand UO_1011 (O_1011,N_24817,N_24846);
and UO_1012 (O_1012,N_24819,N_24909);
nor UO_1013 (O_1013,N_24943,N_24812);
nor UO_1014 (O_1014,N_24941,N_24859);
and UO_1015 (O_1015,N_24824,N_24994);
or UO_1016 (O_1016,N_24775,N_24992);
and UO_1017 (O_1017,N_24913,N_24860);
or UO_1018 (O_1018,N_24990,N_24824);
nand UO_1019 (O_1019,N_24755,N_24805);
nand UO_1020 (O_1020,N_24821,N_24985);
and UO_1021 (O_1021,N_24886,N_24826);
nand UO_1022 (O_1022,N_24950,N_24918);
xor UO_1023 (O_1023,N_24884,N_24845);
xor UO_1024 (O_1024,N_24825,N_24986);
nand UO_1025 (O_1025,N_24948,N_24953);
nor UO_1026 (O_1026,N_24877,N_24799);
and UO_1027 (O_1027,N_24872,N_24981);
nor UO_1028 (O_1028,N_24994,N_24760);
nor UO_1029 (O_1029,N_24920,N_24954);
nor UO_1030 (O_1030,N_24885,N_24812);
nand UO_1031 (O_1031,N_24777,N_24861);
nor UO_1032 (O_1032,N_24838,N_24957);
nor UO_1033 (O_1033,N_24797,N_24987);
xor UO_1034 (O_1034,N_24871,N_24841);
or UO_1035 (O_1035,N_24844,N_24972);
or UO_1036 (O_1036,N_24978,N_24770);
nor UO_1037 (O_1037,N_24933,N_24960);
and UO_1038 (O_1038,N_24883,N_24882);
nor UO_1039 (O_1039,N_24814,N_24802);
or UO_1040 (O_1040,N_24919,N_24855);
nand UO_1041 (O_1041,N_24966,N_24936);
or UO_1042 (O_1042,N_24795,N_24951);
xor UO_1043 (O_1043,N_24964,N_24896);
nor UO_1044 (O_1044,N_24790,N_24896);
xor UO_1045 (O_1045,N_24771,N_24913);
and UO_1046 (O_1046,N_24958,N_24975);
nand UO_1047 (O_1047,N_24805,N_24919);
nor UO_1048 (O_1048,N_24915,N_24978);
xnor UO_1049 (O_1049,N_24830,N_24753);
xor UO_1050 (O_1050,N_24802,N_24992);
xnor UO_1051 (O_1051,N_24994,N_24904);
xor UO_1052 (O_1052,N_24903,N_24901);
nand UO_1053 (O_1053,N_24837,N_24787);
xor UO_1054 (O_1054,N_24965,N_24946);
nand UO_1055 (O_1055,N_24901,N_24933);
or UO_1056 (O_1056,N_24836,N_24769);
nand UO_1057 (O_1057,N_24983,N_24938);
and UO_1058 (O_1058,N_24758,N_24841);
or UO_1059 (O_1059,N_24757,N_24801);
nand UO_1060 (O_1060,N_24816,N_24834);
nor UO_1061 (O_1061,N_24849,N_24990);
nand UO_1062 (O_1062,N_24973,N_24879);
xor UO_1063 (O_1063,N_24825,N_24974);
or UO_1064 (O_1064,N_24782,N_24810);
nand UO_1065 (O_1065,N_24970,N_24801);
or UO_1066 (O_1066,N_24870,N_24771);
nand UO_1067 (O_1067,N_24856,N_24779);
xnor UO_1068 (O_1068,N_24933,N_24817);
and UO_1069 (O_1069,N_24785,N_24888);
xor UO_1070 (O_1070,N_24810,N_24867);
or UO_1071 (O_1071,N_24999,N_24856);
or UO_1072 (O_1072,N_24876,N_24945);
xnor UO_1073 (O_1073,N_24895,N_24993);
and UO_1074 (O_1074,N_24762,N_24818);
xor UO_1075 (O_1075,N_24769,N_24768);
xor UO_1076 (O_1076,N_24817,N_24929);
nand UO_1077 (O_1077,N_24907,N_24958);
nor UO_1078 (O_1078,N_24996,N_24757);
nor UO_1079 (O_1079,N_24793,N_24865);
nor UO_1080 (O_1080,N_24940,N_24858);
xor UO_1081 (O_1081,N_24945,N_24861);
and UO_1082 (O_1082,N_24922,N_24799);
nand UO_1083 (O_1083,N_24956,N_24968);
and UO_1084 (O_1084,N_24785,N_24914);
or UO_1085 (O_1085,N_24924,N_24782);
nor UO_1086 (O_1086,N_24814,N_24875);
nand UO_1087 (O_1087,N_24910,N_24864);
xor UO_1088 (O_1088,N_24993,N_24879);
xnor UO_1089 (O_1089,N_24796,N_24936);
nor UO_1090 (O_1090,N_24834,N_24996);
nor UO_1091 (O_1091,N_24986,N_24885);
xnor UO_1092 (O_1092,N_24881,N_24760);
or UO_1093 (O_1093,N_24783,N_24973);
nor UO_1094 (O_1094,N_24882,N_24800);
nand UO_1095 (O_1095,N_24762,N_24910);
xor UO_1096 (O_1096,N_24825,N_24766);
or UO_1097 (O_1097,N_24757,N_24759);
xor UO_1098 (O_1098,N_24782,N_24917);
nand UO_1099 (O_1099,N_24826,N_24986);
nor UO_1100 (O_1100,N_24774,N_24850);
or UO_1101 (O_1101,N_24834,N_24772);
and UO_1102 (O_1102,N_24829,N_24834);
nor UO_1103 (O_1103,N_24907,N_24936);
nand UO_1104 (O_1104,N_24957,N_24976);
and UO_1105 (O_1105,N_24876,N_24994);
nor UO_1106 (O_1106,N_24896,N_24967);
or UO_1107 (O_1107,N_24999,N_24939);
nand UO_1108 (O_1108,N_24765,N_24844);
nand UO_1109 (O_1109,N_24825,N_24983);
or UO_1110 (O_1110,N_24862,N_24951);
and UO_1111 (O_1111,N_24806,N_24917);
nor UO_1112 (O_1112,N_24786,N_24945);
xnor UO_1113 (O_1113,N_24979,N_24990);
xnor UO_1114 (O_1114,N_24795,N_24937);
and UO_1115 (O_1115,N_24802,N_24895);
and UO_1116 (O_1116,N_24998,N_24825);
nand UO_1117 (O_1117,N_24804,N_24836);
xnor UO_1118 (O_1118,N_24831,N_24800);
or UO_1119 (O_1119,N_24822,N_24899);
and UO_1120 (O_1120,N_24940,N_24818);
and UO_1121 (O_1121,N_24958,N_24834);
xnor UO_1122 (O_1122,N_24796,N_24957);
xnor UO_1123 (O_1123,N_24872,N_24881);
and UO_1124 (O_1124,N_24857,N_24973);
nand UO_1125 (O_1125,N_24917,N_24792);
and UO_1126 (O_1126,N_24916,N_24969);
or UO_1127 (O_1127,N_24884,N_24951);
or UO_1128 (O_1128,N_24946,N_24854);
and UO_1129 (O_1129,N_24976,N_24763);
nor UO_1130 (O_1130,N_24900,N_24754);
nor UO_1131 (O_1131,N_24990,N_24799);
nor UO_1132 (O_1132,N_24938,N_24862);
nor UO_1133 (O_1133,N_24878,N_24768);
nand UO_1134 (O_1134,N_24915,N_24928);
and UO_1135 (O_1135,N_24984,N_24924);
and UO_1136 (O_1136,N_24773,N_24799);
nor UO_1137 (O_1137,N_24928,N_24956);
xnor UO_1138 (O_1138,N_24987,N_24982);
and UO_1139 (O_1139,N_24999,N_24786);
nand UO_1140 (O_1140,N_24873,N_24870);
nand UO_1141 (O_1141,N_24822,N_24832);
or UO_1142 (O_1142,N_24923,N_24762);
or UO_1143 (O_1143,N_24961,N_24913);
nand UO_1144 (O_1144,N_24852,N_24752);
or UO_1145 (O_1145,N_24837,N_24916);
or UO_1146 (O_1146,N_24973,N_24902);
and UO_1147 (O_1147,N_24955,N_24872);
and UO_1148 (O_1148,N_24970,N_24938);
nand UO_1149 (O_1149,N_24762,N_24981);
and UO_1150 (O_1150,N_24994,N_24980);
nor UO_1151 (O_1151,N_24965,N_24801);
nor UO_1152 (O_1152,N_24878,N_24844);
or UO_1153 (O_1153,N_24834,N_24823);
or UO_1154 (O_1154,N_24768,N_24794);
or UO_1155 (O_1155,N_24956,N_24992);
or UO_1156 (O_1156,N_24761,N_24796);
nor UO_1157 (O_1157,N_24880,N_24839);
and UO_1158 (O_1158,N_24917,N_24758);
and UO_1159 (O_1159,N_24770,N_24872);
and UO_1160 (O_1160,N_24778,N_24955);
and UO_1161 (O_1161,N_24936,N_24915);
xnor UO_1162 (O_1162,N_24781,N_24980);
nand UO_1163 (O_1163,N_24936,N_24949);
nand UO_1164 (O_1164,N_24777,N_24915);
nor UO_1165 (O_1165,N_24773,N_24938);
nand UO_1166 (O_1166,N_24978,N_24834);
or UO_1167 (O_1167,N_24888,N_24955);
xnor UO_1168 (O_1168,N_24864,N_24775);
or UO_1169 (O_1169,N_24988,N_24773);
nor UO_1170 (O_1170,N_24893,N_24824);
and UO_1171 (O_1171,N_24908,N_24943);
nor UO_1172 (O_1172,N_24904,N_24890);
nor UO_1173 (O_1173,N_24986,N_24968);
and UO_1174 (O_1174,N_24924,N_24998);
xnor UO_1175 (O_1175,N_24919,N_24911);
nor UO_1176 (O_1176,N_24967,N_24926);
and UO_1177 (O_1177,N_24791,N_24861);
nor UO_1178 (O_1178,N_24986,N_24907);
xnor UO_1179 (O_1179,N_24848,N_24829);
xor UO_1180 (O_1180,N_24995,N_24828);
xnor UO_1181 (O_1181,N_24905,N_24867);
and UO_1182 (O_1182,N_24879,N_24803);
xor UO_1183 (O_1183,N_24950,N_24793);
nor UO_1184 (O_1184,N_24939,N_24826);
and UO_1185 (O_1185,N_24794,N_24752);
nor UO_1186 (O_1186,N_24825,N_24879);
or UO_1187 (O_1187,N_24796,N_24880);
or UO_1188 (O_1188,N_24938,N_24847);
xor UO_1189 (O_1189,N_24799,N_24805);
or UO_1190 (O_1190,N_24811,N_24882);
nor UO_1191 (O_1191,N_24913,N_24937);
nor UO_1192 (O_1192,N_24841,N_24995);
or UO_1193 (O_1193,N_24825,N_24896);
nand UO_1194 (O_1194,N_24895,N_24834);
nand UO_1195 (O_1195,N_24884,N_24994);
or UO_1196 (O_1196,N_24874,N_24823);
xor UO_1197 (O_1197,N_24962,N_24776);
or UO_1198 (O_1198,N_24842,N_24820);
xnor UO_1199 (O_1199,N_24879,N_24785);
nand UO_1200 (O_1200,N_24773,N_24968);
nand UO_1201 (O_1201,N_24864,N_24947);
or UO_1202 (O_1202,N_24861,N_24803);
xor UO_1203 (O_1203,N_24919,N_24870);
nor UO_1204 (O_1204,N_24906,N_24907);
and UO_1205 (O_1205,N_24757,N_24952);
xor UO_1206 (O_1206,N_24958,N_24961);
xor UO_1207 (O_1207,N_24899,N_24796);
nand UO_1208 (O_1208,N_24963,N_24793);
xor UO_1209 (O_1209,N_24994,N_24831);
xnor UO_1210 (O_1210,N_24862,N_24778);
or UO_1211 (O_1211,N_24909,N_24968);
or UO_1212 (O_1212,N_24990,N_24957);
xor UO_1213 (O_1213,N_24929,N_24819);
or UO_1214 (O_1214,N_24956,N_24840);
and UO_1215 (O_1215,N_24911,N_24780);
xor UO_1216 (O_1216,N_24974,N_24863);
nor UO_1217 (O_1217,N_24816,N_24807);
nor UO_1218 (O_1218,N_24953,N_24913);
or UO_1219 (O_1219,N_24847,N_24967);
or UO_1220 (O_1220,N_24756,N_24997);
or UO_1221 (O_1221,N_24843,N_24897);
nor UO_1222 (O_1222,N_24785,N_24834);
and UO_1223 (O_1223,N_24992,N_24779);
or UO_1224 (O_1224,N_24782,N_24795);
xor UO_1225 (O_1225,N_24935,N_24849);
nand UO_1226 (O_1226,N_24773,N_24786);
nand UO_1227 (O_1227,N_24903,N_24854);
nand UO_1228 (O_1228,N_24782,N_24817);
or UO_1229 (O_1229,N_24851,N_24776);
nand UO_1230 (O_1230,N_24755,N_24906);
nand UO_1231 (O_1231,N_24924,N_24963);
nor UO_1232 (O_1232,N_24990,N_24908);
nor UO_1233 (O_1233,N_24762,N_24992);
and UO_1234 (O_1234,N_24840,N_24970);
and UO_1235 (O_1235,N_24861,N_24914);
nor UO_1236 (O_1236,N_24752,N_24806);
nor UO_1237 (O_1237,N_24840,N_24790);
nor UO_1238 (O_1238,N_24855,N_24842);
and UO_1239 (O_1239,N_24896,N_24861);
nand UO_1240 (O_1240,N_24901,N_24996);
xnor UO_1241 (O_1241,N_24962,N_24955);
xor UO_1242 (O_1242,N_24984,N_24967);
or UO_1243 (O_1243,N_24827,N_24879);
or UO_1244 (O_1244,N_24769,N_24790);
nor UO_1245 (O_1245,N_24847,N_24809);
and UO_1246 (O_1246,N_24791,N_24890);
or UO_1247 (O_1247,N_24876,N_24840);
or UO_1248 (O_1248,N_24906,N_24809);
nor UO_1249 (O_1249,N_24941,N_24905);
nand UO_1250 (O_1250,N_24769,N_24860);
or UO_1251 (O_1251,N_24764,N_24993);
or UO_1252 (O_1252,N_24954,N_24851);
and UO_1253 (O_1253,N_24783,N_24834);
xor UO_1254 (O_1254,N_24956,N_24797);
xor UO_1255 (O_1255,N_24769,N_24950);
or UO_1256 (O_1256,N_24840,N_24803);
and UO_1257 (O_1257,N_24884,N_24995);
nand UO_1258 (O_1258,N_24838,N_24827);
nand UO_1259 (O_1259,N_24846,N_24813);
nor UO_1260 (O_1260,N_24800,N_24994);
or UO_1261 (O_1261,N_24778,N_24865);
or UO_1262 (O_1262,N_24889,N_24940);
nand UO_1263 (O_1263,N_24771,N_24780);
and UO_1264 (O_1264,N_24788,N_24791);
or UO_1265 (O_1265,N_24811,N_24866);
or UO_1266 (O_1266,N_24874,N_24758);
nand UO_1267 (O_1267,N_24843,N_24858);
and UO_1268 (O_1268,N_24836,N_24822);
nor UO_1269 (O_1269,N_24830,N_24994);
nor UO_1270 (O_1270,N_24961,N_24808);
or UO_1271 (O_1271,N_24768,N_24950);
or UO_1272 (O_1272,N_24884,N_24865);
nor UO_1273 (O_1273,N_24847,N_24753);
nand UO_1274 (O_1274,N_24952,N_24948);
nand UO_1275 (O_1275,N_24926,N_24818);
xor UO_1276 (O_1276,N_24934,N_24940);
nand UO_1277 (O_1277,N_24774,N_24925);
xor UO_1278 (O_1278,N_24998,N_24835);
xor UO_1279 (O_1279,N_24979,N_24793);
and UO_1280 (O_1280,N_24808,N_24846);
or UO_1281 (O_1281,N_24891,N_24976);
nor UO_1282 (O_1282,N_24944,N_24982);
or UO_1283 (O_1283,N_24941,N_24780);
and UO_1284 (O_1284,N_24776,N_24855);
and UO_1285 (O_1285,N_24992,N_24909);
xnor UO_1286 (O_1286,N_24936,N_24782);
and UO_1287 (O_1287,N_24837,N_24985);
nand UO_1288 (O_1288,N_24952,N_24800);
nor UO_1289 (O_1289,N_24946,N_24935);
nor UO_1290 (O_1290,N_24881,N_24975);
and UO_1291 (O_1291,N_24988,N_24883);
nand UO_1292 (O_1292,N_24847,N_24952);
nand UO_1293 (O_1293,N_24887,N_24784);
or UO_1294 (O_1294,N_24917,N_24960);
xor UO_1295 (O_1295,N_24893,N_24867);
nand UO_1296 (O_1296,N_24839,N_24958);
xnor UO_1297 (O_1297,N_24752,N_24805);
nor UO_1298 (O_1298,N_24934,N_24855);
and UO_1299 (O_1299,N_24875,N_24921);
and UO_1300 (O_1300,N_24887,N_24760);
nand UO_1301 (O_1301,N_24977,N_24908);
nor UO_1302 (O_1302,N_24871,N_24759);
xnor UO_1303 (O_1303,N_24883,N_24826);
xor UO_1304 (O_1304,N_24898,N_24921);
nand UO_1305 (O_1305,N_24806,N_24790);
and UO_1306 (O_1306,N_24865,N_24844);
nor UO_1307 (O_1307,N_24956,N_24977);
xnor UO_1308 (O_1308,N_24877,N_24761);
and UO_1309 (O_1309,N_24826,N_24960);
xnor UO_1310 (O_1310,N_24876,N_24962);
nand UO_1311 (O_1311,N_24930,N_24979);
nand UO_1312 (O_1312,N_24756,N_24967);
nand UO_1313 (O_1313,N_24910,N_24854);
and UO_1314 (O_1314,N_24810,N_24870);
nand UO_1315 (O_1315,N_24751,N_24886);
or UO_1316 (O_1316,N_24966,N_24826);
or UO_1317 (O_1317,N_24972,N_24841);
nand UO_1318 (O_1318,N_24969,N_24757);
nor UO_1319 (O_1319,N_24851,N_24992);
and UO_1320 (O_1320,N_24788,N_24854);
nor UO_1321 (O_1321,N_24949,N_24953);
and UO_1322 (O_1322,N_24868,N_24970);
or UO_1323 (O_1323,N_24783,N_24945);
or UO_1324 (O_1324,N_24855,N_24957);
nor UO_1325 (O_1325,N_24784,N_24999);
xnor UO_1326 (O_1326,N_24783,N_24776);
nand UO_1327 (O_1327,N_24862,N_24871);
and UO_1328 (O_1328,N_24850,N_24924);
nand UO_1329 (O_1329,N_24895,N_24805);
xnor UO_1330 (O_1330,N_24849,N_24885);
and UO_1331 (O_1331,N_24798,N_24780);
or UO_1332 (O_1332,N_24788,N_24994);
and UO_1333 (O_1333,N_24806,N_24968);
and UO_1334 (O_1334,N_24906,N_24820);
nor UO_1335 (O_1335,N_24945,N_24780);
xnor UO_1336 (O_1336,N_24752,N_24818);
or UO_1337 (O_1337,N_24906,N_24851);
nor UO_1338 (O_1338,N_24928,N_24750);
or UO_1339 (O_1339,N_24948,N_24758);
nand UO_1340 (O_1340,N_24848,N_24765);
nand UO_1341 (O_1341,N_24898,N_24803);
nand UO_1342 (O_1342,N_24806,N_24777);
nor UO_1343 (O_1343,N_24819,N_24861);
xor UO_1344 (O_1344,N_24802,N_24905);
nand UO_1345 (O_1345,N_24872,N_24755);
or UO_1346 (O_1346,N_24769,N_24933);
or UO_1347 (O_1347,N_24781,N_24901);
or UO_1348 (O_1348,N_24895,N_24840);
and UO_1349 (O_1349,N_24869,N_24762);
xor UO_1350 (O_1350,N_24834,N_24999);
or UO_1351 (O_1351,N_24802,N_24773);
xor UO_1352 (O_1352,N_24896,N_24809);
xnor UO_1353 (O_1353,N_24931,N_24858);
or UO_1354 (O_1354,N_24781,N_24792);
xnor UO_1355 (O_1355,N_24892,N_24813);
nor UO_1356 (O_1356,N_24920,N_24774);
and UO_1357 (O_1357,N_24963,N_24752);
and UO_1358 (O_1358,N_24973,N_24848);
or UO_1359 (O_1359,N_24758,N_24961);
nor UO_1360 (O_1360,N_24868,N_24893);
and UO_1361 (O_1361,N_24796,N_24883);
and UO_1362 (O_1362,N_24864,N_24828);
xnor UO_1363 (O_1363,N_24881,N_24852);
and UO_1364 (O_1364,N_24922,N_24950);
nand UO_1365 (O_1365,N_24907,N_24750);
xor UO_1366 (O_1366,N_24899,N_24966);
nor UO_1367 (O_1367,N_24782,N_24809);
or UO_1368 (O_1368,N_24806,N_24763);
nand UO_1369 (O_1369,N_24875,N_24821);
and UO_1370 (O_1370,N_24894,N_24775);
or UO_1371 (O_1371,N_24952,N_24988);
nor UO_1372 (O_1372,N_24895,N_24921);
nand UO_1373 (O_1373,N_24945,N_24829);
nand UO_1374 (O_1374,N_24759,N_24927);
xor UO_1375 (O_1375,N_24894,N_24817);
or UO_1376 (O_1376,N_24896,N_24832);
nand UO_1377 (O_1377,N_24960,N_24844);
or UO_1378 (O_1378,N_24790,N_24768);
xor UO_1379 (O_1379,N_24937,N_24940);
nand UO_1380 (O_1380,N_24920,N_24962);
and UO_1381 (O_1381,N_24806,N_24992);
and UO_1382 (O_1382,N_24868,N_24866);
nand UO_1383 (O_1383,N_24780,N_24762);
nand UO_1384 (O_1384,N_24931,N_24764);
and UO_1385 (O_1385,N_24790,N_24864);
nand UO_1386 (O_1386,N_24909,N_24850);
nand UO_1387 (O_1387,N_24974,N_24817);
nand UO_1388 (O_1388,N_24987,N_24902);
nand UO_1389 (O_1389,N_24917,N_24956);
or UO_1390 (O_1390,N_24851,N_24924);
nand UO_1391 (O_1391,N_24977,N_24834);
or UO_1392 (O_1392,N_24872,N_24772);
or UO_1393 (O_1393,N_24965,N_24975);
nand UO_1394 (O_1394,N_24787,N_24782);
or UO_1395 (O_1395,N_24975,N_24933);
xnor UO_1396 (O_1396,N_24962,N_24872);
or UO_1397 (O_1397,N_24831,N_24912);
nor UO_1398 (O_1398,N_24911,N_24894);
nor UO_1399 (O_1399,N_24789,N_24986);
xor UO_1400 (O_1400,N_24754,N_24800);
nand UO_1401 (O_1401,N_24798,N_24938);
nand UO_1402 (O_1402,N_24785,N_24814);
and UO_1403 (O_1403,N_24881,N_24966);
or UO_1404 (O_1404,N_24872,N_24987);
or UO_1405 (O_1405,N_24797,N_24829);
and UO_1406 (O_1406,N_24893,N_24947);
nand UO_1407 (O_1407,N_24909,N_24832);
and UO_1408 (O_1408,N_24959,N_24869);
or UO_1409 (O_1409,N_24918,N_24809);
nand UO_1410 (O_1410,N_24865,N_24840);
nand UO_1411 (O_1411,N_24976,N_24885);
nor UO_1412 (O_1412,N_24751,N_24997);
and UO_1413 (O_1413,N_24872,N_24752);
xnor UO_1414 (O_1414,N_24792,N_24982);
or UO_1415 (O_1415,N_24803,N_24917);
nor UO_1416 (O_1416,N_24922,N_24902);
xor UO_1417 (O_1417,N_24808,N_24912);
nor UO_1418 (O_1418,N_24869,N_24751);
or UO_1419 (O_1419,N_24957,N_24763);
and UO_1420 (O_1420,N_24849,N_24938);
nor UO_1421 (O_1421,N_24797,N_24979);
or UO_1422 (O_1422,N_24988,N_24903);
nand UO_1423 (O_1423,N_24920,N_24990);
or UO_1424 (O_1424,N_24832,N_24994);
nand UO_1425 (O_1425,N_24837,N_24834);
or UO_1426 (O_1426,N_24996,N_24923);
nor UO_1427 (O_1427,N_24779,N_24875);
nand UO_1428 (O_1428,N_24862,N_24918);
or UO_1429 (O_1429,N_24953,N_24966);
and UO_1430 (O_1430,N_24863,N_24846);
and UO_1431 (O_1431,N_24843,N_24814);
nand UO_1432 (O_1432,N_24796,N_24879);
nand UO_1433 (O_1433,N_24762,N_24890);
nor UO_1434 (O_1434,N_24954,N_24893);
or UO_1435 (O_1435,N_24916,N_24778);
or UO_1436 (O_1436,N_24872,N_24934);
and UO_1437 (O_1437,N_24988,N_24993);
nor UO_1438 (O_1438,N_24871,N_24894);
or UO_1439 (O_1439,N_24774,N_24895);
nor UO_1440 (O_1440,N_24888,N_24866);
or UO_1441 (O_1441,N_24950,N_24949);
nand UO_1442 (O_1442,N_24880,N_24992);
nor UO_1443 (O_1443,N_24925,N_24910);
nand UO_1444 (O_1444,N_24879,N_24957);
nor UO_1445 (O_1445,N_24817,N_24836);
nand UO_1446 (O_1446,N_24861,N_24853);
and UO_1447 (O_1447,N_24934,N_24826);
or UO_1448 (O_1448,N_24924,N_24835);
nand UO_1449 (O_1449,N_24824,N_24848);
xor UO_1450 (O_1450,N_24935,N_24783);
or UO_1451 (O_1451,N_24754,N_24780);
and UO_1452 (O_1452,N_24888,N_24831);
nand UO_1453 (O_1453,N_24857,N_24879);
or UO_1454 (O_1454,N_24920,N_24767);
or UO_1455 (O_1455,N_24770,N_24809);
or UO_1456 (O_1456,N_24853,N_24984);
or UO_1457 (O_1457,N_24995,N_24818);
nand UO_1458 (O_1458,N_24880,N_24752);
nor UO_1459 (O_1459,N_24840,N_24993);
nor UO_1460 (O_1460,N_24901,N_24790);
nand UO_1461 (O_1461,N_24970,N_24903);
nor UO_1462 (O_1462,N_24825,N_24866);
xor UO_1463 (O_1463,N_24818,N_24805);
or UO_1464 (O_1464,N_24992,N_24817);
xor UO_1465 (O_1465,N_24766,N_24763);
or UO_1466 (O_1466,N_24790,N_24870);
nand UO_1467 (O_1467,N_24911,N_24835);
nand UO_1468 (O_1468,N_24858,N_24855);
nor UO_1469 (O_1469,N_24919,N_24980);
nor UO_1470 (O_1470,N_24957,N_24995);
or UO_1471 (O_1471,N_24957,N_24865);
xnor UO_1472 (O_1472,N_24966,N_24750);
or UO_1473 (O_1473,N_24765,N_24988);
nor UO_1474 (O_1474,N_24950,N_24772);
nor UO_1475 (O_1475,N_24826,N_24772);
nand UO_1476 (O_1476,N_24988,N_24874);
or UO_1477 (O_1477,N_24951,N_24790);
nand UO_1478 (O_1478,N_24845,N_24843);
xor UO_1479 (O_1479,N_24835,N_24761);
xor UO_1480 (O_1480,N_24884,N_24769);
nor UO_1481 (O_1481,N_24945,N_24811);
nand UO_1482 (O_1482,N_24935,N_24755);
or UO_1483 (O_1483,N_24751,N_24998);
or UO_1484 (O_1484,N_24755,N_24813);
or UO_1485 (O_1485,N_24974,N_24791);
nor UO_1486 (O_1486,N_24919,N_24935);
nor UO_1487 (O_1487,N_24787,N_24846);
or UO_1488 (O_1488,N_24853,N_24788);
and UO_1489 (O_1489,N_24840,N_24986);
nand UO_1490 (O_1490,N_24773,N_24980);
nand UO_1491 (O_1491,N_24807,N_24902);
and UO_1492 (O_1492,N_24963,N_24881);
or UO_1493 (O_1493,N_24893,N_24930);
and UO_1494 (O_1494,N_24896,N_24869);
or UO_1495 (O_1495,N_24829,N_24955);
and UO_1496 (O_1496,N_24783,N_24807);
nand UO_1497 (O_1497,N_24995,N_24821);
and UO_1498 (O_1498,N_24817,N_24783);
nor UO_1499 (O_1499,N_24935,N_24983);
and UO_1500 (O_1500,N_24976,N_24920);
xnor UO_1501 (O_1501,N_24869,N_24829);
xor UO_1502 (O_1502,N_24917,N_24774);
xor UO_1503 (O_1503,N_24988,N_24871);
xor UO_1504 (O_1504,N_24948,N_24779);
or UO_1505 (O_1505,N_24841,N_24797);
and UO_1506 (O_1506,N_24966,N_24802);
and UO_1507 (O_1507,N_24959,N_24942);
nor UO_1508 (O_1508,N_24997,N_24911);
and UO_1509 (O_1509,N_24802,N_24912);
nand UO_1510 (O_1510,N_24766,N_24822);
nand UO_1511 (O_1511,N_24800,N_24993);
or UO_1512 (O_1512,N_24771,N_24914);
xor UO_1513 (O_1513,N_24868,N_24994);
nor UO_1514 (O_1514,N_24767,N_24990);
nor UO_1515 (O_1515,N_24851,N_24934);
nor UO_1516 (O_1516,N_24788,N_24972);
nor UO_1517 (O_1517,N_24809,N_24810);
xnor UO_1518 (O_1518,N_24812,N_24945);
and UO_1519 (O_1519,N_24937,N_24883);
and UO_1520 (O_1520,N_24860,N_24957);
and UO_1521 (O_1521,N_24944,N_24996);
or UO_1522 (O_1522,N_24948,N_24879);
or UO_1523 (O_1523,N_24927,N_24851);
nand UO_1524 (O_1524,N_24961,N_24978);
xnor UO_1525 (O_1525,N_24975,N_24986);
xor UO_1526 (O_1526,N_24819,N_24808);
nand UO_1527 (O_1527,N_24809,N_24795);
nor UO_1528 (O_1528,N_24986,N_24881);
or UO_1529 (O_1529,N_24918,N_24850);
nor UO_1530 (O_1530,N_24899,N_24831);
or UO_1531 (O_1531,N_24952,N_24928);
and UO_1532 (O_1532,N_24801,N_24868);
nor UO_1533 (O_1533,N_24901,N_24874);
and UO_1534 (O_1534,N_24831,N_24941);
nand UO_1535 (O_1535,N_24854,N_24772);
or UO_1536 (O_1536,N_24863,N_24935);
nand UO_1537 (O_1537,N_24964,N_24991);
xnor UO_1538 (O_1538,N_24966,N_24987);
nand UO_1539 (O_1539,N_24963,N_24794);
and UO_1540 (O_1540,N_24851,N_24898);
or UO_1541 (O_1541,N_24839,N_24918);
nor UO_1542 (O_1542,N_24917,N_24935);
nor UO_1543 (O_1543,N_24968,N_24829);
nor UO_1544 (O_1544,N_24980,N_24759);
or UO_1545 (O_1545,N_24875,N_24984);
nand UO_1546 (O_1546,N_24813,N_24873);
or UO_1547 (O_1547,N_24875,N_24905);
nand UO_1548 (O_1548,N_24904,N_24819);
nand UO_1549 (O_1549,N_24988,N_24855);
nor UO_1550 (O_1550,N_24830,N_24945);
nor UO_1551 (O_1551,N_24857,N_24789);
xnor UO_1552 (O_1552,N_24854,N_24985);
nor UO_1553 (O_1553,N_24979,N_24756);
xor UO_1554 (O_1554,N_24882,N_24942);
and UO_1555 (O_1555,N_24804,N_24816);
nor UO_1556 (O_1556,N_24957,N_24830);
or UO_1557 (O_1557,N_24955,N_24901);
and UO_1558 (O_1558,N_24872,N_24751);
nor UO_1559 (O_1559,N_24970,N_24942);
nor UO_1560 (O_1560,N_24901,N_24854);
or UO_1561 (O_1561,N_24750,N_24879);
nor UO_1562 (O_1562,N_24999,N_24849);
nor UO_1563 (O_1563,N_24812,N_24984);
nand UO_1564 (O_1564,N_24970,N_24802);
xnor UO_1565 (O_1565,N_24916,N_24843);
and UO_1566 (O_1566,N_24774,N_24846);
nor UO_1567 (O_1567,N_24851,N_24857);
xnor UO_1568 (O_1568,N_24819,N_24821);
xnor UO_1569 (O_1569,N_24889,N_24759);
nand UO_1570 (O_1570,N_24868,N_24902);
nand UO_1571 (O_1571,N_24852,N_24822);
nand UO_1572 (O_1572,N_24790,N_24913);
and UO_1573 (O_1573,N_24827,N_24903);
nand UO_1574 (O_1574,N_24776,N_24968);
and UO_1575 (O_1575,N_24849,N_24786);
xnor UO_1576 (O_1576,N_24943,N_24773);
and UO_1577 (O_1577,N_24802,N_24794);
nor UO_1578 (O_1578,N_24901,N_24763);
xnor UO_1579 (O_1579,N_24853,N_24973);
and UO_1580 (O_1580,N_24835,N_24862);
and UO_1581 (O_1581,N_24802,N_24771);
or UO_1582 (O_1582,N_24852,N_24767);
and UO_1583 (O_1583,N_24863,N_24977);
xnor UO_1584 (O_1584,N_24753,N_24918);
nand UO_1585 (O_1585,N_24939,N_24835);
nor UO_1586 (O_1586,N_24896,N_24780);
xor UO_1587 (O_1587,N_24916,N_24920);
or UO_1588 (O_1588,N_24949,N_24990);
nand UO_1589 (O_1589,N_24825,N_24953);
nor UO_1590 (O_1590,N_24972,N_24897);
nand UO_1591 (O_1591,N_24849,N_24809);
and UO_1592 (O_1592,N_24848,N_24919);
nor UO_1593 (O_1593,N_24912,N_24924);
xor UO_1594 (O_1594,N_24847,N_24878);
nand UO_1595 (O_1595,N_24753,N_24752);
or UO_1596 (O_1596,N_24819,N_24988);
nor UO_1597 (O_1597,N_24877,N_24893);
nor UO_1598 (O_1598,N_24987,N_24910);
and UO_1599 (O_1599,N_24778,N_24796);
or UO_1600 (O_1600,N_24785,N_24988);
or UO_1601 (O_1601,N_24806,N_24983);
or UO_1602 (O_1602,N_24790,N_24763);
and UO_1603 (O_1603,N_24978,N_24970);
nor UO_1604 (O_1604,N_24930,N_24754);
and UO_1605 (O_1605,N_24807,N_24920);
and UO_1606 (O_1606,N_24965,N_24888);
xnor UO_1607 (O_1607,N_24764,N_24787);
nor UO_1608 (O_1608,N_24814,N_24788);
xnor UO_1609 (O_1609,N_24994,N_24927);
and UO_1610 (O_1610,N_24943,N_24914);
nor UO_1611 (O_1611,N_24972,N_24826);
or UO_1612 (O_1612,N_24841,N_24755);
or UO_1613 (O_1613,N_24778,N_24860);
xor UO_1614 (O_1614,N_24785,N_24954);
xor UO_1615 (O_1615,N_24946,N_24886);
nor UO_1616 (O_1616,N_24967,N_24976);
or UO_1617 (O_1617,N_24788,N_24808);
nor UO_1618 (O_1618,N_24991,N_24949);
nor UO_1619 (O_1619,N_24950,N_24882);
nand UO_1620 (O_1620,N_24786,N_24893);
or UO_1621 (O_1621,N_24943,N_24837);
xnor UO_1622 (O_1622,N_24996,N_24885);
or UO_1623 (O_1623,N_24889,N_24761);
xor UO_1624 (O_1624,N_24807,N_24929);
xnor UO_1625 (O_1625,N_24975,N_24875);
or UO_1626 (O_1626,N_24834,N_24930);
nor UO_1627 (O_1627,N_24770,N_24862);
nand UO_1628 (O_1628,N_24829,N_24812);
xnor UO_1629 (O_1629,N_24771,N_24980);
nor UO_1630 (O_1630,N_24778,N_24837);
and UO_1631 (O_1631,N_24842,N_24802);
xnor UO_1632 (O_1632,N_24937,N_24854);
and UO_1633 (O_1633,N_24888,N_24966);
and UO_1634 (O_1634,N_24764,N_24772);
nand UO_1635 (O_1635,N_24927,N_24950);
and UO_1636 (O_1636,N_24877,N_24759);
nand UO_1637 (O_1637,N_24890,N_24764);
nor UO_1638 (O_1638,N_24786,N_24882);
or UO_1639 (O_1639,N_24773,N_24891);
and UO_1640 (O_1640,N_24920,N_24793);
xnor UO_1641 (O_1641,N_24983,N_24888);
and UO_1642 (O_1642,N_24780,N_24997);
xnor UO_1643 (O_1643,N_24910,N_24777);
xnor UO_1644 (O_1644,N_24789,N_24798);
or UO_1645 (O_1645,N_24958,N_24924);
xnor UO_1646 (O_1646,N_24940,N_24752);
nand UO_1647 (O_1647,N_24874,N_24906);
or UO_1648 (O_1648,N_24778,N_24849);
xor UO_1649 (O_1649,N_24986,N_24933);
and UO_1650 (O_1650,N_24842,N_24968);
xor UO_1651 (O_1651,N_24986,N_24822);
nor UO_1652 (O_1652,N_24837,N_24922);
nor UO_1653 (O_1653,N_24769,N_24765);
xor UO_1654 (O_1654,N_24792,N_24973);
and UO_1655 (O_1655,N_24914,N_24865);
xnor UO_1656 (O_1656,N_24800,N_24750);
or UO_1657 (O_1657,N_24982,N_24978);
nor UO_1658 (O_1658,N_24786,N_24851);
nand UO_1659 (O_1659,N_24989,N_24762);
or UO_1660 (O_1660,N_24961,N_24949);
nor UO_1661 (O_1661,N_24782,N_24989);
xnor UO_1662 (O_1662,N_24839,N_24760);
nand UO_1663 (O_1663,N_24887,N_24926);
or UO_1664 (O_1664,N_24863,N_24872);
and UO_1665 (O_1665,N_24764,N_24780);
nand UO_1666 (O_1666,N_24853,N_24843);
or UO_1667 (O_1667,N_24950,N_24783);
or UO_1668 (O_1668,N_24977,N_24838);
nand UO_1669 (O_1669,N_24870,N_24867);
xor UO_1670 (O_1670,N_24769,N_24760);
nand UO_1671 (O_1671,N_24799,N_24754);
or UO_1672 (O_1672,N_24923,N_24797);
nor UO_1673 (O_1673,N_24860,N_24962);
or UO_1674 (O_1674,N_24870,N_24830);
nand UO_1675 (O_1675,N_24838,N_24966);
xor UO_1676 (O_1676,N_24839,N_24750);
nor UO_1677 (O_1677,N_24962,N_24855);
nor UO_1678 (O_1678,N_24898,N_24883);
nand UO_1679 (O_1679,N_24750,N_24799);
and UO_1680 (O_1680,N_24912,N_24812);
and UO_1681 (O_1681,N_24769,N_24830);
xor UO_1682 (O_1682,N_24925,N_24985);
nand UO_1683 (O_1683,N_24986,N_24927);
nand UO_1684 (O_1684,N_24981,N_24961);
and UO_1685 (O_1685,N_24814,N_24922);
xnor UO_1686 (O_1686,N_24903,N_24964);
nand UO_1687 (O_1687,N_24778,N_24812);
xor UO_1688 (O_1688,N_24861,N_24847);
or UO_1689 (O_1689,N_24762,N_24874);
or UO_1690 (O_1690,N_24894,N_24984);
or UO_1691 (O_1691,N_24792,N_24989);
nand UO_1692 (O_1692,N_24966,N_24754);
and UO_1693 (O_1693,N_24905,N_24814);
or UO_1694 (O_1694,N_24818,N_24892);
and UO_1695 (O_1695,N_24863,N_24911);
xor UO_1696 (O_1696,N_24985,N_24769);
or UO_1697 (O_1697,N_24891,N_24817);
or UO_1698 (O_1698,N_24883,N_24925);
or UO_1699 (O_1699,N_24938,N_24874);
nand UO_1700 (O_1700,N_24884,N_24966);
nor UO_1701 (O_1701,N_24940,N_24905);
and UO_1702 (O_1702,N_24924,N_24997);
xnor UO_1703 (O_1703,N_24908,N_24947);
or UO_1704 (O_1704,N_24946,N_24834);
xor UO_1705 (O_1705,N_24975,N_24859);
or UO_1706 (O_1706,N_24990,N_24791);
or UO_1707 (O_1707,N_24965,N_24922);
nor UO_1708 (O_1708,N_24812,N_24952);
and UO_1709 (O_1709,N_24835,N_24920);
nor UO_1710 (O_1710,N_24975,N_24805);
xor UO_1711 (O_1711,N_24839,N_24864);
nand UO_1712 (O_1712,N_24872,N_24939);
nand UO_1713 (O_1713,N_24890,N_24906);
or UO_1714 (O_1714,N_24942,N_24923);
nand UO_1715 (O_1715,N_24829,N_24842);
nand UO_1716 (O_1716,N_24872,N_24958);
nand UO_1717 (O_1717,N_24813,N_24811);
nor UO_1718 (O_1718,N_24985,N_24773);
xor UO_1719 (O_1719,N_24955,N_24798);
nand UO_1720 (O_1720,N_24993,N_24798);
xor UO_1721 (O_1721,N_24852,N_24758);
xnor UO_1722 (O_1722,N_24897,N_24834);
nor UO_1723 (O_1723,N_24914,N_24901);
nor UO_1724 (O_1724,N_24900,N_24764);
and UO_1725 (O_1725,N_24977,N_24928);
nand UO_1726 (O_1726,N_24855,N_24795);
nor UO_1727 (O_1727,N_24844,N_24764);
nor UO_1728 (O_1728,N_24954,N_24773);
xor UO_1729 (O_1729,N_24764,N_24919);
and UO_1730 (O_1730,N_24858,N_24755);
nand UO_1731 (O_1731,N_24754,N_24817);
or UO_1732 (O_1732,N_24869,N_24805);
xnor UO_1733 (O_1733,N_24943,N_24839);
or UO_1734 (O_1734,N_24903,N_24828);
xnor UO_1735 (O_1735,N_24953,N_24808);
nor UO_1736 (O_1736,N_24809,N_24998);
nand UO_1737 (O_1737,N_24961,N_24777);
nand UO_1738 (O_1738,N_24789,N_24859);
nand UO_1739 (O_1739,N_24904,N_24757);
nand UO_1740 (O_1740,N_24952,N_24959);
xnor UO_1741 (O_1741,N_24951,N_24974);
and UO_1742 (O_1742,N_24833,N_24852);
nor UO_1743 (O_1743,N_24764,N_24980);
xor UO_1744 (O_1744,N_24866,N_24911);
xor UO_1745 (O_1745,N_24944,N_24869);
and UO_1746 (O_1746,N_24786,N_24821);
nor UO_1747 (O_1747,N_24912,N_24848);
xnor UO_1748 (O_1748,N_24752,N_24765);
or UO_1749 (O_1749,N_24953,N_24869);
nor UO_1750 (O_1750,N_24847,N_24819);
or UO_1751 (O_1751,N_24869,N_24877);
and UO_1752 (O_1752,N_24859,N_24782);
or UO_1753 (O_1753,N_24915,N_24773);
nor UO_1754 (O_1754,N_24820,N_24817);
nor UO_1755 (O_1755,N_24992,N_24935);
and UO_1756 (O_1756,N_24886,N_24807);
or UO_1757 (O_1757,N_24851,N_24921);
and UO_1758 (O_1758,N_24916,N_24790);
xnor UO_1759 (O_1759,N_24823,N_24750);
xnor UO_1760 (O_1760,N_24820,N_24859);
and UO_1761 (O_1761,N_24798,N_24914);
xor UO_1762 (O_1762,N_24948,N_24868);
nor UO_1763 (O_1763,N_24786,N_24890);
xnor UO_1764 (O_1764,N_24777,N_24821);
xor UO_1765 (O_1765,N_24889,N_24830);
and UO_1766 (O_1766,N_24803,N_24858);
or UO_1767 (O_1767,N_24780,N_24885);
or UO_1768 (O_1768,N_24793,N_24851);
or UO_1769 (O_1769,N_24954,N_24839);
or UO_1770 (O_1770,N_24913,N_24985);
or UO_1771 (O_1771,N_24927,N_24914);
xnor UO_1772 (O_1772,N_24812,N_24904);
nor UO_1773 (O_1773,N_24869,N_24991);
nor UO_1774 (O_1774,N_24948,N_24881);
nor UO_1775 (O_1775,N_24863,N_24778);
xor UO_1776 (O_1776,N_24911,N_24850);
and UO_1777 (O_1777,N_24855,N_24954);
nor UO_1778 (O_1778,N_24850,N_24962);
and UO_1779 (O_1779,N_24878,N_24953);
or UO_1780 (O_1780,N_24930,N_24951);
nor UO_1781 (O_1781,N_24965,N_24905);
and UO_1782 (O_1782,N_24959,N_24911);
or UO_1783 (O_1783,N_24832,N_24974);
or UO_1784 (O_1784,N_24985,N_24971);
or UO_1785 (O_1785,N_24888,N_24787);
xor UO_1786 (O_1786,N_24837,N_24781);
and UO_1787 (O_1787,N_24897,N_24874);
nor UO_1788 (O_1788,N_24992,N_24888);
nand UO_1789 (O_1789,N_24918,N_24826);
nand UO_1790 (O_1790,N_24800,N_24997);
and UO_1791 (O_1791,N_24981,N_24993);
nor UO_1792 (O_1792,N_24860,N_24902);
or UO_1793 (O_1793,N_24940,N_24790);
xor UO_1794 (O_1794,N_24831,N_24939);
nand UO_1795 (O_1795,N_24756,N_24821);
or UO_1796 (O_1796,N_24962,N_24904);
or UO_1797 (O_1797,N_24757,N_24896);
or UO_1798 (O_1798,N_24808,N_24774);
and UO_1799 (O_1799,N_24836,N_24756);
xnor UO_1800 (O_1800,N_24864,N_24879);
xnor UO_1801 (O_1801,N_24871,N_24915);
xnor UO_1802 (O_1802,N_24755,N_24762);
nor UO_1803 (O_1803,N_24886,N_24797);
and UO_1804 (O_1804,N_24876,N_24804);
or UO_1805 (O_1805,N_24808,N_24861);
xor UO_1806 (O_1806,N_24906,N_24828);
and UO_1807 (O_1807,N_24925,N_24831);
and UO_1808 (O_1808,N_24776,N_24822);
or UO_1809 (O_1809,N_24943,N_24810);
nand UO_1810 (O_1810,N_24983,N_24752);
nand UO_1811 (O_1811,N_24788,N_24755);
xor UO_1812 (O_1812,N_24865,N_24767);
nor UO_1813 (O_1813,N_24843,N_24808);
or UO_1814 (O_1814,N_24853,N_24929);
or UO_1815 (O_1815,N_24851,N_24936);
xor UO_1816 (O_1816,N_24965,N_24779);
nand UO_1817 (O_1817,N_24958,N_24860);
or UO_1818 (O_1818,N_24975,N_24756);
and UO_1819 (O_1819,N_24766,N_24805);
or UO_1820 (O_1820,N_24859,N_24834);
nand UO_1821 (O_1821,N_24966,N_24980);
xnor UO_1822 (O_1822,N_24825,N_24758);
and UO_1823 (O_1823,N_24821,N_24800);
nand UO_1824 (O_1824,N_24932,N_24783);
and UO_1825 (O_1825,N_24983,N_24780);
nand UO_1826 (O_1826,N_24857,N_24903);
xnor UO_1827 (O_1827,N_24759,N_24804);
xor UO_1828 (O_1828,N_24939,N_24914);
and UO_1829 (O_1829,N_24927,N_24971);
nor UO_1830 (O_1830,N_24883,N_24831);
nand UO_1831 (O_1831,N_24896,N_24918);
and UO_1832 (O_1832,N_24752,N_24873);
nand UO_1833 (O_1833,N_24838,N_24769);
nor UO_1834 (O_1834,N_24906,N_24799);
and UO_1835 (O_1835,N_24907,N_24991);
nor UO_1836 (O_1836,N_24838,N_24940);
nand UO_1837 (O_1837,N_24925,N_24956);
nor UO_1838 (O_1838,N_24765,N_24925);
xnor UO_1839 (O_1839,N_24815,N_24842);
or UO_1840 (O_1840,N_24994,N_24983);
nand UO_1841 (O_1841,N_24959,N_24854);
or UO_1842 (O_1842,N_24777,N_24886);
nand UO_1843 (O_1843,N_24984,N_24835);
or UO_1844 (O_1844,N_24988,N_24902);
and UO_1845 (O_1845,N_24850,N_24791);
and UO_1846 (O_1846,N_24809,N_24949);
or UO_1847 (O_1847,N_24930,N_24880);
and UO_1848 (O_1848,N_24869,N_24766);
nor UO_1849 (O_1849,N_24883,N_24842);
nor UO_1850 (O_1850,N_24837,N_24760);
and UO_1851 (O_1851,N_24819,N_24843);
nor UO_1852 (O_1852,N_24816,N_24963);
and UO_1853 (O_1853,N_24891,N_24968);
nand UO_1854 (O_1854,N_24966,N_24918);
xor UO_1855 (O_1855,N_24909,N_24769);
xor UO_1856 (O_1856,N_24994,N_24796);
nand UO_1857 (O_1857,N_24953,N_24783);
nand UO_1858 (O_1858,N_24887,N_24759);
nand UO_1859 (O_1859,N_24941,N_24921);
or UO_1860 (O_1860,N_24808,N_24892);
or UO_1861 (O_1861,N_24852,N_24970);
xor UO_1862 (O_1862,N_24962,N_24782);
nand UO_1863 (O_1863,N_24889,N_24928);
nand UO_1864 (O_1864,N_24801,N_24856);
and UO_1865 (O_1865,N_24916,N_24898);
xor UO_1866 (O_1866,N_24998,N_24931);
and UO_1867 (O_1867,N_24885,N_24880);
and UO_1868 (O_1868,N_24844,N_24942);
xor UO_1869 (O_1869,N_24921,N_24809);
nor UO_1870 (O_1870,N_24791,N_24981);
xor UO_1871 (O_1871,N_24892,N_24875);
xnor UO_1872 (O_1872,N_24786,N_24857);
nand UO_1873 (O_1873,N_24838,N_24927);
nand UO_1874 (O_1874,N_24922,N_24787);
nor UO_1875 (O_1875,N_24973,N_24971);
nand UO_1876 (O_1876,N_24899,N_24996);
nor UO_1877 (O_1877,N_24823,N_24959);
and UO_1878 (O_1878,N_24953,N_24909);
nand UO_1879 (O_1879,N_24904,N_24922);
nand UO_1880 (O_1880,N_24890,N_24839);
or UO_1881 (O_1881,N_24786,N_24956);
xor UO_1882 (O_1882,N_24976,N_24769);
nand UO_1883 (O_1883,N_24795,N_24820);
xnor UO_1884 (O_1884,N_24766,N_24910);
or UO_1885 (O_1885,N_24953,N_24856);
or UO_1886 (O_1886,N_24851,N_24874);
and UO_1887 (O_1887,N_24971,N_24782);
nor UO_1888 (O_1888,N_24844,N_24839);
or UO_1889 (O_1889,N_24958,N_24942);
nand UO_1890 (O_1890,N_24754,N_24870);
nor UO_1891 (O_1891,N_24891,N_24827);
and UO_1892 (O_1892,N_24877,N_24756);
and UO_1893 (O_1893,N_24982,N_24896);
or UO_1894 (O_1894,N_24785,N_24849);
xor UO_1895 (O_1895,N_24893,N_24757);
nor UO_1896 (O_1896,N_24940,N_24859);
xor UO_1897 (O_1897,N_24831,N_24902);
xor UO_1898 (O_1898,N_24897,N_24942);
xor UO_1899 (O_1899,N_24901,N_24934);
nand UO_1900 (O_1900,N_24901,N_24834);
or UO_1901 (O_1901,N_24773,N_24976);
and UO_1902 (O_1902,N_24860,N_24923);
xor UO_1903 (O_1903,N_24947,N_24964);
xor UO_1904 (O_1904,N_24971,N_24816);
nor UO_1905 (O_1905,N_24951,N_24798);
nor UO_1906 (O_1906,N_24879,N_24869);
and UO_1907 (O_1907,N_24843,N_24841);
nor UO_1908 (O_1908,N_24902,N_24877);
xnor UO_1909 (O_1909,N_24770,N_24780);
nand UO_1910 (O_1910,N_24862,N_24910);
and UO_1911 (O_1911,N_24945,N_24791);
xnor UO_1912 (O_1912,N_24872,N_24789);
or UO_1913 (O_1913,N_24767,N_24834);
or UO_1914 (O_1914,N_24770,N_24860);
and UO_1915 (O_1915,N_24950,N_24880);
or UO_1916 (O_1916,N_24838,N_24951);
and UO_1917 (O_1917,N_24803,N_24790);
xnor UO_1918 (O_1918,N_24764,N_24939);
xnor UO_1919 (O_1919,N_24885,N_24835);
or UO_1920 (O_1920,N_24761,N_24815);
and UO_1921 (O_1921,N_24751,N_24784);
and UO_1922 (O_1922,N_24970,N_24885);
and UO_1923 (O_1923,N_24938,N_24949);
xor UO_1924 (O_1924,N_24946,N_24952);
or UO_1925 (O_1925,N_24949,N_24930);
and UO_1926 (O_1926,N_24980,N_24889);
nor UO_1927 (O_1927,N_24990,N_24781);
and UO_1928 (O_1928,N_24822,N_24892);
or UO_1929 (O_1929,N_24925,N_24915);
xnor UO_1930 (O_1930,N_24960,N_24940);
nor UO_1931 (O_1931,N_24923,N_24754);
nand UO_1932 (O_1932,N_24856,N_24977);
or UO_1933 (O_1933,N_24993,N_24874);
xnor UO_1934 (O_1934,N_24885,N_24932);
nor UO_1935 (O_1935,N_24761,N_24882);
nand UO_1936 (O_1936,N_24810,N_24967);
nor UO_1937 (O_1937,N_24868,N_24864);
nor UO_1938 (O_1938,N_24895,N_24793);
nor UO_1939 (O_1939,N_24832,N_24757);
and UO_1940 (O_1940,N_24999,N_24970);
nor UO_1941 (O_1941,N_24848,N_24791);
nor UO_1942 (O_1942,N_24788,N_24907);
xnor UO_1943 (O_1943,N_24752,N_24934);
and UO_1944 (O_1944,N_24828,N_24822);
xnor UO_1945 (O_1945,N_24928,N_24873);
nand UO_1946 (O_1946,N_24981,N_24995);
nand UO_1947 (O_1947,N_24891,N_24809);
and UO_1948 (O_1948,N_24949,N_24833);
xor UO_1949 (O_1949,N_24927,N_24846);
nand UO_1950 (O_1950,N_24781,N_24806);
and UO_1951 (O_1951,N_24817,N_24841);
xor UO_1952 (O_1952,N_24808,N_24915);
and UO_1953 (O_1953,N_24843,N_24922);
nor UO_1954 (O_1954,N_24822,N_24936);
and UO_1955 (O_1955,N_24949,N_24911);
or UO_1956 (O_1956,N_24753,N_24751);
xnor UO_1957 (O_1957,N_24781,N_24959);
xnor UO_1958 (O_1958,N_24933,N_24915);
nor UO_1959 (O_1959,N_24804,N_24880);
nand UO_1960 (O_1960,N_24845,N_24868);
nand UO_1961 (O_1961,N_24816,N_24917);
xor UO_1962 (O_1962,N_24832,N_24869);
xnor UO_1963 (O_1963,N_24828,N_24859);
nand UO_1964 (O_1964,N_24872,N_24786);
xnor UO_1965 (O_1965,N_24763,N_24912);
or UO_1966 (O_1966,N_24943,N_24877);
or UO_1967 (O_1967,N_24977,N_24911);
nor UO_1968 (O_1968,N_24821,N_24758);
xor UO_1969 (O_1969,N_24801,N_24807);
nand UO_1970 (O_1970,N_24817,N_24792);
xnor UO_1971 (O_1971,N_24845,N_24876);
or UO_1972 (O_1972,N_24757,N_24842);
and UO_1973 (O_1973,N_24811,N_24812);
xnor UO_1974 (O_1974,N_24825,N_24812);
xnor UO_1975 (O_1975,N_24788,N_24835);
and UO_1976 (O_1976,N_24877,N_24923);
xnor UO_1977 (O_1977,N_24952,N_24755);
xor UO_1978 (O_1978,N_24829,N_24971);
and UO_1979 (O_1979,N_24970,N_24770);
nand UO_1980 (O_1980,N_24979,N_24776);
xor UO_1981 (O_1981,N_24783,N_24921);
xor UO_1982 (O_1982,N_24872,N_24963);
nor UO_1983 (O_1983,N_24873,N_24966);
nand UO_1984 (O_1984,N_24867,N_24791);
nand UO_1985 (O_1985,N_24919,N_24857);
or UO_1986 (O_1986,N_24887,N_24815);
nor UO_1987 (O_1987,N_24931,N_24863);
and UO_1988 (O_1988,N_24931,N_24877);
nand UO_1989 (O_1989,N_24845,N_24961);
xnor UO_1990 (O_1990,N_24896,N_24770);
or UO_1991 (O_1991,N_24947,N_24903);
and UO_1992 (O_1992,N_24913,N_24973);
or UO_1993 (O_1993,N_24804,N_24766);
nor UO_1994 (O_1994,N_24754,N_24795);
nor UO_1995 (O_1995,N_24997,N_24899);
xnor UO_1996 (O_1996,N_24941,N_24870);
nand UO_1997 (O_1997,N_24927,N_24755);
xor UO_1998 (O_1998,N_24976,N_24799);
nor UO_1999 (O_1999,N_24942,N_24909);
xor UO_2000 (O_2000,N_24955,N_24806);
nand UO_2001 (O_2001,N_24810,N_24905);
and UO_2002 (O_2002,N_24801,N_24996);
and UO_2003 (O_2003,N_24980,N_24818);
nor UO_2004 (O_2004,N_24902,N_24949);
xnor UO_2005 (O_2005,N_24845,N_24840);
xor UO_2006 (O_2006,N_24865,N_24785);
or UO_2007 (O_2007,N_24870,N_24979);
nand UO_2008 (O_2008,N_24763,N_24871);
nand UO_2009 (O_2009,N_24846,N_24897);
and UO_2010 (O_2010,N_24794,N_24843);
nand UO_2011 (O_2011,N_24948,N_24820);
and UO_2012 (O_2012,N_24814,N_24888);
or UO_2013 (O_2013,N_24989,N_24942);
xor UO_2014 (O_2014,N_24868,N_24940);
xnor UO_2015 (O_2015,N_24756,N_24835);
nor UO_2016 (O_2016,N_24899,N_24946);
nand UO_2017 (O_2017,N_24941,N_24890);
and UO_2018 (O_2018,N_24817,N_24921);
or UO_2019 (O_2019,N_24798,N_24763);
nand UO_2020 (O_2020,N_24771,N_24776);
or UO_2021 (O_2021,N_24822,N_24792);
nand UO_2022 (O_2022,N_24782,N_24834);
or UO_2023 (O_2023,N_24971,N_24822);
xor UO_2024 (O_2024,N_24981,N_24970);
nor UO_2025 (O_2025,N_24952,N_24911);
nor UO_2026 (O_2026,N_24896,N_24791);
nand UO_2027 (O_2027,N_24800,N_24850);
xnor UO_2028 (O_2028,N_24813,N_24808);
and UO_2029 (O_2029,N_24830,N_24944);
xor UO_2030 (O_2030,N_24928,N_24927);
xnor UO_2031 (O_2031,N_24816,N_24883);
or UO_2032 (O_2032,N_24836,N_24750);
xor UO_2033 (O_2033,N_24830,N_24923);
xnor UO_2034 (O_2034,N_24973,N_24860);
xor UO_2035 (O_2035,N_24919,N_24810);
nor UO_2036 (O_2036,N_24969,N_24913);
or UO_2037 (O_2037,N_24772,N_24832);
xnor UO_2038 (O_2038,N_24904,N_24817);
xor UO_2039 (O_2039,N_24814,N_24934);
nand UO_2040 (O_2040,N_24911,N_24773);
and UO_2041 (O_2041,N_24890,N_24900);
xnor UO_2042 (O_2042,N_24923,N_24960);
nand UO_2043 (O_2043,N_24781,N_24918);
and UO_2044 (O_2044,N_24858,N_24910);
nand UO_2045 (O_2045,N_24766,N_24811);
xor UO_2046 (O_2046,N_24917,N_24753);
nor UO_2047 (O_2047,N_24763,N_24981);
nor UO_2048 (O_2048,N_24927,N_24894);
xnor UO_2049 (O_2049,N_24754,N_24794);
xnor UO_2050 (O_2050,N_24805,N_24800);
nand UO_2051 (O_2051,N_24754,N_24952);
or UO_2052 (O_2052,N_24833,N_24821);
nand UO_2053 (O_2053,N_24810,N_24858);
xor UO_2054 (O_2054,N_24788,N_24771);
nand UO_2055 (O_2055,N_24893,N_24981);
nor UO_2056 (O_2056,N_24785,N_24772);
xor UO_2057 (O_2057,N_24901,N_24806);
nor UO_2058 (O_2058,N_24844,N_24905);
nor UO_2059 (O_2059,N_24764,N_24806);
nand UO_2060 (O_2060,N_24805,N_24900);
nand UO_2061 (O_2061,N_24885,N_24846);
and UO_2062 (O_2062,N_24909,N_24937);
or UO_2063 (O_2063,N_24794,N_24779);
and UO_2064 (O_2064,N_24762,N_24921);
nor UO_2065 (O_2065,N_24950,N_24851);
nand UO_2066 (O_2066,N_24811,N_24891);
or UO_2067 (O_2067,N_24802,N_24950);
nand UO_2068 (O_2068,N_24829,N_24820);
nand UO_2069 (O_2069,N_24789,N_24914);
nor UO_2070 (O_2070,N_24920,N_24751);
or UO_2071 (O_2071,N_24896,N_24955);
and UO_2072 (O_2072,N_24918,N_24933);
or UO_2073 (O_2073,N_24849,N_24994);
and UO_2074 (O_2074,N_24779,N_24913);
nand UO_2075 (O_2075,N_24905,N_24901);
nor UO_2076 (O_2076,N_24877,N_24758);
or UO_2077 (O_2077,N_24991,N_24998);
or UO_2078 (O_2078,N_24958,N_24980);
and UO_2079 (O_2079,N_24832,N_24946);
or UO_2080 (O_2080,N_24873,N_24780);
and UO_2081 (O_2081,N_24932,N_24774);
and UO_2082 (O_2082,N_24824,N_24863);
nor UO_2083 (O_2083,N_24921,N_24996);
or UO_2084 (O_2084,N_24928,N_24993);
and UO_2085 (O_2085,N_24825,N_24928);
xnor UO_2086 (O_2086,N_24966,N_24983);
nor UO_2087 (O_2087,N_24906,N_24889);
nand UO_2088 (O_2088,N_24792,N_24772);
and UO_2089 (O_2089,N_24823,N_24853);
xnor UO_2090 (O_2090,N_24779,N_24819);
or UO_2091 (O_2091,N_24918,N_24931);
nand UO_2092 (O_2092,N_24918,N_24824);
nand UO_2093 (O_2093,N_24872,N_24829);
or UO_2094 (O_2094,N_24928,N_24858);
and UO_2095 (O_2095,N_24764,N_24942);
and UO_2096 (O_2096,N_24901,N_24800);
or UO_2097 (O_2097,N_24755,N_24834);
xnor UO_2098 (O_2098,N_24820,N_24759);
or UO_2099 (O_2099,N_24943,N_24937);
nor UO_2100 (O_2100,N_24770,N_24949);
and UO_2101 (O_2101,N_24774,N_24814);
and UO_2102 (O_2102,N_24953,N_24990);
or UO_2103 (O_2103,N_24831,N_24768);
nor UO_2104 (O_2104,N_24751,N_24809);
and UO_2105 (O_2105,N_24849,N_24890);
or UO_2106 (O_2106,N_24944,N_24885);
nor UO_2107 (O_2107,N_24856,N_24944);
nor UO_2108 (O_2108,N_24754,N_24825);
nor UO_2109 (O_2109,N_24766,N_24908);
nor UO_2110 (O_2110,N_24799,N_24775);
xor UO_2111 (O_2111,N_24854,N_24821);
or UO_2112 (O_2112,N_24932,N_24895);
or UO_2113 (O_2113,N_24994,N_24791);
xor UO_2114 (O_2114,N_24928,N_24826);
xnor UO_2115 (O_2115,N_24822,N_24865);
nor UO_2116 (O_2116,N_24961,N_24875);
nor UO_2117 (O_2117,N_24931,N_24845);
nor UO_2118 (O_2118,N_24792,N_24908);
and UO_2119 (O_2119,N_24863,N_24805);
xnor UO_2120 (O_2120,N_24900,N_24864);
nand UO_2121 (O_2121,N_24991,N_24997);
nor UO_2122 (O_2122,N_24973,N_24832);
and UO_2123 (O_2123,N_24979,N_24900);
and UO_2124 (O_2124,N_24810,N_24861);
xnor UO_2125 (O_2125,N_24768,N_24853);
and UO_2126 (O_2126,N_24962,N_24869);
xor UO_2127 (O_2127,N_24840,N_24750);
nor UO_2128 (O_2128,N_24786,N_24923);
nand UO_2129 (O_2129,N_24997,N_24897);
nor UO_2130 (O_2130,N_24894,N_24844);
and UO_2131 (O_2131,N_24818,N_24814);
xnor UO_2132 (O_2132,N_24792,N_24949);
nor UO_2133 (O_2133,N_24821,N_24961);
and UO_2134 (O_2134,N_24934,N_24899);
xnor UO_2135 (O_2135,N_24841,N_24811);
xor UO_2136 (O_2136,N_24887,N_24770);
and UO_2137 (O_2137,N_24780,N_24895);
and UO_2138 (O_2138,N_24946,N_24955);
xor UO_2139 (O_2139,N_24836,N_24925);
nand UO_2140 (O_2140,N_24919,N_24788);
and UO_2141 (O_2141,N_24827,N_24965);
or UO_2142 (O_2142,N_24798,N_24779);
and UO_2143 (O_2143,N_24797,N_24991);
and UO_2144 (O_2144,N_24902,N_24751);
and UO_2145 (O_2145,N_24853,N_24827);
or UO_2146 (O_2146,N_24793,N_24912);
and UO_2147 (O_2147,N_24918,N_24861);
xor UO_2148 (O_2148,N_24852,N_24962);
or UO_2149 (O_2149,N_24884,N_24789);
and UO_2150 (O_2150,N_24877,N_24881);
or UO_2151 (O_2151,N_24832,N_24846);
nand UO_2152 (O_2152,N_24850,N_24853);
nand UO_2153 (O_2153,N_24861,N_24892);
and UO_2154 (O_2154,N_24846,N_24996);
xor UO_2155 (O_2155,N_24819,N_24865);
nor UO_2156 (O_2156,N_24779,N_24878);
or UO_2157 (O_2157,N_24788,N_24938);
nor UO_2158 (O_2158,N_24905,N_24890);
nor UO_2159 (O_2159,N_24757,N_24805);
nand UO_2160 (O_2160,N_24934,N_24970);
and UO_2161 (O_2161,N_24775,N_24836);
nor UO_2162 (O_2162,N_24865,N_24880);
and UO_2163 (O_2163,N_24767,N_24859);
nand UO_2164 (O_2164,N_24990,N_24809);
xor UO_2165 (O_2165,N_24902,N_24806);
nor UO_2166 (O_2166,N_24787,N_24751);
nand UO_2167 (O_2167,N_24947,N_24981);
nor UO_2168 (O_2168,N_24846,N_24977);
or UO_2169 (O_2169,N_24854,N_24943);
nand UO_2170 (O_2170,N_24983,N_24934);
and UO_2171 (O_2171,N_24949,N_24973);
or UO_2172 (O_2172,N_24928,N_24792);
nor UO_2173 (O_2173,N_24908,N_24905);
nand UO_2174 (O_2174,N_24902,N_24830);
and UO_2175 (O_2175,N_24978,N_24869);
nor UO_2176 (O_2176,N_24948,N_24834);
nand UO_2177 (O_2177,N_24789,N_24951);
and UO_2178 (O_2178,N_24855,N_24888);
and UO_2179 (O_2179,N_24830,N_24962);
nand UO_2180 (O_2180,N_24948,N_24941);
and UO_2181 (O_2181,N_24954,N_24860);
nor UO_2182 (O_2182,N_24753,N_24865);
or UO_2183 (O_2183,N_24983,N_24981);
or UO_2184 (O_2184,N_24985,N_24977);
xnor UO_2185 (O_2185,N_24998,N_24954);
nand UO_2186 (O_2186,N_24976,N_24947);
and UO_2187 (O_2187,N_24868,N_24943);
or UO_2188 (O_2188,N_24914,N_24984);
xor UO_2189 (O_2189,N_24980,N_24847);
and UO_2190 (O_2190,N_24944,N_24834);
nand UO_2191 (O_2191,N_24922,N_24830);
xor UO_2192 (O_2192,N_24967,N_24796);
nor UO_2193 (O_2193,N_24823,N_24953);
and UO_2194 (O_2194,N_24863,N_24806);
nand UO_2195 (O_2195,N_24770,N_24844);
and UO_2196 (O_2196,N_24908,N_24940);
xor UO_2197 (O_2197,N_24993,N_24990);
nor UO_2198 (O_2198,N_24881,N_24807);
and UO_2199 (O_2199,N_24831,N_24851);
nand UO_2200 (O_2200,N_24886,N_24855);
nor UO_2201 (O_2201,N_24851,N_24778);
and UO_2202 (O_2202,N_24997,N_24837);
nand UO_2203 (O_2203,N_24927,N_24884);
nand UO_2204 (O_2204,N_24963,N_24817);
and UO_2205 (O_2205,N_24881,N_24794);
and UO_2206 (O_2206,N_24753,N_24866);
and UO_2207 (O_2207,N_24919,N_24813);
nand UO_2208 (O_2208,N_24964,N_24898);
or UO_2209 (O_2209,N_24980,N_24970);
or UO_2210 (O_2210,N_24869,N_24811);
or UO_2211 (O_2211,N_24787,N_24781);
nand UO_2212 (O_2212,N_24840,N_24811);
xor UO_2213 (O_2213,N_24991,N_24810);
and UO_2214 (O_2214,N_24905,N_24752);
and UO_2215 (O_2215,N_24850,N_24899);
nor UO_2216 (O_2216,N_24943,N_24788);
nand UO_2217 (O_2217,N_24761,N_24953);
or UO_2218 (O_2218,N_24779,N_24755);
or UO_2219 (O_2219,N_24891,N_24930);
or UO_2220 (O_2220,N_24979,N_24953);
and UO_2221 (O_2221,N_24822,N_24891);
nand UO_2222 (O_2222,N_24899,N_24867);
or UO_2223 (O_2223,N_24892,N_24959);
xnor UO_2224 (O_2224,N_24803,N_24775);
nor UO_2225 (O_2225,N_24963,N_24852);
nand UO_2226 (O_2226,N_24962,N_24936);
or UO_2227 (O_2227,N_24996,N_24780);
nand UO_2228 (O_2228,N_24792,N_24861);
xnor UO_2229 (O_2229,N_24849,N_24755);
nand UO_2230 (O_2230,N_24940,N_24834);
nor UO_2231 (O_2231,N_24841,N_24764);
or UO_2232 (O_2232,N_24992,N_24838);
xor UO_2233 (O_2233,N_24860,N_24874);
nor UO_2234 (O_2234,N_24884,N_24914);
nand UO_2235 (O_2235,N_24761,N_24865);
nand UO_2236 (O_2236,N_24939,N_24770);
nand UO_2237 (O_2237,N_24962,N_24968);
or UO_2238 (O_2238,N_24821,N_24784);
nand UO_2239 (O_2239,N_24878,N_24880);
and UO_2240 (O_2240,N_24985,N_24795);
and UO_2241 (O_2241,N_24984,N_24969);
nand UO_2242 (O_2242,N_24862,N_24771);
nand UO_2243 (O_2243,N_24917,N_24807);
nor UO_2244 (O_2244,N_24927,N_24766);
xor UO_2245 (O_2245,N_24811,N_24949);
nor UO_2246 (O_2246,N_24773,N_24896);
nor UO_2247 (O_2247,N_24995,N_24937);
nand UO_2248 (O_2248,N_24905,N_24882);
xnor UO_2249 (O_2249,N_24815,N_24865);
and UO_2250 (O_2250,N_24814,N_24930);
nor UO_2251 (O_2251,N_24801,N_24900);
nor UO_2252 (O_2252,N_24989,N_24997);
xnor UO_2253 (O_2253,N_24911,N_24897);
nand UO_2254 (O_2254,N_24848,N_24758);
nand UO_2255 (O_2255,N_24788,N_24899);
and UO_2256 (O_2256,N_24769,N_24876);
and UO_2257 (O_2257,N_24947,N_24843);
or UO_2258 (O_2258,N_24796,N_24866);
nand UO_2259 (O_2259,N_24825,N_24950);
nand UO_2260 (O_2260,N_24842,N_24921);
xnor UO_2261 (O_2261,N_24781,N_24938);
and UO_2262 (O_2262,N_24753,N_24771);
nor UO_2263 (O_2263,N_24990,N_24939);
nor UO_2264 (O_2264,N_24750,N_24761);
nor UO_2265 (O_2265,N_24993,N_24776);
or UO_2266 (O_2266,N_24991,N_24978);
nand UO_2267 (O_2267,N_24848,N_24940);
nand UO_2268 (O_2268,N_24938,N_24751);
or UO_2269 (O_2269,N_24937,N_24778);
xnor UO_2270 (O_2270,N_24763,N_24775);
and UO_2271 (O_2271,N_24910,N_24849);
or UO_2272 (O_2272,N_24843,N_24882);
and UO_2273 (O_2273,N_24786,N_24816);
and UO_2274 (O_2274,N_24786,N_24848);
nand UO_2275 (O_2275,N_24911,N_24752);
nand UO_2276 (O_2276,N_24936,N_24989);
xor UO_2277 (O_2277,N_24794,N_24903);
nand UO_2278 (O_2278,N_24794,N_24950);
nor UO_2279 (O_2279,N_24991,N_24782);
nand UO_2280 (O_2280,N_24791,N_24998);
nor UO_2281 (O_2281,N_24933,N_24810);
nand UO_2282 (O_2282,N_24822,N_24925);
and UO_2283 (O_2283,N_24938,N_24835);
or UO_2284 (O_2284,N_24812,N_24916);
or UO_2285 (O_2285,N_24765,N_24863);
nor UO_2286 (O_2286,N_24787,N_24880);
xnor UO_2287 (O_2287,N_24990,N_24856);
xor UO_2288 (O_2288,N_24922,N_24944);
nor UO_2289 (O_2289,N_24892,N_24799);
and UO_2290 (O_2290,N_24973,N_24985);
nor UO_2291 (O_2291,N_24911,N_24799);
and UO_2292 (O_2292,N_24944,N_24793);
nand UO_2293 (O_2293,N_24993,N_24795);
nand UO_2294 (O_2294,N_24805,N_24980);
nor UO_2295 (O_2295,N_24880,N_24834);
or UO_2296 (O_2296,N_24942,N_24901);
or UO_2297 (O_2297,N_24924,N_24751);
nor UO_2298 (O_2298,N_24937,N_24863);
nand UO_2299 (O_2299,N_24849,N_24919);
and UO_2300 (O_2300,N_24961,N_24817);
xnor UO_2301 (O_2301,N_24991,N_24856);
xor UO_2302 (O_2302,N_24970,N_24861);
xnor UO_2303 (O_2303,N_24956,N_24937);
or UO_2304 (O_2304,N_24753,N_24813);
and UO_2305 (O_2305,N_24869,N_24808);
nor UO_2306 (O_2306,N_24872,N_24952);
nor UO_2307 (O_2307,N_24882,N_24906);
and UO_2308 (O_2308,N_24821,N_24764);
xor UO_2309 (O_2309,N_24889,N_24892);
nor UO_2310 (O_2310,N_24778,N_24910);
nand UO_2311 (O_2311,N_24974,N_24924);
xnor UO_2312 (O_2312,N_24957,N_24961);
nand UO_2313 (O_2313,N_24780,N_24806);
or UO_2314 (O_2314,N_24925,N_24766);
or UO_2315 (O_2315,N_24818,N_24991);
nand UO_2316 (O_2316,N_24893,N_24835);
nor UO_2317 (O_2317,N_24862,N_24874);
xnor UO_2318 (O_2318,N_24955,N_24846);
and UO_2319 (O_2319,N_24903,N_24868);
and UO_2320 (O_2320,N_24919,N_24829);
nor UO_2321 (O_2321,N_24881,N_24957);
or UO_2322 (O_2322,N_24872,N_24964);
and UO_2323 (O_2323,N_24864,N_24824);
nand UO_2324 (O_2324,N_24818,N_24793);
nand UO_2325 (O_2325,N_24941,N_24966);
xor UO_2326 (O_2326,N_24863,N_24852);
or UO_2327 (O_2327,N_24920,N_24790);
nand UO_2328 (O_2328,N_24935,N_24889);
xor UO_2329 (O_2329,N_24979,N_24961);
and UO_2330 (O_2330,N_24968,N_24881);
or UO_2331 (O_2331,N_24891,N_24973);
nand UO_2332 (O_2332,N_24839,N_24870);
xor UO_2333 (O_2333,N_24817,N_24804);
xor UO_2334 (O_2334,N_24830,N_24815);
nor UO_2335 (O_2335,N_24997,N_24956);
or UO_2336 (O_2336,N_24955,N_24781);
nor UO_2337 (O_2337,N_24901,N_24927);
or UO_2338 (O_2338,N_24863,N_24869);
and UO_2339 (O_2339,N_24807,N_24981);
xnor UO_2340 (O_2340,N_24939,N_24874);
and UO_2341 (O_2341,N_24859,N_24788);
nor UO_2342 (O_2342,N_24924,N_24934);
xor UO_2343 (O_2343,N_24927,N_24771);
or UO_2344 (O_2344,N_24785,N_24780);
nor UO_2345 (O_2345,N_24780,N_24781);
and UO_2346 (O_2346,N_24958,N_24807);
or UO_2347 (O_2347,N_24840,N_24782);
or UO_2348 (O_2348,N_24775,N_24814);
or UO_2349 (O_2349,N_24832,N_24861);
or UO_2350 (O_2350,N_24913,N_24916);
xnor UO_2351 (O_2351,N_24876,N_24778);
and UO_2352 (O_2352,N_24794,N_24860);
and UO_2353 (O_2353,N_24971,N_24890);
nor UO_2354 (O_2354,N_24769,N_24882);
nand UO_2355 (O_2355,N_24793,N_24760);
xnor UO_2356 (O_2356,N_24997,N_24925);
nor UO_2357 (O_2357,N_24856,N_24874);
nand UO_2358 (O_2358,N_24885,N_24989);
or UO_2359 (O_2359,N_24932,N_24965);
xnor UO_2360 (O_2360,N_24845,N_24871);
nand UO_2361 (O_2361,N_24845,N_24979);
and UO_2362 (O_2362,N_24762,N_24915);
and UO_2363 (O_2363,N_24984,N_24754);
nor UO_2364 (O_2364,N_24875,N_24901);
nand UO_2365 (O_2365,N_24858,N_24885);
and UO_2366 (O_2366,N_24799,N_24794);
or UO_2367 (O_2367,N_24958,N_24756);
nand UO_2368 (O_2368,N_24971,N_24914);
nor UO_2369 (O_2369,N_24874,N_24919);
and UO_2370 (O_2370,N_24914,N_24782);
nor UO_2371 (O_2371,N_24788,N_24998);
nand UO_2372 (O_2372,N_24909,N_24751);
xor UO_2373 (O_2373,N_24768,N_24988);
nor UO_2374 (O_2374,N_24911,N_24760);
nor UO_2375 (O_2375,N_24996,N_24811);
or UO_2376 (O_2376,N_24889,N_24900);
xor UO_2377 (O_2377,N_24988,N_24847);
nor UO_2378 (O_2378,N_24975,N_24940);
nor UO_2379 (O_2379,N_24968,N_24880);
nor UO_2380 (O_2380,N_24763,N_24961);
or UO_2381 (O_2381,N_24931,N_24916);
nor UO_2382 (O_2382,N_24751,N_24911);
xor UO_2383 (O_2383,N_24881,N_24892);
and UO_2384 (O_2384,N_24881,N_24828);
nor UO_2385 (O_2385,N_24815,N_24771);
nor UO_2386 (O_2386,N_24929,N_24848);
xnor UO_2387 (O_2387,N_24957,N_24999);
nor UO_2388 (O_2388,N_24801,N_24995);
or UO_2389 (O_2389,N_24779,N_24957);
and UO_2390 (O_2390,N_24894,N_24967);
or UO_2391 (O_2391,N_24877,N_24884);
nand UO_2392 (O_2392,N_24753,N_24804);
and UO_2393 (O_2393,N_24872,N_24846);
and UO_2394 (O_2394,N_24900,N_24921);
xor UO_2395 (O_2395,N_24949,N_24979);
nand UO_2396 (O_2396,N_24931,N_24973);
or UO_2397 (O_2397,N_24861,N_24978);
nand UO_2398 (O_2398,N_24909,N_24961);
or UO_2399 (O_2399,N_24752,N_24871);
xnor UO_2400 (O_2400,N_24794,N_24921);
nor UO_2401 (O_2401,N_24917,N_24865);
nor UO_2402 (O_2402,N_24809,N_24978);
or UO_2403 (O_2403,N_24881,N_24753);
and UO_2404 (O_2404,N_24787,N_24792);
xor UO_2405 (O_2405,N_24900,N_24809);
nand UO_2406 (O_2406,N_24791,N_24801);
xor UO_2407 (O_2407,N_24853,N_24863);
xnor UO_2408 (O_2408,N_24995,N_24986);
nand UO_2409 (O_2409,N_24908,N_24872);
or UO_2410 (O_2410,N_24852,N_24870);
xnor UO_2411 (O_2411,N_24899,N_24799);
nor UO_2412 (O_2412,N_24861,N_24981);
and UO_2413 (O_2413,N_24859,N_24863);
nor UO_2414 (O_2414,N_24942,N_24780);
or UO_2415 (O_2415,N_24981,N_24862);
and UO_2416 (O_2416,N_24836,N_24931);
nor UO_2417 (O_2417,N_24996,N_24842);
and UO_2418 (O_2418,N_24852,N_24948);
nor UO_2419 (O_2419,N_24798,N_24959);
nand UO_2420 (O_2420,N_24956,N_24999);
or UO_2421 (O_2421,N_24958,N_24812);
or UO_2422 (O_2422,N_24956,N_24932);
xor UO_2423 (O_2423,N_24862,N_24788);
nand UO_2424 (O_2424,N_24890,N_24776);
and UO_2425 (O_2425,N_24811,N_24938);
xor UO_2426 (O_2426,N_24969,N_24949);
nor UO_2427 (O_2427,N_24897,N_24814);
and UO_2428 (O_2428,N_24917,N_24989);
nand UO_2429 (O_2429,N_24897,N_24824);
xor UO_2430 (O_2430,N_24928,N_24912);
and UO_2431 (O_2431,N_24805,N_24939);
or UO_2432 (O_2432,N_24798,N_24962);
nand UO_2433 (O_2433,N_24995,N_24898);
or UO_2434 (O_2434,N_24818,N_24848);
nor UO_2435 (O_2435,N_24957,N_24910);
xnor UO_2436 (O_2436,N_24927,N_24963);
or UO_2437 (O_2437,N_24835,N_24797);
nor UO_2438 (O_2438,N_24803,N_24863);
xnor UO_2439 (O_2439,N_24818,N_24950);
or UO_2440 (O_2440,N_24878,N_24886);
nor UO_2441 (O_2441,N_24852,N_24845);
nand UO_2442 (O_2442,N_24868,N_24817);
or UO_2443 (O_2443,N_24993,N_24907);
or UO_2444 (O_2444,N_24901,N_24845);
or UO_2445 (O_2445,N_24904,N_24823);
xnor UO_2446 (O_2446,N_24957,N_24938);
or UO_2447 (O_2447,N_24859,N_24943);
nor UO_2448 (O_2448,N_24960,N_24919);
nand UO_2449 (O_2449,N_24836,N_24940);
nand UO_2450 (O_2450,N_24957,N_24775);
and UO_2451 (O_2451,N_24769,N_24863);
nor UO_2452 (O_2452,N_24859,N_24897);
nand UO_2453 (O_2453,N_24914,N_24966);
xor UO_2454 (O_2454,N_24772,N_24800);
nand UO_2455 (O_2455,N_24753,N_24988);
nand UO_2456 (O_2456,N_24889,N_24931);
xnor UO_2457 (O_2457,N_24963,N_24920);
or UO_2458 (O_2458,N_24975,N_24931);
nor UO_2459 (O_2459,N_24764,N_24751);
and UO_2460 (O_2460,N_24936,N_24934);
or UO_2461 (O_2461,N_24766,N_24887);
nor UO_2462 (O_2462,N_24760,N_24761);
xor UO_2463 (O_2463,N_24909,N_24934);
xnor UO_2464 (O_2464,N_24960,N_24884);
or UO_2465 (O_2465,N_24841,N_24822);
and UO_2466 (O_2466,N_24768,N_24894);
or UO_2467 (O_2467,N_24897,N_24803);
and UO_2468 (O_2468,N_24837,N_24782);
nand UO_2469 (O_2469,N_24825,N_24926);
and UO_2470 (O_2470,N_24803,N_24960);
and UO_2471 (O_2471,N_24899,N_24895);
and UO_2472 (O_2472,N_24767,N_24866);
and UO_2473 (O_2473,N_24920,N_24758);
nand UO_2474 (O_2474,N_24989,N_24821);
nand UO_2475 (O_2475,N_24822,N_24795);
and UO_2476 (O_2476,N_24750,N_24900);
nand UO_2477 (O_2477,N_24828,N_24991);
xor UO_2478 (O_2478,N_24779,N_24916);
nand UO_2479 (O_2479,N_24847,N_24851);
nand UO_2480 (O_2480,N_24916,N_24963);
and UO_2481 (O_2481,N_24919,N_24896);
or UO_2482 (O_2482,N_24839,N_24848);
xor UO_2483 (O_2483,N_24994,N_24802);
nor UO_2484 (O_2484,N_24882,N_24801);
or UO_2485 (O_2485,N_24899,N_24793);
nor UO_2486 (O_2486,N_24920,N_24979);
nor UO_2487 (O_2487,N_24970,N_24818);
nor UO_2488 (O_2488,N_24951,N_24833);
nor UO_2489 (O_2489,N_24904,N_24873);
nand UO_2490 (O_2490,N_24868,N_24807);
and UO_2491 (O_2491,N_24992,N_24849);
nor UO_2492 (O_2492,N_24915,N_24935);
or UO_2493 (O_2493,N_24843,N_24958);
and UO_2494 (O_2494,N_24891,N_24892);
and UO_2495 (O_2495,N_24909,N_24907);
and UO_2496 (O_2496,N_24901,N_24804);
and UO_2497 (O_2497,N_24954,N_24899);
nor UO_2498 (O_2498,N_24953,N_24925);
nor UO_2499 (O_2499,N_24823,N_24800);
and UO_2500 (O_2500,N_24810,N_24843);
or UO_2501 (O_2501,N_24806,N_24845);
nor UO_2502 (O_2502,N_24968,N_24995);
nor UO_2503 (O_2503,N_24967,N_24763);
nor UO_2504 (O_2504,N_24830,N_24849);
xor UO_2505 (O_2505,N_24853,N_24826);
or UO_2506 (O_2506,N_24788,N_24877);
xnor UO_2507 (O_2507,N_24838,N_24785);
xnor UO_2508 (O_2508,N_24830,N_24897);
and UO_2509 (O_2509,N_24777,N_24774);
or UO_2510 (O_2510,N_24845,N_24820);
nor UO_2511 (O_2511,N_24860,N_24755);
or UO_2512 (O_2512,N_24885,N_24873);
nor UO_2513 (O_2513,N_24992,N_24822);
xnor UO_2514 (O_2514,N_24868,N_24928);
and UO_2515 (O_2515,N_24973,N_24941);
and UO_2516 (O_2516,N_24820,N_24781);
or UO_2517 (O_2517,N_24846,N_24795);
and UO_2518 (O_2518,N_24885,N_24905);
xnor UO_2519 (O_2519,N_24908,N_24758);
nor UO_2520 (O_2520,N_24990,N_24931);
nand UO_2521 (O_2521,N_24969,N_24935);
or UO_2522 (O_2522,N_24900,N_24837);
nor UO_2523 (O_2523,N_24957,N_24991);
and UO_2524 (O_2524,N_24937,N_24970);
nand UO_2525 (O_2525,N_24999,N_24930);
and UO_2526 (O_2526,N_24989,N_24847);
xor UO_2527 (O_2527,N_24918,N_24923);
or UO_2528 (O_2528,N_24987,N_24760);
and UO_2529 (O_2529,N_24859,N_24854);
nor UO_2530 (O_2530,N_24989,N_24972);
nand UO_2531 (O_2531,N_24801,N_24982);
and UO_2532 (O_2532,N_24854,N_24950);
or UO_2533 (O_2533,N_24963,N_24994);
xnor UO_2534 (O_2534,N_24867,N_24969);
xor UO_2535 (O_2535,N_24893,N_24779);
or UO_2536 (O_2536,N_24830,N_24852);
and UO_2537 (O_2537,N_24918,N_24965);
nor UO_2538 (O_2538,N_24774,N_24802);
or UO_2539 (O_2539,N_24967,N_24987);
nor UO_2540 (O_2540,N_24954,N_24791);
and UO_2541 (O_2541,N_24890,N_24889);
nand UO_2542 (O_2542,N_24769,N_24934);
nand UO_2543 (O_2543,N_24804,N_24964);
or UO_2544 (O_2544,N_24758,N_24911);
nor UO_2545 (O_2545,N_24989,N_24837);
nand UO_2546 (O_2546,N_24965,N_24816);
nand UO_2547 (O_2547,N_24785,N_24857);
nand UO_2548 (O_2548,N_24971,N_24852);
or UO_2549 (O_2549,N_24760,N_24974);
xnor UO_2550 (O_2550,N_24881,N_24778);
and UO_2551 (O_2551,N_24801,N_24904);
nor UO_2552 (O_2552,N_24902,N_24762);
nor UO_2553 (O_2553,N_24942,N_24846);
xor UO_2554 (O_2554,N_24768,N_24828);
and UO_2555 (O_2555,N_24774,N_24838);
nor UO_2556 (O_2556,N_24991,N_24969);
nor UO_2557 (O_2557,N_24999,N_24758);
nand UO_2558 (O_2558,N_24925,N_24963);
xor UO_2559 (O_2559,N_24865,N_24841);
or UO_2560 (O_2560,N_24956,N_24794);
and UO_2561 (O_2561,N_24952,N_24982);
xor UO_2562 (O_2562,N_24943,N_24774);
nand UO_2563 (O_2563,N_24987,N_24750);
and UO_2564 (O_2564,N_24770,N_24921);
nor UO_2565 (O_2565,N_24927,N_24813);
nand UO_2566 (O_2566,N_24855,N_24770);
nor UO_2567 (O_2567,N_24856,N_24774);
and UO_2568 (O_2568,N_24995,N_24750);
and UO_2569 (O_2569,N_24844,N_24911);
nand UO_2570 (O_2570,N_24806,N_24838);
nand UO_2571 (O_2571,N_24786,N_24808);
nand UO_2572 (O_2572,N_24946,N_24846);
nand UO_2573 (O_2573,N_24878,N_24763);
xnor UO_2574 (O_2574,N_24958,N_24889);
and UO_2575 (O_2575,N_24900,N_24912);
and UO_2576 (O_2576,N_24979,N_24779);
and UO_2577 (O_2577,N_24948,N_24837);
nand UO_2578 (O_2578,N_24867,N_24849);
xnor UO_2579 (O_2579,N_24787,N_24985);
or UO_2580 (O_2580,N_24830,N_24785);
nor UO_2581 (O_2581,N_24835,N_24759);
nand UO_2582 (O_2582,N_24985,N_24866);
nand UO_2583 (O_2583,N_24871,N_24893);
xor UO_2584 (O_2584,N_24914,N_24922);
or UO_2585 (O_2585,N_24877,N_24970);
nor UO_2586 (O_2586,N_24900,N_24924);
nor UO_2587 (O_2587,N_24845,N_24759);
or UO_2588 (O_2588,N_24756,N_24980);
and UO_2589 (O_2589,N_24787,N_24996);
or UO_2590 (O_2590,N_24970,N_24864);
xnor UO_2591 (O_2591,N_24770,N_24800);
and UO_2592 (O_2592,N_24919,N_24789);
nor UO_2593 (O_2593,N_24840,N_24923);
xnor UO_2594 (O_2594,N_24812,N_24764);
or UO_2595 (O_2595,N_24832,N_24939);
xor UO_2596 (O_2596,N_24996,N_24950);
nor UO_2597 (O_2597,N_24824,N_24971);
or UO_2598 (O_2598,N_24820,N_24848);
xor UO_2599 (O_2599,N_24751,N_24921);
nand UO_2600 (O_2600,N_24964,N_24763);
nor UO_2601 (O_2601,N_24905,N_24833);
and UO_2602 (O_2602,N_24968,N_24781);
nor UO_2603 (O_2603,N_24759,N_24843);
xor UO_2604 (O_2604,N_24907,N_24982);
nor UO_2605 (O_2605,N_24900,N_24852);
or UO_2606 (O_2606,N_24970,N_24961);
xor UO_2607 (O_2607,N_24943,N_24940);
xnor UO_2608 (O_2608,N_24994,N_24753);
or UO_2609 (O_2609,N_24860,N_24858);
and UO_2610 (O_2610,N_24916,N_24984);
xor UO_2611 (O_2611,N_24765,N_24879);
nand UO_2612 (O_2612,N_24943,N_24901);
xnor UO_2613 (O_2613,N_24976,N_24791);
nand UO_2614 (O_2614,N_24966,N_24948);
or UO_2615 (O_2615,N_24848,N_24941);
nand UO_2616 (O_2616,N_24961,N_24923);
nand UO_2617 (O_2617,N_24765,N_24970);
xor UO_2618 (O_2618,N_24803,N_24895);
xnor UO_2619 (O_2619,N_24976,N_24925);
nand UO_2620 (O_2620,N_24975,N_24851);
xnor UO_2621 (O_2621,N_24945,N_24993);
xor UO_2622 (O_2622,N_24907,N_24984);
xnor UO_2623 (O_2623,N_24958,N_24934);
nor UO_2624 (O_2624,N_24818,N_24891);
or UO_2625 (O_2625,N_24990,N_24786);
xor UO_2626 (O_2626,N_24886,N_24973);
nand UO_2627 (O_2627,N_24876,N_24777);
or UO_2628 (O_2628,N_24831,N_24818);
xor UO_2629 (O_2629,N_24936,N_24827);
nor UO_2630 (O_2630,N_24947,N_24837);
or UO_2631 (O_2631,N_24780,N_24817);
or UO_2632 (O_2632,N_24967,N_24866);
nor UO_2633 (O_2633,N_24977,N_24777);
xor UO_2634 (O_2634,N_24894,N_24883);
and UO_2635 (O_2635,N_24893,N_24906);
nand UO_2636 (O_2636,N_24898,N_24809);
or UO_2637 (O_2637,N_24980,N_24904);
nor UO_2638 (O_2638,N_24969,N_24871);
or UO_2639 (O_2639,N_24949,N_24767);
or UO_2640 (O_2640,N_24948,N_24995);
nor UO_2641 (O_2641,N_24911,N_24774);
nor UO_2642 (O_2642,N_24886,N_24919);
xor UO_2643 (O_2643,N_24859,N_24992);
nor UO_2644 (O_2644,N_24763,N_24955);
xnor UO_2645 (O_2645,N_24928,N_24769);
and UO_2646 (O_2646,N_24955,N_24885);
nand UO_2647 (O_2647,N_24938,N_24850);
or UO_2648 (O_2648,N_24922,N_24862);
nor UO_2649 (O_2649,N_24830,N_24842);
nand UO_2650 (O_2650,N_24868,N_24781);
nand UO_2651 (O_2651,N_24862,N_24925);
or UO_2652 (O_2652,N_24828,N_24808);
xor UO_2653 (O_2653,N_24769,N_24892);
nor UO_2654 (O_2654,N_24788,N_24999);
and UO_2655 (O_2655,N_24864,N_24876);
nand UO_2656 (O_2656,N_24766,N_24772);
nand UO_2657 (O_2657,N_24853,N_24883);
xnor UO_2658 (O_2658,N_24900,N_24836);
xnor UO_2659 (O_2659,N_24940,N_24776);
nor UO_2660 (O_2660,N_24875,N_24853);
and UO_2661 (O_2661,N_24912,N_24809);
nand UO_2662 (O_2662,N_24786,N_24797);
nand UO_2663 (O_2663,N_24884,N_24862);
and UO_2664 (O_2664,N_24982,N_24909);
nand UO_2665 (O_2665,N_24989,N_24766);
nand UO_2666 (O_2666,N_24809,N_24963);
or UO_2667 (O_2667,N_24810,N_24868);
xnor UO_2668 (O_2668,N_24787,N_24895);
nor UO_2669 (O_2669,N_24851,N_24974);
and UO_2670 (O_2670,N_24776,N_24954);
nand UO_2671 (O_2671,N_24763,N_24875);
nand UO_2672 (O_2672,N_24839,N_24937);
or UO_2673 (O_2673,N_24997,N_24850);
and UO_2674 (O_2674,N_24842,N_24941);
xor UO_2675 (O_2675,N_24848,N_24997);
xnor UO_2676 (O_2676,N_24992,N_24900);
and UO_2677 (O_2677,N_24773,N_24947);
or UO_2678 (O_2678,N_24872,N_24961);
xor UO_2679 (O_2679,N_24878,N_24981);
and UO_2680 (O_2680,N_24770,N_24768);
xnor UO_2681 (O_2681,N_24847,N_24820);
nor UO_2682 (O_2682,N_24874,N_24768);
nor UO_2683 (O_2683,N_24976,N_24804);
nand UO_2684 (O_2684,N_24927,N_24973);
nand UO_2685 (O_2685,N_24904,N_24919);
nand UO_2686 (O_2686,N_24903,N_24876);
or UO_2687 (O_2687,N_24858,N_24763);
xor UO_2688 (O_2688,N_24945,N_24759);
and UO_2689 (O_2689,N_24882,N_24758);
and UO_2690 (O_2690,N_24876,N_24794);
nand UO_2691 (O_2691,N_24861,N_24948);
nand UO_2692 (O_2692,N_24938,N_24997);
xor UO_2693 (O_2693,N_24925,N_24864);
nand UO_2694 (O_2694,N_24801,N_24768);
xnor UO_2695 (O_2695,N_24990,N_24776);
nand UO_2696 (O_2696,N_24760,N_24775);
xor UO_2697 (O_2697,N_24942,N_24933);
and UO_2698 (O_2698,N_24860,N_24828);
xor UO_2699 (O_2699,N_24929,N_24766);
and UO_2700 (O_2700,N_24939,N_24769);
or UO_2701 (O_2701,N_24916,N_24802);
xnor UO_2702 (O_2702,N_24784,N_24942);
nor UO_2703 (O_2703,N_24838,N_24948);
nor UO_2704 (O_2704,N_24781,N_24872);
or UO_2705 (O_2705,N_24888,N_24943);
nor UO_2706 (O_2706,N_24978,N_24942);
or UO_2707 (O_2707,N_24895,N_24783);
and UO_2708 (O_2708,N_24928,N_24771);
and UO_2709 (O_2709,N_24830,N_24915);
nand UO_2710 (O_2710,N_24789,N_24839);
nor UO_2711 (O_2711,N_24796,N_24995);
nand UO_2712 (O_2712,N_24953,N_24888);
and UO_2713 (O_2713,N_24781,N_24907);
xnor UO_2714 (O_2714,N_24809,N_24823);
and UO_2715 (O_2715,N_24836,N_24893);
nor UO_2716 (O_2716,N_24802,N_24918);
or UO_2717 (O_2717,N_24941,N_24853);
nand UO_2718 (O_2718,N_24917,N_24958);
xor UO_2719 (O_2719,N_24905,N_24774);
xor UO_2720 (O_2720,N_24819,N_24862);
nor UO_2721 (O_2721,N_24892,N_24845);
xor UO_2722 (O_2722,N_24817,N_24824);
xor UO_2723 (O_2723,N_24858,N_24863);
nor UO_2724 (O_2724,N_24811,N_24874);
nand UO_2725 (O_2725,N_24922,N_24984);
xnor UO_2726 (O_2726,N_24792,N_24828);
nor UO_2727 (O_2727,N_24920,N_24770);
xor UO_2728 (O_2728,N_24906,N_24921);
or UO_2729 (O_2729,N_24798,N_24790);
nand UO_2730 (O_2730,N_24765,N_24960);
and UO_2731 (O_2731,N_24995,N_24751);
xnor UO_2732 (O_2732,N_24891,N_24825);
and UO_2733 (O_2733,N_24822,N_24831);
and UO_2734 (O_2734,N_24884,N_24842);
nor UO_2735 (O_2735,N_24964,N_24943);
nor UO_2736 (O_2736,N_24788,N_24929);
nor UO_2737 (O_2737,N_24957,N_24965);
nor UO_2738 (O_2738,N_24989,N_24778);
and UO_2739 (O_2739,N_24826,N_24835);
and UO_2740 (O_2740,N_24913,N_24910);
nand UO_2741 (O_2741,N_24822,N_24758);
xnor UO_2742 (O_2742,N_24977,N_24801);
or UO_2743 (O_2743,N_24846,N_24777);
nor UO_2744 (O_2744,N_24859,N_24837);
or UO_2745 (O_2745,N_24825,N_24923);
or UO_2746 (O_2746,N_24910,N_24983);
nand UO_2747 (O_2747,N_24985,N_24897);
nand UO_2748 (O_2748,N_24838,N_24791);
or UO_2749 (O_2749,N_24874,N_24854);
or UO_2750 (O_2750,N_24968,N_24780);
and UO_2751 (O_2751,N_24956,N_24809);
xor UO_2752 (O_2752,N_24918,N_24913);
or UO_2753 (O_2753,N_24790,N_24923);
nand UO_2754 (O_2754,N_24807,N_24967);
and UO_2755 (O_2755,N_24890,N_24821);
nor UO_2756 (O_2756,N_24971,N_24851);
nor UO_2757 (O_2757,N_24982,N_24788);
xor UO_2758 (O_2758,N_24778,N_24803);
or UO_2759 (O_2759,N_24863,N_24871);
xnor UO_2760 (O_2760,N_24971,N_24905);
or UO_2761 (O_2761,N_24801,N_24934);
xnor UO_2762 (O_2762,N_24888,N_24782);
xor UO_2763 (O_2763,N_24867,N_24861);
xnor UO_2764 (O_2764,N_24986,N_24764);
or UO_2765 (O_2765,N_24921,N_24837);
xnor UO_2766 (O_2766,N_24937,N_24888);
nor UO_2767 (O_2767,N_24966,N_24816);
nand UO_2768 (O_2768,N_24777,N_24792);
nand UO_2769 (O_2769,N_24963,N_24873);
nand UO_2770 (O_2770,N_24832,N_24800);
nor UO_2771 (O_2771,N_24969,N_24972);
xnor UO_2772 (O_2772,N_24891,N_24783);
nor UO_2773 (O_2773,N_24810,N_24807);
nor UO_2774 (O_2774,N_24953,N_24947);
nand UO_2775 (O_2775,N_24836,N_24854);
and UO_2776 (O_2776,N_24759,N_24754);
nand UO_2777 (O_2777,N_24946,N_24991);
xor UO_2778 (O_2778,N_24824,N_24842);
nand UO_2779 (O_2779,N_24755,N_24928);
and UO_2780 (O_2780,N_24946,N_24777);
nor UO_2781 (O_2781,N_24895,N_24986);
or UO_2782 (O_2782,N_24835,N_24764);
or UO_2783 (O_2783,N_24763,N_24752);
or UO_2784 (O_2784,N_24904,N_24777);
nor UO_2785 (O_2785,N_24953,N_24751);
nand UO_2786 (O_2786,N_24821,N_24953);
and UO_2787 (O_2787,N_24949,N_24819);
nor UO_2788 (O_2788,N_24948,N_24947);
xnor UO_2789 (O_2789,N_24826,N_24901);
xor UO_2790 (O_2790,N_24860,N_24803);
nand UO_2791 (O_2791,N_24862,N_24841);
nor UO_2792 (O_2792,N_24841,N_24768);
and UO_2793 (O_2793,N_24827,N_24850);
or UO_2794 (O_2794,N_24774,N_24962);
xor UO_2795 (O_2795,N_24771,N_24993);
and UO_2796 (O_2796,N_24831,N_24796);
nor UO_2797 (O_2797,N_24799,N_24968);
and UO_2798 (O_2798,N_24864,N_24844);
nor UO_2799 (O_2799,N_24879,N_24967);
or UO_2800 (O_2800,N_24799,N_24795);
xnor UO_2801 (O_2801,N_24926,N_24938);
nand UO_2802 (O_2802,N_24785,N_24764);
or UO_2803 (O_2803,N_24911,N_24852);
nand UO_2804 (O_2804,N_24885,N_24925);
xor UO_2805 (O_2805,N_24876,N_24999);
and UO_2806 (O_2806,N_24991,N_24967);
xnor UO_2807 (O_2807,N_24896,N_24940);
or UO_2808 (O_2808,N_24838,N_24816);
xor UO_2809 (O_2809,N_24963,N_24788);
nor UO_2810 (O_2810,N_24769,N_24910);
or UO_2811 (O_2811,N_24761,N_24822);
and UO_2812 (O_2812,N_24766,N_24990);
nor UO_2813 (O_2813,N_24878,N_24821);
and UO_2814 (O_2814,N_24896,N_24806);
nor UO_2815 (O_2815,N_24861,N_24766);
xnor UO_2816 (O_2816,N_24912,N_24935);
nor UO_2817 (O_2817,N_24775,N_24884);
nand UO_2818 (O_2818,N_24824,N_24970);
and UO_2819 (O_2819,N_24980,N_24809);
xnor UO_2820 (O_2820,N_24892,N_24836);
and UO_2821 (O_2821,N_24940,N_24918);
or UO_2822 (O_2822,N_24871,N_24797);
xor UO_2823 (O_2823,N_24979,N_24786);
xnor UO_2824 (O_2824,N_24792,N_24938);
nand UO_2825 (O_2825,N_24859,N_24755);
and UO_2826 (O_2826,N_24820,N_24862);
and UO_2827 (O_2827,N_24972,N_24965);
nor UO_2828 (O_2828,N_24926,N_24853);
and UO_2829 (O_2829,N_24938,N_24765);
nand UO_2830 (O_2830,N_24857,N_24954);
and UO_2831 (O_2831,N_24856,N_24881);
and UO_2832 (O_2832,N_24920,N_24883);
nand UO_2833 (O_2833,N_24985,N_24918);
or UO_2834 (O_2834,N_24797,N_24790);
nor UO_2835 (O_2835,N_24841,N_24969);
nor UO_2836 (O_2836,N_24787,N_24774);
xnor UO_2837 (O_2837,N_24915,N_24851);
nand UO_2838 (O_2838,N_24779,N_24756);
nand UO_2839 (O_2839,N_24947,N_24782);
nand UO_2840 (O_2840,N_24897,N_24925);
or UO_2841 (O_2841,N_24940,N_24967);
nor UO_2842 (O_2842,N_24889,N_24895);
and UO_2843 (O_2843,N_24998,N_24888);
nand UO_2844 (O_2844,N_24834,N_24833);
or UO_2845 (O_2845,N_24934,N_24800);
nand UO_2846 (O_2846,N_24832,N_24954);
nand UO_2847 (O_2847,N_24865,N_24922);
xnor UO_2848 (O_2848,N_24781,N_24811);
nand UO_2849 (O_2849,N_24784,N_24794);
or UO_2850 (O_2850,N_24971,N_24751);
xor UO_2851 (O_2851,N_24868,N_24955);
nor UO_2852 (O_2852,N_24959,N_24962);
xor UO_2853 (O_2853,N_24963,N_24834);
nand UO_2854 (O_2854,N_24793,N_24932);
nand UO_2855 (O_2855,N_24804,N_24818);
xor UO_2856 (O_2856,N_24813,N_24918);
and UO_2857 (O_2857,N_24859,N_24973);
xnor UO_2858 (O_2858,N_24752,N_24907);
nor UO_2859 (O_2859,N_24836,N_24869);
nand UO_2860 (O_2860,N_24762,N_24849);
and UO_2861 (O_2861,N_24805,N_24873);
and UO_2862 (O_2862,N_24862,N_24765);
nor UO_2863 (O_2863,N_24907,N_24875);
nand UO_2864 (O_2864,N_24845,N_24872);
or UO_2865 (O_2865,N_24988,N_24767);
xnor UO_2866 (O_2866,N_24874,N_24915);
or UO_2867 (O_2867,N_24773,N_24917);
nand UO_2868 (O_2868,N_24894,N_24836);
nor UO_2869 (O_2869,N_24874,N_24824);
xnor UO_2870 (O_2870,N_24873,N_24890);
or UO_2871 (O_2871,N_24858,N_24841);
nor UO_2872 (O_2872,N_24794,N_24844);
xor UO_2873 (O_2873,N_24828,N_24827);
nor UO_2874 (O_2874,N_24858,N_24890);
nand UO_2875 (O_2875,N_24844,N_24866);
nand UO_2876 (O_2876,N_24864,N_24793);
nor UO_2877 (O_2877,N_24908,N_24765);
or UO_2878 (O_2878,N_24877,N_24832);
nor UO_2879 (O_2879,N_24836,N_24878);
or UO_2880 (O_2880,N_24897,N_24855);
nand UO_2881 (O_2881,N_24760,N_24984);
nor UO_2882 (O_2882,N_24975,N_24837);
or UO_2883 (O_2883,N_24767,N_24882);
xor UO_2884 (O_2884,N_24970,N_24827);
or UO_2885 (O_2885,N_24885,N_24945);
nand UO_2886 (O_2886,N_24898,N_24932);
xnor UO_2887 (O_2887,N_24769,N_24773);
and UO_2888 (O_2888,N_24788,N_24931);
or UO_2889 (O_2889,N_24853,N_24939);
and UO_2890 (O_2890,N_24794,N_24877);
nand UO_2891 (O_2891,N_24983,N_24817);
nand UO_2892 (O_2892,N_24809,N_24981);
and UO_2893 (O_2893,N_24827,N_24823);
xor UO_2894 (O_2894,N_24985,N_24988);
and UO_2895 (O_2895,N_24793,N_24978);
and UO_2896 (O_2896,N_24865,N_24783);
or UO_2897 (O_2897,N_24840,N_24971);
nor UO_2898 (O_2898,N_24835,N_24914);
or UO_2899 (O_2899,N_24996,N_24932);
nor UO_2900 (O_2900,N_24863,N_24877);
nand UO_2901 (O_2901,N_24938,N_24939);
nand UO_2902 (O_2902,N_24929,N_24780);
or UO_2903 (O_2903,N_24904,N_24884);
and UO_2904 (O_2904,N_24769,N_24971);
or UO_2905 (O_2905,N_24926,N_24976);
nor UO_2906 (O_2906,N_24822,N_24966);
and UO_2907 (O_2907,N_24759,N_24832);
nand UO_2908 (O_2908,N_24998,N_24946);
or UO_2909 (O_2909,N_24854,N_24804);
nor UO_2910 (O_2910,N_24943,N_24961);
nor UO_2911 (O_2911,N_24754,N_24881);
and UO_2912 (O_2912,N_24866,N_24905);
and UO_2913 (O_2913,N_24932,N_24815);
or UO_2914 (O_2914,N_24862,N_24991);
nor UO_2915 (O_2915,N_24897,N_24889);
nand UO_2916 (O_2916,N_24890,N_24822);
xor UO_2917 (O_2917,N_24841,N_24942);
or UO_2918 (O_2918,N_24962,N_24909);
and UO_2919 (O_2919,N_24925,N_24907);
xnor UO_2920 (O_2920,N_24992,N_24906);
nand UO_2921 (O_2921,N_24913,N_24810);
xnor UO_2922 (O_2922,N_24895,N_24766);
nand UO_2923 (O_2923,N_24918,N_24807);
and UO_2924 (O_2924,N_24954,N_24992);
and UO_2925 (O_2925,N_24877,N_24851);
nand UO_2926 (O_2926,N_24895,N_24896);
or UO_2927 (O_2927,N_24887,N_24916);
nand UO_2928 (O_2928,N_24877,N_24991);
nand UO_2929 (O_2929,N_24844,N_24841);
and UO_2930 (O_2930,N_24872,N_24800);
xor UO_2931 (O_2931,N_24914,N_24881);
xnor UO_2932 (O_2932,N_24909,N_24947);
nor UO_2933 (O_2933,N_24888,N_24854);
or UO_2934 (O_2934,N_24845,N_24942);
nor UO_2935 (O_2935,N_24884,N_24799);
or UO_2936 (O_2936,N_24794,N_24856);
and UO_2937 (O_2937,N_24839,N_24905);
nand UO_2938 (O_2938,N_24885,N_24892);
or UO_2939 (O_2939,N_24784,N_24899);
or UO_2940 (O_2940,N_24949,N_24827);
nand UO_2941 (O_2941,N_24956,N_24766);
or UO_2942 (O_2942,N_24994,N_24922);
and UO_2943 (O_2943,N_24955,N_24900);
or UO_2944 (O_2944,N_24894,N_24777);
or UO_2945 (O_2945,N_24907,N_24975);
nor UO_2946 (O_2946,N_24899,N_24751);
and UO_2947 (O_2947,N_24864,N_24782);
xnor UO_2948 (O_2948,N_24797,N_24830);
or UO_2949 (O_2949,N_24949,N_24972);
nor UO_2950 (O_2950,N_24963,N_24921);
nor UO_2951 (O_2951,N_24925,N_24929);
and UO_2952 (O_2952,N_24772,N_24858);
or UO_2953 (O_2953,N_24887,N_24856);
and UO_2954 (O_2954,N_24945,N_24950);
or UO_2955 (O_2955,N_24949,N_24873);
nand UO_2956 (O_2956,N_24919,N_24937);
xnor UO_2957 (O_2957,N_24990,N_24977);
nor UO_2958 (O_2958,N_24803,N_24992);
nor UO_2959 (O_2959,N_24857,N_24750);
xor UO_2960 (O_2960,N_24843,N_24859);
nand UO_2961 (O_2961,N_24878,N_24952);
nor UO_2962 (O_2962,N_24923,N_24959);
nor UO_2963 (O_2963,N_24972,N_24775);
xnor UO_2964 (O_2964,N_24891,N_24931);
or UO_2965 (O_2965,N_24763,N_24918);
and UO_2966 (O_2966,N_24840,N_24862);
or UO_2967 (O_2967,N_24890,N_24855);
xnor UO_2968 (O_2968,N_24920,N_24971);
nand UO_2969 (O_2969,N_24797,N_24934);
nor UO_2970 (O_2970,N_24818,N_24976);
and UO_2971 (O_2971,N_24824,N_24996);
and UO_2972 (O_2972,N_24819,N_24927);
or UO_2973 (O_2973,N_24817,N_24932);
nor UO_2974 (O_2974,N_24933,N_24936);
xor UO_2975 (O_2975,N_24791,N_24790);
or UO_2976 (O_2976,N_24977,N_24803);
nand UO_2977 (O_2977,N_24752,N_24767);
and UO_2978 (O_2978,N_24765,N_24964);
xor UO_2979 (O_2979,N_24767,N_24789);
nor UO_2980 (O_2980,N_24797,N_24975);
xor UO_2981 (O_2981,N_24840,N_24927);
nor UO_2982 (O_2982,N_24781,N_24894);
nand UO_2983 (O_2983,N_24781,N_24870);
and UO_2984 (O_2984,N_24829,N_24757);
nand UO_2985 (O_2985,N_24858,N_24915);
and UO_2986 (O_2986,N_24765,N_24931);
and UO_2987 (O_2987,N_24901,N_24827);
xor UO_2988 (O_2988,N_24778,N_24903);
and UO_2989 (O_2989,N_24784,N_24852);
or UO_2990 (O_2990,N_24881,N_24895);
and UO_2991 (O_2991,N_24893,N_24827);
and UO_2992 (O_2992,N_24806,N_24771);
xnor UO_2993 (O_2993,N_24958,N_24950);
nand UO_2994 (O_2994,N_24833,N_24898);
and UO_2995 (O_2995,N_24922,N_24776);
and UO_2996 (O_2996,N_24913,N_24912);
nor UO_2997 (O_2997,N_24872,N_24893);
nand UO_2998 (O_2998,N_24967,N_24869);
xor UO_2999 (O_2999,N_24983,N_24948);
endmodule